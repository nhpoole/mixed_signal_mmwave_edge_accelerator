magic
tech sky130A
magscale 1 2
timestamp 1624494425
<< locali >>
rect 0 5639 2354 5673
rect 138 5369 1754 5403
rect 262 5121 1854 5155
rect 2165 4970 2199 5004
rect 0 4225 2354 4259
rect 2165 3480 2199 3514
rect 1374 3329 1854 3363
rect 1002 3081 1754 3115
rect 0 2811 2354 2845
rect 1250 2541 1754 2575
rect 1126 2293 1854 2327
rect 262 2142 594 2176
rect 2165 2142 2199 2176
rect 0 1397 2354 1431
rect 138 652 594 686
rect 2165 652 2199 686
rect 1126 501 1854 535
rect 1002 253 1754 287
rect 0 -17 2354 17
<< metal1 >>
rect 374 5630 438 5682
rect 1486 5630 1550 5682
rect 124 698 152 5532
rect 248 2188 276 5532
rect 374 4216 438 4268
rect 374 2802 438 2854
rect 239 2130 285 2188
rect 677 2133 741 2185
rect 115 640 161 698
rect 124 124 152 640
rect 248 124 276 2130
rect 374 1388 438 1440
rect 677 643 741 695
rect 988 124 1016 5532
rect 1112 124 1140 5532
rect 1236 124 1264 5532
rect 1360 124 1388 5532
rect 1486 4216 1550 4268
rect 1486 2802 1550 2854
rect 1486 1388 1550 1440
rect 374 -26 438 26
rect 1486 -26 1550 26
<< metal2 >>
rect 378 5632 434 5680
rect 1490 5632 1546 5680
rect 378 4218 434 4266
rect 1490 4218 1546 4266
rect 378 2804 434 2852
rect 1490 2804 1546 2852
rect 850 2730 1126 2758
rect 850 2173 878 2730
rect 709 2145 878 2173
rect 378 1390 434 1438
rect 1490 1390 1546 1438
rect 850 1316 1002 1344
rect 850 683 878 1316
rect 709 655 878 683
rect 378 -24 434 24
rect 1490 -24 1546 24
<< metal3 >>
rect 357 5607 455 5705
rect 1469 5607 1567 5705
rect 357 4193 455 4291
rect 1469 4193 1567 4291
rect 357 2779 455 2877
rect 1469 2779 1567 2877
rect 357 1365 455 1463
rect 1469 1365 1567 1463
rect 357 -49 455 49
rect 1469 -49 1567 49
use contact_16  contact_16_9
timestamp 1624494425
transform 1 0 105 0 1 640
box 0 0 66 58
use contact_9  contact_9_13
timestamp 1624494425
transform 1 0 373 0 1 -37
box 0 0 66 74
use contact_8  contact_8_13
timestamp 1624494425
transform 1 0 374 0 1 -32
box 0 0 64 64
use contact_7  contact_7_13
timestamp 1624494425
transform 1 0 377 0 1 -33
box 0 0 58 66
use contact_8  contact_8_17
timestamp 1624494425
transform 1 0 677 0 1 637
box 0 0 64 64
use contact_7  contact_7_21
timestamp 1624494425
transform 1 0 680 0 1 636
box 0 0 58 66
use contact_9  contact_9_11
timestamp 1624494425
transform 1 0 373 0 1 1377
box 0 0 66 74
use contact_8  contact_8_11
timestamp 1624494425
transform 1 0 374 0 1 1382
box 0 0 64 64
use contact_7  contact_7_11
timestamp 1624494425
transform 1 0 377 0 1 1381
box 0 0 58 66
use contact_9  contact_9_15
timestamp 1624494425
transform 1 0 373 0 1 1377
box 0 0 66 74
use contact_8  contact_8_15
timestamp 1624494425
transform 1 0 374 0 1 1382
box 0 0 64 64
use contact_7  contact_7_15
timestamp 1624494425
transform 1 0 377 0 1 1381
box 0 0 58 66
use pinv_1  pinv_1_1
timestamp 1624494425
transform 1 0 496 0 1 0
box -36 -17 404 1471
use pinv_1  pinv_1_0
timestamp 1624494425
transform 1 0 496 0 -1 2828
box -36 -17 404 1471
use contact_16  contact_16_7
timestamp 1624494425
transform 1 0 969 0 1 241
box 0 0 66 58
use contact_16  contact_16_6
timestamp 1624494425
transform 1 0 1093 0 1 489
box 0 0 66 58
use contact_9  contact_9_12
timestamp 1624494425
transform 1 0 1485 0 1 -37
box 0 0 66 74
use contact_8  contact_8_12
timestamp 1624494425
transform 1 0 1486 0 1 -32
box 0 0 64 64
use contact_7  contact_7_12
timestamp 1624494425
transform 1 0 1489 0 1 -33
box 0 0 58 66
use contact_17  contact_17_1
timestamp 1624494425
transform 1 0 970 0 1 1298
box 0 0 64 64
use contact_9  contact_9_10
timestamp 1624494425
transform 1 0 1485 0 1 1377
box 0 0 66 74
use contact_8  contact_8_10
timestamp 1624494425
transform 1 0 1486 0 1 1382
box 0 0 64 64
use contact_7  contact_7_10
timestamp 1624494425
transform 1 0 1489 0 1 1381
box 0 0 58 66
use contact_9  contact_9_14
timestamp 1624494425
transform 1 0 1485 0 1 1377
box 0 0 66 74
use contact_8  contact_8_14
timestamp 1624494425
transform 1 0 1486 0 1 1382
box 0 0 64 64
use contact_7  contact_7_14
timestamp 1624494425
transform 1 0 1489 0 1 1381
box 0 0 58 66
use pand2_0  pand2_0_3
timestamp 1624494425
transform 1 0 1608 0 1 0
box -36 -17 782 1471
use pand2_0  pand2_0_2
timestamp 1624494425
transform 1 0 1608 0 -1 2828
box -36 -17 782 1471
use contact_7  contact_7_20
timestamp 1624494425
transform 1 0 680 0 1 2126
box 0 0 58 66
use contact_8  contact_8_16
timestamp 1624494425
transform 1 0 677 0 1 2127
box 0 0 64 64
use contact_7  contact_7_9
timestamp 1624494425
transform 1 0 377 0 1 2795
box 0 0 58 66
use contact_8  contact_8_9
timestamp 1624494425
transform 1 0 374 0 1 2796
box 0 0 64 64
use contact_9  contact_9_9
timestamp 1624494425
transform 1 0 373 0 1 2791
box 0 0 66 74
use contact_7  contact_7_5
timestamp 1624494425
transform 1 0 377 0 1 2795
box 0 0 58 66
use contact_8  contact_8_5
timestamp 1624494425
transform 1 0 374 0 1 2796
box 0 0 64 64
use contact_9  contact_9_5
timestamp 1624494425
transform 1 0 373 0 1 2791
box 0 0 66 74
use contact_16  contact_16_8
timestamp 1624494425
transform 1 0 229 0 1 2130
box 0 0 66 58
use contact_17  contact_17_0
timestamp 1624494425
transform 1 0 1094 0 1 2712
box 0 0 64 64
use contact_16  contact_16_5
timestamp 1624494425
transform 1 0 1217 0 1 2529
box 0 0 66 58
use contact_16  contact_16_4
timestamp 1624494425
transform 1 0 1093 0 1 2281
box 0 0 66 58
use contact_9  contact_9_4
timestamp 1624494425
transform 1 0 1485 0 1 2791
box 0 0 66 74
use contact_8  contact_8_4
timestamp 1624494425
transform 1 0 1486 0 1 2796
box 0 0 64 64
use contact_7  contact_7_4
timestamp 1624494425
transform 1 0 1489 0 1 2795
box 0 0 58 66
use contact_9  contact_9_8
timestamp 1624494425
transform 1 0 1485 0 1 2791
box 0 0 66 74
use contact_8  contact_8_8
timestamp 1624494425
transform 1 0 1486 0 1 2796
box 0 0 64 64
use contact_7  contact_7_8
timestamp 1624494425
transform 1 0 1489 0 1 2795
box 0 0 58 66
use pand2_0  pand2_0_1
timestamp 1624494425
transform 1 0 1608 0 1 2828
box -36 -17 782 1471
use contact_7  contact_7_7
timestamp 1624494425
transform 1 0 377 0 1 4209
box 0 0 58 66
use contact_8  contact_8_7
timestamp 1624494425
transform 1 0 374 0 1 4210
box 0 0 64 64
use contact_9  contact_9_7
timestamp 1624494425
transform 1 0 373 0 1 4205
box 0 0 66 74
use contact_7  contact_7_3
timestamp 1624494425
transform 1 0 377 0 1 4209
box 0 0 58 66
use contact_8  contact_8_3
timestamp 1624494425
transform 1 0 374 0 1 4210
box 0 0 64 64
use contact_9  contact_9_3
timestamp 1624494425
transform 1 0 373 0 1 4205
box 0 0 66 74
use contact_7  contact_7_6
timestamp 1624494425
transform 1 0 1489 0 1 4209
box 0 0 58 66
use contact_8  contact_8_6
timestamp 1624494425
transform 1 0 1486 0 1 4210
box 0 0 64 64
use contact_9  contact_9_6
timestamp 1624494425
transform 1 0 1485 0 1 4205
box 0 0 66 74
use contact_7  contact_7_2
timestamp 1624494425
transform 1 0 1489 0 1 4209
box 0 0 58 66
use contact_8  contact_8_2
timestamp 1624494425
transform 1 0 1486 0 1 4210
box 0 0 64 64
use contact_9  contact_9_2
timestamp 1624494425
transform 1 0 1485 0 1 4205
box 0 0 66 74
use contact_16  contact_16_2
timestamp 1624494425
transform 1 0 1341 0 1 3317
box 0 0 66 58
use contact_16  contact_16_3
timestamp 1624494425
transform 1 0 969 0 1 3069
box 0 0 66 58
use pand2_0  pand2_0_0
timestamp 1624494425
transform 1 0 1608 0 -1 5656
box -36 -17 782 1471
use contact_7  contact_7_19
timestamp 1624494425
transform 1 0 109 0 1 5353
box 0 0 58 66
use contact_7  contact_7_17
timestamp 1624494425
transform 1 0 233 0 1 5105
box 0 0 58 66
use contact_7  contact_7_1
timestamp 1624494425
transform 1 0 377 0 1 5623
box 0 0 58 66
use contact_8  contact_8_1
timestamp 1624494425
transform 1 0 374 0 1 5624
box 0 0 64 64
use contact_9  contact_9_1
timestamp 1624494425
transform 1 0 373 0 1 5619
box 0 0 66 74
use contact_7  contact_7_18
timestamp 1624494425
transform 1 0 1221 0 1 5353
box 0 0 58 66
use contact_7  contact_7_16
timestamp 1624494425
transform 1 0 1345 0 1 5105
box 0 0 58 66
use contact_7  contact_7_0
timestamp 1624494425
transform 1 0 1489 0 1 5623
box 0 0 58 66
use contact_8  contact_8_0
timestamp 1624494425
transform 1 0 1486 0 1 5624
box 0 0 64 64
use contact_9  contact_9_0
timestamp 1624494425
transform 1 0 1485 0 1 5619
box 0 0 66 74
use contact_16  contact_16_0
timestamp 1624494425
transform 1 0 1341 0 1 5109
box 0 0 66 58
use contact_16  contact_16_1
timestamp 1624494425
transform 1 0 1217 0 1 5357
box 0 0 66 58
<< labels >>
rlabel metal1 s 115 640 161 698 4 in_0
rlabel metal1 s 239 2130 285 2188 4 in_1
rlabel locali s 2182 669 2182 669 4 out_0
rlabel locali s 2182 2159 2182 2159 4 out_1
rlabel locali s 2182 3497 2182 3497 4 out_2
rlabel locali s 2182 4987 2182 4987 4 out_3
rlabel metal3 s 357 1365 455 1463 4 vdd
rlabel metal3 s 357 4193 455 4291 4 vdd
rlabel metal3 s 1469 1365 1567 1463 4 vdd
rlabel metal3 s 1469 4193 1567 4291 4 vdd
rlabel metal3 s 1469 2779 1567 2877 4 gnd
rlabel metal3 s 357 2779 455 2877 4 gnd
rlabel metal3 s 1469 5607 1567 5705 4 gnd
rlabel metal3 s 357 -49 455 49 4 gnd
rlabel metal3 s 357 5607 455 5705 4 gnd
rlabel metal3 s 1469 -49 1567 49 4 gnd
<< properties >>
string FIXED_BBOX 0 0 2354 5656
<< end >>
