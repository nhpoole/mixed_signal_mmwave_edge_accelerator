magic
tech sky130A
magscale 1 2
timestamp 1623981280
<< nwell >>
rect 23294 14174 32818 17540
rect 12924 4730 22020 8734
rect 30172 8677 36115 8998
rect 30340 8676 36115 8677
rect 23506 8653 29390 8654
rect 23506 4730 29850 8653
rect 30172 7588 36114 8156
rect 30172 6500 36114 7068
rect 30172 5658 36114 5980
rect 8316 -1644 18832 4432
rect 23316 -1644 33832 4432
rect 12270 -13188 22786 -7112
rect 27270 -13188 37786 -7112
rect 8316 -19644 18832 -13568
rect 23316 -19644 33832 -13568
<< pwell >>
rect 23296 11020 32814 14118
rect 12924 8898 22020 10844
rect 29000 10770 29804 10774
rect 23506 8824 29804 10770
rect 23506 8818 29802 8824
rect 28994 8710 29802 8818
rect 30212 8212 36074 8620
rect 30212 7124 36074 7532
rect 30212 6036 36074 6444
rect 8316 -4174 18832 -1808
rect 23316 -4174 33832 -1808
rect 12270 -6948 22786 -4582
rect 27270 -6948 37786 -4582
rect 8316 -22174 18832 -19808
rect 23316 -22174 33832 -19808
<< nmos >>
rect 25331 13707 25531 13907
rect 25589 13707 25789 13907
rect 25847 13707 26047 13907
rect 26105 13707 26305 13907
rect 26363 13707 26563 13907
rect 26621 13707 26821 13907
rect 24296 12654 25096 12854
rect 25154 12654 25954 12854
rect 26012 12654 26812 12854
rect 26870 12654 27670 12854
rect 27728 12654 28528 12854
rect 28586 12654 29386 12854
rect 29444 12654 30244 12854
rect 30302 12654 31102 12854
rect 31160 12654 31960 12854
rect 24296 12072 25096 12272
rect 25154 12072 25954 12272
rect 26012 12072 26812 12272
rect 26870 12072 27670 12272
rect 27728 12072 28528 12272
rect 28586 12072 29386 12272
rect 29444 12072 30244 12272
rect 30302 12072 31102 12272
rect 31160 12072 31960 12272
rect 15214 9468 15614 9668
rect 15672 9468 16072 9668
rect 16130 9468 16530 9668
rect 16588 9468 16988 9668
rect 17046 9468 17446 9668
rect 17504 9468 17904 9668
rect 17962 9468 18362 9668
rect 18420 9468 18820 9668
rect 18878 9468 19278 9668
rect 19336 9468 19736 9668
rect 23976 9468 24376 9668
rect 24434 9468 24834 9668
rect 24892 9468 25292 9668
rect 25350 9468 25750 9668
rect 25808 9468 26208 9668
rect 26266 9468 26666 9668
rect 26724 9468 27124 9668
rect 27182 9468 27582 9668
rect 27640 9468 28040 9668
rect 28098 9468 28498 9668
rect 8824 -2414 9224 -2214
rect 9282 -2414 9682 -2214
rect 9740 -2414 10140 -2214
rect 10198 -2414 10598 -2214
rect 10656 -2414 11056 -2214
rect 11114 -2414 11514 -2214
rect 11572 -2414 11972 -2214
rect 12030 -2414 12430 -2214
rect 12488 -2414 12888 -2214
rect 12946 -2414 13346 -2214
rect 13824 -2414 14224 -2214
rect 14282 -2414 14682 -2214
rect 14740 -2414 15140 -2214
rect 15198 -2414 15598 -2214
rect 15656 -2414 16056 -2214
rect 16114 -2414 16514 -2214
rect 16572 -2414 16972 -2214
rect 17030 -2414 17430 -2214
rect 17488 -2414 17888 -2214
rect 17946 -2414 18346 -2214
rect 8824 -3082 9224 -2882
rect 9282 -3082 9682 -2882
rect 9740 -3082 10140 -2882
rect 10198 -3082 10598 -2882
rect 10656 -3082 11056 -2882
rect 11114 -3082 11514 -2882
rect 11572 -3082 11972 -2882
rect 12030 -3082 12430 -2882
rect 12488 -3082 12888 -2882
rect 12946 -3082 13346 -2882
rect 23824 -2414 24224 -2214
rect 24282 -2414 24682 -2214
rect 24740 -2414 25140 -2214
rect 25198 -2414 25598 -2214
rect 25656 -2414 26056 -2214
rect 26114 -2414 26514 -2214
rect 26572 -2414 26972 -2214
rect 27030 -2414 27430 -2214
rect 27488 -2414 27888 -2214
rect 27946 -2414 28346 -2214
rect 28824 -2414 29224 -2214
rect 29282 -2414 29682 -2214
rect 29740 -2414 30140 -2214
rect 30198 -2414 30598 -2214
rect 30656 -2414 31056 -2214
rect 31114 -2414 31514 -2214
rect 31572 -2414 31972 -2214
rect 32030 -2414 32430 -2214
rect 32488 -2414 32888 -2214
rect 32946 -2414 33346 -2214
rect 23824 -3082 24224 -2882
rect 24282 -3082 24682 -2882
rect 24740 -3082 25140 -2882
rect 25198 -3082 25598 -2882
rect 25656 -3082 26056 -2882
rect 26114 -3082 26514 -2882
rect 26572 -3082 26972 -2882
rect 27030 -3082 27430 -2882
rect 27488 -3082 27888 -2882
rect 27946 -3082 28346 -2882
rect 17756 -5874 18156 -5674
rect 18214 -5874 18614 -5674
rect 18672 -5874 19072 -5674
rect 19130 -5874 19530 -5674
rect 19588 -5874 19988 -5674
rect 20046 -5874 20446 -5674
rect 20504 -5874 20904 -5674
rect 20962 -5874 21362 -5674
rect 21420 -5874 21820 -5674
rect 21878 -5874 22278 -5674
rect 12756 -6542 13156 -6342
rect 13214 -6542 13614 -6342
rect 13672 -6542 14072 -6342
rect 14130 -6542 14530 -6342
rect 14588 -6542 14988 -6342
rect 15046 -6542 15446 -6342
rect 15504 -6542 15904 -6342
rect 15962 -6542 16362 -6342
rect 16420 -6542 16820 -6342
rect 16878 -6542 17278 -6342
rect 17756 -6542 18156 -6342
rect 18214 -6542 18614 -6342
rect 18672 -6542 19072 -6342
rect 19130 -6542 19530 -6342
rect 19588 -6542 19988 -6342
rect 20046 -6542 20446 -6342
rect 20504 -6542 20904 -6342
rect 20962 -6542 21362 -6342
rect 21420 -6542 21820 -6342
rect 21878 -6542 22278 -6342
rect 32756 -5874 33156 -5674
rect 33214 -5874 33614 -5674
rect 33672 -5874 34072 -5674
rect 34130 -5874 34530 -5674
rect 34588 -5874 34988 -5674
rect 35046 -5874 35446 -5674
rect 35504 -5874 35904 -5674
rect 35962 -5874 36362 -5674
rect 36420 -5874 36820 -5674
rect 36878 -5874 37278 -5674
rect 27756 -6542 28156 -6342
rect 28214 -6542 28614 -6342
rect 28672 -6542 29072 -6342
rect 29130 -6542 29530 -6342
rect 29588 -6542 29988 -6342
rect 30046 -6542 30446 -6342
rect 30504 -6542 30904 -6342
rect 30962 -6542 31362 -6342
rect 31420 -6542 31820 -6342
rect 31878 -6542 32278 -6342
rect 32756 -6542 33156 -6342
rect 33214 -6542 33614 -6342
rect 33672 -6542 34072 -6342
rect 34130 -6542 34530 -6342
rect 34588 -6542 34988 -6342
rect 35046 -6542 35446 -6342
rect 35504 -6542 35904 -6342
rect 35962 -6542 36362 -6342
rect 36420 -6542 36820 -6342
rect 36878 -6542 37278 -6342
rect 8824 -20414 9224 -20214
rect 9282 -20414 9682 -20214
rect 9740 -20414 10140 -20214
rect 10198 -20414 10598 -20214
rect 10656 -20414 11056 -20214
rect 11114 -20414 11514 -20214
rect 11572 -20414 11972 -20214
rect 12030 -20414 12430 -20214
rect 12488 -20414 12888 -20214
rect 12946 -20414 13346 -20214
rect 13824 -20414 14224 -20214
rect 14282 -20414 14682 -20214
rect 14740 -20414 15140 -20214
rect 15198 -20414 15598 -20214
rect 15656 -20414 16056 -20214
rect 16114 -20414 16514 -20214
rect 16572 -20414 16972 -20214
rect 17030 -20414 17430 -20214
rect 17488 -20414 17888 -20214
rect 17946 -20414 18346 -20214
rect 8824 -21082 9224 -20882
rect 9282 -21082 9682 -20882
rect 9740 -21082 10140 -20882
rect 10198 -21082 10598 -20882
rect 10656 -21082 11056 -20882
rect 11114 -21082 11514 -20882
rect 11572 -21082 11972 -20882
rect 12030 -21082 12430 -20882
rect 12488 -21082 12888 -20882
rect 12946 -21082 13346 -20882
rect 23824 -20414 24224 -20214
rect 24282 -20414 24682 -20214
rect 24740 -20414 25140 -20214
rect 25198 -20414 25598 -20214
rect 25656 -20414 26056 -20214
rect 26114 -20414 26514 -20214
rect 26572 -20414 26972 -20214
rect 27030 -20414 27430 -20214
rect 27488 -20414 27888 -20214
rect 27946 -20414 28346 -20214
rect 28824 -20414 29224 -20214
rect 29282 -20414 29682 -20214
rect 29740 -20414 30140 -20214
rect 30198 -20414 30598 -20214
rect 30656 -20414 31056 -20214
rect 31114 -20414 31514 -20214
rect 31572 -20414 31972 -20214
rect 32030 -20414 32430 -20214
rect 32488 -20414 32888 -20214
rect 32946 -20414 33346 -20214
rect 23824 -21082 24224 -20882
rect 24282 -21082 24682 -20882
rect 24740 -21082 25140 -20882
rect 25198 -21082 25598 -20882
rect 25656 -21082 26056 -20882
rect 26114 -21082 26514 -20882
rect 26572 -21082 26972 -20882
rect 27030 -21082 27430 -20882
rect 27488 -21082 27888 -20882
rect 27946 -21082 28346 -20882
<< scnmos >>
rect 27339 13961 27369 14045
rect 27423 13961 27453 14045
rect 27678 13961 27708 14045
rect 27773 13961 27803 14033
rect 27869 13961 27899 14033
rect 28035 13961 28065 14045
rect 28107 13961 28137 14045
rect 28239 13961 28269 14089
rect 28338 13961 28368 14033
rect 28447 13961 28477 14033
rect 28543 13961 28573 14045
rect 28692 13961 28722 14045
rect 28783 13961 28813 14045
rect 28971 13961 29001 14091
rect 29159 13961 29189 14045
rect 29256 13961 29286 14091
rect 29496 13961 29526 14091
rect 29735 13961 29765 14091
rect 29819 13961 29849 14091
rect 30054 13961 30084 14091
rect 30294 13961 30324 14091
rect 30391 13961 30421 14045
rect 30579 13961 30609 14091
rect 30767 13961 30797 14045
rect 30858 13961 30888 14045
rect 31007 13961 31037 14045
rect 31103 13961 31133 14033
rect 31212 13961 31242 14033
rect 31311 13961 31341 14089
rect 31443 13961 31473 14045
rect 31515 13961 31545 14045
rect 31681 13961 31711 14033
rect 31777 13961 31807 14033
rect 31872 13961 31902 14045
rect 32127 13961 32157 14045
rect 32211 13961 32241 14045
rect 29196 8737 29226 8867
rect 29441 8737 29471 8867
rect 29525 8737 29555 8867
rect 29609 8737 29639 8867
rect 29693 8737 29723 8867
rect 30631 8463 30661 8547
rect 30715 8463 30745 8547
rect 30903 8463 30933 8547
rect 31015 8463 31045 8535
rect 31114 8463 31144 8535
rect 31213 8463 31243 8547
rect 31332 8463 31362 8591
rect 31433 8463 31463 8535
rect 31539 8463 31569 8535
rect 31634 8463 31664 8547
rect 31824 8463 31854 8593
rect 31908 8463 31938 8593
rect 32096 8463 32126 8547
rect 32191 8463 32221 8593
rect 32420 8463 32450 8593
rect 32665 8463 32695 8593
rect 32749 8463 32779 8593
rect 32833 8463 32863 8593
rect 32917 8463 32947 8593
rect 30631 8285 30661 8369
rect 30715 8285 30745 8369
rect 30903 8285 30933 8369
rect 31015 8297 31045 8369
rect 31114 8297 31144 8369
rect 31213 8285 31243 8369
rect 31332 8241 31362 8369
rect 31433 8297 31463 8369
rect 31539 8297 31569 8369
rect 31634 8285 31664 8369
rect 31824 8239 31854 8369
rect 31908 8239 31938 8369
rect 32096 8285 32126 8369
rect 32191 8239 32221 8369
rect 32420 8239 32450 8369
rect 32665 8239 32695 8369
rect 32749 8239 32779 8369
rect 32833 8239 32863 8369
rect 32917 8239 32947 8369
rect 33329 8285 33359 8369
rect 33413 8285 33443 8369
rect 33601 8285 33631 8369
rect 33713 8297 33743 8369
rect 33812 8297 33842 8369
rect 33911 8285 33941 8369
rect 34030 8241 34060 8369
rect 34131 8297 34161 8369
rect 34237 8297 34267 8369
rect 34332 8285 34362 8369
rect 34522 8239 34552 8369
rect 34606 8239 34636 8369
rect 34794 8285 34824 8369
rect 34889 8239 34919 8369
rect 35118 8239 35148 8369
rect 35363 8239 35393 8369
rect 35447 8239 35477 8369
rect 35531 8239 35561 8369
rect 35615 8239 35645 8369
rect 30631 7375 30661 7459
rect 30715 7375 30745 7459
rect 30903 7375 30933 7459
rect 31015 7375 31045 7447
rect 31114 7375 31144 7447
rect 31213 7375 31243 7459
rect 31332 7375 31362 7503
rect 31433 7375 31463 7447
rect 31539 7375 31569 7447
rect 31634 7375 31664 7459
rect 31824 7375 31854 7505
rect 31908 7375 31938 7505
rect 32096 7375 32126 7459
rect 32191 7375 32221 7505
rect 32420 7375 32450 7505
rect 32665 7375 32695 7505
rect 32749 7375 32779 7505
rect 32833 7375 32863 7505
rect 32917 7375 32947 7505
rect 33329 7375 33359 7459
rect 33413 7375 33443 7459
rect 33601 7375 33631 7459
rect 33713 7375 33743 7447
rect 33812 7375 33842 7447
rect 33911 7375 33941 7459
rect 34030 7375 34060 7503
rect 34131 7375 34161 7447
rect 34237 7375 34267 7447
rect 34332 7375 34362 7459
rect 34522 7375 34552 7505
rect 34606 7375 34636 7505
rect 34794 7375 34824 7459
rect 34889 7375 34919 7505
rect 35118 7375 35148 7505
rect 35363 7375 35393 7505
rect 35447 7375 35477 7505
rect 35531 7375 35561 7505
rect 35615 7375 35645 7505
rect 30631 7197 30661 7281
rect 30715 7197 30745 7281
rect 30903 7197 30933 7281
rect 31015 7209 31045 7281
rect 31114 7209 31144 7281
rect 31213 7197 31243 7281
rect 31332 7153 31362 7281
rect 31433 7209 31463 7281
rect 31539 7209 31569 7281
rect 31634 7197 31664 7281
rect 31824 7151 31854 7281
rect 31908 7151 31938 7281
rect 32096 7197 32126 7281
rect 32191 7151 32221 7281
rect 32420 7151 32450 7281
rect 32665 7151 32695 7281
rect 32749 7151 32779 7281
rect 32833 7151 32863 7281
rect 32917 7151 32947 7281
rect 33329 7197 33359 7281
rect 33413 7197 33443 7281
rect 33601 7197 33631 7281
rect 33713 7209 33743 7281
rect 33812 7209 33842 7281
rect 33911 7197 33941 7281
rect 34030 7153 34060 7281
rect 34131 7209 34161 7281
rect 34237 7209 34267 7281
rect 34332 7197 34362 7281
rect 34522 7151 34552 7281
rect 34606 7151 34636 7281
rect 34794 7197 34824 7281
rect 34889 7151 34919 7281
rect 35118 7151 35148 7281
rect 35363 7151 35393 7281
rect 35447 7151 35477 7281
rect 35531 7151 35561 7281
rect 35615 7151 35645 7281
rect 30631 6287 30661 6371
rect 30715 6287 30745 6371
rect 30903 6287 30933 6371
rect 31015 6287 31045 6359
rect 31114 6287 31144 6359
rect 31213 6287 31243 6371
rect 31332 6287 31362 6415
rect 31433 6287 31463 6359
rect 31539 6287 31569 6359
rect 31634 6287 31664 6371
rect 31824 6287 31854 6417
rect 31908 6287 31938 6417
rect 32096 6287 32126 6371
rect 32191 6287 32221 6417
rect 32420 6287 32450 6417
rect 32665 6287 32695 6417
rect 32749 6287 32779 6417
rect 32833 6287 32863 6417
rect 32917 6287 32947 6417
rect 33329 6287 33359 6371
rect 33413 6287 33443 6371
rect 33601 6287 33631 6371
rect 33713 6287 33743 6359
rect 33812 6287 33842 6359
rect 33911 6287 33941 6371
rect 34030 6287 34060 6415
rect 34131 6287 34161 6359
rect 34237 6287 34267 6359
rect 34332 6287 34362 6371
rect 34522 6287 34552 6417
rect 34606 6287 34636 6417
rect 34794 6287 34824 6371
rect 34889 6287 34919 6417
rect 35118 6287 35148 6417
rect 35363 6287 35393 6417
rect 35447 6287 35477 6417
rect 35531 6287 35561 6417
rect 35615 6287 35645 6417
rect 30631 6109 30661 6193
rect 30715 6109 30745 6193
rect 30903 6109 30933 6193
rect 31015 6121 31045 6193
rect 31114 6121 31144 6193
rect 31213 6109 31243 6193
rect 31332 6065 31362 6193
rect 31433 6121 31463 6193
rect 31539 6121 31569 6193
rect 31634 6109 31664 6193
rect 31824 6063 31854 6193
rect 31908 6063 31938 6193
rect 32096 6109 32126 6193
rect 32191 6063 32221 6193
rect 32420 6063 32450 6193
rect 32665 6063 32695 6193
rect 32749 6063 32779 6193
rect 32833 6063 32863 6193
rect 32917 6063 32947 6193
rect 33329 6109 33359 6193
rect 33413 6109 33443 6193
rect 33601 6109 33631 6193
rect 33713 6121 33743 6193
rect 33812 6121 33842 6193
rect 33911 6109 33941 6193
rect 34030 6065 34060 6193
rect 34131 6121 34161 6193
rect 34237 6121 34267 6193
rect 34332 6109 34362 6193
rect 34522 6063 34552 6193
rect 34606 6063 34636 6193
rect 34794 6109 34824 6193
rect 34889 6063 34919 6193
rect 35118 6063 35148 6193
rect 35363 6063 35393 6193
rect 35447 6063 35477 6193
rect 35531 6063 35561 6193
rect 35615 6063 35645 6193
<< pmos >>
rect 23822 16234 24622 16434
rect 24680 16234 25480 16434
rect 25538 16234 26338 16434
rect 26396 16234 27196 16434
rect 27254 16234 28054 16434
rect 28112 16234 28912 16434
rect 28970 16234 29770 16434
rect 29828 16234 30628 16434
rect 30686 16234 31486 16434
rect 31544 16234 32344 16434
rect 23822 15634 24622 15834
rect 24680 15634 25480 15834
rect 25538 15634 26338 15834
rect 26396 15634 27196 15834
rect 27254 15634 28054 15834
rect 28112 15634 28912 15834
rect 28970 15634 29770 15834
rect 29828 15634 30628 15834
rect 30686 15634 31486 15834
rect 31544 15634 32344 15834
rect 25331 14394 25531 14794
rect 25589 14394 25789 14794
rect 25847 14394 26047 14794
rect 26105 14394 26305 14794
rect 26363 14394 26563 14794
rect 26621 14394 26821 14794
<< scpmoshvt >>
rect 27339 14277 27369 14405
rect 27423 14277 27453 14405
rect 27690 14327 27720 14411
rect 27782 14327 27812 14411
rect 27881 14327 27911 14411
rect 28021 14327 28051 14411
rect 28118 14327 28148 14411
rect 28315 14243 28345 14411
rect 28414 14327 28444 14411
rect 28500 14327 28530 14411
rect 28584 14327 28614 14411
rect 28692 14327 28722 14411
rect 28776 14327 28806 14411
rect 28940 14211 28970 14411
rect 29159 14283 29189 14411
rect 29256 14211 29286 14411
rect 29496 14211 29526 14411
rect 29735 14211 29765 14411
rect 29819 14211 29849 14411
rect 30054 14211 30084 14411
rect 30294 14211 30324 14411
rect 30391 14283 30421 14411
rect 30610 14211 30640 14411
rect 30774 14327 30804 14411
rect 30858 14327 30888 14411
rect 30966 14327 30996 14411
rect 31050 14327 31080 14411
rect 31136 14327 31166 14411
rect 31235 14243 31265 14411
rect 31432 14327 31462 14411
rect 31529 14327 31559 14411
rect 31669 14327 31699 14411
rect 31768 14327 31798 14411
rect 31860 14327 31890 14411
rect 32127 14277 32157 14405
rect 32211 14277 32241 14405
rect 30631 8779 30661 8907
rect 30715 8779 30745 8907
rect 30903 8829 30933 8913
rect 30988 8829 31018 8913
rect 31083 8829 31113 8913
rect 31186 8829 31216 8913
rect 29196 8417 29226 8617
rect 29441 8417 29471 8617
rect 29525 8417 29555 8617
rect 29609 8417 29639 8617
rect 29693 8417 29723 8617
rect 31318 8763 31348 8913
rect 31413 8829 31443 8913
rect 31497 8829 31527 8913
rect 31611 8829 31641 8913
rect 31822 8713 31852 8913
rect 31906 8713 31936 8913
rect 32094 8785 32124 8913
rect 32191 8713 32221 8913
rect 32420 8713 32450 8913
rect 32665 8713 32695 8913
rect 32749 8713 32779 8913
rect 32833 8713 32863 8913
rect 32917 8713 32947 8913
rect 30631 7925 30661 8053
rect 30715 7925 30745 8053
rect 30903 7919 30933 8003
rect 30988 7919 31018 8003
rect 31083 7919 31113 8003
rect 31186 7919 31216 8003
rect 31318 7919 31348 8069
rect 31413 7919 31443 8003
rect 31497 7919 31527 8003
rect 31611 7919 31641 8003
rect 31822 7919 31852 8119
rect 31906 7919 31936 8119
rect 32094 7919 32124 8047
rect 32191 7919 32221 8119
rect 32420 7919 32450 8119
rect 32665 7919 32695 8119
rect 32749 7919 32779 8119
rect 32833 7919 32863 8119
rect 32917 7919 32947 8119
rect 33329 7925 33359 8053
rect 33413 7925 33443 8053
rect 33601 7919 33631 8003
rect 33686 7919 33716 8003
rect 33781 7919 33811 8003
rect 33884 7919 33914 8003
rect 34016 7919 34046 8069
rect 34111 7919 34141 8003
rect 34195 7919 34225 8003
rect 34309 7919 34339 8003
rect 34520 7919 34550 8119
rect 34604 7919 34634 8119
rect 34792 7919 34822 8047
rect 34889 7919 34919 8119
rect 35118 7919 35148 8119
rect 35363 7919 35393 8119
rect 35447 7919 35477 8119
rect 35531 7919 35561 8119
rect 35615 7919 35645 8119
rect 30631 7691 30661 7819
rect 30715 7691 30745 7819
rect 30903 7741 30933 7825
rect 30988 7741 31018 7825
rect 31083 7741 31113 7825
rect 31186 7741 31216 7825
rect 31318 7675 31348 7825
rect 31413 7741 31443 7825
rect 31497 7741 31527 7825
rect 31611 7741 31641 7825
rect 31822 7625 31852 7825
rect 31906 7625 31936 7825
rect 32094 7697 32124 7825
rect 32191 7625 32221 7825
rect 32420 7625 32450 7825
rect 32665 7625 32695 7825
rect 32749 7625 32779 7825
rect 32833 7625 32863 7825
rect 32917 7625 32947 7825
rect 33329 7691 33359 7819
rect 33413 7691 33443 7819
rect 33601 7741 33631 7825
rect 33686 7741 33716 7825
rect 33781 7741 33811 7825
rect 33884 7741 33914 7825
rect 34016 7675 34046 7825
rect 34111 7741 34141 7825
rect 34195 7741 34225 7825
rect 34309 7741 34339 7825
rect 34520 7625 34550 7825
rect 34604 7625 34634 7825
rect 34792 7697 34822 7825
rect 34889 7625 34919 7825
rect 35118 7625 35148 7825
rect 35363 7625 35393 7825
rect 35447 7625 35477 7825
rect 35531 7625 35561 7825
rect 35615 7625 35645 7825
rect 30631 6837 30661 6965
rect 30715 6837 30745 6965
rect 30903 6831 30933 6915
rect 30988 6831 31018 6915
rect 31083 6831 31113 6915
rect 31186 6831 31216 6915
rect 31318 6831 31348 6981
rect 31413 6831 31443 6915
rect 31497 6831 31527 6915
rect 31611 6831 31641 6915
rect 31822 6831 31852 7031
rect 31906 6831 31936 7031
rect 32094 6831 32124 6959
rect 32191 6831 32221 7031
rect 32420 6831 32450 7031
rect 32665 6831 32695 7031
rect 32749 6831 32779 7031
rect 32833 6831 32863 7031
rect 32917 6831 32947 7031
rect 33329 6837 33359 6965
rect 33413 6837 33443 6965
rect 33601 6831 33631 6915
rect 33686 6831 33716 6915
rect 33781 6831 33811 6915
rect 33884 6831 33914 6915
rect 34016 6831 34046 6981
rect 34111 6831 34141 6915
rect 34195 6831 34225 6915
rect 34309 6831 34339 6915
rect 34520 6831 34550 7031
rect 34604 6831 34634 7031
rect 34792 6831 34822 6959
rect 34889 6831 34919 7031
rect 35118 6831 35148 7031
rect 35363 6831 35393 7031
rect 35447 6831 35477 7031
rect 35531 6831 35561 7031
rect 35615 6831 35645 7031
rect 30631 6603 30661 6731
rect 30715 6603 30745 6731
rect 30903 6653 30933 6737
rect 30988 6653 31018 6737
rect 31083 6653 31113 6737
rect 31186 6653 31216 6737
rect 31318 6587 31348 6737
rect 31413 6653 31443 6737
rect 31497 6653 31527 6737
rect 31611 6653 31641 6737
rect 31822 6537 31852 6737
rect 31906 6537 31936 6737
rect 32094 6609 32124 6737
rect 32191 6537 32221 6737
rect 32420 6537 32450 6737
rect 32665 6537 32695 6737
rect 32749 6537 32779 6737
rect 32833 6537 32863 6737
rect 32917 6537 32947 6737
rect 33329 6603 33359 6731
rect 33413 6603 33443 6731
rect 33601 6653 33631 6737
rect 33686 6653 33716 6737
rect 33781 6653 33811 6737
rect 33884 6653 33914 6737
rect 34016 6587 34046 6737
rect 34111 6653 34141 6737
rect 34195 6653 34225 6737
rect 34309 6653 34339 6737
rect 34520 6537 34550 6737
rect 34604 6537 34634 6737
rect 34792 6609 34822 6737
rect 34889 6537 34919 6737
rect 35118 6537 35148 6737
rect 35363 6537 35393 6737
rect 35447 6537 35477 6737
rect 35531 6537 35561 6737
rect 35615 6537 35645 6737
rect 30631 5749 30661 5877
rect 30715 5749 30745 5877
rect 30903 5743 30933 5827
rect 30988 5743 31018 5827
rect 31083 5743 31113 5827
rect 31186 5743 31216 5827
rect 31318 5743 31348 5893
rect 31413 5743 31443 5827
rect 31497 5743 31527 5827
rect 31611 5743 31641 5827
rect 31822 5743 31852 5943
rect 31906 5743 31936 5943
rect 32094 5743 32124 5871
rect 32191 5743 32221 5943
rect 32420 5743 32450 5943
rect 32665 5743 32695 5943
rect 32749 5743 32779 5943
rect 32833 5743 32863 5943
rect 32917 5743 32947 5943
rect 33329 5749 33359 5877
rect 33413 5749 33443 5877
rect 33601 5743 33631 5827
rect 33686 5743 33716 5827
rect 33781 5743 33811 5827
rect 33884 5743 33914 5827
rect 34016 5743 34046 5893
rect 34111 5743 34141 5827
rect 34195 5743 34225 5827
rect 34309 5743 34339 5827
rect 34520 5743 34550 5943
rect 34604 5743 34634 5943
rect 34792 5743 34822 5871
rect 34889 5743 34919 5943
rect 35118 5743 35148 5943
rect 35363 5743 35393 5943
rect 35447 5743 35477 5943
rect 35531 5743 35561 5943
rect 35615 5743 35645 5943
<< pmoslvt >>
rect 24209 14394 24409 14794
rect 24467 14394 24667 14794
rect 24725 14394 24925 14794
<< pmoshvt >>
rect 13382 6217 13782 7817
rect 13840 6217 14240 7817
rect 14298 6217 14698 7817
rect 14756 6217 15156 7817
rect 15214 6217 15614 7817
rect 15672 6217 16072 7817
rect 16130 6217 16530 7817
rect 16588 6217 16988 7817
rect 17046 6217 17446 7817
rect 17504 6217 17904 7817
rect 17962 6217 18362 7817
rect 18420 6217 18820 7817
rect 18878 6217 19278 7817
rect 19336 6217 19736 7817
rect 19794 6217 20194 7817
rect 20252 6217 20652 7817
rect 20710 6217 21110 7817
rect 21168 6217 21568 7817
rect 23977 7037 24377 8237
rect 24435 7037 24835 8237
rect 24893 7037 25293 8237
rect 25351 7037 25751 8237
rect 25809 7037 26209 8237
rect 26267 7037 26667 8237
rect 26725 7037 27125 8237
rect 27183 7037 27583 8237
rect 27641 7037 28041 8237
rect 28099 7037 28499 8237
rect 9384 1344 9784 2944
rect 9842 1344 10242 2944
rect 10300 1344 10700 2944
rect 10758 1344 11158 2944
rect 11216 1344 11616 2944
rect 11674 1344 12074 2944
rect 12132 1344 12532 2944
rect 12590 1344 12990 2944
rect 13048 1344 13448 2944
rect 13506 1344 13906 2944
rect 13964 1344 14364 2944
rect 14422 1344 14822 2944
rect 14880 1344 15280 2944
rect 15338 1344 15738 2944
rect 15796 1344 16196 2944
rect 16254 1344 16654 2944
rect 16712 1344 17112 2944
rect 17170 1344 17570 2944
rect 8825 -921 9225 279
rect 9283 -921 9683 279
rect 9741 -921 10141 279
rect 10199 -921 10599 279
rect 10657 -921 11057 279
rect 11115 -921 11515 279
rect 11573 -921 11973 279
rect 12031 -921 12431 279
rect 12489 -921 12889 279
rect 12947 -921 13347 279
rect 13825 -921 14225 279
rect 14283 -921 14683 279
rect 14741 -921 15141 279
rect 15199 -921 15599 279
rect 15657 -921 16057 279
rect 16115 -921 16515 279
rect 16573 -921 16973 279
rect 17031 -921 17431 279
rect 17489 -921 17889 279
rect 17947 -921 18347 279
rect 24384 1344 24784 2944
rect 24842 1344 25242 2944
rect 25300 1344 25700 2944
rect 25758 1344 26158 2944
rect 26216 1344 26616 2944
rect 26674 1344 27074 2944
rect 27132 1344 27532 2944
rect 27590 1344 27990 2944
rect 28048 1344 28448 2944
rect 28506 1344 28906 2944
rect 28964 1344 29364 2944
rect 29422 1344 29822 2944
rect 29880 1344 30280 2944
rect 30338 1344 30738 2944
rect 30796 1344 31196 2944
rect 31254 1344 31654 2944
rect 31712 1344 32112 2944
rect 32170 1344 32570 2944
rect 23825 -921 24225 279
rect 24283 -921 24683 279
rect 24741 -921 25141 279
rect 25199 -921 25599 279
rect 25657 -921 26057 279
rect 26115 -921 26515 279
rect 26573 -921 26973 279
rect 27031 -921 27431 279
rect 27489 -921 27889 279
rect 27947 -921 28347 279
rect 28825 -921 29225 279
rect 29283 -921 29683 279
rect 29741 -921 30141 279
rect 30199 -921 30599 279
rect 30657 -921 31057 279
rect 31115 -921 31515 279
rect 31573 -921 31973 279
rect 32031 -921 32431 279
rect 32489 -921 32889 279
rect 32947 -921 33347 279
rect 12755 -9035 13155 -7835
rect 13213 -9035 13613 -7835
rect 13671 -9035 14071 -7835
rect 14129 -9035 14529 -7835
rect 14587 -9035 14987 -7835
rect 15045 -9035 15445 -7835
rect 15503 -9035 15903 -7835
rect 15961 -9035 16361 -7835
rect 16419 -9035 16819 -7835
rect 16877 -9035 17277 -7835
rect 17755 -9035 18155 -7835
rect 18213 -9035 18613 -7835
rect 18671 -9035 19071 -7835
rect 19129 -9035 19529 -7835
rect 19587 -9035 19987 -7835
rect 20045 -9035 20445 -7835
rect 20503 -9035 20903 -7835
rect 20961 -9035 21361 -7835
rect 21419 -9035 21819 -7835
rect 21877 -9035 22277 -7835
rect 13532 -11700 13932 -10100
rect 13990 -11700 14390 -10100
rect 14448 -11700 14848 -10100
rect 14906 -11700 15306 -10100
rect 15364 -11700 15764 -10100
rect 15822 -11700 16222 -10100
rect 16280 -11700 16680 -10100
rect 16738 -11700 17138 -10100
rect 17196 -11700 17596 -10100
rect 17654 -11700 18054 -10100
rect 18112 -11700 18512 -10100
rect 18570 -11700 18970 -10100
rect 19028 -11700 19428 -10100
rect 19486 -11700 19886 -10100
rect 19944 -11700 20344 -10100
rect 20402 -11700 20802 -10100
rect 20860 -11700 21260 -10100
rect 21318 -11700 21718 -10100
rect 27755 -9035 28155 -7835
rect 28213 -9035 28613 -7835
rect 28671 -9035 29071 -7835
rect 29129 -9035 29529 -7835
rect 29587 -9035 29987 -7835
rect 30045 -9035 30445 -7835
rect 30503 -9035 30903 -7835
rect 30961 -9035 31361 -7835
rect 31419 -9035 31819 -7835
rect 31877 -9035 32277 -7835
rect 32755 -9035 33155 -7835
rect 33213 -9035 33613 -7835
rect 33671 -9035 34071 -7835
rect 34129 -9035 34529 -7835
rect 34587 -9035 34987 -7835
rect 35045 -9035 35445 -7835
rect 35503 -9035 35903 -7835
rect 35961 -9035 36361 -7835
rect 36419 -9035 36819 -7835
rect 36877 -9035 37277 -7835
rect 28532 -11700 28932 -10100
rect 28990 -11700 29390 -10100
rect 29448 -11700 29848 -10100
rect 29906 -11700 30306 -10100
rect 30364 -11700 30764 -10100
rect 30822 -11700 31222 -10100
rect 31280 -11700 31680 -10100
rect 31738 -11700 32138 -10100
rect 32196 -11700 32596 -10100
rect 32654 -11700 33054 -10100
rect 33112 -11700 33512 -10100
rect 33570 -11700 33970 -10100
rect 34028 -11700 34428 -10100
rect 34486 -11700 34886 -10100
rect 34944 -11700 35344 -10100
rect 35402 -11700 35802 -10100
rect 35860 -11700 36260 -10100
rect 36318 -11700 36718 -10100
rect 9384 -16656 9784 -15056
rect 9842 -16656 10242 -15056
rect 10300 -16656 10700 -15056
rect 10758 -16656 11158 -15056
rect 11216 -16656 11616 -15056
rect 11674 -16656 12074 -15056
rect 12132 -16656 12532 -15056
rect 12590 -16656 12990 -15056
rect 13048 -16656 13448 -15056
rect 13506 -16656 13906 -15056
rect 13964 -16656 14364 -15056
rect 14422 -16656 14822 -15056
rect 14880 -16656 15280 -15056
rect 15338 -16656 15738 -15056
rect 15796 -16656 16196 -15056
rect 16254 -16656 16654 -15056
rect 16712 -16656 17112 -15056
rect 17170 -16656 17570 -15056
rect 8825 -18921 9225 -17721
rect 9283 -18921 9683 -17721
rect 9741 -18921 10141 -17721
rect 10199 -18921 10599 -17721
rect 10657 -18921 11057 -17721
rect 11115 -18921 11515 -17721
rect 11573 -18921 11973 -17721
rect 12031 -18921 12431 -17721
rect 12489 -18921 12889 -17721
rect 12947 -18921 13347 -17721
rect 13825 -18921 14225 -17721
rect 14283 -18921 14683 -17721
rect 14741 -18921 15141 -17721
rect 15199 -18921 15599 -17721
rect 15657 -18921 16057 -17721
rect 16115 -18921 16515 -17721
rect 16573 -18921 16973 -17721
rect 17031 -18921 17431 -17721
rect 17489 -18921 17889 -17721
rect 17947 -18921 18347 -17721
rect 24384 -16656 24784 -15056
rect 24842 -16656 25242 -15056
rect 25300 -16656 25700 -15056
rect 25758 -16656 26158 -15056
rect 26216 -16656 26616 -15056
rect 26674 -16656 27074 -15056
rect 27132 -16656 27532 -15056
rect 27590 -16656 27990 -15056
rect 28048 -16656 28448 -15056
rect 28506 -16656 28906 -15056
rect 28964 -16656 29364 -15056
rect 29422 -16656 29822 -15056
rect 29880 -16656 30280 -15056
rect 30338 -16656 30738 -15056
rect 30796 -16656 31196 -15056
rect 31254 -16656 31654 -15056
rect 31712 -16656 32112 -15056
rect 32170 -16656 32570 -15056
rect 23825 -18921 24225 -17721
rect 24283 -18921 24683 -17721
rect 24741 -18921 25141 -17721
rect 25199 -18921 25599 -17721
rect 25657 -18921 26057 -17721
rect 26115 -18921 26515 -17721
rect 26573 -18921 26973 -17721
rect 27031 -18921 27431 -17721
rect 27489 -18921 27889 -17721
rect 27947 -18921 28347 -17721
rect 28825 -18921 29225 -17721
rect 29283 -18921 29683 -17721
rect 29741 -18921 30141 -17721
rect 30199 -18921 30599 -17721
rect 30657 -18921 31057 -17721
rect 31115 -18921 31515 -17721
rect 31573 -18921 31973 -17721
rect 32031 -18921 32431 -17721
rect 32489 -18921 32889 -17721
rect 32947 -18921 33347 -17721
<< nmoslvt >>
rect 24209 13707 24409 13907
rect 24467 13707 24667 13907
rect 24725 13707 24925 13907
<< ndiff >>
rect 24151 13895 24209 13907
rect 24151 13719 24163 13895
rect 24197 13719 24209 13895
rect 24151 13707 24209 13719
rect 24409 13895 24467 13907
rect 24409 13719 24421 13895
rect 24455 13719 24467 13895
rect 24409 13707 24467 13719
rect 24667 13895 24725 13907
rect 24667 13719 24679 13895
rect 24713 13719 24725 13895
rect 24667 13707 24725 13719
rect 24925 13895 24983 13907
rect 24925 13719 24937 13895
rect 24971 13719 24983 13895
rect 24925 13707 24983 13719
rect 25273 13895 25331 13907
rect 25273 13719 25285 13895
rect 25319 13719 25331 13895
rect 25273 13707 25331 13719
rect 25531 13895 25589 13907
rect 25531 13719 25543 13895
rect 25577 13719 25589 13895
rect 25531 13707 25589 13719
rect 25789 13895 25847 13907
rect 25789 13719 25801 13895
rect 25835 13719 25847 13895
rect 25789 13707 25847 13719
rect 26047 13895 26105 13907
rect 26047 13719 26059 13895
rect 26093 13719 26105 13895
rect 26047 13707 26105 13719
rect 26305 13895 26363 13907
rect 26305 13719 26317 13895
rect 26351 13719 26363 13895
rect 26305 13707 26363 13719
rect 26563 13895 26621 13907
rect 26563 13719 26575 13895
rect 26609 13719 26621 13895
rect 26563 13707 26621 13719
rect 26821 13895 26879 13907
rect 26821 13719 26833 13895
rect 26867 13719 26879 13895
rect 26821 13707 26879 13719
rect 27287 14033 27339 14045
rect 27287 13999 27295 14033
rect 27329 13999 27339 14033
rect 27287 13961 27339 13999
rect 27369 14007 27423 14045
rect 27369 13973 27379 14007
rect 27413 13973 27423 14007
rect 27369 13961 27423 13973
rect 27453 14033 27505 14045
rect 27453 13999 27463 14033
rect 27497 13999 27505 14033
rect 27453 13961 27505 13999
rect 27573 14003 27678 14045
rect 27573 13969 27585 14003
rect 27619 13969 27678 14003
rect 27573 13961 27678 13969
rect 27708 14033 27758 14045
rect 28189 14045 28239 14089
rect 27917 14033 28035 14045
rect 27708 14009 27773 14033
rect 27708 13975 27718 14009
rect 27752 13975 27773 14009
rect 27708 13961 27773 13975
rect 27803 14009 27869 14033
rect 27803 13975 27825 14009
rect 27859 13975 27869 14009
rect 27803 13961 27869 13975
rect 27899 13961 28035 14033
rect 28065 13961 28107 14045
rect 28137 14007 28239 14045
rect 28137 13973 28171 14007
rect 28205 13973 28239 14007
rect 28137 13961 28239 13973
rect 28269 14033 28323 14089
rect 28919 14046 28971 14091
rect 28493 14033 28543 14045
rect 28269 14003 28338 14033
rect 28269 13969 28283 14003
rect 28317 13969 28338 14003
rect 28269 13961 28338 13969
rect 28368 14007 28447 14033
rect 28368 13973 28393 14007
rect 28427 13973 28447 14007
rect 28368 13961 28447 13973
rect 28477 13961 28543 14033
rect 28573 14003 28692 14045
rect 28573 13969 28605 14003
rect 28639 13969 28692 14003
rect 28573 13961 28692 13969
rect 28722 13961 28783 14045
rect 28813 14023 28865 14045
rect 28813 13989 28823 14023
rect 28857 13989 28865 14023
rect 28813 13961 28865 13989
rect 28919 14012 28927 14046
rect 28961 14012 28971 14046
rect 28919 13961 28971 14012
rect 29001 14079 29053 14091
rect 29001 14045 29011 14079
rect 29045 14045 29053 14079
rect 29204 14045 29256 14091
rect 29001 14011 29053 14045
rect 29001 13977 29011 14011
rect 29045 13977 29053 14011
rect 29001 13961 29053 13977
rect 29107 14033 29159 14045
rect 29107 13999 29115 14033
rect 29149 13999 29159 14033
rect 29107 13961 29159 13999
rect 29189 14027 29256 14045
rect 29189 13993 29212 14027
rect 29246 13993 29256 14027
rect 29189 13961 29256 13993
rect 29286 14057 29338 14091
rect 29286 14023 29296 14057
rect 29330 14023 29338 14057
rect 29286 13961 29338 14023
rect 29444 14079 29496 14091
rect 29444 14045 29452 14079
rect 29486 14045 29496 14079
rect 29444 14011 29496 14045
rect 29444 13977 29452 14011
rect 29486 13977 29496 14011
rect 29444 13961 29496 13977
rect 29526 14079 29578 14091
rect 29526 14045 29536 14079
rect 29570 14045 29578 14079
rect 29526 14011 29578 14045
rect 29526 13977 29536 14011
rect 29570 13977 29578 14011
rect 29526 13961 29578 13977
rect 29683 14075 29735 14091
rect 29683 14041 29691 14075
rect 29725 14041 29735 14075
rect 29683 14007 29735 14041
rect 29683 13973 29691 14007
rect 29725 13973 29735 14007
rect 29683 13961 29735 13973
rect 29765 13961 29819 14091
rect 29849 14075 29901 14091
rect 29849 14041 29859 14075
rect 29893 14041 29901 14075
rect 29849 14007 29901 14041
rect 29849 13973 29859 14007
rect 29893 13973 29901 14007
rect 29849 13961 29901 13973
rect 30002 14079 30054 14091
rect 30002 14045 30010 14079
rect 30044 14045 30054 14079
rect 30002 14011 30054 14045
rect 30002 13977 30010 14011
rect 30044 13977 30054 14011
rect 30002 13961 30054 13977
rect 30084 14079 30136 14091
rect 30084 14045 30094 14079
rect 30128 14045 30136 14079
rect 30084 14011 30136 14045
rect 30084 13977 30094 14011
rect 30128 13977 30136 14011
rect 30084 13961 30136 13977
rect 30242 14057 30294 14091
rect 30242 14023 30250 14057
rect 30284 14023 30294 14057
rect 30242 13961 30294 14023
rect 30324 14045 30376 14091
rect 30527 14079 30579 14091
rect 30527 14045 30535 14079
rect 30569 14045 30579 14079
rect 30324 14027 30391 14045
rect 30324 13993 30334 14027
rect 30368 13993 30391 14027
rect 30324 13961 30391 13993
rect 30421 14033 30473 14045
rect 30421 13999 30431 14033
rect 30465 13999 30473 14033
rect 30421 13961 30473 13999
rect 30527 14011 30579 14045
rect 30527 13977 30535 14011
rect 30569 13977 30579 14011
rect 30527 13961 30579 13977
rect 30609 14046 30661 14091
rect 30609 14012 30619 14046
rect 30653 14012 30661 14046
rect 30609 13961 30661 14012
rect 30715 14023 30767 14045
rect 30715 13989 30723 14023
rect 30757 13989 30767 14023
rect 30715 13961 30767 13989
rect 30797 13961 30858 14045
rect 30888 14003 31007 14045
rect 30888 13969 30941 14003
rect 30975 13969 31007 14003
rect 30888 13961 31007 13969
rect 31037 14033 31087 14045
rect 31257 14033 31311 14089
rect 31037 13961 31103 14033
rect 31133 14007 31212 14033
rect 31133 13973 31153 14007
rect 31187 13973 31212 14007
rect 31133 13961 31212 13973
rect 31242 14003 31311 14033
rect 31242 13969 31263 14003
rect 31297 13969 31311 14003
rect 31242 13961 31311 13969
rect 31341 14045 31391 14089
rect 31341 14007 31443 14045
rect 31341 13973 31375 14007
rect 31409 13973 31443 14007
rect 31341 13961 31443 13973
rect 31473 13961 31515 14045
rect 31545 14033 31663 14045
rect 31822 14033 31872 14045
rect 31545 13961 31681 14033
rect 31711 14009 31777 14033
rect 31711 13975 31721 14009
rect 31755 13975 31777 14009
rect 31711 13961 31777 13975
rect 31807 14009 31872 14033
rect 31807 13975 31828 14009
rect 31862 13975 31872 14009
rect 31807 13961 31872 13975
rect 31902 14003 32007 14045
rect 31902 13969 31961 14003
rect 31995 13969 32007 14003
rect 31902 13961 32007 13969
rect 32075 14033 32127 14045
rect 32075 13999 32083 14033
rect 32117 13999 32127 14033
rect 32075 13961 32127 13999
rect 32157 14007 32211 14045
rect 32157 13973 32167 14007
rect 32201 13973 32211 14007
rect 32157 13961 32211 13973
rect 32241 14033 32293 14045
rect 32241 13999 32251 14033
rect 32285 13999 32293 14033
rect 32241 13961 32293 13999
rect 24238 12842 24296 12854
rect 24238 12666 24250 12842
rect 24284 12666 24296 12842
rect 24238 12654 24296 12666
rect 25096 12842 25154 12854
rect 25096 12666 25108 12842
rect 25142 12666 25154 12842
rect 25096 12654 25154 12666
rect 25954 12842 26012 12854
rect 25954 12666 25966 12842
rect 26000 12666 26012 12842
rect 25954 12654 26012 12666
rect 26812 12842 26870 12854
rect 26812 12666 26824 12842
rect 26858 12666 26870 12842
rect 26812 12654 26870 12666
rect 27670 12842 27728 12854
rect 27670 12666 27682 12842
rect 27716 12666 27728 12842
rect 27670 12654 27728 12666
rect 28528 12842 28586 12854
rect 28528 12666 28540 12842
rect 28574 12666 28586 12842
rect 28528 12654 28586 12666
rect 29386 12842 29444 12854
rect 29386 12666 29398 12842
rect 29432 12666 29444 12842
rect 29386 12654 29444 12666
rect 30244 12842 30302 12854
rect 30244 12666 30256 12842
rect 30290 12666 30302 12842
rect 30244 12654 30302 12666
rect 31102 12842 31160 12854
rect 31102 12666 31114 12842
rect 31148 12666 31160 12842
rect 31102 12654 31160 12666
rect 31960 12842 32018 12854
rect 31960 12666 31972 12842
rect 32006 12666 32018 12842
rect 31960 12654 32018 12666
rect 24238 12260 24296 12272
rect 24238 12084 24250 12260
rect 24284 12084 24296 12260
rect 24238 12072 24296 12084
rect 25096 12260 25154 12272
rect 25096 12084 25108 12260
rect 25142 12084 25154 12260
rect 25096 12072 25154 12084
rect 25954 12260 26012 12272
rect 25954 12084 25966 12260
rect 26000 12084 26012 12260
rect 25954 12072 26012 12084
rect 26812 12260 26870 12272
rect 26812 12084 26824 12260
rect 26858 12084 26870 12260
rect 26812 12072 26870 12084
rect 27670 12260 27728 12272
rect 27670 12084 27682 12260
rect 27716 12084 27728 12260
rect 27670 12072 27728 12084
rect 28528 12260 28586 12272
rect 28528 12084 28540 12260
rect 28574 12084 28586 12260
rect 28528 12072 28586 12084
rect 29386 12260 29444 12272
rect 29386 12084 29398 12260
rect 29432 12084 29444 12260
rect 29386 12072 29444 12084
rect 30244 12260 30302 12272
rect 30244 12084 30256 12260
rect 30290 12084 30302 12260
rect 30244 12072 30302 12084
rect 31102 12260 31160 12272
rect 31102 12084 31114 12260
rect 31148 12084 31160 12260
rect 31102 12072 31160 12084
rect 31960 12260 32018 12272
rect 31960 12084 31972 12260
rect 32006 12084 32018 12260
rect 31960 12072 32018 12084
rect 15156 9656 15214 9668
rect 15156 9480 15168 9656
rect 15202 9480 15214 9656
rect 15156 9468 15214 9480
rect 15614 9656 15672 9668
rect 15614 9480 15626 9656
rect 15660 9480 15672 9656
rect 15614 9468 15672 9480
rect 16072 9656 16130 9668
rect 16072 9480 16084 9656
rect 16118 9480 16130 9656
rect 16072 9468 16130 9480
rect 16530 9656 16588 9668
rect 16530 9480 16542 9656
rect 16576 9480 16588 9656
rect 16530 9468 16588 9480
rect 16988 9656 17046 9668
rect 16988 9480 17000 9656
rect 17034 9480 17046 9656
rect 16988 9468 17046 9480
rect 17446 9656 17504 9668
rect 17446 9480 17458 9656
rect 17492 9480 17504 9656
rect 17446 9468 17504 9480
rect 17904 9656 17962 9668
rect 17904 9480 17916 9656
rect 17950 9480 17962 9656
rect 17904 9468 17962 9480
rect 18362 9656 18420 9668
rect 18362 9480 18374 9656
rect 18408 9480 18420 9656
rect 18362 9468 18420 9480
rect 18820 9656 18878 9668
rect 18820 9480 18832 9656
rect 18866 9480 18878 9656
rect 18820 9468 18878 9480
rect 19278 9656 19336 9668
rect 19278 9480 19290 9656
rect 19324 9480 19336 9656
rect 19278 9468 19336 9480
rect 19736 9656 19794 9668
rect 19736 9480 19748 9656
rect 19782 9480 19794 9656
rect 19736 9468 19794 9480
rect 23918 9656 23976 9668
rect 23918 9480 23930 9656
rect 23964 9480 23976 9656
rect 23918 9468 23976 9480
rect 24376 9656 24434 9668
rect 24376 9480 24388 9656
rect 24422 9480 24434 9656
rect 24376 9468 24434 9480
rect 24834 9656 24892 9668
rect 24834 9480 24846 9656
rect 24880 9480 24892 9656
rect 24834 9468 24892 9480
rect 25292 9656 25350 9668
rect 25292 9480 25304 9656
rect 25338 9480 25350 9656
rect 25292 9468 25350 9480
rect 25750 9656 25808 9668
rect 25750 9480 25762 9656
rect 25796 9480 25808 9656
rect 25750 9468 25808 9480
rect 26208 9656 26266 9668
rect 26208 9480 26220 9656
rect 26254 9480 26266 9656
rect 26208 9468 26266 9480
rect 26666 9656 26724 9668
rect 26666 9480 26678 9656
rect 26712 9480 26724 9656
rect 26666 9468 26724 9480
rect 27124 9656 27182 9668
rect 27124 9480 27136 9656
rect 27170 9480 27182 9656
rect 27124 9468 27182 9480
rect 27582 9656 27640 9668
rect 27582 9480 27594 9656
rect 27628 9480 27640 9656
rect 27582 9468 27640 9480
rect 28040 9656 28098 9668
rect 28040 9480 28052 9656
rect 28086 9480 28098 9656
rect 28040 9468 28098 9480
rect 28498 9656 28556 9668
rect 28498 9480 28510 9656
rect 28544 9480 28556 9656
rect 28498 9468 28556 9480
rect 29144 8851 29196 8867
rect 29144 8817 29152 8851
rect 29186 8817 29196 8851
rect 29144 8783 29196 8817
rect 29144 8749 29152 8783
rect 29186 8749 29196 8783
rect 29144 8737 29196 8749
rect 29226 8851 29278 8867
rect 29226 8817 29236 8851
rect 29270 8817 29278 8851
rect 29226 8783 29278 8817
rect 29226 8749 29236 8783
rect 29270 8749 29278 8783
rect 29226 8737 29278 8749
rect 29389 8855 29441 8867
rect 29389 8821 29397 8855
rect 29431 8821 29441 8855
rect 29389 8737 29441 8821
rect 29471 8847 29525 8867
rect 29471 8813 29481 8847
rect 29515 8813 29525 8847
rect 29471 8737 29525 8813
rect 29555 8855 29609 8867
rect 29555 8821 29565 8855
rect 29599 8821 29609 8855
rect 29555 8737 29609 8821
rect 29639 8847 29693 8867
rect 29639 8813 29649 8847
rect 29683 8813 29693 8847
rect 29639 8737 29693 8813
rect 29723 8854 29775 8867
rect 29723 8820 29733 8854
rect 29767 8820 29775 8854
rect 29723 8737 29775 8820
rect 30579 8535 30631 8547
rect 30579 8501 30587 8535
rect 30621 8501 30631 8535
rect 30579 8463 30631 8501
rect 30661 8509 30715 8547
rect 30661 8475 30671 8509
rect 30705 8475 30715 8509
rect 30661 8463 30715 8475
rect 30745 8535 30797 8547
rect 30745 8501 30755 8535
rect 30789 8501 30797 8535
rect 30745 8463 30797 8501
rect 30851 8509 30903 8547
rect 30851 8475 30859 8509
rect 30893 8475 30903 8509
rect 30851 8463 30903 8475
rect 30933 8535 30983 8547
rect 31282 8547 31332 8591
rect 31163 8535 31213 8547
rect 30933 8523 31015 8535
rect 30933 8489 30944 8523
rect 30978 8489 31015 8523
rect 30933 8463 31015 8489
rect 31045 8523 31114 8535
rect 31045 8489 31055 8523
rect 31089 8489 31114 8523
rect 31045 8463 31114 8489
rect 31144 8463 31213 8535
rect 31243 8517 31332 8547
rect 31243 8483 31254 8517
rect 31288 8483 31332 8517
rect 31243 8463 31332 8483
rect 31362 8535 31412 8591
rect 31772 8578 31824 8593
rect 31584 8535 31634 8547
rect 31362 8523 31433 8535
rect 31362 8489 31373 8523
rect 31407 8489 31433 8523
rect 31362 8463 31433 8489
rect 31463 8523 31539 8535
rect 31463 8489 31476 8523
rect 31510 8489 31539 8523
rect 31463 8463 31539 8489
rect 31569 8463 31634 8535
rect 31664 8523 31716 8547
rect 31664 8489 31674 8523
rect 31708 8489 31716 8523
rect 31664 8463 31716 8489
rect 31772 8544 31780 8578
rect 31814 8544 31824 8578
rect 31772 8510 31824 8544
rect 31772 8476 31780 8510
rect 31814 8476 31824 8510
rect 31772 8463 31824 8476
rect 31854 8539 31908 8593
rect 31854 8505 31864 8539
rect 31898 8505 31908 8539
rect 31854 8463 31908 8505
rect 31938 8580 31990 8593
rect 31938 8546 31948 8580
rect 31982 8546 31990 8580
rect 32141 8547 32191 8593
rect 31938 8512 31990 8546
rect 31938 8478 31948 8512
rect 31982 8478 31990 8512
rect 31938 8463 31990 8478
rect 32044 8535 32096 8547
rect 32044 8501 32052 8535
rect 32086 8501 32096 8535
rect 32044 8463 32096 8501
rect 32126 8509 32191 8547
rect 32126 8475 32147 8509
rect 32181 8475 32191 8509
rect 32126 8463 32191 8475
rect 32221 8547 32273 8593
rect 32221 8513 32231 8547
rect 32265 8513 32273 8547
rect 32221 8463 32273 8513
rect 32368 8581 32420 8593
rect 32368 8547 32376 8581
rect 32410 8547 32420 8581
rect 32368 8513 32420 8547
rect 32368 8479 32376 8513
rect 32410 8479 32420 8513
rect 32368 8463 32420 8479
rect 32450 8581 32502 8593
rect 32450 8547 32460 8581
rect 32494 8547 32502 8581
rect 32450 8513 32502 8547
rect 32450 8479 32460 8513
rect 32494 8479 32502 8513
rect 32450 8463 32502 8479
rect 32613 8509 32665 8593
rect 32613 8475 32621 8509
rect 32655 8475 32665 8509
rect 32613 8463 32665 8475
rect 32695 8517 32749 8593
rect 32695 8483 32705 8517
rect 32739 8483 32749 8517
rect 32695 8463 32749 8483
rect 32779 8509 32833 8593
rect 32779 8475 32789 8509
rect 32823 8475 32833 8509
rect 32779 8463 32833 8475
rect 32863 8517 32917 8593
rect 32863 8483 32873 8517
rect 32907 8483 32917 8517
rect 32863 8463 32917 8483
rect 32947 8510 32999 8593
rect 32947 8476 32957 8510
rect 32991 8476 32999 8510
rect 32947 8463 32999 8476
rect 30579 8331 30631 8369
rect 30579 8297 30587 8331
rect 30621 8297 30631 8331
rect 30579 8285 30631 8297
rect 30661 8357 30715 8369
rect 30661 8323 30671 8357
rect 30705 8323 30715 8357
rect 30661 8285 30715 8323
rect 30745 8331 30797 8369
rect 30745 8297 30755 8331
rect 30789 8297 30797 8331
rect 30745 8285 30797 8297
rect 30851 8357 30903 8369
rect 30851 8323 30859 8357
rect 30893 8323 30903 8357
rect 30851 8285 30903 8323
rect 30933 8343 31015 8369
rect 30933 8309 30944 8343
rect 30978 8309 31015 8343
rect 30933 8297 31015 8309
rect 31045 8343 31114 8369
rect 31045 8309 31055 8343
rect 31089 8309 31114 8343
rect 31045 8297 31114 8309
rect 31144 8297 31213 8369
rect 30933 8285 30983 8297
rect 31163 8285 31213 8297
rect 31243 8349 31332 8369
rect 31243 8315 31254 8349
rect 31288 8315 31332 8349
rect 31243 8285 31332 8315
rect 31282 8241 31332 8285
rect 31362 8343 31433 8369
rect 31362 8309 31373 8343
rect 31407 8309 31433 8343
rect 31362 8297 31433 8309
rect 31463 8343 31539 8369
rect 31463 8309 31476 8343
rect 31510 8309 31539 8343
rect 31463 8297 31539 8309
rect 31569 8297 31634 8369
rect 31362 8241 31412 8297
rect 31584 8285 31634 8297
rect 31664 8343 31716 8369
rect 31664 8309 31674 8343
rect 31708 8309 31716 8343
rect 31664 8285 31716 8309
rect 31772 8356 31824 8369
rect 31772 8322 31780 8356
rect 31814 8322 31824 8356
rect 31772 8288 31824 8322
rect 31772 8254 31780 8288
rect 31814 8254 31824 8288
rect 31772 8239 31824 8254
rect 31854 8327 31908 8369
rect 31854 8293 31864 8327
rect 31898 8293 31908 8327
rect 31854 8239 31908 8293
rect 31938 8354 31990 8369
rect 31938 8320 31948 8354
rect 31982 8320 31990 8354
rect 31938 8286 31990 8320
rect 31938 8252 31948 8286
rect 31982 8252 31990 8286
rect 32044 8331 32096 8369
rect 32044 8297 32052 8331
rect 32086 8297 32096 8331
rect 32044 8285 32096 8297
rect 32126 8357 32191 8369
rect 32126 8323 32147 8357
rect 32181 8323 32191 8357
rect 32126 8285 32191 8323
rect 31938 8239 31990 8252
rect 32141 8239 32191 8285
rect 32221 8319 32273 8369
rect 32221 8285 32231 8319
rect 32265 8285 32273 8319
rect 32221 8239 32273 8285
rect 32368 8353 32420 8369
rect 32368 8319 32376 8353
rect 32410 8319 32420 8353
rect 32368 8285 32420 8319
rect 32368 8251 32376 8285
rect 32410 8251 32420 8285
rect 32368 8239 32420 8251
rect 32450 8353 32502 8369
rect 32450 8319 32460 8353
rect 32494 8319 32502 8353
rect 32450 8285 32502 8319
rect 32450 8251 32460 8285
rect 32494 8251 32502 8285
rect 32450 8239 32502 8251
rect 32613 8357 32665 8369
rect 32613 8323 32621 8357
rect 32655 8323 32665 8357
rect 32613 8239 32665 8323
rect 32695 8349 32749 8369
rect 32695 8315 32705 8349
rect 32739 8315 32749 8349
rect 32695 8239 32749 8315
rect 32779 8357 32833 8369
rect 32779 8323 32789 8357
rect 32823 8323 32833 8357
rect 32779 8239 32833 8323
rect 32863 8349 32917 8369
rect 32863 8315 32873 8349
rect 32907 8315 32917 8349
rect 32863 8239 32917 8315
rect 32947 8356 32999 8369
rect 32947 8322 32957 8356
rect 32991 8322 32999 8356
rect 32947 8239 32999 8322
rect 33277 8331 33329 8369
rect 33277 8297 33285 8331
rect 33319 8297 33329 8331
rect 33277 8285 33329 8297
rect 33359 8357 33413 8369
rect 33359 8323 33369 8357
rect 33403 8323 33413 8357
rect 33359 8285 33413 8323
rect 33443 8331 33495 8369
rect 33443 8297 33453 8331
rect 33487 8297 33495 8331
rect 33443 8285 33495 8297
rect 33549 8357 33601 8369
rect 33549 8323 33557 8357
rect 33591 8323 33601 8357
rect 33549 8285 33601 8323
rect 33631 8343 33713 8369
rect 33631 8309 33642 8343
rect 33676 8309 33713 8343
rect 33631 8297 33713 8309
rect 33743 8343 33812 8369
rect 33743 8309 33753 8343
rect 33787 8309 33812 8343
rect 33743 8297 33812 8309
rect 33842 8297 33911 8369
rect 33631 8285 33681 8297
rect 33861 8285 33911 8297
rect 33941 8349 34030 8369
rect 33941 8315 33952 8349
rect 33986 8315 34030 8349
rect 33941 8285 34030 8315
rect 33980 8241 34030 8285
rect 34060 8343 34131 8369
rect 34060 8309 34071 8343
rect 34105 8309 34131 8343
rect 34060 8297 34131 8309
rect 34161 8343 34237 8369
rect 34161 8309 34174 8343
rect 34208 8309 34237 8343
rect 34161 8297 34237 8309
rect 34267 8297 34332 8369
rect 34060 8241 34110 8297
rect 34282 8285 34332 8297
rect 34362 8343 34414 8369
rect 34362 8309 34372 8343
rect 34406 8309 34414 8343
rect 34362 8285 34414 8309
rect 34470 8356 34522 8369
rect 34470 8322 34478 8356
rect 34512 8322 34522 8356
rect 34470 8288 34522 8322
rect 34470 8254 34478 8288
rect 34512 8254 34522 8288
rect 34470 8239 34522 8254
rect 34552 8327 34606 8369
rect 34552 8293 34562 8327
rect 34596 8293 34606 8327
rect 34552 8239 34606 8293
rect 34636 8354 34688 8369
rect 34636 8320 34646 8354
rect 34680 8320 34688 8354
rect 34636 8286 34688 8320
rect 34636 8252 34646 8286
rect 34680 8252 34688 8286
rect 34742 8331 34794 8369
rect 34742 8297 34750 8331
rect 34784 8297 34794 8331
rect 34742 8285 34794 8297
rect 34824 8357 34889 8369
rect 34824 8323 34845 8357
rect 34879 8323 34889 8357
rect 34824 8285 34889 8323
rect 34636 8239 34688 8252
rect 34839 8239 34889 8285
rect 34919 8319 34971 8369
rect 34919 8285 34929 8319
rect 34963 8285 34971 8319
rect 34919 8239 34971 8285
rect 35066 8353 35118 8369
rect 35066 8319 35074 8353
rect 35108 8319 35118 8353
rect 35066 8285 35118 8319
rect 35066 8251 35074 8285
rect 35108 8251 35118 8285
rect 35066 8239 35118 8251
rect 35148 8353 35200 8369
rect 35148 8319 35158 8353
rect 35192 8319 35200 8353
rect 35148 8285 35200 8319
rect 35148 8251 35158 8285
rect 35192 8251 35200 8285
rect 35148 8239 35200 8251
rect 35311 8357 35363 8369
rect 35311 8323 35319 8357
rect 35353 8323 35363 8357
rect 35311 8239 35363 8323
rect 35393 8349 35447 8369
rect 35393 8315 35403 8349
rect 35437 8315 35447 8349
rect 35393 8239 35447 8315
rect 35477 8357 35531 8369
rect 35477 8323 35487 8357
rect 35521 8323 35531 8357
rect 35477 8239 35531 8323
rect 35561 8349 35615 8369
rect 35561 8315 35571 8349
rect 35605 8315 35615 8349
rect 35561 8239 35615 8315
rect 35645 8356 35697 8369
rect 35645 8322 35655 8356
rect 35689 8322 35697 8356
rect 35645 8239 35697 8322
rect 30579 7447 30631 7459
rect 30579 7413 30587 7447
rect 30621 7413 30631 7447
rect 30579 7375 30631 7413
rect 30661 7421 30715 7459
rect 30661 7387 30671 7421
rect 30705 7387 30715 7421
rect 30661 7375 30715 7387
rect 30745 7447 30797 7459
rect 30745 7413 30755 7447
rect 30789 7413 30797 7447
rect 30745 7375 30797 7413
rect 30851 7421 30903 7459
rect 30851 7387 30859 7421
rect 30893 7387 30903 7421
rect 30851 7375 30903 7387
rect 30933 7447 30983 7459
rect 31282 7459 31332 7503
rect 31163 7447 31213 7459
rect 30933 7435 31015 7447
rect 30933 7401 30944 7435
rect 30978 7401 31015 7435
rect 30933 7375 31015 7401
rect 31045 7435 31114 7447
rect 31045 7401 31055 7435
rect 31089 7401 31114 7435
rect 31045 7375 31114 7401
rect 31144 7375 31213 7447
rect 31243 7429 31332 7459
rect 31243 7395 31254 7429
rect 31288 7395 31332 7429
rect 31243 7375 31332 7395
rect 31362 7447 31412 7503
rect 31772 7490 31824 7505
rect 31584 7447 31634 7459
rect 31362 7435 31433 7447
rect 31362 7401 31373 7435
rect 31407 7401 31433 7435
rect 31362 7375 31433 7401
rect 31463 7435 31539 7447
rect 31463 7401 31476 7435
rect 31510 7401 31539 7435
rect 31463 7375 31539 7401
rect 31569 7375 31634 7447
rect 31664 7435 31716 7459
rect 31664 7401 31674 7435
rect 31708 7401 31716 7435
rect 31664 7375 31716 7401
rect 31772 7456 31780 7490
rect 31814 7456 31824 7490
rect 31772 7422 31824 7456
rect 31772 7388 31780 7422
rect 31814 7388 31824 7422
rect 31772 7375 31824 7388
rect 31854 7451 31908 7505
rect 31854 7417 31864 7451
rect 31898 7417 31908 7451
rect 31854 7375 31908 7417
rect 31938 7492 31990 7505
rect 31938 7458 31948 7492
rect 31982 7458 31990 7492
rect 32141 7459 32191 7505
rect 31938 7424 31990 7458
rect 31938 7390 31948 7424
rect 31982 7390 31990 7424
rect 31938 7375 31990 7390
rect 32044 7447 32096 7459
rect 32044 7413 32052 7447
rect 32086 7413 32096 7447
rect 32044 7375 32096 7413
rect 32126 7421 32191 7459
rect 32126 7387 32147 7421
rect 32181 7387 32191 7421
rect 32126 7375 32191 7387
rect 32221 7459 32273 7505
rect 32221 7425 32231 7459
rect 32265 7425 32273 7459
rect 32221 7375 32273 7425
rect 32368 7493 32420 7505
rect 32368 7459 32376 7493
rect 32410 7459 32420 7493
rect 32368 7425 32420 7459
rect 32368 7391 32376 7425
rect 32410 7391 32420 7425
rect 32368 7375 32420 7391
rect 32450 7493 32502 7505
rect 32450 7459 32460 7493
rect 32494 7459 32502 7493
rect 32450 7425 32502 7459
rect 32450 7391 32460 7425
rect 32494 7391 32502 7425
rect 32450 7375 32502 7391
rect 32613 7421 32665 7505
rect 32613 7387 32621 7421
rect 32655 7387 32665 7421
rect 32613 7375 32665 7387
rect 32695 7429 32749 7505
rect 32695 7395 32705 7429
rect 32739 7395 32749 7429
rect 32695 7375 32749 7395
rect 32779 7421 32833 7505
rect 32779 7387 32789 7421
rect 32823 7387 32833 7421
rect 32779 7375 32833 7387
rect 32863 7429 32917 7505
rect 32863 7395 32873 7429
rect 32907 7395 32917 7429
rect 32863 7375 32917 7395
rect 32947 7422 32999 7505
rect 32947 7388 32957 7422
rect 32991 7388 32999 7422
rect 32947 7375 32999 7388
rect 33277 7447 33329 7459
rect 33277 7413 33285 7447
rect 33319 7413 33329 7447
rect 33277 7375 33329 7413
rect 33359 7421 33413 7459
rect 33359 7387 33369 7421
rect 33403 7387 33413 7421
rect 33359 7375 33413 7387
rect 33443 7447 33495 7459
rect 33443 7413 33453 7447
rect 33487 7413 33495 7447
rect 33443 7375 33495 7413
rect 33549 7421 33601 7459
rect 33549 7387 33557 7421
rect 33591 7387 33601 7421
rect 33549 7375 33601 7387
rect 33631 7447 33681 7459
rect 33980 7459 34030 7503
rect 33861 7447 33911 7459
rect 33631 7435 33713 7447
rect 33631 7401 33642 7435
rect 33676 7401 33713 7435
rect 33631 7375 33713 7401
rect 33743 7435 33812 7447
rect 33743 7401 33753 7435
rect 33787 7401 33812 7435
rect 33743 7375 33812 7401
rect 33842 7375 33911 7447
rect 33941 7429 34030 7459
rect 33941 7395 33952 7429
rect 33986 7395 34030 7429
rect 33941 7375 34030 7395
rect 34060 7447 34110 7503
rect 34470 7490 34522 7505
rect 34282 7447 34332 7459
rect 34060 7435 34131 7447
rect 34060 7401 34071 7435
rect 34105 7401 34131 7435
rect 34060 7375 34131 7401
rect 34161 7435 34237 7447
rect 34161 7401 34174 7435
rect 34208 7401 34237 7435
rect 34161 7375 34237 7401
rect 34267 7375 34332 7447
rect 34362 7435 34414 7459
rect 34362 7401 34372 7435
rect 34406 7401 34414 7435
rect 34362 7375 34414 7401
rect 34470 7456 34478 7490
rect 34512 7456 34522 7490
rect 34470 7422 34522 7456
rect 34470 7388 34478 7422
rect 34512 7388 34522 7422
rect 34470 7375 34522 7388
rect 34552 7451 34606 7505
rect 34552 7417 34562 7451
rect 34596 7417 34606 7451
rect 34552 7375 34606 7417
rect 34636 7492 34688 7505
rect 34636 7458 34646 7492
rect 34680 7458 34688 7492
rect 34839 7459 34889 7505
rect 34636 7424 34688 7458
rect 34636 7390 34646 7424
rect 34680 7390 34688 7424
rect 34636 7375 34688 7390
rect 34742 7447 34794 7459
rect 34742 7413 34750 7447
rect 34784 7413 34794 7447
rect 34742 7375 34794 7413
rect 34824 7421 34889 7459
rect 34824 7387 34845 7421
rect 34879 7387 34889 7421
rect 34824 7375 34889 7387
rect 34919 7459 34971 7505
rect 34919 7425 34929 7459
rect 34963 7425 34971 7459
rect 34919 7375 34971 7425
rect 35066 7493 35118 7505
rect 35066 7459 35074 7493
rect 35108 7459 35118 7493
rect 35066 7425 35118 7459
rect 35066 7391 35074 7425
rect 35108 7391 35118 7425
rect 35066 7375 35118 7391
rect 35148 7493 35200 7505
rect 35148 7459 35158 7493
rect 35192 7459 35200 7493
rect 35148 7425 35200 7459
rect 35148 7391 35158 7425
rect 35192 7391 35200 7425
rect 35148 7375 35200 7391
rect 35311 7421 35363 7505
rect 35311 7387 35319 7421
rect 35353 7387 35363 7421
rect 35311 7375 35363 7387
rect 35393 7429 35447 7505
rect 35393 7395 35403 7429
rect 35437 7395 35447 7429
rect 35393 7375 35447 7395
rect 35477 7421 35531 7505
rect 35477 7387 35487 7421
rect 35521 7387 35531 7421
rect 35477 7375 35531 7387
rect 35561 7429 35615 7505
rect 35561 7395 35571 7429
rect 35605 7395 35615 7429
rect 35561 7375 35615 7395
rect 35645 7422 35697 7505
rect 35645 7388 35655 7422
rect 35689 7388 35697 7422
rect 35645 7375 35697 7388
rect 30579 7243 30631 7281
rect 30579 7209 30587 7243
rect 30621 7209 30631 7243
rect 30579 7197 30631 7209
rect 30661 7269 30715 7281
rect 30661 7235 30671 7269
rect 30705 7235 30715 7269
rect 30661 7197 30715 7235
rect 30745 7243 30797 7281
rect 30745 7209 30755 7243
rect 30789 7209 30797 7243
rect 30745 7197 30797 7209
rect 30851 7269 30903 7281
rect 30851 7235 30859 7269
rect 30893 7235 30903 7269
rect 30851 7197 30903 7235
rect 30933 7255 31015 7281
rect 30933 7221 30944 7255
rect 30978 7221 31015 7255
rect 30933 7209 31015 7221
rect 31045 7255 31114 7281
rect 31045 7221 31055 7255
rect 31089 7221 31114 7255
rect 31045 7209 31114 7221
rect 31144 7209 31213 7281
rect 30933 7197 30983 7209
rect 31163 7197 31213 7209
rect 31243 7261 31332 7281
rect 31243 7227 31254 7261
rect 31288 7227 31332 7261
rect 31243 7197 31332 7227
rect 31282 7153 31332 7197
rect 31362 7255 31433 7281
rect 31362 7221 31373 7255
rect 31407 7221 31433 7255
rect 31362 7209 31433 7221
rect 31463 7255 31539 7281
rect 31463 7221 31476 7255
rect 31510 7221 31539 7255
rect 31463 7209 31539 7221
rect 31569 7209 31634 7281
rect 31362 7153 31412 7209
rect 31584 7197 31634 7209
rect 31664 7255 31716 7281
rect 31664 7221 31674 7255
rect 31708 7221 31716 7255
rect 31664 7197 31716 7221
rect 31772 7268 31824 7281
rect 31772 7234 31780 7268
rect 31814 7234 31824 7268
rect 31772 7200 31824 7234
rect 31772 7166 31780 7200
rect 31814 7166 31824 7200
rect 31772 7151 31824 7166
rect 31854 7239 31908 7281
rect 31854 7205 31864 7239
rect 31898 7205 31908 7239
rect 31854 7151 31908 7205
rect 31938 7266 31990 7281
rect 31938 7232 31948 7266
rect 31982 7232 31990 7266
rect 31938 7198 31990 7232
rect 31938 7164 31948 7198
rect 31982 7164 31990 7198
rect 32044 7243 32096 7281
rect 32044 7209 32052 7243
rect 32086 7209 32096 7243
rect 32044 7197 32096 7209
rect 32126 7269 32191 7281
rect 32126 7235 32147 7269
rect 32181 7235 32191 7269
rect 32126 7197 32191 7235
rect 31938 7151 31990 7164
rect 32141 7151 32191 7197
rect 32221 7231 32273 7281
rect 32221 7197 32231 7231
rect 32265 7197 32273 7231
rect 32221 7151 32273 7197
rect 32368 7265 32420 7281
rect 32368 7231 32376 7265
rect 32410 7231 32420 7265
rect 32368 7197 32420 7231
rect 32368 7163 32376 7197
rect 32410 7163 32420 7197
rect 32368 7151 32420 7163
rect 32450 7265 32502 7281
rect 32450 7231 32460 7265
rect 32494 7231 32502 7265
rect 32450 7197 32502 7231
rect 32450 7163 32460 7197
rect 32494 7163 32502 7197
rect 32450 7151 32502 7163
rect 32613 7269 32665 7281
rect 32613 7235 32621 7269
rect 32655 7235 32665 7269
rect 32613 7151 32665 7235
rect 32695 7261 32749 7281
rect 32695 7227 32705 7261
rect 32739 7227 32749 7261
rect 32695 7151 32749 7227
rect 32779 7269 32833 7281
rect 32779 7235 32789 7269
rect 32823 7235 32833 7269
rect 32779 7151 32833 7235
rect 32863 7261 32917 7281
rect 32863 7227 32873 7261
rect 32907 7227 32917 7261
rect 32863 7151 32917 7227
rect 32947 7268 32999 7281
rect 32947 7234 32957 7268
rect 32991 7234 32999 7268
rect 32947 7151 32999 7234
rect 33277 7243 33329 7281
rect 33277 7209 33285 7243
rect 33319 7209 33329 7243
rect 33277 7197 33329 7209
rect 33359 7269 33413 7281
rect 33359 7235 33369 7269
rect 33403 7235 33413 7269
rect 33359 7197 33413 7235
rect 33443 7243 33495 7281
rect 33443 7209 33453 7243
rect 33487 7209 33495 7243
rect 33443 7197 33495 7209
rect 33549 7269 33601 7281
rect 33549 7235 33557 7269
rect 33591 7235 33601 7269
rect 33549 7197 33601 7235
rect 33631 7255 33713 7281
rect 33631 7221 33642 7255
rect 33676 7221 33713 7255
rect 33631 7209 33713 7221
rect 33743 7255 33812 7281
rect 33743 7221 33753 7255
rect 33787 7221 33812 7255
rect 33743 7209 33812 7221
rect 33842 7209 33911 7281
rect 33631 7197 33681 7209
rect 33861 7197 33911 7209
rect 33941 7261 34030 7281
rect 33941 7227 33952 7261
rect 33986 7227 34030 7261
rect 33941 7197 34030 7227
rect 33980 7153 34030 7197
rect 34060 7255 34131 7281
rect 34060 7221 34071 7255
rect 34105 7221 34131 7255
rect 34060 7209 34131 7221
rect 34161 7255 34237 7281
rect 34161 7221 34174 7255
rect 34208 7221 34237 7255
rect 34161 7209 34237 7221
rect 34267 7209 34332 7281
rect 34060 7153 34110 7209
rect 34282 7197 34332 7209
rect 34362 7255 34414 7281
rect 34362 7221 34372 7255
rect 34406 7221 34414 7255
rect 34362 7197 34414 7221
rect 34470 7268 34522 7281
rect 34470 7234 34478 7268
rect 34512 7234 34522 7268
rect 34470 7200 34522 7234
rect 34470 7166 34478 7200
rect 34512 7166 34522 7200
rect 34470 7151 34522 7166
rect 34552 7239 34606 7281
rect 34552 7205 34562 7239
rect 34596 7205 34606 7239
rect 34552 7151 34606 7205
rect 34636 7266 34688 7281
rect 34636 7232 34646 7266
rect 34680 7232 34688 7266
rect 34636 7198 34688 7232
rect 34636 7164 34646 7198
rect 34680 7164 34688 7198
rect 34742 7243 34794 7281
rect 34742 7209 34750 7243
rect 34784 7209 34794 7243
rect 34742 7197 34794 7209
rect 34824 7269 34889 7281
rect 34824 7235 34845 7269
rect 34879 7235 34889 7269
rect 34824 7197 34889 7235
rect 34636 7151 34688 7164
rect 34839 7151 34889 7197
rect 34919 7231 34971 7281
rect 34919 7197 34929 7231
rect 34963 7197 34971 7231
rect 34919 7151 34971 7197
rect 35066 7265 35118 7281
rect 35066 7231 35074 7265
rect 35108 7231 35118 7265
rect 35066 7197 35118 7231
rect 35066 7163 35074 7197
rect 35108 7163 35118 7197
rect 35066 7151 35118 7163
rect 35148 7265 35200 7281
rect 35148 7231 35158 7265
rect 35192 7231 35200 7265
rect 35148 7197 35200 7231
rect 35148 7163 35158 7197
rect 35192 7163 35200 7197
rect 35148 7151 35200 7163
rect 35311 7269 35363 7281
rect 35311 7235 35319 7269
rect 35353 7235 35363 7269
rect 35311 7151 35363 7235
rect 35393 7261 35447 7281
rect 35393 7227 35403 7261
rect 35437 7227 35447 7261
rect 35393 7151 35447 7227
rect 35477 7269 35531 7281
rect 35477 7235 35487 7269
rect 35521 7235 35531 7269
rect 35477 7151 35531 7235
rect 35561 7261 35615 7281
rect 35561 7227 35571 7261
rect 35605 7227 35615 7261
rect 35561 7151 35615 7227
rect 35645 7268 35697 7281
rect 35645 7234 35655 7268
rect 35689 7234 35697 7268
rect 35645 7151 35697 7234
rect 30579 6359 30631 6371
rect 30579 6325 30587 6359
rect 30621 6325 30631 6359
rect 30579 6287 30631 6325
rect 30661 6333 30715 6371
rect 30661 6299 30671 6333
rect 30705 6299 30715 6333
rect 30661 6287 30715 6299
rect 30745 6359 30797 6371
rect 30745 6325 30755 6359
rect 30789 6325 30797 6359
rect 30745 6287 30797 6325
rect 30851 6333 30903 6371
rect 30851 6299 30859 6333
rect 30893 6299 30903 6333
rect 30851 6287 30903 6299
rect 30933 6359 30983 6371
rect 31282 6371 31332 6415
rect 31163 6359 31213 6371
rect 30933 6347 31015 6359
rect 30933 6313 30944 6347
rect 30978 6313 31015 6347
rect 30933 6287 31015 6313
rect 31045 6347 31114 6359
rect 31045 6313 31055 6347
rect 31089 6313 31114 6347
rect 31045 6287 31114 6313
rect 31144 6287 31213 6359
rect 31243 6341 31332 6371
rect 31243 6307 31254 6341
rect 31288 6307 31332 6341
rect 31243 6287 31332 6307
rect 31362 6359 31412 6415
rect 31772 6402 31824 6417
rect 31584 6359 31634 6371
rect 31362 6347 31433 6359
rect 31362 6313 31373 6347
rect 31407 6313 31433 6347
rect 31362 6287 31433 6313
rect 31463 6347 31539 6359
rect 31463 6313 31476 6347
rect 31510 6313 31539 6347
rect 31463 6287 31539 6313
rect 31569 6287 31634 6359
rect 31664 6347 31716 6371
rect 31664 6313 31674 6347
rect 31708 6313 31716 6347
rect 31664 6287 31716 6313
rect 31772 6368 31780 6402
rect 31814 6368 31824 6402
rect 31772 6334 31824 6368
rect 31772 6300 31780 6334
rect 31814 6300 31824 6334
rect 31772 6287 31824 6300
rect 31854 6363 31908 6417
rect 31854 6329 31864 6363
rect 31898 6329 31908 6363
rect 31854 6287 31908 6329
rect 31938 6404 31990 6417
rect 31938 6370 31948 6404
rect 31982 6370 31990 6404
rect 32141 6371 32191 6417
rect 31938 6336 31990 6370
rect 31938 6302 31948 6336
rect 31982 6302 31990 6336
rect 31938 6287 31990 6302
rect 32044 6359 32096 6371
rect 32044 6325 32052 6359
rect 32086 6325 32096 6359
rect 32044 6287 32096 6325
rect 32126 6333 32191 6371
rect 32126 6299 32147 6333
rect 32181 6299 32191 6333
rect 32126 6287 32191 6299
rect 32221 6371 32273 6417
rect 32221 6337 32231 6371
rect 32265 6337 32273 6371
rect 32221 6287 32273 6337
rect 32368 6405 32420 6417
rect 32368 6371 32376 6405
rect 32410 6371 32420 6405
rect 32368 6337 32420 6371
rect 32368 6303 32376 6337
rect 32410 6303 32420 6337
rect 32368 6287 32420 6303
rect 32450 6405 32502 6417
rect 32450 6371 32460 6405
rect 32494 6371 32502 6405
rect 32450 6337 32502 6371
rect 32450 6303 32460 6337
rect 32494 6303 32502 6337
rect 32450 6287 32502 6303
rect 32613 6333 32665 6417
rect 32613 6299 32621 6333
rect 32655 6299 32665 6333
rect 32613 6287 32665 6299
rect 32695 6341 32749 6417
rect 32695 6307 32705 6341
rect 32739 6307 32749 6341
rect 32695 6287 32749 6307
rect 32779 6333 32833 6417
rect 32779 6299 32789 6333
rect 32823 6299 32833 6333
rect 32779 6287 32833 6299
rect 32863 6341 32917 6417
rect 32863 6307 32873 6341
rect 32907 6307 32917 6341
rect 32863 6287 32917 6307
rect 32947 6334 32999 6417
rect 32947 6300 32957 6334
rect 32991 6300 32999 6334
rect 32947 6287 32999 6300
rect 33277 6359 33329 6371
rect 33277 6325 33285 6359
rect 33319 6325 33329 6359
rect 33277 6287 33329 6325
rect 33359 6333 33413 6371
rect 33359 6299 33369 6333
rect 33403 6299 33413 6333
rect 33359 6287 33413 6299
rect 33443 6359 33495 6371
rect 33443 6325 33453 6359
rect 33487 6325 33495 6359
rect 33443 6287 33495 6325
rect 33549 6333 33601 6371
rect 33549 6299 33557 6333
rect 33591 6299 33601 6333
rect 33549 6287 33601 6299
rect 33631 6359 33681 6371
rect 33980 6371 34030 6415
rect 33861 6359 33911 6371
rect 33631 6347 33713 6359
rect 33631 6313 33642 6347
rect 33676 6313 33713 6347
rect 33631 6287 33713 6313
rect 33743 6347 33812 6359
rect 33743 6313 33753 6347
rect 33787 6313 33812 6347
rect 33743 6287 33812 6313
rect 33842 6287 33911 6359
rect 33941 6341 34030 6371
rect 33941 6307 33952 6341
rect 33986 6307 34030 6341
rect 33941 6287 34030 6307
rect 34060 6359 34110 6415
rect 34470 6402 34522 6417
rect 34282 6359 34332 6371
rect 34060 6347 34131 6359
rect 34060 6313 34071 6347
rect 34105 6313 34131 6347
rect 34060 6287 34131 6313
rect 34161 6347 34237 6359
rect 34161 6313 34174 6347
rect 34208 6313 34237 6347
rect 34161 6287 34237 6313
rect 34267 6287 34332 6359
rect 34362 6347 34414 6371
rect 34362 6313 34372 6347
rect 34406 6313 34414 6347
rect 34362 6287 34414 6313
rect 34470 6368 34478 6402
rect 34512 6368 34522 6402
rect 34470 6334 34522 6368
rect 34470 6300 34478 6334
rect 34512 6300 34522 6334
rect 34470 6287 34522 6300
rect 34552 6363 34606 6417
rect 34552 6329 34562 6363
rect 34596 6329 34606 6363
rect 34552 6287 34606 6329
rect 34636 6404 34688 6417
rect 34636 6370 34646 6404
rect 34680 6370 34688 6404
rect 34839 6371 34889 6417
rect 34636 6336 34688 6370
rect 34636 6302 34646 6336
rect 34680 6302 34688 6336
rect 34636 6287 34688 6302
rect 34742 6359 34794 6371
rect 34742 6325 34750 6359
rect 34784 6325 34794 6359
rect 34742 6287 34794 6325
rect 34824 6333 34889 6371
rect 34824 6299 34845 6333
rect 34879 6299 34889 6333
rect 34824 6287 34889 6299
rect 34919 6371 34971 6417
rect 34919 6337 34929 6371
rect 34963 6337 34971 6371
rect 34919 6287 34971 6337
rect 35066 6405 35118 6417
rect 35066 6371 35074 6405
rect 35108 6371 35118 6405
rect 35066 6337 35118 6371
rect 35066 6303 35074 6337
rect 35108 6303 35118 6337
rect 35066 6287 35118 6303
rect 35148 6405 35200 6417
rect 35148 6371 35158 6405
rect 35192 6371 35200 6405
rect 35148 6337 35200 6371
rect 35148 6303 35158 6337
rect 35192 6303 35200 6337
rect 35148 6287 35200 6303
rect 35311 6333 35363 6417
rect 35311 6299 35319 6333
rect 35353 6299 35363 6333
rect 35311 6287 35363 6299
rect 35393 6341 35447 6417
rect 35393 6307 35403 6341
rect 35437 6307 35447 6341
rect 35393 6287 35447 6307
rect 35477 6333 35531 6417
rect 35477 6299 35487 6333
rect 35521 6299 35531 6333
rect 35477 6287 35531 6299
rect 35561 6341 35615 6417
rect 35561 6307 35571 6341
rect 35605 6307 35615 6341
rect 35561 6287 35615 6307
rect 35645 6334 35697 6417
rect 35645 6300 35655 6334
rect 35689 6300 35697 6334
rect 35645 6287 35697 6300
rect 30579 6155 30631 6193
rect 30579 6121 30587 6155
rect 30621 6121 30631 6155
rect 30579 6109 30631 6121
rect 30661 6181 30715 6193
rect 30661 6147 30671 6181
rect 30705 6147 30715 6181
rect 30661 6109 30715 6147
rect 30745 6155 30797 6193
rect 30745 6121 30755 6155
rect 30789 6121 30797 6155
rect 30745 6109 30797 6121
rect 30851 6181 30903 6193
rect 30851 6147 30859 6181
rect 30893 6147 30903 6181
rect 30851 6109 30903 6147
rect 30933 6167 31015 6193
rect 30933 6133 30944 6167
rect 30978 6133 31015 6167
rect 30933 6121 31015 6133
rect 31045 6167 31114 6193
rect 31045 6133 31055 6167
rect 31089 6133 31114 6167
rect 31045 6121 31114 6133
rect 31144 6121 31213 6193
rect 30933 6109 30983 6121
rect 31163 6109 31213 6121
rect 31243 6173 31332 6193
rect 31243 6139 31254 6173
rect 31288 6139 31332 6173
rect 31243 6109 31332 6139
rect 31282 6065 31332 6109
rect 31362 6167 31433 6193
rect 31362 6133 31373 6167
rect 31407 6133 31433 6167
rect 31362 6121 31433 6133
rect 31463 6167 31539 6193
rect 31463 6133 31476 6167
rect 31510 6133 31539 6167
rect 31463 6121 31539 6133
rect 31569 6121 31634 6193
rect 31362 6065 31412 6121
rect 31584 6109 31634 6121
rect 31664 6167 31716 6193
rect 31664 6133 31674 6167
rect 31708 6133 31716 6167
rect 31664 6109 31716 6133
rect 31772 6180 31824 6193
rect 31772 6146 31780 6180
rect 31814 6146 31824 6180
rect 31772 6112 31824 6146
rect 31772 6078 31780 6112
rect 31814 6078 31824 6112
rect 31772 6063 31824 6078
rect 31854 6151 31908 6193
rect 31854 6117 31864 6151
rect 31898 6117 31908 6151
rect 31854 6063 31908 6117
rect 31938 6178 31990 6193
rect 31938 6144 31948 6178
rect 31982 6144 31990 6178
rect 31938 6110 31990 6144
rect 31938 6076 31948 6110
rect 31982 6076 31990 6110
rect 32044 6155 32096 6193
rect 32044 6121 32052 6155
rect 32086 6121 32096 6155
rect 32044 6109 32096 6121
rect 32126 6181 32191 6193
rect 32126 6147 32147 6181
rect 32181 6147 32191 6181
rect 32126 6109 32191 6147
rect 31938 6063 31990 6076
rect 32141 6063 32191 6109
rect 32221 6143 32273 6193
rect 32221 6109 32231 6143
rect 32265 6109 32273 6143
rect 32221 6063 32273 6109
rect 32368 6177 32420 6193
rect 32368 6143 32376 6177
rect 32410 6143 32420 6177
rect 32368 6109 32420 6143
rect 32368 6075 32376 6109
rect 32410 6075 32420 6109
rect 32368 6063 32420 6075
rect 32450 6177 32502 6193
rect 32450 6143 32460 6177
rect 32494 6143 32502 6177
rect 32450 6109 32502 6143
rect 32450 6075 32460 6109
rect 32494 6075 32502 6109
rect 32450 6063 32502 6075
rect 32613 6181 32665 6193
rect 32613 6147 32621 6181
rect 32655 6147 32665 6181
rect 32613 6063 32665 6147
rect 32695 6173 32749 6193
rect 32695 6139 32705 6173
rect 32739 6139 32749 6173
rect 32695 6063 32749 6139
rect 32779 6181 32833 6193
rect 32779 6147 32789 6181
rect 32823 6147 32833 6181
rect 32779 6063 32833 6147
rect 32863 6173 32917 6193
rect 32863 6139 32873 6173
rect 32907 6139 32917 6173
rect 32863 6063 32917 6139
rect 32947 6180 32999 6193
rect 32947 6146 32957 6180
rect 32991 6146 32999 6180
rect 32947 6063 32999 6146
rect 33277 6155 33329 6193
rect 33277 6121 33285 6155
rect 33319 6121 33329 6155
rect 33277 6109 33329 6121
rect 33359 6181 33413 6193
rect 33359 6147 33369 6181
rect 33403 6147 33413 6181
rect 33359 6109 33413 6147
rect 33443 6155 33495 6193
rect 33443 6121 33453 6155
rect 33487 6121 33495 6155
rect 33443 6109 33495 6121
rect 33549 6181 33601 6193
rect 33549 6147 33557 6181
rect 33591 6147 33601 6181
rect 33549 6109 33601 6147
rect 33631 6167 33713 6193
rect 33631 6133 33642 6167
rect 33676 6133 33713 6167
rect 33631 6121 33713 6133
rect 33743 6167 33812 6193
rect 33743 6133 33753 6167
rect 33787 6133 33812 6167
rect 33743 6121 33812 6133
rect 33842 6121 33911 6193
rect 33631 6109 33681 6121
rect 33861 6109 33911 6121
rect 33941 6173 34030 6193
rect 33941 6139 33952 6173
rect 33986 6139 34030 6173
rect 33941 6109 34030 6139
rect 33980 6065 34030 6109
rect 34060 6167 34131 6193
rect 34060 6133 34071 6167
rect 34105 6133 34131 6167
rect 34060 6121 34131 6133
rect 34161 6167 34237 6193
rect 34161 6133 34174 6167
rect 34208 6133 34237 6167
rect 34161 6121 34237 6133
rect 34267 6121 34332 6193
rect 34060 6065 34110 6121
rect 34282 6109 34332 6121
rect 34362 6167 34414 6193
rect 34362 6133 34372 6167
rect 34406 6133 34414 6167
rect 34362 6109 34414 6133
rect 34470 6180 34522 6193
rect 34470 6146 34478 6180
rect 34512 6146 34522 6180
rect 34470 6112 34522 6146
rect 34470 6078 34478 6112
rect 34512 6078 34522 6112
rect 34470 6063 34522 6078
rect 34552 6151 34606 6193
rect 34552 6117 34562 6151
rect 34596 6117 34606 6151
rect 34552 6063 34606 6117
rect 34636 6178 34688 6193
rect 34636 6144 34646 6178
rect 34680 6144 34688 6178
rect 34636 6110 34688 6144
rect 34636 6076 34646 6110
rect 34680 6076 34688 6110
rect 34742 6155 34794 6193
rect 34742 6121 34750 6155
rect 34784 6121 34794 6155
rect 34742 6109 34794 6121
rect 34824 6181 34889 6193
rect 34824 6147 34845 6181
rect 34879 6147 34889 6181
rect 34824 6109 34889 6147
rect 34636 6063 34688 6076
rect 34839 6063 34889 6109
rect 34919 6143 34971 6193
rect 34919 6109 34929 6143
rect 34963 6109 34971 6143
rect 34919 6063 34971 6109
rect 35066 6177 35118 6193
rect 35066 6143 35074 6177
rect 35108 6143 35118 6177
rect 35066 6109 35118 6143
rect 35066 6075 35074 6109
rect 35108 6075 35118 6109
rect 35066 6063 35118 6075
rect 35148 6177 35200 6193
rect 35148 6143 35158 6177
rect 35192 6143 35200 6177
rect 35148 6109 35200 6143
rect 35148 6075 35158 6109
rect 35192 6075 35200 6109
rect 35148 6063 35200 6075
rect 35311 6181 35363 6193
rect 35311 6147 35319 6181
rect 35353 6147 35363 6181
rect 35311 6063 35363 6147
rect 35393 6173 35447 6193
rect 35393 6139 35403 6173
rect 35437 6139 35447 6173
rect 35393 6063 35447 6139
rect 35477 6181 35531 6193
rect 35477 6147 35487 6181
rect 35521 6147 35531 6181
rect 35477 6063 35531 6147
rect 35561 6173 35615 6193
rect 35561 6139 35571 6173
rect 35605 6139 35615 6173
rect 35561 6063 35615 6139
rect 35645 6180 35697 6193
rect 35645 6146 35655 6180
rect 35689 6146 35697 6180
rect 35645 6063 35697 6146
rect 8766 -2226 8824 -2214
rect 8766 -2402 8778 -2226
rect 8812 -2402 8824 -2226
rect 8766 -2414 8824 -2402
rect 9224 -2226 9282 -2214
rect 9224 -2402 9236 -2226
rect 9270 -2402 9282 -2226
rect 9224 -2414 9282 -2402
rect 9682 -2226 9740 -2214
rect 9682 -2402 9694 -2226
rect 9728 -2402 9740 -2226
rect 9682 -2414 9740 -2402
rect 10140 -2226 10198 -2214
rect 10140 -2402 10152 -2226
rect 10186 -2402 10198 -2226
rect 10140 -2414 10198 -2402
rect 10598 -2226 10656 -2214
rect 10598 -2402 10610 -2226
rect 10644 -2402 10656 -2226
rect 10598 -2414 10656 -2402
rect 11056 -2226 11114 -2214
rect 11056 -2402 11068 -2226
rect 11102 -2402 11114 -2226
rect 11056 -2414 11114 -2402
rect 11514 -2226 11572 -2214
rect 11514 -2402 11526 -2226
rect 11560 -2402 11572 -2226
rect 11514 -2414 11572 -2402
rect 11972 -2226 12030 -2214
rect 11972 -2402 11984 -2226
rect 12018 -2402 12030 -2226
rect 11972 -2414 12030 -2402
rect 12430 -2226 12488 -2214
rect 12430 -2402 12442 -2226
rect 12476 -2402 12488 -2226
rect 12430 -2414 12488 -2402
rect 12888 -2226 12946 -2214
rect 12888 -2402 12900 -2226
rect 12934 -2402 12946 -2226
rect 12888 -2414 12946 -2402
rect 13346 -2226 13404 -2214
rect 13346 -2402 13358 -2226
rect 13392 -2402 13404 -2226
rect 13346 -2414 13404 -2402
rect 13766 -2226 13824 -2214
rect 13766 -2402 13778 -2226
rect 13812 -2402 13824 -2226
rect 13766 -2414 13824 -2402
rect 14224 -2226 14282 -2214
rect 14224 -2402 14236 -2226
rect 14270 -2402 14282 -2226
rect 14224 -2414 14282 -2402
rect 14682 -2226 14740 -2214
rect 14682 -2402 14694 -2226
rect 14728 -2402 14740 -2226
rect 14682 -2414 14740 -2402
rect 15140 -2226 15198 -2214
rect 15140 -2402 15152 -2226
rect 15186 -2402 15198 -2226
rect 15140 -2414 15198 -2402
rect 15598 -2226 15656 -2214
rect 15598 -2402 15610 -2226
rect 15644 -2402 15656 -2226
rect 15598 -2414 15656 -2402
rect 16056 -2226 16114 -2214
rect 16056 -2402 16068 -2226
rect 16102 -2402 16114 -2226
rect 16056 -2414 16114 -2402
rect 16514 -2226 16572 -2214
rect 16514 -2402 16526 -2226
rect 16560 -2402 16572 -2226
rect 16514 -2414 16572 -2402
rect 16972 -2226 17030 -2214
rect 16972 -2402 16984 -2226
rect 17018 -2402 17030 -2226
rect 16972 -2414 17030 -2402
rect 17430 -2226 17488 -2214
rect 17430 -2402 17442 -2226
rect 17476 -2402 17488 -2226
rect 17430 -2414 17488 -2402
rect 17888 -2226 17946 -2214
rect 17888 -2402 17900 -2226
rect 17934 -2402 17946 -2226
rect 17888 -2414 17946 -2402
rect 18346 -2226 18404 -2214
rect 18346 -2402 18358 -2226
rect 18392 -2402 18404 -2226
rect 18346 -2414 18404 -2402
rect 8766 -2894 8824 -2882
rect 8766 -3070 8778 -2894
rect 8812 -3070 8824 -2894
rect 8766 -3082 8824 -3070
rect 9224 -2894 9282 -2882
rect 9224 -3070 9236 -2894
rect 9270 -3070 9282 -2894
rect 9224 -3082 9282 -3070
rect 9682 -2894 9740 -2882
rect 9682 -3070 9694 -2894
rect 9728 -3070 9740 -2894
rect 9682 -3082 9740 -3070
rect 10140 -2894 10198 -2882
rect 10140 -3070 10152 -2894
rect 10186 -3070 10198 -2894
rect 10140 -3082 10198 -3070
rect 10598 -2894 10656 -2882
rect 10598 -3070 10610 -2894
rect 10644 -3070 10656 -2894
rect 10598 -3082 10656 -3070
rect 11056 -2894 11114 -2882
rect 11056 -3070 11068 -2894
rect 11102 -3070 11114 -2894
rect 11056 -3082 11114 -3070
rect 11514 -2894 11572 -2882
rect 11514 -3070 11526 -2894
rect 11560 -3070 11572 -2894
rect 11514 -3082 11572 -3070
rect 11972 -2894 12030 -2882
rect 11972 -3070 11984 -2894
rect 12018 -3070 12030 -2894
rect 11972 -3082 12030 -3070
rect 12430 -2894 12488 -2882
rect 12430 -3070 12442 -2894
rect 12476 -3070 12488 -2894
rect 12430 -3082 12488 -3070
rect 12888 -2894 12946 -2882
rect 12888 -3070 12900 -2894
rect 12934 -3070 12946 -2894
rect 12888 -3082 12946 -3070
rect 13346 -2894 13404 -2882
rect 13346 -3070 13358 -2894
rect 13392 -3070 13404 -2894
rect 13346 -3082 13404 -3070
rect 23766 -2226 23824 -2214
rect 23766 -2402 23778 -2226
rect 23812 -2402 23824 -2226
rect 23766 -2414 23824 -2402
rect 24224 -2226 24282 -2214
rect 24224 -2402 24236 -2226
rect 24270 -2402 24282 -2226
rect 24224 -2414 24282 -2402
rect 24682 -2226 24740 -2214
rect 24682 -2402 24694 -2226
rect 24728 -2402 24740 -2226
rect 24682 -2414 24740 -2402
rect 25140 -2226 25198 -2214
rect 25140 -2402 25152 -2226
rect 25186 -2402 25198 -2226
rect 25140 -2414 25198 -2402
rect 25598 -2226 25656 -2214
rect 25598 -2402 25610 -2226
rect 25644 -2402 25656 -2226
rect 25598 -2414 25656 -2402
rect 26056 -2226 26114 -2214
rect 26056 -2402 26068 -2226
rect 26102 -2402 26114 -2226
rect 26056 -2414 26114 -2402
rect 26514 -2226 26572 -2214
rect 26514 -2402 26526 -2226
rect 26560 -2402 26572 -2226
rect 26514 -2414 26572 -2402
rect 26972 -2226 27030 -2214
rect 26972 -2402 26984 -2226
rect 27018 -2402 27030 -2226
rect 26972 -2414 27030 -2402
rect 27430 -2226 27488 -2214
rect 27430 -2402 27442 -2226
rect 27476 -2402 27488 -2226
rect 27430 -2414 27488 -2402
rect 27888 -2226 27946 -2214
rect 27888 -2402 27900 -2226
rect 27934 -2402 27946 -2226
rect 27888 -2414 27946 -2402
rect 28346 -2226 28404 -2214
rect 28346 -2402 28358 -2226
rect 28392 -2402 28404 -2226
rect 28346 -2414 28404 -2402
rect 28766 -2226 28824 -2214
rect 28766 -2402 28778 -2226
rect 28812 -2402 28824 -2226
rect 28766 -2414 28824 -2402
rect 29224 -2226 29282 -2214
rect 29224 -2402 29236 -2226
rect 29270 -2402 29282 -2226
rect 29224 -2414 29282 -2402
rect 29682 -2226 29740 -2214
rect 29682 -2402 29694 -2226
rect 29728 -2402 29740 -2226
rect 29682 -2414 29740 -2402
rect 30140 -2226 30198 -2214
rect 30140 -2402 30152 -2226
rect 30186 -2402 30198 -2226
rect 30140 -2414 30198 -2402
rect 30598 -2226 30656 -2214
rect 30598 -2402 30610 -2226
rect 30644 -2402 30656 -2226
rect 30598 -2414 30656 -2402
rect 31056 -2226 31114 -2214
rect 31056 -2402 31068 -2226
rect 31102 -2402 31114 -2226
rect 31056 -2414 31114 -2402
rect 31514 -2226 31572 -2214
rect 31514 -2402 31526 -2226
rect 31560 -2402 31572 -2226
rect 31514 -2414 31572 -2402
rect 31972 -2226 32030 -2214
rect 31972 -2402 31984 -2226
rect 32018 -2402 32030 -2226
rect 31972 -2414 32030 -2402
rect 32430 -2226 32488 -2214
rect 32430 -2402 32442 -2226
rect 32476 -2402 32488 -2226
rect 32430 -2414 32488 -2402
rect 32888 -2226 32946 -2214
rect 32888 -2402 32900 -2226
rect 32934 -2402 32946 -2226
rect 32888 -2414 32946 -2402
rect 33346 -2226 33404 -2214
rect 33346 -2402 33358 -2226
rect 33392 -2402 33404 -2226
rect 33346 -2414 33404 -2402
rect 23766 -2894 23824 -2882
rect 23766 -3070 23778 -2894
rect 23812 -3070 23824 -2894
rect 23766 -3082 23824 -3070
rect 24224 -2894 24282 -2882
rect 24224 -3070 24236 -2894
rect 24270 -3070 24282 -2894
rect 24224 -3082 24282 -3070
rect 24682 -2894 24740 -2882
rect 24682 -3070 24694 -2894
rect 24728 -3070 24740 -2894
rect 24682 -3082 24740 -3070
rect 25140 -2894 25198 -2882
rect 25140 -3070 25152 -2894
rect 25186 -3070 25198 -2894
rect 25140 -3082 25198 -3070
rect 25598 -2894 25656 -2882
rect 25598 -3070 25610 -2894
rect 25644 -3070 25656 -2894
rect 25598 -3082 25656 -3070
rect 26056 -2894 26114 -2882
rect 26056 -3070 26068 -2894
rect 26102 -3070 26114 -2894
rect 26056 -3082 26114 -3070
rect 26514 -2894 26572 -2882
rect 26514 -3070 26526 -2894
rect 26560 -3070 26572 -2894
rect 26514 -3082 26572 -3070
rect 26972 -2894 27030 -2882
rect 26972 -3070 26984 -2894
rect 27018 -3070 27030 -2894
rect 26972 -3082 27030 -3070
rect 27430 -2894 27488 -2882
rect 27430 -3070 27442 -2894
rect 27476 -3070 27488 -2894
rect 27430 -3082 27488 -3070
rect 27888 -2894 27946 -2882
rect 27888 -3070 27900 -2894
rect 27934 -3070 27946 -2894
rect 27888 -3082 27946 -3070
rect 28346 -2894 28404 -2882
rect 28346 -3070 28358 -2894
rect 28392 -3070 28404 -2894
rect 28346 -3082 28404 -3070
rect 17698 -5686 17756 -5674
rect 17698 -5862 17710 -5686
rect 17744 -5862 17756 -5686
rect 17698 -5874 17756 -5862
rect 18156 -5686 18214 -5674
rect 18156 -5862 18168 -5686
rect 18202 -5862 18214 -5686
rect 18156 -5874 18214 -5862
rect 18614 -5686 18672 -5674
rect 18614 -5862 18626 -5686
rect 18660 -5862 18672 -5686
rect 18614 -5874 18672 -5862
rect 19072 -5686 19130 -5674
rect 19072 -5862 19084 -5686
rect 19118 -5862 19130 -5686
rect 19072 -5874 19130 -5862
rect 19530 -5686 19588 -5674
rect 19530 -5862 19542 -5686
rect 19576 -5862 19588 -5686
rect 19530 -5874 19588 -5862
rect 19988 -5686 20046 -5674
rect 19988 -5862 20000 -5686
rect 20034 -5862 20046 -5686
rect 19988 -5874 20046 -5862
rect 20446 -5686 20504 -5674
rect 20446 -5862 20458 -5686
rect 20492 -5862 20504 -5686
rect 20446 -5874 20504 -5862
rect 20904 -5686 20962 -5674
rect 20904 -5862 20916 -5686
rect 20950 -5862 20962 -5686
rect 20904 -5874 20962 -5862
rect 21362 -5686 21420 -5674
rect 21362 -5862 21374 -5686
rect 21408 -5862 21420 -5686
rect 21362 -5874 21420 -5862
rect 21820 -5686 21878 -5674
rect 21820 -5862 21832 -5686
rect 21866 -5862 21878 -5686
rect 21820 -5874 21878 -5862
rect 22278 -5686 22336 -5674
rect 22278 -5862 22290 -5686
rect 22324 -5862 22336 -5686
rect 22278 -5874 22336 -5862
rect 12698 -6354 12756 -6342
rect 12698 -6530 12710 -6354
rect 12744 -6530 12756 -6354
rect 12698 -6542 12756 -6530
rect 13156 -6354 13214 -6342
rect 13156 -6530 13168 -6354
rect 13202 -6530 13214 -6354
rect 13156 -6542 13214 -6530
rect 13614 -6354 13672 -6342
rect 13614 -6530 13626 -6354
rect 13660 -6530 13672 -6354
rect 13614 -6542 13672 -6530
rect 14072 -6354 14130 -6342
rect 14072 -6530 14084 -6354
rect 14118 -6530 14130 -6354
rect 14072 -6542 14130 -6530
rect 14530 -6354 14588 -6342
rect 14530 -6530 14542 -6354
rect 14576 -6530 14588 -6354
rect 14530 -6542 14588 -6530
rect 14988 -6354 15046 -6342
rect 14988 -6530 15000 -6354
rect 15034 -6530 15046 -6354
rect 14988 -6542 15046 -6530
rect 15446 -6354 15504 -6342
rect 15446 -6530 15458 -6354
rect 15492 -6530 15504 -6354
rect 15446 -6542 15504 -6530
rect 15904 -6354 15962 -6342
rect 15904 -6530 15916 -6354
rect 15950 -6530 15962 -6354
rect 15904 -6542 15962 -6530
rect 16362 -6354 16420 -6342
rect 16362 -6530 16374 -6354
rect 16408 -6530 16420 -6354
rect 16362 -6542 16420 -6530
rect 16820 -6354 16878 -6342
rect 16820 -6530 16832 -6354
rect 16866 -6530 16878 -6354
rect 16820 -6542 16878 -6530
rect 17278 -6354 17336 -6342
rect 17278 -6530 17290 -6354
rect 17324 -6530 17336 -6354
rect 17278 -6542 17336 -6530
rect 17698 -6354 17756 -6342
rect 17698 -6530 17710 -6354
rect 17744 -6530 17756 -6354
rect 17698 -6542 17756 -6530
rect 18156 -6354 18214 -6342
rect 18156 -6530 18168 -6354
rect 18202 -6530 18214 -6354
rect 18156 -6542 18214 -6530
rect 18614 -6354 18672 -6342
rect 18614 -6530 18626 -6354
rect 18660 -6530 18672 -6354
rect 18614 -6542 18672 -6530
rect 19072 -6354 19130 -6342
rect 19072 -6530 19084 -6354
rect 19118 -6530 19130 -6354
rect 19072 -6542 19130 -6530
rect 19530 -6354 19588 -6342
rect 19530 -6530 19542 -6354
rect 19576 -6530 19588 -6354
rect 19530 -6542 19588 -6530
rect 19988 -6354 20046 -6342
rect 19988 -6530 20000 -6354
rect 20034 -6530 20046 -6354
rect 19988 -6542 20046 -6530
rect 20446 -6354 20504 -6342
rect 20446 -6530 20458 -6354
rect 20492 -6530 20504 -6354
rect 20446 -6542 20504 -6530
rect 20904 -6354 20962 -6342
rect 20904 -6530 20916 -6354
rect 20950 -6530 20962 -6354
rect 20904 -6542 20962 -6530
rect 21362 -6354 21420 -6342
rect 21362 -6530 21374 -6354
rect 21408 -6530 21420 -6354
rect 21362 -6542 21420 -6530
rect 21820 -6354 21878 -6342
rect 21820 -6530 21832 -6354
rect 21866 -6530 21878 -6354
rect 21820 -6542 21878 -6530
rect 22278 -6354 22336 -6342
rect 22278 -6530 22290 -6354
rect 22324 -6530 22336 -6354
rect 22278 -6542 22336 -6530
rect 32698 -5686 32756 -5674
rect 32698 -5862 32710 -5686
rect 32744 -5862 32756 -5686
rect 32698 -5874 32756 -5862
rect 33156 -5686 33214 -5674
rect 33156 -5862 33168 -5686
rect 33202 -5862 33214 -5686
rect 33156 -5874 33214 -5862
rect 33614 -5686 33672 -5674
rect 33614 -5862 33626 -5686
rect 33660 -5862 33672 -5686
rect 33614 -5874 33672 -5862
rect 34072 -5686 34130 -5674
rect 34072 -5862 34084 -5686
rect 34118 -5862 34130 -5686
rect 34072 -5874 34130 -5862
rect 34530 -5686 34588 -5674
rect 34530 -5862 34542 -5686
rect 34576 -5862 34588 -5686
rect 34530 -5874 34588 -5862
rect 34988 -5686 35046 -5674
rect 34988 -5862 35000 -5686
rect 35034 -5862 35046 -5686
rect 34988 -5874 35046 -5862
rect 35446 -5686 35504 -5674
rect 35446 -5862 35458 -5686
rect 35492 -5862 35504 -5686
rect 35446 -5874 35504 -5862
rect 35904 -5686 35962 -5674
rect 35904 -5862 35916 -5686
rect 35950 -5862 35962 -5686
rect 35904 -5874 35962 -5862
rect 36362 -5686 36420 -5674
rect 36362 -5862 36374 -5686
rect 36408 -5862 36420 -5686
rect 36362 -5874 36420 -5862
rect 36820 -5686 36878 -5674
rect 36820 -5862 36832 -5686
rect 36866 -5862 36878 -5686
rect 36820 -5874 36878 -5862
rect 37278 -5686 37336 -5674
rect 37278 -5862 37290 -5686
rect 37324 -5862 37336 -5686
rect 37278 -5874 37336 -5862
rect 27698 -6354 27756 -6342
rect 27698 -6530 27710 -6354
rect 27744 -6530 27756 -6354
rect 27698 -6542 27756 -6530
rect 28156 -6354 28214 -6342
rect 28156 -6530 28168 -6354
rect 28202 -6530 28214 -6354
rect 28156 -6542 28214 -6530
rect 28614 -6354 28672 -6342
rect 28614 -6530 28626 -6354
rect 28660 -6530 28672 -6354
rect 28614 -6542 28672 -6530
rect 29072 -6354 29130 -6342
rect 29072 -6530 29084 -6354
rect 29118 -6530 29130 -6354
rect 29072 -6542 29130 -6530
rect 29530 -6354 29588 -6342
rect 29530 -6530 29542 -6354
rect 29576 -6530 29588 -6354
rect 29530 -6542 29588 -6530
rect 29988 -6354 30046 -6342
rect 29988 -6530 30000 -6354
rect 30034 -6530 30046 -6354
rect 29988 -6542 30046 -6530
rect 30446 -6354 30504 -6342
rect 30446 -6530 30458 -6354
rect 30492 -6530 30504 -6354
rect 30446 -6542 30504 -6530
rect 30904 -6354 30962 -6342
rect 30904 -6530 30916 -6354
rect 30950 -6530 30962 -6354
rect 30904 -6542 30962 -6530
rect 31362 -6354 31420 -6342
rect 31362 -6530 31374 -6354
rect 31408 -6530 31420 -6354
rect 31362 -6542 31420 -6530
rect 31820 -6354 31878 -6342
rect 31820 -6530 31832 -6354
rect 31866 -6530 31878 -6354
rect 31820 -6542 31878 -6530
rect 32278 -6354 32336 -6342
rect 32278 -6530 32290 -6354
rect 32324 -6530 32336 -6354
rect 32278 -6542 32336 -6530
rect 32698 -6354 32756 -6342
rect 32698 -6530 32710 -6354
rect 32744 -6530 32756 -6354
rect 32698 -6542 32756 -6530
rect 33156 -6354 33214 -6342
rect 33156 -6530 33168 -6354
rect 33202 -6530 33214 -6354
rect 33156 -6542 33214 -6530
rect 33614 -6354 33672 -6342
rect 33614 -6530 33626 -6354
rect 33660 -6530 33672 -6354
rect 33614 -6542 33672 -6530
rect 34072 -6354 34130 -6342
rect 34072 -6530 34084 -6354
rect 34118 -6530 34130 -6354
rect 34072 -6542 34130 -6530
rect 34530 -6354 34588 -6342
rect 34530 -6530 34542 -6354
rect 34576 -6530 34588 -6354
rect 34530 -6542 34588 -6530
rect 34988 -6354 35046 -6342
rect 34988 -6530 35000 -6354
rect 35034 -6530 35046 -6354
rect 34988 -6542 35046 -6530
rect 35446 -6354 35504 -6342
rect 35446 -6530 35458 -6354
rect 35492 -6530 35504 -6354
rect 35446 -6542 35504 -6530
rect 35904 -6354 35962 -6342
rect 35904 -6530 35916 -6354
rect 35950 -6530 35962 -6354
rect 35904 -6542 35962 -6530
rect 36362 -6354 36420 -6342
rect 36362 -6530 36374 -6354
rect 36408 -6530 36420 -6354
rect 36362 -6542 36420 -6530
rect 36820 -6354 36878 -6342
rect 36820 -6530 36832 -6354
rect 36866 -6530 36878 -6354
rect 36820 -6542 36878 -6530
rect 37278 -6354 37336 -6342
rect 37278 -6530 37290 -6354
rect 37324 -6530 37336 -6354
rect 37278 -6542 37336 -6530
rect 8766 -20226 8824 -20214
rect 8766 -20402 8778 -20226
rect 8812 -20402 8824 -20226
rect 8766 -20414 8824 -20402
rect 9224 -20226 9282 -20214
rect 9224 -20402 9236 -20226
rect 9270 -20402 9282 -20226
rect 9224 -20414 9282 -20402
rect 9682 -20226 9740 -20214
rect 9682 -20402 9694 -20226
rect 9728 -20402 9740 -20226
rect 9682 -20414 9740 -20402
rect 10140 -20226 10198 -20214
rect 10140 -20402 10152 -20226
rect 10186 -20402 10198 -20226
rect 10140 -20414 10198 -20402
rect 10598 -20226 10656 -20214
rect 10598 -20402 10610 -20226
rect 10644 -20402 10656 -20226
rect 10598 -20414 10656 -20402
rect 11056 -20226 11114 -20214
rect 11056 -20402 11068 -20226
rect 11102 -20402 11114 -20226
rect 11056 -20414 11114 -20402
rect 11514 -20226 11572 -20214
rect 11514 -20402 11526 -20226
rect 11560 -20402 11572 -20226
rect 11514 -20414 11572 -20402
rect 11972 -20226 12030 -20214
rect 11972 -20402 11984 -20226
rect 12018 -20402 12030 -20226
rect 11972 -20414 12030 -20402
rect 12430 -20226 12488 -20214
rect 12430 -20402 12442 -20226
rect 12476 -20402 12488 -20226
rect 12430 -20414 12488 -20402
rect 12888 -20226 12946 -20214
rect 12888 -20402 12900 -20226
rect 12934 -20402 12946 -20226
rect 12888 -20414 12946 -20402
rect 13346 -20226 13404 -20214
rect 13346 -20402 13358 -20226
rect 13392 -20402 13404 -20226
rect 13346 -20414 13404 -20402
rect 13766 -20226 13824 -20214
rect 13766 -20402 13778 -20226
rect 13812 -20402 13824 -20226
rect 13766 -20414 13824 -20402
rect 14224 -20226 14282 -20214
rect 14224 -20402 14236 -20226
rect 14270 -20402 14282 -20226
rect 14224 -20414 14282 -20402
rect 14682 -20226 14740 -20214
rect 14682 -20402 14694 -20226
rect 14728 -20402 14740 -20226
rect 14682 -20414 14740 -20402
rect 15140 -20226 15198 -20214
rect 15140 -20402 15152 -20226
rect 15186 -20402 15198 -20226
rect 15140 -20414 15198 -20402
rect 15598 -20226 15656 -20214
rect 15598 -20402 15610 -20226
rect 15644 -20402 15656 -20226
rect 15598 -20414 15656 -20402
rect 16056 -20226 16114 -20214
rect 16056 -20402 16068 -20226
rect 16102 -20402 16114 -20226
rect 16056 -20414 16114 -20402
rect 16514 -20226 16572 -20214
rect 16514 -20402 16526 -20226
rect 16560 -20402 16572 -20226
rect 16514 -20414 16572 -20402
rect 16972 -20226 17030 -20214
rect 16972 -20402 16984 -20226
rect 17018 -20402 17030 -20226
rect 16972 -20414 17030 -20402
rect 17430 -20226 17488 -20214
rect 17430 -20402 17442 -20226
rect 17476 -20402 17488 -20226
rect 17430 -20414 17488 -20402
rect 17888 -20226 17946 -20214
rect 17888 -20402 17900 -20226
rect 17934 -20402 17946 -20226
rect 17888 -20414 17946 -20402
rect 18346 -20226 18404 -20214
rect 18346 -20402 18358 -20226
rect 18392 -20402 18404 -20226
rect 18346 -20414 18404 -20402
rect 8766 -20894 8824 -20882
rect 8766 -21070 8778 -20894
rect 8812 -21070 8824 -20894
rect 8766 -21082 8824 -21070
rect 9224 -20894 9282 -20882
rect 9224 -21070 9236 -20894
rect 9270 -21070 9282 -20894
rect 9224 -21082 9282 -21070
rect 9682 -20894 9740 -20882
rect 9682 -21070 9694 -20894
rect 9728 -21070 9740 -20894
rect 9682 -21082 9740 -21070
rect 10140 -20894 10198 -20882
rect 10140 -21070 10152 -20894
rect 10186 -21070 10198 -20894
rect 10140 -21082 10198 -21070
rect 10598 -20894 10656 -20882
rect 10598 -21070 10610 -20894
rect 10644 -21070 10656 -20894
rect 10598 -21082 10656 -21070
rect 11056 -20894 11114 -20882
rect 11056 -21070 11068 -20894
rect 11102 -21070 11114 -20894
rect 11056 -21082 11114 -21070
rect 11514 -20894 11572 -20882
rect 11514 -21070 11526 -20894
rect 11560 -21070 11572 -20894
rect 11514 -21082 11572 -21070
rect 11972 -20894 12030 -20882
rect 11972 -21070 11984 -20894
rect 12018 -21070 12030 -20894
rect 11972 -21082 12030 -21070
rect 12430 -20894 12488 -20882
rect 12430 -21070 12442 -20894
rect 12476 -21070 12488 -20894
rect 12430 -21082 12488 -21070
rect 12888 -20894 12946 -20882
rect 12888 -21070 12900 -20894
rect 12934 -21070 12946 -20894
rect 12888 -21082 12946 -21070
rect 13346 -20894 13404 -20882
rect 13346 -21070 13358 -20894
rect 13392 -21070 13404 -20894
rect 13346 -21082 13404 -21070
rect 23766 -20226 23824 -20214
rect 23766 -20402 23778 -20226
rect 23812 -20402 23824 -20226
rect 23766 -20414 23824 -20402
rect 24224 -20226 24282 -20214
rect 24224 -20402 24236 -20226
rect 24270 -20402 24282 -20226
rect 24224 -20414 24282 -20402
rect 24682 -20226 24740 -20214
rect 24682 -20402 24694 -20226
rect 24728 -20402 24740 -20226
rect 24682 -20414 24740 -20402
rect 25140 -20226 25198 -20214
rect 25140 -20402 25152 -20226
rect 25186 -20402 25198 -20226
rect 25140 -20414 25198 -20402
rect 25598 -20226 25656 -20214
rect 25598 -20402 25610 -20226
rect 25644 -20402 25656 -20226
rect 25598 -20414 25656 -20402
rect 26056 -20226 26114 -20214
rect 26056 -20402 26068 -20226
rect 26102 -20402 26114 -20226
rect 26056 -20414 26114 -20402
rect 26514 -20226 26572 -20214
rect 26514 -20402 26526 -20226
rect 26560 -20402 26572 -20226
rect 26514 -20414 26572 -20402
rect 26972 -20226 27030 -20214
rect 26972 -20402 26984 -20226
rect 27018 -20402 27030 -20226
rect 26972 -20414 27030 -20402
rect 27430 -20226 27488 -20214
rect 27430 -20402 27442 -20226
rect 27476 -20402 27488 -20226
rect 27430 -20414 27488 -20402
rect 27888 -20226 27946 -20214
rect 27888 -20402 27900 -20226
rect 27934 -20402 27946 -20226
rect 27888 -20414 27946 -20402
rect 28346 -20226 28404 -20214
rect 28346 -20402 28358 -20226
rect 28392 -20402 28404 -20226
rect 28346 -20414 28404 -20402
rect 28766 -20226 28824 -20214
rect 28766 -20402 28778 -20226
rect 28812 -20402 28824 -20226
rect 28766 -20414 28824 -20402
rect 29224 -20226 29282 -20214
rect 29224 -20402 29236 -20226
rect 29270 -20402 29282 -20226
rect 29224 -20414 29282 -20402
rect 29682 -20226 29740 -20214
rect 29682 -20402 29694 -20226
rect 29728 -20402 29740 -20226
rect 29682 -20414 29740 -20402
rect 30140 -20226 30198 -20214
rect 30140 -20402 30152 -20226
rect 30186 -20402 30198 -20226
rect 30140 -20414 30198 -20402
rect 30598 -20226 30656 -20214
rect 30598 -20402 30610 -20226
rect 30644 -20402 30656 -20226
rect 30598 -20414 30656 -20402
rect 31056 -20226 31114 -20214
rect 31056 -20402 31068 -20226
rect 31102 -20402 31114 -20226
rect 31056 -20414 31114 -20402
rect 31514 -20226 31572 -20214
rect 31514 -20402 31526 -20226
rect 31560 -20402 31572 -20226
rect 31514 -20414 31572 -20402
rect 31972 -20226 32030 -20214
rect 31972 -20402 31984 -20226
rect 32018 -20402 32030 -20226
rect 31972 -20414 32030 -20402
rect 32430 -20226 32488 -20214
rect 32430 -20402 32442 -20226
rect 32476 -20402 32488 -20226
rect 32430 -20414 32488 -20402
rect 32888 -20226 32946 -20214
rect 32888 -20402 32900 -20226
rect 32934 -20402 32946 -20226
rect 32888 -20414 32946 -20402
rect 33346 -20226 33404 -20214
rect 33346 -20402 33358 -20226
rect 33392 -20402 33404 -20226
rect 33346 -20414 33404 -20402
rect 23766 -20894 23824 -20882
rect 23766 -21070 23778 -20894
rect 23812 -21070 23824 -20894
rect 23766 -21082 23824 -21070
rect 24224 -20894 24282 -20882
rect 24224 -21070 24236 -20894
rect 24270 -21070 24282 -20894
rect 24224 -21082 24282 -21070
rect 24682 -20894 24740 -20882
rect 24682 -21070 24694 -20894
rect 24728 -21070 24740 -20894
rect 24682 -21082 24740 -21070
rect 25140 -20894 25198 -20882
rect 25140 -21070 25152 -20894
rect 25186 -21070 25198 -20894
rect 25140 -21082 25198 -21070
rect 25598 -20894 25656 -20882
rect 25598 -21070 25610 -20894
rect 25644 -21070 25656 -20894
rect 25598 -21082 25656 -21070
rect 26056 -20894 26114 -20882
rect 26056 -21070 26068 -20894
rect 26102 -21070 26114 -20894
rect 26056 -21082 26114 -21070
rect 26514 -20894 26572 -20882
rect 26514 -21070 26526 -20894
rect 26560 -21070 26572 -20894
rect 26514 -21082 26572 -21070
rect 26972 -20894 27030 -20882
rect 26972 -21070 26984 -20894
rect 27018 -21070 27030 -20894
rect 26972 -21082 27030 -21070
rect 27430 -20894 27488 -20882
rect 27430 -21070 27442 -20894
rect 27476 -21070 27488 -20894
rect 27430 -21082 27488 -21070
rect 27888 -20894 27946 -20882
rect 27888 -21070 27900 -20894
rect 27934 -21070 27946 -20894
rect 27888 -21082 27946 -21070
rect 28346 -20894 28404 -20882
rect 28346 -21070 28358 -20894
rect 28392 -21070 28404 -20894
rect 28346 -21082 28404 -21070
<< pdiff >>
rect 23764 16422 23822 16434
rect 23764 16246 23776 16422
rect 23810 16246 23822 16422
rect 23764 16234 23822 16246
rect 24622 16422 24680 16434
rect 24622 16246 24634 16422
rect 24668 16246 24680 16422
rect 24622 16234 24680 16246
rect 25480 16422 25538 16434
rect 25480 16246 25492 16422
rect 25526 16246 25538 16422
rect 25480 16234 25538 16246
rect 26338 16422 26396 16434
rect 26338 16246 26350 16422
rect 26384 16246 26396 16422
rect 26338 16234 26396 16246
rect 27196 16422 27254 16434
rect 27196 16246 27208 16422
rect 27242 16246 27254 16422
rect 27196 16234 27254 16246
rect 28054 16422 28112 16434
rect 28054 16246 28066 16422
rect 28100 16246 28112 16422
rect 28054 16234 28112 16246
rect 28912 16422 28970 16434
rect 28912 16246 28924 16422
rect 28958 16246 28970 16422
rect 28912 16234 28970 16246
rect 29770 16422 29828 16434
rect 29770 16246 29782 16422
rect 29816 16246 29828 16422
rect 29770 16234 29828 16246
rect 30628 16422 30686 16434
rect 30628 16246 30640 16422
rect 30674 16246 30686 16422
rect 30628 16234 30686 16246
rect 31486 16422 31544 16434
rect 31486 16246 31498 16422
rect 31532 16246 31544 16422
rect 31486 16234 31544 16246
rect 32344 16422 32402 16434
rect 32344 16246 32356 16422
rect 32390 16246 32402 16422
rect 32344 16234 32402 16246
rect 23764 15822 23822 15834
rect 23764 15646 23776 15822
rect 23810 15646 23822 15822
rect 23764 15634 23822 15646
rect 24622 15822 24680 15834
rect 24622 15646 24634 15822
rect 24668 15646 24680 15822
rect 24622 15634 24680 15646
rect 25480 15822 25538 15834
rect 25480 15646 25492 15822
rect 25526 15646 25538 15822
rect 25480 15634 25538 15646
rect 26338 15822 26396 15834
rect 26338 15646 26350 15822
rect 26384 15646 26396 15822
rect 26338 15634 26396 15646
rect 27196 15822 27254 15834
rect 27196 15646 27208 15822
rect 27242 15646 27254 15822
rect 27196 15634 27254 15646
rect 28054 15822 28112 15834
rect 28054 15646 28066 15822
rect 28100 15646 28112 15822
rect 28054 15634 28112 15646
rect 28912 15822 28970 15834
rect 28912 15646 28924 15822
rect 28958 15646 28970 15822
rect 28912 15634 28970 15646
rect 29770 15822 29828 15834
rect 29770 15646 29782 15822
rect 29816 15646 29828 15822
rect 29770 15634 29828 15646
rect 30628 15822 30686 15834
rect 30628 15646 30640 15822
rect 30674 15646 30686 15822
rect 30628 15634 30686 15646
rect 31486 15822 31544 15834
rect 31486 15646 31498 15822
rect 31532 15646 31544 15822
rect 31486 15634 31544 15646
rect 32344 15822 32402 15834
rect 32344 15646 32356 15822
rect 32390 15646 32402 15822
rect 32344 15634 32402 15646
rect 24151 14782 24209 14794
rect 24151 14406 24163 14782
rect 24197 14406 24209 14782
rect 24151 14394 24209 14406
rect 24409 14782 24467 14794
rect 24409 14406 24421 14782
rect 24455 14406 24467 14782
rect 24409 14394 24467 14406
rect 24667 14782 24725 14794
rect 24667 14406 24679 14782
rect 24713 14406 24725 14782
rect 24667 14394 24725 14406
rect 24925 14782 24983 14794
rect 24925 14406 24937 14782
rect 24971 14406 24983 14782
rect 24925 14394 24983 14406
rect 25273 14782 25331 14794
rect 25273 14406 25285 14782
rect 25319 14406 25331 14782
rect 25273 14394 25331 14406
rect 25531 14782 25589 14794
rect 25531 14406 25543 14782
rect 25577 14406 25589 14782
rect 25531 14394 25589 14406
rect 25789 14782 25847 14794
rect 25789 14406 25801 14782
rect 25835 14406 25847 14782
rect 25789 14394 25847 14406
rect 26047 14782 26105 14794
rect 26047 14406 26059 14782
rect 26093 14406 26105 14782
rect 26047 14394 26105 14406
rect 26305 14782 26363 14794
rect 26305 14406 26317 14782
rect 26351 14406 26363 14782
rect 26305 14394 26363 14406
rect 26563 14782 26621 14794
rect 26563 14406 26575 14782
rect 26609 14406 26621 14782
rect 26563 14394 26621 14406
rect 26821 14782 26879 14794
rect 26821 14406 26833 14782
rect 26867 14406 26879 14782
rect 26821 14394 26879 14406
rect 27287 14391 27339 14405
rect 27287 14357 27295 14391
rect 27329 14357 27339 14391
rect 27287 14323 27339 14357
rect 27287 14289 27295 14323
rect 27329 14289 27339 14323
rect 27287 14277 27339 14289
rect 27369 14375 27423 14405
rect 27369 14341 27379 14375
rect 27413 14341 27423 14375
rect 27369 14277 27423 14341
rect 27453 14391 27505 14405
rect 27453 14357 27463 14391
rect 27497 14357 27505 14391
rect 27453 14323 27505 14357
rect 27638 14399 27690 14411
rect 27638 14365 27646 14399
rect 27680 14365 27690 14399
rect 27638 14327 27690 14365
rect 27720 14391 27782 14411
rect 27720 14357 27730 14391
rect 27764 14357 27782 14391
rect 27720 14327 27782 14357
rect 27812 14397 27881 14411
rect 27812 14363 27823 14397
rect 27857 14363 27881 14397
rect 27812 14327 27881 14363
rect 27911 14373 28021 14411
rect 27911 14339 27977 14373
rect 28011 14339 28021 14373
rect 27911 14327 28021 14339
rect 28051 14389 28118 14411
rect 28051 14355 28074 14389
rect 28108 14355 28118 14389
rect 28051 14327 28118 14355
rect 28148 14373 28200 14411
rect 28148 14339 28158 14373
rect 28192 14339 28200 14373
rect 28148 14327 28200 14339
rect 28263 14399 28315 14411
rect 28263 14365 28271 14399
rect 28305 14365 28315 14399
rect 27453 14289 27463 14323
rect 27497 14289 27505 14323
rect 27453 14277 27505 14289
rect 28263 14243 28315 14365
rect 28345 14391 28414 14411
rect 28345 14357 28359 14391
rect 28393 14357 28414 14391
rect 28345 14327 28414 14357
rect 28444 14398 28500 14411
rect 28444 14364 28456 14398
rect 28490 14364 28500 14398
rect 28444 14327 28500 14364
rect 28530 14327 28584 14411
rect 28614 14399 28692 14411
rect 28614 14365 28648 14399
rect 28682 14365 28692 14399
rect 28614 14327 28692 14365
rect 28722 14373 28776 14411
rect 28722 14339 28732 14373
rect 28766 14339 28776 14373
rect 28722 14327 28776 14339
rect 28806 14399 28940 14411
rect 28806 14365 28818 14399
rect 28852 14365 28896 14399
rect 28930 14365 28940 14399
rect 28806 14327 28940 14365
rect 28345 14243 28399 14327
rect 28890 14211 28940 14327
rect 28970 14391 29026 14411
rect 28970 14357 28980 14391
rect 29014 14357 29026 14391
rect 28970 14323 29026 14357
rect 28970 14289 28980 14323
rect 29014 14289 29026 14323
rect 28970 14255 29026 14289
rect 29107 14399 29159 14411
rect 29107 14365 29115 14399
rect 29149 14365 29159 14399
rect 29107 14331 29159 14365
rect 29107 14297 29115 14331
rect 29149 14297 29159 14331
rect 29107 14283 29159 14297
rect 29189 14399 29256 14411
rect 29189 14365 29212 14399
rect 29246 14365 29256 14399
rect 29189 14331 29256 14365
rect 29189 14297 29212 14331
rect 29246 14297 29256 14331
rect 29189 14283 29256 14297
rect 28970 14221 28980 14255
rect 29014 14221 29026 14255
rect 28970 14211 29026 14221
rect 29204 14263 29256 14283
rect 29204 14229 29212 14263
rect 29246 14229 29256 14263
rect 29204 14211 29256 14229
rect 29286 14363 29338 14411
rect 29286 14329 29296 14363
rect 29330 14329 29338 14363
rect 29286 14295 29338 14329
rect 29286 14261 29296 14295
rect 29330 14261 29338 14295
rect 29286 14211 29338 14261
rect 29444 14399 29496 14411
rect 29444 14365 29452 14399
rect 29486 14365 29496 14399
rect 29444 14331 29496 14365
rect 29444 14297 29452 14331
rect 29486 14297 29496 14331
rect 29444 14263 29496 14297
rect 29444 14229 29452 14263
rect 29486 14229 29496 14263
rect 29444 14211 29496 14229
rect 29526 14399 29578 14411
rect 29526 14365 29536 14399
rect 29570 14365 29578 14399
rect 29526 14331 29578 14365
rect 29526 14297 29536 14331
rect 29570 14297 29578 14331
rect 29526 14263 29578 14297
rect 29526 14229 29536 14263
rect 29570 14229 29578 14263
rect 29526 14211 29578 14229
rect 29683 14399 29735 14411
rect 29683 14365 29691 14399
rect 29725 14365 29735 14399
rect 29683 14331 29735 14365
rect 29683 14297 29691 14331
rect 29725 14297 29735 14331
rect 29683 14263 29735 14297
rect 29683 14229 29691 14263
rect 29725 14229 29735 14263
rect 29683 14211 29735 14229
rect 29765 14399 29819 14411
rect 29765 14365 29775 14399
rect 29809 14365 29819 14399
rect 29765 14331 29819 14365
rect 29765 14297 29775 14331
rect 29809 14297 29819 14331
rect 29765 14263 29819 14297
rect 29765 14229 29775 14263
rect 29809 14229 29819 14263
rect 29765 14211 29819 14229
rect 29849 14399 29901 14411
rect 29849 14365 29859 14399
rect 29893 14365 29901 14399
rect 29849 14331 29901 14365
rect 29849 14297 29859 14331
rect 29893 14297 29901 14331
rect 29849 14263 29901 14297
rect 29849 14229 29859 14263
rect 29893 14229 29901 14263
rect 29849 14211 29901 14229
rect 30002 14399 30054 14411
rect 30002 14365 30010 14399
rect 30044 14365 30054 14399
rect 30002 14331 30054 14365
rect 30002 14297 30010 14331
rect 30044 14297 30054 14331
rect 30002 14263 30054 14297
rect 30002 14229 30010 14263
rect 30044 14229 30054 14263
rect 30002 14211 30054 14229
rect 30084 14399 30136 14411
rect 30084 14365 30094 14399
rect 30128 14365 30136 14399
rect 30084 14331 30136 14365
rect 30084 14297 30094 14331
rect 30128 14297 30136 14331
rect 30084 14263 30136 14297
rect 30084 14229 30094 14263
rect 30128 14229 30136 14263
rect 30084 14211 30136 14229
rect 30242 14363 30294 14411
rect 30242 14329 30250 14363
rect 30284 14329 30294 14363
rect 30242 14295 30294 14329
rect 30242 14261 30250 14295
rect 30284 14261 30294 14295
rect 30242 14211 30294 14261
rect 30324 14399 30391 14411
rect 30324 14365 30334 14399
rect 30368 14365 30391 14399
rect 30324 14331 30391 14365
rect 30324 14297 30334 14331
rect 30368 14297 30391 14331
rect 30324 14283 30391 14297
rect 30421 14399 30473 14411
rect 30421 14365 30431 14399
rect 30465 14365 30473 14399
rect 30421 14331 30473 14365
rect 30421 14297 30431 14331
rect 30465 14297 30473 14331
rect 30421 14283 30473 14297
rect 30554 14391 30610 14411
rect 30554 14357 30566 14391
rect 30600 14357 30610 14391
rect 30554 14323 30610 14357
rect 30554 14289 30566 14323
rect 30600 14289 30610 14323
rect 30324 14263 30376 14283
rect 30324 14229 30334 14263
rect 30368 14229 30376 14263
rect 30324 14211 30376 14229
rect 30554 14255 30610 14289
rect 30554 14221 30566 14255
rect 30600 14221 30610 14255
rect 30554 14211 30610 14221
rect 30640 14399 30774 14411
rect 30640 14365 30650 14399
rect 30684 14365 30728 14399
rect 30762 14365 30774 14399
rect 30640 14327 30774 14365
rect 30804 14373 30858 14411
rect 30804 14339 30814 14373
rect 30848 14339 30858 14373
rect 30804 14327 30858 14339
rect 30888 14399 30966 14411
rect 30888 14365 30898 14399
rect 30932 14365 30966 14399
rect 30888 14327 30966 14365
rect 30996 14327 31050 14411
rect 31080 14398 31136 14411
rect 31080 14364 31090 14398
rect 31124 14364 31136 14398
rect 31080 14327 31136 14364
rect 31166 14391 31235 14411
rect 31166 14357 31187 14391
rect 31221 14357 31235 14391
rect 31166 14327 31235 14357
rect 30640 14211 30690 14327
rect 31181 14243 31235 14327
rect 31265 14399 31317 14411
rect 31265 14365 31275 14399
rect 31309 14365 31317 14399
rect 31265 14243 31317 14365
rect 31380 14373 31432 14411
rect 31380 14339 31388 14373
rect 31422 14339 31432 14373
rect 31380 14327 31432 14339
rect 31462 14389 31529 14411
rect 31462 14355 31472 14389
rect 31506 14355 31529 14389
rect 31462 14327 31529 14355
rect 31559 14373 31669 14411
rect 31559 14339 31569 14373
rect 31603 14339 31669 14373
rect 31559 14327 31669 14339
rect 31699 14397 31768 14411
rect 31699 14363 31723 14397
rect 31757 14363 31768 14397
rect 31699 14327 31768 14363
rect 31798 14391 31860 14411
rect 31798 14357 31816 14391
rect 31850 14357 31860 14391
rect 31798 14327 31860 14357
rect 31890 14399 31942 14411
rect 31890 14365 31900 14399
rect 31934 14365 31942 14399
rect 31890 14327 31942 14365
rect 32075 14391 32127 14405
rect 32075 14357 32083 14391
rect 32117 14357 32127 14391
rect 32075 14323 32127 14357
rect 32075 14289 32083 14323
rect 32117 14289 32127 14323
rect 32075 14277 32127 14289
rect 32157 14375 32211 14405
rect 32157 14341 32167 14375
rect 32201 14341 32211 14375
rect 32157 14277 32211 14341
rect 32241 14391 32293 14405
rect 32241 14357 32251 14391
rect 32285 14357 32293 14391
rect 32241 14323 32293 14357
rect 32241 14289 32251 14323
rect 32285 14289 32293 14323
rect 32241 14277 32293 14289
rect 30579 8893 30631 8907
rect 30579 8859 30587 8893
rect 30621 8859 30631 8893
rect 30579 8825 30631 8859
rect 30579 8791 30587 8825
rect 30621 8791 30631 8825
rect 30579 8779 30631 8791
rect 30661 8877 30715 8907
rect 30661 8843 30671 8877
rect 30705 8843 30715 8877
rect 30661 8779 30715 8843
rect 30745 8893 30797 8907
rect 30745 8859 30755 8893
rect 30789 8859 30797 8893
rect 30745 8825 30797 8859
rect 30851 8901 30903 8913
rect 30851 8867 30859 8901
rect 30893 8867 30903 8901
rect 30851 8829 30903 8867
rect 30933 8893 30988 8913
rect 30933 8859 30943 8893
rect 30977 8859 30988 8893
rect 30933 8829 30988 8859
rect 31018 8888 31083 8913
rect 31018 8854 31035 8888
rect 31069 8854 31083 8888
rect 31018 8829 31083 8854
rect 31113 8829 31186 8913
rect 31216 8901 31318 8913
rect 31216 8867 31274 8901
rect 31308 8867 31318 8901
rect 31216 8833 31318 8867
rect 31216 8829 31274 8833
rect 30745 8791 30755 8825
rect 30789 8791 30797 8825
rect 30745 8779 30797 8791
rect 13324 7805 13382 7817
rect 13324 6229 13336 7805
rect 13370 6229 13382 7805
rect 13324 6217 13382 6229
rect 13782 7805 13840 7817
rect 13782 6229 13794 7805
rect 13828 6229 13840 7805
rect 13782 6217 13840 6229
rect 14240 7805 14298 7817
rect 14240 6229 14252 7805
rect 14286 6229 14298 7805
rect 14240 6217 14298 6229
rect 14698 7805 14756 7817
rect 14698 6229 14710 7805
rect 14744 6229 14756 7805
rect 14698 6217 14756 6229
rect 15156 7805 15214 7817
rect 15156 6229 15168 7805
rect 15202 6229 15214 7805
rect 15156 6217 15214 6229
rect 15614 7805 15672 7817
rect 15614 6229 15626 7805
rect 15660 6229 15672 7805
rect 15614 6217 15672 6229
rect 16072 7805 16130 7817
rect 16072 6229 16084 7805
rect 16118 6229 16130 7805
rect 16072 6217 16130 6229
rect 16530 7805 16588 7817
rect 16530 6229 16542 7805
rect 16576 6229 16588 7805
rect 16530 6217 16588 6229
rect 16988 7805 17046 7817
rect 16988 6229 17000 7805
rect 17034 6229 17046 7805
rect 16988 6217 17046 6229
rect 17446 7805 17504 7817
rect 17446 6229 17458 7805
rect 17492 6229 17504 7805
rect 17446 6217 17504 6229
rect 17904 7805 17962 7817
rect 17904 6229 17916 7805
rect 17950 6229 17962 7805
rect 17904 6217 17962 6229
rect 18362 7805 18420 7817
rect 18362 6229 18374 7805
rect 18408 6229 18420 7805
rect 18362 6217 18420 6229
rect 18820 7805 18878 7817
rect 18820 6229 18832 7805
rect 18866 6229 18878 7805
rect 18820 6217 18878 6229
rect 19278 7805 19336 7817
rect 19278 6229 19290 7805
rect 19324 6229 19336 7805
rect 19278 6217 19336 6229
rect 19736 7805 19794 7817
rect 19736 6229 19748 7805
rect 19782 6229 19794 7805
rect 19736 6217 19794 6229
rect 20194 7805 20252 7817
rect 20194 6229 20206 7805
rect 20240 6229 20252 7805
rect 20194 6217 20252 6229
rect 20652 7805 20710 7817
rect 20652 6229 20664 7805
rect 20698 6229 20710 7805
rect 20652 6217 20710 6229
rect 21110 7805 21168 7817
rect 21110 6229 21122 7805
rect 21156 6229 21168 7805
rect 21110 6217 21168 6229
rect 21568 7805 21626 7817
rect 21568 6229 21580 7805
rect 21614 6229 21626 7805
rect 21568 6217 21626 6229
rect 23919 8225 23977 8237
rect 23919 7049 23931 8225
rect 23965 7049 23977 8225
rect 23919 7037 23977 7049
rect 24377 8225 24435 8237
rect 24377 7049 24389 8225
rect 24423 7049 24435 8225
rect 24377 7037 24435 7049
rect 24835 8225 24893 8237
rect 24835 7049 24847 8225
rect 24881 7049 24893 8225
rect 24835 7037 24893 7049
rect 25293 8225 25351 8237
rect 25293 7049 25305 8225
rect 25339 7049 25351 8225
rect 25293 7037 25351 7049
rect 25751 8225 25809 8237
rect 25751 7049 25763 8225
rect 25797 7049 25809 8225
rect 25751 7037 25809 7049
rect 26209 8225 26267 8237
rect 26209 7049 26221 8225
rect 26255 7049 26267 8225
rect 26209 7037 26267 7049
rect 26667 8225 26725 8237
rect 26667 7049 26679 8225
rect 26713 7049 26725 8225
rect 26667 7037 26725 7049
rect 27125 8225 27183 8237
rect 27125 7049 27137 8225
rect 27171 7049 27183 8225
rect 27125 7037 27183 7049
rect 27583 8225 27641 8237
rect 27583 7049 27595 8225
rect 27629 7049 27641 8225
rect 27583 7037 27641 7049
rect 28041 8225 28099 8237
rect 28041 7049 28053 8225
rect 28087 7049 28099 8225
rect 28041 7037 28099 7049
rect 28499 8225 28557 8237
rect 28499 7049 28511 8225
rect 28545 7049 28557 8225
rect 28499 7037 28557 7049
rect 29144 8599 29196 8617
rect 29144 8565 29152 8599
rect 29186 8565 29196 8599
rect 29144 8531 29196 8565
rect 29144 8497 29152 8531
rect 29186 8497 29196 8531
rect 29144 8463 29196 8497
rect 29144 8429 29152 8463
rect 29186 8429 29196 8463
rect 29144 8417 29196 8429
rect 29226 8599 29278 8617
rect 29226 8565 29236 8599
rect 29270 8565 29278 8599
rect 29226 8531 29278 8565
rect 29226 8497 29236 8531
rect 29270 8497 29278 8531
rect 29226 8463 29278 8497
rect 29226 8429 29236 8463
rect 29270 8429 29278 8463
rect 29226 8417 29278 8429
rect 29389 8599 29441 8617
rect 29389 8565 29397 8599
rect 29431 8565 29441 8599
rect 29389 8531 29441 8565
rect 29389 8497 29397 8531
rect 29431 8497 29441 8531
rect 29389 8463 29441 8497
rect 29389 8429 29397 8463
rect 29431 8429 29441 8463
rect 29389 8417 29441 8429
rect 29471 8599 29525 8617
rect 29471 8565 29481 8599
rect 29515 8565 29525 8599
rect 29471 8531 29525 8565
rect 29471 8497 29481 8531
rect 29515 8497 29525 8531
rect 29471 8463 29525 8497
rect 29471 8429 29481 8463
rect 29515 8429 29525 8463
rect 29471 8417 29525 8429
rect 29555 8531 29609 8617
rect 29555 8497 29565 8531
rect 29599 8497 29609 8531
rect 29555 8463 29609 8497
rect 29555 8429 29565 8463
rect 29599 8429 29609 8463
rect 29555 8417 29609 8429
rect 29639 8599 29693 8617
rect 29639 8565 29649 8599
rect 29683 8565 29693 8599
rect 29639 8531 29693 8565
rect 29639 8497 29649 8531
rect 29683 8497 29693 8531
rect 29639 8463 29693 8497
rect 29639 8429 29649 8463
rect 29683 8429 29693 8463
rect 29639 8417 29693 8429
rect 29723 8463 29775 8617
rect 31231 8799 31274 8829
rect 31308 8799 31318 8833
rect 31231 8763 31318 8799
rect 31348 8893 31413 8913
rect 31348 8859 31358 8893
rect 31392 8859 31413 8893
rect 31348 8829 31413 8859
rect 31443 8883 31497 8913
rect 31443 8849 31453 8883
rect 31487 8849 31497 8883
rect 31443 8829 31497 8849
rect 31527 8829 31611 8913
rect 31641 8893 31694 8913
rect 31641 8859 31652 8893
rect 31686 8859 31694 8893
rect 31641 8829 31694 8859
rect 31768 8901 31822 8913
rect 31768 8867 31776 8901
rect 31810 8867 31822 8901
rect 31768 8830 31822 8867
rect 31348 8763 31398 8829
rect 31768 8796 31776 8830
rect 31810 8796 31822 8830
rect 31768 8759 31822 8796
rect 31768 8725 31776 8759
rect 31810 8725 31822 8759
rect 31768 8713 31822 8725
rect 31852 8871 31906 8913
rect 31852 8837 31862 8871
rect 31896 8837 31906 8871
rect 31852 8791 31906 8837
rect 31852 8757 31862 8791
rect 31896 8757 31906 8791
rect 31852 8713 31906 8757
rect 31936 8895 31988 8913
rect 31936 8861 31946 8895
rect 31980 8861 31988 8895
rect 31936 8827 31988 8861
rect 31936 8793 31946 8827
rect 31980 8793 31988 8827
rect 31936 8759 31988 8793
rect 32042 8901 32094 8913
rect 32042 8867 32050 8901
rect 32084 8867 32094 8901
rect 32042 8833 32094 8867
rect 32042 8799 32050 8833
rect 32084 8799 32094 8833
rect 32042 8785 32094 8799
rect 32124 8901 32191 8913
rect 32124 8867 32147 8901
rect 32181 8867 32191 8901
rect 32124 8833 32191 8867
rect 32124 8799 32147 8833
rect 32181 8799 32191 8833
rect 32124 8785 32191 8799
rect 31936 8725 31946 8759
rect 31980 8725 31988 8759
rect 31936 8713 31988 8725
rect 32139 8765 32191 8785
rect 32139 8731 32147 8765
rect 32181 8731 32191 8765
rect 32139 8713 32191 8731
rect 32221 8901 32273 8913
rect 32221 8867 32231 8901
rect 32265 8867 32273 8901
rect 32221 8830 32273 8867
rect 32221 8796 32231 8830
rect 32265 8796 32273 8830
rect 32221 8759 32273 8796
rect 32221 8725 32231 8759
rect 32265 8725 32273 8759
rect 32221 8713 32273 8725
rect 32368 8901 32420 8913
rect 32368 8867 32376 8901
rect 32410 8867 32420 8901
rect 32368 8833 32420 8867
rect 32368 8799 32376 8833
rect 32410 8799 32420 8833
rect 32368 8765 32420 8799
rect 32368 8731 32376 8765
rect 32410 8731 32420 8765
rect 32368 8713 32420 8731
rect 32450 8901 32502 8913
rect 32450 8867 32460 8901
rect 32494 8867 32502 8901
rect 32450 8833 32502 8867
rect 32450 8799 32460 8833
rect 32494 8799 32502 8833
rect 32450 8765 32502 8799
rect 32450 8731 32460 8765
rect 32494 8731 32502 8765
rect 32450 8713 32502 8731
rect 32613 8901 32665 8913
rect 32613 8867 32621 8901
rect 32655 8867 32665 8901
rect 32613 8833 32665 8867
rect 32613 8799 32621 8833
rect 32655 8799 32665 8833
rect 32613 8765 32665 8799
rect 32613 8731 32621 8765
rect 32655 8731 32665 8765
rect 32613 8713 32665 8731
rect 32695 8901 32749 8913
rect 32695 8867 32705 8901
rect 32739 8867 32749 8901
rect 32695 8833 32749 8867
rect 32695 8799 32705 8833
rect 32739 8799 32749 8833
rect 32695 8765 32749 8799
rect 32695 8731 32705 8765
rect 32739 8731 32749 8765
rect 32695 8713 32749 8731
rect 32779 8901 32833 8913
rect 32779 8867 32789 8901
rect 32823 8867 32833 8901
rect 32779 8833 32833 8867
rect 32779 8799 32789 8833
rect 32823 8799 32833 8833
rect 32779 8713 32833 8799
rect 32863 8901 32917 8913
rect 32863 8867 32873 8901
rect 32907 8867 32917 8901
rect 32863 8833 32917 8867
rect 32863 8799 32873 8833
rect 32907 8799 32917 8833
rect 32863 8765 32917 8799
rect 32863 8731 32873 8765
rect 32907 8731 32917 8765
rect 32863 8713 32917 8731
rect 32947 8901 32999 8913
rect 32947 8867 32957 8901
rect 32991 8867 32999 8901
rect 32947 8713 32999 8867
rect 29723 8429 29733 8463
rect 29767 8429 29775 8463
rect 29723 8417 29775 8429
rect 30579 8041 30631 8053
rect 30579 8007 30587 8041
rect 30621 8007 30631 8041
rect 30579 7973 30631 8007
rect 30579 7939 30587 7973
rect 30621 7939 30631 7973
rect 30579 7925 30631 7939
rect 30661 7989 30715 8053
rect 30661 7955 30671 7989
rect 30705 7955 30715 7989
rect 30661 7925 30715 7955
rect 30745 8041 30797 8053
rect 30745 8007 30755 8041
rect 30789 8007 30797 8041
rect 30745 7973 30797 8007
rect 31768 8107 31822 8119
rect 31231 8033 31318 8069
rect 31231 8003 31274 8033
rect 30745 7939 30755 7973
rect 30789 7939 30797 7973
rect 30745 7925 30797 7939
rect 30851 7965 30903 8003
rect 30851 7931 30859 7965
rect 30893 7931 30903 7965
rect 30851 7919 30903 7931
rect 30933 7973 30988 8003
rect 30933 7939 30943 7973
rect 30977 7939 30988 7973
rect 30933 7919 30988 7939
rect 31018 7978 31083 8003
rect 31018 7944 31035 7978
rect 31069 7944 31083 7978
rect 31018 7919 31083 7944
rect 31113 7919 31186 8003
rect 31216 7999 31274 8003
rect 31308 7999 31318 8033
rect 31216 7965 31318 7999
rect 31216 7931 31274 7965
rect 31308 7931 31318 7965
rect 31216 7919 31318 7931
rect 31348 8003 31398 8069
rect 31768 8073 31776 8107
rect 31810 8073 31822 8107
rect 31768 8036 31822 8073
rect 31348 7973 31413 8003
rect 31348 7939 31358 7973
rect 31392 7939 31413 7973
rect 31348 7919 31413 7939
rect 31443 7983 31497 8003
rect 31443 7949 31453 7983
rect 31487 7949 31497 7983
rect 31443 7919 31497 7949
rect 31527 7919 31611 8003
rect 31641 7973 31694 8003
rect 31641 7939 31652 7973
rect 31686 7939 31694 7973
rect 31641 7919 31694 7939
rect 31768 8002 31776 8036
rect 31810 8002 31822 8036
rect 31768 7965 31822 8002
rect 31768 7931 31776 7965
rect 31810 7931 31822 7965
rect 31768 7919 31822 7931
rect 31852 8075 31906 8119
rect 31852 8041 31862 8075
rect 31896 8041 31906 8075
rect 31852 7995 31906 8041
rect 31852 7961 31862 7995
rect 31896 7961 31906 7995
rect 31852 7919 31906 7961
rect 31936 8107 31988 8119
rect 31936 8073 31946 8107
rect 31980 8073 31988 8107
rect 31936 8039 31988 8073
rect 32139 8101 32191 8119
rect 32139 8067 32147 8101
rect 32181 8067 32191 8101
rect 32139 8047 32191 8067
rect 31936 8005 31946 8039
rect 31980 8005 31988 8039
rect 31936 7971 31988 8005
rect 31936 7937 31946 7971
rect 31980 7937 31988 7971
rect 31936 7919 31988 7937
rect 32042 8033 32094 8047
rect 32042 7999 32050 8033
rect 32084 7999 32094 8033
rect 32042 7965 32094 7999
rect 32042 7931 32050 7965
rect 32084 7931 32094 7965
rect 32042 7919 32094 7931
rect 32124 8033 32191 8047
rect 32124 7999 32147 8033
rect 32181 7999 32191 8033
rect 32124 7965 32191 7999
rect 32124 7931 32147 7965
rect 32181 7931 32191 7965
rect 32124 7919 32191 7931
rect 32221 8107 32273 8119
rect 32221 8073 32231 8107
rect 32265 8073 32273 8107
rect 32221 8036 32273 8073
rect 32221 8002 32231 8036
rect 32265 8002 32273 8036
rect 32221 7965 32273 8002
rect 32221 7931 32231 7965
rect 32265 7931 32273 7965
rect 32221 7919 32273 7931
rect 32368 8101 32420 8119
rect 32368 8067 32376 8101
rect 32410 8067 32420 8101
rect 32368 8033 32420 8067
rect 32368 7999 32376 8033
rect 32410 7999 32420 8033
rect 32368 7965 32420 7999
rect 32368 7931 32376 7965
rect 32410 7931 32420 7965
rect 32368 7919 32420 7931
rect 32450 8101 32502 8119
rect 32450 8067 32460 8101
rect 32494 8067 32502 8101
rect 32450 8033 32502 8067
rect 32450 7999 32460 8033
rect 32494 7999 32502 8033
rect 32450 7965 32502 7999
rect 32450 7931 32460 7965
rect 32494 7931 32502 7965
rect 32450 7919 32502 7931
rect 32613 8101 32665 8119
rect 32613 8067 32621 8101
rect 32655 8067 32665 8101
rect 32613 8033 32665 8067
rect 32613 7999 32621 8033
rect 32655 7999 32665 8033
rect 32613 7965 32665 7999
rect 32613 7931 32621 7965
rect 32655 7931 32665 7965
rect 32613 7919 32665 7931
rect 32695 8101 32749 8119
rect 32695 8067 32705 8101
rect 32739 8067 32749 8101
rect 32695 8033 32749 8067
rect 32695 7999 32705 8033
rect 32739 7999 32749 8033
rect 32695 7965 32749 7999
rect 32695 7931 32705 7965
rect 32739 7931 32749 7965
rect 32695 7919 32749 7931
rect 32779 8033 32833 8119
rect 32779 7999 32789 8033
rect 32823 7999 32833 8033
rect 32779 7965 32833 7999
rect 32779 7931 32789 7965
rect 32823 7931 32833 7965
rect 32779 7919 32833 7931
rect 32863 8101 32917 8119
rect 32863 8067 32873 8101
rect 32907 8067 32917 8101
rect 32863 8033 32917 8067
rect 32863 7999 32873 8033
rect 32907 7999 32917 8033
rect 32863 7965 32917 7999
rect 32863 7931 32873 7965
rect 32907 7931 32917 7965
rect 32863 7919 32917 7931
rect 32947 7965 32999 8119
rect 32947 7931 32957 7965
rect 32991 7931 32999 7965
rect 32947 7919 32999 7931
rect 33277 8041 33329 8053
rect 33277 8007 33285 8041
rect 33319 8007 33329 8041
rect 33277 7973 33329 8007
rect 33277 7939 33285 7973
rect 33319 7939 33329 7973
rect 33277 7925 33329 7939
rect 33359 7989 33413 8053
rect 33359 7955 33369 7989
rect 33403 7955 33413 7989
rect 33359 7925 33413 7955
rect 33443 8041 33495 8053
rect 33443 8007 33453 8041
rect 33487 8007 33495 8041
rect 33443 7973 33495 8007
rect 34466 8107 34520 8119
rect 33929 8033 34016 8069
rect 33929 8003 33972 8033
rect 33443 7939 33453 7973
rect 33487 7939 33495 7973
rect 33443 7925 33495 7939
rect 33549 7965 33601 8003
rect 33549 7931 33557 7965
rect 33591 7931 33601 7965
rect 33549 7919 33601 7931
rect 33631 7973 33686 8003
rect 33631 7939 33641 7973
rect 33675 7939 33686 7973
rect 33631 7919 33686 7939
rect 33716 7978 33781 8003
rect 33716 7944 33733 7978
rect 33767 7944 33781 7978
rect 33716 7919 33781 7944
rect 33811 7919 33884 8003
rect 33914 7999 33972 8003
rect 34006 7999 34016 8033
rect 33914 7965 34016 7999
rect 33914 7931 33972 7965
rect 34006 7931 34016 7965
rect 33914 7919 34016 7931
rect 34046 8003 34096 8069
rect 34466 8073 34474 8107
rect 34508 8073 34520 8107
rect 34466 8036 34520 8073
rect 34046 7973 34111 8003
rect 34046 7939 34056 7973
rect 34090 7939 34111 7973
rect 34046 7919 34111 7939
rect 34141 7983 34195 8003
rect 34141 7949 34151 7983
rect 34185 7949 34195 7983
rect 34141 7919 34195 7949
rect 34225 7919 34309 8003
rect 34339 7973 34392 8003
rect 34339 7939 34350 7973
rect 34384 7939 34392 7973
rect 34339 7919 34392 7939
rect 34466 8002 34474 8036
rect 34508 8002 34520 8036
rect 34466 7965 34520 8002
rect 34466 7931 34474 7965
rect 34508 7931 34520 7965
rect 34466 7919 34520 7931
rect 34550 8075 34604 8119
rect 34550 8041 34560 8075
rect 34594 8041 34604 8075
rect 34550 7995 34604 8041
rect 34550 7961 34560 7995
rect 34594 7961 34604 7995
rect 34550 7919 34604 7961
rect 34634 8107 34686 8119
rect 34634 8073 34644 8107
rect 34678 8073 34686 8107
rect 34634 8039 34686 8073
rect 34837 8101 34889 8119
rect 34837 8067 34845 8101
rect 34879 8067 34889 8101
rect 34837 8047 34889 8067
rect 34634 8005 34644 8039
rect 34678 8005 34686 8039
rect 34634 7971 34686 8005
rect 34634 7937 34644 7971
rect 34678 7937 34686 7971
rect 34634 7919 34686 7937
rect 34740 8033 34792 8047
rect 34740 7999 34748 8033
rect 34782 7999 34792 8033
rect 34740 7965 34792 7999
rect 34740 7931 34748 7965
rect 34782 7931 34792 7965
rect 34740 7919 34792 7931
rect 34822 8033 34889 8047
rect 34822 7999 34845 8033
rect 34879 7999 34889 8033
rect 34822 7965 34889 7999
rect 34822 7931 34845 7965
rect 34879 7931 34889 7965
rect 34822 7919 34889 7931
rect 34919 8107 34971 8119
rect 34919 8073 34929 8107
rect 34963 8073 34971 8107
rect 34919 8036 34971 8073
rect 34919 8002 34929 8036
rect 34963 8002 34971 8036
rect 34919 7965 34971 8002
rect 34919 7931 34929 7965
rect 34963 7931 34971 7965
rect 34919 7919 34971 7931
rect 35066 8101 35118 8119
rect 35066 8067 35074 8101
rect 35108 8067 35118 8101
rect 35066 8033 35118 8067
rect 35066 7999 35074 8033
rect 35108 7999 35118 8033
rect 35066 7965 35118 7999
rect 35066 7931 35074 7965
rect 35108 7931 35118 7965
rect 35066 7919 35118 7931
rect 35148 8101 35200 8119
rect 35148 8067 35158 8101
rect 35192 8067 35200 8101
rect 35148 8033 35200 8067
rect 35148 7999 35158 8033
rect 35192 7999 35200 8033
rect 35148 7965 35200 7999
rect 35148 7931 35158 7965
rect 35192 7931 35200 7965
rect 35148 7919 35200 7931
rect 35311 8101 35363 8119
rect 35311 8067 35319 8101
rect 35353 8067 35363 8101
rect 35311 8033 35363 8067
rect 35311 7999 35319 8033
rect 35353 7999 35363 8033
rect 35311 7965 35363 7999
rect 35311 7931 35319 7965
rect 35353 7931 35363 7965
rect 35311 7919 35363 7931
rect 35393 8101 35447 8119
rect 35393 8067 35403 8101
rect 35437 8067 35447 8101
rect 35393 8033 35447 8067
rect 35393 7999 35403 8033
rect 35437 7999 35447 8033
rect 35393 7965 35447 7999
rect 35393 7931 35403 7965
rect 35437 7931 35447 7965
rect 35393 7919 35447 7931
rect 35477 8033 35531 8119
rect 35477 7999 35487 8033
rect 35521 7999 35531 8033
rect 35477 7965 35531 7999
rect 35477 7931 35487 7965
rect 35521 7931 35531 7965
rect 35477 7919 35531 7931
rect 35561 8101 35615 8119
rect 35561 8067 35571 8101
rect 35605 8067 35615 8101
rect 35561 8033 35615 8067
rect 35561 7999 35571 8033
rect 35605 7999 35615 8033
rect 35561 7965 35615 7999
rect 35561 7931 35571 7965
rect 35605 7931 35615 7965
rect 35561 7919 35615 7931
rect 35645 7965 35697 8119
rect 35645 7931 35655 7965
rect 35689 7931 35697 7965
rect 35645 7919 35697 7931
rect 30579 7805 30631 7819
rect 30579 7771 30587 7805
rect 30621 7771 30631 7805
rect 30579 7737 30631 7771
rect 30579 7703 30587 7737
rect 30621 7703 30631 7737
rect 30579 7691 30631 7703
rect 30661 7789 30715 7819
rect 30661 7755 30671 7789
rect 30705 7755 30715 7789
rect 30661 7691 30715 7755
rect 30745 7805 30797 7819
rect 30745 7771 30755 7805
rect 30789 7771 30797 7805
rect 30745 7737 30797 7771
rect 30851 7813 30903 7825
rect 30851 7779 30859 7813
rect 30893 7779 30903 7813
rect 30851 7741 30903 7779
rect 30933 7805 30988 7825
rect 30933 7771 30943 7805
rect 30977 7771 30988 7805
rect 30933 7741 30988 7771
rect 31018 7800 31083 7825
rect 31018 7766 31035 7800
rect 31069 7766 31083 7800
rect 31018 7741 31083 7766
rect 31113 7741 31186 7825
rect 31216 7813 31318 7825
rect 31216 7779 31274 7813
rect 31308 7779 31318 7813
rect 31216 7745 31318 7779
rect 31216 7741 31274 7745
rect 30745 7703 30755 7737
rect 30789 7703 30797 7737
rect 30745 7691 30797 7703
rect 31231 7711 31274 7741
rect 31308 7711 31318 7745
rect 31231 7675 31318 7711
rect 31348 7805 31413 7825
rect 31348 7771 31358 7805
rect 31392 7771 31413 7805
rect 31348 7741 31413 7771
rect 31443 7795 31497 7825
rect 31443 7761 31453 7795
rect 31487 7761 31497 7795
rect 31443 7741 31497 7761
rect 31527 7741 31611 7825
rect 31641 7805 31694 7825
rect 31641 7771 31652 7805
rect 31686 7771 31694 7805
rect 31641 7741 31694 7771
rect 31768 7813 31822 7825
rect 31768 7779 31776 7813
rect 31810 7779 31822 7813
rect 31768 7742 31822 7779
rect 31348 7675 31398 7741
rect 31768 7708 31776 7742
rect 31810 7708 31822 7742
rect 31768 7671 31822 7708
rect 31768 7637 31776 7671
rect 31810 7637 31822 7671
rect 31768 7625 31822 7637
rect 31852 7783 31906 7825
rect 31852 7749 31862 7783
rect 31896 7749 31906 7783
rect 31852 7703 31906 7749
rect 31852 7669 31862 7703
rect 31896 7669 31906 7703
rect 31852 7625 31906 7669
rect 31936 7807 31988 7825
rect 31936 7773 31946 7807
rect 31980 7773 31988 7807
rect 31936 7739 31988 7773
rect 31936 7705 31946 7739
rect 31980 7705 31988 7739
rect 31936 7671 31988 7705
rect 32042 7813 32094 7825
rect 32042 7779 32050 7813
rect 32084 7779 32094 7813
rect 32042 7745 32094 7779
rect 32042 7711 32050 7745
rect 32084 7711 32094 7745
rect 32042 7697 32094 7711
rect 32124 7813 32191 7825
rect 32124 7779 32147 7813
rect 32181 7779 32191 7813
rect 32124 7745 32191 7779
rect 32124 7711 32147 7745
rect 32181 7711 32191 7745
rect 32124 7697 32191 7711
rect 31936 7637 31946 7671
rect 31980 7637 31988 7671
rect 31936 7625 31988 7637
rect 32139 7677 32191 7697
rect 32139 7643 32147 7677
rect 32181 7643 32191 7677
rect 32139 7625 32191 7643
rect 32221 7813 32273 7825
rect 32221 7779 32231 7813
rect 32265 7779 32273 7813
rect 32221 7742 32273 7779
rect 32221 7708 32231 7742
rect 32265 7708 32273 7742
rect 32221 7671 32273 7708
rect 32221 7637 32231 7671
rect 32265 7637 32273 7671
rect 32221 7625 32273 7637
rect 32368 7813 32420 7825
rect 32368 7779 32376 7813
rect 32410 7779 32420 7813
rect 32368 7745 32420 7779
rect 32368 7711 32376 7745
rect 32410 7711 32420 7745
rect 32368 7677 32420 7711
rect 32368 7643 32376 7677
rect 32410 7643 32420 7677
rect 32368 7625 32420 7643
rect 32450 7813 32502 7825
rect 32450 7779 32460 7813
rect 32494 7779 32502 7813
rect 32450 7745 32502 7779
rect 32450 7711 32460 7745
rect 32494 7711 32502 7745
rect 32450 7677 32502 7711
rect 32450 7643 32460 7677
rect 32494 7643 32502 7677
rect 32450 7625 32502 7643
rect 32613 7813 32665 7825
rect 32613 7779 32621 7813
rect 32655 7779 32665 7813
rect 32613 7745 32665 7779
rect 32613 7711 32621 7745
rect 32655 7711 32665 7745
rect 32613 7677 32665 7711
rect 32613 7643 32621 7677
rect 32655 7643 32665 7677
rect 32613 7625 32665 7643
rect 32695 7813 32749 7825
rect 32695 7779 32705 7813
rect 32739 7779 32749 7813
rect 32695 7745 32749 7779
rect 32695 7711 32705 7745
rect 32739 7711 32749 7745
rect 32695 7677 32749 7711
rect 32695 7643 32705 7677
rect 32739 7643 32749 7677
rect 32695 7625 32749 7643
rect 32779 7813 32833 7825
rect 32779 7779 32789 7813
rect 32823 7779 32833 7813
rect 32779 7745 32833 7779
rect 32779 7711 32789 7745
rect 32823 7711 32833 7745
rect 32779 7625 32833 7711
rect 32863 7813 32917 7825
rect 32863 7779 32873 7813
rect 32907 7779 32917 7813
rect 32863 7745 32917 7779
rect 32863 7711 32873 7745
rect 32907 7711 32917 7745
rect 32863 7677 32917 7711
rect 32863 7643 32873 7677
rect 32907 7643 32917 7677
rect 32863 7625 32917 7643
rect 32947 7813 32999 7825
rect 32947 7779 32957 7813
rect 32991 7779 32999 7813
rect 32947 7625 32999 7779
rect 33277 7805 33329 7819
rect 33277 7771 33285 7805
rect 33319 7771 33329 7805
rect 33277 7737 33329 7771
rect 33277 7703 33285 7737
rect 33319 7703 33329 7737
rect 33277 7691 33329 7703
rect 33359 7789 33413 7819
rect 33359 7755 33369 7789
rect 33403 7755 33413 7789
rect 33359 7691 33413 7755
rect 33443 7805 33495 7819
rect 33443 7771 33453 7805
rect 33487 7771 33495 7805
rect 33443 7737 33495 7771
rect 33549 7813 33601 7825
rect 33549 7779 33557 7813
rect 33591 7779 33601 7813
rect 33549 7741 33601 7779
rect 33631 7805 33686 7825
rect 33631 7771 33641 7805
rect 33675 7771 33686 7805
rect 33631 7741 33686 7771
rect 33716 7800 33781 7825
rect 33716 7766 33733 7800
rect 33767 7766 33781 7800
rect 33716 7741 33781 7766
rect 33811 7741 33884 7825
rect 33914 7813 34016 7825
rect 33914 7779 33972 7813
rect 34006 7779 34016 7813
rect 33914 7745 34016 7779
rect 33914 7741 33972 7745
rect 33443 7703 33453 7737
rect 33487 7703 33495 7737
rect 33443 7691 33495 7703
rect 33929 7711 33972 7741
rect 34006 7711 34016 7745
rect 33929 7675 34016 7711
rect 34046 7805 34111 7825
rect 34046 7771 34056 7805
rect 34090 7771 34111 7805
rect 34046 7741 34111 7771
rect 34141 7795 34195 7825
rect 34141 7761 34151 7795
rect 34185 7761 34195 7795
rect 34141 7741 34195 7761
rect 34225 7741 34309 7825
rect 34339 7805 34392 7825
rect 34339 7771 34350 7805
rect 34384 7771 34392 7805
rect 34339 7741 34392 7771
rect 34466 7813 34520 7825
rect 34466 7779 34474 7813
rect 34508 7779 34520 7813
rect 34466 7742 34520 7779
rect 34046 7675 34096 7741
rect 34466 7708 34474 7742
rect 34508 7708 34520 7742
rect 34466 7671 34520 7708
rect 34466 7637 34474 7671
rect 34508 7637 34520 7671
rect 34466 7625 34520 7637
rect 34550 7783 34604 7825
rect 34550 7749 34560 7783
rect 34594 7749 34604 7783
rect 34550 7703 34604 7749
rect 34550 7669 34560 7703
rect 34594 7669 34604 7703
rect 34550 7625 34604 7669
rect 34634 7807 34686 7825
rect 34634 7773 34644 7807
rect 34678 7773 34686 7807
rect 34634 7739 34686 7773
rect 34634 7705 34644 7739
rect 34678 7705 34686 7739
rect 34634 7671 34686 7705
rect 34740 7813 34792 7825
rect 34740 7779 34748 7813
rect 34782 7779 34792 7813
rect 34740 7745 34792 7779
rect 34740 7711 34748 7745
rect 34782 7711 34792 7745
rect 34740 7697 34792 7711
rect 34822 7813 34889 7825
rect 34822 7779 34845 7813
rect 34879 7779 34889 7813
rect 34822 7745 34889 7779
rect 34822 7711 34845 7745
rect 34879 7711 34889 7745
rect 34822 7697 34889 7711
rect 34634 7637 34644 7671
rect 34678 7637 34686 7671
rect 34634 7625 34686 7637
rect 34837 7677 34889 7697
rect 34837 7643 34845 7677
rect 34879 7643 34889 7677
rect 34837 7625 34889 7643
rect 34919 7813 34971 7825
rect 34919 7779 34929 7813
rect 34963 7779 34971 7813
rect 34919 7742 34971 7779
rect 34919 7708 34929 7742
rect 34963 7708 34971 7742
rect 34919 7671 34971 7708
rect 34919 7637 34929 7671
rect 34963 7637 34971 7671
rect 34919 7625 34971 7637
rect 35066 7813 35118 7825
rect 35066 7779 35074 7813
rect 35108 7779 35118 7813
rect 35066 7745 35118 7779
rect 35066 7711 35074 7745
rect 35108 7711 35118 7745
rect 35066 7677 35118 7711
rect 35066 7643 35074 7677
rect 35108 7643 35118 7677
rect 35066 7625 35118 7643
rect 35148 7813 35200 7825
rect 35148 7779 35158 7813
rect 35192 7779 35200 7813
rect 35148 7745 35200 7779
rect 35148 7711 35158 7745
rect 35192 7711 35200 7745
rect 35148 7677 35200 7711
rect 35148 7643 35158 7677
rect 35192 7643 35200 7677
rect 35148 7625 35200 7643
rect 35311 7813 35363 7825
rect 35311 7779 35319 7813
rect 35353 7779 35363 7813
rect 35311 7745 35363 7779
rect 35311 7711 35319 7745
rect 35353 7711 35363 7745
rect 35311 7677 35363 7711
rect 35311 7643 35319 7677
rect 35353 7643 35363 7677
rect 35311 7625 35363 7643
rect 35393 7813 35447 7825
rect 35393 7779 35403 7813
rect 35437 7779 35447 7813
rect 35393 7745 35447 7779
rect 35393 7711 35403 7745
rect 35437 7711 35447 7745
rect 35393 7677 35447 7711
rect 35393 7643 35403 7677
rect 35437 7643 35447 7677
rect 35393 7625 35447 7643
rect 35477 7813 35531 7825
rect 35477 7779 35487 7813
rect 35521 7779 35531 7813
rect 35477 7745 35531 7779
rect 35477 7711 35487 7745
rect 35521 7711 35531 7745
rect 35477 7625 35531 7711
rect 35561 7813 35615 7825
rect 35561 7779 35571 7813
rect 35605 7779 35615 7813
rect 35561 7745 35615 7779
rect 35561 7711 35571 7745
rect 35605 7711 35615 7745
rect 35561 7677 35615 7711
rect 35561 7643 35571 7677
rect 35605 7643 35615 7677
rect 35561 7625 35615 7643
rect 35645 7813 35697 7825
rect 35645 7779 35655 7813
rect 35689 7779 35697 7813
rect 35645 7625 35697 7779
rect 30579 6953 30631 6965
rect 30579 6919 30587 6953
rect 30621 6919 30631 6953
rect 30579 6885 30631 6919
rect 30579 6851 30587 6885
rect 30621 6851 30631 6885
rect 30579 6837 30631 6851
rect 30661 6901 30715 6965
rect 30661 6867 30671 6901
rect 30705 6867 30715 6901
rect 30661 6837 30715 6867
rect 30745 6953 30797 6965
rect 30745 6919 30755 6953
rect 30789 6919 30797 6953
rect 30745 6885 30797 6919
rect 31768 7019 31822 7031
rect 31231 6945 31318 6981
rect 31231 6915 31274 6945
rect 30745 6851 30755 6885
rect 30789 6851 30797 6885
rect 30745 6837 30797 6851
rect 30851 6877 30903 6915
rect 30851 6843 30859 6877
rect 30893 6843 30903 6877
rect 30851 6831 30903 6843
rect 30933 6885 30988 6915
rect 30933 6851 30943 6885
rect 30977 6851 30988 6885
rect 30933 6831 30988 6851
rect 31018 6890 31083 6915
rect 31018 6856 31035 6890
rect 31069 6856 31083 6890
rect 31018 6831 31083 6856
rect 31113 6831 31186 6915
rect 31216 6911 31274 6915
rect 31308 6911 31318 6945
rect 31216 6877 31318 6911
rect 31216 6843 31274 6877
rect 31308 6843 31318 6877
rect 31216 6831 31318 6843
rect 31348 6915 31398 6981
rect 31768 6985 31776 7019
rect 31810 6985 31822 7019
rect 31768 6948 31822 6985
rect 31348 6885 31413 6915
rect 31348 6851 31358 6885
rect 31392 6851 31413 6885
rect 31348 6831 31413 6851
rect 31443 6895 31497 6915
rect 31443 6861 31453 6895
rect 31487 6861 31497 6895
rect 31443 6831 31497 6861
rect 31527 6831 31611 6915
rect 31641 6885 31694 6915
rect 31641 6851 31652 6885
rect 31686 6851 31694 6885
rect 31641 6831 31694 6851
rect 31768 6914 31776 6948
rect 31810 6914 31822 6948
rect 31768 6877 31822 6914
rect 31768 6843 31776 6877
rect 31810 6843 31822 6877
rect 31768 6831 31822 6843
rect 31852 6987 31906 7031
rect 31852 6953 31862 6987
rect 31896 6953 31906 6987
rect 31852 6907 31906 6953
rect 31852 6873 31862 6907
rect 31896 6873 31906 6907
rect 31852 6831 31906 6873
rect 31936 7019 31988 7031
rect 31936 6985 31946 7019
rect 31980 6985 31988 7019
rect 31936 6951 31988 6985
rect 32139 7013 32191 7031
rect 32139 6979 32147 7013
rect 32181 6979 32191 7013
rect 32139 6959 32191 6979
rect 31936 6917 31946 6951
rect 31980 6917 31988 6951
rect 31936 6883 31988 6917
rect 31936 6849 31946 6883
rect 31980 6849 31988 6883
rect 31936 6831 31988 6849
rect 32042 6945 32094 6959
rect 32042 6911 32050 6945
rect 32084 6911 32094 6945
rect 32042 6877 32094 6911
rect 32042 6843 32050 6877
rect 32084 6843 32094 6877
rect 32042 6831 32094 6843
rect 32124 6945 32191 6959
rect 32124 6911 32147 6945
rect 32181 6911 32191 6945
rect 32124 6877 32191 6911
rect 32124 6843 32147 6877
rect 32181 6843 32191 6877
rect 32124 6831 32191 6843
rect 32221 7019 32273 7031
rect 32221 6985 32231 7019
rect 32265 6985 32273 7019
rect 32221 6948 32273 6985
rect 32221 6914 32231 6948
rect 32265 6914 32273 6948
rect 32221 6877 32273 6914
rect 32221 6843 32231 6877
rect 32265 6843 32273 6877
rect 32221 6831 32273 6843
rect 32368 7013 32420 7031
rect 32368 6979 32376 7013
rect 32410 6979 32420 7013
rect 32368 6945 32420 6979
rect 32368 6911 32376 6945
rect 32410 6911 32420 6945
rect 32368 6877 32420 6911
rect 32368 6843 32376 6877
rect 32410 6843 32420 6877
rect 32368 6831 32420 6843
rect 32450 7013 32502 7031
rect 32450 6979 32460 7013
rect 32494 6979 32502 7013
rect 32450 6945 32502 6979
rect 32450 6911 32460 6945
rect 32494 6911 32502 6945
rect 32450 6877 32502 6911
rect 32450 6843 32460 6877
rect 32494 6843 32502 6877
rect 32450 6831 32502 6843
rect 32613 7013 32665 7031
rect 32613 6979 32621 7013
rect 32655 6979 32665 7013
rect 32613 6945 32665 6979
rect 32613 6911 32621 6945
rect 32655 6911 32665 6945
rect 32613 6877 32665 6911
rect 32613 6843 32621 6877
rect 32655 6843 32665 6877
rect 32613 6831 32665 6843
rect 32695 7013 32749 7031
rect 32695 6979 32705 7013
rect 32739 6979 32749 7013
rect 32695 6945 32749 6979
rect 32695 6911 32705 6945
rect 32739 6911 32749 6945
rect 32695 6877 32749 6911
rect 32695 6843 32705 6877
rect 32739 6843 32749 6877
rect 32695 6831 32749 6843
rect 32779 6945 32833 7031
rect 32779 6911 32789 6945
rect 32823 6911 32833 6945
rect 32779 6877 32833 6911
rect 32779 6843 32789 6877
rect 32823 6843 32833 6877
rect 32779 6831 32833 6843
rect 32863 7013 32917 7031
rect 32863 6979 32873 7013
rect 32907 6979 32917 7013
rect 32863 6945 32917 6979
rect 32863 6911 32873 6945
rect 32907 6911 32917 6945
rect 32863 6877 32917 6911
rect 32863 6843 32873 6877
rect 32907 6843 32917 6877
rect 32863 6831 32917 6843
rect 32947 6877 32999 7031
rect 32947 6843 32957 6877
rect 32991 6843 32999 6877
rect 32947 6831 32999 6843
rect 33277 6953 33329 6965
rect 33277 6919 33285 6953
rect 33319 6919 33329 6953
rect 33277 6885 33329 6919
rect 33277 6851 33285 6885
rect 33319 6851 33329 6885
rect 33277 6837 33329 6851
rect 33359 6901 33413 6965
rect 33359 6867 33369 6901
rect 33403 6867 33413 6901
rect 33359 6837 33413 6867
rect 33443 6953 33495 6965
rect 33443 6919 33453 6953
rect 33487 6919 33495 6953
rect 33443 6885 33495 6919
rect 34466 7019 34520 7031
rect 33929 6945 34016 6981
rect 33929 6915 33972 6945
rect 33443 6851 33453 6885
rect 33487 6851 33495 6885
rect 33443 6837 33495 6851
rect 33549 6877 33601 6915
rect 33549 6843 33557 6877
rect 33591 6843 33601 6877
rect 33549 6831 33601 6843
rect 33631 6885 33686 6915
rect 33631 6851 33641 6885
rect 33675 6851 33686 6885
rect 33631 6831 33686 6851
rect 33716 6890 33781 6915
rect 33716 6856 33733 6890
rect 33767 6856 33781 6890
rect 33716 6831 33781 6856
rect 33811 6831 33884 6915
rect 33914 6911 33972 6915
rect 34006 6911 34016 6945
rect 33914 6877 34016 6911
rect 33914 6843 33972 6877
rect 34006 6843 34016 6877
rect 33914 6831 34016 6843
rect 34046 6915 34096 6981
rect 34466 6985 34474 7019
rect 34508 6985 34520 7019
rect 34466 6948 34520 6985
rect 34046 6885 34111 6915
rect 34046 6851 34056 6885
rect 34090 6851 34111 6885
rect 34046 6831 34111 6851
rect 34141 6895 34195 6915
rect 34141 6861 34151 6895
rect 34185 6861 34195 6895
rect 34141 6831 34195 6861
rect 34225 6831 34309 6915
rect 34339 6885 34392 6915
rect 34339 6851 34350 6885
rect 34384 6851 34392 6885
rect 34339 6831 34392 6851
rect 34466 6914 34474 6948
rect 34508 6914 34520 6948
rect 34466 6877 34520 6914
rect 34466 6843 34474 6877
rect 34508 6843 34520 6877
rect 34466 6831 34520 6843
rect 34550 6987 34604 7031
rect 34550 6953 34560 6987
rect 34594 6953 34604 6987
rect 34550 6907 34604 6953
rect 34550 6873 34560 6907
rect 34594 6873 34604 6907
rect 34550 6831 34604 6873
rect 34634 7019 34686 7031
rect 34634 6985 34644 7019
rect 34678 6985 34686 7019
rect 34634 6951 34686 6985
rect 34837 7013 34889 7031
rect 34837 6979 34845 7013
rect 34879 6979 34889 7013
rect 34837 6959 34889 6979
rect 34634 6917 34644 6951
rect 34678 6917 34686 6951
rect 34634 6883 34686 6917
rect 34634 6849 34644 6883
rect 34678 6849 34686 6883
rect 34634 6831 34686 6849
rect 34740 6945 34792 6959
rect 34740 6911 34748 6945
rect 34782 6911 34792 6945
rect 34740 6877 34792 6911
rect 34740 6843 34748 6877
rect 34782 6843 34792 6877
rect 34740 6831 34792 6843
rect 34822 6945 34889 6959
rect 34822 6911 34845 6945
rect 34879 6911 34889 6945
rect 34822 6877 34889 6911
rect 34822 6843 34845 6877
rect 34879 6843 34889 6877
rect 34822 6831 34889 6843
rect 34919 7019 34971 7031
rect 34919 6985 34929 7019
rect 34963 6985 34971 7019
rect 34919 6948 34971 6985
rect 34919 6914 34929 6948
rect 34963 6914 34971 6948
rect 34919 6877 34971 6914
rect 34919 6843 34929 6877
rect 34963 6843 34971 6877
rect 34919 6831 34971 6843
rect 35066 7013 35118 7031
rect 35066 6979 35074 7013
rect 35108 6979 35118 7013
rect 35066 6945 35118 6979
rect 35066 6911 35074 6945
rect 35108 6911 35118 6945
rect 35066 6877 35118 6911
rect 35066 6843 35074 6877
rect 35108 6843 35118 6877
rect 35066 6831 35118 6843
rect 35148 7013 35200 7031
rect 35148 6979 35158 7013
rect 35192 6979 35200 7013
rect 35148 6945 35200 6979
rect 35148 6911 35158 6945
rect 35192 6911 35200 6945
rect 35148 6877 35200 6911
rect 35148 6843 35158 6877
rect 35192 6843 35200 6877
rect 35148 6831 35200 6843
rect 35311 7013 35363 7031
rect 35311 6979 35319 7013
rect 35353 6979 35363 7013
rect 35311 6945 35363 6979
rect 35311 6911 35319 6945
rect 35353 6911 35363 6945
rect 35311 6877 35363 6911
rect 35311 6843 35319 6877
rect 35353 6843 35363 6877
rect 35311 6831 35363 6843
rect 35393 7013 35447 7031
rect 35393 6979 35403 7013
rect 35437 6979 35447 7013
rect 35393 6945 35447 6979
rect 35393 6911 35403 6945
rect 35437 6911 35447 6945
rect 35393 6877 35447 6911
rect 35393 6843 35403 6877
rect 35437 6843 35447 6877
rect 35393 6831 35447 6843
rect 35477 6945 35531 7031
rect 35477 6911 35487 6945
rect 35521 6911 35531 6945
rect 35477 6877 35531 6911
rect 35477 6843 35487 6877
rect 35521 6843 35531 6877
rect 35477 6831 35531 6843
rect 35561 7013 35615 7031
rect 35561 6979 35571 7013
rect 35605 6979 35615 7013
rect 35561 6945 35615 6979
rect 35561 6911 35571 6945
rect 35605 6911 35615 6945
rect 35561 6877 35615 6911
rect 35561 6843 35571 6877
rect 35605 6843 35615 6877
rect 35561 6831 35615 6843
rect 35645 6877 35697 7031
rect 35645 6843 35655 6877
rect 35689 6843 35697 6877
rect 35645 6831 35697 6843
rect 30579 6717 30631 6731
rect 30579 6683 30587 6717
rect 30621 6683 30631 6717
rect 30579 6649 30631 6683
rect 30579 6615 30587 6649
rect 30621 6615 30631 6649
rect 30579 6603 30631 6615
rect 30661 6701 30715 6731
rect 30661 6667 30671 6701
rect 30705 6667 30715 6701
rect 30661 6603 30715 6667
rect 30745 6717 30797 6731
rect 30745 6683 30755 6717
rect 30789 6683 30797 6717
rect 30745 6649 30797 6683
rect 30851 6725 30903 6737
rect 30851 6691 30859 6725
rect 30893 6691 30903 6725
rect 30851 6653 30903 6691
rect 30933 6717 30988 6737
rect 30933 6683 30943 6717
rect 30977 6683 30988 6717
rect 30933 6653 30988 6683
rect 31018 6712 31083 6737
rect 31018 6678 31035 6712
rect 31069 6678 31083 6712
rect 31018 6653 31083 6678
rect 31113 6653 31186 6737
rect 31216 6725 31318 6737
rect 31216 6691 31274 6725
rect 31308 6691 31318 6725
rect 31216 6657 31318 6691
rect 31216 6653 31274 6657
rect 30745 6615 30755 6649
rect 30789 6615 30797 6649
rect 30745 6603 30797 6615
rect 31231 6623 31274 6653
rect 31308 6623 31318 6657
rect 31231 6587 31318 6623
rect 31348 6717 31413 6737
rect 31348 6683 31358 6717
rect 31392 6683 31413 6717
rect 31348 6653 31413 6683
rect 31443 6707 31497 6737
rect 31443 6673 31453 6707
rect 31487 6673 31497 6707
rect 31443 6653 31497 6673
rect 31527 6653 31611 6737
rect 31641 6717 31694 6737
rect 31641 6683 31652 6717
rect 31686 6683 31694 6717
rect 31641 6653 31694 6683
rect 31768 6725 31822 6737
rect 31768 6691 31776 6725
rect 31810 6691 31822 6725
rect 31768 6654 31822 6691
rect 31348 6587 31398 6653
rect 31768 6620 31776 6654
rect 31810 6620 31822 6654
rect 31768 6583 31822 6620
rect 31768 6549 31776 6583
rect 31810 6549 31822 6583
rect 31768 6537 31822 6549
rect 31852 6695 31906 6737
rect 31852 6661 31862 6695
rect 31896 6661 31906 6695
rect 31852 6615 31906 6661
rect 31852 6581 31862 6615
rect 31896 6581 31906 6615
rect 31852 6537 31906 6581
rect 31936 6719 31988 6737
rect 31936 6685 31946 6719
rect 31980 6685 31988 6719
rect 31936 6651 31988 6685
rect 31936 6617 31946 6651
rect 31980 6617 31988 6651
rect 31936 6583 31988 6617
rect 32042 6725 32094 6737
rect 32042 6691 32050 6725
rect 32084 6691 32094 6725
rect 32042 6657 32094 6691
rect 32042 6623 32050 6657
rect 32084 6623 32094 6657
rect 32042 6609 32094 6623
rect 32124 6725 32191 6737
rect 32124 6691 32147 6725
rect 32181 6691 32191 6725
rect 32124 6657 32191 6691
rect 32124 6623 32147 6657
rect 32181 6623 32191 6657
rect 32124 6609 32191 6623
rect 31936 6549 31946 6583
rect 31980 6549 31988 6583
rect 31936 6537 31988 6549
rect 32139 6589 32191 6609
rect 32139 6555 32147 6589
rect 32181 6555 32191 6589
rect 32139 6537 32191 6555
rect 32221 6725 32273 6737
rect 32221 6691 32231 6725
rect 32265 6691 32273 6725
rect 32221 6654 32273 6691
rect 32221 6620 32231 6654
rect 32265 6620 32273 6654
rect 32221 6583 32273 6620
rect 32221 6549 32231 6583
rect 32265 6549 32273 6583
rect 32221 6537 32273 6549
rect 32368 6725 32420 6737
rect 32368 6691 32376 6725
rect 32410 6691 32420 6725
rect 32368 6657 32420 6691
rect 32368 6623 32376 6657
rect 32410 6623 32420 6657
rect 32368 6589 32420 6623
rect 32368 6555 32376 6589
rect 32410 6555 32420 6589
rect 32368 6537 32420 6555
rect 32450 6725 32502 6737
rect 32450 6691 32460 6725
rect 32494 6691 32502 6725
rect 32450 6657 32502 6691
rect 32450 6623 32460 6657
rect 32494 6623 32502 6657
rect 32450 6589 32502 6623
rect 32450 6555 32460 6589
rect 32494 6555 32502 6589
rect 32450 6537 32502 6555
rect 32613 6725 32665 6737
rect 32613 6691 32621 6725
rect 32655 6691 32665 6725
rect 32613 6657 32665 6691
rect 32613 6623 32621 6657
rect 32655 6623 32665 6657
rect 32613 6589 32665 6623
rect 32613 6555 32621 6589
rect 32655 6555 32665 6589
rect 32613 6537 32665 6555
rect 32695 6725 32749 6737
rect 32695 6691 32705 6725
rect 32739 6691 32749 6725
rect 32695 6657 32749 6691
rect 32695 6623 32705 6657
rect 32739 6623 32749 6657
rect 32695 6589 32749 6623
rect 32695 6555 32705 6589
rect 32739 6555 32749 6589
rect 32695 6537 32749 6555
rect 32779 6725 32833 6737
rect 32779 6691 32789 6725
rect 32823 6691 32833 6725
rect 32779 6657 32833 6691
rect 32779 6623 32789 6657
rect 32823 6623 32833 6657
rect 32779 6537 32833 6623
rect 32863 6725 32917 6737
rect 32863 6691 32873 6725
rect 32907 6691 32917 6725
rect 32863 6657 32917 6691
rect 32863 6623 32873 6657
rect 32907 6623 32917 6657
rect 32863 6589 32917 6623
rect 32863 6555 32873 6589
rect 32907 6555 32917 6589
rect 32863 6537 32917 6555
rect 32947 6725 32999 6737
rect 32947 6691 32957 6725
rect 32991 6691 32999 6725
rect 32947 6537 32999 6691
rect 33277 6717 33329 6731
rect 33277 6683 33285 6717
rect 33319 6683 33329 6717
rect 33277 6649 33329 6683
rect 33277 6615 33285 6649
rect 33319 6615 33329 6649
rect 33277 6603 33329 6615
rect 33359 6701 33413 6731
rect 33359 6667 33369 6701
rect 33403 6667 33413 6701
rect 33359 6603 33413 6667
rect 33443 6717 33495 6731
rect 33443 6683 33453 6717
rect 33487 6683 33495 6717
rect 33443 6649 33495 6683
rect 33549 6725 33601 6737
rect 33549 6691 33557 6725
rect 33591 6691 33601 6725
rect 33549 6653 33601 6691
rect 33631 6717 33686 6737
rect 33631 6683 33641 6717
rect 33675 6683 33686 6717
rect 33631 6653 33686 6683
rect 33716 6712 33781 6737
rect 33716 6678 33733 6712
rect 33767 6678 33781 6712
rect 33716 6653 33781 6678
rect 33811 6653 33884 6737
rect 33914 6725 34016 6737
rect 33914 6691 33972 6725
rect 34006 6691 34016 6725
rect 33914 6657 34016 6691
rect 33914 6653 33972 6657
rect 33443 6615 33453 6649
rect 33487 6615 33495 6649
rect 33443 6603 33495 6615
rect 33929 6623 33972 6653
rect 34006 6623 34016 6657
rect 33929 6587 34016 6623
rect 34046 6717 34111 6737
rect 34046 6683 34056 6717
rect 34090 6683 34111 6717
rect 34046 6653 34111 6683
rect 34141 6707 34195 6737
rect 34141 6673 34151 6707
rect 34185 6673 34195 6707
rect 34141 6653 34195 6673
rect 34225 6653 34309 6737
rect 34339 6717 34392 6737
rect 34339 6683 34350 6717
rect 34384 6683 34392 6717
rect 34339 6653 34392 6683
rect 34466 6725 34520 6737
rect 34466 6691 34474 6725
rect 34508 6691 34520 6725
rect 34466 6654 34520 6691
rect 34046 6587 34096 6653
rect 34466 6620 34474 6654
rect 34508 6620 34520 6654
rect 34466 6583 34520 6620
rect 34466 6549 34474 6583
rect 34508 6549 34520 6583
rect 34466 6537 34520 6549
rect 34550 6695 34604 6737
rect 34550 6661 34560 6695
rect 34594 6661 34604 6695
rect 34550 6615 34604 6661
rect 34550 6581 34560 6615
rect 34594 6581 34604 6615
rect 34550 6537 34604 6581
rect 34634 6719 34686 6737
rect 34634 6685 34644 6719
rect 34678 6685 34686 6719
rect 34634 6651 34686 6685
rect 34634 6617 34644 6651
rect 34678 6617 34686 6651
rect 34634 6583 34686 6617
rect 34740 6725 34792 6737
rect 34740 6691 34748 6725
rect 34782 6691 34792 6725
rect 34740 6657 34792 6691
rect 34740 6623 34748 6657
rect 34782 6623 34792 6657
rect 34740 6609 34792 6623
rect 34822 6725 34889 6737
rect 34822 6691 34845 6725
rect 34879 6691 34889 6725
rect 34822 6657 34889 6691
rect 34822 6623 34845 6657
rect 34879 6623 34889 6657
rect 34822 6609 34889 6623
rect 34634 6549 34644 6583
rect 34678 6549 34686 6583
rect 34634 6537 34686 6549
rect 34837 6589 34889 6609
rect 34837 6555 34845 6589
rect 34879 6555 34889 6589
rect 34837 6537 34889 6555
rect 34919 6725 34971 6737
rect 34919 6691 34929 6725
rect 34963 6691 34971 6725
rect 34919 6654 34971 6691
rect 34919 6620 34929 6654
rect 34963 6620 34971 6654
rect 34919 6583 34971 6620
rect 34919 6549 34929 6583
rect 34963 6549 34971 6583
rect 34919 6537 34971 6549
rect 35066 6725 35118 6737
rect 35066 6691 35074 6725
rect 35108 6691 35118 6725
rect 35066 6657 35118 6691
rect 35066 6623 35074 6657
rect 35108 6623 35118 6657
rect 35066 6589 35118 6623
rect 35066 6555 35074 6589
rect 35108 6555 35118 6589
rect 35066 6537 35118 6555
rect 35148 6725 35200 6737
rect 35148 6691 35158 6725
rect 35192 6691 35200 6725
rect 35148 6657 35200 6691
rect 35148 6623 35158 6657
rect 35192 6623 35200 6657
rect 35148 6589 35200 6623
rect 35148 6555 35158 6589
rect 35192 6555 35200 6589
rect 35148 6537 35200 6555
rect 35311 6725 35363 6737
rect 35311 6691 35319 6725
rect 35353 6691 35363 6725
rect 35311 6657 35363 6691
rect 35311 6623 35319 6657
rect 35353 6623 35363 6657
rect 35311 6589 35363 6623
rect 35311 6555 35319 6589
rect 35353 6555 35363 6589
rect 35311 6537 35363 6555
rect 35393 6725 35447 6737
rect 35393 6691 35403 6725
rect 35437 6691 35447 6725
rect 35393 6657 35447 6691
rect 35393 6623 35403 6657
rect 35437 6623 35447 6657
rect 35393 6589 35447 6623
rect 35393 6555 35403 6589
rect 35437 6555 35447 6589
rect 35393 6537 35447 6555
rect 35477 6725 35531 6737
rect 35477 6691 35487 6725
rect 35521 6691 35531 6725
rect 35477 6657 35531 6691
rect 35477 6623 35487 6657
rect 35521 6623 35531 6657
rect 35477 6537 35531 6623
rect 35561 6725 35615 6737
rect 35561 6691 35571 6725
rect 35605 6691 35615 6725
rect 35561 6657 35615 6691
rect 35561 6623 35571 6657
rect 35605 6623 35615 6657
rect 35561 6589 35615 6623
rect 35561 6555 35571 6589
rect 35605 6555 35615 6589
rect 35561 6537 35615 6555
rect 35645 6725 35697 6737
rect 35645 6691 35655 6725
rect 35689 6691 35697 6725
rect 35645 6537 35697 6691
rect 30579 5865 30631 5877
rect 30579 5831 30587 5865
rect 30621 5831 30631 5865
rect 30579 5797 30631 5831
rect 30579 5763 30587 5797
rect 30621 5763 30631 5797
rect 30579 5749 30631 5763
rect 30661 5813 30715 5877
rect 30661 5779 30671 5813
rect 30705 5779 30715 5813
rect 30661 5749 30715 5779
rect 30745 5865 30797 5877
rect 30745 5831 30755 5865
rect 30789 5831 30797 5865
rect 30745 5797 30797 5831
rect 31768 5931 31822 5943
rect 31231 5857 31318 5893
rect 31231 5827 31274 5857
rect 30745 5763 30755 5797
rect 30789 5763 30797 5797
rect 30745 5749 30797 5763
rect 30851 5789 30903 5827
rect 30851 5755 30859 5789
rect 30893 5755 30903 5789
rect 30851 5743 30903 5755
rect 30933 5797 30988 5827
rect 30933 5763 30943 5797
rect 30977 5763 30988 5797
rect 30933 5743 30988 5763
rect 31018 5802 31083 5827
rect 31018 5768 31035 5802
rect 31069 5768 31083 5802
rect 31018 5743 31083 5768
rect 31113 5743 31186 5827
rect 31216 5823 31274 5827
rect 31308 5823 31318 5857
rect 31216 5789 31318 5823
rect 31216 5755 31274 5789
rect 31308 5755 31318 5789
rect 31216 5743 31318 5755
rect 31348 5827 31398 5893
rect 31768 5897 31776 5931
rect 31810 5897 31822 5931
rect 31768 5860 31822 5897
rect 31348 5797 31413 5827
rect 31348 5763 31358 5797
rect 31392 5763 31413 5797
rect 31348 5743 31413 5763
rect 31443 5807 31497 5827
rect 31443 5773 31453 5807
rect 31487 5773 31497 5807
rect 31443 5743 31497 5773
rect 31527 5743 31611 5827
rect 31641 5797 31694 5827
rect 31641 5763 31652 5797
rect 31686 5763 31694 5797
rect 31641 5743 31694 5763
rect 31768 5826 31776 5860
rect 31810 5826 31822 5860
rect 31768 5789 31822 5826
rect 31768 5755 31776 5789
rect 31810 5755 31822 5789
rect 31768 5743 31822 5755
rect 31852 5899 31906 5943
rect 31852 5865 31862 5899
rect 31896 5865 31906 5899
rect 31852 5819 31906 5865
rect 31852 5785 31862 5819
rect 31896 5785 31906 5819
rect 31852 5743 31906 5785
rect 31936 5931 31988 5943
rect 31936 5897 31946 5931
rect 31980 5897 31988 5931
rect 31936 5863 31988 5897
rect 32139 5925 32191 5943
rect 32139 5891 32147 5925
rect 32181 5891 32191 5925
rect 32139 5871 32191 5891
rect 31936 5829 31946 5863
rect 31980 5829 31988 5863
rect 31936 5795 31988 5829
rect 31936 5761 31946 5795
rect 31980 5761 31988 5795
rect 31936 5743 31988 5761
rect 32042 5857 32094 5871
rect 32042 5823 32050 5857
rect 32084 5823 32094 5857
rect 32042 5789 32094 5823
rect 32042 5755 32050 5789
rect 32084 5755 32094 5789
rect 32042 5743 32094 5755
rect 32124 5857 32191 5871
rect 32124 5823 32147 5857
rect 32181 5823 32191 5857
rect 32124 5789 32191 5823
rect 32124 5755 32147 5789
rect 32181 5755 32191 5789
rect 32124 5743 32191 5755
rect 32221 5931 32273 5943
rect 32221 5897 32231 5931
rect 32265 5897 32273 5931
rect 32221 5860 32273 5897
rect 32221 5826 32231 5860
rect 32265 5826 32273 5860
rect 32221 5789 32273 5826
rect 32221 5755 32231 5789
rect 32265 5755 32273 5789
rect 32221 5743 32273 5755
rect 32368 5925 32420 5943
rect 32368 5891 32376 5925
rect 32410 5891 32420 5925
rect 32368 5857 32420 5891
rect 32368 5823 32376 5857
rect 32410 5823 32420 5857
rect 32368 5789 32420 5823
rect 32368 5755 32376 5789
rect 32410 5755 32420 5789
rect 32368 5743 32420 5755
rect 32450 5925 32502 5943
rect 32450 5891 32460 5925
rect 32494 5891 32502 5925
rect 32450 5857 32502 5891
rect 32450 5823 32460 5857
rect 32494 5823 32502 5857
rect 32450 5789 32502 5823
rect 32450 5755 32460 5789
rect 32494 5755 32502 5789
rect 32450 5743 32502 5755
rect 32613 5925 32665 5943
rect 32613 5891 32621 5925
rect 32655 5891 32665 5925
rect 32613 5857 32665 5891
rect 32613 5823 32621 5857
rect 32655 5823 32665 5857
rect 32613 5789 32665 5823
rect 32613 5755 32621 5789
rect 32655 5755 32665 5789
rect 32613 5743 32665 5755
rect 32695 5925 32749 5943
rect 32695 5891 32705 5925
rect 32739 5891 32749 5925
rect 32695 5857 32749 5891
rect 32695 5823 32705 5857
rect 32739 5823 32749 5857
rect 32695 5789 32749 5823
rect 32695 5755 32705 5789
rect 32739 5755 32749 5789
rect 32695 5743 32749 5755
rect 32779 5857 32833 5943
rect 32779 5823 32789 5857
rect 32823 5823 32833 5857
rect 32779 5789 32833 5823
rect 32779 5755 32789 5789
rect 32823 5755 32833 5789
rect 32779 5743 32833 5755
rect 32863 5925 32917 5943
rect 32863 5891 32873 5925
rect 32907 5891 32917 5925
rect 32863 5857 32917 5891
rect 32863 5823 32873 5857
rect 32907 5823 32917 5857
rect 32863 5789 32917 5823
rect 32863 5755 32873 5789
rect 32907 5755 32917 5789
rect 32863 5743 32917 5755
rect 32947 5789 32999 5943
rect 32947 5755 32957 5789
rect 32991 5755 32999 5789
rect 32947 5743 32999 5755
rect 33277 5865 33329 5877
rect 33277 5831 33285 5865
rect 33319 5831 33329 5865
rect 33277 5797 33329 5831
rect 33277 5763 33285 5797
rect 33319 5763 33329 5797
rect 33277 5749 33329 5763
rect 33359 5813 33413 5877
rect 33359 5779 33369 5813
rect 33403 5779 33413 5813
rect 33359 5749 33413 5779
rect 33443 5865 33495 5877
rect 33443 5831 33453 5865
rect 33487 5831 33495 5865
rect 33443 5797 33495 5831
rect 34466 5931 34520 5943
rect 33929 5857 34016 5893
rect 33929 5827 33972 5857
rect 33443 5763 33453 5797
rect 33487 5763 33495 5797
rect 33443 5749 33495 5763
rect 33549 5789 33601 5827
rect 33549 5755 33557 5789
rect 33591 5755 33601 5789
rect 33549 5743 33601 5755
rect 33631 5797 33686 5827
rect 33631 5763 33641 5797
rect 33675 5763 33686 5797
rect 33631 5743 33686 5763
rect 33716 5802 33781 5827
rect 33716 5768 33733 5802
rect 33767 5768 33781 5802
rect 33716 5743 33781 5768
rect 33811 5743 33884 5827
rect 33914 5823 33972 5827
rect 34006 5823 34016 5857
rect 33914 5789 34016 5823
rect 33914 5755 33972 5789
rect 34006 5755 34016 5789
rect 33914 5743 34016 5755
rect 34046 5827 34096 5893
rect 34466 5897 34474 5931
rect 34508 5897 34520 5931
rect 34466 5860 34520 5897
rect 34046 5797 34111 5827
rect 34046 5763 34056 5797
rect 34090 5763 34111 5797
rect 34046 5743 34111 5763
rect 34141 5807 34195 5827
rect 34141 5773 34151 5807
rect 34185 5773 34195 5807
rect 34141 5743 34195 5773
rect 34225 5743 34309 5827
rect 34339 5797 34392 5827
rect 34339 5763 34350 5797
rect 34384 5763 34392 5797
rect 34339 5743 34392 5763
rect 34466 5826 34474 5860
rect 34508 5826 34520 5860
rect 34466 5789 34520 5826
rect 34466 5755 34474 5789
rect 34508 5755 34520 5789
rect 34466 5743 34520 5755
rect 34550 5899 34604 5943
rect 34550 5865 34560 5899
rect 34594 5865 34604 5899
rect 34550 5819 34604 5865
rect 34550 5785 34560 5819
rect 34594 5785 34604 5819
rect 34550 5743 34604 5785
rect 34634 5931 34686 5943
rect 34634 5897 34644 5931
rect 34678 5897 34686 5931
rect 34634 5863 34686 5897
rect 34837 5925 34889 5943
rect 34837 5891 34845 5925
rect 34879 5891 34889 5925
rect 34837 5871 34889 5891
rect 34634 5829 34644 5863
rect 34678 5829 34686 5863
rect 34634 5795 34686 5829
rect 34634 5761 34644 5795
rect 34678 5761 34686 5795
rect 34634 5743 34686 5761
rect 34740 5857 34792 5871
rect 34740 5823 34748 5857
rect 34782 5823 34792 5857
rect 34740 5789 34792 5823
rect 34740 5755 34748 5789
rect 34782 5755 34792 5789
rect 34740 5743 34792 5755
rect 34822 5857 34889 5871
rect 34822 5823 34845 5857
rect 34879 5823 34889 5857
rect 34822 5789 34889 5823
rect 34822 5755 34845 5789
rect 34879 5755 34889 5789
rect 34822 5743 34889 5755
rect 34919 5931 34971 5943
rect 34919 5897 34929 5931
rect 34963 5897 34971 5931
rect 34919 5860 34971 5897
rect 34919 5826 34929 5860
rect 34963 5826 34971 5860
rect 34919 5789 34971 5826
rect 34919 5755 34929 5789
rect 34963 5755 34971 5789
rect 34919 5743 34971 5755
rect 35066 5925 35118 5943
rect 35066 5891 35074 5925
rect 35108 5891 35118 5925
rect 35066 5857 35118 5891
rect 35066 5823 35074 5857
rect 35108 5823 35118 5857
rect 35066 5789 35118 5823
rect 35066 5755 35074 5789
rect 35108 5755 35118 5789
rect 35066 5743 35118 5755
rect 35148 5925 35200 5943
rect 35148 5891 35158 5925
rect 35192 5891 35200 5925
rect 35148 5857 35200 5891
rect 35148 5823 35158 5857
rect 35192 5823 35200 5857
rect 35148 5789 35200 5823
rect 35148 5755 35158 5789
rect 35192 5755 35200 5789
rect 35148 5743 35200 5755
rect 35311 5925 35363 5943
rect 35311 5891 35319 5925
rect 35353 5891 35363 5925
rect 35311 5857 35363 5891
rect 35311 5823 35319 5857
rect 35353 5823 35363 5857
rect 35311 5789 35363 5823
rect 35311 5755 35319 5789
rect 35353 5755 35363 5789
rect 35311 5743 35363 5755
rect 35393 5925 35447 5943
rect 35393 5891 35403 5925
rect 35437 5891 35447 5925
rect 35393 5857 35447 5891
rect 35393 5823 35403 5857
rect 35437 5823 35447 5857
rect 35393 5789 35447 5823
rect 35393 5755 35403 5789
rect 35437 5755 35447 5789
rect 35393 5743 35447 5755
rect 35477 5857 35531 5943
rect 35477 5823 35487 5857
rect 35521 5823 35531 5857
rect 35477 5789 35531 5823
rect 35477 5755 35487 5789
rect 35521 5755 35531 5789
rect 35477 5743 35531 5755
rect 35561 5925 35615 5943
rect 35561 5891 35571 5925
rect 35605 5891 35615 5925
rect 35561 5857 35615 5891
rect 35561 5823 35571 5857
rect 35605 5823 35615 5857
rect 35561 5789 35615 5823
rect 35561 5755 35571 5789
rect 35605 5755 35615 5789
rect 35561 5743 35615 5755
rect 35645 5789 35697 5943
rect 35645 5755 35655 5789
rect 35689 5755 35697 5789
rect 35645 5743 35697 5755
rect 9326 2932 9384 2944
rect 9326 1356 9338 2932
rect 9372 1356 9384 2932
rect 9326 1344 9384 1356
rect 9784 2932 9842 2944
rect 9784 1356 9796 2932
rect 9830 1356 9842 2932
rect 9784 1344 9842 1356
rect 10242 2932 10300 2944
rect 10242 1356 10254 2932
rect 10288 1356 10300 2932
rect 10242 1344 10300 1356
rect 10700 2932 10758 2944
rect 10700 1356 10712 2932
rect 10746 1356 10758 2932
rect 10700 1344 10758 1356
rect 11158 2932 11216 2944
rect 11158 1356 11170 2932
rect 11204 1356 11216 2932
rect 11158 1344 11216 1356
rect 11616 2932 11674 2944
rect 11616 1356 11628 2932
rect 11662 1356 11674 2932
rect 11616 1344 11674 1356
rect 12074 2932 12132 2944
rect 12074 1356 12086 2932
rect 12120 1356 12132 2932
rect 12074 1344 12132 1356
rect 12532 2932 12590 2944
rect 12532 1356 12544 2932
rect 12578 1356 12590 2932
rect 12532 1344 12590 1356
rect 12990 2932 13048 2944
rect 12990 1356 13002 2932
rect 13036 1356 13048 2932
rect 12990 1344 13048 1356
rect 13448 2932 13506 2944
rect 13448 1356 13460 2932
rect 13494 1356 13506 2932
rect 13448 1344 13506 1356
rect 13906 2932 13964 2944
rect 13906 1356 13918 2932
rect 13952 1356 13964 2932
rect 13906 1344 13964 1356
rect 14364 2932 14422 2944
rect 14364 1356 14376 2932
rect 14410 1356 14422 2932
rect 14364 1344 14422 1356
rect 14822 2932 14880 2944
rect 14822 1356 14834 2932
rect 14868 1356 14880 2932
rect 14822 1344 14880 1356
rect 15280 2932 15338 2944
rect 15280 1356 15292 2932
rect 15326 1356 15338 2932
rect 15280 1344 15338 1356
rect 15738 2932 15796 2944
rect 15738 1356 15750 2932
rect 15784 1356 15796 2932
rect 15738 1344 15796 1356
rect 16196 2932 16254 2944
rect 16196 1356 16208 2932
rect 16242 1356 16254 2932
rect 16196 1344 16254 1356
rect 16654 2932 16712 2944
rect 16654 1356 16666 2932
rect 16700 1356 16712 2932
rect 16654 1344 16712 1356
rect 17112 2932 17170 2944
rect 17112 1356 17124 2932
rect 17158 1356 17170 2932
rect 17112 1344 17170 1356
rect 17570 2932 17628 2944
rect 17570 1356 17582 2932
rect 17616 1356 17628 2932
rect 17570 1344 17628 1356
rect 8767 267 8825 279
rect 8767 -909 8779 267
rect 8813 -909 8825 267
rect 8767 -921 8825 -909
rect 9225 267 9283 279
rect 9225 -909 9237 267
rect 9271 -909 9283 267
rect 9225 -921 9283 -909
rect 9683 267 9741 279
rect 9683 -909 9695 267
rect 9729 -909 9741 267
rect 9683 -921 9741 -909
rect 10141 267 10199 279
rect 10141 -909 10153 267
rect 10187 -909 10199 267
rect 10141 -921 10199 -909
rect 10599 267 10657 279
rect 10599 -909 10611 267
rect 10645 -909 10657 267
rect 10599 -921 10657 -909
rect 11057 267 11115 279
rect 11057 -909 11069 267
rect 11103 -909 11115 267
rect 11057 -921 11115 -909
rect 11515 267 11573 279
rect 11515 -909 11527 267
rect 11561 -909 11573 267
rect 11515 -921 11573 -909
rect 11973 267 12031 279
rect 11973 -909 11985 267
rect 12019 -909 12031 267
rect 11973 -921 12031 -909
rect 12431 267 12489 279
rect 12431 -909 12443 267
rect 12477 -909 12489 267
rect 12431 -921 12489 -909
rect 12889 267 12947 279
rect 12889 -909 12901 267
rect 12935 -909 12947 267
rect 12889 -921 12947 -909
rect 13347 267 13405 279
rect 13347 -909 13359 267
rect 13393 -909 13405 267
rect 13347 -921 13405 -909
rect 13767 267 13825 279
rect 13767 -909 13779 267
rect 13813 -909 13825 267
rect 13767 -921 13825 -909
rect 14225 267 14283 279
rect 14225 -909 14237 267
rect 14271 -909 14283 267
rect 14225 -921 14283 -909
rect 14683 267 14741 279
rect 14683 -909 14695 267
rect 14729 -909 14741 267
rect 14683 -921 14741 -909
rect 15141 267 15199 279
rect 15141 -909 15153 267
rect 15187 -909 15199 267
rect 15141 -921 15199 -909
rect 15599 267 15657 279
rect 15599 -909 15611 267
rect 15645 -909 15657 267
rect 15599 -921 15657 -909
rect 16057 267 16115 279
rect 16057 -909 16069 267
rect 16103 -909 16115 267
rect 16057 -921 16115 -909
rect 16515 267 16573 279
rect 16515 -909 16527 267
rect 16561 -909 16573 267
rect 16515 -921 16573 -909
rect 16973 267 17031 279
rect 16973 -909 16985 267
rect 17019 -909 17031 267
rect 16973 -921 17031 -909
rect 17431 267 17489 279
rect 17431 -909 17443 267
rect 17477 -909 17489 267
rect 17431 -921 17489 -909
rect 17889 267 17947 279
rect 17889 -909 17901 267
rect 17935 -909 17947 267
rect 17889 -921 17947 -909
rect 18347 267 18405 279
rect 18347 -909 18359 267
rect 18393 -909 18405 267
rect 18347 -921 18405 -909
rect 24326 2932 24384 2944
rect 24326 1356 24338 2932
rect 24372 1356 24384 2932
rect 24326 1344 24384 1356
rect 24784 2932 24842 2944
rect 24784 1356 24796 2932
rect 24830 1356 24842 2932
rect 24784 1344 24842 1356
rect 25242 2932 25300 2944
rect 25242 1356 25254 2932
rect 25288 1356 25300 2932
rect 25242 1344 25300 1356
rect 25700 2932 25758 2944
rect 25700 1356 25712 2932
rect 25746 1356 25758 2932
rect 25700 1344 25758 1356
rect 26158 2932 26216 2944
rect 26158 1356 26170 2932
rect 26204 1356 26216 2932
rect 26158 1344 26216 1356
rect 26616 2932 26674 2944
rect 26616 1356 26628 2932
rect 26662 1356 26674 2932
rect 26616 1344 26674 1356
rect 27074 2932 27132 2944
rect 27074 1356 27086 2932
rect 27120 1356 27132 2932
rect 27074 1344 27132 1356
rect 27532 2932 27590 2944
rect 27532 1356 27544 2932
rect 27578 1356 27590 2932
rect 27532 1344 27590 1356
rect 27990 2932 28048 2944
rect 27990 1356 28002 2932
rect 28036 1356 28048 2932
rect 27990 1344 28048 1356
rect 28448 2932 28506 2944
rect 28448 1356 28460 2932
rect 28494 1356 28506 2932
rect 28448 1344 28506 1356
rect 28906 2932 28964 2944
rect 28906 1356 28918 2932
rect 28952 1356 28964 2932
rect 28906 1344 28964 1356
rect 29364 2932 29422 2944
rect 29364 1356 29376 2932
rect 29410 1356 29422 2932
rect 29364 1344 29422 1356
rect 29822 2932 29880 2944
rect 29822 1356 29834 2932
rect 29868 1356 29880 2932
rect 29822 1344 29880 1356
rect 30280 2932 30338 2944
rect 30280 1356 30292 2932
rect 30326 1356 30338 2932
rect 30280 1344 30338 1356
rect 30738 2932 30796 2944
rect 30738 1356 30750 2932
rect 30784 1356 30796 2932
rect 30738 1344 30796 1356
rect 31196 2932 31254 2944
rect 31196 1356 31208 2932
rect 31242 1356 31254 2932
rect 31196 1344 31254 1356
rect 31654 2932 31712 2944
rect 31654 1356 31666 2932
rect 31700 1356 31712 2932
rect 31654 1344 31712 1356
rect 32112 2932 32170 2944
rect 32112 1356 32124 2932
rect 32158 1356 32170 2932
rect 32112 1344 32170 1356
rect 32570 2932 32628 2944
rect 32570 1356 32582 2932
rect 32616 1356 32628 2932
rect 32570 1344 32628 1356
rect 23767 267 23825 279
rect 23767 -909 23779 267
rect 23813 -909 23825 267
rect 23767 -921 23825 -909
rect 24225 267 24283 279
rect 24225 -909 24237 267
rect 24271 -909 24283 267
rect 24225 -921 24283 -909
rect 24683 267 24741 279
rect 24683 -909 24695 267
rect 24729 -909 24741 267
rect 24683 -921 24741 -909
rect 25141 267 25199 279
rect 25141 -909 25153 267
rect 25187 -909 25199 267
rect 25141 -921 25199 -909
rect 25599 267 25657 279
rect 25599 -909 25611 267
rect 25645 -909 25657 267
rect 25599 -921 25657 -909
rect 26057 267 26115 279
rect 26057 -909 26069 267
rect 26103 -909 26115 267
rect 26057 -921 26115 -909
rect 26515 267 26573 279
rect 26515 -909 26527 267
rect 26561 -909 26573 267
rect 26515 -921 26573 -909
rect 26973 267 27031 279
rect 26973 -909 26985 267
rect 27019 -909 27031 267
rect 26973 -921 27031 -909
rect 27431 267 27489 279
rect 27431 -909 27443 267
rect 27477 -909 27489 267
rect 27431 -921 27489 -909
rect 27889 267 27947 279
rect 27889 -909 27901 267
rect 27935 -909 27947 267
rect 27889 -921 27947 -909
rect 28347 267 28405 279
rect 28347 -909 28359 267
rect 28393 -909 28405 267
rect 28347 -921 28405 -909
rect 28767 267 28825 279
rect 28767 -909 28779 267
rect 28813 -909 28825 267
rect 28767 -921 28825 -909
rect 29225 267 29283 279
rect 29225 -909 29237 267
rect 29271 -909 29283 267
rect 29225 -921 29283 -909
rect 29683 267 29741 279
rect 29683 -909 29695 267
rect 29729 -909 29741 267
rect 29683 -921 29741 -909
rect 30141 267 30199 279
rect 30141 -909 30153 267
rect 30187 -909 30199 267
rect 30141 -921 30199 -909
rect 30599 267 30657 279
rect 30599 -909 30611 267
rect 30645 -909 30657 267
rect 30599 -921 30657 -909
rect 31057 267 31115 279
rect 31057 -909 31069 267
rect 31103 -909 31115 267
rect 31057 -921 31115 -909
rect 31515 267 31573 279
rect 31515 -909 31527 267
rect 31561 -909 31573 267
rect 31515 -921 31573 -909
rect 31973 267 32031 279
rect 31973 -909 31985 267
rect 32019 -909 32031 267
rect 31973 -921 32031 -909
rect 32431 267 32489 279
rect 32431 -909 32443 267
rect 32477 -909 32489 267
rect 32431 -921 32489 -909
rect 32889 267 32947 279
rect 32889 -909 32901 267
rect 32935 -909 32947 267
rect 32889 -921 32947 -909
rect 33347 267 33405 279
rect 33347 -909 33359 267
rect 33393 -909 33405 267
rect 33347 -921 33405 -909
rect 12697 -7847 12755 -7835
rect 12697 -9023 12709 -7847
rect 12743 -9023 12755 -7847
rect 12697 -9035 12755 -9023
rect 13155 -7847 13213 -7835
rect 13155 -9023 13167 -7847
rect 13201 -9023 13213 -7847
rect 13155 -9035 13213 -9023
rect 13613 -7847 13671 -7835
rect 13613 -9023 13625 -7847
rect 13659 -9023 13671 -7847
rect 13613 -9035 13671 -9023
rect 14071 -7847 14129 -7835
rect 14071 -9023 14083 -7847
rect 14117 -9023 14129 -7847
rect 14071 -9035 14129 -9023
rect 14529 -7847 14587 -7835
rect 14529 -9023 14541 -7847
rect 14575 -9023 14587 -7847
rect 14529 -9035 14587 -9023
rect 14987 -7847 15045 -7835
rect 14987 -9023 14999 -7847
rect 15033 -9023 15045 -7847
rect 14987 -9035 15045 -9023
rect 15445 -7847 15503 -7835
rect 15445 -9023 15457 -7847
rect 15491 -9023 15503 -7847
rect 15445 -9035 15503 -9023
rect 15903 -7847 15961 -7835
rect 15903 -9023 15915 -7847
rect 15949 -9023 15961 -7847
rect 15903 -9035 15961 -9023
rect 16361 -7847 16419 -7835
rect 16361 -9023 16373 -7847
rect 16407 -9023 16419 -7847
rect 16361 -9035 16419 -9023
rect 16819 -7847 16877 -7835
rect 16819 -9023 16831 -7847
rect 16865 -9023 16877 -7847
rect 16819 -9035 16877 -9023
rect 17277 -7847 17335 -7835
rect 17277 -9023 17289 -7847
rect 17323 -9023 17335 -7847
rect 17277 -9035 17335 -9023
rect 17697 -7847 17755 -7835
rect 17697 -9023 17709 -7847
rect 17743 -9023 17755 -7847
rect 17697 -9035 17755 -9023
rect 18155 -7847 18213 -7835
rect 18155 -9023 18167 -7847
rect 18201 -9023 18213 -7847
rect 18155 -9035 18213 -9023
rect 18613 -7847 18671 -7835
rect 18613 -9023 18625 -7847
rect 18659 -9023 18671 -7847
rect 18613 -9035 18671 -9023
rect 19071 -7847 19129 -7835
rect 19071 -9023 19083 -7847
rect 19117 -9023 19129 -7847
rect 19071 -9035 19129 -9023
rect 19529 -7847 19587 -7835
rect 19529 -9023 19541 -7847
rect 19575 -9023 19587 -7847
rect 19529 -9035 19587 -9023
rect 19987 -7847 20045 -7835
rect 19987 -9023 19999 -7847
rect 20033 -9023 20045 -7847
rect 19987 -9035 20045 -9023
rect 20445 -7847 20503 -7835
rect 20445 -9023 20457 -7847
rect 20491 -9023 20503 -7847
rect 20445 -9035 20503 -9023
rect 20903 -7847 20961 -7835
rect 20903 -9023 20915 -7847
rect 20949 -9023 20961 -7847
rect 20903 -9035 20961 -9023
rect 21361 -7847 21419 -7835
rect 21361 -9023 21373 -7847
rect 21407 -9023 21419 -7847
rect 21361 -9035 21419 -9023
rect 21819 -7847 21877 -7835
rect 21819 -9023 21831 -7847
rect 21865 -9023 21877 -7847
rect 21819 -9035 21877 -9023
rect 22277 -7847 22335 -7835
rect 22277 -9023 22289 -7847
rect 22323 -9023 22335 -7847
rect 22277 -9035 22335 -9023
rect 13474 -10112 13532 -10100
rect 13474 -11688 13486 -10112
rect 13520 -11688 13532 -10112
rect 13474 -11700 13532 -11688
rect 13932 -10112 13990 -10100
rect 13932 -11688 13944 -10112
rect 13978 -11688 13990 -10112
rect 13932 -11700 13990 -11688
rect 14390 -10112 14448 -10100
rect 14390 -11688 14402 -10112
rect 14436 -11688 14448 -10112
rect 14390 -11700 14448 -11688
rect 14848 -10112 14906 -10100
rect 14848 -11688 14860 -10112
rect 14894 -11688 14906 -10112
rect 14848 -11700 14906 -11688
rect 15306 -10112 15364 -10100
rect 15306 -11688 15318 -10112
rect 15352 -11688 15364 -10112
rect 15306 -11700 15364 -11688
rect 15764 -10112 15822 -10100
rect 15764 -11688 15776 -10112
rect 15810 -11688 15822 -10112
rect 15764 -11700 15822 -11688
rect 16222 -10112 16280 -10100
rect 16222 -11688 16234 -10112
rect 16268 -11688 16280 -10112
rect 16222 -11700 16280 -11688
rect 16680 -10112 16738 -10100
rect 16680 -11688 16692 -10112
rect 16726 -11688 16738 -10112
rect 16680 -11700 16738 -11688
rect 17138 -10112 17196 -10100
rect 17138 -11688 17150 -10112
rect 17184 -11688 17196 -10112
rect 17138 -11700 17196 -11688
rect 17596 -10112 17654 -10100
rect 17596 -11688 17608 -10112
rect 17642 -11688 17654 -10112
rect 17596 -11700 17654 -11688
rect 18054 -10112 18112 -10100
rect 18054 -11688 18066 -10112
rect 18100 -11688 18112 -10112
rect 18054 -11700 18112 -11688
rect 18512 -10112 18570 -10100
rect 18512 -11688 18524 -10112
rect 18558 -11688 18570 -10112
rect 18512 -11700 18570 -11688
rect 18970 -10112 19028 -10100
rect 18970 -11688 18982 -10112
rect 19016 -11688 19028 -10112
rect 18970 -11700 19028 -11688
rect 19428 -10112 19486 -10100
rect 19428 -11688 19440 -10112
rect 19474 -11688 19486 -10112
rect 19428 -11700 19486 -11688
rect 19886 -10112 19944 -10100
rect 19886 -11688 19898 -10112
rect 19932 -11688 19944 -10112
rect 19886 -11700 19944 -11688
rect 20344 -10112 20402 -10100
rect 20344 -11688 20356 -10112
rect 20390 -11688 20402 -10112
rect 20344 -11700 20402 -11688
rect 20802 -10112 20860 -10100
rect 20802 -11688 20814 -10112
rect 20848 -11688 20860 -10112
rect 20802 -11700 20860 -11688
rect 21260 -10112 21318 -10100
rect 21260 -11688 21272 -10112
rect 21306 -11688 21318 -10112
rect 21260 -11700 21318 -11688
rect 21718 -10112 21776 -10100
rect 21718 -11688 21730 -10112
rect 21764 -11688 21776 -10112
rect 21718 -11700 21776 -11688
rect 27697 -7847 27755 -7835
rect 27697 -9023 27709 -7847
rect 27743 -9023 27755 -7847
rect 27697 -9035 27755 -9023
rect 28155 -7847 28213 -7835
rect 28155 -9023 28167 -7847
rect 28201 -9023 28213 -7847
rect 28155 -9035 28213 -9023
rect 28613 -7847 28671 -7835
rect 28613 -9023 28625 -7847
rect 28659 -9023 28671 -7847
rect 28613 -9035 28671 -9023
rect 29071 -7847 29129 -7835
rect 29071 -9023 29083 -7847
rect 29117 -9023 29129 -7847
rect 29071 -9035 29129 -9023
rect 29529 -7847 29587 -7835
rect 29529 -9023 29541 -7847
rect 29575 -9023 29587 -7847
rect 29529 -9035 29587 -9023
rect 29987 -7847 30045 -7835
rect 29987 -9023 29999 -7847
rect 30033 -9023 30045 -7847
rect 29987 -9035 30045 -9023
rect 30445 -7847 30503 -7835
rect 30445 -9023 30457 -7847
rect 30491 -9023 30503 -7847
rect 30445 -9035 30503 -9023
rect 30903 -7847 30961 -7835
rect 30903 -9023 30915 -7847
rect 30949 -9023 30961 -7847
rect 30903 -9035 30961 -9023
rect 31361 -7847 31419 -7835
rect 31361 -9023 31373 -7847
rect 31407 -9023 31419 -7847
rect 31361 -9035 31419 -9023
rect 31819 -7847 31877 -7835
rect 31819 -9023 31831 -7847
rect 31865 -9023 31877 -7847
rect 31819 -9035 31877 -9023
rect 32277 -7847 32335 -7835
rect 32277 -9023 32289 -7847
rect 32323 -9023 32335 -7847
rect 32277 -9035 32335 -9023
rect 32697 -7847 32755 -7835
rect 32697 -9023 32709 -7847
rect 32743 -9023 32755 -7847
rect 32697 -9035 32755 -9023
rect 33155 -7847 33213 -7835
rect 33155 -9023 33167 -7847
rect 33201 -9023 33213 -7847
rect 33155 -9035 33213 -9023
rect 33613 -7847 33671 -7835
rect 33613 -9023 33625 -7847
rect 33659 -9023 33671 -7847
rect 33613 -9035 33671 -9023
rect 34071 -7847 34129 -7835
rect 34071 -9023 34083 -7847
rect 34117 -9023 34129 -7847
rect 34071 -9035 34129 -9023
rect 34529 -7847 34587 -7835
rect 34529 -9023 34541 -7847
rect 34575 -9023 34587 -7847
rect 34529 -9035 34587 -9023
rect 34987 -7847 35045 -7835
rect 34987 -9023 34999 -7847
rect 35033 -9023 35045 -7847
rect 34987 -9035 35045 -9023
rect 35445 -7847 35503 -7835
rect 35445 -9023 35457 -7847
rect 35491 -9023 35503 -7847
rect 35445 -9035 35503 -9023
rect 35903 -7847 35961 -7835
rect 35903 -9023 35915 -7847
rect 35949 -9023 35961 -7847
rect 35903 -9035 35961 -9023
rect 36361 -7847 36419 -7835
rect 36361 -9023 36373 -7847
rect 36407 -9023 36419 -7847
rect 36361 -9035 36419 -9023
rect 36819 -7847 36877 -7835
rect 36819 -9023 36831 -7847
rect 36865 -9023 36877 -7847
rect 36819 -9035 36877 -9023
rect 37277 -7847 37335 -7835
rect 37277 -9023 37289 -7847
rect 37323 -9023 37335 -7847
rect 37277 -9035 37335 -9023
rect 28474 -10112 28532 -10100
rect 28474 -11688 28486 -10112
rect 28520 -11688 28532 -10112
rect 28474 -11700 28532 -11688
rect 28932 -10112 28990 -10100
rect 28932 -11688 28944 -10112
rect 28978 -11688 28990 -10112
rect 28932 -11700 28990 -11688
rect 29390 -10112 29448 -10100
rect 29390 -11688 29402 -10112
rect 29436 -11688 29448 -10112
rect 29390 -11700 29448 -11688
rect 29848 -10112 29906 -10100
rect 29848 -11688 29860 -10112
rect 29894 -11688 29906 -10112
rect 29848 -11700 29906 -11688
rect 30306 -10112 30364 -10100
rect 30306 -11688 30318 -10112
rect 30352 -11688 30364 -10112
rect 30306 -11700 30364 -11688
rect 30764 -10112 30822 -10100
rect 30764 -11688 30776 -10112
rect 30810 -11688 30822 -10112
rect 30764 -11700 30822 -11688
rect 31222 -10112 31280 -10100
rect 31222 -11688 31234 -10112
rect 31268 -11688 31280 -10112
rect 31222 -11700 31280 -11688
rect 31680 -10112 31738 -10100
rect 31680 -11688 31692 -10112
rect 31726 -11688 31738 -10112
rect 31680 -11700 31738 -11688
rect 32138 -10112 32196 -10100
rect 32138 -11688 32150 -10112
rect 32184 -11688 32196 -10112
rect 32138 -11700 32196 -11688
rect 32596 -10112 32654 -10100
rect 32596 -11688 32608 -10112
rect 32642 -11688 32654 -10112
rect 32596 -11700 32654 -11688
rect 33054 -10112 33112 -10100
rect 33054 -11688 33066 -10112
rect 33100 -11688 33112 -10112
rect 33054 -11700 33112 -11688
rect 33512 -10112 33570 -10100
rect 33512 -11688 33524 -10112
rect 33558 -11688 33570 -10112
rect 33512 -11700 33570 -11688
rect 33970 -10112 34028 -10100
rect 33970 -11688 33982 -10112
rect 34016 -11688 34028 -10112
rect 33970 -11700 34028 -11688
rect 34428 -10112 34486 -10100
rect 34428 -11688 34440 -10112
rect 34474 -11688 34486 -10112
rect 34428 -11700 34486 -11688
rect 34886 -10112 34944 -10100
rect 34886 -11688 34898 -10112
rect 34932 -11688 34944 -10112
rect 34886 -11700 34944 -11688
rect 35344 -10112 35402 -10100
rect 35344 -11688 35356 -10112
rect 35390 -11688 35402 -10112
rect 35344 -11700 35402 -11688
rect 35802 -10112 35860 -10100
rect 35802 -11688 35814 -10112
rect 35848 -11688 35860 -10112
rect 35802 -11700 35860 -11688
rect 36260 -10112 36318 -10100
rect 36260 -11688 36272 -10112
rect 36306 -11688 36318 -10112
rect 36260 -11700 36318 -11688
rect 36718 -10112 36776 -10100
rect 36718 -11688 36730 -10112
rect 36764 -11688 36776 -10112
rect 36718 -11700 36776 -11688
rect 9326 -15068 9384 -15056
rect 9326 -16644 9338 -15068
rect 9372 -16644 9384 -15068
rect 9326 -16656 9384 -16644
rect 9784 -15068 9842 -15056
rect 9784 -16644 9796 -15068
rect 9830 -16644 9842 -15068
rect 9784 -16656 9842 -16644
rect 10242 -15068 10300 -15056
rect 10242 -16644 10254 -15068
rect 10288 -16644 10300 -15068
rect 10242 -16656 10300 -16644
rect 10700 -15068 10758 -15056
rect 10700 -16644 10712 -15068
rect 10746 -16644 10758 -15068
rect 10700 -16656 10758 -16644
rect 11158 -15068 11216 -15056
rect 11158 -16644 11170 -15068
rect 11204 -16644 11216 -15068
rect 11158 -16656 11216 -16644
rect 11616 -15068 11674 -15056
rect 11616 -16644 11628 -15068
rect 11662 -16644 11674 -15068
rect 11616 -16656 11674 -16644
rect 12074 -15068 12132 -15056
rect 12074 -16644 12086 -15068
rect 12120 -16644 12132 -15068
rect 12074 -16656 12132 -16644
rect 12532 -15068 12590 -15056
rect 12532 -16644 12544 -15068
rect 12578 -16644 12590 -15068
rect 12532 -16656 12590 -16644
rect 12990 -15068 13048 -15056
rect 12990 -16644 13002 -15068
rect 13036 -16644 13048 -15068
rect 12990 -16656 13048 -16644
rect 13448 -15068 13506 -15056
rect 13448 -16644 13460 -15068
rect 13494 -16644 13506 -15068
rect 13448 -16656 13506 -16644
rect 13906 -15068 13964 -15056
rect 13906 -16644 13918 -15068
rect 13952 -16644 13964 -15068
rect 13906 -16656 13964 -16644
rect 14364 -15068 14422 -15056
rect 14364 -16644 14376 -15068
rect 14410 -16644 14422 -15068
rect 14364 -16656 14422 -16644
rect 14822 -15068 14880 -15056
rect 14822 -16644 14834 -15068
rect 14868 -16644 14880 -15068
rect 14822 -16656 14880 -16644
rect 15280 -15068 15338 -15056
rect 15280 -16644 15292 -15068
rect 15326 -16644 15338 -15068
rect 15280 -16656 15338 -16644
rect 15738 -15068 15796 -15056
rect 15738 -16644 15750 -15068
rect 15784 -16644 15796 -15068
rect 15738 -16656 15796 -16644
rect 16196 -15068 16254 -15056
rect 16196 -16644 16208 -15068
rect 16242 -16644 16254 -15068
rect 16196 -16656 16254 -16644
rect 16654 -15068 16712 -15056
rect 16654 -16644 16666 -15068
rect 16700 -16644 16712 -15068
rect 16654 -16656 16712 -16644
rect 17112 -15068 17170 -15056
rect 17112 -16644 17124 -15068
rect 17158 -16644 17170 -15068
rect 17112 -16656 17170 -16644
rect 17570 -15068 17628 -15056
rect 17570 -16644 17582 -15068
rect 17616 -16644 17628 -15068
rect 17570 -16656 17628 -16644
rect 8767 -17733 8825 -17721
rect 8767 -18909 8779 -17733
rect 8813 -18909 8825 -17733
rect 8767 -18921 8825 -18909
rect 9225 -17733 9283 -17721
rect 9225 -18909 9237 -17733
rect 9271 -18909 9283 -17733
rect 9225 -18921 9283 -18909
rect 9683 -17733 9741 -17721
rect 9683 -18909 9695 -17733
rect 9729 -18909 9741 -17733
rect 9683 -18921 9741 -18909
rect 10141 -17733 10199 -17721
rect 10141 -18909 10153 -17733
rect 10187 -18909 10199 -17733
rect 10141 -18921 10199 -18909
rect 10599 -17733 10657 -17721
rect 10599 -18909 10611 -17733
rect 10645 -18909 10657 -17733
rect 10599 -18921 10657 -18909
rect 11057 -17733 11115 -17721
rect 11057 -18909 11069 -17733
rect 11103 -18909 11115 -17733
rect 11057 -18921 11115 -18909
rect 11515 -17733 11573 -17721
rect 11515 -18909 11527 -17733
rect 11561 -18909 11573 -17733
rect 11515 -18921 11573 -18909
rect 11973 -17733 12031 -17721
rect 11973 -18909 11985 -17733
rect 12019 -18909 12031 -17733
rect 11973 -18921 12031 -18909
rect 12431 -17733 12489 -17721
rect 12431 -18909 12443 -17733
rect 12477 -18909 12489 -17733
rect 12431 -18921 12489 -18909
rect 12889 -17733 12947 -17721
rect 12889 -18909 12901 -17733
rect 12935 -18909 12947 -17733
rect 12889 -18921 12947 -18909
rect 13347 -17733 13405 -17721
rect 13347 -18909 13359 -17733
rect 13393 -18909 13405 -17733
rect 13347 -18921 13405 -18909
rect 13767 -17733 13825 -17721
rect 13767 -18909 13779 -17733
rect 13813 -18909 13825 -17733
rect 13767 -18921 13825 -18909
rect 14225 -17733 14283 -17721
rect 14225 -18909 14237 -17733
rect 14271 -18909 14283 -17733
rect 14225 -18921 14283 -18909
rect 14683 -17733 14741 -17721
rect 14683 -18909 14695 -17733
rect 14729 -18909 14741 -17733
rect 14683 -18921 14741 -18909
rect 15141 -17733 15199 -17721
rect 15141 -18909 15153 -17733
rect 15187 -18909 15199 -17733
rect 15141 -18921 15199 -18909
rect 15599 -17733 15657 -17721
rect 15599 -18909 15611 -17733
rect 15645 -18909 15657 -17733
rect 15599 -18921 15657 -18909
rect 16057 -17733 16115 -17721
rect 16057 -18909 16069 -17733
rect 16103 -18909 16115 -17733
rect 16057 -18921 16115 -18909
rect 16515 -17733 16573 -17721
rect 16515 -18909 16527 -17733
rect 16561 -18909 16573 -17733
rect 16515 -18921 16573 -18909
rect 16973 -17733 17031 -17721
rect 16973 -18909 16985 -17733
rect 17019 -18909 17031 -17733
rect 16973 -18921 17031 -18909
rect 17431 -17733 17489 -17721
rect 17431 -18909 17443 -17733
rect 17477 -18909 17489 -17733
rect 17431 -18921 17489 -18909
rect 17889 -17733 17947 -17721
rect 17889 -18909 17901 -17733
rect 17935 -18909 17947 -17733
rect 17889 -18921 17947 -18909
rect 18347 -17733 18405 -17721
rect 18347 -18909 18359 -17733
rect 18393 -18909 18405 -17733
rect 18347 -18921 18405 -18909
rect 24326 -15068 24384 -15056
rect 24326 -16644 24338 -15068
rect 24372 -16644 24384 -15068
rect 24326 -16656 24384 -16644
rect 24784 -15068 24842 -15056
rect 24784 -16644 24796 -15068
rect 24830 -16644 24842 -15068
rect 24784 -16656 24842 -16644
rect 25242 -15068 25300 -15056
rect 25242 -16644 25254 -15068
rect 25288 -16644 25300 -15068
rect 25242 -16656 25300 -16644
rect 25700 -15068 25758 -15056
rect 25700 -16644 25712 -15068
rect 25746 -16644 25758 -15068
rect 25700 -16656 25758 -16644
rect 26158 -15068 26216 -15056
rect 26158 -16644 26170 -15068
rect 26204 -16644 26216 -15068
rect 26158 -16656 26216 -16644
rect 26616 -15068 26674 -15056
rect 26616 -16644 26628 -15068
rect 26662 -16644 26674 -15068
rect 26616 -16656 26674 -16644
rect 27074 -15068 27132 -15056
rect 27074 -16644 27086 -15068
rect 27120 -16644 27132 -15068
rect 27074 -16656 27132 -16644
rect 27532 -15068 27590 -15056
rect 27532 -16644 27544 -15068
rect 27578 -16644 27590 -15068
rect 27532 -16656 27590 -16644
rect 27990 -15068 28048 -15056
rect 27990 -16644 28002 -15068
rect 28036 -16644 28048 -15068
rect 27990 -16656 28048 -16644
rect 28448 -15068 28506 -15056
rect 28448 -16644 28460 -15068
rect 28494 -16644 28506 -15068
rect 28448 -16656 28506 -16644
rect 28906 -15068 28964 -15056
rect 28906 -16644 28918 -15068
rect 28952 -16644 28964 -15068
rect 28906 -16656 28964 -16644
rect 29364 -15068 29422 -15056
rect 29364 -16644 29376 -15068
rect 29410 -16644 29422 -15068
rect 29364 -16656 29422 -16644
rect 29822 -15068 29880 -15056
rect 29822 -16644 29834 -15068
rect 29868 -16644 29880 -15068
rect 29822 -16656 29880 -16644
rect 30280 -15068 30338 -15056
rect 30280 -16644 30292 -15068
rect 30326 -16644 30338 -15068
rect 30280 -16656 30338 -16644
rect 30738 -15068 30796 -15056
rect 30738 -16644 30750 -15068
rect 30784 -16644 30796 -15068
rect 30738 -16656 30796 -16644
rect 31196 -15068 31254 -15056
rect 31196 -16644 31208 -15068
rect 31242 -16644 31254 -15068
rect 31196 -16656 31254 -16644
rect 31654 -15068 31712 -15056
rect 31654 -16644 31666 -15068
rect 31700 -16644 31712 -15068
rect 31654 -16656 31712 -16644
rect 32112 -15068 32170 -15056
rect 32112 -16644 32124 -15068
rect 32158 -16644 32170 -15068
rect 32112 -16656 32170 -16644
rect 32570 -15068 32628 -15056
rect 32570 -16644 32582 -15068
rect 32616 -16644 32628 -15068
rect 32570 -16656 32628 -16644
rect 23767 -17733 23825 -17721
rect 23767 -18909 23779 -17733
rect 23813 -18909 23825 -17733
rect 23767 -18921 23825 -18909
rect 24225 -17733 24283 -17721
rect 24225 -18909 24237 -17733
rect 24271 -18909 24283 -17733
rect 24225 -18921 24283 -18909
rect 24683 -17733 24741 -17721
rect 24683 -18909 24695 -17733
rect 24729 -18909 24741 -17733
rect 24683 -18921 24741 -18909
rect 25141 -17733 25199 -17721
rect 25141 -18909 25153 -17733
rect 25187 -18909 25199 -17733
rect 25141 -18921 25199 -18909
rect 25599 -17733 25657 -17721
rect 25599 -18909 25611 -17733
rect 25645 -18909 25657 -17733
rect 25599 -18921 25657 -18909
rect 26057 -17733 26115 -17721
rect 26057 -18909 26069 -17733
rect 26103 -18909 26115 -17733
rect 26057 -18921 26115 -18909
rect 26515 -17733 26573 -17721
rect 26515 -18909 26527 -17733
rect 26561 -18909 26573 -17733
rect 26515 -18921 26573 -18909
rect 26973 -17733 27031 -17721
rect 26973 -18909 26985 -17733
rect 27019 -18909 27031 -17733
rect 26973 -18921 27031 -18909
rect 27431 -17733 27489 -17721
rect 27431 -18909 27443 -17733
rect 27477 -18909 27489 -17733
rect 27431 -18921 27489 -18909
rect 27889 -17733 27947 -17721
rect 27889 -18909 27901 -17733
rect 27935 -18909 27947 -17733
rect 27889 -18921 27947 -18909
rect 28347 -17733 28405 -17721
rect 28347 -18909 28359 -17733
rect 28393 -18909 28405 -17733
rect 28347 -18921 28405 -18909
rect 28767 -17733 28825 -17721
rect 28767 -18909 28779 -17733
rect 28813 -18909 28825 -17733
rect 28767 -18921 28825 -18909
rect 29225 -17733 29283 -17721
rect 29225 -18909 29237 -17733
rect 29271 -18909 29283 -17733
rect 29225 -18921 29283 -18909
rect 29683 -17733 29741 -17721
rect 29683 -18909 29695 -17733
rect 29729 -18909 29741 -17733
rect 29683 -18921 29741 -18909
rect 30141 -17733 30199 -17721
rect 30141 -18909 30153 -17733
rect 30187 -18909 30199 -17733
rect 30141 -18921 30199 -18909
rect 30599 -17733 30657 -17721
rect 30599 -18909 30611 -17733
rect 30645 -18909 30657 -17733
rect 30599 -18921 30657 -18909
rect 31057 -17733 31115 -17721
rect 31057 -18909 31069 -17733
rect 31103 -18909 31115 -17733
rect 31057 -18921 31115 -18909
rect 31515 -17733 31573 -17721
rect 31515 -18909 31527 -17733
rect 31561 -18909 31573 -17733
rect 31515 -18921 31573 -18909
rect 31973 -17733 32031 -17721
rect 31973 -18909 31985 -17733
rect 32019 -18909 32031 -17733
rect 31973 -18921 32031 -18909
rect 32431 -17733 32489 -17721
rect 32431 -18909 32443 -17733
rect 32477 -18909 32489 -17733
rect 32431 -18921 32489 -18909
rect 32889 -17733 32947 -17721
rect 32889 -18909 32901 -17733
rect 32935 -18909 32947 -17733
rect 32889 -18921 32947 -18909
rect 33347 -17733 33405 -17721
rect 33347 -18909 33359 -17733
rect 33393 -18909 33405 -17733
rect 33347 -18921 33405 -18909
<< ndiffc >>
rect 24163 13719 24197 13895
rect 24421 13719 24455 13895
rect 24679 13719 24713 13895
rect 24937 13719 24971 13895
rect 25285 13719 25319 13895
rect 25543 13719 25577 13895
rect 25801 13719 25835 13895
rect 26059 13719 26093 13895
rect 26317 13719 26351 13895
rect 26575 13719 26609 13895
rect 26833 13719 26867 13895
rect 27295 13999 27329 14033
rect 27379 13973 27413 14007
rect 27463 13999 27497 14033
rect 27585 13969 27619 14003
rect 27718 13975 27752 14009
rect 27825 13975 27859 14009
rect 28171 13973 28205 14007
rect 28283 13969 28317 14003
rect 28393 13973 28427 14007
rect 28605 13969 28639 14003
rect 28823 13989 28857 14023
rect 28927 14012 28961 14046
rect 29011 14045 29045 14079
rect 29011 13977 29045 14011
rect 29115 13999 29149 14033
rect 29212 13993 29246 14027
rect 29296 14023 29330 14057
rect 29452 14045 29486 14079
rect 29452 13977 29486 14011
rect 29536 14045 29570 14079
rect 29536 13977 29570 14011
rect 29691 14041 29725 14075
rect 29691 13973 29725 14007
rect 29859 14041 29893 14075
rect 29859 13973 29893 14007
rect 30010 14045 30044 14079
rect 30010 13977 30044 14011
rect 30094 14045 30128 14079
rect 30094 13977 30128 14011
rect 30250 14023 30284 14057
rect 30535 14045 30569 14079
rect 30334 13993 30368 14027
rect 30431 13999 30465 14033
rect 30535 13977 30569 14011
rect 30619 14012 30653 14046
rect 30723 13989 30757 14023
rect 30941 13969 30975 14003
rect 31153 13973 31187 14007
rect 31263 13969 31297 14003
rect 31375 13973 31409 14007
rect 31721 13975 31755 14009
rect 31828 13975 31862 14009
rect 31961 13969 31995 14003
rect 32083 13999 32117 14033
rect 32167 13973 32201 14007
rect 32251 13999 32285 14033
rect 24250 12666 24284 12842
rect 25108 12666 25142 12842
rect 25966 12666 26000 12842
rect 26824 12666 26858 12842
rect 27682 12666 27716 12842
rect 28540 12666 28574 12842
rect 29398 12666 29432 12842
rect 30256 12666 30290 12842
rect 31114 12666 31148 12842
rect 31972 12666 32006 12842
rect 24250 12084 24284 12260
rect 25108 12084 25142 12260
rect 25966 12084 26000 12260
rect 26824 12084 26858 12260
rect 27682 12084 27716 12260
rect 28540 12084 28574 12260
rect 29398 12084 29432 12260
rect 30256 12084 30290 12260
rect 31114 12084 31148 12260
rect 31972 12084 32006 12260
rect 15168 9480 15202 9656
rect 15626 9480 15660 9656
rect 16084 9480 16118 9656
rect 16542 9480 16576 9656
rect 17000 9480 17034 9656
rect 17458 9480 17492 9656
rect 17916 9480 17950 9656
rect 18374 9480 18408 9656
rect 18832 9480 18866 9656
rect 19290 9480 19324 9656
rect 19748 9480 19782 9656
rect 23930 9480 23964 9656
rect 24388 9480 24422 9656
rect 24846 9480 24880 9656
rect 25304 9480 25338 9656
rect 25762 9480 25796 9656
rect 26220 9480 26254 9656
rect 26678 9480 26712 9656
rect 27136 9480 27170 9656
rect 27594 9480 27628 9656
rect 28052 9480 28086 9656
rect 28510 9480 28544 9656
rect 29152 8817 29186 8851
rect 29152 8749 29186 8783
rect 29236 8817 29270 8851
rect 29236 8749 29270 8783
rect 29397 8821 29431 8855
rect 29481 8813 29515 8847
rect 29565 8821 29599 8855
rect 29649 8813 29683 8847
rect 29733 8820 29767 8854
rect 30587 8501 30621 8535
rect 30671 8475 30705 8509
rect 30755 8501 30789 8535
rect 30859 8475 30893 8509
rect 30944 8489 30978 8523
rect 31055 8489 31089 8523
rect 31254 8483 31288 8517
rect 31373 8489 31407 8523
rect 31476 8489 31510 8523
rect 31674 8489 31708 8523
rect 31780 8544 31814 8578
rect 31780 8476 31814 8510
rect 31864 8505 31898 8539
rect 31948 8546 31982 8580
rect 31948 8478 31982 8512
rect 32052 8501 32086 8535
rect 32147 8475 32181 8509
rect 32231 8513 32265 8547
rect 32376 8547 32410 8581
rect 32376 8479 32410 8513
rect 32460 8547 32494 8581
rect 32460 8479 32494 8513
rect 32621 8475 32655 8509
rect 32705 8483 32739 8517
rect 32789 8475 32823 8509
rect 32873 8483 32907 8517
rect 32957 8476 32991 8510
rect 30587 8297 30621 8331
rect 30671 8323 30705 8357
rect 30755 8297 30789 8331
rect 30859 8323 30893 8357
rect 30944 8309 30978 8343
rect 31055 8309 31089 8343
rect 31254 8315 31288 8349
rect 31373 8309 31407 8343
rect 31476 8309 31510 8343
rect 31674 8309 31708 8343
rect 31780 8322 31814 8356
rect 31780 8254 31814 8288
rect 31864 8293 31898 8327
rect 31948 8320 31982 8354
rect 31948 8252 31982 8286
rect 32052 8297 32086 8331
rect 32147 8323 32181 8357
rect 32231 8285 32265 8319
rect 32376 8319 32410 8353
rect 32376 8251 32410 8285
rect 32460 8319 32494 8353
rect 32460 8251 32494 8285
rect 32621 8323 32655 8357
rect 32705 8315 32739 8349
rect 32789 8323 32823 8357
rect 32873 8315 32907 8349
rect 32957 8322 32991 8356
rect 33285 8297 33319 8331
rect 33369 8323 33403 8357
rect 33453 8297 33487 8331
rect 33557 8323 33591 8357
rect 33642 8309 33676 8343
rect 33753 8309 33787 8343
rect 33952 8315 33986 8349
rect 34071 8309 34105 8343
rect 34174 8309 34208 8343
rect 34372 8309 34406 8343
rect 34478 8322 34512 8356
rect 34478 8254 34512 8288
rect 34562 8293 34596 8327
rect 34646 8320 34680 8354
rect 34646 8252 34680 8286
rect 34750 8297 34784 8331
rect 34845 8323 34879 8357
rect 34929 8285 34963 8319
rect 35074 8319 35108 8353
rect 35074 8251 35108 8285
rect 35158 8319 35192 8353
rect 35158 8251 35192 8285
rect 35319 8323 35353 8357
rect 35403 8315 35437 8349
rect 35487 8323 35521 8357
rect 35571 8315 35605 8349
rect 35655 8322 35689 8356
rect 30587 7413 30621 7447
rect 30671 7387 30705 7421
rect 30755 7413 30789 7447
rect 30859 7387 30893 7421
rect 30944 7401 30978 7435
rect 31055 7401 31089 7435
rect 31254 7395 31288 7429
rect 31373 7401 31407 7435
rect 31476 7401 31510 7435
rect 31674 7401 31708 7435
rect 31780 7456 31814 7490
rect 31780 7388 31814 7422
rect 31864 7417 31898 7451
rect 31948 7458 31982 7492
rect 31948 7390 31982 7424
rect 32052 7413 32086 7447
rect 32147 7387 32181 7421
rect 32231 7425 32265 7459
rect 32376 7459 32410 7493
rect 32376 7391 32410 7425
rect 32460 7459 32494 7493
rect 32460 7391 32494 7425
rect 32621 7387 32655 7421
rect 32705 7395 32739 7429
rect 32789 7387 32823 7421
rect 32873 7395 32907 7429
rect 32957 7388 32991 7422
rect 33285 7413 33319 7447
rect 33369 7387 33403 7421
rect 33453 7413 33487 7447
rect 33557 7387 33591 7421
rect 33642 7401 33676 7435
rect 33753 7401 33787 7435
rect 33952 7395 33986 7429
rect 34071 7401 34105 7435
rect 34174 7401 34208 7435
rect 34372 7401 34406 7435
rect 34478 7456 34512 7490
rect 34478 7388 34512 7422
rect 34562 7417 34596 7451
rect 34646 7458 34680 7492
rect 34646 7390 34680 7424
rect 34750 7413 34784 7447
rect 34845 7387 34879 7421
rect 34929 7425 34963 7459
rect 35074 7459 35108 7493
rect 35074 7391 35108 7425
rect 35158 7459 35192 7493
rect 35158 7391 35192 7425
rect 35319 7387 35353 7421
rect 35403 7395 35437 7429
rect 35487 7387 35521 7421
rect 35571 7395 35605 7429
rect 35655 7388 35689 7422
rect 30587 7209 30621 7243
rect 30671 7235 30705 7269
rect 30755 7209 30789 7243
rect 30859 7235 30893 7269
rect 30944 7221 30978 7255
rect 31055 7221 31089 7255
rect 31254 7227 31288 7261
rect 31373 7221 31407 7255
rect 31476 7221 31510 7255
rect 31674 7221 31708 7255
rect 31780 7234 31814 7268
rect 31780 7166 31814 7200
rect 31864 7205 31898 7239
rect 31948 7232 31982 7266
rect 31948 7164 31982 7198
rect 32052 7209 32086 7243
rect 32147 7235 32181 7269
rect 32231 7197 32265 7231
rect 32376 7231 32410 7265
rect 32376 7163 32410 7197
rect 32460 7231 32494 7265
rect 32460 7163 32494 7197
rect 32621 7235 32655 7269
rect 32705 7227 32739 7261
rect 32789 7235 32823 7269
rect 32873 7227 32907 7261
rect 32957 7234 32991 7268
rect 33285 7209 33319 7243
rect 33369 7235 33403 7269
rect 33453 7209 33487 7243
rect 33557 7235 33591 7269
rect 33642 7221 33676 7255
rect 33753 7221 33787 7255
rect 33952 7227 33986 7261
rect 34071 7221 34105 7255
rect 34174 7221 34208 7255
rect 34372 7221 34406 7255
rect 34478 7234 34512 7268
rect 34478 7166 34512 7200
rect 34562 7205 34596 7239
rect 34646 7232 34680 7266
rect 34646 7164 34680 7198
rect 34750 7209 34784 7243
rect 34845 7235 34879 7269
rect 34929 7197 34963 7231
rect 35074 7231 35108 7265
rect 35074 7163 35108 7197
rect 35158 7231 35192 7265
rect 35158 7163 35192 7197
rect 35319 7235 35353 7269
rect 35403 7227 35437 7261
rect 35487 7235 35521 7269
rect 35571 7227 35605 7261
rect 35655 7234 35689 7268
rect 30587 6325 30621 6359
rect 30671 6299 30705 6333
rect 30755 6325 30789 6359
rect 30859 6299 30893 6333
rect 30944 6313 30978 6347
rect 31055 6313 31089 6347
rect 31254 6307 31288 6341
rect 31373 6313 31407 6347
rect 31476 6313 31510 6347
rect 31674 6313 31708 6347
rect 31780 6368 31814 6402
rect 31780 6300 31814 6334
rect 31864 6329 31898 6363
rect 31948 6370 31982 6404
rect 31948 6302 31982 6336
rect 32052 6325 32086 6359
rect 32147 6299 32181 6333
rect 32231 6337 32265 6371
rect 32376 6371 32410 6405
rect 32376 6303 32410 6337
rect 32460 6371 32494 6405
rect 32460 6303 32494 6337
rect 32621 6299 32655 6333
rect 32705 6307 32739 6341
rect 32789 6299 32823 6333
rect 32873 6307 32907 6341
rect 32957 6300 32991 6334
rect 33285 6325 33319 6359
rect 33369 6299 33403 6333
rect 33453 6325 33487 6359
rect 33557 6299 33591 6333
rect 33642 6313 33676 6347
rect 33753 6313 33787 6347
rect 33952 6307 33986 6341
rect 34071 6313 34105 6347
rect 34174 6313 34208 6347
rect 34372 6313 34406 6347
rect 34478 6368 34512 6402
rect 34478 6300 34512 6334
rect 34562 6329 34596 6363
rect 34646 6370 34680 6404
rect 34646 6302 34680 6336
rect 34750 6325 34784 6359
rect 34845 6299 34879 6333
rect 34929 6337 34963 6371
rect 35074 6371 35108 6405
rect 35074 6303 35108 6337
rect 35158 6371 35192 6405
rect 35158 6303 35192 6337
rect 35319 6299 35353 6333
rect 35403 6307 35437 6341
rect 35487 6299 35521 6333
rect 35571 6307 35605 6341
rect 35655 6300 35689 6334
rect 30587 6121 30621 6155
rect 30671 6147 30705 6181
rect 30755 6121 30789 6155
rect 30859 6147 30893 6181
rect 30944 6133 30978 6167
rect 31055 6133 31089 6167
rect 31254 6139 31288 6173
rect 31373 6133 31407 6167
rect 31476 6133 31510 6167
rect 31674 6133 31708 6167
rect 31780 6146 31814 6180
rect 31780 6078 31814 6112
rect 31864 6117 31898 6151
rect 31948 6144 31982 6178
rect 31948 6076 31982 6110
rect 32052 6121 32086 6155
rect 32147 6147 32181 6181
rect 32231 6109 32265 6143
rect 32376 6143 32410 6177
rect 32376 6075 32410 6109
rect 32460 6143 32494 6177
rect 32460 6075 32494 6109
rect 32621 6147 32655 6181
rect 32705 6139 32739 6173
rect 32789 6147 32823 6181
rect 32873 6139 32907 6173
rect 32957 6146 32991 6180
rect 33285 6121 33319 6155
rect 33369 6147 33403 6181
rect 33453 6121 33487 6155
rect 33557 6147 33591 6181
rect 33642 6133 33676 6167
rect 33753 6133 33787 6167
rect 33952 6139 33986 6173
rect 34071 6133 34105 6167
rect 34174 6133 34208 6167
rect 34372 6133 34406 6167
rect 34478 6146 34512 6180
rect 34478 6078 34512 6112
rect 34562 6117 34596 6151
rect 34646 6144 34680 6178
rect 34646 6076 34680 6110
rect 34750 6121 34784 6155
rect 34845 6147 34879 6181
rect 34929 6109 34963 6143
rect 35074 6143 35108 6177
rect 35074 6075 35108 6109
rect 35158 6143 35192 6177
rect 35158 6075 35192 6109
rect 35319 6147 35353 6181
rect 35403 6139 35437 6173
rect 35487 6147 35521 6181
rect 35571 6139 35605 6173
rect 35655 6146 35689 6180
rect 8778 -2402 8812 -2226
rect 9236 -2402 9270 -2226
rect 9694 -2402 9728 -2226
rect 10152 -2402 10186 -2226
rect 10610 -2402 10644 -2226
rect 11068 -2402 11102 -2226
rect 11526 -2402 11560 -2226
rect 11984 -2402 12018 -2226
rect 12442 -2402 12476 -2226
rect 12900 -2402 12934 -2226
rect 13358 -2402 13392 -2226
rect 13778 -2402 13812 -2226
rect 14236 -2402 14270 -2226
rect 14694 -2402 14728 -2226
rect 15152 -2402 15186 -2226
rect 15610 -2402 15644 -2226
rect 16068 -2402 16102 -2226
rect 16526 -2402 16560 -2226
rect 16984 -2402 17018 -2226
rect 17442 -2402 17476 -2226
rect 17900 -2402 17934 -2226
rect 18358 -2402 18392 -2226
rect 8778 -3070 8812 -2894
rect 9236 -3070 9270 -2894
rect 9694 -3070 9728 -2894
rect 10152 -3070 10186 -2894
rect 10610 -3070 10644 -2894
rect 11068 -3070 11102 -2894
rect 11526 -3070 11560 -2894
rect 11984 -3070 12018 -2894
rect 12442 -3070 12476 -2894
rect 12900 -3070 12934 -2894
rect 13358 -3070 13392 -2894
rect 23778 -2402 23812 -2226
rect 24236 -2402 24270 -2226
rect 24694 -2402 24728 -2226
rect 25152 -2402 25186 -2226
rect 25610 -2402 25644 -2226
rect 26068 -2402 26102 -2226
rect 26526 -2402 26560 -2226
rect 26984 -2402 27018 -2226
rect 27442 -2402 27476 -2226
rect 27900 -2402 27934 -2226
rect 28358 -2402 28392 -2226
rect 28778 -2402 28812 -2226
rect 29236 -2402 29270 -2226
rect 29694 -2402 29728 -2226
rect 30152 -2402 30186 -2226
rect 30610 -2402 30644 -2226
rect 31068 -2402 31102 -2226
rect 31526 -2402 31560 -2226
rect 31984 -2402 32018 -2226
rect 32442 -2402 32476 -2226
rect 32900 -2402 32934 -2226
rect 33358 -2402 33392 -2226
rect 23778 -3070 23812 -2894
rect 24236 -3070 24270 -2894
rect 24694 -3070 24728 -2894
rect 25152 -3070 25186 -2894
rect 25610 -3070 25644 -2894
rect 26068 -3070 26102 -2894
rect 26526 -3070 26560 -2894
rect 26984 -3070 27018 -2894
rect 27442 -3070 27476 -2894
rect 27900 -3070 27934 -2894
rect 28358 -3070 28392 -2894
rect 17710 -5862 17744 -5686
rect 18168 -5862 18202 -5686
rect 18626 -5862 18660 -5686
rect 19084 -5862 19118 -5686
rect 19542 -5862 19576 -5686
rect 20000 -5862 20034 -5686
rect 20458 -5862 20492 -5686
rect 20916 -5862 20950 -5686
rect 21374 -5862 21408 -5686
rect 21832 -5862 21866 -5686
rect 22290 -5862 22324 -5686
rect 12710 -6530 12744 -6354
rect 13168 -6530 13202 -6354
rect 13626 -6530 13660 -6354
rect 14084 -6530 14118 -6354
rect 14542 -6530 14576 -6354
rect 15000 -6530 15034 -6354
rect 15458 -6530 15492 -6354
rect 15916 -6530 15950 -6354
rect 16374 -6530 16408 -6354
rect 16832 -6530 16866 -6354
rect 17290 -6530 17324 -6354
rect 17710 -6530 17744 -6354
rect 18168 -6530 18202 -6354
rect 18626 -6530 18660 -6354
rect 19084 -6530 19118 -6354
rect 19542 -6530 19576 -6354
rect 20000 -6530 20034 -6354
rect 20458 -6530 20492 -6354
rect 20916 -6530 20950 -6354
rect 21374 -6530 21408 -6354
rect 21832 -6530 21866 -6354
rect 22290 -6530 22324 -6354
rect 32710 -5862 32744 -5686
rect 33168 -5862 33202 -5686
rect 33626 -5862 33660 -5686
rect 34084 -5862 34118 -5686
rect 34542 -5862 34576 -5686
rect 35000 -5862 35034 -5686
rect 35458 -5862 35492 -5686
rect 35916 -5862 35950 -5686
rect 36374 -5862 36408 -5686
rect 36832 -5862 36866 -5686
rect 37290 -5862 37324 -5686
rect 27710 -6530 27744 -6354
rect 28168 -6530 28202 -6354
rect 28626 -6530 28660 -6354
rect 29084 -6530 29118 -6354
rect 29542 -6530 29576 -6354
rect 30000 -6530 30034 -6354
rect 30458 -6530 30492 -6354
rect 30916 -6530 30950 -6354
rect 31374 -6530 31408 -6354
rect 31832 -6530 31866 -6354
rect 32290 -6530 32324 -6354
rect 32710 -6530 32744 -6354
rect 33168 -6530 33202 -6354
rect 33626 -6530 33660 -6354
rect 34084 -6530 34118 -6354
rect 34542 -6530 34576 -6354
rect 35000 -6530 35034 -6354
rect 35458 -6530 35492 -6354
rect 35916 -6530 35950 -6354
rect 36374 -6530 36408 -6354
rect 36832 -6530 36866 -6354
rect 37290 -6530 37324 -6354
rect 8778 -20402 8812 -20226
rect 9236 -20402 9270 -20226
rect 9694 -20402 9728 -20226
rect 10152 -20402 10186 -20226
rect 10610 -20402 10644 -20226
rect 11068 -20402 11102 -20226
rect 11526 -20402 11560 -20226
rect 11984 -20402 12018 -20226
rect 12442 -20402 12476 -20226
rect 12900 -20402 12934 -20226
rect 13358 -20402 13392 -20226
rect 13778 -20402 13812 -20226
rect 14236 -20402 14270 -20226
rect 14694 -20402 14728 -20226
rect 15152 -20402 15186 -20226
rect 15610 -20402 15644 -20226
rect 16068 -20402 16102 -20226
rect 16526 -20402 16560 -20226
rect 16984 -20402 17018 -20226
rect 17442 -20402 17476 -20226
rect 17900 -20402 17934 -20226
rect 18358 -20402 18392 -20226
rect 8778 -21070 8812 -20894
rect 9236 -21070 9270 -20894
rect 9694 -21070 9728 -20894
rect 10152 -21070 10186 -20894
rect 10610 -21070 10644 -20894
rect 11068 -21070 11102 -20894
rect 11526 -21070 11560 -20894
rect 11984 -21070 12018 -20894
rect 12442 -21070 12476 -20894
rect 12900 -21070 12934 -20894
rect 13358 -21070 13392 -20894
rect 23778 -20402 23812 -20226
rect 24236 -20402 24270 -20226
rect 24694 -20402 24728 -20226
rect 25152 -20402 25186 -20226
rect 25610 -20402 25644 -20226
rect 26068 -20402 26102 -20226
rect 26526 -20402 26560 -20226
rect 26984 -20402 27018 -20226
rect 27442 -20402 27476 -20226
rect 27900 -20402 27934 -20226
rect 28358 -20402 28392 -20226
rect 28778 -20402 28812 -20226
rect 29236 -20402 29270 -20226
rect 29694 -20402 29728 -20226
rect 30152 -20402 30186 -20226
rect 30610 -20402 30644 -20226
rect 31068 -20402 31102 -20226
rect 31526 -20402 31560 -20226
rect 31984 -20402 32018 -20226
rect 32442 -20402 32476 -20226
rect 32900 -20402 32934 -20226
rect 33358 -20402 33392 -20226
rect 23778 -21070 23812 -20894
rect 24236 -21070 24270 -20894
rect 24694 -21070 24728 -20894
rect 25152 -21070 25186 -20894
rect 25610 -21070 25644 -20894
rect 26068 -21070 26102 -20894
rect 26526 -21070 26560 -20894
rect 26984 -21070 27018 -20894
rect 27442 -21070 27476 -20894
rect 27900 -21070 27934 -20894
rect 28358 -21070 28392 -20894
<< pdiffc >>
rect 23776 16246 23810 16422
rect 24634 16246 24668 16422
rect 25492 16246 25526 16422
rect 26350 16246 26384 16422
rect 27208 16246 27242 16422
rect 28066 16246 28100 16422
rect 28924 16246 28958 16422
rect 29782 16246 29816 16422
rect 30640 16246 30674 16422
rect 31498 16246 31532 16422
rect 32356 16246 32390 16422
rect 23776 15646 23810 15822
rect 24634 15646 24668 15822
rect 25492 15646 25526 15822
rect 26350 15646 26384 15822
rect 27208 15646 27242 15822
rect 28066 15646 28100 15822
rect 28924 15646 28958 15822
rect 29782 15646 29816 15822
rect 30640 15646 30674 15822
rect 31498 15646 31532 15822
rect 32356 15646 32390 15822
rect 24163 14406 24197 14782
rect 24421 14406 24455 14782
rect 24679 14406 24713 14782
rect 24937 14406 24971 14782
rect 25285 14406 25319 14782
rect 25543 14406 25577 14782
rect 25801 14406 25835 14782
rect 26059 14406 26093 14782
rect 26317 14406 26351 14782
rect 26575 14406 26609 14782
rect 26833 14406 26867 14782
rect 27295 14357 27329 14391
rect 27295 14289 27329 14323
rect 27379 14341 27413 14375
rect 27463 14357 27497 14391
rect 27646 14365 27680 14399
rect 27730 14357 27764 14391
rect 27823 14363 27857 14397
rect 27977 14339 28011 14373
rect 28074 14355 28108 14389
rect 28158 14339 28192 14373
rect 28271 14365 28305 14399
rect 27463 14289 27497 14323
rect 28359 14357 28393 14391
rect 28456 14364 28490 14398
rect 28648 14365 28682 14399
rect 28732 14339 28766 14373
rect 28818 14365 28852 14399
rect 28896 14365 28930 14399
rect 28980 14357 29014 14391
rect 28980 14289 29014 14323
rect 29115 14365 29149 14399
rect 29115 14297 29149 14331
rect 29212 14365 29246 14399
rect 29212 14297 29246 14331
rect 28980 14221 29014 14255
rect 29212 14229 29246 14263
rect 29296 14329 29330 14363
rect 29296 14261 29330 14295
rect 29452 14365 29486 14399
rect 29452 14297 29486 14331
rect 29452 14229 29486 14263
rect 29536 14365 29570 14399
rect 29536 14297 29570 14331
rect 29536 14229 29570 14263
rect 29691 14365 29725 14399
rect 29691 14297 29725 14331
rect 29691 14229 29725 14263
rect 29775 14365 29809 14399
rect 29775 14297 29809 14331
rect 29775 14229 29809 14263
rect 29859 14365 29893 14399
rect 29859 14297 29893 14331
rect 29859 14229 29893 14263
rect 30010 14365 30044 14399
rect 30010 14297 30044 14331
rect 30010 14229 30044 14263
rect 30094 14365 30128 14399
rect 30094 14297 30128 14331
rect 30094 14229 30128 14263
rect 30250 14329 30284 14363
rect 30250 14261 30284 14295
rect 30334 14365 30368 14399
rect 30334 14297 30368 14331
rect 30431 14365 30465 14399
rect 30431 14297 30465 14331
rect 30566 14357 30600 14391
rect 30566 14289 30600 14323
rect 30334 14229 30368 14263
rect 30566 14221 30600 14255
rect 30650 14365 30684 14399
rect 30728 14365 30762 14399
rect 30814 14339 30848 14373
rect 30898 14365 30932 14399
rect 31090 14364 31124 14398
rect 31187 14357 31221 14391
rect 31275 14365 31309 14399
rect 31388 14339 31422 14373
rect 31472 14355 31506 14389
rect 31569 14339 31603 14373
rect 31723 14363 31757 14397
rect 31816 14357 31850 14391
rect 31900 14365 31934 14399
rect 32083 14357 32117 14391
rect 32083 14289 32117 14323
rect 32167 14341 32201 14375
rect 32251 14357 32285 14391
rect 32251 14289 32285 14323
rect 30587 8859 30621 8893
rect 30587 8791 30621 8825
rect 30671 8843 30705 8877
rect 30755 8859 30789 8893
rect 30859 8867 30893 8901
rect 30943 8859 30977 8893
rect 31035 8854 31069 8888
rect 31274 8867 31308 8901
rect 30755 8791 30789 8825
rect 13336 6229 13370 7805
rect 13794 6229 13828 7805
rect 14252 6229 14286 7805
rect 14710 6229 14744 7805
rect 15168 6229 15202 7805
rect 15626 6229 15660 7805
rect 16084 6229 16118 7805
rect 16542 6229 16576 7805
rect 17000 6229 17034 7805
rect 17458 6229 17492 7805
rect 17916 6229 17950 7805
rect 18374 6229 18408 7805
rect 18832 6229 18866 7805
rect 19290 6229 19324 7805
rect 19748 6229 19782 7805
rect 20206 6229 20240 7805
rect 20664 6229 20698 7805
rect 21122 6229 21156 7805
rect 21580 6229 21614 7805
rect 23931 7049 23965 8225
rect 24389 7049 24423 8225
rect 24847 7049 24881 8225
rect 25305 7049 25339 8225
rect 25763 7049 25797 8225
rect 26221 7049 26255 8225
rect 26679 7049 26713 8225
rect 27137 7049 27171 8225
rect 27595 7049 27629 8225
rect 28053 7049 28087 8225
rect 28511 7049 28545 8225
rect 29152 8565 29186 8599
rect 29152 8497 29186 8531
rect 29152 8429 29186 8463
rect 29236 8565 29270 8599
rect 29236 8497 29270 8531
rect 29236 8429 29270 8463
rect 29397 8565 29431 8599
rect 29397 8497 29431 8531
rect 29397 8429 29431 8463
rect 29481 8565 29515 8599
rect 29481 8497 29515 8531
rect 29481 8429 29515 8463
rect 29565 8497 29599 8531
rect 29565 8429 29599 8463
rect 29649 8565 29683 8599
rect 29649 8497 29683 8531
rect 29649 8429 29683 8463
rect 31274 8799 31308 8833
rect 31358 8859 31392 8893
rect 31453 8849 31487 8883
rect 31652 8859 31686 8893
rect 31776 8867 31810 8901
rect 31776 8796 31810 8830
rect 31776 8725 31810 8759
rect 31862 8837 31896 8871
rect 31862 8757 31896 8791
rect 31946 8861 31980 8895
rect 31946 8793 31980 8827
rect 32050 8867 32084 8901
rect 32050 8799 32084 8833
rect 32147 8867 32181 8901
rect 32147 8799 32181 8833
rect 31946 8725 31980 8759
rect 32147 8731 32181 8765
rect 32231 8867 32265 8901
rect 32231 8796 32265 8830
rect 32231 8725 32265 8759
rect 32376 8867 32410 8901
rect 32376 8799 32410 8833
rect 32376 8731 32410 8765
rect 32460 8867 32494 8901
rect 32460 8799 32494 8833
rect 32460 8731 32494 8765
rect 32621 8867 32655 8901
rect 32621 8799 32655 8833
rect 32621 8731 32655 8765
rect 32705 8867 32739 8901
rect 32705 8799 32739 8833
rect 32705 8731 32739 8765
rect 32789 8867 32823 8901
rect 32789 8799 32823 8833
rect 32873 8867 32907 8901
rect 32873 8799 32907 8833
rect 32873 8731 32907 8765
rect 32957 8867 32991 8901
rect 29733 8429 29767 8463
rect 30587 8007 30621 8041
rect 30587 7939 30621 7973
rect 30671 7955 30705 7989
rect 30755 8007 30789 8041
rect 30755 7939 30789 7973
rect 30859 7931 30893 7965
rect 30943 7939 30977 7973
rect 31035 7944 31069 7978
rect 31274 7999 31308 8033
rect 31274 7931 31308 7965
rect 31776 8073 31810 8107
rect 31358 7939 31392 7973
rect 31453 7949 31487 7983
rect 31652 7939 31686 7973
rect 31776 8002 31810 8036
rect 31776 7931 31810 7965
rect 31862 8041 31896 8075
rect 31862 7961 31896 7995
rect 31946 8073 31980 8107
rect 32147 8067 32181 8101
rect 31946 8005 31980 8039
rect 31946 7937 31980 7971
rect 32050 7999 32084 8033
rect 32050 7931 32084 7965
rect 32147 7999 32181 8033
rect 32147 7931 32181 7965
rect 32231 8073 32265 8107
rect 32231 8002 32265 8036
rect 32231 7931 32265 7965
rect 32376 8067 32410 8101
rect 32376 7999 32410 8033
rect 32376 7931 32410 7965
rect 32460 8067 32494 8101
rect 32460 7999 32494 8033
rect 32460 7931 32494 7965
rect 32621 8067 32655 8101
rect 32621 7999 32655 8033
rect 32621 7931 32655 7965
rect 32705 8067 32739 8101
rect 32705 7999 32739 8033
rect 32705 7931 32739 7965
rect 32789 7999 32823 8033
rect 32789 7931 32823 7965
rect 32873 8067 32907 8101
rect 32873 7999 32907 8033
rect 32873 7931 32907 7965
rect 32957 7931 32991 7965
rect 33285 8007 33319 8041
rect 33285 7939 33319 7973
rect 33369 7955 33403 7989
rect 33453 8007 33487 8041
rect 33453 7939 33487 7973
rect 33557 7931 33591 7965
rect 33641 7939 33675 7973
rect 33733 7944 33767 7978
rect 33972 7999 34006 8033
rect 33972 7931 34006 7965
rect 34474 8073 34508 8107
rect 34056 7939 34090 7973
rect 34151 7949 34185 7983
rect 34350 7939 34384 7973
rect 34474 8002 34508 8036
rect 34474 7931 34508 7965
rect 34560 8041 34594 8075
rect 34560 7961 34594 7995
rect 34644 8073 34678 8107
rect 34845 8067 34879 8101
rect 34644 8005 34678 8039
rect 34644 7937 34678 7971
rect 34748 7999 34782 8033
rect 34748 7931 34782 7965
rect 34845 7999 34879 8033
rect 34845 7931 34879 7965
rect 34929 8073 34963 8107
rect 34929 8002 34963 8036
rect 34929 7931 34963 7965
rect 35074 8067 35108 8101
rect 35074 7999 35108 8033
rect 35074 7931 35108 7965
rect 35158 8067 35192 8101
rect 35158 7999 35192 8033
rect 35158 7931 35192 7965
rect 35319 8067 35353 8101
rect 35319 7999 35353 8033
rect 35319 7931 35353 7965
rect 35403 8067 35437 8101
rect 35403 7999 35437 8033
rect 35403 7931 35437 7965
rect 35487 7999 35521 8033
rect 35487 7931 35521 7965
rect 35571 8067 35605 8101
rect 35571 7999 35605 8033
rect 35571 7931 35605 7965
rect 35655 7931 35689 7965
rect 30587 7771 30621 7805
rect 30587 7703 30621 7737
rect 30671 7755 30705 7789
rect 30755 7771 30789 7805
rect 30859 7779 30893 7813
rect 30943 7771 30977 7805
rect 31035 7766 31069 7800
rect 31274 7779 31308 7813
rect 30755 7703 30789 7737
rect 31274 7711 31308 7745
rect 31358 7771 31392 7805
rect 31453 7761 31487 7795
rect 31652 7771 31686 7805
rect 31776 7779 31810 7813
rect 31776 7708 31810 7742
rect 31776 7637 31810 7671
rect 31862 7749 31896 7783
rect 31862 7669 31896 7703
rect 31946 7773 31980 7807
rect 31946 7705 31980 7739
rect 32050 7779 32084 7813
rect 32050 7711 32084 7745
rect 32147 7779 32181 7813
rect 32147 7711 32181 7745
rect 31946 7637 31980 7671
rect 32147 7643 32181 7677
rect 32231 7779 32265 7813
rect 32231 7708 32265 7742
rect 32231 7637 32265 7671
rect 32376 7779 32410 7813
rect 32376 7711 32410 7745
rect 32376 7643 32410 7677
rect 32460 7779 32494 7813
rect 32460 7711 32494 7745
rect 32460 7643 32494 7677
rect 32621 7779 32655 7813
rect 32621 7711 32655 7745
rect 32621 7643 32655 7677
rect 32705 7779 32739 7813
rect 32705 7711 32739 7745
rect 32705 7643 32739 7677
rect 32789 7779 32823 7813
rect 32789 7711 32823 7745
rect 32873 7779 32907 7813
rect 32873 7711 32907 7745
rect 32873 7643 32907 7677
rect 32957 7779 32991 7813
rect 33285 7771 33319 7805
rect 33285 7703 33319 7737
rect 33369 7755 33403 7789
rect 33453 7771 33487 7805
rect 33557 7779 33591 7813
rect 33641 7771 33675 7805
rect 33733 7766 33767 7800
rect 33972 7779 34006 7813
rect 33453 7703 33487 7737
rect 33972 7711 34006 7745
rect 34056 7771 34090 7805
rect 34151 7761 34185 7795
rect 34350 7771 34384 7805
rect 34474 7779 34508 7813
rect 34474 7708 34508 7742
rect 34474 7637 34508 7671
rect 34560 7749 34594 7783
rect 34560 7669 34594 7703
rect 34644 7773 34678 7807
rect 34644 7705 34678 7739
rect 34748 7779 34782 7813
rect 34748 7711 34782 7745
rect 34845 7779 34879 7813
rect 34845 7711 34879 7745
rect 34644 7637 34678 7671
rect 34845 7643 34879 7677
rect 34929 7779 34963 7813
rect 34929 7708 34963 7742
rect 34929 7637 34963 7671
rect 35074 7779 35108 7813
rect 35074 7711 35108 7745
rect 35074 7643 35108 7677
rect 35158 7779 35192 7813
rect 35158 7711 35192 7745
rect 35158 7643 35192 7677
rect 35319 7779 35353 7813
rect 35319 7711 35353 7745
rect 35319 7643 35353 7677
rect 35403 7779 35437 7813
rect 35403 7711 35437 7745
rect 35403 7643 35437 7677
rect 35487 7779 35521 7813
rect 35487 7711 35521 7745
rect 35571 7779 35605 7813
rect 35571 7711 35605 7745
rect 35571 7643 35605 7677
rect 35655 7779 35689 7813
rect 30587 6919 30621 6953
rect 30587 6851 30621 6885
rect 30671 6867 30705 6901
rect 30755 6919 30789 6953
rect 30755 6851 30789 6885
rect 30859 6843 30893 6877
rect 30943 6851 30977 6885
rect 31035 6856 31069 6890
rect 31274 6911 31308 6945
rect 31274 6843 31308 6877
rect 31776 6985 31810 7019
rect 31358 6851 31392 6885
rect 31453 6861 31487 6895
rect 31652 6851 31686 6885
rect 31776 6914 31810 6948
rect 31776 6843 31810 6877
rect 31862 6953 31896 6987
rect 31862 6873 31896 6907
rect 31946 6985 31980 7019
rect 32147 6979 32181 7013
rect 31946 6917 31980 6951
rect 31946 6849 31980 6883
rect 32050 6911 32084 6945
rect 32050 6843 32084 6877
rect 32147 6911 32181 6945
rect 32147 6843 32181 6877
rect 32231 6985 32265 7019
rect 32231 6914 32265 6948
rect 32231 6843 32265 6877
rect 32376 6979 32410 7013
rect 32376 6911 32410 6945
rect 32376 6843 32410 6877
rect 32460 6979 32494 7013
rect 32460 6911 32494 6945
rect 32460 6843 32494 6877
rect 32621 6979 32655 7013
rect 32621 6911 32655 6945
rect 32621 6843 32655 6877
rect 32705 6979 32739 7013
rect 32705 6911 32739 6945
rect 32705 6843 32739 6877
rect 32789 6911 32823 6945
rect 32789 6843 32823 6877
rect 32873 6979 32907 7013
rect 32873 6911 32907 6945
rect 32873 6843 32907 6877
rect 32957 6843 32991 6877
rect 33285 6919 33319 6953
rect 33285 6851 33319 6885
rect 33369 6867 33403 6901
rect 33453 6919 33487 6953
rect 33453 6851 33487 6885
rect 33557 6843 33591 6877
rect 33641 6851 33675 6885
rect 33733 6856 33767 6890
rect 33972 6911 34006 6945
rect 33972 6843 34006 6877
rect 34474 6985 34508 7019
rect 34056 6851 34090 6885
rect 34151 6861 34185 6895
rect 34350 6851 34384 6885
rect 34474 6914 34508 6948
rect 34474 6843 34508 6877
rect 34560 6953 34594 6987
rect 34560 6873 34594 6907
rect 34644 6985 34678 7019
rect 34845 6979 34879 7013
rect 34644 6917 34678 6951
rect 34644 6849 34678 6883
rect 34748 6911 34782 6945
rect 34748 6843 34782 6877
rect 34845 6911 34879 6945
rect 34845 6843 34879 6877
rect 34929 6985 34963 7019
rect 34929 6914 34963 6948
rect 34929 6843 34963 6877
rect 35074 6979 35108 7013
rect 35074 6911 35108 6945
rect 35074 6843 35108 6877
rect 35158 6979 35192 7013
rect 35158 6911 35192 6945
rect 35158 6843 35192 6877
rect 35319 6979 35353 7013
rect 35319 6911 35353 6945
rect 35319 6843 35353 6877
rect 35403 6979 35437 7013
rect 35403 6911 35437 6945
rect 35403 6843 35437 6877
rect 35487 6911 35521 6945
rect 35487 6843 35521 6877
rect 35571 6979 35605 7013
rect 35571 6911 35605 6945
rect 35571 6843 35605 6877
rect 35655 6843 35689 6877
rect 30587 6683 30621 6717
rect 30587 6615 30621 6649
rect 30671 6667 30705 6701
rect 30755 6683 30789 6717
rect 30859 6691 30893 6725
rect 30943 6683 30977 6717
rect 31035 6678 31069 6712
rect 31274 6691 31308 6725
rect 30755 6615 30789 6649
rect 31274 6623 31308 6657
rect 31358 6683 31392 6717
rect 31453 6673 31487 6707
rect 31652 6683 31686 6717
rect 31776 6691 31810 6725
rect 31776 6620 31810 6654
rect 31776 6549 31810 6583
rect 31862 6661 31896 6695
rect 31862 6581 31896 6615
rect 31946 6685 31980 6719
rect 31946 6617 31980 6651
rect 32050 6691 32084 6725
rect 32050 6623 32084 6657
rect 32147 6691 32181 6725
rect 32147 6623 32181 6657
rect 31946 6549 31980 6583
rect 32147 6555 32181 6589
rect 32231 6691 32265 6725
rect 32231 6620 32265 6654
rect 32231 6549 32265 6583
rect 32376 6691 32410 6725
rect 32376 6623 32410 6657
rect 32376 6555 32410 6589
rect 32460 6691 32494 6725
rect 32460 6623 32494 6657
rect 32460 6555 32494 6589
rect 32621 6691 32655 6725
rect 32621 6623 32655 6657
rect 32621 6555 32655 6589
rect 32705 6691 32739 6725
rect 32705 6623 32739 6657
rect 32705 6555 32739 6589
rect 32789 6691 32823 6725
rect 32789 6623 32823 6657
rect 32873 6691 32907 6725
rect 32873 6623 32907 6657
rect 32873 6555 32907 6589
rect 32957 6691 32991 6725
rect 33285 6683 33319 6717
rect 33285 6615 33319 6649
rect 33369 6667 33403 6701
rect 33453 6683 33487 6717
rect 33557 6691 33591 6725
rect 33641 6683 33675 6717
rect 33733 6678 33767 6712
rect 33972 6691 34006 6725
rect 33453 6615 33487 6649
rect 33972 6623 34006 6657
rect 34056 6683 34090 6717
rect 34151 6673 34185 6707
rect 34350 6683 34384 6717
rect 34474 6691 34508 6725
rect 34474 6620 34508 6654
rect 34474 6549 34508 6583
rect 34560 6661 34594 6695
rect 34560 6581 34594 6615
rect 34644 6685 34678 6719
rect 34644 6617 34678 6651
rect 34748 6691 34782 6725
rect 34748 6623 34782 6657
rect 34845 6691 34879 6725
rect 34845 6623 34879 6657
rect 34644 6549 34678 6583
rect 34845 6555 34879 6589
rect 34929 6691 34963 6725
rect 34929 6620 34963 6654
rect 34929 6549 34963 6583
rect 35074 6691 35108 6725
rect 35074 6623 35108 6657
rect 35074 6555 35108 6589
rect 35158 6691 35192 6725
rect 35158 6623 35192 6657
rect 35158 6555 35192 6589
rect 35319 6691 35353 6725
rect 35319 6623 35353 6657
rect 35319 6555 35353 6589
rect 35403 6691 35437 6725
rect 35403 6623 35437 6657
rect 35403 6555 35437 6589
rect 35487 6691 35521 6725
rect 35487 6623 35521 6657
rect 35571 6691 35605 6725
rect 35571 6623 35605 6657
rect 35571 6555 35605 6589
rect 35655 6691 35689 6725
rect 30587 5831 30621 5865
rect 30587 5763 30621 5797
rect 30671 5779 30705 5813
rect 30755 5831 30789 5865
rect 30755 5763 30789 5797
rect 30859 5755 30893 5789
rect 30943 5763 30977 5797
rect 31035 5768 31069 5802
rect 31274 5823 31308 5857
rect 31274 5755 31308 5789
rect 31776 5897 31810 5931
rect 31358 5763 31392 5797
rect 31453 5773 31487 5807
rect 31652 5763 31686 5797
rect 31776 5826 31810 5860
rect 31776 5755 31810 5789
rect 31862 5865 31896 5899
rect 31862 5785 31896 5819
rect 31946 5897 31980 5931
rect 32147 5891 32181 5925
rect 31946 5829 31980 5863
rect 31946 5761 31980 5795
rect 32050 5823 32084 5857
rect 32050 5755 32084 5789
rect 32147 5823 32181 5857
rect 32147 5755 32181 5789
rect 32231 5897 32265 5931
rect 32231 5826 32265 5860
rect 32231 5755 32265 5789
rect 32376 5891 32410 5925
rect 32376 5823 32410 5857
rect 32376 5755 32410 5789
rect 32460 5891 32494 5925
rect 32460 5823 32494 5857
rect 32460 5755 32494 5789
rect 32621 5891 32655 5925
rect 32621 5823 32655 5857
rect 32621 5755 32655 5789
rect 32705 5891 32739 5925
rect 32705 5823 32739 5857
rect 32705 5755 32739 5789
rect 32789 5823 32823 5857
rect 32789 5755 32823 5789
rect 32873 5891 32907 5925
rect 32873 5823 32907 5857
rect 32873 5755 32907 5789
rect 32957 5755 32991 5789
rect 33285 5831 33319 5865
rect 33285 5763 33319 5797
rect 33369 5779 33403 5813
rect 33453 5831 33487 5865
rect 33453 5763 33487 5797
rect 33557 5755 33591 5789
rect 33641 5763 33675 5797
rect 33733 5768 33767 5802
rect 33972 5823 34006 5857
rect 33972 5755 34006 5789
rect 34474 5897 34508 5931
rect 34056 5763 34090 5797
rect 34151 5773 34185 5807
rect 34350 5763 34384 5797
rect 34474 5826 34508 5860
rect 34474 5755 34508 5789
rect 34560 5865 34594 5899
rect 34560 5785 34594 5819
rect 34644 5897 34678 5931
rect 34845 5891 34879 5925
rect 34644 5829 34678 5863
rect 34644 5761 34678 5795
rect 34748 5823 34782 5857
rect 34748 5755 34782 5789
rect 34845 5823 34879 5857
rect 34845 5755 34879 5789
rect 34929 5897 34963 5931
rect 34929 5826 34963 5860
rect 34929 5755 34963 5789
rect 35074 5891 35108 5925
rect 35074 5823 35108 5857
rect 35074 5755 35108 5789
rect 35158 5891 35192 5925
rect 35158 5823 35192 5857
rect 35158 5755 35192 5789
rect 35319 5891 35353 5925
rect 35319 5823 35353 5857
rect 35319 5755 35353 5789
rect 35403 5891 35437 5925
rect 35403 5823 35437 5857
rect 35403 5755 35437 5789
rect 35487 5823 35521 5857
rect 35487 5755 35521 5789
rect 35571 5891 35605 5925
rect 35571 5823 35605 5857
rect 35571 5755 35605 5789
rect 35655 5755 35689 5789
rect 9338 1356 9372 2932
rect 9796 1356 9830 2932
rect 10254 1356 10288 2932
rect 10712 1356 10746 2932
rect 11170 1356 11204 2932
rect 11628 1356 11662 2932
rect 12086 1356 12120 2932
rect 12544 1356 12578 2932
rect 13002 1356 13036 2932
rect 13460 1356 13494 2932
rect 13918 1356 13952 2932
rect 14376 1356 14410 2932
rect 14834 1356 14868 2932
rect 15292 1356 15326 2932
rect 15750 1356 15784 2932
rect 16208 1356 16242 2932
rect 16666 1356 16700 2932
rect 17124 1356 17158 2932
rect 17582 1356 17616 2932
rect 8779 -909 8813 267
rect 9237 -909 9271 267
rect 9695 -909 9729 267
rect 10153 -909 10187 267
rect 10611 -909 10645 267
rect 11069 -909 11103 267
rect 11527 -909 11561 267
rect 11985 -909 12019 267
rect 12443 -909 12477 267
rect 12901 -909 12935 267
rect 13359 -909 13393 267
rect 13779 -909 13813 267
rect 14237 -909 14271 267
rect 14695 -909 14729 267
rect 15153 -909 15187 267
rect 15611 -909 15645 267
rect 16069 -909 16103 267
rect 16527 -909 16561 267
rect 16985 -909 17019 267
rect 17443 -909 17477 267
rect 17901 -909 17935 267
rect 18359 -909 18393 267
rect 24338 1356 24372 2932
rect 24796 1356 24830 2932
rect 25254 1356 25288 2932
rect 25712 1356 25746 2932
rect 26170 1356 26204 2932
rect 26628 1356 26662 2932
rect 27086 1356 27120 2932
rect 27544 1356 27578 2932
rect 28002 1356 28036 2932
rect 28460 1356 28494 2932
rect 28918 1356 28952 2932
rect 29376 1356 29410 2932
rect 29834 1356 29868 2932
rect 30292 1356 30326 2932
rect 30750 1356 30784 2932
rect 31208 1356 31242 2932
rect 31666 1356 31700 2932
rect 32124 1356 32158 2932
rect 32582 1356 32616 2932
rect 23779 -909 23813 267
rect 24237 -909 24271 267
rect 24695 -909 24729 267
rect 25153 -909 25187 267
rect 25611 -909 25645 267
rect 26069 -909 26103 267
rect 26527 -909 26561 267
rect 26985 -909 27019 267
rect 27443 -909 27477 267
rect 27901 -909 27935 267
rect 28359 -909 28393 267
rect 28779 -909 28813 267
rect 29237 -909 29271 267
rect 29695 -909 29729 267
rect 30153 -909 30187 267
rect 30611 -909 30645 267
rect 31069 -909 31103 267
rect 31527 -909 31561 267
rect 31985 -909 32019 267
rect 32443 -909 32477 267
rect 32901 -909 32935 267
rect 33359 -909 33393 267
rect 12709 -9023 12743 -7847
rect 13167 -9023 13201 -7847
rect 13625 -9023 13659 -7847
rect 14083 -9023 14117 -7847
rect 14541 -9023 14575 -7847
rect 14999 -9023 15033 -7847
rect 15457 -9023 15491 -7847
rect 15915 -9023 15949 -7847
rect 16373 -9023 16407 -7847
rect 16831 -9023 16865 -7847
rect 17289 -9023 17323 -7847
rect 17709 -9023 17743 -7847
rect 18167 -9023 18201 -7847
rect 18625 -9023 18659 -7847
rect 19083 -9023 19117 -7847
rect 19541 -9023 19575 -7847
rect 19999 -9023 20033 -7847
rect 20457 -9023 20491 -7847
rect 20915 -9023 20949 -7847
rect 21373 -9023 21407 -7847
rect 21831 -9023 21865 -7847
rect 22289 -9023 22323 -7847
rect 13486 -11688 13520 -10112
rect 13944 -11688 13978 -10112
rect 14402 -11688 14436 -10112
rect 14860 -11688 14894 -10112
rect 15318 -11688 15352 -10112
rect 15776 -11688 15810 -10112
rect 16234 -11688 16268 -10112
rect 16692 -11688 16726 -10112
rect 17150 -11688 17184 -10112
rect 17608 -11688 17642 -10112
rect 18066 -11688 18100 -10112
rect 18524 -11688 18558 -10112
rect 18982 -11688 19016 -10112
rect 19440 -11688 19474 -10112
rect 19898 -11688 19932 -10112
rect 20356 -11688 20390 -10112
rect 20814 -11688 20848 -10112
rect 21272 -11688 21306 -10112
rect 21730 -11688 21764 -10112
rect 27709 -9023 27743 -7847
rect 28167 -9023 28201 -7847
rect 28625 -9023 28659 -7847
rect 29083 -9023 29117 -7847
rect 29541 -9023 29575 -7847
rect 29999 -9023 30033 -7847
rect 30457 -9023 30491 -7847
rect 30915 -9023 30949 -7847
rect 31373 -9023 31407 -7847
rect 31831 -9023 31865 -7847
rect 32289 -9023 32323 -7847
rect 32709 -9023 32743 -7847
rect 33167 -9023 33201 -7847
rect 33625 -9023 33659 -7847
rect 34083 -9023 34117 -7847
rect 34541 -9023 34575 -7847
rect 34999 -9023 35033 -7847
rect 35457 -9023 35491 -7847
rect 35915 -9023 35949 -7847
rect 36373 -9023 36407 -7847
rect 36831 -9023 36865 -7847
rect 37289 -9023 37323 -7847
rect 28486 -11688 28520 -10112
rect 28944 -11688 28978 -10112
rect 29402 -11688 29436 -10112
rect 29860 -11688 29894 -10112
rect 30318 -11688 30352 -10112
rect 30776 -11688 30810 -10112
rect 31234 -11688 31268 -10112
rect 31692 -11688 31726 -10112
rect 32150 -11688 32184 -10112
rect 32608 -11688 32642 -10112
rect 33066 -11688 33100 -10112
rect 33524 -11688 33558 -10112
rect 33982 -11688 34016 -10112
rect 34440 -11688 34474 -10112
rect 34898 -11688 34932 -10112
rect 35356 -11688 35390 -10112
rect 35814 -11688 35848 -10112
rect 36272 -11688 36306 -10112
rect 36730 -11688 36764 -10112
rect 9338 -16644 9372 -15068
rect 9796 -16644 9830 -15068
rect 10254 -16644 10288 -15068
rect 10712 -16644 10746 -15068
rect 11170 -16644 11204 -15068
rect 11628 -16644 11662 -15068
rect 12086 -16644 12120 -15068
rect 12544 -16644 12578 -15068
rect 13002 -16644 13036 -15068
rect 13460 -16644 13494 -15068
rect 13918 -16644 13952 -15068
rect 14376 -16644 14410 -15068
rect 14834 -16644 14868 -15068
rect 15292 -16644 15326 -15068
rect 15750 -16644 15784 -15068
rect 16208 -16644 16242 -15068
rect 16666 -16644 16700 -15068
rect 17124 -16644 17158 -15068
rect 17582 -16644 17616 -15068
rect 8779 -18909 8813 -17733
rect 9237 -18909 9271 -17733
rect 9695 -18909 9729 -17733
rect 10153 -18909 10187 -17733
rect 10611 -18909 10645 -17733
rect 11069 -18909 11103 -17733
rect 11527 -18909 11561 -17733
rect 11985 -18909 12019 -17733
rect 12443 -18909 12477 -17733
rect 12901 -18909 12935 -17733
rect 13359 -18909 13393 -17733
rect 13779 -18909 13813 -17733
rect 14237 -18909 14271 -17733
rect 14695 -18909 14729 -17733
rect 15153 -18909 15187 -17733
rect 15611 -18909 15645 -17733
rect 16069 -18909 16103 -17733
rect 16527 -18909 16561 -17733
rect 16985 -18909 17019 -17733
rect 17443 -18909 17477 -17733
rect 17901 -18909 17935 -17733
rect 18359 -18909 18393 -17733
rect 24338 -16644 24372 -15068
rect 24796 -16644 24830 -15068
rect 25254 -16644 25288 -15068
rect 25712 -16644 25746 -15068
rect 26170 -16644 26204 -15068
rect 26628 -16644 26662 -15068
rect 27086 -16644 27120 -15068
rect 27544 -16644 27578 -15068
rect 28002 -16644 28036 -15068
rect 28460 -16644 28494 -15068
rect 28918 -16644 28952 -15068
rect 29376 -16644 29410 -15068
rect 29834 -16644 29868 -15068
rect 30292 -16644 30326 -15068
rect 30750 -16644 30784 -15068
rect 31208 -16644 31242 -15068
rect 31666 -16644 31700 -15068
rect 32124 -16644 32158 -15068
rect 32582 -16644 32616 -15068
rect 23779 -18909 23813 -17733
rect 24237 -18909 24271 -17733
rect 24695 -18909 24729 -17733
rect 25153 -18909 25187 -17733
rect 25611 -18909 25645 -17733
rect 26069 -18909 26103 -17733
rect 26527 -18909 26561 -17733
rect 26985 -18909 27019 -17733
rect 27443 -18909 27477 -17733
rect 27901 -18909 27935 -17733
rect 28359 -18909 28393 -17733
rect 28779 -18909 28813 -17733
rect 29237 -18909 29271 -17733
rect 29695 -18909 29729 -17733
rect 30153 -18909 30187 -17733
rect 30611 -18909 30645 -17733
rect 31069 -18909 31103 -17733
rect 31527 -18909 31561 -17733
rect 31985 -18909 32019 -17733
rect 32443 -18909 32477 -17733
rect 32901 -18909 32935 -17733
rect 33359 -18909 33393 -17733
<< psubdiff >>
rect 24049 14047 24145 14081
rect 24989 14047 25085 14081
rect 24049 13985 24083 14047
rect 25051 13985 25085 14047
rect 24049 13567 24083 13629
rect 25051 13567 25085 13629
rect 24049 13533 24145 13567
rect 24989 13533 25085 13567
rect 25171 14047 25267 14081
rect 26885 14047 26981 14081
rect 25171 13985 25205 14047
rect 26947 13985 26981 14047
rect 25171 13567 25205 13629
rect 26947 13567 26981 13629
rect 25171 13533 25267 13567
rect 26885 13533 26981 13567
rect 23334 13220 23496 13320
rect 32616 13220 32778 13320
rect 23334 13158 23434 13220
rect 32678 13158 32778 13220
rect 23334 11156 23434 11218
rect 32678 11156 32778 11218
rect 23334 11056 23496 11156
rect 32616 11056 32778 11156
rect 12960 10634 13122 10734
rect 21822 10634 21984 10734
rect 12960 10572 13060 10634
rect 21884 10572 21984 10634
rect 12960 9034 13060 9096
rect 21884 9034 21984 9096
rect 12960 8934 13122 9034
rect 21822 8934 21984 9034
rect 23542 10634 23704 10734
rect 28824 10634 28986 10734
rect 23542 10572 23642 10634
rect 28886 10572 28986 10634
rect 23542 8954 23642 9016
rect 28886 8954 28986 9016
rect 23542 8854 23704 8954
rect 28824 8854 28986 8954
rect 30239 8561 30273 8585
rect 30239 8480 30273 8527
rect 33139 8561 33173 8585
rect 33139 8480 33173 8527
rect 36013 8561 36047 8585
rect 36013 8480 36047 8527
rect 30239 8305 30273 8352
rect 30239 8247 30273 8271
rect 36013 8305 36047 8352
rect 36013 8247 36047 8271
rect 30239 7473 30273 7497
rect 30239 7392 30273 7439
rect 36013 7473 36047 7497
rect 36013 7392 36047 7439
rect 30239 7217 30273 7264
rect 30239 7159 30273 7183
rect 36013 7217 36047 7264
rect 36013 7159 36047 7183
rect 30239 6385 30273 6409
rect 30239 6304 30273 6351
rect 36013 6385 36047 6409
rect 36013 6304 36047 6351
rect 30239 6129 30273 6176
rect 30239 6071 30273 6095
rect 36013 6129 36047 6176
rect 36013 6071 36047 6095
rect 8352 -1784 8514 -1684
rect 18634 -1784 18796 -1684
rect 8352 -1846 8452 -1784
rect 18696 -1846 18796 -1784
rect 8352 -4048 8452 -3986
rect 18696 -4048 18796 -3986
rect 8352 -4148 8514 -4048
rect 18634 -4148 18796 -4048
rect 23352 -1784 23514 -1684
rect 33634 -1784 33796 -1684
rect 23352 -1846 23452 -1784
rect 33696 -1846 33796 -1784
rect 23352 -4048 23452 -3986
rect 33696 -4048 33796 -3986
rect 23352 -4148 23514 -4048
rect 33634 -4148 33796 -4048
rect 12306 -4708 12468 -4608
rect 22588 -4708 22750 -4608
rect 12306 -4770 12406 -4708
rect 22650 -4770 22750 -4708
rect 12306 -6972 12406 -6910
rect 22650 -6972 22750 -6910
rect 12306 -7072 12468 -6972
rect 22588 -7072 22750 -6972
rect 27306 -4708 27468 -4608
rect 37588 -4708 37750 -4608
rect 27306 -4770 27406 -4708
rect 37650 -4770 37750 -4708
rect 27306 -6972 27406 -6910
rect 37650 -6972 37750 -6910
rect 27306 -7072 27468 -6972
rect 37588 -7072 37750 -6972
rect 8352 -19784 8514 -19684
rect 18634 -19784 18796 -19684
rect 8352 -19846 8452 -19784
rect 18696 -19846 18796 -19784
rect 8352 -22048 8452 -21986
rect 18696 -22048 18796 -21986
rect 8352 -22148 8514 -22048
rect 18634 -22148 18796 -22048
rect 23352 -19784 23514 -19684
rect 33634 -19784 33796 -19684
rect 23352 -19846 23452 -19784
rect 33696 -19846 33796 -19784
rect 23352 -22048 23452 -21986
rect 33696 -22048 33796 -21986
rect 23352 -22148 23514 -22048
rect 33634 -22148 33796 -22048
<< nsubdiff >>
rect 23334 17400 23496 17500
rect 32616 17400 32778 17500
rect 23334 17338 23434 17400
rect 32678 17338 32778 17400
rect 23334 15296 23434 15358
rect 32678 15296 32778 15358
rect 23334 15196 23496 15296
rect 32616 15196 32778 15296
rect 24049 14943 24145 14977
rect 24989 14943 25085 14977
rect 24049 14881 24083 14943
rect 25051 14881 25085 14943
rect 24049 14245 24083 14307
rect 25051 14245 25085 14307
rect 24049 14211 24145 14245
rect 24989 14211 25085 14245
rect 25171 14943 25267 14977
rect 26885 14943 26981 14977
rect 25171 14881 25205 14943
rect 26947 14881 26981 14943
rect 25171 14245 25205 14307
rect 26947 14245 26981 14307
rect 25171 14211 25267 14245
rect 26885 14211 26981 14245
rect 30239 8872 30273 8896
rect 30239 8779 30273 8838
rect 30239 8721 30273 8745
rect 12960 8598 13122 8698
rect 21822 8598 21984 8698
rect 12960 8536 13060 8598
rect 21884 8536 21984 8598
rect 12960 4866 13060 4928
rect 21884 4866 21984 4928
rect 12960 4766 13122 4866
rect 21822 4766 21984 4866
rect 23542 8518 23704 8618
rect 28824 8518 28986 8618
rect 23542 8456 23642 8518
rect 28886 8456 28986 8518
rect 23542 4866 23642 4928
rect 33139 8872 33173 8896
rect 33139 8779 33173 8838
rect 33139 8721 33173 8745
rect 36013 8872 36047 8896
rect 36013 8779 36047 8838
rect 36013 8721 36047 8745
rect 30239 8087 30273 8111
rect 30239 7994 30273 8053
rect 30239 7936 30273 7960
rect 36013 8087 36047 8111
rect 36013 7994 36047 8053
rect 36013 7936 36047 7960
rect 30239 7784 30273 7808
rect 30239 7691 30273 7750
rect 30239 7633 30273 7657
rect 36013 7784 36047 7808
rect 36013 7691 36047 7750
rect 36013 7633 36047 7657
rect 30239 6999 30273 7023
rect 30239 6906 30273 6965
rect 30239 6848 30273 6872
rect 36013 6999 36047 7023
rect 36013 6906 36047 6965
rect 36013 6848 36047 6872
rect 30239 6696 30273 6720
rect 30239 6603 30273 6662
rect 30239 6545 30273 6569
rect 36013 6696 36047 6720
rect 36013 6603 36047 6662
rect 36013 6545 36047 6569
rect 30239 5911 30273 5935
rect 30239 5818 30273 5877
rect 30239 5760 30273 5784
rect 36013 5911 36047 5935
rect 36013 5818 36047 5877
rect 36013 5760 36047 5784
rect 28886 4866 28986 4928
rect 23542 4766 23704 4866
rect 28824 4766 28986 4866
rect 8352 4296 8514 4396
rect 18634 4296 18796 4396
rect 8352 4234 8452 4296
rect 18696 4234 18796 4296
rect 8352 -1348 8452 -1286
rect 18696 -1348 18796 -1286
rect 8352 -1448 8514 -1348
rect 18634 -1448 18796 -1348
rect 23352 4296 23514 4396
rect 33634 4296 33796 4396
rect 23352 4234 23452 4296
rect 33696 4234 33796 4296
rect 23352 -1348 23452 -1286
rect 33696 -1348 33796 -1286
rect 23352 -1448 23514 -1348
rect 33634 -1448 33796 -1348
rect 12306 -7408 12468 -7308
rect 22588 -7408 22750 -7308
rect 12306 -7470 12406 -7408
rect 22650 -7470 22750 -7408
rect 12306 -13052 12406 -12990
rect 22650 -13052 22750 -12990
rect 12306 -13152 12468 -13052
rect 22588 -13152 22750 -13052
rect 27306 -7408 27468 -7308
rect 37588 -7408 37750 -7308
rect 27306 -7470 27406 -7408
rect 37650 -7470 37750 -7408
rect 27306 -13052 27406 -12990
rect 37650 -13052 37750 -12990
rect 27306 -13152 27468 -13052
rect 37588 -13152 37750 -13052
rect 8352 -13704 8514 -13604
rect 18634 -13704 18796 -13604
rect 8352 -13766 8452 -13704
rect 18696 -13766 18796 -13704
rect 8352 -19348 8452 -19286
rect 18696 -19348 18796 -19286
rect 8352 -19448 8514 -19348
rect 18634 -19448 18796 -19348
rect 23352 -13704 23514 -13604
rect 33634 -13704 33796 -13604
rect 23352 -13766 23452 -13704
rect 33696 -13766 33796 -13704
rect 23352 -19348 23452 -19286
rect 33696 -19348 33796 -19286
rect 23352 -19448 23514 -19348
rect 33634 -19448 33796 -19348
<< psubdiffcont >>
rect 24145 14047 24989 14081
rect 24049 13629 24083 13985
rect 25051 13629 25085 13985
rect 24145 13533 24989 13567
rect 25267 14047 26885 14081
rect 25171 13629 25205 13985
rect 26947 13629 26981 13985
rect 25267 13533 26885 13567
rect 23496 13220 32616 13320
rect 23334 11218 23434 13158
rect 32678 11218 32778 13158
rect 23496 11056 32616 11156
rect 13122 10634 21822 10734
rect 12960 9096 13060 10572
rect 21884 9096 21984 10572
rect 13122 8934 21822 9034
rect 23704 10634 28824 10734
rect 23542 9016 23642 10572
rect 28886 9016 28986 10572
rect 23704 8854 28824 8954
rect 30239 8527 30273 8561
rect 33139 8527 33173 8561
rect 36013 8527 36047 8561
rect 30239 8271 30273 8305
rect 36013 8271 36047 8305
rect 30239 7439 30273 7473
rect 36013 7439 36047 7473
rect 30239 7183 30273 7217
rect 36013 7183 36047 7217
rect 30239 6351 30273 6385
rect 36013 6351 36047 6385
rect 30239 6095 30273 6129
rect 36013 6095 36047 6129
rect 8514 -1784 18634 -1684
rect 8352 -3986 8452 -1846
rect 18696 -3986 18796 -1846
rect 8514 -4148 18634 -4048
rect 23514 -1784 33634 -1684
rect 23352 -3986 23452 -1846
rect 33696 -3986 33796 -1846
rect 23514 -4148 33634 -4048
rect 12468 -4708 22588 -4608
rect 12306 -6910 12406 -4770
rect 22650 -6910 22750 -4770
rect 12468 -7072 22588 -6972
rect 27468 -4708 37588 -4608
rect 27306 -6910 27406 -4770
rect 37650 -6910 37750 -4770
rect 27468 -7072 37588 -6972
rect 8514 -19784 18634 -19684
rect 8352 -21986 8452 -19846
rect 18696 -21986 18796 -19846
rect 8514 -22148 18634 -22048
rect 23514 -19784 33634 -19684
rect 23352 -21986 23452 -19846
rect 33696 -21986 33796 -19846
rect 23514 -22148 33634 -22048
<< nsubdiffcont >>
rect 23496 17400 32616 17500
rect 23334 15358 23434 17338
rect 32678 15358 32778 17338
rect 23496 15196 32616 15296
rect 24145 14943 24989 14977
rect 24049 14307 24083 14881
rect 25051 14307 25085 14881
rect 24145 14211 24989 14245
rect 25267 14943 26885 14977
rect 25171 14307 25205 14881
rect 26947 14307 26981 14881
rect 25267 14211 26885 14245
rect 30239 8838 30273 8872
rect 30239 8745 30273 8779
rect 13122 8598 21822 8698
rect 12960 4928 13060 8536
rect 21884 4928 21984 8536
rect 13122 4766 21822 4866
rect 23704 8518 28824 8618
rect 23542 4928 23642 8456
rect 28886 4928 28986 8456
rect 33139 8838 33173 8872
rect 33139 8745 33173 8779
rect 36013 8838 36047 8872
rect 36013 8745 36047 8779
rect 30239 8053 30273 8087
rect 30239 7960 30273 7994
rect 36013 8053 36047 8087
rect 36013 7960 36047 7994
rect 30239 7750 30273 7784
rect 30239 7657 30273 7691
rect 36013 7750 36047 7784
rect 36013 7657 36047 7691
rect 30239 6965 30273 6999
rect 30239 6872 30273 6906
rect 36013 6965 36047 6999
rect 36013 6872 36047 6906
rect 30239 6662 30273 6696
rect 30239 6569 30273 6603
rect 36013 6662 36047 6696
rect 36013 6569 36047 6603
rect 30239 5877 30273 5911
rect 30239 5784 30273 5818
rect 36013 5877 36047 5911
rect 36013 5784 36047 5818
rect 23704 4766 28824 4866
rect 8514 4296 18634 4396
rect 8352 -1286 8452 4234
rect 18696 -1286 18796 4234
rect 8514 -1448 18634 -1348
rect 23514 4296 33634 4396
rect 23352 -1286 23452 4234
rect 33696 -1286 33796 4234
rect 23514 -1448 33634 -1348
rect 12468 -7408 22588 -7308
rect 12306 -12990 12406 -7470
rect 22650 -12990 22750 -7470
rect 12468 -13152 22588 -13052
rect 27468 -7408 37588 -7308
rect 27306 -12990 27406 -7470
rect 37650 -12990 37750 -7470
rect 27468 -13152 37588 -13052
rect 8514 -13704 18634 -13604
rect 8352 -19286 8452 -13766
rect 18696 -19286 18796 -13766
rect 8514 -19448 18634 -19348
rect 23514 -13704 33634 -13604
rect 23352 -19286 23452 -13766
rect 33696 -19286 33796 -13766
rect 23514 -19448 33634 -19348
<< poly >>
rect 24014 16515 24430 16531
rect 24014 16498 24030 16515
rect 23822 16481 24030 16498
rect 24414 16498 24430 16515
rect 24872 16515 25288 16531
rect 24872 16498 24888 16515
rect 24414 16481 24622 16498
rect 23822 16434 24622 16481
rect 24680 16481 24888 16498
rect 25272 16498 25288 16515
rect 25730 16515 26146 16531
rect 25730 16498 25746 16515
rect 25272 16481 25480 16498
rect 24680 16434 25480 16481
rect 25538 16481 25746 16498
rect 26130 16498 26146 16515
rect 26588 16515 27004 16531
rect 26588 16498 26604 16515
rect 26130 16481 26338 16498
rect 25538 16434 26338 16481
rect 26396 16481 26604 16498
rect 26988 16498 27004 16515
rect 27446 16515 27862 16531
rect 27446 16498 27462 16515
rect 26988 16481 27196 16498
rect 26396 16434 27196 16481
rect 27254 16481 27462 16498
rect 27846 16498 27862 16515
rect 28304 16515 28720 16531
rect 28304 16498 28320 16515
rect 27846 16481 28054 16498
rect 27254 16434 28054 16481
rect 28112 16481 28320 16498
rect 28704 16498 28720 16515
rect 29162 16515 29578 16531
rect 29162 16498 29178 16515
rect 28704 16481 28912 16498
rect 28112 16434 28912 16481
rect 28970 16481 29178 16498
rect 29562 16498 29578 16515
rect 30020 16515 30436 16531
rect 30020 16498 30036 16515
rect 29562 16481 29770 16498
rect 28970 16434 29770 16481
rect 29828 16481 30036 16498
rect 30420 16498 30436 16515
rect 30878 16515 31294 16531
rect 30878 16498 30894 16515
rect 30420 16481 30628 16498
rect 29828 16434 30628 16481
rect 30686 16481 30894 16498
rect 31278 16498 31294 16515
rect 31736 16515 32152 16531
rect 31736 16498 31752 16515
rect 31278 16481 31486 16498
rect 30686 16434 31486 16481
rect 31544 16481 31752 16498
rect 32136 16498 32152 16515
rect 32136 16481 32344 16498
rect 31544 16434 32344 16481
rect 23822 16187 24622 16234
rect 23822 16170 24030 16187
rect 24014 16153 24030 16170
rect 24414 16170 24622 16187
rect 24680 16187 25480 16234
rect 24680 16170 24888 16187
rect 24414 16153 24430 16170
rect 24014 16137 24430 16153
rect 24872 16153 24888 16170
rect 25272 16170 25480 16187
rect 25538 16187 26338 16234
rect 25538 16170 25746 16187
rect 25272 16153 25288 16170
rect 24872 16137 25288 16153
rect 25730 16153 25746 16170
rect 26130 16170 26338 16187
rect 26396 16187 27196 16234
rect 26396 16170 26604 16187
rect 26130 16153 26146 16170
rect 25730 16137 26146 16153
rect 26588 16153 26604 16170
rect 26988 16170 27196 16187
rect 27254 16187 28054 16234
rect 27254 16170 27462 16187
rect 26988 16153 27004 16170
rect 26588 16137 27004 16153
rect 27446 16153 27462 16170
rect 27846 16170 28054 16187
rect 28112 16187 28912 16234
rect 28112 16170 28320 16187
rect 27846 16153 27862 16170
rect 27446 16137 27862 16153
rect 28304 16153 28320 16170
rect 28704 16170 28912 16187
rect 28970 16187 29770 16234
rect 28970 16170 29178 16187
rect 28704 16153 28720 16170
rect 28304 16137 28720 16153
rect 29162 16153 29178 16170
rect 29562 16170 29770 16187
rect 29828 16187 30628 16234
rect 29828 16170 30036 16187
rect 29562 16153 29578 16170
rect 29162 16137 29578 16153
rect 30020 16153 30036 16170
rect 30420 16170 30628 16187
rect 30686 16187 31486 16234
rect 30686 16170 30894 16187
rect 30420 16153 30436 16170
rect 30020 16137 30436 16153
rect 30878 16153 30894 16170
rect 31278 16170 31486 16187
rect 31544 16187 32344 16234
rect 31544 16170 31752 16187
rect 31278 16153 31294 16170
rect 30878 16137 31294 16153
rect 31736 16153 31752 16170
rect 32136 16170 32344 16187
rect 32136 16153 32152 16170
rect 31736 16137 32152 16153
rect 24014 15915 24430 15931
rect 24014 15898 24030 15915
rect 23822 15881 24030 15898
rect 24414 15898 24430 15915
rect 24872 15915 25288 15931
rect 24872 15898 24888 15915
rect 24414 15881 24622 15898
rect 23822 15834 24622 15881
rect 24680 15881 24888 15898
rect 25272 15898 25288 15915
rect 25730 15915 26146 15931
rect 25730 15898 25746 15915
rect 25272 15881 25480 15898
rect 24680 15834 25480 15881
rect 25538 15881 25746 15898
rect 26130 15898 26146 15915
rect 26588 15915 27004 15931
rect 26588 15898 26604 15915
rect 26130 15881 26338 15898
rect 25538 15834 26338 15881
rect 26396 15881 26604 15898
rect 26988 15898 27004 15915
rect 27446 15915 27862 15931
rect 27446 15898 27462 15915
rect 26988 15881 27196 15898
rect 26396 15834 27196 15881
rect 27254 15881 27462 15898
rect 27846 15898 27862 15915
rect 28304 15915 28720 15931
rect 28304 15898 28320 15915
rect 27846 15881 28054 15898
rect 27254 15834 28054 15881
rect 28112 15881 28320 15898
rect 28704 15898 28720 15915
rect 29162 15915 29578 15931
rect 29162 15898 29178 15915
rect 28704 15881 28912 15898
rect 28112 15834 28912 15881
rect 28970 15881 29178 15898
rect 29562 15898 29578 15915
rect 30020 15915 30436 15931
rect 30020 15898 30036 15915
rect 29562 15881 29770 15898
rect 28970 15834 29770 15881
rect 29828 15881 30036 15898
rect 30420 15898 30436 15915
rect 30878 15915 31294 15931
rect 30878 15898 30894 15915
rect 30420 15881 30628 15898
rect 29828 15834 30628 15881
rect 30686 15881 30894 15898
rect 31278 15898 31294 15915
rect 31736 15915 32152 15931
rect 31736 15898 31752 15915
rect 31278 15881 31486 15898
rect 30686 15834 31486 15881
rect 31544 15881 31752 15898
rect 32136 15898 32152 15915
rect 32136 15881 32344 15898
rect 31544 15834 32344 15881
rect 23822 15587 24622 15634
rect 23822 15570 24030 15587
rect 24014 15553 24030 15570
rect 24414 15570 24622 15587
rect 24680 15587 25480 15634
rect 24680 15570 24888 15587
rect 24414 15553 24430 15570
rect 24014 15537 24430 15553
rect 24872 15553 24888 15570
rect 25272 15570 25480 15587
rect 25538 15587 26338 15634
rect 25538 15570 25746 15587
rect 25272 15553 25288 15570
rect 24872 15537 25288 15553
rect 25730 15553 25746 15570
rect 26130 15570 26338 15587
rect 26396 15587 27196 15634
rect 26396 15570 26604 15587
rect 26130 15553 26146 15570
rect 25730 15537 26146 15553
rect 26588 15553 26604 15570
rect 26988 15570 27196 15587
rect 27254 15587 28054 15634
rect 27254 15570 27462 15587
rect 26988 15553 27004 15570
rect 26588 15537 27004 15553
rect 27446 15553 27462 15570
rect 27846 15570 28054 15587
rect 28112 15587 28912 15634
rect 28112 15570 28320 15587
rect 27846 15553 27862 15570
rect 27446 15537 27862 15553
rect 28304 15553 28320 15570
rect 28704 15570 28912 15587
rect 28970 15587 29770 15634
rect 28970 15570 29178 15587
rect 28704 15553 28720 15570
rect 28304 15537 28720 15553
rect 29162 15553 29178 15570
rect 29562 15570 29770 15587
rect 29828 15587 30628 15634
rect 29828 15570 30036 15587
rect 29562 15553 29578 15570
rect 29162 15537 29578 15553
rect 30020 15553 30036 15570
rect 30420 15570 30628 15587
rect 30686 15587 31486 15634
rect 30686 15570 30894 15587
rect 30420 15553 30436 15570
rect 30020 15537 30436 15553
rect 30878 15553 30894 15570
rect 31278 15570 31486 15587
rect 31544 15587 32344 15634
rect 31544 15570 31752 15587
rect 31278 15553 31294 15570
rect 30878 15537 31294 15553
rect 31736 15553 31752 15570
rect 32136 15570 32344 15587
rect 32136 15553 32152 15570
rect 31736 15537 32152 15553
rect 24243 14875 24375 14891
rect 24243 14858 24259 14875
rect 24209 14841 24259 14858
rect 24359 14858 24375 14875
rect 24501 14875 24633 14891
rect 24501 14858 24517 14875
rect 24359 14841 24409 14858
rect 24209 14794 24409 14841
rect 24467 14841 24517 14858
rect 24617 14858 24633 14875
rect 24759 14875 24891 14891
rect 24759 14858 24775 14875
rect 24617 14841 24667 14858
rect 24467 14794 24667 14841
rect 24725 14841 24775 14858
rect 24875 14858 24891 14875
rect 24875 14841 24925 14858
rect 24725 14794 24925 14841
rect 24209 14347 24409 14394
rect 24209 14330 24259 14347
rect 24243 14313 24259 14330
rect 24359 14330 24409 14347
rect 24467 14347 24667 14394
rect 24467 14330 24517 14347
rect 24359 14313 24375 14330
rect 24243 14297 24375 14313
rect 24501 14313 24517 14330
rect 24617 14330 24667 14347
rect 24725 14347 24925 14394
rect 24725 14330 24775 14347
rect 24617 14313 24633 14330
rect 24501 14297 24633 14313
rect 24759 14313 24775 14330
rect 24875 14330 24925 14347
rect 24875 14313 24891 14330
rect 24759 14297 24891 14313
rect 25365 14875 25497 14891
rect 25365 14858 25381 14875
rect 25331 14841 25381 14858
rect 25481 14858 25497 14875
rect 25623 14875 25755 14891
rect 25623 14858 25639 14875
rect 25481 14841 25531 14858
rect 25331 14794 25531 14841
rect 25589 14841 25639 14858
rect 25739 14858 25755 14875
rect 25881 14875 26013 14891
rect 25881 14858 25897 14875
rect 25739 14841 25789 14858
rect 25589 14794 25789 14841
rect 25847 14841 25897 14858
rect 25997 14858 26013 14875
rect 26139 14875 26271 14891
rect 26139 14858 26155 14875
rect 25997 14841 26047 14858
rect 25847 14794 26047 14841
rect 26105 14841 26155 14858
rect 26255 14858 26271 14875
rect 26397 14875 26529 14891
rect 26397 14858 26413 14875
rect 26255 14841 26305 14858
rect 26105 14794 26305 14841
rect 26363 14841 26413 14858
rect 26513 14858 26529 14875
rect 26655 14875 26787 14891
rect 26655 14858 26671 14875
rect 26513 14841 26563 14858
rect 26363 14794 26563 14841
rect 26621 14841 26671 14858
rect 26771 14858 26787 14875
rect 26771 14841 26821 14858
rect 26621 14794 26821 14841
rect 25331 14347 25531 14394
rect 25331 14330 25381 14347
rect 25365 14313 25381 14330
rect 25481 14330 25531 14347
rect 25589 14347 25789 14394
rect 25589 14330 25639 14347
rect 25481 14313 25497 14330
rect 25365 14297 25497 14313
rect 25623 14313 25639 14330
rect 25739 14330 25789 14347
rect 25847 14347 26047 14394
rect 25847 14330 25897 14347
rect 25739 14313 25755 14330
rect 25623 14297 25755 14313
rect 25881 14313 25897 14330
rect 25997 14330 26047 14347
rect 26105 14347 26305 14394
rect 26105 14330 26155 14347
rect 25997 14313 26013 14330
rect 25881 14297 26013 14313
rect 26139 14313 26155 14330
rect 26255 14330 26305 14347
rect 26363 14347 26563 14394
rect 26363 14330 26413 14347
rect 26255 14313 26271 14330
rect 26139 14297 26271 14313
rect 26397 14313 26413 14330
rect 26513 14330 26563 14347
rect 26621 14347 26821 14394
rect 26621 14330 26671 14347
rect 26513 14313 26529 14330
rect 26397 14297 26529 14313
rect 26655 14313 26671 14330
rect 26771 14330 26821 14347
rect 26771 14313 26787 14330
rect 26655 14297 26787 14313
rect 27339 14405 27369 14431
rect 27423 14405 27453 14431
rect 27690 14411 27720 14437
rect 27782 14411 27812 14437
rect 27881 14411 27911 14437
rect 28021 14411 28051 14437
rect 28118 14411 28148 14437
rect 28315 14411 28345 14437
rect 28414 14411 28444 14437
rect 28500 14411 28530 14437
rect 28584 14411 28614 14437
rect 28692 14411 28722 14437
rect 28776 14411 28806 14437
rect 28940 14411 28970 14437
rect 29159 14411 29189 14437
rect 29256 14411 29286 14437
rect 29496 14411 29526 14437
rect 29735 14411 29765 14437
rect 29819 14411 29849 14437
rect 30054 14411 30084 14437
rect 30294 14411 30324 14437
rect 30391 14411 30421 14437
rect 30610 14411 30640 14437
rect 30774 14411 30804 14437
rect 30858 14411 30888 14437
rect 30966 14411 30996 14437
rect 31050 14411 31080 14437
rect 31136 14411 31166 14437
rect 31235 14411 31265 14437
rect 31432 14411 31462 14437
rect 31529 14411 31559 14437
rect 31669 14411 31699 14437
rect 31768 14411 31798 14437
rect 31860 14411 31890 14437
rect 27339 14262 27369 14277
rect 27306 14232 27369 14262
rect 27306 14179 27336 14232
rect 27423 14188 27453 14277
rect 27690 14240 27720 14327
rect 27782 14289 27812 14327
rect 27282 14163 27336 14179
rect 27282 14129 27292 14163
rect 27326 14129 27336 14163
rect 27378 14178 27453 14188
rect 27378 14144 27394 14178
rect 27428 14144 27453 14178
rect 27591 14224 27720 14240
rect 27766 14279 27832 14289
rect 27766 14245 27782 14279
rect 27816 14245 27832 14279
rect 27766 14235 27832 14245
rect 27591 14190 27601 14224
rect 27635 14210 27720 14224
rect 27635 14190 27708 14210
rect 27881 14193 27911 14327
rect 28021 14269 28051 14327
rect 28021 14253 28076 14269
rect 28021 14219 28031 14253
rect 28065 14219 28076 14253
rect 28021 14203 28076 14219
rect 27591 14174 27708 14190
rect 27378 14134 27453 14144
rect 27282 14113 27336 14129
rect 27306 14090 27336 14113
rect 24243 13979 24375 13995
rect 24243 13962 24259 13979
rect 24209 13945 24259 13962
rect 24359 13962 24375 13979
rect 24501 13979 24633 13995
rect 24501 13962 24517 13979
rect 24359 13945 24409 13962
rect 24209 13907 24409 13945
rect 24467 13945 24517 13962
rect 24617 13962 24633 13979
rect 24759 13979 24891 13995
rect 24759 13962 24775 13979
rect 24617 13945 24667 13962
rect 24467 13907 24667 13945
rect 24725 13945 24775 13962
rect 24875 13962 24891 13979
rect 24875 13945 24925 13962
rect 24725 13907 24925 13945
rect 24209 13669 24409 13707
rect 24209 13652 24259 13669
rect 24243 13635 24259 13652
rect 24359 13652 24409 13669
rect 24467 13669 24667 13707
rect 24467 13652 24517 13669
rect 24359 13635 24375 13652
rect 24243 13619 24375 13635
rect 24501 13635 24517 13652
rect 24617 13652 24667 13669
rect 24725 13669 24925 13707
rect 24725 13652 24775 13669
rect 24617 13635 24633 13652
rect 24501 13619 24633 13635
rect 24759 13635 24775 13652
rect 24875 13652 24925 13669
rect 24875 13635 24891 13652
rect 24759 13619 24891 13635
rect 27306 14060 27369 14090
rect 25365 13979 25497 13995
rect 25365 13962 25381 13979
rect 25331 13945 25381 13962
rect 25481 13962 25497 13979
rect 25623 13979 25755 13995
rect 25623 13962 25639 13979
rect 25481 13945 25531 13962
rect 25331 13907 25531 13945
rect 25589 13945 25639 13962
rect 25739 13962 25755 13979
rect 25881 13979 26013 13995
rect 25881 13962 25897 13979
rect 25739 13945 25789 13962
rect 25589 13907 25789 13945
rect 25847 13945 25897 13962
rect 25997 13962 26013 13979
rect 26139 13979 26271 13995
rect 26139 13962 26155 13979
rect 25997 13945 26047 13962
rect 25847 13907 26047 13945
rect 26105 13945 26155 13962
rect 26255 13962 26271 13979
rect 26397 13979 26529 13995
rect 26397 13962 26413 13979
rect 26255 13945 26305 13962
rect 26105 13907 26305 13945
rect 26363 13945 26413 13962
rect 26513 13962 26529 13979
rect 26655 13979 26787 13995
rect 26655 13962 26671 13979
rect 26513 13945 26563 13962
rect 26363 13907 26563 13945
rect 26621 13945 26671 13962
rect 26771 13962 26787 13979
rect 27339 14045 27369 14060
rect 27423 14045 27453 14134
rect 27678 14045 27708 14174
rect 27773 14163 27911 14193
rect 27773 14133 27804 14163
rect 27750 14117 27804 14133
rect 27750 14083 27760 14117
rect 27794 14083 27804 14117
rect 27750 14067 27804 14083
rect 27846 14111 27912 14121
rect 27846 14077 27862 14111
rect 27896 14077 27912 14111
rect 27846 14067 27912 14077
rect 26771 13945 26821 13962
rect 26621 13907 26821 13945
rect 25331 13669 25531 13707
rect 25331 13652 25381 13669
rect 25365 13635 25381 13652
rect 25481 13652 25531 13669
rect 25589 13669 25789 13707
rect 25589 13652 25639 13669
rect 25481 13635 25497 13652
rect 25365 13619 25497 13635
rect 25623 13635 25639 13652
rect 25739 13652 25789 13669
rect 25847 13669 26047 13707
rect 25847 13652 25897 13669
rect 25739 13635 25755 13652
rect 25623 13619 25755 13635
rect 25881 13635 25897 13652
rect 25997 13652 26047 13669
rect 26105 13669 26305 13707
rect 26105 13652 26155 13669
rect 25997 13635 26013 13652
rect 25881 13619 26013 13635
rect 26139 13635 26155 13652
rect 26255 13652 26305 13669
rect 26363 13669 26563 13707
rect 26363 13652 26413 13669
rect 26255 13635 26271 13652
rect 26139 13619 26271 13635
rect 26397 13635 26413 13652
rect 26513 13652 26563 13669
rect 26621 13669 26821 13707
rect 26621 13652 26671 13669
rect 26513 13635 26529 13652
rect 26397 13619 26529 13635
rect 26655 13635 26671 13652
rect 26771 13652 26821 13669
rect 26771 13635 26787 13652
rect 26655 13619 26787 13635
rect 27773 14033 27803 14067
rect 27869 14033 27899 14067
rect 28035 14045 28065 14203
rect 28118 14133 28148 14327
rect 28315 14228 28345 14243
rect 28239 14198 28345 14228
rect 28239 14181 28269 14198
rect 28203 14165 28269 14181
rect 28107 14117 28161 14133
rect 28107 14083 28117 14117
rect 28151 14083 28161 14117
rect 28203 14131 28213 14165
rect 28247 14131 28269 14165
rect 28414 14193 28444 14327
rect 28500 14295 28530 14327
rect 28486 14279 28540 14295
rect 28486 14245 28496 14279
rect 28530 14245 28540 14279
rect 28486 14229 28540 14245
rect 28414 14181 28464 14193
rect 28414 14169 28477 14181
rect 28414 14163 28501 14169
rect 28435 14153 28501 14163
rect 28435 14151 28457 14153
rect 28203 14115 28269 14131
rect 28239 14089 28269 14115
rect 28338 14105 28405 14121
rect 28107 14067 28161 14083
rect 28107 14045 28137 14067
rect 28338 14071 28361 14105
rect 28395 14071 28405 14105
rect 28338 14055 28405 14071
rect 28447 14119 28457 14151
rect 28491 14119 28501 14153
rect 28447 14103 28501 14119
rect 28584 14143 28614 14327
rect 28692 14171 28722 14327
rect 28776 14279 28806 14327
rect 28764 14263 28818 14279
rect 28764 14229 28774 14263
rect 28808 14229 28818 14263
rect 28764 14213 28818 14229
rect 28687 14155 28741 14171
rect 28584 14127 28645 14143
rect 28584 14107 28601 14127
rect 28338 14033 28368 14055
rect 28447 14033 28477 14103
rect 28543 14093 28601 14107
rect 28635 14093 28645 14127
rect 28687 14121 28697 14155
rect 28731 14121 28741 14155
rect 28687 14105 28741 14121
rect 28543 14077 28645 14093
rect 28543 14045 28573 14077
rect 28692 14045 28722 14105
rect 28783 14045 28813 14213
rect 29159 14247 29189 14283
rect 29148 14217 29189 14247
rect 28940 14179 28970 14211
rect 29148 14179 29178 14217
rect 30391 14247 30421 14283
rect 30391 14217 30432 14247
rect 29256 14179 29286 14211
rect 29496 14179 29526 14211
rect 29735 14179 29765 14211
rect 28869 14163 29178 14179
rect 28869 14129 28897 14163
rect 28931 14129 29178 14163
rect 28869 14113 29178 14129
rect 29227 14163 29286 14179
rect 29227 14129 29237 14163
rect 29271 14129 29286 14163
rect 29227 14113 29286 14129
rect 29440 14163 29526 14179
rect 29440 14129 29456 14163
rect 29490 14129 29526 14163
rect 29440 14113 29526 14129
rect 29673 14163 29765 14179
rect 29673 14129 29688 14163
rect 29722 14129 29765 14163
rect 29673 14113 29765 14129
rect 28971 14091 29001 14113
rect 29148 14090 29178 14113
rect 29256 14091 29286 14113
rect 29496 14091 29526 14113
rect 29735 14091 29765 14113
rect 29819 14179 29849 14211
rect 30054 14179 30084 14211
rect 30294 14179 30324 14211
rect 30402 14179 30432 14217
rect 30774 14279 30804 14327
rect 30762 14263 30816 14279
rect 30762 14229 30772 14263
rect 30806 14229 30816 14263
rect 30762 14213 30816 14229
rect 30610 14179 30640 14211
rect 29819 14163 29907 14179
rect 29819 14129 29856 14163
rect 29890 14129 29907 14163
rect 29819 14113 29907 14129
rect 30054 14163 30140 14179
rect 30054 14129 30090 14163
rect 30124 14129 30140 14163
rect 30054 14113 30140 14129
rect 30294 14163 30353 14179
rect 30294 14129 30309 14163
rect 30343 14129 30353 14163
rect 30294 14113 30353 14129
rect 30402 14163 30711 14179
rect 30402 14129 30649 14163
rect 30683 14129 30711 14163
rect 30402 14113 30711 14129
rect 29819 14091 29849 14113
rect 30054 14091 30084 14113
rect 30294 14091 30324 14113
rect 29148 14060 29189 14090
rect 29159 14045 29189 14060
rect 30402 14090 30432 14113
rect 30579 14091 30609 14113
rect 30391 14060 30432 14090
rect 30391 14045 30421 14060
rect 30767 14045 30797 14213
rect 30858 14171 30888 14327
rect 30839 14155 30893 14171
rect 30839 14121 30849 14155
rect 30883 14121 30893 14155
rect 30966 14143 30996 14327
rect 31050 14295 31080 14327
rect 31040 14279 31094 14295
rect 31040 14245 31050 14279
rect 31084 14245 31094 14279
rect 31040 14229 31094 14245
rect 31136 14193 31166 14327
rect 32127 14405 32157 14431
rect 32211 14405 32241 14431
rect 31235 14228 31265 14243
rect 31235 14198 31341 14228
rect 31116 14181 31166 14193
rect 31103 14169 31166 14181
rect 30839 14105 30893 14121
rect 30935 14127 30996 14143
rect 30858 14045 30888 14105
rect 30935 14093 30945 14127
rect 30979 14107 30996 14127
rect 31079 14163 31166 14169
rect 31311 14181 31341 14198
rect 31311 14165 31377 14181
rect 31079 14153 31145 14163
rect 31079 14119 31089 14153
rect 31123 14151 31145 14153
rect 31123 14119 31133 14151
rect 31311 14131 31333 14165
rect 31367 14131 31377 14165
rect 31432 14133 31462 14327
rect 31529 14269 31559 14327
rect 31504 14253 31559 14269
rect 31504 14219 31515 14253
rect 31549 14219 31559 14253
rect 31504 14203 31559 14219
rect 30979 14093 31037 14107
rect 31079 14103 31133 14119
rect 30935 14077 31037 14093
rect 31007 14045 31037 14077
rect 31103 14033 31133 14103
rect 31175 14105 31242 14121
rect 31175 14071 31185 14105
rect 31219 14071 31242 14105
rect 31311 14115 31377 14131
rect 31419 14117 31473 14133
rect 31311 14089 31341 14115
rect 31175 14055 31242 14071
rect 31212 14033 31242 14055
rect 31419 14083 31429 14117
rect 31463 14083 31473 14117
rect 31419 14067 31473 14083
rect 31443 14045 31473 14067
rect 31515 14045 31545 14203
rect 31669 14193 31699 14327
rect 31768 14289 31798 14327
rect 31748 14279 31814 14289
rect 31748 14245 31764 14279
rect 31798 14245 31814 14279
rect 31748 14235 31814 14245
rect 31860 14240 31890 14327
rect 31860 14224 31989 14240
rect 31860 14210 31945 14224
rect 31669 14163 31807 14193
rect 31776 14133 31807 14163
rect 31872 14190 31945 14210
rect 31979 14190 31989 14224
rect 31872 14174 31989 14190
rect 32127 14188 32157 14277
rect 32211 14262 32241 14277
rect 32211 14232 32274 14262
rect 32127 14178 32202 14188
rect 31668 14111 31734 14121
rect 31668 14077 31684 14111
rect 31718 14077 31734 14111
rect 31668 14067 31734 14077
rect 31776 14117 31830 14133
rect 31776 14083 31786 14117
rect 31820 14083 31830 14117
rect 31776 14067 31830 14083
rect 31681 14033 31711 14067
rect 31777 14033 31807 14067
rect 31872 14045 31902 14174
rect 32127 14144 32152 14178
rect 32186 14144 32202 14178
rect 32127 14134 32202 14144
rect 32244 14179 32274 14232
rect 32244 14163 32298 14179
rect 32127 14045 32157 14134
rect 32244 14129 32254 14163
rect 32288 14129 32298 14163
rect 32244 14113 32298 14129
rect 32244 14090 32274 14113
rect 32211 14060 32274 14090
rect 32211 14045 32241 14060
rect 27339 13935 27369 13961
rect 27423 13935 27453 13961
rect 27678 13935 27708 13961
rect 27773 13935 27803 13961
rect 27869 13935 27899 13961
rect 28035 13935 28065 13961
rect 28107 13935 28137 13961
rect 28239 13935 28269 13961
rect 28338 13935 28368 13961
rect 28447 13935 28477 13961
rect 28543 13935 28573 13961
rect 28692 13935 28722 13961
rect 28783 13935 28813 13961
rect 28971 13935 29001 13961
rect 29159 13935 29189 13961
rect 29256 13935 29286 13961
rect 29496 13935 29526 13961
rect 29735 13935 29765 13961
rect 29819 13935 29849 13961
rect 30054 13935 30084 13961
rect 30294 13935 30324 13961
rect 30391 13935 30421 13961
rect 30579 13935 30609 13961
rect 30767 13935 30797 13961
rect 30858 13935 30888 13961
rect 31007 13935 31037 13961
rect 31103 13935 31133 13961
rect 31212 13935 31242 13961
rect 31311 13935 31341 13961
rect 31443 13935 31473 13961
rect 31515 13935 31545 13961
rect 31681 13935 31711 13961
rect 31777 13935 31807 13961
rect 31872 13935 31902 13961
rect 32127 13935 32157 13961
rect 32211 13935 32241 13961
rect 24450 12926 24942 12942
rect 24450 12909 24466 12926
rect 24296 12892 24466 12909
rect 24926 12909 24942 12926
rect 25308 12926 25800 12942
rect 25308 12909 25324 12926
rect 24926 12892 25096 12909
rect 24296 12854 25096 12892
rect 25154 12892 25324 12909
rect 25784 12909 25800 12926
rect 26166 12926 26658 12942
rect 26166 12909 26182 12926
rect 25784 12892 25954 12909
rect 25154 12854 25954 12892
rect 26012 12892 26182 12909
rect 26642 12909 26658 12926
rect 27024 12926 27516 12942
rect 27024 12909 27040 12926
rect 26642 12892 26812 12909
rect 26012 12854 26812 12892
rect 26870 12892 27040 12909
rect 27500 12909 27516 12926
rect 27882 12926 28374 12942
rect 27882 12909 27898 12926
rect 27500 12892 27670 12909
rect 26870 12854 27670 12892
rect 27728 12892 27898 12909
rect 28358 12909 28374 12926
rect 28740 12926 29232 12942
rect 28740 12909 28756 12926
rect 28358 12892 28528 12909
rect 27728 12854 28528 12892
rect 28586 12892 28756 12909
rect 29216 12909 29232 12926
rect 29598 12926 30090 12942
rect 29598 12909 29614 12926
rect 29216 12892 29386 12909
rect 28586 12854 29386 12892
rect 29444 12892 29614 12909
rect 30074 12909 30090 12926
rect 30456 12926 30948 12942
rect 30456 12909 30472 12926
rect 30074 12892 30244 12909
rect 29444 12854 30244 12892
rect 30302 12892 30472 12909
rect 30932 12909 30948 12926
rect 31314 12926 31806 12942
rect 31314 12909 31330 12926
rect 30932 12892 31102 12909
rect 30302 12854 31102 12892
rect 31160 12892 31330 12909
rect 31790 12909 31806 12926
rect 31790 12892 31960 12909
rect 31160 12854 31960 12892
rect 24296 12616 25096 12654
rect 24296 12599 24466 12616
rect 24450 12582 24466 12599
rect 24926 12599 25096 12616
rect 25154 12616 25954 12654
rect 25154 12599 25324 12616
rect 24926 12582 24942 12599
rect 24450 12566 24942 12582
rect 25308 12582 25324 12599
rect 25784 12599 25954 12616
rect 26012 12616 26812 12654
rect 26012 12599 26182 12616
rect 25784 12582 25800 12599
rect 25308 12566 25800 12582
rect 26166 12582 26182 12599
rect 26642 12599 26812 12616
rect 26870 12616 27670 12654
rect 26870 12599 27040 12616
rect 26642 12582 26658 12599
rect 26166 12566 26658 12582
rect 27024 12582 27040 12599
rect 27500 12599 27670 12616
rect 27728 12616 28528 12654
rect 27728 12599 27898 12616
rect 27500 12582 27516 12599
rect 27024 12566 27516 12582
rect 27882 12582 27898 12599
rect 28358 12599 28528 12616
rect 28586 12616 29386 12654
rect 28586 12599 28756 12616
rect 28358 12582 28374 12599
rect 27882 12566 28374 12582
rect 28740 12582 28756 12599
rect 29216 12599 29386 12616
rect 29444 12616 30244 12654
rect 29444 12599 29614 12616
rect 29216 12582 29232 12599
rect 28740 12566 29232 12582
rect 29598 12582 29614 12599
rect 30074 12599 30244 12616
rect 30302 12616 31102 12654
rect 30302 12599 30472 12616
rect 30074 12582 30090 12599
rect 29598 12566 30090 12582
rect 30456 12582 30472 12599
rect 30932 12599 31102 12616
rect 31160 12616 31960 12654
rect 31160 12599 31330 12616
rect 30932 12582 30948 12599
rect 30456 12566 30948 12582
rect 31314 12582 31330 12599
rect 31790 12599 31960 12616
rect 31790 12582 31806 12599
rect 31314 12566 31806 12582
rect 24450 12344 24942 12360
rect 24450 12327 24466 12344
rect 24296 12310 24466 12327
rect 24926 12327 24942 12344
rect 25308 12344 25800 12360
rect 25308 12327 25324 12344
rect 24926 12310 25096 12327
rect 24296 12272 25096 12310
rect 25154 12310 25324 12327
rect 25784 12327 25800 12344
rect 26166 12344 26658 12360
rect 26166 12327 26182 12344
rect 25784 12310 25954 12327
rect 25154 12272 25954 12310
rect 26012 12310 26182 12327
rect 26642 12327 26658 12344
rect 27024 12344 27516 12360
rect 27024 12327 27040 12344
rect 26642 12310 26812 12327
rect 26012 12272 26812 12310
rect 26870 12310 27040 12327
rect 27500 12327 27516 12344
rect 27882 12344 28374 12360
rect 27882 12327 27898 12344
rect 27500 12310 27670 12327
rect 26870 12272 27670 12310
rect 27728 12310 27898 12327
rect 28358 12327 28374 12344
rect 28740 12344 29232 12360
rect 28740 12327 28756 12344
rect 28358 12310 28528 12327
rect 27728 12272 28528 12310
rect 28586 12310 28756 12327
rect 29216 12327 29232 12344
rect 29598 12344 30090 12360
rect 29598 12327 29614 12344
rect 29216 12310 29386 12327
rect 28586 12272 29386 12310
rect 29444 12310 29614 12327
rect 30074 12327 30090 12344
rect 30456 12344 30948 12360
rect 30456 12327 30472 12344
rect 30074 12310 30244 12327
rect 29444 12272 30244 12310
rect 30302 12310 30472 12327
rect 30932 12327 30948 12344
rect 31314 12344 31806 12360
rect 31314 12327 31330 12344
rect 30932 12310 31102 12327
rect 30302 12272 31102 12310
rect 31160 12310 31330 12327
rect 31790 12327 31806 12344
rect 31790 12310 31960 12327
rect 31160 12272 31960 12310
rect 24296 12034 25096 12072
rect 24296 12017 24466 12034
rect 24450 12000 24466 12017
rect 24926 12017 25096 12034
rect 25154 12034 25954 12072
rect 25154 12017 25324 12034
rect 24926 12000 24942 12017
rect 24450 11984 24942 12000
rect 25308 12000 25324 12017
rect 25784 12017 25954 12034
rect 26012 12034 26812 12072
rect 26012 12017 26182 12034
rect 25784 12000 25800 12017
rect 25308 11984 25800 12000
rect 26166 12000 26182 12017
rect 26642 12017 26812 12034
rect 26870 12034 27670 12072
rect 26870 12017 27040 12034
rect 26642 12000 26658 12017
rect 26166 11984 26658 12000
rect 27024 12000 27040 12017
rect 27500 12017 27670 12034
rect 27728 12034 28528 12072
rect 27728 12017 27898 12034
rect 27500 12000 27516 12017
rect 27024 11984 27516 12000
rect 27882 12000 27898 12017
rect 28358 12017 28528 12034
rect 28586 12034 29386 12072
rect 28586 12017 28756 12034
rect 28358 12000 28374 12017
rect 27882 11984 28374 12000
rect 28740 12000 28756 12017
rect 29216 12017 29386 12034
rect 29444 12034 30244 12072
rect 29444 12017 29614 12034
rect 29216 12000 29232 12017
rect 28740 11984 29232 12000
rect 29598 12000 29614 12017
rect 30074 12017 30244 12034
rect 30302 12034 31102 12072
rect 30302 12017 30472 12034
rect 30074 12000 30090 12017
rect 29598 11984 30090 12000
rect 30456 12000 30472 12017
rect 30932 12017 31102 12034
rect 31160 12034 31960 12072
rect 31160 12017 31330 12034
rect 30932 12000 30948 12017
rect 30456 11984 30948 12000
rect 31314 12000 31330 12017
rect 31790 12017 31960 12034
rect 31790 12000 31806 12017
rect 31314 11984 31806 12000
rect 15288 9740 15540 9756
rect 15288 9723 15304 9740
rect 15214 9706 15304 9723
rect 15524 9723 15540 9740
rect 15746 9740 15998 9756
rect 15746 9723 15762 9740
rect 15524 9706 15614 9723
rect 15214 9668 15614 9706
rect 15672 9706 15762 9723
rect 15982 9723 15998 9740
rect 16204 9740 16456 9756
rect 16204 9723 16220 9740
rect 15982 9706 16072 9723
rect 15672 9668 16072 9706
rect 16130 9706 16220 9723
rect 16440 9723 16456 9740
rect 16662 9740 16914 9756
rect 16662 9723 16678 9740
rect 16440 9706 16530 9723
rect 16130 9668 16530 9706
rect 16588 9706 16678 9723
rect 16898 9723 16914 9740
rect 17120 9740 17372 9756
rect 17120 9723 17136 9740
rect 16898 9706 16988 9723
rect 16588 9668 16988 9706
rect 17046 9706 17136 9723
rect 17356 9723 17372 9740
rect 17578 9740 17830 9756
rect 17578 9723 17594 9740
rect 17356 9706 17446 9723
rect 17046 9668 17446 9706
rect 17504 9706 17594 9723
rect 17814 9723 17830 9740
rect 18036 9740 18288 9756
rect 18036 9723 18052 9740
rect 17814 9706 17904 9723
rect 17504 9668 17904 9706
rect 17962 9706 18052 9723
rect 18272 9723 18288 9740
rect 18494 9740 18746 9756
rect 18494 9723 18510 9740
rect 18272 9706 18362 9723
rect 17962 9668 18362 9706
rect 18420 9706 18510 9723
rect 18730 9723 18746 9740
rect 18952 9740 19204 9756
rect 18952 9723 18968 9740
rect 18730 9706 18820 9723
rect 18420 9668 18820 9706
rect 18878 9706 18968 9723
rect 19188 9723 19204 9740
rect 19410 9740 19662 9756
rect 19410 9723 19426 9740
rect 19188 9706 19278 9723
rect 18878 9668 19278 9706
rect 19336 9706 19426 9723
rect 19646 9723 19662 9740
rect 19646 9706 19736 9723
rect 19336 9668 19736 9706
rect 15214 9430 15614 9468
rect 15214 9413 15304 9430
rect 15288 9396 15304 9413
rect 15524 9413 15614 9430
rect 15672 9430 16072 9468
rect 15672 9413 15762 9430
rect 15524 9396 15540 9413
rect 15288 9380 15540 9396
rect 15746 9396 15762 9413
rect 15982 9413 16072 9430
rect 16130 9430 16530 9468
rect 16130 9413 16220 9430
rect 15982 9396 15998 9413
rect 15746 9380 15998 9396
rect 16204 9396 16220 9413
rect 16440 9413 16530 9430
rect 16588 9430 16988 9468
rect 16588 9413 16678 9430
rect 16440 9396 16456 9413
rect 16204 9380 16456 9396
rect 16662 9396 16678 9413
rect 16898 9413 16988 9430
rect 17046 9430 17446 9468
rect 17046 9413 17136 9430
rect 16898 9396 16914 9413
rect 16662 9380 16914 9396
rect 17120 9396 17136 9413
rect 17356 9413 17446 9430
rect 17504 9430 17904 9468
rect 17504 9413 17594 9430
rect 17356 9396 17372 9413
rect 17120 9380 17372 9396
rect 17578 9396 17594 9413
rect 17814 9413 17904 9430
rect 17962 9430 18362 9468
rect 17962 9413 18052 9430
rect 17814 9396 17830 9413
rect 17578 9380 17830 9396
rect 18036 9396 18052 9413
rect 18272 9413 18362 9430
rect 18420 9430 18820 9468
rect 18420 9413 18510 9430
rect 18272 9396 18288 9413
rect 18036 9380 18288 9396
rect 18494 9396 18510 9413
rect 18730 9413 18820 9430
rect 18878 9430 19278 9468
rect 18878 9413 18968 9430
rect 18730 9396 18746 9413
rect 18494 9380 18746 9396
rect 18952 9396 18968 9413
rect 19188 9413 19278 9430
rect 19336 9430 19736 9468
rect 19336 9413 19426 9430
rect 19188 9396 19204 9413
rect 18952 9380 19204 9396
rect 19410 9396 19426 9413
rect 19646 9413 19736 9430
rect 19646 9396 19662 9413
rect 19410 9380 19662 9396
rect 24050 9740 24302 9756
rect 24050 9723 24066 9740
rect 23976 9706 24066 9723
rect 24286 9723 24302 9740
rect 24508 9740 24760 9756
rect 24508 9723 24524 9740
rect 24286 9706 24376 9723
rect 23976 9668 24376 9706
rect 24434 9706 24524 9723
rect 24744 9723 24760 9740
rect 24966 9740 25218 9756
rect 24966 9723 24982 9740
rect 24744 9706 24834 9723
rect 24434 9668 24834 9706
rect 24892 9706 24982 9723
rect 25202 9723 25218 9740
rect 25424 9740 25676 9756
rect 25424 9723 25440 9740
rect 25202 9706 25292 9723
rect 24892 9668 25292 9706
rect 25350 9706 25440 9723
rect 25660 9723 25676 9740
rect 25882 9740 26134 9756
rect 25882 9723 25898 9740
rect 25660 9706 25750 9723
rect 25350 9668 25750 9706
rect 25808 9706 25898 9723
rect 26118 9723 26134 9740
rect 26340 9740 26592 9756
rect 26340 9723 26356 9740
rect 26118 9706 26208 9723
rect 25808 9668 26208 9706
rect 26266 9706 26356 9723
rect 26576 9723 26592 9740
rect 26798 9740 27050 9756
rect 26798 9723 26814 9740
rect 26576 9706 26666 9723
rect 26266 9668 26666 9706
rect 26724 9706 26814 9723
rect 27034 9723 27050 9740
rect 27256 9740 27508 9756
rect 27256 9723 27272 9740
rect 27034 9706 27124 9723
rect 26724 9668 27124 9706
rect 27182 9706 27272 9723
rect 27492 9723 27508 9740
rect 27714 9740 27966 9756
rect 27714 9723 27730 9740
rect 27492 9706 27582 9723
rect 27182 9668 27582 9706
rect 27640 9706 27730 9723
rect 27950 9723 27966 9740
rect 28172 9740 28424 9756
rect 28172 9723 28188 9740
rect 27950 9706 28040 9723
rect 27640 9668 28040 9706
rect 28098 9706 28188 9723
rect 28408 9723 28424 9740
rect 28408 9706 28498 9723
rect 28098 9668 28498 9706
rect 23976 9430 24376 9468
rect 23976 9413 24066 9430
rect 24050 9396 24066 9413
rect 24286 9413 24376 9430
rect 24434 9430 24834 9468
rect 24434 9413 24524 9430
rect 24286 9396 24302 9413
rect 24050 9380 24302 9396
rect 24508 9396 24524 9413
rect 24744 9413 24834 9430
rect 24892 9430 25292 9468
rect 24892 9413 24982 9430
rect 24744 9396 24760 9413
rect 24508 9380 24760 9396
rect 24966 9396 24982 9413
rect 25202 9413 25292 9430
rect 25350 9430 25750 9468
rect 25350 9413 25440 9430
rect 25202 9396 25218 9413
rect 24966 9380 25218 9396
rect 25424 9396 25440 9413
rect 25660 9413 25750 9430
rect 25808 9430 26208 9468
rect 25808 9413 25898 9430
rect 25660 9396 25676 9413
rect 25424 9380 25676 9396
rect 25882 9396 25898 9413
rect 26118 9413 26208 9430
rect 26266 9430 26666 9468
rect 26266 9413 26356 9430
rect 26118 9396 26134 9413
rect 25882 9380 26134 9396
rect 26340 9396 26356 9413
rect 26576 9413 26666 9430
rect 26724 9430 27124 9468
rect 26724 9413 26814 9430
rect 26576 9396 26592 9413
rect 26340 9380 26592 9396
rect 26798 9396 26814 9413
rect 27034 9413 27124 9430
rect 27182 9430 27582 9468
rect 27182 9413 27272 9430
rect 27034 9396 27050 9413
rect 26798 9380 27050 9396
rect 27256 9396 27272 9413
rect 27492 9413 27582 9430
rect 27640 9430 28040 9468
rect 27640 9413 27730 9430
rect 27492 9396 27508 9413
rect 27256 9380 27508 9396
rect 27714 9396 27730 9413
rect 27950 9413 28040 9430
rect 28098 9430 28498 9468
rect 28098 9413 28188 9430
rect 27950 9396 27966 9413
rect 27714 9380 27966 9396
rect 28172 9396 28188 9413
rect 28408 9413 28498 9430
rect 28408 9396 28424 9413
rect 28172 9380 28424 9396
rect 30631 8907 30661 8933
rect 30715 8907 30745 8933
rect 30903 8913 30933 8939
rect 30988 8913 31018 8939
rect 31083 8913 31113 8939
rect 31186 8913 31216 8939
rect 31318 8913 31348 8939
rect 31413 8913 31443 8939
rect 31497 8913 31527 8939
rect 31611 8913 31641 8939
rect 31822 8913 31852 8939
rect 31906 8913 31936 8939
rect 32094 8913 32124 8939
rect 32191 8913 32221 8939
rect 32420 8913 32450 8939
rect 32665 8913 32695 8939
rect 32749 8913 32779 8939
rect 32833 8913 32863 8939
rect 32917 8913 32947 8939
rect 29196 8867 29226 8893
rect 29441 8867 29471 8893
rect 29525 8867 29555 8893
rect 29609 8867 29639 8893
rect 29693 8867 29723 8893
rect 30631 8764 30661 8779
rect 29196 8715 29226 8737
rect 29441 8715 29471 8737
rect 29525 8715 29555 8737
rect 29609 8715 29639 8737
rect 29693 8715 29723 8737
rect 30598 8734 30661 8764
rect 29140 8699 29226 8715
rect 29140 8665 29156 8699
rect 29190 8665 29226 8699
rect 29140 8649 29226 8665
rect 29373 8699 29723 8715
rect 29373 8665 29389 8699
rect 29423 8665 29481 8699
rect 29515 8665 29565 8699
rect 29599 8665 29649 8699
rect 29683 8665 29723 8699
rect 30598 8681 30628 8734
rect 30715 8690 30745 8779
rect 30903 8749 30933 8829
rect 29373 8649 29723 8665
rect 13456 7898 13708 7914
rect 13456 7881 13472 7898
rect 13382 7864 13472 7881
rect 13692 7881 13708 7898
rect 13914 7898 14166 7914
rect 13914 7881 13930 7898
rect 13692 7864 13782 7881
rect 13382 7817 13782 7864
rect 13840 7864 13930 7881
rect 14150 7881 14166 7898
rect 14372 7898 14624 7914
rect 14372 7881 14388 7898
rect 14150 7864 14240 7881
rect 13840 7817 14240 7864
rect 14298 7864 14388 7881
rect 14608 7881 14624 7898
rect 14830 7898 15082 7914
rect 14830 7881 14846 7898
rect 14608 7864 14698 7881
rect 14298 7817 14698 7864
rect 14756 7864 14846 7881
rect 15066 7881 15082 7898
rect 15288 7898 15540 7914
rect 15288 7881 15304 7898
rect 15066 7864 15156 7881
rect 14756 7817 15156 7864
rect 15214 7864 15304 7881
rect 15524 7881 15540 7898
rect 15746 7898 15998 7914
rect 15746 7881 15762 7898
rect 15524 7864 15614 7881
rect 15214 7817 15614 7864
rect 15672 7864 15762 7881
rect 15982 7881 15998 7898
rect 16204 7898 16456 7914
rect 16204 7881 16220 7898
rect 15982 7864 16072 7881
rect 15672 7817 16072 7864
rect 16130 7864 16220 7881
rect 16440 7881 16456 7898
rect 16662 7898 16914 7914
rect 16662 7881 16678 7898
rect 16440 7864 16530 7881
rect 16130 7817 16530 7864
rect 16588 7864 16678 7881
rect 16898 7881 16914 7898
rect 17120 7898 17372 7914
rect 17120 7881 17136 7898
rect 16898 7864 16988 7881
rect 16588 7817 16988 7864
rect 17046 7864 17136 7881
rect 17356 7881 17372 7898
rect 17578 7898 17830 7914
rect 17578 7881 17594 7898
rect 17356 7864 17446 7881
rect 17046 7817 17446 7864
rect 17504 7864 17594 7881
rect 17814 7881 17830 7898
rect 18036 7898 18288 7914
rect 18036 7881 18052 7898
rect 17814 7864 17904 7881
rect 17504 7817 17904 7864
rect 17962 7864 18052 7881
rect 18272 7881 18288 7898
rect 18494 7898 18746 7914
rect 18494 7881 18510 7898
rect 18272 7864 18362 7881
rect 17962 7817 18362 7864
rect 18420 7864 18510 7881
rect 18730 7881 18746 7898
rect 18952 7898 19204 7914
rect 18952 7881 18968 7898
rect 18730 7864 18820 7881
rect 18420 7817 18820 7864
rect 18878 7864 18968 7881
rect 19188 7881 19204 7898
rect 19410 7898 19662 7914
rect 19410 7881 19426 7898
rect 19188 7864 19278 7881
rect 18878 7817 19278 7864
rect 19336 7864 19426 7881
rect 19646 7881 19662 7898
rect 19868 7898 20120 7914
rect 19868 7881 19884 7898
rect 19646 7864 19736 7881
rect 19336 7817 19736 7864
rect 19794 7864 19884 7881
rect 20104 7881 20120 7898
rect 20326 7898 20578 7914
rect 20326 7881 20342 7898
rect 20104 7864 20194 7881
rect 19794 7817 20194 7864
rect 20252 7864 20342 7881
rect 20562 7881 20578 7898
rect 20784 7898 21036 7914
rect 20784 7881 20800 7898
rect 20562 7864 20652 7881
rect 20252 7817 20652 7864
rect 20710 7864 20800 7881
rect 21020 7881 21036 7898
rect 21242 7898 21494 7914
rect 21242 7881 21258 7898
rect 21020 7864 21110 7881
rect 20710 7817 21110 7864
rect 21168 7864 21258 7881
rect 21478 7881 21494 7898
rect 21478 7864 21568 7881
rect 21168 7817 21568 7864
rect 13382 6170 13782 6217
rect 13382 6153 13472 6170
rect 13456 6136 13472 6153
rect 13692 6153 13782 6170
rect 13840 6170 14240 6217
rect 13840 6153 13930 6170
rect 13692 6136 13708 6153
rect 13456 6120 13708 6136
rect 13914 6136 13930 6153
rect 14150 6153 14240 6170
rect 14298 6170 14698 6217
rect 14298 6153 14388 6170
rect 14150 6136 14166 6153
rect 13914 6120 14166 6136
rect 14372 6136 14388 6153
rect 14608 6153 14698 6170
rect 14756 6170 15156 6217
rect 14756 6153 14846 6170
rect 14608 6136 14624 6153
rect 14372 6120 14624 6136
rect 14830 6136 14846 6153
rect 15066 6153 15156 6170
rect 15214 6170 15614 6217
rect 15214 6153 15304 6170
rect 15066 6136 15082 6153
rect 14830 6120 15082 6136
rect 15288 6136 15304 6153
rect 15524 6153 15614 6170
rect 15672 6170 16072 6217
rect 15672 6153 15762 6170
rect 15524 6136 15540 6153
rect 15288 6120 15540 6136
rect 15746 6136 15762 6153
rect 15982 6153 16072 6170
rect 16130 6170 16530 6217
rect 16130 6153 16220 6170
rect 15982 6136 15998 6153
rect 15746 6120 15998 6136
rect 16204 6136 16220 6153
rect 16440 6153 16530 6170
rect 16588 6170 16988 6217
rect 16588 6153 16678 6170
rect 16440 6136 16456 6153
rect 16204 6120 16456 6136
rect 16662 6136 16678 6153
rect 16898 6153 16988 6170
rect 17046 6170 17446 6217
rect 17046 6153 17136 6170
rect 16898 6136 16914 6153
rect 16662 6120 16914 6136
rect 17120 6136 17136 6153
rect 17356 6153 17446 6170
rect 17504 6170 17904 6217
rect 17504 6153 17594 6170
rect 17356 6136 17372 6153
rect 17120 6120 17372 6136
rect 17578 6136 17594 6153
rect 17814 6153 17904 6170
rect 17962 6170 18362 6217
rect 17962 6153 18052 6170
rect 17814 6136 17830 6153
rect 17578 6120 17830 6136
rect 18036 6136 18052 6153
rect 18272 6153 18362 6170
rect 18420 6170 18820 6217
rect 18420 6153 18510 6170
rect 18272 6136 18288 6153
rect 18036 6120 18288 6136
rect 18494 6136 18510 6153
rect 18730 6153 18820 6170
rect 18878 6170 19278 6217
rect 18878 6153 18968 6170
rect 18730 6136 18746 6153
rect 18494 6120 18746 6136
rect 18952 6136 18968 6153
rect 19188 6153 19278 6170
rect 19336 6170 19736 6217
rect 19336 6153 19426 6170
rect 19188 6136 19204 6153
rect 18952 6120 19204 6136
rect 19410 6136 19426 6153
rect 19646 6153 19736 6170
rect 19794 6170 20194 6217
rect 19794 6153 19884 6170
rect 19646 6136 19662 6153
rect 19410 6120 19662 6136
rect 19868 6136 19884 6153
rect 20104 6153 20194 6170
rect 20252 6170 20652 6217
rect 20252 6153 20342 6170
rect 20104 6136 20120 6153
rect 19868 6120 20120 6136
rect 20326 6136 20342 6153
rect 20562 6153 20652 6170
rect 20710 6170 21110 6217
rect 20710 6153 20800 6170
rect 20562 6136 20578 6153
rect 20326 6120 20578 6136
rect 20784 6136 20800 6153
rect 21020 6153 21110 6170
rect 21168 6170 21568 6217
rect 21168 6153 21258 6170
rect 21020 6136 21036 6153
rect 20784 6120 21036 6136
rect 21242 6136 21258 6153
rect 21478 6153 21568 6170
rect 21478 6136 21494 6153
rect 21242 6120 21494 6136
rect 29196 8617 29226 8649
rect 29441 8617 29471 8649
rect 29525 8617 29555 8649
rect 29609 8617 29639 8649
rect 29693 8617 29723 8649
rect 30574 8665 30628 8681
rect 30574 8631 30584 8665
rect 30618 8631 30628 8665
rect 30670 8680 30745 8690
rect 30838 8733 30933 8749
rect 30838 8699 30848 8733
rect 30882 8699 30933 8733
rect 30988 8713 31018 8829
rect 31083 8797 31113 8829
rect 31083 8781 31144 8797
rect 31083 8747 31100 8781
rect 31134 8747 31144 8781
rect 31083 8731 31144 8747
rect 30838 8683 30933 8699
rect 30670 8646 30686 8680
rect 30720 8646 30745 8680
rect 30670 8636 30745 8646
rect 24051 8318 24303 8334
rect 24051 8301 24067 8318
rect 23977 8284 24067 8301
rect 24287 8301 24303 8318
rect 24509 8318 24761 8334
rect 24509 8301 24525 8318
rect 24287 8284 24377 8301
rect 23977 8237 24377 8284
rect 24435 8284 24525 8301
rect 24745 8301 24761 8318
rect 24967 8318 25219 8334
rect 24967 8301 24983 8318
rect 24745 8284 24835 8301
rect 24435 8237 24835 8284
rect 24893 8284 24983 8301
rect 25203 8301 25219 8318
rect 25425 8318 25677 8334
rect 25425 8301 25441 8318
rect 25203 8284 25293 8301
rect 24893 8237 25293 8284
rect 25351 8284 25441 8301
rect 25661 8301 25677 8318
rect 25883 8318 26135 8334
rect 25883 8301 25899 8318
rect 25661 8284 25751 8301
rect 25351 8237 25751 8284
rect 25809 8284 25899 8301
rect 26119 8301 26135 8318
rect 26341 8318 26593 8334
rect 26341 8301 26357 8318
rect 26119 8284 26209 8301
rect 25809 8237 26209 8284
rect 26267 8284 26357 8301
rect 26577 8301 26593 8318
rect 26799 8318 27051 8334
rect 26799 8301 26815 8318
rect 26577 8284 26667 8301
rect 26267 8237 26667 8284
rect 26725 8284 26815 8301
rect 27035 8301 27051 8318
rect 27257 8318 27509 8334
rect 27257 8301 27273 8318
rect 27035 8284 27125 8301
rect 26725 8237 27125 8284
rect 27183 8284 27273 8301
rect 27493 8301 27509 8318
rect 27715 8318 27967 8334
rect 27715 8301 27731 8318
rect 27493 8284 27583 8301
rect 27183 8237 27583 8284
rect 27641 8284 27731 8301
rect 27951 8301 27967 8318
rect 28173 8318 28425 8334
rect 28173 8301 28189 8318
rect 27951 8284 28041 8301
rect 27641 8237 28041 8284
rect 28099 8284 28189 8301
rect 28409 8301 28425 8318
rect 28409 8284 28499 8301
rect 28099 8237 28499 8284
rect 23977 6990 24377 7037
rect 23977 6973 24067 6990
rect 24051 6956 24067 6973
rect 24287 6973 24377 6990
rect 24435 6990 24835 7037
rect 24435 6973 24525 6990
rect 24287 6956 24303 6973
rect 24051 6940 24303 6956
rect 24509 6956 24525 6973
rect 24745 6973 24835 6990
rect 24893 6990 25293 7037
rect 24893 6973 24983 6990
rect 24745 6956 24761 6973
rect 24509 6940 24761 6956
rect 24967 6956 24983 6973
rect 25203 6973 25293 6990
rect 25351 6990 25751 7037
rect 25351 6973 25441 6990
rect 25203 6956 25219 6973
rect 24967 6940 25219 6956
rect 25425 6956 25441 6973
rect 25661 6973 25751 6990
rect 25809 6990 26209 7037
rect 25809 6973 25899 6990
rect 25661 6956 25677 6973
rect 25425 6940 25677 6956
rect 25883 6956 25899 6973
rect 26119 6973 26209 6990
rect 26267 6990 26667 7037
rect 26267 6973 26357 6990
rect 26119 6956 26135 6973
rect 25883 6940 26135 6956
rect 26341 6956 26357 6973
rect 26577 6973 26667 6990
rect 26725 6990 27125 7037
rect 26725 6973 26815 6990
rect 26577 6956 26593 6973
rect 26341 6940 26593 6956
rect 26799 6956 26815 6973
rect 27035 6973 27125 6990
rect 27183 6990 27583 7037
rect 27183 6973 27273 6990
rect 27035 6956 27051 6973
rect 26799 6940 27051 6956
rect 27257 6956 27273 6973
rect 27493 6973 27583 6990
rect 27641 6990 28041 7037
rect 27641 6973 27731 6990
rect 27493 6956 27509 6973
rect 27257 6940 27509 6956
rect 27715 6956 27731 6973
rect 27951 6973 28041 6990
rect 28099 6990 28499 7037
rect 28099 6973 28189 6990
rect 27951 6956 27967 6973
rect 27715 6940 27967 6956
rect 28173 6956 28189 6973
rect 28409 6973 28499 6990
rect 28409 6956 28425 6973
rect 28173 6940 28425 6956
rect 30574 8615 30628 8631
rect 30598 8592 30628 8615
rect 30598 8562 30661 8592
rect 30631 8547 30661 8562
rect 30715 8547 30745 8636
rect 30903 8547 30933 8683
rect 30975 8703 31041 8713
rect 30975 8669 30991 8703
rect 31025 8689 31041 8703
rect 31025 8669 31144 8689
rect 30975 8659 31144 8669
rect 30995 8607 31061 8617
rect 30995 8573 31011 8607
rect 31045 8573 31061 8607
rect 30995 8563 31061 8573
rect 31015 8535 31045 8563
rect 31114 8535 31144 8659
rect 31186 8629 31216 8829
rect 31318 8725 31348 8763
rect 31413 8731 31443 8829
rect 31497 8791 31527 8829
rect 31611 8797 31641 8829
rect 31496 8781 31562 8791
rect 31496 8747 31512 8781
rect 31546 8747 31562 8781
rect 31496 8737 31562 8747
rect 31611 8781 31692 8797
rect 31611 8747 31648 8781
rect 31682 8747 31692 8781
rect 31611 8731 31692 8747
rect 31258 8715 31348 8725
rect 31258 8681 31274 8715
rect 31308 8681 31348 8715
rect 31258 8671 31348 8681
rect 31318 8636 31348 8671
rect 31400 8715 31454 8731
rect 31400 8681 31410 8715
rect 31444 8695 31454 8715
rect 31444 8681 31569 8695
rect 31400 8665 31569 8681
rect 31186 8619 31260 8629
rect 31186 8585 31210 8619
rect 31244 8585 31260 8619
rect 31318 8606 31362 8636
rect 31332 8591 31362 8606
rect 31433 8607 31497 8623
rect 31186 8575 31260 8585
rect 31213 8547 31243 8575
rect 31433 8573 31453 8607
rect 31487 8573 31497 8607
rect 31433 8557 31497 8573
rect 31433 8535 31463 8557
rect 31539 8535 31569 8665
rect 31634 8547 31664 8731
rect 32094 8749 32124 8785
rect 32085 8719 32124 8749
rect 31822 8681 31852 8713
rect 31906 8681 31936 8713
rect 32085 8681 32115 8719
rect 32191 8681 32221 8713
rect 32420 8681 32450 8713
rect 32665 8681 32695 8713
rect 32749 8681 32779 8713
rect 32833 8681 32863 8713
rect 32917 8681 32947 8713
rect 31712 8665 31854 8681
rect 31712 8631 31722 8665
rect 31756 8631 31854 8665
rect 31712 8615 31854 8631
rect 31896 8665 32115 8681
rect 31896 8631 31906 8665
rect 31940 8631 32115 8665
rect 31896 8615 32115 8631
rect 32157 8665 32221 8681
rect 32157 8631 32167 8665
rect 32201 8631 32221 8665
rect 32157 8615 32221 8631
rect 32364 8665 32450 8681
rect 32364 8631 32380 8665
rect 32414 8631 32450 8665
rect 32364 8615 32450 8631
rect 32597 8665 32947 8681
rect 32597 8631 32613 8665
rect 32647 8631 32705 8665
rect 32739 8631 32789 8665
rect 32823 8631 32873 8665
rect 32907 8631 32947 8665
rect 32597 8615 32947 8631
rect 31824 8593 31854 8615
rect 31908 8593 31938 8615
rect 32085 8586 32115 8615
rect 32191 8593 32221 8615
rect 32420 8593 32450 8615
rect 32665 8593 32695 8615
rect 32749 8593 32779 8615
rect 32833 8593 32863 8615
rect 32917 8593 32947 8615
rect 32085 8562 32126 8586
rect 32096 8547 32126 8562
rect 30631 8437 30661 8463
rect 30715 8437 30745 8463
rect 30903 8437 30933 8463
rect 31015 8437 31045 8463
rect 31114 8437 31144 8463
rect 31213 8437 31243 8463
rect 31332 8437 31362 8463
rect 31433 8437 31463 8463
rect 31539 8437 31569 8463
rect 31634 8437 31664 8463
rect 31824 8437 31854 8463
rect 31908 8437 31938 8463
rect 32096 8437 32126 8463
rect 32191 8437 32221 8463
rect 32420 8437 32450 8463
rect 32665 8437 32695 8463
rect 32749 8437 32779 8463
rect 32833 8437 32863 8463
rect 32917 8437 32947 8463
rect 29196 8391 29226 8417
rect 29441 8391 29471 8417
rect 29525 8391 29555 8417
rect 29609 8391 29639 8417
rect 29693 8391 29723 8417
rect 30631 8369 30661 8395
rect 30715 8369 30745 8395
rect 30903 8369 30933 8395
rect 31015 8369 31045 8395
rect 31114 8369 31144 8395
rect 31213 8369 31243 8395
rect 31332 8369 31362 8395
rect 31433 8369 31463 8395
rect 31539 8369 31569 8395
rect 31634 8369 31664 8395
rect 31824 8369 31854 8395
rect 31908 8369 31938 8395
rect 32096 8369 32126 8395
rect 32191 8369 32221 8395
rect 32420 8369 32450 8395
rect 32665 8369 32695 8395
rect 32749 8369 32779 8395
rect 32833 8369 32863 8395
rect 32917 8369 32947 8395
rect 33329 8369 33359 8395
rect 33413 8369 33443 8395
rect 33601 8369 33631 8395
rect 33713 8369 33743 8395
rect 33812 8369 33842 8395
rect 33911 8369 33941 8395
rect 34030 8369 34060 8395
rect 34131 8369 34161 8395
rect 34237 8369 34267 8395
rect 34332 8369 34362 8395
rect 34522 8369 34552 8395
rect 34606 8369 34636 8395
rect 34794 8369 34824 8395
rect 34889 8369 34919 8395
rect 35118 8369 35148 8395
rect 35363 8369 35393 8395
rect 35447 8369 35477 8395
rect 35531 8369 35561 8395
rect 35615 8369 35645 8395
rect 30631 8270 30661 8285
rect 30598 8240 30661 8270
rect 30598 8217 30628 8240
rect 30574 8201 30628 8217
rect 30574 8167 30584 8201
rect 30618 8167 30628 8201
rect 30715 8196 30745 8285
rect 30574 8151 30628 8167
rect 30598 8098 30628 8151
rect 30670 8186 30745 8196
rect 30670 8152 30686 8186
rect 30720 8152 30745 8186
rect 30670 8142 30745 8152
rect 30903 8149 30933 8285
rect 31015 8269 31045 8297
rect 30995 8259 31061 8269
rect 30995 8225 31011 8259
rect 31045 8225 31061 8259
rect 30995 8215 31061 8225
rect 31114 8173 31144 8297
rect 31213 8257 31243 8285
rect 30598 8068 30661 8098
rect 30631 8053 30661 8068
rect 30715 8053 30745 8142
rect 30838 8133 30933 8149
rect 30838 8099 30848 8133
rect 30882 8099 30933 8133
rect 30975 8163 31144 8173
rect 30975 8129 30991 8163
rect 31025 8143 31144 8163
rect 31186 8247 31260 8257
rect 31186 8213 31210 8247
rect 31244 8213 31260 8247
rect 31433 8275 31463 8297
rect 31433 8259 31497 8275
rect 31332 8226 31362 8241
rect 31186 8203 31260 8213
rect 31025 8129 31041 8143
rect 30975 8119 31041 8129
rect 30838 8083 30933 8099
rect 30903 8003 30933 8083
rect 30988 8003 31018 8119
rect 31083 8085 31144 8101
rect 31083 8051 31100 8085
rect 31134 8051 31144 8085
rect 31083 8035 31144 8051
rect 31083 8003 31113 8035
rect 31186 8003 31216 8203
rect 31318 8196 31362 8226
rect 31433 8225 31453 8259
rect 31487 8225 31497 8259
rect 31433 8209 31497 8225
rect 31318 8161 31348 8196
rect 31539 8167 31569 8297
rect 31258 8151 31348 8161
rect 31258 8117 31274 8151
rect 31308 8117 31348 8151
rect 31258 8107 31348 8117
rect 31318 8069 31348 8107
rect 31400 8151 31569 8167
rect 31400 8117 31410 8151
rect 31444 8137 31569 8151
rect 31444 8117 31454 8137
rect 31400 8101 31454 8117
rect 31634 8101 31664 8285
rect 32096 8270 32126 8285
rect 32085 8246 32126 8270
rect 31824 8217 31854 8239
rect 31908 8217 31938 8239
rect 32085 8217 32115 8246
rect 33329 8270 33359 8285
rect 33296 8240 33359 8270
rect 32191 8217 32221 8239
rect 32420 8217 32450 8239
rect 32665 8217 32695 8239
rect 32749 8217 32779 8239
rect 32833 8217 32863 8239
rect 32917 8217 32947 8239
rect 33296 8217 33326 8240
rect 31712 8201 31854 8217
rect 31712 8167 31722 8201
rect 31756 8167 31854 8201
rect 31712 8151 31854 8167
rect 31896 8201 32115 8217
rect 31896 8167 31906 8201
rect 31940 8167 32115 8201
rect 31896 8151 32115 8167
rect 32157 8201 32221 8217
rect 32157 8167 32167 8201
rect 32201 8167 32221 8201
rect 32157 8151 32221 8167
rect 32364 8201 32450 8217
rect 32364 8167 32380 8201
rect 32414 8167 32450 8201
rect 32364 8151 32450 8167
rect 32597 8201 32947 8217
rect 32597 8167 32613 8201
rect 32647 8167 32705 8201
rect 32739 8167 32789 8201
rect 32823 8167 32873 8201
rect 32907 8167 32947 8201
rect 32597 8151 32947 8167
rect 33272 8201 33326 8217
rect 33272 8167 33282 8201
rect 33316 8167 33326 8201
rect 33413 8196 33443 8285
rect 33272 8151 33326 8167
rect 31822 8119 31852 8151
rect 31906 8119 31936 8151
rect 30631 7899 30661 7925
rect 30715 7899 30745 7925
rect 31413 8003 31443 8101
rect 31496 8085 31562 8095
rect 31496 8051 31512 8085
rect 31546 8051 31562 8085
rect 31496 8041 31562 8051
rect 31611 8085 31692 8101
rect 31611 8051 31648 8085
rect 31682 8051 31692 8085
rect 31497 8003 31527 8041
rect 31611 8035 31692 8051
rect 31611 8003 31641 8035
rect 32085 8113 32115 8151
rect 32191 8119 32221 8151
rect 32420 8119 32450 8151
rect 32665 8119 32695 8151
rect 32749 8119 32779 8151
rect 32833 8119 32863 8151
rect 32917 8119 32947 8151
rect 32085 8083 32124 8113
rect 32094 8047 32124 8083
rect 33296 8098 33326 8151
rect 33368 8186 33443 8196
rect 33368 8152 33384 8186
rect 33418 8152 33443 8186
rect 33368 8142 33443 8152
rect 33601 8149 33631 8285
rect 33713 8269 33743 8297
rect 33693 8259 33759 8269
rect 33693 8225 33709 8259
rect 33743 8225 33759 8259
rect 33693 8215 33759 8225
rect 33812 8173 33842 8297
rect 33911 8257 33941 8285
rect 33296 8068 33359 8098
rect 33329 8053 33359 8068
rect 33413 8053 33443 8142
rect 33536 8133 33631 8149
rect 33536 8099 33546 8133
rect 33580 8099 33631 8133
rect 33673 8163 33842 8173
rect 33673 8129 33689 8163
rect 33723 8143 33842 8163
rect 33884 8247 33958 8257
rect 33884 8213 33908 8247
rect 33942 8213 33958 8247
rect 34131 8275 34161 8297
rect 34131 8259 34195 8275
rect 34030 8226 34060 8241
rect 33884 8203 33958 8213
rect 33723 8129 33739 8143
rect 33673 8119 33739 8129
rect 33536 8083 33631 8099
rect 33601 8003 33631 8083
rect 33686 8003 33716 8119
rect 33781 8085 33842 8101
rect 33781 8051 33798 8085
rect 33832 8051 33842 8085
rect 33781 8035 33842 8051
rect 33781 8003 33811 8035
rect 33884 8003 33914 8203
rect 34016 8196 34060 8226
rect 34131 8225 34151 8259
rect 34185 8225 34195 8259
rect 34131 8209 34195 8225
rect 34016 8161 34046 8196
rect 34237 8167 34267 8297
rect 33956 8151 34046 8161
rect 33956 8117 33972 8151
rect 34006 8117 34046 8151
rect 33956 8107 34046 8117
rect 34016 8069 34046 8107
rect 34098 8151 34267 8167
rect 34098 8117 34108 8151
rect 34142 8137 34267 8151
rect 34142 8117 34152 8137
rect 34098 8101 34152 8117
rect 34332 8101 34362 8285
rect 34794 8270 34824 8285
rect 34783 8246 34824 8270
rect 34522 8217 34552 8239
rect 34606 8217 34636 8239
rect 34783 8217 34813 8246
rect 34889 8217 34919 8239
rect 35118 8217 35148 8239
rect 35363 8217 35393 8239
rect 35447 8217 35477 8239
rect 35531 8217 35561 8239
rect 35615 8217 35645 8239
rect 34410 8201 34552 8217
rect 34410 8167 34420 8201
rect 34454 8167 34552 8201
rect 34410 8151 34552 8167
rect 34594 8201 34813 8217
rect 34594 8167 34604 8201
rect 34638 8167 34813 8201
rect 34594 8151 34813 8167
rect 34855 8201 34919 8217
rect 34855 8167 34865 8201
rect 34899 8167 34919 8201
rect 34855 8151 34919 8167
rect 35062 8201 35148 8217
rect 35062 8167 35078 8201
rect 35112 8167 35148 8201
rect 35062 8151 35148 8167
rect 35295 8201 35645 8217
rect 35295 8167 35311 8201
rect 35345 8167 35403 8201
rect 35437 8167 35487 8201
rect 35521 8167 35571 8201
rect 35605 8167 35645 8201
rect 35295 8151 35645 8167
rect 34520 8119 34550 8151
rect 34604 8119 34634 8151
rect 30903 7893 30933 7919
rect 30988 7893 31018 7919
rect 31083 7893 31113 7919
rect 31186 7893 31216 7919
rect 31318 7893 31348 7919
rect 31413 7893 31443 7919
rect 31497 7893 31527 7919
rect 31611 7893 31641 7919
rect 31822 7893 31852 7919
rect 31906 7893 31936 7919
rect 32094 7893 32124 7919
rect 32191 7893 32221 7919
rect 32420 7893 32450 7919
rect 32665 7893 32695 7919
rect 32749 7893 32779 7919
rect 32833 7893 32863 7919
rect 32917 7893 32947 7919
rect 33329 7899 33359 7925
rect 33413 7899 33443 7925
rect 34111 8003 34141 8101
rect 34194 8085 34260 8095
rect 34194 8051 34210 8085
rect 34244 8051 34260 8085
rect 34194 8041 34260 8051
rect 34309 8085 34390 8101
rect 34309 8051 34346 8085
rect 34380 8051 34390 8085
rect 34195 8003 34225 8041
rect 34309 8035 34390 8051
rect 34309 8003 34339 8035
rect 34783 8113 34813 8151
rect 34889 8119 34919 8151
rect 35118 8119 35148 8151
rect 35363 8119 35393 8151
rect 35447 8119 35477 8151
rect 35531 8119 35561 8151
rect 35615 8119 35645 8151
rect 34783 8083 34822 8113
rect 34792 8047 34822 8083
rect 33601 7893 33631 7919
rect 33686 7893 33716 7919
rect 33781 7893 33811 7919
rect 33884 7893 33914 7919
rect 34016 7893 34046 7919
rect 34111 7893 34141 7919
rect 34195 7893 34225 7919
rect 34309 7893 34339 7919
rect 34520 7893 34550 7919
rect 34604 7893 34634 7919
rect 34792 7893 34822 7919
rect 34889 7893 34919 7919
rect 35118 7893 35148 7919
rect 35363 7893 35393 7919
rect 35447 7893 35477 7919
rect 35531 7893 35561 7919
rect 35615 7893 35645 7919
rect 30631 7819 30661 7845
rect 30715 7819 30745 7845
rect 30903 7825 30933 7851
rect 30988 7825 31018 7851
rect 31083 7825 31113 7851
rect 31186 7825 31216 7851
rect 31318 7825 31348 7851
rect 31413 7825 31443 7851
rect 31497 7825 31527 7851
rect 31611 7825 31641 7851
rect 31822 7825 31852 7851
rect 31906 7825 31936 7851
rect 32094 7825 32124 7851
rect 32191 7825 32221 7851
rect 32420 7825 32450 7851
rect 32665 7825 32695 7851
rect 32749 7825 32779 7851
rect 32833 7825 32863 7851
rect 32917 7825 32947 7851
rect 30631 7676 30661 7691
rect 30598 7646 30661 7676
rect 30598 7593 30628 7646
rect 30715 7602 30745 7691
rect 30903 7661 30933 7741
rect 30574 7577 30628 7593
rect 30574 7543 30584 7577
rect 30618 7543 30628 7577
rect 30670 7592 30745 7602
rect 30838 7645 30933 7661
rect 30838 7611 30848 7645
rect 30882 7611 30933 7645
rect 30988 7625 31018 7741
rect 31083 7709 31113 7741
rect 31083 7693 31144 7709
rect 31083 7659 31100 7693
rect 31134 7659 31144 7693
rect 31083 7643 31144 7659
rect 30838 7595 30933 7611
rect 30670 7558 30686 7592
rect 30720 7558 30745 7592
rect 30670 7548 30745 7558
rect 30574 7527 30628 7543
rect 30598 7504 30628 7527
rect 30598 7474 30661 7504
rect 30631 7459 30661 7474
rect 30715 7459 30745 7548
rect 30903 7459 30933 7595
rect 30975 7615 31041 7625
rect 30975 7581 30991 7615
rect 31025 7601 31041 7615
rect 31025 7581 31144 7601
rect 30975 7571 31144 7581
rect 30995 7519 31061 7529
rect 30995 7485 31011 7519
rect 31045 7485 31061 7519
rect 30995 7475 31061 7485
rect 31015 7447 31045 7475
rect 31114 7447 31144 7571
rect 31186 7541 31216 7741
rect 31318 7637 31348 7675
rect 31413 7643 31443 7741
rect 31497 7703 31527 7741
rect 31611 7709 31641 7741
rect 31496 7693 31562 7703
rect 31496 7659 31512 7693
rect 31546 7659 31562 7693
rect 31496 7649 31562 7659
rect 31611 7693 31692 7709
rect 31611 7659 31648 7693
rect 31682 7659 31692 7693
rect 31611 7643 31692 7659
rect 31258 7627 31348 7637
rect 31258 7593 31274 7627
rect 31308 7593 31348 7627
rect 31258 7583 31348 7593
rect 31318 7548 31348 7583
rect 31400 7627 31454 7643
rect 31400 7593 31410 7627
rect 31444 7607 31454 7627
rect 31444 7593 31569 7607
rect 31400 7577 31569 7593
rect 31186 7531 31260 7541
rect 31186 7497 31210 7531
rect 31244 7497 31260 7531
rect 31318 7518 31362 7548
rect 31332 7503 31362 7518
rect 31433 7519 31497 7535
rect 31186 7487 31260 7497
rect 31213 7459 31243 7487
rect 31433 7485 31453 7519
rect 31487 7485 31497 7519
rect 31433 7469 31497 7485
rect 31433 7447 31463 7469
rect 31539 7447 31569 7577
rect 31634 7459 31664 7643
rect 32094 7661 32124 7697
rect 32085 7631 32124 7661
rect 31822 7593 31852 7625
rect 31906 7593 31936 7625
rect 32085 7593 32115 7631
rect 33329 7819 33359 7845
rect 33413 7819 33443 7845
rect 33601 7825 33631 7851
rect 33686 7825 33716 7851
rect 33781 7825 33811 7851
rect 33884 7825 33914 7851
rect 34016 7825 34046 7851
rect 34111 7825 34141 7851
rect 34195 7825 34225 7851
rect 34309 7825 34339 7851
rect 34520 7825 34550 7851
rect 34604 7825 34634 7851
rect 34792 7825 34822 7851
rect 34889 7825 34919 7851
rect 35118 7825 35148 7851
rect 35363 7825 35393 7851
rect 35447 7825 35477 7851
rect 35531 7825 35561 7851
rect 35615 7825 35645 7851
rect 33329 7676 33359 7691
rect 33296 7646 33359 7676
rect 32191 7593 32221 7625
rect 32420 7593 32450 7625
rect 32665 7593 32695 7625
rect 32749 7593 32779 7625
rect 32833 7593 32863 7625
rect 32917 7593 32947 7625
rect 33296 7593 33326 7646
rect 33413 7602 33443 7691
rect 33601 7661 33631 7741
rect 31712 7577 31854 7593
rect 31712 7543 31722 7577
rect 31756 7543 31854 7577
rect 31712 7527 31854 7543
rect 31896 7577 32115 7593
rect 31896 7543 31906 7577
rect 31940 7543 32115 7577
rect 31896 7527 32115 7543
rect 32157 7577 32221 7593
rect 32157 7543 32167 7577
rect 32201 7543 32221 7577
rect 32157 7527 32221 7543
rect 32364 7577 32450 7593
rect 32364 7543 32380 7577
rect 32414 7543 32450 7577
rect 32364 7527 32450 7543
rect 32597 7577 32947 7593
rect 32597 7543 32613 7577
rect 32647 7543 32705 7577
rect 32739 7543 32789 7577
rect 32823 7543 32873 7577
rect 32907 7543 32947 7577
rect 32597 7527 32947 7543
rect 33272 7577 33326 7593
rect 33272 7543 33282 7577
rect 33316 7543 33326 7577
rect 33368 7592 33443 7602
rect 33536 7645 33631 7661
rect 33536 7611 33546 7645
rect 33580 7611 33631 7645
rect 33686 7625 33716 7741
rect 33781 7709 33811 7741
rect 33781 7693 33842 7709
rect 33781 7659 33798 7693
rect 33832 7659 33842 7693
rect 33781 7643 33842 7659
rect 33536 7595 33631 7611
rect 33368 7558 33384 7592
rect 33418 7558 33443 7592
rect 33368 7548 33443 7558
rect 33272 7527 33326 7543
rect 31824 7505 31854 7527
rect 31908 7505 31938 7527
rect 32085 7498 32115 7527
rect 32191 7505 32221 7527
rect 32420 7505 32450 7527
rect 32665 7505 32695 7527
rect 32749 7505 32779 7527
rect 32833 7505 32863 7527
rect 32917 7505 32947 7527
rect 32085 7474 32126 7498
rect 32096 7459 32126 7474
rect 33296 7504 33326 7527
rect 33296 7474 33359 7504
rect 33329 7459 33359 7474
rect 33413 7459 33443 7548
rect 33601 7459 33631 7595
rect 33673 7615 33739 7625
rect 33673 7581 33689 7615
rect 33723 7601 33739 7615
rect 33723 7581 33842 7601
rect 33673 7571 33842 7581
rect 33693 7519 33759 7529
rect 33693 7485 33709 7519
rect 33743 7485 33759 7519
rect 33693 7475 33759 7485
rect 33713 7447 33743 7475
rect 33812 7447 33842 7571
rect 33884 7541 33914 7741
rect 34016 7637 34046 7675
rect 34111 7643 34141 7741
rect 34195 7703 34225 7741
rect 34309 7709 34339 7741
rect 34194 7693 34260 7703
rect 34194 7659 34210 7693
rect 34244 7659 34260 7693
rect 34194 7649 34260 7659
rect 34309 7693 34390 7709
rect 34309 7659 34346 7693
rect 34380 7659 34390 7693
rect 34309 7643 34390 7659
rect 33956 7627 34046 7637
rect 33956 7593 33972 7627
rect 34006 7593 34046 7627
rect 33956 7583 34046 7593
rect 34016 7548 34046 7583
rect 34098 7627 34152 7643
rect 34098 7593 34108 7627
rect 34142 7607 34152 7627
rect 34142 7593 34267 7607
rect 34098 7577 34267 7593
rect 33884 7531 33958 7541
rect 33884 7497 33908 7531
rect 33942 7497 33958 7531
rect 34016 7518 34060 7548
rect 34030 7503 34060 7518
rect 34131 7519 34195 7535
rect 33884 7487 33958 7497
rect 33911 7459 33941 7487
rect 34131 7485 34151 7519
rect 34185 7485 34195 7519
rect 34131 7469 34195 7485
rect 34131 7447 34161 7469
rect 34237 7447 34267 7577
rect 34332 7459 34362 7643
rect 34792 7661 34822 7697
rect 34783 7631 34822 7661
rect 34520 7593 34550 7625
rect 34604 7593 34634 7625
rect 34783 7593 34813 7631
rect 34889 7593 34919 7625
rect 35118 7593 35148 7625
rect 35363 7593 35393 7625
rect 35447 7593 35477 7625
rect 35531 7593 35561 7625
rect 35615 7593 35645 7625
rect 34410 7577 34552 7593
rect 34410 7543 34420 7577
rect 34454 7543 34552 7577
rect 34410 7527 34552 7543
rect 34594 7577 34813 7593
rect 34594 7543 34604 7577
rect 34638 7543 34813 7577
rect 34594 7527 34813 7543
rect 34855 7577 34919 7593
rect 34855 7543 34865 7577
rect 34899 7543 34919 7577
rect 34855 7527 34919 7543
rect 35062 7577 35148 7593
rect 35062 7543 35078 7577
rect 35112 7543 35148 7577
rect 35062 7527 35148 7543
rect 35295 7577 35645 7593
rect 35295 7543 35311 7577
rect 35345 7543 35403 7577
rect 35437 7543 35487 7577
rect 35521 7543 35571 7577
rect 35605 7543 35645 7577
rect 35295 7527 35645 7543
rect 34522 7505 34552 7527
rect 34606 7505 34636 7527
rect 34783 7498 34813 7527
rect 34889 7505 34919 7527
rect 35118 7505 35148 7527
rect 35363 7505 35393 7527
rect 35447 7505 35477 7527
rect 35531 7505 35561 7527
rect 35615 7505 35645 7527
rect 34783 7474 34824 7498
rect 34794 7459 34824 7474
rect 30631 7349 30661 7375
rect 30715 7349 30745 7375
rect 30903 7349 30933 7375
rect 31015 7349 31045 7375
rect 31114 7349 31144 7375
rect 31213 7349 31243 7375
rect 31332 7349 31362 7375
rect 31433 7349 31463 7375
rect 31539 7349 31569 7375
rect 31634 7349 31664 7375
rect 31824 7349 31854 7375
rect 31908 7349 31938 7375
rect 32096 7349 32126 7375
rect 32191 7349 32221 7375
rect 32420 7349 32450 7375
rect 32665 7349 32695 7375
rect 32749 7349 32779 7375
rect 32833 7349 32863 7375
rect 32917 7349 32947 7375
rect 33329 7349 33359 7375
rect 33413 7349 33443 7375
rect 33601 7349 33631 7375
rect 33713 7349 33743 7375
rect 33812 7349 33842 7375
rect 33911 7349 33941 7375
rect 34030 7349 34060 7375
rect 34131 7349 34161 7375
rect 34237 7349 34267 7375
rect 34332 7349 34362 7375
rect 34522 7349 34552 7375
rect 34606 7349 34636 7375
rect 34794 7349 34824 7375
rect 34889 7349 34919 7375
rect 35118 7349 35148 7375
rect 35363 7349 35393 7375
rect 35447 7349 35477 7375
rect 35531 7349 35561 7375
rect 35615 7349 35645 7375
rect 30631 7281 30661 7307
rect 30715 7281 30745 7307
rect 30903 7281 30933 7307
rect 31015 7281 31045 7307
rect 31114 7281 31144 7307
rect 31213 7281 31243 7307
rect 31332 7281 31362 7307
rect 31433 7281 31463 7307
rect 31539 7281 31569 7307
rect 31634 7281 31664 7307
rect 31824 7281 31854 7307
rect 31908 7281 31938 7307
rect 32096 7281 32126 7307
rect 32191 7281 32221 7307
rect 32420 7281 32450 7307
rect 32665 7281 32695 7307
rect 32749 7281 32779 7307
rect 32833 7281 32863 7307
rect 32917 7281 32947 7307
rect 33329 7281 33359 7307
rect 33413 7281 33443 7307
rect 33601 7281 33631 7307
rect 33713 7281 33743 7307
rect 33812 7281 33842 7307
rect 33911 7281 33941 7307
rect 34030 7281 34060 7307
rect 34131 7281 34161 7307
rect 34237 7281 34267 7307
rect 34332 7281 34362 7307
rect 34522 7281 34552 7307
rect 34606 7281 34636 7307
rect 34794 7281 34824 7307
rect 34889 7281 34919 7307
rect 35118 7281 35148 7307
rect 35363 7281 35393 7307
rect 35447 7281 35477 7307
rect 35531 7281 35561 7307
rect 35615 7281 35645 7307
rect 30631 7182 30661 7197
rect 30598 7152 30661 7182
rect 30598 7129 30628 7152
rect 30574 7113 30628 7129
rect 30574 7079 30584 7113
rect 30618 7079 30628 7113
rect 30715 7108 30745 7197
rect 30574 7063 30628 7079
rect 30598 7010 30628 7063
rect 30670 7098 30745 7108
rect 30670 7064 30686 7098
rect 30720 7064 30745 7098
rect 30670 7054 30745 7064
rect 30903 7061 30933 7197
rect 31015 7181 31045 7209
rect 30995 7171 31061 7181
rect 30995 7137 31011 7171
rect 31045 7137 31061 7171
rect 30995 7127 31061 7137
rect 31114 7085 31144 7209
rect 31213 7169 31243 7197
rect 30598 6980 30661 7010
rect 30631 6965 30661 6980
rect 30715 6965 30745 7054
rect 30838 7045 30933 7061
rect 30838 7011 30848 7045
rect 30882 7011 30933 7045
rect 30975 7075 31144 7085
rect 30975 7041 30991 7075
rect 31025 7055 31144 7075
rect 31186 7159 31260 7169
rect 31186 7125 31210 7159
rect 31244 7125 31260 7159
rect 31433 7187 31463 7209
rect 31433 7171 31497 7187
rect 31332 7138 31362 7153
rect 31186 7115 31260 7125
rect 31025 7041 31041 7055
rect 30975 7031 31041 7041
rect 30838 6995 30933 7011
rect 30903 6915 30933 6995
rect 30988 6915 31018 7031
rect 31083 6997 31144 7013
rect 31083 6963 31100 6997
rect 31134 6963 31144 6997
rect 31083 6947 31144 6963
rect 31083 6915 31113 6947
rect 31186 6915 31216 7115
rect 31318 7108 31362 7138
rect 31433 7137 31453 7171
rect 31487 7137 31497 7171
rect 31433 7121 31497 7137
rect 31318 7073 31348 7108
rect 31539 7079 31569 7209
rect 31258 7063 31348 7073
rect 31258 7029 31274 7063
rect 31308 7029 31348 7063
rect 31258 7019 31348 7029
rect 31318 6981 31348 7019
rect 31400 7063 31569 7079
rect 31400 7029 31410 7063
rect 31444 7049 31569 7063
rect 31444 7029 31454 7049
rect 31400 7013 31454 7029
rect 31634 7013 31664 7197
rect 32096 7182 32126 7197
rect 32085 7158 32126 7182
rect 31824 7129 31854 7151
rect 31908 7129 31938 7151
rect 32085 7129 32115 7158
rect 33329 7182 33359 7197
rect 33296 7152 33359 7182
rect 32191 7129 32221 7151
rect 32420 7129 32450 7151
rect 32665 7129 32695 7151
rect 32749 7129 32779 7151
rect 32833 7129 32863 7151
rect 32917 7129 32947 7151
rect 33296 7129 33326 7152
rect 31712 7113 31854 7129
rect 31712 7079 31722 7113
rect 31756 7079 31854 7113
rect 31712 7063 31854 7079
rect 31896 7113 32115 7129
rect 31896 7079 31906 7113
rect 31940 7079 32115 7113
rect 31896 7063 32115 7079
rect 32157 7113 32221 7129
rect 32157 7079 32167 7113
rect 32201 7079 32221 7113
rect 32157 7063 32221 7079
rect 32364 7113 32450 7129
rect 32364 7079 32380 7113
rect 32414 7079 32450 7113
rect 32364 7063 32450 7079
rect 32597 7113 32947 7129
rect 32597 7079 32613 7113
rect 32647 7079 32705 7113
rect 32739 7079 32789 7113
rect 32823 7079 32873 7113
rect 32907 7079 32947 7113
rect 32597 7063 32947 7079
rect 33272 7113 33326 7129
rect 33272 7079 33282 7113
rect 33316 7079 33326 7113
rect 33413 7108 33443 7197
rect 33272 7063 33326 7079
rect 31822 7031 31852 7063
rect 31906 7031 31936 7063
rect 30631 6811 30661 6837
rect 30715 6811 30745 6837
rect 31413 6915 31443 7013
rect 31496 6997 31562 7007
rect 31496 6963 31512 6997
rect 31546 6963 31562 6997
rect 31496 6953 31562 6963
rect 31611 6997 31692 7013
rect 31611 6963 31648 6997
rect 31682 6963 31692 6997
rect 31497 6915 31527 6953
rect 31611 6947 31692 6963
rect 31611 6915 31641 6947
rect 32085 7025 32115 7063
rect 32191 7031 32221 7063
rect 32420 7031 32450 7063
rect 32665 7031 32695 7063
rect 32749 7031 32779 7063
rect 32833 7031 32863 7063
rect 32917 7031 32947 7063
rect 32085 6995 32124 7025
rect 32094 6959 32124 6995
rect 33296 7010 33326 7063
rect 33368 7098 33443 7108
rect 33368 7064 33384 7098
rect 33418 7064 33443 7098
rect 33368 7054 33443 7064
rect 33601 7061 33631 7197
rect 33713 7181 33743 7209
rect 33693 7171 33759 7181
rect 33693 7137 33709 7171
rect 33743 7137 33759 7171
rect 33693 7127 33759 7137
rect 33812 7085 33842 7209
rect 33911 7169 33941 7197
rect 33296 6980 33359 7010
rect 33329 6965 33359 6980
rect 33413 6965 33443 7054
rect 33536 7045 33631 7061
rect 33536 7011 33546 7045
rect 33580 7011 33631 7045
rect 33673 7075 33842 7085
rect 33673 7041 33689 7075
rect 33723 7055 33842 7075
rect 33884 7159 33958 7169
rect 33884 7125 33908 7159
rect 33942 7125 33958 7159
rect 34131 7187 34161 7209
rect 34131 7171 34195 7187
rect 34030 7138 34060 7153
rect 33884 7115 33958 7125
rect 33723 7041 33739 7055
rect 33673 7031 33739 7041
rect 33536 6995 33631 7011
rect 33601 6915 33631 6995
rect 33686 6915 33716 7031
rect 33781 6997 33842 7013
rect 33781 6963 33798 6997
rect 33832 6963 33842 6997
rect 33781 6947 33842 6963
rect 33781 6915 33811 6947
rect 33884 6915 33914 7115
rect 34016 7108 34060 7138
rect 34131 7137 34151 7171
rect 34185 7137 34195 7171
rect 34131 7121 34195 7137
rect 34016 7073 34046 7108
rect 34237 7079 34267 7209
rect 33956 7063 34046 7073
rect 33956 7029 33972 7063
rect 34006 7029 34046 7063
rect 33956 7019 34046 7029
rect 34016 6981 34046 7019
rect 34098 7063 34267 7079
rect 34098 7029 34108 7063
rect 34142 7049 34267 7063
rect 34142 7029 34152 7049
rect 34098 7013 34152 7029
rect 34332 7013 34362 7197
rect 34794 7182 34824 7197
rect 34783 7158 34824 7182
rect 34522 7129 34552 7151
rect 34606 7129 34636 7151
rect 34783 7129 34813 7158
rect 34889 7129 34919 7151
rect 35118 7129 35148 7151
rect 35363 7129 35393 7151
rect 35447 7129 35477 7151
rect 35531 7129 35561 7151
rect 35615 7129 35645 7151
rect 34410 7113 34552 7129
rect 34410 7079 34420 7113
rect 34454 7079 34552 7113
rect 34410 7063 34552 7079
rect 34594 7113 34813 7129
rect 34594 7079 34604 7113
rect 34638 7079 34813 7113
rect 34594 7063 34813 7079
rect 34855 7113 34919 7129
rect 34855 7079 34865 7113
rect 34899 7079 34919 7113
rect 34855 7063 34919 7079
rect 35062 7113 35148 7129
rect 35062 7079 35078 7113
rect 35112 7079 35148 7113
rect 35062 7063 35148 7079
rect 35295 7113 35645 7129
rect 35295 7079 35311 7113
rect 35345 7079 35403 7113
rect 35437 7079 35487 7113
rect 35521 7079 35571 7113
rect 35605 7079 35645 7113
rect 35295 7063 35645 7079
rect 34520 7031 34550 7063
rect 34604 7031 34634 7063
rect 30903 6805 30933 6831
rect 30988 6805 31018 6831
rect 31083 6805 31113 6831
rect 31186 6805 31216 6831
rect 31318 6805 31348 6831
rect 31413 6805 31443 6831
rect 31497 6805 31527 6831
rect 31611 6805 31641 6831
rect 31822 6805 31852 6831
rect 31906 6805 31936 6831
rect 32094 6805 32124 6831
rect 32191 6805 32221 6831
rect 32420 6805 32450 6831
rect 32665 6805 32695 6831
rect 32749 6805 32779 6831
rect 32833 6805 32863 6831
rect 32917 6805 32947 6831
rect 33329 6811 33359 6837
rect 33413 6811 33443 6837
rect 34111 6915 34141 7013
rect 34194 6997 34260 7007
rect 34194 6963 34210 6997
rect 34244 6963 34260 6997
rect 34194 6953 34260 6963
rect 34309 6997 34390 7013
rect 34309 6963 34346 6997
rect 34380 6963 34390 6997
rect 34195 6915 34225 6953
rect 34309 6947 34390 6963
rect 34309 6915 34339 6947
rect 34783 7025 34813 7063
rect 34889 7031 34919 7063
rect 35118 7031 35148 7063
rect 35363 7031 35393 7063
rect 35447 7031 35477 7063
rect 35531 7031 35561 7063
rect 35615 7031 35645 7063
rect 34783 6995 34822 7025
rect 34792 6959 34822 6995
rect 33601 6805 33631 6831
rect 33686 6805 33716 6831
rect 33781 6805 33811 6831
rect 33884 6805 33914 6831
rect 34016 6805 34046 6831
rect 34111 6805 34141 6831
rect 34195 6805 34225 6831
rect 34309 6805 34339 6831
rect 34520 6805 34550 6831
rect 34604 6805 34634 6831
rect 34792 6805 34822 6831
rect 34889 6805 34919 6831
rect 35118 6805 35148 6831
rect 35363 6805 35393 6831
rect 35447 6805 35477 6831
rect 35531 6805 35561 6831
rect 35615 6805 35645 6831
rect 30631 6731 30661 6757
rect 30715 6731 30745 6757
rect 30903 6737 30933 6763
rect 30988 6737 31018 6763
rect 31083 6737 31113 6763
rect 31186 6737 31216 6763
rect 31318 6737 31348 6763
rect 31413 6737 31443 6763
rect 31497 6737 31527 6763
rect 31611 6737 31641 6763
rect 31822 6737 31852 6763
rect 31906 6737 31936 6763
rect 32094 6737 32124 6763
rect 32191 6737 32221 6763
rect 32420 6737 32450 6763
rect 32665 6737 32695 6763
rect 32749 6737 32779 6763
rect 32833 6737 32863 6763
rect 32917 6737 32947 6763
rect 30631 6588 30661 6603
rect 30598 6558 30661 6588
rect 30598 6505 30628 6558
rect 30715 6514 30745 6603
rect 30903 6573 30933 6653
rect 30574 6489 30628 6505
rect 30574 6455 30584 6489
rect 30618 6455 30628 6489
rect 30670 6504 30745 6514
rect 30838 6557 30933 6573
rect 30838 6523 30848 6557
rect 30882 6523 30933 6557
rect 30988 6537 31018 6653
rect 31083 6621 31113 6653
rect 31083 6605 31144 6621
rect 31083 6571 31100 6605
rect 31134 6571 31144 6605
rect 31083 6555 31144 6571
rect 30838 6507 30933 6523
rect 30670 6470 30686 6504
rect 30720 6470 30745 6504
rect 30670 6460 30745 6470
rect 30574 6439 30628 6455
rect 30598 6416 30628 6439
rect 30598 6386 30661 6416
rect 30631 6371 30661 6386
rect 30715 6371 30745 6460
rect 30903 6371 30933 6507
rect 30975 6527 31041 6537
rect 30975 6493 30991 6527
rect 31025 6513 31041 6527
rect 31025 6493 31144 6513
rect 30975 6483 31144 6493
rect 30995 6431 31061 6441
rect 30995 6397 31011 6431
rect 31045 6397 31061 6431
rect 30995 6387 31061 6397
rect 31015 6359 31045 6387
rect 31114 6359 31144 6483
rect 31186 6453 31216 6653
rect 31318 6549 31348 6587
rect 31413 6555 31443 6653
rect 31497 6615 31527 6653
rect 31611 6621 31641 6653
rect 31496 6605 31562 6615
rect 31496 6571 31512 6605
rect 31546 6571 31562 6605
rect 31496 6561 31562 6571
rect 31611 6605 31692 6621
rect 31611 6571 31648 6605
rect 31682 6571 31692 6605
rect 31611 6555 31692 6571
rect 31258 6539 31348 6549
rect 31258 6505 31274 6539
rect 31308 6505 31348 6539
rect 31258 6495 31348 6505
rect 31318 6460 31348 6495
rect 31400 6539 31454 6555
rect 31400 6505 31410 6539
rect 31444 6519 31454 6539
rect 31444 6505 31569 6519
rect 31400 6489 31569 6505
rect 31186 6443 31260 6453
rect 31186 6409 31210 6443
rect 31244 6409 31260 6443
rect 31318 6430 31362 6460
rect 31332 6415 31362 6430
rect 31433 6431 31497 6447
rect 31186 6399 31260 6409
rect 31213 6371 31243 6399
rect 31433 6397 31453 6431
rect 31487 6397 31497 6431
rect 31433 6381 31497 6397
rect 31433 6359 31463 6381
rect 31539 6359 31569 6489
rect 31634 6371 31664 6555
rect 32094 6573 32124 6609
rect 32085 6543 32124 6573
rect 31822 6505 31852 6537
rect 31906 6505 31936 6537
rect 32085 6505 32115 6543
rect 33329 6731 33359 6757
rect 33413 6731 33443 6757
rect 33601 6737 33631 6763
rect 33686 6737 33716 6763
rect 33781 6737 33811 6763
rect 33884 6737 33914 6763
rect 34016 6737 34046 6763
rect 34111 6737 34141 6763
rect 34195 6737 34225 6763
rect 34309 6737 34339 6763
rect 34520 6737 34550 6763
rect 34604 6737 34634 6763
rect 34792 6737 34822 6763
rect 34889 6737 34919 6763
rect 35118 6737 35148 6763
rect 35363 6737 35393 6763
rect 35447 6737 35477 6763
rect 35531 6737 35561 6763
rect 35615 6737 35645 6763
rect 33329 6588 33359 6603
rect 33296 6558 33359 6588
rect 32191 6505 32221 6537
rect 32420 6505 32450 6537
rect 32665 6505 32695 6537
rect 32749 6505 32779 6537
rect 32833 6505 32863 6537
rect 32917 6505 32947 6537
rect 33296 6505 33326 6558
rect 33413 6514 33443 6603
rect 33601 6573 33631 6653
rect 31712 6489 31854 6505
rect 31712 6455 31722 6489
rect 31756 6455 31854 6489
rect 31712 6439 31854 6455
rect 31896 6489 32115 6505
rect 31896 6455 31906 6489
rect 31940 6455 32115 6489
rect 31896 6439 32115 6455
rect 32157 6489 32221 6505
rect 32157 6455 32167 6489
rect 32201 6455 32221 6489
rect 32157 6439 32221 6455
rect 32364 6489 32450 6505
rect 32364 6455 32380 6489
rect 32414 6455 32450 6489
rect 32364 6439 32450 6455
rect 32597 6489 32947 6505
rect 32597 6455 32613 6489
rect 32647 6455 32705 6489
rect 32739 6455 32789 6489
rect 32823 6455 32873 6489
rect 32907 6455 32947 6489
rect 32597 6439 32947 6455
rect 33272 6489 33326 6505
rect 33272 6455 33282 6489
rect 33316 6455 33326 6489
rect 33368 6504 33443 6514
rect 33536 6557 33631 6573
rect 33536 6523 33546 6557
rect 33580 6523 33631 6557
rect 33686 6537 33716 6653
rect 33781 6621 33811 6653
rect 33781 6605 33842 6621
rect 33781 6571 33798 6605
rect 33832 6571 33842 6605
rect 33781 6555 33842 6571
rect 33536 6507 33631 6523
rect 33368 6470 33384 6504
rect 33418 6470 33443 6504
rect 33368 6460 33443 6470
rect 33272 6439 33326 6455
rect 31824 6417 31854 6439
rect 31908 6417 31938 6439
rect 32085 6410 32115 6439
rect 32191 6417 32221 6439
rect 32420 6417 32450 6439
rect 32665 6417 32695 6439
rect 32749 6417 32779 6439
rect 32833 6417 32863 6439
rect 32917 6417 32947 6439
rect 32085 6386 32126 6410
rect 32096 6371 32126 6386
rect 33296 6416 33326 6439
rect 33296 6386 33359 6416
rect 33329 6371 33359 6386
rect 33413 6371 33443 6460
rect 33601 6371 33631 6507
rect 33673 6527 33739 6537
rect 33673 6493 33689 6527
rect 33723 6513 33739 6527
rect 33723 6493 33842 6513
rect 33673 6483 33842 6493
rect 33693 6431 33759 6441
rect 33693 6397 33709 6431
rect 33743 6397 33759 6431
rect 33693 6387 33759 6397
rect 33713 6359 33743 6387
rect 33812 6359 33842 6483
rect 33884 6453 33914 6653
rect 34016 6549 34046 6587
rect 34111 6555 34141 6653
rect 34195 6615 34225 6653
rect 34309 6621 34339 6653
rect 34194 6605 34260 6615
rect 34194 6571 34210 6605
rect 34244 6571 34260 6605
rect 34194 6561 34260 6571
rect 34309 6605 34390 6621
rect 34309 6571 34346 6605
rect 34380 6571 34390 6605
rect 34309 6555 34390 6571
rect 33956 6539 34046 6549
rect 33956 6505 33972 6539
rect 34006 6505 34046 6539
rect 33956 6495 34046 6505
rect 34016 6460 34046 6495
rect 34098 6539 34152 6555
rect 34098 6505 34108 6539
rect 34142 6519 34152 6539
rect 34142 6505 34267 6519
rect 34098 6489 34267 6505
rect 33884 6443 33958 6453
rect 33884 6409 33908 6443
rect 33942 6409 33958 6443
rect 34016 6430 34060 6460
rect 34030 6415 34060 6430
rect 34131 6431 34195 6447
rect 33884 6399 33958 6409
rect 33911 6371 33941 6399
rect 34131 6397 34151 6431
rect 34185 6397 34195 6431
rect 34131 6381 34195 6397
rect 34131 6359 34161 6381
rect 34237 6359 34267 6489
rect 34332 6371 34362 6555
rect 34792 6573 34822 6609
rect 34783 6543 34822 6573
rect 34520 6505 34550 6537
rect 34604 6505 34634 6537
rect 34783 6505 34813 6543
rect 34889 6505 34919 6537
rect 35118 6505 35148 6537
rect 35363 6505 35393 6537
rect 35447 6505 35477 6537
rect 35531 6505 35561 6537
rect 35615 6505 35645 6537
rect 34410 6489 34552 6505
rect 34410 6455 34420 6489
rect 34454 6455 34552 6489
rect 34410 6439 34552 6455
rect 34594 6489 34813 6505
rect 34594 6455 34604 6489
rect 34638 6455 34813 6489
rect 34594 6439 34813 6455
rect 34855 6489 34919 6505
rect 34855 6455 34865 6489
rect 34899 6455 34919 6489
rect 34855 6439 34919 6455
rect 35062 6489 35148 6505
rect 35062 6455 35078 6489
rect 35112 6455 35148 6489
rect 35062 6439 35148 6455
rect 35295 6489 35645 6505
rect 35295 6455 35311 6489
rect 35345 6455 35403 6489
rect 35437 6455 35487 6489
rect 35521 6455 35571 6489
rect 35605 6455 35645 6489
rect 35295 6439 35645 6455
rect 34522 6417 34552 6439
rect 34606 6417 34636 6439
rect 34783 6410 34813 6439
rect 34889 6417 34919 6439
rect 35118 6417 35148 6439
rect 35363 6417 35393 6439
rect 35447 6417 35477 6439
rect 35531 6417 35561 6439
rect 35615 6417 35645 6439
rect 34783 6386 34824 6410
rect 34794 6371 34824 6386
rect 30631 6261 30661 6287
rect 30715 6261 30745 6287
rect 30903 6261 30933 6287
rect 31015 6261 31045 6287
rect 31114 6261 31144 6287
rect 31213 6261 31243 6287
rect 31332 6261 31362 6287
rect 31433 6261 31463 6287
rect 31539 6261 31569 6287
rect 31634 6261 31664 6287
rect 31824 6261 31854 6287
rect 31908 6261 31938 6287
rect 32096 6261 32126 6287
rect 32191 6261 32221 6287
rect 32420 6261 32450 6287
rect 32665 6261 32695 6287
rect 32749 6261 32779 6287
rect 32833 6261 32863 6287
rect 32917 6261 32947 6287
rect 33329 6261 33359 6287
rect 33413 6261 33443 6287
rect 33601 6261 33631 6287
rect 33713 6261 33743 6287
rect 33812 6261 33842 6287
rect 33911 6261 33941 6287
rect 34030 6261 34060 6287
rect 34131 6261 34161 6287
rect 34237 6261 34267 6287
rect 34332 6261 34362 6287
rect 34522 6261 34552 6287
rect 34606 6261 34636 6287
rect 34794 6261 34824 6287
rect 34889 6261 34919 6287
rect 35118 6261 35148 6287
rect 35363 6261 35393 6287
rect 35447 6261 35477 6287
rect 35531 6261 35561 6287
rect 35615 6261 35645 6287
rect 30631 6193 30661 6219
rect 30715 6193 30745 6219
rect 30903 6193 30933 6219
rect 31015 6193 31045 6219
rect 31114 6193 31144 6219
rect 31213 6193 31243 6219
rect 31332 6193 31362 6219
rect 31433 6193 31463 6219
rect 31539 6193 31569 6219
rect 31634 6193 31664 6219
rect 31824 6193 31854 6219
rect 31908 6193 31938 6219
rect 32096 6193 32126 6219
rect 32191 6193 32221 6219
rect 32420 6193 32450 6219
rect 32665 6193 32695 6219
rect 32749 6193 32779 6219
rect 32833 6193 32863 6219
rect 32917 6193 32947 6219
rect 33329 6193 33359 6219
rect 33413 6193 33443 6219
rect 33601 6193 33631 6219
rect 33713 6193 33743 6219
rect 33812 6193 33842 6219
rect 33911 6193 33941 6219
rect 34030 6193 34060 6219
rect 34131 6193 34161 6219
rect 34237 6193 34267 6219
rect 34332 6193 34362 6219
rect 34522 6193 34552 6219
rect 34606 6193 34636 6219
rect 34794 6193 34824 6219
rect 34889 6193 34919 6219
rect 35118 6193 35148 6219
rect 35363 6193 35393 6219
rect 35447 6193 35477 6219
rect 35531 6193 35561 6219
rect 35615 6193 35645 6219
rect 30631 6094 30661 6109
rect 30598 6064 30661 6094
rect 30598 6041 30628 6064
rect 30574 6025 30628 6041
rect 30574 5991 30584 6025
rect 30618 5991 30628 6025
rect 30715 6020 30745 6109
rect 30574 5975 30628 5991
rect 30598 5922 30628 5975
rect 30670 6010 30745 6020
rect 30670 5976 30686 6010
rect 30720 5976 30745 6010
rect 30670 5966 30745 5976
rect 30903 5973 30933 6109
rect 31015 6093 31045 6121
rect 30995 6083 31061 6093
rect 30995 6049 31011 6083
rect 31045 6049 31061 6083
rect 30995 6039 31061 6049
rect 31114 5997 31144 6121
rect 31213 6081 31243 6109
rect 30598 5892 30661 5922
rect 30631 5877 30661 5892
rect 30715 5877 30745 5966
rect 30838 5957 30933 5973
rect 30838 5923 30848 5957
rect 30882 5923 30933 5957
rect 30975 5987 31144 5997
rect 30975 5953 30991 5987
rect 31025 5967 31144 5987
rect 31186 6071 31260 6081
rect 31186 6037 31210 6071
rect 31244 6037 31260 6071
rect 31433 6099 31463 6121
rect 31433 6083 31497 6099
rect 31332 6050 31362 6065
rect 31186 6027 31260 6037
rect 31025 5953 31041 5967
rect 30975 5943 31041 5953
rect 30838 5907 30933 5923
rect 30903 5827 30933 5907
rect 30988 5827 31018 5943
rect 31083 5909 31144 5925
rect 31083 5875 31100 5909
rect 31134 5875 31144 5909
rect 31083 5859 31144 5875
rect 31083 5827 31113 5859
rect 31186 5827 31216 6027
rect 31318 6020 31362 6050
rect 31433 6049 31453 6083
rect 31487 6049 31497 6083
rect 31433 6033 31497 6049
rect 31318 5985 31348 6020
rect 31539 5991 31569 6121
rect 31258 5975 31348 5985
rect 31258 5941 31274 5975
rect 31308 5941 31348 5975
rect 31258 5931 31348 5941
rect 31318 5893 31348 5931
rect 31400 5975 31569 5991
rect 31400 5941 31410 5975
rect 31444 5961 31569 5975
rect 31444 5941 31454 5961
rect 31400 5925 31454 5941
rect 31634 5925 31664 6109
rect 32096 6094 32126 6109
rect 32085 6070 32126 6094
rect 31824 6041 31854 6063
rect 31908 6041 31938 6063
rect 32085 6041 32115 6070
rect 33329 6094 33359 6109
rect 33296 6064 33359 6094
rect 32191 6041 32221 6063
rect 32420 6041 32450 6063
rect 32665 6041 32695 6063
rect 32749 6041 32779 6063
rect 32833 6041 32863 6063
rect 32917 6041 32947 6063
rect 33296 6041 33326 6064
rect 31712 6025 31854 6041
rect 31712 5991 31722 6025
rect 31756 5991 31854 6025
rect 31712 5975 31854 5991
rect 31896 6025 32115 6041
rect 31896 5991 31906 6025
rect 31940 5991 32115 6025
rect 31896 5975 32115 5991
rect 32157 6025 32221 6041
rect 32157 5991 32167 6025
rect 32201 5991 32221 6025
rect 32157 5975 32221 5991
rect 32364 6025 32450 6041
rect 32364 5991 32380 6025
rect 32414 5991 32450 6025
rect 32364 5975 32450 5991
rect 32597 6025 32947 6041
rect 32597 5991 32613 6025
rect 32647 5991 32705 6025
rect 32739 5991 32789 6025
rect 32823 5991 32873 6025
rect 32907 5991 32947 6025
rect 32597 5975 32947 5991
rect 33272 6025 33326 6041
rect 33272 5991 33282 6025
rect 33316 5991 33326 6025
rect 33413 6020 33443 6109
rect 33272 5975 33326 5991
rect 31822 5943 31852 5975
rect 31906 5943 31936 5975
rect 30631 5723 30661 5749
rect 30715 5723 30745 5749
rect 31413 5827 31443 5925
rect 31496 5909 31562 5919
rect 31496 5875 31512 5909
rect 31546 5875 31562 5909
rect 31496 5865 31562 5875
rect 31611 5909 31692 5925
rect 31611 5875 31648 5909
rect 31682 5875 31692 5909
rect 31497 5827 31527 5865
rect 31611 5859 31692 5875
rect 31611 5827 31641 5859
rect 32085 5937 32115 5975
rect 32191 5943 32221 5975
rect 32420 5943 32450 5975
rect 32665 5943 32695 5975
rect 32749 5943 32779 5975
rect 32833 5943 32863 5975
rect 32917 5943 32947 5975
rect 32085 5907 32124 5937
rect 32094 5871 32124 5907
rect 33296 5922 33326 5975
rect 33368 6010 33443 6020
rect 33368 5976 33384 6010
rect 33418 5976 33443 6010
rect 33368 5966 33443 5976
rect 33601 5973 33631 6109
rect 33713 6093 33743 6121
rect 33693 6083 33759 6093
rect 33693 6049 33709 6083
rect 33743 6049 33759 6083
rect 33693 6039 33759 6049
rect 33812 5997 33842 6121
rect 33911 6081 33941 6109
rect 33296 5892 33359 5922
rect 33329 5877 33359 5892
rect 33413 5877 33443 5966
rect 33536 5957 33631 5973
rect 33536 5923 33546 5957
rect 33580 5923 33631 5957
rect 33673 5987 33842 5997
rect 33673 5953 33689 5987
rect 33723 5967 33842 5987
rect 33884 6071 33958 6081
rect 33884 6037 33908 6071
rect 33942 6037 33958 6071
rect 34131 6099 34161 6121
rect 34131 6083 34195 6099
rect 34030 6050 34060 6065
rect 33884 6027 33958 6037
rect 33723 5953 33739 5967
rect 33673 5943 33739 5953
rect 33536 5907 33631 5923
rect 33601 5827 33631 5907
rect 33686 5827 33716 5943
rect 33781 5909 33842 5925
rect 33781 5875 33798 5909
rect 33832 5875 33842 5909
rect 33781 5859 33842 5875
rect 33781 5827 33811 5859
rect 33884 5827 33914 6027
rect 34016 6020 34060 6050
rect 34131 6049 34151 6083
rect 34185 6049 34195 6083
rect 34131 6033 34195 6049
rect 34016 5985 34046 6020
rect 34237 5991 34267 6121
rect 33956 5975 34046 5985
rect 33956 5941 33972 5975
rect 34006 5941 34046 5975
rect 33956 5931 34046 5941
rect 34016 5893 34046 5931
rect 34098 5975 34267 5991
rect 34098 5941 34108 5975
rect 34142 5961 34267 5975
rect 34142 5941 34152 5961
rect 34098 5925 34152 5941
rect 34332 5925 34362 6109
rect 34794 6094 34824 6109
rect 34783 6070 34824 6094
rect 34522 6041 34552 6063
rect 34606 6041 34636 6063
rect 34783 6041 34813 6070
rect 34889 6041 34919 6063
rect 35118 6041 35148 6063
rect 35363 6041 35393 6063
rect 35447 6041 35477 6063
rect 35531 6041 35561 6063
rect 35615 6041 35645 6063
rect 34410 6025 34552 6041
rect 34410 5991 34420 6025
rect 34454 5991 34552 6025
rect 34410 5975 34552 5991
rect 34594 6025 34813 6041
rect 34594 5991 34604 6025
rect 34638 5991 34813 6025
rect 34594 5975 34813 5991
rect 34855 6025 34919 6041
rect 34855 5991 34865 6025
rect 34899 5991 34919 6025
rect 34855 5975 34919 5991
rect 35062 6025 35148 6041
rect 35062 5991 35078 6025
rect 35112 5991 35148 6025
rect 35062 5975 35148 5991
rect 35295 6025 35645 6041
rect 35295 5991 35311 6025
rect 35345 5991 35403 6025
rect 35437 5991 35487 6025
rect 35521 5991 35571 6025
rect 35605 5991 35645 6025
rect 35295 5975 35645 5991
rect 34520 5943 34550 5975
rect 34604 5943 34634 5975
rect 30903 5717 30933 5743
rect 30988 5717 31018 5743
rect 31083 5717 31113 5743
rect 31186 5717 31216 5743
rect 31318 5717 31348 5743
rect 31413 5717 31443 5743
rect 31497 5717 31527 5743
rect 31611 5717 31641 5743
rect 31822 5717 31852 5743
rect 31906 5717 31936 5743
rect 32094 5717 32124 5743
rect 32191 5717 32221 5743
rect 32420 5717 32450 5743
rect 32665 5717 32695 5743
rect 32749 5717 32779 5743
rect 32833 5717 32863 5743
rect 32917 5717 32947 5743
rect 33329 5723 33359 5749
rect 33413 5723 33443 5749
rect 34111 5827 34141 5925
rect 34194 5909 34260 5919
rect 34194 5875 34210 5909
rect 34244 5875 34260 5909
rect 34194 5865 34260 5875
rect 34309 5909 34390 5925
rect 34309 5875 34346 5909
rect 34380 5875 34390 5909
rect 34195 5827 34225 5865
rect 34309 5859 34390 5875
rect 34309 5827 34339 5859
rect 34783 5937 34813 5975
rect 34889 5943 34919 5975
rect 35118 5943 35148 5975
rect 35363 5943 35393 5975
rect 35447 5943 35477 5975
rect 35531 5943 35561 5975
rect 35615 5943 35645 5975
rect 34783 5907 34822 5937
rect 34792 5871 34822 5907
rect 33601 5717 33631 5743
rect 33686 5717 33716 5743
rect 33781 5717 33811 5743
rect 33884 5717 33914 5743
rect 34016 5717 34046 5743
rect 34111 5717 34141 5743
rect 34195 5717 34225 5743
rect 34309 5717 34339 5743
rect 34520 5717 34550 5743
rect 34604 5717 34634 5743
rect 34792 5717 34822 5743
rect 34889 5717 34919 5743
rect 35118 5717 35148 5743
rect 35363 5717 35393 5743
rect 35447 5717 35477 5743
rect 35531 5717 35561 5743
rect 35615 5717 35645 5743
rect 9458 3025 9710 3041
rect 9458 3008 9474 3025
rect 9384 2991 9474 3008
rect 9694 3008 9710 3025
rect 9916 3025 10168 3041
rect 9916 3008 9932 3025
rect 9694 2991 9784 3008
rect 9384 2944 9784 2991
rect 9842 2991 9932 3008
rect 10152 3008 10168 3025
rect 10374 3025 10626 3041
rect 10374 3008 10390 3025
rect 10152 2991 10242 3008
rect 9842 2944 10242 2991
rect 10300 2991 10390 3008
rect 10610 3008 10626 3025
rect 10832 3025 11084 3041
rect 10832 3008 10848 3025
rect 10610 2991 10700 3008
rect 10300 2944 10700 2991
rect 10758 2991 10848 3008
rect 11068 3008 11084 3025
rect 11290 3025 11542 3041
rect 11290 3008 11306 3025
rect 11068 2991 11158 3008
rect 10758 2944 11158 2991
rect 11216 2991 11306 3008
rect 11526 3008 11542 3025
rect 11748 3025 12000 3041
rect 11748 3008 11764 3025
rect 11526 2991 11616 3008
rect 11216 2944 11616 2991
rect 11674 2991 11764 3008
rect 11984 3008 12000 3025
rect 12206 3025 12458 3041
rect 12206 3008 12222 3025
rect 11984 2991 12074 3008
rect 11674 2944 12074 2991
rect 12132 2991 12222 3008
rect 12442 3008 12458 3025
rect 12664 3025 12916 3041
rect 12664 3008 12680 3025
rect 12442 2991 12532 3008
rect 12132 2944 12532 2991
rect 12590 2991 12680 3008
rect 12900 3008 12916 3025
rect 13122 3025 13374 3041
rect 13122 3008 13138 3025
rect 12900 2991 12990 3008
rect 12590 2944 12990 2991
rect 13048 2991 13138 3008
rect 13358 3008 13374 3025
rect 13580 3025 13832 3041
rect 13580 3008 13596 3025
rect 13358 2991 13448 3008
rect 13048 2944 13448 2991
rect 13506 2991 13596 3008
rect 13816 3008 13832 3025
rect 14038 3025 14290 3041
rect 14038 3008 14054 3025
rect 13816 2991 13906 3008
rect 13506 2944 13906 2991
rect 13964 2991 14054 3008
rect 14274 3008 14290 3025
rect 14496 3025 14748 3041
rect 14496 3008 14512 3025
rect 14274 2991 14364 3008
rect 13964 2944 14364 2991
rect 14422 2991 14512 3008
rect 14732 3008 14748 3025
rect 14954 3025 15206 3041
rect 14954 3008 14970 3025
rect 14732 2991 14822 3008
rect 14422 2944 14822 2991
rect 14880 2991 14970 3008
rect 15190 3008 15206 3025
rect 15412 3025 15664 3041
rect 15412 3008 15428 3025
rect 15190 2991 15280 3008
rect 14880 2944 15280 2991
rect 15338 2991 15428 3008
rect 15648 3008 15664 3025
rect 15870 3025 16122 3041
rect 15870 3008 15886 3025
rect 15648 2991 15738 3008
rect 15338 2944 15738 2991
rect 15796 2991 15886 3008
rect 16106 3008 16122 3025
rect 16328 3025 16580 3041
rect 16328 3008 16344 3025
rect 16106 2991 16196 3008
rect 15796 2944 16196 2991
rect 16254 2991 16344 3008
rect 16564 3008 16580 3025
rect 16786 3025 17038 3041
rect 16786 3008 16802 3025
rect 16564 2991 16654 3008
rect 16254 2944 16654 2991
rect 16712 2991 16802 3008
rect 17022 3008 17038 3025
rect 17244 3025 17496 3041
rect 17244 3008 17260 3025
rect 17022 2991 17112 3008
rect 16712 2944 17112 2991
rect 17170 2991 17260 3008
rect 17480 3008 17496 3025
rect 17480 2991 17570 3008
rect 17170 2944 17570 2991
rect 9384 1297 9784 1344
rect 9384 1280 9474 1297
rect 9458 1263 9474 1280
rect 9694 1280 9784 1297
rect 9842 1297 10242 1344
rect 9842 1280 9932 1297
rect 9694 1263 9710 1280
rect 9458 1247 9710 1263
rect 9916 1263 9932 1280
rect 10152 1280 10242 1297
rect 10300 1297 10700 1344
rect 10300 1280 10390 1297
rect 10152 1263 10168 1280
rect 9916 1247 10168 1263
rect 10374 1263 10390 1280
rect 10610 1280 10700 1297
rect 10758 1297 11158 1344
rect 10758 1280 10848 1297
rect 10610 1263 10626 1280
rect 10374 1247 10626 1263
rect 10832 1263 10848 1280
rect 11068 1280 11158 1297
rect 11216 1297 11616 1344
rect 11216 1280 11306 1297
rect 11068 1263 11084 1280
rect 10832 1247 11084 1263
rect 11290 1263 11306 1280
rect 11526 1280 11616 1297
rect 11674 1297 12074 1344
rect 11674 1280 11764 1297
rect 11526 1263 11542 1280
rect 11290 1247 11542 1263
rect 11748 1263 11764 1280
rect 11984 1280 12074 1297
rect 12132 1297 12532 1344
rect 12132 1280 12222 1297
rect 11984 1263 12000 1280
rect 11748 1247 12000 1263
rect 12206 1263 12222 1280
rect 12442 1280 12532 1297
rect 12590 1297 12990 1344
rect 12590 1280 12680 1297
rect 12442 1263 12458 1280
rect 12206 1247 12458 1263
rect 12664 1263 12680 1280
rect 12900 1280 12990 1297
rect 13048 1297 13448 1344
rect 13048 1280 13138 1297
rect 12900 1263 12916 1280
rect 12664 1247 12916 1263
rect 13122 1263 13138 1280
rect 13358 1280 13448 1297
rect 13506 1297 13906 1344
rect 13506 1280 13596 1297
rect 13358 1263 13374 1280
rect 13122 1247 13374 1263
rect 13580 1263 13596 1280
rect 13816 1280 13906 1297
rect 13964 1297 14364 1344
rect 13964 1280 14054 1297
rect 13816 1263 13832 1280
rect 13580 1247 13832 1263
rect 14038 1263 14054 1280
rect 14274 1280 14364 1297
rect 14422 1297 14822 1344
rect 14422 1280 14512 1297
rect 14274 1263 14290 1280
rect 14038 1247 14290 1263
rect 14496 1263 14512 1280
rect 14732 1280 14822 1297
rect 14880 1297 15280 1344
rect 14880 1280 14970 1297
rect 14732 1263 14748 1280
rect 14496 1247 14748 1263
rect 14954 1263 14970 1280
rect 15190 1280 15280 1297
rect 15338 1297 15738 1344
rect 15338 1280 15428 1297
rect 15190 1263 15206 1280
rect 14954 1247 15206 1263
rect 15412 1263 15428 1280
rect 15648 1280 15738 1297
rect 15796 1297 16196 1344
rect 15796 1280 15886 1297
rect 15648 1263 15664 1280
rect 15412 1247 15664 1263
rect 15870 1263 15886 1280
rect 16106 1280 16196 1297
rect 16254 1297 16654 1344
rect 16254 1280 16344 1297
rect 16106 1263 16122 1280
rect 15870 1247 16122 1263
rect 16328 1263 16344 1280
rect 16564 1280 16654 1297
rect 16712 1297 17112 1344
rect 16712 1280 16802 1297
rect 16564 1263 16580 1280
rect 16328 1247 16580 1263
rect 16786 1263 16802 1280
rect 17022 1280 17112 1297
rect 17170 1297 17570 1344
rect 17170 1280 17260 1297
rect 17022 1263 17038 1280
rect 16786 1247 17038 1263
rect 17244 1263 17260 1280
rect 17480 1280 17570 1297
rect 17480 1263 17496 1280
rect 17244 1247 17496 1263
rect 8899 360 9151 376
rect 8899 343 8915 360
rect 8825 326 8915 343
rect 9135 343 9151 360
rect 9357 360 9609 376
rect 9357 343 9373 360
rect 9135 326 9225 343
rect 8825 279 9225 326
rect 9283 326 9373 343
rect 9593 343 9609 360
rect 9815 360 10067 376
rect 9815 343 9831 360
rect 9593 326 9683 343
rect 9283 279 9683 326
rect 9741 326 9831 343
rect 10051 343 10067 360
rect 10273 360 10525 376
rect 10273 343 10289 360
rect 10051 326 10141 343
rect 9741 279 10141 326
rect 10199 326 10289 343
rect 10509 343 10525 360
rect 10731 360 10983 376
rect 10731 343 10747 360
rect 10509 326 10599 343
rect 10199 279 10599 326
rect 10657 326 10747 343
rect 10967 343 10983 360
rect 11189 360 11441 376
rect 11189 343 11205 360
rect 10967 326 11057 343
rect 10657 279 11057 326
rect 11115 326 11205 343
rect 11425 343 11441 360
rect 11647 360 11899 376
rect 11647 343 11663 360
rect 11425 326 11515 343
rect 11115 279 11515 326
rect 11573 326 11663 343
rect 11883 343 11899 360
rect 12105 360 12357 376
rect 12105 343 12121 360
rect 11883 326 11973 343
rect 11573 279 11973 326
rect 12031 326 12121 343
rect 12341 343 12357 360
rect 12563 360 12815 376
rect 12563 343 12579 360
rect 12341 326 12431 343
rect 12031 279 12431 326
rect 12489 326 12579 343
rect 12799 343 12815 360
rect 13021 360 13273 376
rect 13021 343 13037 360
rect 12799 326 12889 343
rect 12489 279 12889 326
rect 12947 326 13037 343
rect 13257 343 13273 360
rect 13899 360 14151 376
rect 13899 343 13915 360
rect 13257 326 13347 343
rect 12947 279 13347 326
rect 13825 326 13915 343
rect 14135 343 14151 360
rect 14357 360 14609 376
rect 14357 343 14373 360
rect 14135 326 14225 343
rect 13825 279 14225 326
rect 14283 326 14373 343
rect 14593 343 14609 360
rect 14815 360 15067 376
rect 14815 343 14831 360
rect 14593 326 14683 343
rect 14283 279 14683 326
rect 14741 326 14831 343
rect 15051 343 15067 360
rect 15273 360 15525 376
rect 15273 343 15289 360
rect 15051 326 15141 343
rect 14741 279 15141 326
rect 15199 326 15289 343
rect 15509 343 15525 360
rect 15731 360 15983 376
rect 15731 343 15747 360
rect 15509 326 15599 343
rect 15199 279 15599 326
rect 15657 326 15747 343
rect 15967 343 15983 360
rect 16189 360 16441 376
rect 16189 343 16205 360
rect 15967 326 16057 343
rect 15657 279 16057 326
rect 16115 326 16205 343
rect 16425 343 16441 360
rect 16647 360 16899 376
rect 16647 343 16663 360
rect 16425 326 16515 343
rect 16115 279 16515 326
rect 16573 326 16663 343
rect 16883 343 16899 360
rect 17105 360 17357 376
rect 17105 343 17121 360
rect 16883 326 16973 343
rect 16573 279 16973 326
rect 17031 326 17121 343
rect 17341 343 17357 360
rect 17563 360 17815 376
rect 17563 343 17579 360
rect 17341 326 17431 343
rect 17031 279 17431 326
rect 17489 326 17579 343
rect 17799 343 17815 360
rect 18021 360 18273 376
rect 18021 343 18037 360
rect 17799 326 17889 343
rect 17489 279 17889 326
rect 17947 326 18037 343
rect 18257 343 18273 360
rect 18257 326 18347 343
rect 17947 279 18347 326
rect 8825 -968 9225 -921
rect 8825 -985 8915 -968
rect 8899 -1002 8915 -985
rect 9135 -985 9225 -968
rect 9283 -968 9683 -921
rect 9283 -985 9373 -968
rect 9135 -1002 9151 -985
rect 8899 -1018 9151 -1002
rect 9357 -1002 9373 -985
rect 9593 -985 9683 -968
rect 9741 -968 10141 -921
rect 9741 -985 9831 -968
rect 9593 -1002 9609 -985
rect 9357 -1018 9609 -1002
rect 9815 -1002 9831 -985
rect 10051 -985 10141 -968
rect 10199 -968 10599 -921
rect 10199 -985 10289 -968
rect 10051 -1002 10067 -985
rect 9815 -1018 10067 -1002
rect 10273 -1002 10289 -985
rect 10509 -985 10599 -968
rect 10657 -968 11057 -921
rect 10657 -985 10747 -968
rect 10509 -1002 10525 -985
rect 10273 -1018 10525 -1002
rect 10731 -1002 10747 -985
rect 10967 -985 11057 -968
rect 11115 -968 11515 -921
rect 11115 -985 11205 -968
rect 10967 -1002 10983 -985
rect 10731 -1018 10983 -1002
rect 11189 -1002 11205 -985
rect 11425 -985 11515 -968
rect 11573 -968 11973 -921
rect 11573 -985 11663 -968
rect 11425 -1002 11441 -985
rect 11189 -1018 11441 -1002
rect 11647 -1002 11663 -985
rect 11883 -985 11973 -968
rect 12031 -968 12431 -921
rect 12031 -985 12121 -968
rect 11883 -1002 11899 -985
rect 11647 -1018 11899 -1002
rect 12105 -1002 12121 -985
rect 12341 -985 12431 -968
rect 12489 -968 12889 -921
rect 12489 -985 12579 -968
rect 12341 -1002 12357 -985
rect 12105 -1018 12357 -1002
rect 12563 -1002 12579 -985
rect 12799 -985 12889 -968
rect 12947 -968 13347 -921
rect 12947 -985 13037 -968
rect 12799 -1002 12815 -985
rect 12563 -1018 12815 -1002
rect 13021 -1002 13037 -985
rect 13257 -985 13347 -968
rect 13825 -968 14225 -921
rect 13825 -985 13915 -968
rect 13257 -1002 13273 -985
rect 13021 -1018 13273 -1002
rect 13899 -1002 13915 -985
rect 14135 -985 14225 -968
rect 14283 -968 14683 -921
rect 14283 -985 14373 -968
rect 14135 -1002 14151 -985
rect 13899 -1018 14151 -1002
rect 14357 -1002 14373 -985
rect 14593 -985 14683 -968
rect 14741 -968 15141 -921
rect 14741 -985 14831 -968
rect 14593 -1002 14609 -985
rect 14357 -1018 14609 -1002
rect 14815 -1002 14831 -985
rect 15051 -985 15141 -968
rect 15199 -968 15599 -921
rect 15199 -985 15289 -968
rect 15051 -1002 15067 -985
rect 14815 -1018 15067 -1002
rect 15273 -1002 15289 -985
rect 15509 -985 15599 -968
rect 15657 -968 16057 -921
rect 15657 -985 15747 -968
rect 15509 -1002 15525 -985
rect 15273 -1018 15525 -1002
rect 15731 -1002 15747 -985
rect 15967 -985 16057 -968
rect 16115 -968 16515 -921
rect 16115 -985 16205 -968
rect 15967 -1002 15983 -985
rect 15731 -1018 15983 -1002
rect 16189 -1002 16205 -985
rect 16425 -985 16515 -968
rect 16573 -968 16973 -921
rect 16573 -985 16663 -968
rect 16425 -1002 16441 -985
rect 16189 -1018 16441 -1002
rect 16647 -1002 16663 -985
rect 16883 -985 16973 -968
rect 17031 -968 17431 -921
rect 17031 -985 17121 -968
rect 16883 -1002 16899 -985
rect 16647 -1018 16899 -1002
rect 17105 -1002 17121 -985
rect 17341 -985 17431 -968
rect 17489 -968 17889 -921
rect 17489 -985 17579 -968
rect 17341 -1002 17357 -985
rect 17105 -1018 17357 -1002
rect 17563 -1002 17579 -985
rect 17799 -985 17889 -968
rect 17947 -968 18347 -921
rect 17947 -985 18037 -968
rect 17799 -1002 17815 -985
rect 17563 -1018 17815 -1002
rect 18021 -1002 18037 -985
rect 18257 -985 18347 -968
rect 18257 -1002 18273 -985
rect 18021 -1018 18273 -1002
rect 24458 3025 24710 3041
rect 24458 3008 24474 3025
rect 24384 2991 24474 3008
rect 24694 3008 24710 3025
rect 24916 3025 25168 3041
rect 24916 3008 24932 3025
rect 24694 2991 24784 3008
rect 24384 2944 24784 2991
rect 24842 2991 24932 3008
rect 25152 3008 25168 3025
rect 25374 3025 25626 3041
rect 25374 3008 25390 3025
rect 25152 2991 25242 3008
rect 24842 2944 25242 2991
rect 25300 2991 25390 3008
rect 25610 3008 25626 3025
rect 25832 3025 26084 3041
rect 25832 3008 25848 3025
rect 25610 2991 25700 3008
rect 25300 2944 25700 2991
rect 25758 2991 25848 3008
rect 26068 3008 26084 3025
rect 26290 3025 26542 3041
rect 26290 3008 26306 3025
rect 26068 2991 26158 3008
rect 25758 2944 26158 2991
rect 26216 2991 26306 3008
rect 26526 3008 26542 3025
rect 26748 3025 27000 3041
rect 26748 3008 26764 3025
rect 26526 2991 26616 3008
rect 26216 2944 26616 2991
rect 26674 2991 26764 3008
rect 26984 3008 27000 3025
rect 27206 3025 27458 3041
rect 27206 3008 27222 3025
rect 26984 2991 27074 3008
rect 26674 2944 27074 2991
rect 27132 2991 27222 3008
rect 27442 3008 27458 3025
rect 27664 3025 27916 3041
rect 27664 3008 27680 3025
rect 27442 2991 27532 3008
rect 27132 2944 27532 2991
rect 27590 2991 27680 3008
rect 27900 3008 27916 3025
rect 28122 3025 28374 3041
rect 28122 3008 28138 3025
rect 27900 2991 27990 3008
rect 27590 2944 27990 2991
rect 28048 2991 28138 3008
rect 28358 3008 28374 3025
rect 28580 3025 28832 3041
rect 28580 3008 28596 3025
rect 28358 2991 28448 3008
rect 28048 2944 28448 2991
rect 28506 2991 28596 3008
rect 28816 3008 28832 3025
rect 29038 3025 29290 3041
rect 29038 3008 29054 3025
rect 28816 2991 28906 3008
rect 28506 2944 28906 2991
rect 28964 2991 29054 3008
rect 29274 3008 29290 3025
rect 29496 3025 29748 3041
rect 29496 3008 29512 3025
rect 29274 2991 29364 3008
rect 28964 2944 29364 2991
rect 29422 2991 29512 3008
rect 29732 3008 29748 3025
rect 29954 3025 30206 3041
rect 29954 3008 29970 3025
rect 29732 2991 29822 3008
rect 29422 2944 29822 2991
rect 29880 2991 29970 3008
rect 30190 3008 30206 3025
rect 30412 3025 30664 3041
rect 30412 3008 30428 3025
rect 30190 2991 30280 3008
rect 29880 2944 30280 2991
rect 30338 2991 30428 3008
rect 30648 3008 30664 3025
rect 30870 3025 31122 3041
rect 30870 3008 30886 3025
rect 30648 2991 30738 3008
rect 30338 2944 30738 2991
rect 30796 2991 30886 3008
rect 31106 3008 31122 3025
rect 31328 3025 31580 3041
rect 31328 3008 31344 3025
rect 31106 2991 31196 3008
rect 30796 2944 31196 2991
rect 31254 2991 31344 3008
rect 31564 3008 31580 3025
rect 31786 3025 32038 3041
rect 31786 3008 31802 3025
rect 31564 2991 31654 3008
rect 31254 2944 31654 2991
rect 31712 2991 31802 3008
rect 32022 3008 32038 3025
rect 32244 3025 32496 3041
rect 32244 3008 32260 3025
rect 32022 2991 32112 3008
rect 31712 2944 32112 2991
rect 32170 2991 32260 3008
rect 32480 3008 32496 3025
rect 32480 2991 32570 3008
rect 32170 2944 32570 2991
rect 24384 1297 24784 1344
rect 24384 1280 24474 1297
rect 24458 1263 24474 1280
rect 24694 1280 24784 1297
rect 24842 1297 25242 1344
rect 24842 1280 24932 1297
rect 24694 1263 24710 1280
rect 24458 1247 24710 1263
rect 24916 1263 24932 1280
rect 25152 1280 25242 1297
rect 25300 1297 25700 1344
rect 25300 1280 25390 1297
rect 25152 1263 25168 1280
rect 24916 1247 25168 1263
rect 25374 1263 25390 1280
rect 25610 1280 25700 1297
rect 25758 1297 26158 1344
rect 25758 1280 25848 1297
rect 25610 1263 25626 1280
rect 25374 1247 25626 1263
rect 25832 1263 25848 1280
rect 26068 1280 26158 1297
rect 26216 1297 26616 1344
rect 26216 1280 26306 1297
rect 26068 1263 26084 1280
rect 25832 1247 26084 1263
rect 26290 1263 26306 1280
rect 26526 1280 26616 1297
rect 26674 1297 27074 1344
rect 26674 1280 26764 1297
rect 26526 1263 26542 1280
rect 26290 1247 26542 1263
rect 26748 1263 26764 1280
rect 26984 1280 27074 1297
rect 27132 1297 27532 1344
rect 27132 1280 27222 1297
rect 26984 1263 27000 1280
rect 26748 1247 27000 1263
rect 27206 1263 27222 1280
rect 27442 1280 27532 1297
rect 27590 1297 27990 1344
rect 27590 1280 27680 1297
rect 27442 1263 27458 1280
rect 27206 1247 27458 1263
rect 27664 1263 27680 1280
rect 27900 1280 27990 1297
rect 28048 1297 28448 1344
rect 28048 1280 28138 1297
rect 27900 1263 27916 1280
rect 27664 1247 27916 1263
rect 28122 1263 28138 1280
rect 28358 1280 28448 1297
rect 28506 1297 28906 1344
rect 28506 1280 28596 1297
rect 28358 1263 28374 1280
rect 28122 1247 28374 1263
rect 28580 1263 28596 1280
rect 28816 1280 28906 1297
rect 28964 1297 29364 1344
rect 28964 1280 29054 1297
rect 28816 1263 28832 1280
rect 28580 1247 28832 1263
rect 29038 1263 29054 1280
rect 29274 1280 29364 1297
rect 29422 1297 29822 1344
rect 29422 1280 29512 1297
rect 29274 1263 29290 1280
rect 29038 1247 29290 1263
rect 29496 1263 29512 1280
rect 29732 1280 29822 1297
rect 29880 1297 30280 1344
rect 29880 1280 29970 1297
rect 29732 1263 29748 1280
rect 29496 1247 29748 1263
rect 29954 1263 29970 1280
rect 30190 1280 30280 1297
rect 30338 1297 30738 1344
rect 30338 1280 30428 1297
rect 30190 1263 30206 1280
rect 29954 1247 30206 1263
rect 30412 1263 30428 1280
rect 30648 1280 30738 1297
rect 30796 1297 31196 1344
rect 30796 1280 30886 1297
rect 30648 1263 30664 1280
rect 30412 1247 30664 1263
rect 30870 1263 30886 1280
rect 31106 1280 31196 1297
rect 31254 1297 31654 1344
rect 31254 1280 31344 1297
rect 31106 1263 31122 1280
rect 30870 1247 31122 1263
rect 31328 1263 31344 1280
rect 31564 1280 31654 1297
rect 31712 1297 32112 1344
rect 31712 1280 31802 1297
rect 31564 1263 31580 1280
rect 31328 1247 31580 1263
rect 31786 1263 31802 1280
rect 32022 1280 32112 1297
rect 32170 1297 32570 1344
rect 32170 1280 32260 1297
rect 32022 1263 32038 1280
rect 31786 1247 32038 1263
rect 32244 1263 32260 1280
rect 32480 1280 32570 1297
rect 32480 1263 32496 1280
rect 32244 1247 32496 1263
rect 23899 360 24151 376
rect 23899 343 23915 360
rect 23825 326 23915 343
rect 24135 343 24151 360
rect 24357 360 24609 376
rect 24357 343 24373 360
rect 24135 326 24225 343
rect 23825 279 24225 326
rect 24283 326 24373 343
rect 24593 343 24609 360
rect 24815 360 25067 376
rect 24815 343 24831 360
rect 24593 326 24683 343
rect 24283 279 24683 326
rect 24741 326 24831 343
rect 25051 343 25067 360
rect 25273 360 25525 376
rect 25273 343 25289 360
rect 25051 326 25141 343
rect 24741 279 25141 326
rect 25199 326 25289 343
rect 25509 343 25525 360
rect 25731 360 25983 376
rect 25731 343 25747 360
rect 25509 326 25599 343
rect 25199 279 25599 326
rect 25657 326 25747 343
rect 25967 343 25983 360
rect 26189 360 26441 376
rect 26189 343 26205 360
rect 25967 326 26057 343
rect 25657 279 26057 326
rect 26115 326 26205 343
rect 26425 343 26441 360
rect 26647 360 26899 376
rect 26647 343 26663 360
rect 26425 326 26515 343
rect 26115 279 26515 326
rect 26573 326 26663 343
rect 26883 343 26899 360
rect 27105 360 27357 376
rect 27105 343 27121 360
rect 26883 326 26973 343
rect 26573 279 26973 326
rect 27031 326 27121 343
rect 27341 343 27357 360
rect 27563 360 27815 376
rect 27563 343 27579 360
rect 27341 326 27431 343
rect 27031 279 27431 326
rect 27489 326 27579 343
rect 27799 343 27815 360
rect 28021 360 28273 376
rect 28021 343 28037 360
rect 27799 326 27889 343
rect 27489 279 27889 326
rect 27947 326 28037 343
rect 28257 343 28273 360
rect 28899 360 29151 376
rect 28899 343 28915 360
rect 28257 326 28347 343
rect 27947 279 28347 326
rect 28825 326 28915 343
rect 29135 343 29151 360
rect 29357 360 29609 376
rect 29357 343 29373 360
rect 29135 326 29225 343
rect 28825 279 29225 326
rect 29283 326 29373 343
rect 29593 343 29609 360
rect 29815 360 30067 376
rect 29815 343 29831 360
rect 29593 326 29683 343
rect 29283 279 29683 326
rect 29741 326 29831 343
rect 30051 343 30067 360
rect 30273 360 30525 376
rect 30273 343 30289 360
rect 30051 326 30141 343
rect 29741 279 30141 326
rect 30199 326 30289 343
rect 30509 343 30525 360
rect 30731 360 30983 376
rect 30731 343 30747 360
rect 30509 326 30599 343
rect 30199 279 30599 326
rect 30657 326 30747 343
rect 30967 343 30983 360
rect 31189 360 31441 376
rect 31189 343 31205 360
rect 30967 326 31057 343
rect 30657 279 31057 326
rect 31115 326 31205 343
rect 31425 343 31441 360
rect 31647 360 31899 376
rect 31647 343 31663 360
rect 31425 326 31515 343
rect 31115 279 31515 326
rect 31573 326 31663 343
rect 31883 343 31899 360
rect 32105 360 32357 376
rect 32105 343 32121 360
rect 31883 326 31973 343
rect 31573 279 31973 326
rect 32031 326 32121 343
rect 32341 343 32357 360
rect 32563 360 32815 376
rect 32563 343 32579 360
rect 32341 326 32431 343
rect 32031 279 32431 326
rect 32489 326 32579 343
rect 32799 343 32815 360
rect 33021 360 33273 376
rect 33021 343 33037 360
rect 32799 326 32889 343
rect 32489 279 32889 326
rect 32947 326 33037 343
rect 33257 343 33273 360
rect 33257 326 33347 343
rect 32947 279 33347 326
rect 23825 -968 24225 -921
rect 23825 -985 23915 -968
rect 23899 -1002 23915 -985
rect 24135 -985 24225 -968
rect 24283 -968 24683 -921
rect 24283 -985 24373 -968
rect 24135 -1002 24151 -985
rect 23899 -1018 24151 -1002
rect 24357 -1002 24373 -985
rect 24593 -985 24683 -968
rect 24741 -968 25141 -921
rect 24741 -985 24831 -968
rect 24593 -1002 24609 -985
rect 24357 -1018 24609 -1002
rect 24815 -1002 24831 -985
rect 25051 -985 25141 -968
rect 25199 -968 25599 -921
rect 25199 -985 25289 -968
rect 25051 -1002 25067 -985
rect 24815 -1018 25067 -1002
rect 25273 -1002 25289 -985
rect 25509 -985 25599 -968
rect 25657 -968 26057 -921
rect 25657 -985 25747 -968
rect 25509 -1002 25525 -985
rect 25273 -1018 25525 -1002
rect 25731 -1002 25747 -985
rect 25967 -985 26057 -968
rect 26115 -968 26515 -921
rect 26115 -985 26205 -968
rect 25967 -1002 25983 -985
rect 25731 -1018 25983 -1002
rect 26189 -1002 26205 -985
rect 26425 -985 26515 -968
rect 26573 -968 26973 -921
rect 26573 -985 26663 -968
rect 26425 -1002 26441 -985
rect 26189 -1018 26441 -1002
rect 26647 -1002 26663 -985
rect 26883 -985 26973 -968
rect 27031 -968 27431 -921
rect 27031 -985 27121 -968
rect 26883 -1002 26899 -985
rect 26647 -1018 26899 -1002
rect 27105 -1002 27121 -985
rect 27341 -985 27431 -968
rect 27489 -968 27889 -921
rect 27489 -985 27579 -968
rect 27341 -1002 27357 -985
rect 27105 -1018 27357 -1002
rect 27563 -1002 27579 -985
rect 27799 -985 27889 -968
rect 27947 -968 28347 -921
rect 27947 -985 28037 -968
rect 27799 -1002 27815 -985
rect 27563 -1018 27815 -1002
rect 28021 -1002 28037 -985
rect 28257 -985 28347 -968
rect 28825 -968 29225 -921
rect 28825 -985 28915 -968
rect 28257 -1002 28273 -985
rect 28021 -1018 28273 -1002
rect 28899 -1002 28915 -985
rect 29135 -985 29225 -968
rect 29283 -968 29683 -921
rect 29283 -985 29373 -968
rect 29135 -1002 29151 -985
rect 28899 -1018 29151 -1002
rect 29357 -1002 29373 -985
rect 29593 -985 29683 -968
rect 29741 -968 30141 -921
rect 29741 -985 29831 -968
rect 29593 -1002 29609 -985
rect 29357 -1018 29609 -1002
rect 29815 -1002 29831 -985
rect 30051 -985 30141 -968
rect 30199 -968 30599 -921
rect 30199 -985 30289 -968
rect 30051 -1002 30067 -985
rect 29815 -1018 30067 -1002
rect 30273 -1002 30289 -985
rect 30509 -985 30599 -968
rect 30657 -968 31057 -921
rect 30657 -985 30747 -968
rect 30509 -1002 30525 -985
rect 30273 -1018 30525 -1002
rect 30731 -1002 30747 -985
rect 30967 -985 31057 -968
rect 31115 -968 31515 -921
rect 31115 -985 31205 -968
rect 30967 -1002 30983 -985
rect 30731 -1018 30983 -1002
rect 31189 -1002 31205 -985
rect 31425 -985 31515 -968
rect 31573 -968 31973 -921
rect 31573 -985 31663 -968
rect 31425 -1002 31441 -985
rect 31189 -1018 31441 -1002
rect 31647 -1002 31663 -985
rect 31883 -985 31973 -968
rect 32031 -968 32431 -921
rect 32031 -985 32121 -968
rect 31883 -1002 31899 -985
rect 31647 -1018 31899 -1002
rect 32105 -1002 32121 -985
rect 32341 -985 32431 -968
rect 32489 -968 32889 -921
rect 32489 -985 32579 -968
rect 32341 -1002 32357 -985
rect 32105 -1018 32357 -1002
rect 32563 -1002 32579 -985
rect 32799 -985 32889 -968
rect 32947 -968 33347 -921
rect 32947 -985 33037 -968
rect 32799 -1002 32815 -985
rect 32563 -1018 32815 -1002
rect 33021 -1002 33037 -985
rect 33257 -985 33347 -968
rect 33257 -1002 33273 -985
rect 33021 -1018 33273 -1002
rect 8898 -2142 9150 -2126
rect 8898 -2159 8914 -2142
rect 8824 -2176 8914 -2159
rect 9134 -2159 9150 -2142
rect 9356 -2142 9608 -2126
rect 9356 -2159 9372 -2142
rect 9134 -2176 9224 -2159
rect 8824 -2214 9224 -2176
rect 9282 -2176 9372 -2159
rect 9592 -2159 9608 -2142
rect 9814 -2142 10066 -2126
rect 9814 -2159 9830 -2142
rect 9592 -2176 9682 -2159
rect 9282 -2214 9682 -2176
rect 9740 -2176 9830 -2159
rect 10050 -2159 10066 -2142
rect 10272 -2142 10524 -2126
rect 10272 -2159 10288 -2142
rect 10050 -2176 10140 -2159
rect 9740 -2214 10140 -2176
rect 10198 -2176 10288 -2159
rect 10508 -2159 10524 -2142
rect 10730 -2142 10982 -2126
rect 10730 -2159 10746 -2142
rect 10508 -2176 10598 -2159
rect 10198 -2214 10598 -2176
rect 10656 -2176 10746 -2159
rect 10966 -2159 10982 -2142
rect 11188 -2142 11440 -2126
rect 11188 -2159 11204 -2142
rect 10966 -2176 11056 -2159
rect 10656 -2214 11056 -2176
rect 11114 -2176 11204 -2159
rect 11424 -2159 11440 -2142
rect 11646 -2142 11898 -2126
rect 11646 -2159 11662 -2142
rect 11424 -2176 11514 -2159
rect 11114 -2214 11514 -2176
rect 11572 -2176 11662 -2159
rect 11882 -2159 11898 -2142
rect 12104 -2142 12356 -2126
rect 12104 -2159 12120 -2142
rect 11882 -2176 11972 -2159
rect 11572 -2214 11972 -2176
rect 12030 -2176 12120 -2159
rect 12340 -2159 12356 -2142
rect 12562 -2142 12814 -2126
rect 12562 -2159 12578 -2142
rect 12340 -2176 12430 -2159
rect 12030 -2214 12430 -2176
rect 12488 -2176 12578 -2159
rect 12798 -2159 12814 -2142
rect 13020 -2142 13272 -2126
rect 13020 -2159 13036 -2142
rect 12798 -2176 12888 -2159
rect 12488 -2214 12888 -2176
rect 12946 -2176 13036 -2159
rect 13256 -2159 13272 -2142
rect 13898 -2142 14150 -2126
rect 13898 -2159 13914 -2142
rect 13256 -2176 13346 -2159
rect 12946 -2214 13346 -2176
rect 13824 -2176 13914 -2159
rect 14134 -2159 14150 -2142
rect 14356 -2142 14608 -2126
rect 14356 -2159 14372 -2142
rect 14134 -2176 14224 -2159
rect 13824 -2214 14224 -2176
rect 14282 -2176 14372 -2159
rect 14592 -2159 14608 -2142
rect 14814 -2142 15066 -2126
rect 14814 -2159 14830 -2142
rect 14592 -2176 14682 -2159
rect 14282 -2214 14682 -2176
rect 14740 -2176 14830 -2159
rect 15050 -2159 15066 -2142
rect 15272 -2142 15524 -2126
rect 15272 -2159 15288 -2142
rect 15050 -2176 15140 -2159
rect 14740 -2214 15140 -2176
rect 15198 -2176 15288 -2159
rect 15508 -2159 15524 -2142
rect 15730 -2142 15982 -2126
rect 15730 -2159 15746 -2142
rect 15508 -2176 15598 -2159
rect 15198 -2214 15598 -2176
rect 15656 -2176 15746 -2159
rect 15966 -2159 15982 -2142
rect 16188 -2142 16440 -2126
rect 16188 -2159 16204 -2142
rect 15966 -2176 16056 -2159
rect 15656 -2214 16056 -2176
rect 16114 -2176 16204 -2159
rect 16424 -2159 16440 -2142
rect 16646 -2142 16898 -2126
rect 16646 -2159 16662 -2142
rect 16424 -2176 16514 -2159
rect 16114 -2214 16514 -2176
rect 16572 -2176 16662 -2159
rect 16882 -2159 16898 -2142
rect 17104 -2142 17356 -2126
rect 17104 -2159 17120 -2142
rect 16882 -2176 16972 -2159
rect 16572 -2214 16972 -2176
rect 17030 -2176 17120 -2159
rect 17340 -2159 17356 -2142
rect 17562 -2142 17814 -2126
rect 17562 -2159 17578 -2142
rect 17340 -2176 17430 -2159
rect 17030 -2214 17430 -2176
rect 17488 -2176 17578 -2159
rect 17798 -2159 17814 -2142
rect 18020 -2142 18272 -2126
rect 18020 -2159 18036 -2142
rect 17798 -2176 17888 -2159
rect 17488 -2214 17888 -2176
rect 17946 -2176 18036 -2159
rect 18256 -2159 18272 -2142
rect 18256 -2176 18346 -2159
rect 17946 -2214 18346 -2176
rect 8824 -2452 9224 -2414
rect 8824 -2469 8914 -2452
rect 8898 -2486 8914 -2469
rect 9134 -2469 9224 -2452
rect 9282 -2452 9682 -2414
rect 9282 -2469 9372 -2452
rect 9134 -2486 9150 -2469
rect 8898 -2502 9150 -2486
rect 9356 -2486 9372 -2469
rect 9592 -2469 9682 -2452
rect 9740 -2452 10140 -2414
rect 9740 -2469 9830 -2452
rect 9592 -2486 9608 -2469
rect 9356 -2502 9608 -2486
rect 9814 -2486 9830 -2469
rect 10050 -2469 10140 -2452
rect 10198 -2452 10598 -2414
rect 10198 -2469 10288 -2452
rect 10050 -2486 10066 -2469
rect 9814 -2502 10066 -2486
rect 10272 -2486 10288 -2469
rect 10508 -2469 10598 -2452
rect 10656 -2452 11056 -2414
rect 10656 -2469 10746 -2452
rect 10508 -2486 10524 -2469
rect 10272 -2502 10524 -2486
rect 10730 -2486 10746 -2469
rect 10966 -2469 11056 -2452
rect 11114 -2452 11514 -2414
rect 11114 -2469 11204 -2452
rect 10966 -2486 10982 -2469
rect 10730 -2502 10982 -2486
rect 11188 -2486 11204 -2469
rect 11424 -2469 11514 -2452
rect 11572 -2452 11972 -2414
rect 11572 -2469 11662 -2452
rect 11424 -2486 11440 -2469
rect 11188 -2502 11440 -2486
rect 11646 -2486 11662 -2469
rect 11882 -2469 11972 -2452
rect 12030 -2452 12430 -2414
rect 12030 -2469 12120 -2452
rect 11882 -2486 11898 -2469
rect 11646 -2502 11898 -2486
rect 12104 -2486 12120 -2469
rect 12340 -2469 12430 -2452
rect 12488 -2452 12888 -2414
rect 12488 -2469 12578 -2452
rect 12340 -2486 12356 -2469
rect 12104 -2502 12356 -2486
rect 12562 -2486 12578 -2469
rect 12798 -2469 12888 -2452
rect 12946 -2452 13346 -2414
rect 12946 -2469 13036 -2452
rect 12798 -2486 12814 -2469
rect 12562 -2502 12814 -2486
rect 13020 -2486 13036 -2469
rect 13256 -2469 13346 -2452
rect 13824 -2452 14224 -2414
rect 13824 -2469 13914 -2452
rect 13256 -2486 13272 -2469
rect 13020 -2502 13272 -2486
rect 13898 -2486 13914 -2469
rect 14134 -2469 14224 -2452
rect 14282 -2452 14682 -2414
rect 14282 -2469 14372 -2452
rect 14134 -2486 14150 -2469
rect 13898 -2502 14150 -2486
rect 14356 -2486 14372 -2469
rect 14592 -2469 14682 -2452
rect 14740 -2452 15140 -2414
rect 14740 -2469 14830 -2452
rect 14592 -2486 14608 -2469
rect 14356 -2502 14608 -2486
rect 14814 -2486 14830 -2469
rect 15050 -2469 15140 -2452
rect 15198 -2452 15598 -2414
rect 15198 -2469 15288 -2452
rect 15050 -2486 15066 -2469
rect 14814 -2502 15066 -2486
rect 15272 -2486 15288 -2469
rect 15508 -2469 15598 -2452
rect 15656 -2452 16056 -2414
rect 15656 -2469 15746 -2452
rect 15508 -2486 15524 -2469
rect 15272 -2502 15524 -2486
rect 15730 -2486 15746 -2469
rect 15966 -2469 16056 -2452
rect 16114 -2452 16514 -2414
rect 16114 -2469 16204 -2452
rect 15966 -2486 15982 -2469
rect 15730 -2502 15982 -2486
rect 16188 -2486 16204 -2469
rect 16424 -2469 16514 -2452
rect 16572 -2452 16972 -2414
rect 16572 -2469 16662 -2452
rect 16424 -2486 16440 -2469
rect 16188 -2502 16440 -2486
rect 16646 -2486 16662 -2469
rect 16882 -2469 16972 -2452
rect 17030 -2452 17430 -2414
rect 17030 -2469 17120 -2452
rect 16882 -2486 16898 -2469
rect 16646 -2502 16898 -2486
rect 17104 -2486 17120 -2469
rect 17340 -2469 17430 -2452
rect 17488 -2452 17888 -2414
rect 17488 -2469 17578 -2452
rect 17340 -2486 17356 -2469
rect 17104 -2502 17356 -2486
rect 17562 -2486 17578 -2469
rect 17798 -2469 17888 -2452
rect 17946 -2452 18346 -2414
rect 17946 -2469 18036 -2452
rect 17798 -2486 17814 -2469
rect 17562 -2502 17814 -2486
rect 18020 -2486 18036 -2469
rect 18256 -2469 18346 -2452
rect 18256 -2486 18272 -2469
rect 18020 -2502 18272 -2486
rect 8898 -2810 9150 -2794
rect 8898 -2827 8914 -2810
rect 8824 -2844 8914 -2827
rect 9134 -2827 9150 -2810
rect 9356 -2810 9608 -2794
rect 9356 -2827 9372 -2810
rect 9134 -2844 9224 -2827
rect 8824 -2882 9224 -2844
rect 9282 -2844 9372 -2827
rect 9592 -2827 9608 -2810
rect 9814 -2810 10066 -2794
rect 9814 -2827 9830 -2810
rect 9592 -2844 9682 -2827
rect 9282 -2882 9682 -2844
rect 9740 -2844 9830 -2827
rect 10050 -2827 10066 -2810
rect 10272 -2810 10524 -2794
rect 10272 -2827 10288 -2810
rect 10050 -2844 10140 -2827
rect 9740 -2882 10140 -2844
rect 10198 -2844 10288 -2827
rect 10508 -2827 10524 -2810
rect 10730 -2810 10982 -2794
rect 10730 -2827 10746 -2810
rect 10508 -2844 10598 -2827
rect 10198 -2882 10598 -2844
rect 10656 -2844 10746 -2827
rect 10966 -2827 10982 -2810
rect 11188 -2810 11440 -2794
rect 11188 -2827 11204 -2810
rect 10966 -2844 11056 -2827
rect 10656 -2882 11056 -2844
rect 11114 -2844 11204 -2827
rect 11424 -2827 11440 -2810
rect 11646 -2810 11898 -2794
rect 11646 -2827 11662 -2810
rect 11424 -2844 11514 -2827
rect 11114 -2882 11514 -2844
rect 11572 -2844 11662 -2827
rect 11882 -2827 11898 -2810
rect 12104 -2810 12356 -2794
rect 12104 -2827 12120 -2810
rect 11882 -2844 11972 -2827
rect 11572 -2882 11972 -2844
rect 12030 -2844 12120 -2827
rect 12340 -2827 12356 -2810
rect 12562 -2810 12814 -2794
rect 12562 -2827 12578 -2810
rect 12340 -2844 12430 -2827
rect 12030 -2882 12430 -2844
rect 12488 -2844 12578 -2827
rect 12798 -2827 12814 -2810
rect 13020 -2810 13272 -2794
rect 13020 -2827 13036 -2810
rect 12798 -2844 12888 -2827
rect 12488 -2882 12888 -2844
rect 12946 -2844 13036 -2827
rect 13256 -2827 13272 -2810
rect 13256 -2844 13346 -2827
rect 12946 -2882 13346 -2844
rect 8824 -3120 9224 -3082
rect 8824 -3137 8914 -3120
rect 8898 -3154 8914 -3137
rect 9134 -3137 9224 -3120
rect 9282 -3120 9682 -3082
rect 9282 -3137 9372 -3120
rect 9134 -3154 9150 -3137
rect 8898 -3170 9150 -3154
rect 9356 -3154 9372 -3137
rect 9592 -3137 9682 -3120
rect 9740 -3120 10140 -3082
rect 9740 -3137 9830 -3120
rect 9592 -3154 9608 -3137
rect 9356 -3170 9608 -3154
rect 9814 -3154 9830 -3137
rect 10050 -3137 10140 -3120
rect 10198 -3120 10598 -3082
rect 10198 -3137 10288 -3120
rect 10050 -3154 10066 -3137
rect 9814 -3170 10066 -3154
rect 10272 -3154 10288 -3137
rect 10508 -3137 10598 -3120
rect 10656 -3120 11056 -3082
rect 10656 -3137 10746 -3120
rect 10508 -3154 10524 -3137
rect 10272 -3170 10524 -3154
rect 10730 -3154 10746 -3137
rect 10966 -3137 11056 -3120
rect 11114 -3120 11514 -3082
rect 11114 -3137 11204 -3120
rect 10966 -3154 10982 -3137
rect 10730 -3170 10982 -3154
rect 11188 -3154 11204 -3137
rect 11424 -3137 11514 -3120
rect 11572 -3120 11972 -3082
rect 11572 -3137 11662 -3120
rect 11424 -3154 11440 -3137
rect 11188 -3170 11440 -3154
rect 11646 -3154 11662 -3137
rect 11882 -3137 11972 -3120
rect 12030 -3120 12430 -3082
rect 12030 -3137 12120 -3120
rect 11882 -3154 11898 -3137
rect 11646 -3170 11898 -3154
rect 12104 -3154 12120 -3137
rect 12340 -3137 12430 -3120
rect 12488 -3120 12888 -3082
rect 12488 -3137 12578 -3120
rect 12340 -3154 12356 -3137
rect 12104 -3170 12356 -3154
rect 12562 -3154 12578 -3137
rect 12798 -3137 12888 -3120
rect 12946 -3120 13346 -3082
rect 12946 -3137 13036 -3120
rect 12798 -3154 12814 -3137
rect 12562 -3170 12814 -3154
rect 13020 -3154 13036 -3137
rect 13256 -3137 13346 -3120
rect 13256 -3154 13272 -3137
rect 13020 -3170 13272 -3154
rect 23898 -2142 24150 -2126
rect 23898 -2159 23914 -2142
rect 23824 -2176 23914 -2159
rect 24134 -2159 24150 -2142
rect 24356 -2142 24608 -2126
rect 24356 -2159 24372 -2142
rect 24134 -2176 24224 -2159
rect 23824 -2214 24224 -2176
rect 24282 -2176 24372 -2159
rect 24592 -2159 24608 -2142
rect 24814 -2142 25066 -2126
rect 24814 -2159 24830 -2142
rect 24592 -2176 24682 -2159
rect 24282 -2214 24682 -2176
rect 24740 -2176 24830 -2159
rect 25050 -2159 25066 -2142
rect 25272 -2142 25524 -2126
rect 25272 -2159 25288 -2142
rect 25050 -2176 25140 -2159
rect 24740 -2214 25140 -2176
rect 25198 -2176 25288 -2159
rect 25508 -2159 25524 -2142
rect 25730 -2142 25982 -2126
rect 25730 -2159 25746 -2142
rect 25508 -2176 25598 -2159
rect 25198 -2214 25598 -2176
rect 25656 -2176 25746 -2159
rect 25966 -2159 25982 -2142
rect 26188 -2142 26440 -2126
rect 26188 -2159 26204 -2142
rect 25966 -2176 26056 -2159
rect 25656 -2214 26056 -2176
rect 26114 -2176 26204 -2159
rect 26424 -2159 26440 -2142
rect 26646 -2142 26898 -2126
rect 26646 -2159 26662 -2142
rect 26424 -2176 26514 -2159
rect 26114 -2214 26514 -2176
rect 26572 -2176 26662 -2159
rect 26882 -2159 26898 -2142
rect 27104 -2142 27356 -2126
rect 27104 -2159 27120 -2142
rect 26882 -2176 26972 -2159
rect 26572 -2214 26972 -2176
rect 27030 -2176 27120 -2159
rect 27340 -2159 27356 -2142
rect 27562 -2142 27814 -2126
rect 27562 -2159 27578 -2142
rect 27340 -2176 27430 -2159
rect 27030 -2214 27430 -2176
rect 27488 -2176 27578 -2159
rect 27798 -2159 27814 -2142
rect 28020 -2142 28272 -2126
rect 28020 -2159 28036 -2142
rect 27798 -2176 27888 -2159
rect 27488 -2214 27888 -2176
rect 27946 -2176 28036 -2159
rect 28256 -2159 28272 -2142
rect 28898 -2142 29150 -2126
rect 28898 -2159 28914 -2142
rect 28256 -2176 28346 -2159
rect 27946 -2214 28346 -2176
rect 28824 -2176 28914 -2159
rect 29134 -2159 29150 -2142
rect 29356 -2142 29608 -2126
rect 29356 -2159 29372 -2142
rect 29134 -2176 29224 -2159
rect 28824 -2214 29224 -2176
rect 29282 -2176 29372 -2159
rect 29592 -2159 29608 -2142
rect 29814 -2142 30066 -2126
rect 29814 -2159 29830 -2142
rect 29592 -2176 29682 -2159
rect 29282 -2214 29682 -2176
rect 29740 -2176 29830 -2159
rect 30050 -2159 30066 -2142
rect 30272 -2142 30524 -2126
rect 30272 -2159 30288 -2142
rect 30050 -2176 30140 -2159
rect 29740 -2214 30140 -2176
rect 30198 -2176 30288 -2159
rect 30508 -2159 30524 -2142
rect 30730 -2142 30982 -2126
rect 30730 -2159 30746 -2142
rect 30508 -2176 30598 -2159
rect 30198 -2214 30598 -2176
rect 30656 -2176 30746 -2159
rect 30966 -2159 30982 -2142
rect 31188 -2142 31440 -2126
rect 31188 -2159 31204 -2142
rect 30966 -2176 31056 -2159
rect 30656 -2214 31056 -2176
rect 31114 -2176 31204 -2159
rect 31424 -2159 31440 -2142
rect 31646 -2142 31898 -2126
rect 31646 -2159 31662 -2142
rect 31424 -2176 31514 -2159
rect 31114 -2214 31514 -2176
rect 31572 -2176 31662 -2159
rect 31882 -2159 31898 -2142
rect 32104 -2142 32356 -2126
rect 32104 -2159 32120 -2142
rect 31882 -2176 31972 -2159
rect 31572 -2214 31972 -2176
rect 32030 -2176 32120 -2159
rect 32340 -2159 32356 -2142
rect 32562 -2142 32814 -2126
rect 32562 -2159 32578 -2142
rect 32340 -2176 32430 -2159
rect 32030 -2214 32430 -2176
rect 32488 -2176 32578 -2159
rect 32798 -2159 32814 -2142
rect 33020 -2142 33272 -2126
rect 33020 -2159 33036 -2142
rect 32798 -2176 32888 -2159
rect 32488 -2214 32888 -2176
rect 32946 -2176 33036 -2159
rect 33256 -2159 33272 -2142
rect 33256 -2176 33346 -2159
rect 32946 -2214 33346 -2176
rect 23824 -2452 24224 -2414
rect 23824 -2469 23914 -2452
rect 23898 -2486 23914 -2469
rect 24134 -2469 24224 -2452
rect 24282 -2452 24682 -2414
rect 24282 -2469 24372 -2452
rect 24134 -2486 24150 -2469
rect 23898 -2502 24150 -2486
rect 24356 -2486 24372 -2469
rect 24592 -2469 24682 -2452
rect 24740 -2452 25140 -2414
rect 24740 -2469 24830 -2452
rect 24592 -2486 24608 -2469
rect 24356 -2502 24608 -2486
rect 24814 -2486 24830 -2469
rect 25050 -2469 25140 -2452
rect 25198 -2452 25598 -2414
rect 25198 -2469 25288 -2452
rect 25050 -2486 25066 -2469
rect 24814 -2502 25066 -2486
rect 25272 -2486 25288 -2469
rect 25508 -2469 25598 -2452
rect 25656 -2452 26056 -2414
rect 25656 -2469 25746 -2452
rect 25508 -2486 25524 -2469
rect 25272 -2502 25524 -2486
rect 25730 -2486 25746 -2469
rect 25966 -2469 26056 -2452
rect 26114 -2452 26514 -2414
rect 26114 -2469 26204 -2452
rect 25966 -2486 25982 -2469
rect 25730 -2502 25982 -2486
rect 26188 -2486 26204 -2469
rect 26424 -2469 26514 -2452
rect 26572 -2452 26972 -2414
rect 26572 -2469 26662 -2452
rect 26424 -2486 26440 -2469
rect 26188 -2502 26440 -2486
rect 26646 -2486 26662 -2469
rect 26882 -2469 26972 -2452
rect 27030 -2452 27430 -2414
rect 27030 -2469 27120 -2452
rect 26882 -2486 26898 -2469
rect 26646 -2502 26898 -2486
rect 27104 -2486 27120 -2469
rect 27340 -2469 27430 -2452
rect 27488 -2452 27888 -2414
rect 27488 -2469 27578 -2452
rect 27340 -2486 27356 -2469
rect 27104 -2502 27356 -2486
rect 27562 -2486 27578 -2469
rect 27798 -2469 27888 -2452
rect 27946 -2452 28346 -2414
rect 27946 -2469 28036 -2452
rect 27798 -2486 27814 -2469
rect 27562 -2502 27814 -2486
rect 28020 -2486 28036 -2469
rect 28256 -2469 28346 -2452
rect 28824 -2452 29224 -2414
rect 28824 -2469 28914 -2452
rect 28256 -2486 28272 -2469
rect 28020 -2502 28272 -2486
rect 28898 -2486 28914 -2469
rect 29134 -2469 29224 -2452
rect 29282 -2452 29682 -2414
rect 29282 -2469 29372 -2452
rect 29134 -2486 29150 -2469
rect 28898 -2502 29150 -2486
rect 29356 -2486 29372 -2469
rect 29592 -2469 29682 -2452
rect 29740 -2452 30140 -2414
rect 29740 -2469 29830 -2452
rect 29592 -2486 29608 -2469
rect 29356 -2502 29608 -2486
rect 29814 -2486 29830 -2469
rect 30050 -2469 30140 -2452
rect 30198 -2452 30598 -2414
rect 30198 -2469 30288 -2452
rect 30050 -2486 30066 -2469
rect 29814 -2502 30066 -2486
rect 30272 -2486 30288 -2469
rect 30508 -2469 30598 -2452
rect 30656 -2452 31056 -2414
rect 30656 -2469 30746 -2452
rect 30508 -2486 30524 -2469
rect 30272 -2502 30524 -2486
rect 30730 -2486 30746 -2469
rect 30966 -2469 31056 -2452
rect 31114 -2452 31514 -2414
rect 31114 -2469 31204 -2452
rect 30966 -2486 30982 -2469
rect 30730 -2502 30982 -2486
rect 31188 -2486 31204 -2469
rect 31424 -2469 31514 -2452
rect 31572 -2452 31972 -2414
rect 31572 -2469 31662 -2452
rect 31424 -2486 31440 -2469
rect 31188 -2502 31440 -2486
rect 31646 -2486 31662 -2469
rect 31882 -2469 31972 -2452
rect 32030 -2452 32430 -2414
rect 32030 -2469 32120 -2452
rect 31882 -2486 31898 -2469
rect 31646 -2502 31898 -2486
rect 32104 -2486 32120 -2469
rect 32340 -2469 32430 -2452
rect 32488 -2452 32888 -2414
rect 32488 -2469 32578 -2452
rect 32340 -2486 32356 -2469
rect 32104 -2502 32356 -2486
rect 32562 -2486 32578 -2469
rect 32798 -2469 32888 -2452
rect 32946 -2452 33346 -2414
rect 32946 -2469 33036 -2452
rect 32798 -2486 32814 -2469
rect 32562 -2502 32814 -2486
rect 33020 -2486 33036 -2469
rect 33256 -2469 33346 -2452
rect 33256 -2486 33272 -2469
rect 33020 -2502 33272 -2486
rect 23898 -2810 24150 -2794
rect 23898 -2827 23914 -2810
rect 23824 -2844 23914 -2827
rect 24134 -2827 24150 -2810
rect 24356 -2810 24608 -2794
rect 24356 -2827 24372 -2810
rect 24134 -2844 24224 -2827
rect 23824 -2882 24224 -2844
rect 24282 -2844 24372 -2827
rect 24592 -2827 24608 -2810
rect 24814 -2810 25066 -2794
rect 24814 -2827 24830 -2810
rect 24592 -2844 24682 -2827
rect 24282 -2882 24682 -2844
rect 24740 -2844 24830 -2827
rect 25050 -2827 25066 -2810
rect 25272 -2810 25524 -2794
rect 25272 -2827 25288 -2810
rect 25050 -2844 25140 -2827
rect 24740 -2882 25140 -2844
rect 25198 -2844 25288 -2827
rect 25508 -2827 25524 -2810
rect 25730 -2810 25982 -2794
rect 25730 -2827 25746 -2810
rect 25508 -2844 25598 -2827
rect 25198 -2882 25598 -2844
rect 25656 -2844 25746 -2827
rect 25966 -2827 25982 -2810
rect 26188 -2810 26440 -2794
rect 26188 -2827 26204 -2810
rect 25966 -2844 26056 -2827
rect 25656 -2882 26056 -2844
rect 26114 -2844 26204 -2827
rect 26424 -2827 26440 -2810
rect 26646 -2810 26898 -2794
rect 26646 -2827 26662 -2810
rect 26424 -2844 26514 -2827
rect 26114 -2882 26514 -2844
rect 26572 -2844 26662 -2827
rect 26882 -2827 26898 -2810
rect 27104 -2810 27356 -2794
rect 27104 -2827 27120 -2810
rect 26882 -2844 26972 -2827
rect 26572 -2882 26972 -2844
rect 27030 -2844 27120 -2827
rect 27340 -2827 27356 -2810
rect 27562 -2810 27814 -2794
rect 27562 -2827 27578 -2810
rect 27340 -2844 27430 -2827
rect 27030 -2882 27430 -2844
rect 27488 -2844 27578 -2827
rect 27798 -2827 27814 -2810
rect 28020 -2810 28272 -2794
rect 28020 -2827 28036 -2810
rect 27798 -2844 27888 -2827
rect 27488 -2882 27888 -2844
rect 27946 -2844 28036 -2827
rect 28256 -2827 28272 -2810
rect 28256 -2844 28346 -2827
rect 27946 -2882 28346 -2844
rect 23824 -3120 24224 -3082
rect 23824 -3137 23914 -3120
rect 23898 -3154 23914 -3137
rect 24134 -3137 24224 -3120
rect 24282 -3120 24682 -3082
rect 24282 -3137 24372 -3120
rect 24134 -3154 24150 -3137
rect 23898 -3170 24150 -3154
rect 24356 -3154 24372 -3137
rect 24592 -3137 24682 -3120
rect 24740 -3120 25140 -3082
rect 24740 -3137 24830 -3120
rect 24592 -3154 24608 -3137
rect 24356 -3170 24608 -3154
rect 24814 -3154 24830 -3137
rect 25050 -3137 25140 -3120
rect 25198 -3120 25598 -3082
rect 25198 -3137 25288 -3120
rect 25050 -3154 25066 -3137
rect 24814 -3170 25066 -3154
rect 25272 -3154 25288 -3137
rect 25508 -3137 25598 -3120
rect 25656 -3120 26056 -3082
rect 25656 -3137 25746 -3120
rect 25508 -3154 25524 -3137
rect 25272 -3170 25524 -3154
rect 25730 -3154 25746 -3137
rect 25966 -3137 26056 -3120
rect 26114 -3120 26514 -3082
rect 26114 -3137 26204 -3120
rect 25966 -3154 25982 -3137
rect 25730 -3170 25982 -3154
rect 26188 -3154 26204 -3137
rect 26424 -3137 26514 -3120
rect 26572 -3120 26972 -3082
rect 26572 -3137 26662 -3120
rect 26424 -3154 26440 -3137
rect 26188 -3170 26440 -3154
rect 26646 -3154 26662 -3137
rect 26882 -3137 26972 -3120
rect 27030 -3120 27430 -3082
rect 27030 -3137 27120 -3120
rect 26882 -3154 26898 -3137
rect 26646 -3170 26898 -3154
rect 27104 -3154 27120 -3137
rect 27340 -3137 27430 -3120
rect 27488 -3120 27888 -3082
rect 27488 -3137 27578 -3120
rect 27340 -3154 27356 -3137
rect 27104 -3170 27356 -3154
rect 27562 -3154 27578 -3137
rect 27798 -3137 27888 -3120
rect 27946 -3120 28346 -3082
rect 27946 -3137 28036 -3120
rect 27798 -3154 27814 -3137
rect 27562 -3170 27814 -3154
rect 28020 -3154 28036 -3137
rect 28256 -3137 28346 -3120
rect 28256 -3154 28272 -3137
rect 28020 -3170 28272 -3154
rect 17830 -5602 18082 -5586
rect 17830 -5619 17846 -5602
rect 17756 -5636 17846 -5619
rect 18066 -5619 18082 -5602
rect 18288 -5602 18540 -5586
rect 18288 -5619 18304 -5602
rect 18066 -5636 18156 -5619
rect 17756 -5674 18156 -5636
rect 18214 -5636 18304 -5619
rect 18524 -5619 18540 -5602
rect 18746 -5602 18998 -5586
rect 18746 -5619 18762 -5602
rect 18524 -5636 18614 -5619
rect 18214 -5674 18614 -5636
rect 18672 -5636 18762 -5619
rect 18982 -5619 18998 -5602
rect 19204 -5602 19456 -5586
rect 19204 -5619 19220 -5602
rect 18982 -5636 19072 -5619
rect 18672 -5674 19072 -5636
rect 19130 -5636 19220 -5619
rect 19440 -5619 19456 -5602
rect 19662 -5602 19914 -5586
rect 19662 -5619 19678 -5602
rect 19440 -5636 19530 -5619
rect 19130 -5674 19530 -5636
rect 19588 -5636 19678 -5619
rect 19898 -5619 19914 -5602
rect 20120 -5602 20372 -5586
rect 20120 -5619 20136 -5602
rect 19898 -5636 19988 -5619
rect 19588 -5674 19988 -5636
rect 20046 -5636 20136 -5619
rect 20356 -5619 20372 -5602
rect 20578 -5602 20830 -5586
rect 20578 -5619 20594 -5602
rect 20356 -5636 20446 -5619
rect 20046 -5674 20446 -5636
rect 20504 -5636 20594 -5619
rect 20814 -5619 20830 -5602
rect 21036 -5602 21288 -5586
rect 21036 -5619 21052 -5602
rect 20814 -5636 20904 -5619
rect 20504 -5674 20904 -5636
rect 20962 -5636 21052 -5619
rect 21272 -5619 21288 -5602
rect 21494 -5602 21746 -5586
rect 21494 -5619 21510 -5602
rect 21272 -5636 21362 -5619
rect 20962 -5674 21362 -5636
rect 21420 -5636 21510 -5619
rect 21730 -5619 21746 -5602
rect 21952 -5602 22204 -5586
rect 21952 -5619 21968 -5602
rect 21730 -5636 21820 -5619
rect 21420 -5674 21820 -5636
rect 21878 -5636 21968 -5619
rect 22188 -5619 22204 -5602
rect 22188 -5636 22278 -5619
rect 21878 -5674 22278 -5636
rect 17756 -5912 18156 -5874
rect 17756 -5929 17846 -5912
rect 17830 -5946 17846 -5929
rect 18066 -5929 18156 -5912
rect 18214 -5912 18614 -5874
rect 18214 -5929 18304 -5912
rect 18066 -5946 18082 -5929
rect 17830 -5962 18082 -5946
rect 18288 -5946 18304 -5929
rect 18524 -5929 18614 -5912
rect 18672 -5912 19072 -5874
rect 18672 -5929 18762 -5912
rect 18524 -5946 18540 -5929
rect 18288 -5962 18540 -5946
rect 18746 -5946 18762 -5929
rect 18982 -5929 19072 -5912
rect 19130 -5912 19530 -5874
rect 19130 -5929 19220 -5912
rect 18982 -5946 18998 -5929
rect 18746 -5962 18998 -5946
rect 19204 -5946 19220 -5929
rect 19440 -5929 19530 -5912
rect 19588 -5912 19988 -5874
rect 19588 -5929 19678 -5912
rect 19440 -5946 19456 -5929
rect 19204 -5962 19456 -5946
rect 19662 -5946 19678 -5929
rect 19898 -5929 19988 -5912
rect 20046 -5912 20446 -5874
rect 20046 -5929 20136 -5912
rect 19898 -5946 19914 -5929
rect 19662 -5962 19914 -5946
rect 20120 -5946 20136 -5929
rect 20356 -5929 20446 -5912
rect 20504 -5912 20904 -5874
rect 20504 -5929 20594 -5912
rect 20356 -5946 20372 -5929
rect 20120 -5962 20372 -5946
rect 20578 -5946 20594 -5929
rect 20814 -5929 20904 -5912
rect 20962 -5912 21362 -5874
rect 20962 -5929 21052 -5912
rect 20814 -5946 20830 -5929
rect 20578 -5962 20830 -5946
rect 21036 -5946 21052 -5929
rect 21272 -5929 21362 -5912
rect 21420 -5912 21820 -5874
rect 21420 -5929 21510 -5912
rect 21272 -5946 21288 -5929
rect 21036 -5962 21288 -5946
rect 21494 -5946 21510 -5929
rect 21730 -5929 21820 -5912
rect 21878 -5912 22278 -5874
rect 21878 -5929 21968 -5912
rect 21730 -5946 21746 -5929
rect 21494 -5962 21746 -5946
rect 21952 -5946 21968 -5929
rect 22188 -5929 22278 -5912
rect 22188 -5946 22204 -5929
rect 21952 -5962 22204 -5946
rect 12830 -6270 13082 -6254
rect 12830 -6287 12846 -6270
rect 12756 -6304 12846 -6287
rect 13066 -6287 13082 -6270
rect 13288 -6270 13540 -6254
rect 13288 -6287 13304 -6270
rect 13066 -6304 13156 -6287
rect 12756 -6342 13156 -6304
rect 13214 -6304 13304 -6287
rect 13524 -6287 13540 -6270
rect 13746 -6270 13998 -6254
rect 13746 -6287 13762 -6270
rect 13524 -6304 13614 -6287
rect 13214 -6342 13614 -6304
rect 13672 -6304 13762 -6287
rect 13982 -6287 13998 -6270
rect 14204 -6270 14456 -6254
rect 14204 -6287 14220 -6270
rect 13982 -6304 14072 -6287
rect 13672 -6342 14072 -6304
rect 14130 -6304 14220 -6287
rect 14440 -6287 14456 -6270
rect 14662 -6270 14914 -6254
rect 14662 -6287 14678 -6270
rect 14440 -6304 14530 -6287
rect 14130 -6342 14530 -6304
rect 14588 -6304 14678 -6287
rect 14898 -6287 14914 -6270
rect 15120 -6270 15372 -6254
rect 15120 -6287 15136 -6270
rect 14898 -6304 14988 -6287
rect 14588 -6342 14988 -6304
rect 15046 -6304 15136 -6287
rect 15356 -6287 15372 -6270
rect 15578 -6270 15830 -6254
rect 15578 -6287 15594 -6270
rect 15356 -6304 15446 -6287
rect 15046 -6342 15446 -6304
rect 15504 -6304 15594 -6287
rect 15814 -6287 15830 -6270
rect 16036 -6270 16288 -6254
rect 16036 -6287 16052 -6270
rect 15814 -6304 15904 -6287
rect 15504 -6342 15904 -6304
rect 15962 -6304 16052 -6287
rect 16272 -6287 16288 -6270
rect 16494 -6270 16746 -6254
rect 16494 -6287 16510 -6270
rect 16272 -6304 16362 -6287
rect 15962 -6342 16362 -6304
rect 16420 -6304 16510 -6287
rect 16730 -6287 16746 -6270
rect 16952 -6270 17204 -6254
rect 16952 -6287 16968 -6270
rect 16730 -6304 16820 -6287
rect 16420 -6342 16820 -6304
rect 16878 -6304 16968 -6287
rect 17188 -6287 17204 -6270
rect 17830 -6270 18082 -6254
rect 17830 -6287 17846 -6270
rect 17188 -6304 17278 -6287
rect 16878 -6342 17278 -6304
rect 17756 -6304 17846 -6287
rect 18066 -6287 18082 -6270
rect 18288 -6270 18540 -6254
rect 18288 -6287 18304 -6270
rect 18066 -6304 18156 -6287
rect 17756 -6342 18156 -6304
rect 18214 -6304 18304 -6287
rect 18524 -6287 18540 -6270
rect 18746 -6270 18998 -6254
rect 18746 -6287 18762 -6270
rect 18524 -6304 18614 -6287
rect 18214 -6342 18614 -6304
rect 18672 -6304 18762 -6287
rect 18982 -6287 18998 -6270
rect 19204 -6270 19456 -6254
rect 19204 -6287 19220 -6270
rect 18982 -6304 19072 -6287
rect 18672 -6342 19072 -6304
rect 19130 -6304 19220 -6287
rect 19440 -6287 19456 -6270
rect 19662 -6270 19914 -6254
rect 19662 -6287 19678 -6270
rect 19440 -6304 19530 -6287
rect 19130 -6342 19530 -6304
rect 19588 -6304 19678 -6287
rect 19898 -6287 19914 -6270
rect 20120 -6270 20372 -6254
rect 20120 -6287 20136 -6270
rect 19898 -6304 19988 -6287
rect 19588 -6342 19988 -6304
rect 20046 -6304 20136 -6287
rect 20356 -6287 20372 -6270
rect 20578 -6270 20830 -6254
rect 20578 -6287 20594 -6270
rect 20356 -6304 20446 -6287
rect 20046 -6342 20446 -6304
rect 20504 -6304 20594 -6287
rect 20814 -6287 20830 -6270
rect 21036 -6270 21288 -6254
rect 21036 -6287 21052 -6270
rect 20814 -6304 20904 -6287
rect 20504 -6342 20904 -6304
rect 20962 -6304 21052 -6287
rect 21272 -6287 21288 -6270
rect 21494 -6270 21746 -6254
rect 21494 -6287 21510 -6270
rect 21272 -6304 21362 -6287
rect 20962 -6342 21362 -6304
rect 21420 -6304 21510 -6287
rect 21730 -6287 21746 -6270
rect 21952 -6270 22204 -6254
rect 21952 -6287 21968 -6270
rect 21730 -6304 21820 -6287
rect 21420 -6342 21820 -6304
rect 21878 -6304 21968 -6287
rect 22188 -6287 22204 -6270
rect 22188 -6304 22278 -6287
rect 21878 -6342 22278 -6304
rect 12756 -6580 13156 -6542
rect 12756 -6597 12846 -6580
rect 12830 -6614 12846 -6597
rect 13066 -6597 13156 -6580
rect 13214 -6580 13614 -6542
rect 13214 -6597 13304 -6580
rect 13066 -6614 13082 -6597
rect 12830 -6630 13082 -6614
rect 13288 -6614 13304 -6597
rect 13524 -6597 13614 -6580
rect 13672 -6580 14072 -6542
rect 13672 -6597 13762 -6580
rect 13524 -6614 13540 -6597
rect 13288 -6630 13540 -6614
rect 13746 -6614 13762 -6597
rect 13982 -6597 14072 -6580
rect 14130 -6580 14530 -6542
rect 14130 -6597 14220 -6580
rect 13982 -6614 13998 -6597
rect 13746 -6630 13998 -6614
rect 14204 -6614 14220 -6597
rect 14440 -6597 14530 -6580
rect 14588 -6580 14988 -6542
rect 14588 -6597 14678 -6580
rect 14440 -6614 14456 -6597
rect 14204 -6630 14456 -6614
rect 14662 -6614 14678 -6597
rect 14898 -6597 14988 -6580
rect 15046 -6580 15446 -6542
rect 15046 -6597 15136 -6580
rect 14898 -6614 14914 -6597
rect 14662 -6630 14914 -6614
rect 15120 -6614 15136 -6597
rect 15356 -6597 15446 -6580
rect 15504 -6580 15904 -6542
rect 15504 -6597 15594 -6580
rect 15356 -6614 15372 -6597
rect 15120 -6630 15372 -6614
rect 15578 -6614 15594 -6597
rect 15814 -6597 15904 -6580
rect 15962 -6580 16362 -6542
rect 15962 -6597 16052 -6580
rect 15814 -6614 15830 -6597
rect 15578 -6630 15830 -6614
rect 16036 -6614 16052 -6597
rect 16272 -6597 16362 -6580
rect 16420 -6580 16820 -6542
rect 16420 -6597 16510 -6580
rect 16272 -6614 16288 -6597
rect 16036 -6630 16288 -6614
rect 16494 -6614 16510 -6597
rect 16730 -6597 16820 -6580
rect 16878 -6580 17278 -6542
rect 16878 -6597 16968 -6580
rect 16730 -6614 16746 -6597
rect 16494 -6630 16746 -6614
rect 16952 -6614 16968 -6597
rect 17188 -6597 17278 -6580
rect 17756 -6580 18156 -6542
rect 17756 -6597 17846 -6580
rect 17188 -6614 17204 -6597
rect 16952 -6630 17204 -6614
rect 17830 -6614 17846 -6597
rect 18066 -6597 18156 -6580
rect 18214 -6580 18614 -6542
rect 18214 -6597 18304 -6580
rect 18066 -6614 18082 -6597
rect 17830 -6630 18082 -6614
rect 18288 -6614 18304 -6597
rect 18524 -6597 18614 -6580
rect 18672 -6580 19072 -6542
rect 18672 -6597 18762 -6580
rect 18524 -6614 18540 -6597
rect 18288 -6630 18540 -6614
rect 18746 -6614 18762 -6597
rect 18982 -6597 19072 -6580
rect 19130 -6580 19530 -6542
rect 19130 -6597 19220 -6580
rect 18982 -6614 18998 -6597
rect 18746 -6630 18998 -6614
rect 19204 -6614 19220 -6597
rect 19440 -6597 19530 -6580
rect 19588 -6580 19988 -6542
rect 19588 -6597 19678 -6580
rect 19440 -6614 19456 -6597
rect 19204 -6630 19456 -6614
rect 19662 -6614 19678 -6597
rect 19898 -6597 19988 -6580
rect 20046 -6580 20446 -6542
rect 20046 -6597 20136 -6580
rect 19898 -6614 19914 -6597
rect 19662 -6630 19914 -6614
rect 20120 -6614 20136 -6597
rect 20356 -6597 20446 -6580
rect 20504 -6580 20904 -6542
rect 20504 -6597 20594 -6580
rect 20356 -6614 20372 -6597
rect 20120 -6630 20372 -6614
rect 20578 -6614 20594 -6597
rect 20814 -6597 20904 -6580
rect 20962 -6580 21362 -6542
rect 20962 -6597 21052 -6580
rect 20814 -6614 20830 -6597
rect 20578 -6630 20830 -6614
rect 21036 -6614 21052 -6597
rect 21272 -6597 21362 -6580
rect 21420 -6580 21820 -6542
rect 21420 -6597 21510 -6580
rect 21272 -6614 21288 -6597
rect 21036 -6630 21288 -6614
rect 21494 -6614 21510 -6597
rect 21730 -6597 21820 -6580
rect 21878 -6580 22278 -6542
rect 21878 -6597 21968 -6580
rect 21730 -6614 21746 -6597
rect 21494 -6630 21746 -6614
rect 21952 -6614 21968 -6597
rect 22188 -6597 22278 -6580
rect 22188 -6614 22204 -6597
rect 21952 -6630 22204 -6614
rect 32830 -5602 33082 -5586
rect 32830 -5619 32846 -5602
rect 32756 -5636 32846 -5619
rect 33066 -5619 33082 -5602
rect 33288 -5602 33540 -5586
rect 33288 -5619 33304 -5602
rect 33066 -5636 33156 -5619
rect 32756 -5674 33156 -5636
rect 33214 -5636 33304 -5619
rect 33524 -5619 33540 -5602
rect 33746 -5602 33998 -5586
rect 33746 -5619 33762 -5602
rect 33524 -5636 33614 -5619
rect 33214 -5674 33614 -5636
rect 33672 -5636 33762 -5619
rect 33982 -5619 33998 -5602
rect 34204 -5602 34456 -5586
rect 34204 -5619 34220 -5602
rect 33982 -5636 34072 -5619
rect 33672 -5674 34072 -5636
rect 34130 -5636 34220 -5619
rect 34440 -5619 34456 -5602
rect 34662 -5602 34914 -5586
rect 34662 -5619 34678 -5602
rect 34440 -5636 34530 -5619
rect 34130 -5674 34530 -5636
rect 34588 -5636 34678 -5619
rect 34898 -5619 34914 -5602
rect 35120 -5602 35372 -5586
rect 35120 -5619 35136 -5602
rect 34898 -5636 34988 -5619
rect 34588 -5674 34988 -5636
rect 35046 -5636 35136 -5619
rect 35356 -5619 35372 -5602
rect 35578 -5602 35830 -5586
rect 35578 -5619 35594 -5602
rect 35356 -5636 35446 -5619
rect 35046 -5674 35446 -5636
rect 35504 -5636 35594 -5619
rect 35814 -5619 35830 -5602
rect 36036 -5602 36288 -5586
rect 36036 -5619 36052 -5602
rect 35814 -5636 35904 -5619
rect 35504 -5674 35904 -5636
rect 35962 -5636 36052 -5619
rect 36272 -5619 36288 -5602
rect 36494 -5602 36746 -5586
rect 36494 -5619 36510 -5602
rect 36272 -5636 36362 -5619
rect 35962 -5674 36362 -5636
rect 36420 -5636 36510 -5619
rect 36730 -5619 36746 -5602
rect 36952 -5602 37204 -5586
rect 36952 -5619 36968 -5602
rect 36730 -5636 36820 -5619
rect 36420 -5674 36820 -5636
rect 36878 -5636 36968 -5619
rect 37188 -5619 37204 -5602
rect 37188 -5636 37278 -5619
rect 36878 -5674 37278 -5636
rect 32756 -5912 33156 -5874
rect 32756 -5929 32846 -5912
rect 32830 -5946 32846 -5929
rect 33066 -5929 33156 -5912
rect 33214 -5912 33614 -5874
rect 33214 -5929 33304 -5912
rect 33066 -5946 33082 -5929
rect 32830 -5962 33082 -5946
rect 33288 -5946 33304 -5929
rect 33524 -5929 33614 -5912
rect 33672 -5912 34072 -5874
rect 33672 -5929 33762 -5912
rect 33524 -5946 33540 -5929
rect 33288 -5962 33540 -5946
rect 33746 -5946 33762 -5929
rect 33982 -5929 34072 -5912
rect 34130 -5912 34530 -5874
rect 34130 -5929 34220 -5912
rect 33982 -5946 33998 -5929
rect 33746 -5962 33998 -5946
rect 34204 -5946 34220 -5929
rect 34440 -5929 34530 -5912
rect 34588 -5912 34988 -5874
rect 34588 -5929 34678 -5912
rect 34440 -5946 34456 -5929
rect 34204 -5962 34456 -5946
rect 34662 -5946 34678 -5929
rect 34898 -5929 34988 -5912
rect 35046 -5912 35446 -5874
rect 35046 -5929 35136 -5912
rect 34898 -5946 34914 -5929
rect 34662 -5962 34914 -5946
rect 35120 -5946 35136 -5929
rect 35356 -5929 35446 -5912
rect 35504 -5912 35904 -5874
rect 35504 -5929 35594 -5912
rect 35356 -5946 35372 -5929
rect 35120 -5962 35372 -5946
rect 35578 -5946 35594 -5929
rect 35814 -5929 35904 -5912
rect 35962 -5912 36362 -5874
rect 35962 -5929 36052 -5912
rect 35814 -5946 35830 -5929
rect 35578 -5962 35830 -5946
rect 36036 -5946 36052 -5929
rect 36272 -5929 36362 -5912
rect 36420 -5912 36820 -5874
rect 36420 -5929 36510 -5912
rect 36272 -5946 36288 -5929
rect 36036 -5962 36288 -5946
rect 36494 -5946 36510 -5929
rect 36730 -5929 36820 -5912
rect 36878 -5912 37278 -5874
rect 36878 -5929 36968 -5912
rect 36730 -5946 36746 -5929
rect 36494 -5962 36746 -5946
rect 36952 -5946 36968 -5929
rect 37188 -5929 37278 -5912
rect 37188 -5946 37204 -5929
rect 36952 -5962 37204 -5946
rect 27830 -6270 28082 -6254
rect 27830 -6287 27846 -6270
rect 27756 -6304 27846 -6287
rect 28066 -6287 28082 -6270
rect 28288 -6270 28540 -6254
rect 28288 -6287 28304 -6270
rect 28066 -6304 28156 -6287
rect 27756 -6342 28156 -6304
rect 28214 -6304 28304 -6287
rect 28524 -6287 28540 -6270
rect 28746 -6270 28998 -6254
rect 28746 -6287 28762 -6270
rect 28524 -6304 28614 -6287
rect 28214 -6342 28614 -6304
rect 28672 -6304 28762 -6287
rect 28982 -6287 28998 -6270
rect 29204 -6270 29456 -6254
rect 29204 -6287 29220 -6270
rect 28982 -6304 29072 -6287
rect 28672 -6342 29072 -6304
rect 29130 -6304 29220 -6287
rect 29440 -6287 29456 -6270
rect 29662 -6270 29914 -6254
rect 29662 -6287 29678 -6270
rect 29440 -6304 29530 -6287
rect 29130 -6342 29530 -6304
rect 29588 -6304 29678 -6287
rect 29898 -6287 29914 -6270
rect 30120 -6270 30372 -6254
rect 30120 -6287 30136 -6270
rect 29898 -6304 29988 -6287
rect 29588 -6342 29988 -6304
rect 30046 -6304 30136 -6287
rect 30356 -6287 30372 -6270
rect 30578 -6270 30830 -6254
rect 30578 -6287 30594 -6270
rect 30356 -6304 30446 -6287
rect 30046 -6342 30446 -6304
rect 30504 -6304 30594 -6287
rect 30814 -6287 30830 -6270
rect 31036 -6270 31288 -6254
rect 31036 -6287 31052 -6270
rect 30814 -6304 30904 -6287
rect 30504 -6342 30904 -6304
rect 30962 -6304 31052 -6287
rect 31272 -6287 31288 -6270
rect 31494 -6270 31746 -6254
rect 31494 -6287 31510 -6270
rect 31272 -6304 31362 -6287
rect 30962 -6342 31362 -6304
rect 31420 -6304 31510 -6287
rect 31730 -6287 31746 -6270
rect 31952 -6270 32204 -6254
rect 31952 -6287 31968 -6270
rect 31730 -6304 31820 -6287
rect 31420 -6342 31820 -6304
rect 31878 -6304 31968 -6287
rect 32188 -6287 32204 -6270
rect 32830 -6270 33082 -6254
rect 32830 -6287 32846 -6270
rect 32188 -6304 32278 -6287
rect 31878 -6342 32278 -6304
rect 32756 -6304 32846 -6287
rect 33066 -6287 33082 -6270
rect 33288 -6270 33540 -6254
rect 33288 -6287 33304 -6270
rect 33066 -6304 33156 -6287
rect 32756 -6342 33156 -6304
rect 33214 -6304 33304 -6287
rect 33524 -6287 33540 -6270
rect 33746 -6270 33998 -6254
rect 33746 -6287 33762 -6270
rect 33524 -6304 33614 -6287
rect 33214 -6342 33614 -6304
rect 33672 -6304 33762 -6287
rect 33982 -6287 33998 -6270
rect 34204 -6270 34456 -6254
rect 34204 -6287 34220 -6270
rect 33982 -6304 34072 -6287
rect 33672 -6342 34072 -6304
rect 34130 -6304 34220 -6287
rect 34440 -6287 34456 -6270
rect 34662 -6270 34914 -6254
rect 34662 -6287 34678 -6270
rect 34440 -6304 34530 -6287
rect 34130 -6342 34530 -6304
rect 34588 -6304 34678 -6287
rect 34898 -6287 34914 -6270
rect 35120 -6270 35372 -6254
rect 35120 -6287 35136 -6270
rect 34898 -6304 34988 -6287
rect 34588 -6342 34988 -6304
rect 35046 -6304 35136 -6287
rect 35356 -6287 35372 -6270
rect 35578 -6270 35830 -6254
rect 35578 -6287 35594 -6270
rect 35356 -6304 35446 -6287
rect 35046 -6342 35446 -6304
rect 35504 -6304 35594 -6287
rect 35814 -6287 35830 -6270
rect 36036 -6270 36288 -6254
rect 36036 -6287 36052 -6270
rect 35814 -6304 35904 -6287
rect 35504 -6342 35904 -6304
rect 35962 -6304 36052 -6287
rect 36272 -6287 36288 -6270
rect 36494 -6270 36746 -6254
rect 36494 -6287 36510 -6270
rect 36272 -6304 36362 -6287
rect 35962 -6342 36362 -6304
rect 36420 -6304 36510 -6287
rect 36730 -6287 36746 -6270
rect 36952 -6270 37204 -6254
rect 36952 -6287 36968 -6270
rect 36730 -6304 36820 -6287
rect 36420 -6342 36820 -6304
rect 36878 -6304 36968 -6287
rect 37188 -6287 37204 -6270
rect 37188 -6304 37278 -6287
rect 36878 -6342 37278 -6304
rect 27756 -6580 28156 -6542
rect 27756 -6597 27846 -6580
rect 27830 -6614 27846 -6597
rect 28066 -6597 28156 -6580
rect 28214 -6580 28614 -6542
rect 28214 -6597 28304 -6580
rect 28066 -6614 28082 -6597
rect 27830 -6630 28082 -6614
rect 28288 -6614 28304 -6597
rect 28524 -6597 28614 -6580
rect 28672 -6580 29072 -6542
rect 28672 -6597 28762 -6580
rect 28524 -6614 28540 -6597
rect 28288 -6630 28540 -6614
rect 28746 -6614 28762 -6597
rect 28982 -6597 29072 -6580
rect 29130 -6580 29530 -6542
rect 29130 -6597 29220 -6580
rect 28982 -6614 28998 -6597
rect 28746 -6630 28998 -6614
rect 29204 -6614 29220 -6597
rect 29440 -6597 29530 -6580
rect 29588 -6580 29988 -6542
rect 29588 -6597 29678 -6580
rect 29440 -6614 29456 -6597
rect 29204 -6630 29456 -6614
rect 29662 -6614 29678 -6597
rect 29898 -6597 29988 -6580
rect 30046 -6580 30446 -6542
rect 30046 -6597 30136 -6580
rect 29898 -6614 29914 -6597
rect 29662 -6630 29914 -6614
rect 30120 -6614 30136 -6597
rect 30356 -6597 30446 -6580
rect 30504 -6580 30904 -6542
rect 30504 -6597 30594 -6580
rect 30356 -6614 30372 -6597
rect 30120 -6630 30372 -6614
rect 30578 -6614 30594 -6597
rect 30814 -6597 30904 -6580
rect 30962 -6580 31362 -6542
rect 30962 -6597 31052 -6580
rect 30814 -6614 30830 -6597
rect 30578 -6630 30830 -6614
rect 31036 -6614 31052 -6597
rect 31272 -6597 31362 -6580
rect 31420 -6580 31820 -6542
rect 31420 -6597 31510 -6580
rect 31272 -6614 31288 -6597
rect 31036 -6630 31288 -6614
rect 31494 -6614 31510 -6597
rect 31730 -6597 31820 -6580
rect 31878 -6580 32278 -6542
rect 31878 -6597 31968 -6580
rect 31730 -6614 31746 -6597
rect 31494 -6630 31746 -6614
rect 31952 -6614 31968 -6597
rect 32188 -6597 32278 -6580
rect 32756 -6580 33156 -6542
rect 32756 -6597 32846 -6580
rect 32188 -6614 32204 -6597
rect 31952 -6630 32204 -6614
rect 32830 -6614 32846 -6597
rect 33066 -6597 33156 -6580
rect 33214 -6580 33614 -6542
rect 33214 -6597 33304 -6580
rect 33066 -6614 33082 -6597
rect 32830 -6630 33082 -6614
rect 33288 -6614 33304 -6597
rect 33524 -6597 33614 -6580
rect 33672 -6580 34072 -6542
rect 33672 -6597 33762 -6580
rect 33524 -6614 33540 -6597
rect 33288 -6630 33540 -6614
rect 33746 -6614 33762 -6597
rect 33982 -6597 34072 -6580
rect 34130 -6580 34530 -6542
rect 34130 -6597 34220 -6580
rect 33982 -6614 33998 -6597
rect 33746 -6630 33998 -6614
rect 34204 -6614 34220 -6597
rect 34440 -6597 34530 -6580
rect 34588 -6580 34988 -6542
rect 34588 -6597 34678 -6580
rect 34440 -6614 34456 -6597
rect 34204 -6630 34456 -6614
rect 34662 -6614 34678 -6597
rect 34898 -6597 34988 -6580
rect 35046 -6580 35446 -6542
rect 35046 -6597 35136 -6580
rect 34898 -6614 34914 -6597
rect 34662 -6630 34914 -6614
rect 35120 -6614 35136 -6597
rect 35356 -6597 35446 -6580
rect 35504 -6580 35904 -6542
rect 35504 -6597 35594 -6580
rect 35356 -6614 35372 -6597
rect 35120 -6630 35372 -6614
rect 35578 -6614 35594 -6597
rect 35814 -6597 35904 -6580
rect 35962 -6580 36362 -6542
rect 35962 -6597 36052 -6580
rect 35814 -6614 35830 -6597
rect 35578 -6630 35830 -6614
rect 36036 -6614 36052 -6597
rect 36272 -6597 36362 -6580
rect 36420 -6580 36820 -6542
rect 36420 -6597 36510 -6580
rect 36272 -6614 36288 -6597
rect 36036 -6630 36288 -6614
rect 36494 -6614 36510 -6597
rect 36730 -6597 36820 -6580
rect 36878 -6580 37278 -6542
rect 36878 -6597 36968 -6580
rect 36730 -6614 36746 -6597
rect 36494 -6630 36746 -6614
rect 36952 -6614 36968 -6597
rect 37188 -6597 37278 -6580
rect 37188 -6614 37204 -6597
rect 36952 -6630 37204 -6614
rect 12829 -7754 13081 -7738
rect 12829 -7771 12845 -7754
rect 12755 -7788 12845 -7771
rect 13065 -7771 13081 -7754
rect 13287 -7754 13539 -7738
rect 13287 -7771 13303 -7754
rect 13065 -7788 13155 -7771
rect 12755 -7835 13155 -7788
rect 13213 -7788 13303 -7771
rect 13523 -7771 13539 -7754
rect 13745 -7754 13997 -7738
rect 13745 -7771 13761 -7754
rect 13523 -7788 13613 -7771
rect 13213 -7835 13613 -7788
rect 13671 -7788 13761 -7771
rect 13981 -7771 13997 -7754
rect 14203 -7754 14455 -7738
rect 14203 -7771 14219 -7754
rect 13981 -7788 14071 -7771
rect 13671 -7835 14071 -7788
rect 14129 -7788 14219 -7771
rect 14439 -7771 14455 -7754
rect 14661 -7754 14913 -7738
rect 14661 -7771 14677 -7754
rect 14439 -7788 14529 -7771
rect 14129 -7835 14529 -7788
rect 14587 -7788 14677 -7771
rect 14897 -7771 14913 -7754
rect 15119 -7754 15371 -7738
rect 15119 -7771 15135 -7754
rect 14897 -7788 14987 -7771
rect 14587 -7835 14987 -7788
rect 15045 -7788 15135 -7771
rect 15355 -7771 15371 -7754
rect 15577 -7754 15829 -7738
rect 15577 -7771 15593 -7754
rect 15355 -7788 15445 -7771
rect 15045 -7835 15445 -7788
rect 15503 -7788 15593 -7771
rect 15813 -7771 15829 -7754
rect 16035 -7754 16287 -7738
rect 16035 -7771 16051 -7754
rect 15813 -7788 15903 -7771
rect 15503 -7835 15903 -7788
rect 15961 -7788 16051 -7771
rect 16271 -7771 16287 -7754
rect 16493 -7754 16745 -7738
rect 16493 -7771 16509 -7754
rect 16271 -7788 16361 -7771
rect 15961 -7835 16361 -7788
rect 16419 -7788 16509 -7771
rect 16729 -7771 16745 -7754
rect 16951 -7754 17203 -7738
rect 16951 -7771 16967 -7754
rect 16729 -7788 16819 -7771
rect 16419 -7835 16819 -7788
rect 16877 -7788 16967 -7771
rect 17187 -7771 17203 -7754
rect 17829 -7754 18081 -7738
rect 17829 -7771 17845 -7754
rect 17187 -7788 17277 -7771
rect 16877 -7835 17277 -7788
rect 17755 -7788 17845 -7771
rect 18065 -7771 18081 -7754
rect 18287 -7754 18539 -7738
rect 18287 -7771 18303 -7754
rect 18065 -7788 18155 -7771
rect 17755 -7835 18155 -7788
rect 18213 -7788 18303 -7771
rect 18523 -7771 18539 -7754
rect 18745 -7754 18997 -7738
rect 18745 -7771 18761 -7754
rect 18523 -7788 18613 -7771
rect 18213 -7835 18613 -7788
rect 18671 -7788 18761 -7771
rect 18981 -7771 18997 -7754
rect 19203 -7754 19455 -7738
rect 19203 -7771 19219 -7754
rect 18981 -7788 19071 -7771
rect 18671 -7835 19071 -7788
rect 19129 -7788 19219 -7771
rect 19439 -7771 19455 -7754
rect 19661 -7754 19913 -7738
rect 19661 -7771 19677 -7754
rect 19439 -7788 19529 -7771
rect 19129 -7835 19529 -7788
rect 19587 -7788 19677 -7771
rect 19897 -7771 19913 -7754
rect 20119 -7754 20371 -7738
rect 20119 -7771 20135 -7754
rect 19897 -7788 19987 -7771
rect 19587 -7835 19987 -7788
rect 20045 -7788 20135 -7771
rect 20355 -7771 20371 -7754
rect 20577 -7754 20829 -7738
rect 20577 -7771 20593 -7754
rect 20355 -7788 20445 -7771
rect 20045 -7835 20445 -7788
rect 20503 -7788 20593 -7771
rect 20813 -7771 20829 -7754
rect 21035 -7754 21287 -7738
rect 21035 -7771 21051 -7754
rect 20813 -7788 20903 -7771
rect 20503 -7835 20903 -7788
rect 20961 -7788 21051 -7771
rect 21271 -7771 21287 -7754
rect 21493 -7754 21745 -7738
rect 21493 -7771 21509 -7754
rect 21271 -7788 21361 -7771
rect 20961 -7835 21361 -7788
rect 21419 -7788 21509 -7771
rect 21729 -7771 21745 -7754
rect 21951 -7754 22203 -7738
rect 21951 -7771 21967 -7754
rect 21729 -7788 21819 -7771
rect 21419 -7835 21819 -7788
rect 21877 -7788 21967 -7771
rect 22187 -7771 22203 -7754
rect 22187 -7788 22277 -7771
rect 21877 -7835 22277 -7788
rect 12755 -9082 13155 -9035
rect 12755 -9099 12845 -9082
rect 12829 -9116 12845 -9099
rect 13065 -9099 13155 -9082
rect 13213 -9082 13613 -9035
rect 13213 -9099 13303 -9082
rect 13065 -9116 13081 -9099
rect 12829 -9132 13081 -9116
rect 13287 -9116 13303 -9099
rect 13523 -9099 13613 -9082
rect 13671 -9082 14071 -9035
rect 13671 -9099 13761 -9082
rect 13523 -9116 13539 -9099
rect 13287 -9132 13539 -9116
rect 13745 -9116 13761 -9099
rect 13981 -9099 14071 -9082
rect 14129 -9082 14529 -9035
rect 14129 -9099 14219 -9082
rect 13981 -9116 13997 -9099
rect 13745 -9132 13997 -9116
rect 14203 -9116 14219 -9099
rect 14439 -9099 14529 -9082
rect 14587 -9082 14987 -9035
rect 14587 -9099 14677 -9082
rect 14439 -9116 14455 -9099
rect 14203 -9132 14455 -9116
rect 14661 -9116 14677 -9099
rect 14897 -9099 14987 -9082
rect 15045 -9082 15445 -9035
rect 15045 -9099 15135 -9082
rect 14897 -9116 14913 -9099
rect 14661 -9132 14913 -9116
rect 15119 -9116 15135 -9099
rect 15355 -9099 15445 -9082
rect 15503 -9082 15903 -9035
rect 15503 -9099 15593 -9082
rect 15355 -9116 15371 -9099
rect 15119 -9132 15371 -9116
rect 15577 -9116 15593 -9099
rect 15813 -9099 15903 -9082
rect 15961 -9082 16361 -9035
rect 15961 -9099 16051 -9082
rect 15813 -9116 15829 -9099
rect 15577 -9132 15829 -9116
rect 16035 -9116 16051 -9099
rect 16271 -9099 16361 -9082
rect 16419 -9082 16819 -9035
rect 16419 -9099 16509 -9082
rect 16271 -9116 16287 -9099
rect 16035 -9132 16287 -9116
rect 16493 -9116 16509 -9099
rect 16729 -9099 16819 -9082
rect 16877 -9082 17277 -9035
rect 16877 -9099 16967 -9082
rect 16729 -9116 16745 -9099
rect 16493 -9132 16745 -9116
rect 16951 -9116 16967 -9099
rect 17187 -9099 17277 -9082
rect 17755 -9082 18155 -9035
rect 17755 -9099 17845 -9082
rect 17187 -9116 17203 -9099
rect 16951 -9132 17203 -9116
rect 17829 -9116 17845 -9099
rect 18065 -9099 18155 -9082
rect 18213 -9082 18613 -9035
rect 18213 -9099 18303 -9082
rect 18065 -9116 18081 -9099
rect 17829 -9132 18081 -9116
rect 18287 -9116 18303 -9099
rect 18523 -9099 18613 -9082
rect 18671 -9082 19071 -9035
rect 18671 -9099 18761 -9082
rect 18523 -9116 18539 -9099
rect 18287 -9132 18539 -9116
rect 18745 -9116 18761 -9099
rect 18981 -9099 19071 -9082
rect 19129 -9082 19529 -9035
rect 19129 -9099 19219 -9082
rect 18981 -9116 18997 -9099
rect 18745 -9132 18997 -9116
rect 19203 -9116 19219 -9099
rect 19439 -9099 19529 -9082
rect 19587 -9082 19987 -9035
rect 19587 -9099 19677 -9082
rect 19439 -9116 19455 -9099
rect 19203 -9132 19455 -9116
rect 19661 -9116 19677 -9099
rect 19897 -9099 19987 -9082
rect 20045 -9082 20445 -9035
rect 20045 -9099 20135 -9082
rect 19897 -9116 19913 -9099
rect 19661 -9132 19913 -9116
rect 20119 -9116 20135 -9099
rect 20355 -9099 20445 -9082
rect 20503 -9082 20903 -9035
rect 20503 -9099 20593 -9082
rect 20355 -9116 20371 -9099
rect 20119 -9132 20371 -9116
rect 20577 -9116 20593 -9099
rect 20813 -9099 20903 -9082
rect 20961 -9082 21361 -9035
rect 20961 -9099 21051 -9082
rect 20813 -9116 20829 -9099
rect 20577 -9132 20829 -9116
rect 21035 -9116 21051 -9099
rect 21271 -9099 21361 -9082
rect 21419 -9082 21819 -9035
rect 21419 -9099 21509 -9082
rect 21271 -9116 21287 -9099
rect 21035 -9132 21287 -9116
rect 21493 -9116 21509 -9099
rect 21729 -9099 21819 -9082
rect 21877 -9082 22277 -9035
rect 21877 -9099 21967 -9082
rect 21729 -9116 21745 -9099
rect 21493 -9132 21745 -9116
rect 21951 -9116 21967 -9099
rect 22187 -9099 22277 -9082
rect 22187 -9116 22203 -9099
rect 21951 -9132 22203 -9116
rect 13606 -10019 13858 -10003
rect 13606 -10036 13622 -10019
rect 13532 -10053 13622 -10036
rect 13842 -10036 13858 -10019
rect 14064 -10019 14316 -10003
rect 14064 -10036 14080 -10019
rect 13842 -10053 13932 -10036
rect 13532 -10100 13932 -10053
rect 13990 -10053 14080 -10036
rect 14300 -10036 14316 -10019
rect 14522 -10019 14774 -10003
rect 14522 -10036 14538 -10019
rect 14300 -10053 14390 -10036
rect 13990 -10100 14390 -10053
rect 14448 -10053 14538 -10036
rect 14758 -10036 14774 -10019
rect 14980 -10019 15232 -10003
rect 14980 -10036 14996 -10019
rect 14758 -10053 14848 -10036
rect 14448 -10100 14848 -10053
rect 14906 -10053 14996 -10036
rect 15216 -10036 15232 -10019
rect 15438 -10019 15690 -10003
rect 15438 -10036 15454 -10019
rect 15216 -10053 15306 -10036
rect 14906 -10100 15306 -10053
rect 15364 -10053 15454 -10036
rect 15674 -10036 15690 -10019
rect 15896 -10019 16148 -10003
rect 15896 -10036 15912 -10019
rect 15674 -10053 15764 -10036
rect 15364 -10100 15764 -10053
rect 15822 -10053 15912 -10036
rect 16132 -10036 16148 -10019
rect 16354 -10019 16606 -10003
rect 16354 -10036 16370 -10019
rect 16132 -10053 16222 -10036
rect 15822 -10100 16222 -10053
rect 16280 -10053 16370 -10036
rect 16590 -10036 16606 -10019
rect 16812 -10019 17064 -10003
rect 16812 -10036 16828 -10019
rect 16590 -10053 16680 -10036
rect 16280 -10100 16680 -10053
rect 16738 -10053 16828 -10036
rect 17048 -10036 17064 -10019
rect 17270 -10019 17522 -10003
rect 17270 -10036 17286 -10019
rect 17048 -10053 17138 -10036
rect 16738 -10100 17138 -10053
rect 17196 -10053 17286 -10036
rect 17506 -10036 17522 -10019
rect 17728 -10019 17980 -10003
rect 17728 -10036 17744 -10019
rect 17506 -10053 17596 -10036
rect 17196 -10100 17596 -10053
rect 17654 -10053 17744 -10036
rect 17964 -10036 17980 -10019
rect 18186 -10019 18438 -10003
rect 18186 -10036 18202 -10019
rect 17964 -10053 18054 -10036
rect 17654 -10100 18054 -10053
rect 18112 -10053 18202 -10036
rect 18422 -10036 18438 -10019
rect 18644 -10019 18896 -10003
rect 18644 -10036 18660 -10019
rect 18422 -10053 18512 -10036
rect 18112 -10100 18512 -10053
rect 18570 -10053 18660 -10036
rect 18880 -10036 18896 -10019
rect 19102 -10019 19354 -10003
rect 19102 -10036 19118 -10019
rect 18880 -10053 18970 -10036
rect 18570 -10100 18970 -10053
rect 19028 -10053 19118 -10036
rect 19338 -10036 19354 -10019
rect 19560 -10019 19812 -10003
rect 19560 -10036 19576 -10019
rect 19338 -10053 19428 -10036
rect 19028 -10100 19428 -10053
rect 19486 -10053 19576 -10036
rect 19796 -10036 19812 -10019
rect 20018 -10019 20270 -10003
rect 20018 -10036 20034 -10019
rect 19796 -10053 19886 -10036
rect 19486 -10100 19886 -10053
rect 19944 -10053 20034 -10036
rect 20254 -10036 20270 -10019
rect 20476 -10019 20728 -10003
rect 20476 -10036 20492 -10019
rect 20254 -10053 20344 -10036
rect 19944 -10100 20344 -10053
rect 20402 -10053 20492 -10036
rect 20712 -10036 20728 -10019
rect 20934 -10019 21186 -10003
rect 20934 -10036 20950 -10019
rect 20712 -10053 20802 -10036
rect 20402 -10100 20802 -10053
rect 20860 -10053 20950 -10036
rect 21170 -10036 21186 -10019
rect 21392 -10019 21644 -10003
rect 21392 -10036 21408 -10019
rect 21170 -10053 21260 -10036
rect 20860 -10100 21260 -10053
rect 21318 -10053 21408 -10036
rect 21628 -10036 21644 -10019
rect 21628 -10053 21718 -10036
rect 21318 -10100 21718 -10053
rect 13532 -11747 13932 -11700
rect 13532 -11764 13622 -11747
rect 13606 -11781 13622 -11764
rect 13842 -11764 13932 -11747
rect 13990 -11747 14390 -11700
rect 13990 -11764 14080 -11747
rect 13842 -11781 13858 -11764
rect 13606 -11797 13858 -11781
rect 14064 -11781 14080 -11764
rect 14300 -11764 14390 -11747
rect 14448 -11747 14848 -11700
rect 14448 -11764 14538 -11747
rect 14300 -11781 14316 -11764
rect 14064 -11797 14316 -11781
rect 14522 -11781 14538 -11764
rect 14758 -11764 14848 -11747
rect 14906 -11747 15306 -11700
rect 14906 -11764 14996 -11747
rect 14758 -11781 14774 -11764
rect 14522 -11797 14774 -11781
rect 14980 -11781 14996 -11764
rect 15216 -11764 15306 -11747
rect 15364 -11747 15764 -11700
rect 15364 -11764 15454 -11747
rect 15216 -11781 15232 -11764
rect 14980 -11797 15232 -11781
rect 15438 -11781 15454 -11764
rect 15674 -11764 15764 -11747
rect 15822 -11747 16222 -11700
rect 15822 -11764 15912 -11747
rect 15674 -11781 15690 -11764
rect 15438 -11797 15690 -11781
rect 15896 -11781 15912 -11764
rect 16132 -11764 16222 -11747
rect 16280 -11747 16680 -11700
rect 16280 -11764 16370 -11747
rect 16132 -11781 16148 -11764
rect 15896 -11797 16148 -11781
rect 16354 -11781 16370 -11764
rect 16590 -11764 16680 -11747
rect 16738 -11747 17138 -11700
rect 16738 -11764 16828 -11747
rect 16590 -11781 16606 -11764
rect 16354 -11797 16606 -11781
rect 16812 -11781 16828 -11764
rect 17048 -11764 17138 -11747
rect 17196 -11747 17596 -11700
rect 17196 -11764 17286 -11747
rect 17048 -11781 17064 -11764
rect 16812 -11797 17064 -11781
rect 17270 -11781 17286 -11764
rect 17506 -11764 17596 -11747
rect 17654 -11747 18054 -11700
rect 17654 -11764 17744 -11747
rect 17506 -11781 17522 -11764
rect 17270 -11797 17522 -11781
rect 17728 -11781 17744 -11764
rect 17964 -11764 18054 -11747
rect 18112 -11747 18512 -11700
rect 18112 -11764 18202 -11747
rect 17964 -11781 17980 -11764
rect 17728 -11797 17980 -11781
rect 18186 -11781 18202 -11764
rect 18422 -11764 18512 -11747
rect 18570 -11747 18970 -11700
rect 18570 -11764 18660 -11747
rect 18422 -11781 18438 -11764
rect 18186 -11797 18438 -11781
rect 18644 -11781 18660 -11764
rect 18880 -11764 18970 -11747
rect 19028 -11747 19428 -11700
rect 19028 -11764 19118 -11747
rect 18880 -11781 18896 -11764
rect 18644 -11797 18896 -11781
rect 19102 -11781 19118 -11764
rect 19338 -11764 19428 -11747
rect 19486 -11747 19886 -11700
rect 19486 -11764 19576 -11747
rect 19338 -11781 19354 -11764
rect 19102 -11797 19354 -11781
rect 19560 -11781 19576 -11764
rect 19796 -11764 19886 -11747
rect 19944 -11747 20344 -11700
rect 19944 -11764 20034 -11747
rect 19796 -11781 19812 -11764
rect 19560 -11797 19812 -11781
rect 20018 -11781 20034 -11764
rect 20254 -11764 20344 -11747
rect 20402 -11747 20802 -11700
rect 20402 -11764 20492 -11747
rect 20254 -11781 20270 -11764
rect 20018 -11797 20270 -11781
rect 20476 -11781 20492 -11764
rect 20712 -11764 20802 -11747
rect 20860 -11747 21260 -11700
rect 20860 -11764 20950 -11747
rect 20712 -11781 20728 -11764
rect 20476 -11797 20728 -11781
rect 20934 -11781 20950 -11764
rect 21170 -11764 21260 -11747
rect 21318 -11747 21718 -11700
rect 21318 -11764 21408 -11747
rect 21170 -11781 21186 -11764
rect 20934 -11797 21186 -11781
rect 21392 -11781 21408 -11764
rect 21628 -11764 21718 -11747
rect 21628 -11781 21644 -11764
rect 21392 -11797 21644 -11781
rect 27829 -7754 28081 -7738
rect 27829 -7771 27845 -7754
rect 27755 -7788 27845 -7771
rect 28065 -7771 28081 -7754
rect 28287 -7754 28539 -7738
rect 28287 -7771 28303 -7754
rect 28065 -7788 28155 -7771
rect 27755 -7835 28155 -7788
rect 28213 -7788 28303 -7771
rect 28523 -7771 28539 -7754
rect 28745 -7754 28997 -7738
rect 28745 -7771 28761 -7754
rect 28523 -7788 28613 -7771
rect 28213 -7835 28613 -7788
rect 28671 -7788 28761 -7771
rect 28981 -7771 28997 -7754
rect 29203 -7754 29455 -7738
rect 29203 -7771 29219 -7754
rect 28981 -7788 29071 -7771
rect 28671 -7835 29071 -7788
rect 29129 -7788 29219 -7771
rect 29439 -7771 29455 -7754
rect 29661 -7754 29913 -7738
rect 29661 -7771 29677 -7754
rect 29439 -7788 29529 -7771
rect 29129 -7835 29529 -7788
rect 29587 -7788 29677 -7771
rect 29897 -7771 29913 -7754
rect 30119 -7754 30371 -7738
rect 30119 -7771 30135 -7754
rect 29897 -7788 29987 -7771
rect 29587 -7835 29987 -7788
rect 30045 -7788 30135 -7771
rect 30355 -7771 30371 -7754
rect 30577 -7754 30829 -7738
rect 30577 -7771 30593 -7754
rect 30355 -7788 30445 -7771
rect 30045 -7835 30445 -7788
rect 30503 -7788 30593 -7771
rect 30813 -7771 30829 -7754
rect 31035 -7754 31287 -7738
rect 31035 -7771 31051 -7754
rect 30813 -7788 30903 -7771
rect 30503 -7835 30903 -7788
rect 30961 -7788 31051 -7771
rect 31271 -7771 31287 -7754
rect 31493 -7754 31745 -7738
rect 31493 -7771 31509 -7754
rect 31271 -7788 31361 -7771
rect 30961 -7835 31361 -7788
rect 31419 -7788 31509 -7771
rect 31729 -7771 31745 -7754
rect 31951 -7754 32203 -7738
rect 31951 -7771 31967 -7754
rect 31729 -7788 31819 -7771
rect 31419 -7835 31819 -7788
rect 31877 -7788 31967 -7771
rect 32187 -7771 32203 -7754
rect 32829 -7754 33081 -7738
rect 32829 -7771 32845 -7754
rect 32187 -7788 32277 -7771
rect 31877 -7835 32277 -7788
rect 32755 -7788 32845 -7771
rect 33065 -7771 33081 -7754
rect 33287 -7754 33539 -7738
rect 33287 -7771 33303 -7754
rect 33065 -7788 33155 -7771
rect 32755 -7835 33155 -7788
rect 33213 -7788 33303 -7771
rect 33523 -7771 33539 -7754
rect 33745 -7754 33997 -7738
rect 33745 -7771 33761 -7754
rect 33523 -7788 33613 -7771
rect 33213 -7835 33613 -7788
rect 33671 -7788 33761 -7771
rect 33981 -7771 33997 -7754
rect 34203 -7754 34455 -7738
rect 34203 -7771 34219 -7754
rect 33981 -7788 34071 -7771
rect 33671 -7835 34071 -7788
rect 34129 -7788 34219 -7771
rect 34439 -7771 34455 -7754
rect 34661 -7754 34913 -7738
rect 34661 -7771 34677 -7754
rect 34439 -7788 34529 -7771
rect 34129 -7835 34529 -7788
rect 34587 -7788 34677 -7771
rect 34897 -7771 34913 -7754
rect 35119 -7754 35371 -7738
rect 35119 -7771 35135 -7754
rect 34897 -7788 34987 -7771
rect 34587 -7835 34987 -7788
rect 35045 -7788 35135 -7771
rect 35355 -7771 35371 -7754
rect 35577 -7754 35829 -7738
rect 35577 -7771 35593 -7754
rect 35355 -7788 35445 -7771
rect 35045 -7835 35445 -7788
rect 35503 -7788 35593 -7771
rect 35813 -7771 35829 -7754
rect 36035 -7754 36287 -7738
rect 36035 -7771 36051 -7754
rect 35813 -7788 35903 -7771
rect 35503 -7835 35903 -7788
rect 35961 -7788 36051 -7771
rect 36271 -7771 36287 -7754
rect 36493 -7754 36745 -7738
rect 36493 -7771 36509 -7754
rect 36271 -7788 36361 -7771
rect 35961 -7835 36361 -7788
rect 36419 -7788 36509 -7771
rect 36729 -7771 36745 -7754
rect 36951 -7754 37203 -7738
rect 36951 -7771 36967 -7754
rect 36729 -7788 36819 -7771
rect 36419 -7835 36819 -7788
rect 36877 -7788 36967 -7771
rect 37187 -7771 37203 -7754
rect 37187 -7788 37277 -7771
rect 36877 -7835 37277 -7788
rect 27755 -9082 28155 -9035
rect 27755 -9099 27845 -9082
rect 27829 -9116 27845 -9099
rect 28065 -9099 28155 -9082
rect 28213 -9082 28613 -9035
rect 28213 -9099 28303 -9082
rect 28065 -9116 28081 -9099
rect 27829 -9132 28081 -9116
rect 28287 -9116 28303 -9099
rect 28523 -9099 28613 -9082
rect 28671 -9082 29071 -9035
rect 28671 -9099 28761 -9082
rect 28523 -9116 28539 -9099
rect 28287 -9132 28539 -9116
rect 28745 -9116 28761 -9099
rect 28981 -9099 29071 -9082
rect 29129 -9082 29529 -9035
rect 29129 -9099 29219 -9082
rect 28981 -9116 28997 -9099
rect 28745 -9132 28997 -9116
rect 29203 -9116 29219 -9099
rect 29439 -9099 29529 -9082
rect 29587 -9082 29987 -9035
rect 29587 -9099 29677 -9082
rect 29439 -9116 29455 -9099
rect 29203 -9132 29455 -9116
rect 29661 -9116 29677 -9099
rect 29897 -9099 29987 -9082
rect 30045 -9082 30445 -9035
rect 30045 -9099 30135 -9082
rect 29897 -9116 29913 -9099
rect 29661 -9132 29913 -9116
rect 30119 -9116 30135 -9099
rect 30355 -9099 30445 -9082
rect 30503 -9082 30903 -9035
rect 30503 -9099 30593 -9082
rect 30355 -9116 30371 -9099
rect 30119 -9132 30371 -9116
rect 30577 -9116 30593 -9099
rect 30813 -9099 30903 -9082
rect 30961 -9082 31361 -9035
rect 30961 -9099 31051 -9082
rect 30813 -9116 30829 -9099
rect 30577 -9132 30829 -9116
rect 31035 -9116 31051 -9099
rect 31271 -9099 31361 -9082
rect 31419 -9082 31819 -9035
rect 31419 -9099 31509 -9082
rect 31271 -9116 31287 -9099
rect 31035 -9132 31287 -9116
rect 31493 -9116 31509 -9099
rect 31729 -9099 31819 -9082
rect 31877 -9082 32277 -9035
rect 31877 -9099 31967 -9082
rect 31729 -9116 31745 -9099
rect 31493 -9132 31745 -9116
rect 31951 -9116 31967 -9099
rect 32187 -9099 32277 -9082
rect 32755 -9082 33155 -9035
rect 32755 -9099 32845 -9082
rect 32187 -9116 32203 -9099
rect 31951 -9132 32203 -9116
rect 32829 -9116 32845 -9099
rect 33065 -9099 33155 -9082
rect 33213 -9082 33613 -9035
rect 33213 -9099 33303 -9082
rect 33065 -9116 33081 -9099
rect 32829 -9132 33081 -9116
rect 33287 -9116 33303 -9099
rect 33523 -9099 33613 -9082
rect 33671 -9082 34071 -9035
rect 33671 -9099 33761 -9082
rect 33523 -9116 33539 -9099
rect 33287 -9132 33539 -9116
rect 33745 -9116 33761 -9099
rect 33981 -9099 34071 -9082
rect 34129 -9082 34529 -9035
rect 34129 -9099 34219 -9082
rect 33981 -9116 33997 -9099
rect 33745 -9132 33997 -9116
rect 34203 -9116 34219 -9099
rect 34439 -9099 34529 -9082
rect 34587 -9082 34987 -9035
rect 34587 -9099 34677 -9082
rect 34439 -9116 34455 -9099
rect 34203 -9132 34455 -9116
rect 34661 -9116 34677 -9099
rect 34897 -9099 34987 -9082
rect 35045 -9082 35445 -9035
rect 35045 -9099 35135 -9082
rect 34897 -9116 34913 -9099
rect 34661 -9132 34913 -9116
rect 35119 -9116 35135 -9099
rect 35355 -9099 35445 -9082
rect 35503 -9082 35903 -9035
rect 35503 -9099 35593 -9082
rect 35355 -9116 35371 -9099
rect 35119 -9132 35371 -9116
rect 35577 -9116 35593 -9099
rect 35813 -9099 35903 -9082
rect 35961 -9082 36361 -9035
rect 35961 -9099 36051 -9082
rect 35813 -9116 35829 -9099
rect 35577 -9132 35829 -9116
rect 36035 -9116 36051 -9099
rect 36271 -9099 36361 -9082
rect 36419 -9082 36819 -9035
rect 36419 -9099 36509 -9082
rect 36271 -9116 36287 -9099
rect 36035 -9132 36287 -9116
rect 36493 -9116 36509 -9099
rect 36729 -9099 36819 -9082
rect 36877 -9082 37277 -9035
rect 36877 -9099 36967 -9082
rect 36729 -9116 36745 -9099
rect 36493 -9132 36745 -9116
rect 36951 -9116 36967 -9099
rect 37187 -9099 37277 -9082
rect 37187 -9116 37203 -9099
rect 36951 -9132 37203 -9116
rect 28606 -10019 28858 -10003
rect 28606 -10036 28622 -10019
rect 28532 -10053 28622 -10036
rect 28842 -10036 28858 -10019
rect 29064 -10019 29316 -10003
rect 29064 -10036 29080 -10019
rect 28842 -10053 28932 -10036
rect 28532 -10100 28932 -10053
rect 28990 -10053 29080 -10036
rect 29300 -10036 29316 -10019
rect 29522 -10019 29774 -10003
rect 29522 -10036 29538 -10019
rect 29300 -10053 29390 -10036
rect 28990 -10100 29390 -10053
rect 29448 -10053 29538 -10036
rect 29758 -10036 29774 -10019
rect 29980 -10019 30232 -10003
rect 29980 -10036 29996 -10019
rect 29758 -10053 29848 -10036
rect 29448 -10100 29848 -10053
rect 29906 -10053 29996 -10036
rect 30216 -10036 30232 -10019
rect 30438 -10019 30690 -10003
rect 30438 -10036 30454 -10019
rect 30216 -10053 30306 -10036
rect 29906 -10100 30306 -10053
rect 30364 -10053 30454 -10036
rect 30674 -10036 30690 -10019
rect 30896 -10019 31148 -10003
rect 30896 -10036 30912 -10019
rect 30674 -10053 30764 -10036
rect 30364 -10100 30764 -10053
rect 30822 -10053 30912 -10036
rect 31132 -10036 31148 -10019
rect 31354 -10019 31606 -10003
rect 31354 -10036 31370 -10019
rect 31132 -10053 31222 -10036
rect 30822 -10100 31222 -10053
rect 31280 -10053 31370 -10036
rect 31590 -10036 31606 -10019
rect 31812 -10019 32064 -10003
rect 31812 -10036 31828 -10019
rect 31590 -10053 31680 -10036
rect 31280 -10100 31680 -10053
rect 31738 -10053 31828 -10036
rect 32048 -10036 32064 -10019
rect 32270 -10019 32522 -10003
rect 32270 -10036 32286 -10019
rect 32048 -10053 32138 -10036
rect 31738 -10100 32138 -10053
rect 32196 -10053 32286 -10036
rect 32506 -10036 32522 -10019
rect 32728 -10019 32980 -10003
rect 32728 -10036 32744 -10019
rect 32506 -10053 32596 -10036
rect 32196 -10100 32596 -10053
rect 32654 -10053 32744 -10036
rect 32964 -10036 32980 -10019
rect 33186 -10019 33438 -10003
rect 33186 -10036 33202 -10019
rect 32964 -10053 33054 -10036
rect 32654 -10100 33054 -10053
rect 33112 -10053 33202 -10036
rect 33422 -10036 33438 -10019
rect 33644 -10019 33896 -10003
rect 33644 -10036 33660 -10019
rect 33422 -10053 33512 -10036
rect 33112 -10100 33512 -10053
rect 33570 -10053 33660 -10036
rect 33880 -10036 33896 -10019
rect 34102 -10019 34354 -10003
rect 34102 -10036 34118 -10019
rect 33880 -10053 33970 -10036
rect 33570 -10100 33970 -10053
rect 34028 -10053 34118 -10036
rect 34338 -10036 34354 -10019
rect 34560 -10019 34812 -10003
rect 34560 -10036 34576 -10019
rect 34338 -10053 34428 -10036
rect 34028 -10100 34428 -10053
rect 34486 -10053 34576 -10036
rect 34796 -10036 34812 -10019
rect 35018 -10019 35270 -10003
rect 35018 -10036 35034 -10019
rect 34796 -10053 34886 -10036
rect 34486 -10100 34886 -10053
rect 34944 -10053 35034 -10036
rect 35254 -10036 35270 -10019
rect 35476 -10019 35728 -10003
rect 35476 -10036 35492 -10019
rect 35254 -10053 35344 -10036
rect 34944 -10100 35344 -10053
rect 35402 -10053 35492 -10036
rect 35712 -10036 35728 -10019
rect 35934 -10019 36186 -10003
rect 35934 -10036 35950 -10019
rect 35712 -10053 35802 -10036
rect 35402 -10100 35802 -10053
rect 35860 -10053 35950 -10036
rect 36170 -10036 36186 -10019
rect 36392 -10019 36644 -10003
rect 36392 -10036 36408 -10019
rect 36170 -10053 36260 -10036
rect 35860 -10100 36260 -10053
rect 36318 -10053 36408 -10036
rect 36628 -10036 36644 -10019
rect 36628 -10053 36718 -10036
rect 36318 -10100 36718 -10053
rect 28532 -11747 28932 -11700
rect 28532 -11764 28622 -11747
rect 28606 -11781 28622 -11764
rect 28842 -11764 28932 -11747
rect 28990 -11747 29390 -11700
rect 28990 -11764 29080 -11747
rect 28842 -11781 28858 -11764
rect 28606 -11797 28858 -11781
rect 29064 -11781 29080 -11764
rect 29300 -11764 29390 -11747
rect 29448 -11747 29848 -11700
rect 29448 -11764 29538 -11747
rect 29300 -11781 29316 -11764
rect 29064 -11797 29316 -11781
rect 29522 -11781 29538 -11764
rect 29758 -11764 29848 -11747
rect 29906 -11747 30306 -11700
rect 29906 -11764 29996 -11747
rect 29758 -11781 29774 -11764
rect 29522 -11797 29774 -11781
rect 29980 -11781 29996 -11764
rect 30216 -11764 30306 -11747
rect 30364 -11747 30764 -11700
rect 30364 -11764 30454 -11747
rect 30216 -11781 30232 -11764
rect 29980 -11797 30232 -11781
rect 30438 -11781 30454 -11764
rect 30674 -11764 30764 -11747
rect 30822 -11747 31222 -11700
rect 30822 -11764 30912 -11747
rect 30674 -11781 30690 -11764
rect 30438 -11797 30690 -11781
rect 30896 -11781 30912 -11764
rect 31132 -11764 31222 -11747
rect 31280 -11747 31680 -11700
rect 31280 -11764 31370 -11747
rect 31132 -11781 31148 -11764
rect 30896 -11797 31148 -11781
rect 31354 -11781 31370 -11764
rect 31590 -11764 31680 -11747
rect 31738 -11747 32138 -11700
rect 31738 -11764 31828 -11747
rect 31590 -11781 31606 -11764
rect 31354 -11797 31606 -11781
rect 31812 -11781 31828 -11764
rect 32048 -11764 32138 -11747
rect 32196 -11747 32596 -11700
rect 32196 -11764 32286 -11747
rect 32048 -11781 32064 -11764
rect 31812 -11797 32064 -11781
rect 32270 -11781 32286 -11764
rect 32506 -11764 32596 -11747
rect 32654 -11747 33054 -11700
rect 32654 -11764 32744 -11747
rect 32506 -11781 32522 -11764
rect 32270 -11797 32522 -11781
rect 32728 -11781 32744 -11764
rect 32964 -11764 33054 -11747
rect 33112 -11747 33512 -11700
rect 33112 -11764 33202 -11747
rect 32964 -11781 32980 -11764
rect 32728 -11797 32980 -11781
rect 33186 -11781 33202 -11764
rect 33422 -11764 33512 -11747
rect 33570 -11747 33970 -11700
rect 33570 -11764 33660 -11747
rect 33422 -11781 33438 -11764
rect 33186 -11797 33438 -11781
rect 33644 -11781 33660 -11764
rect 33880 -11764 33970 -11747
rect 34028 -11747 34428 -11700
rect 34028 -11764 34118 -11747
rect 33880 -11781 33896 -11764
rect 33644 -11797 33896 -11781
rect 34102 -11781 34118 -11764
rect 34338 -11764 34428 -11747
rect 34486 -11747 34886 -11700
rect 34486 -11764 34576 -11747
rect 34338 -11781 34354 -11764
rect 34102 -11797 34354 -11781
rect 34560 -11781 34576 -11764
rect 34796 -11764 34886 -11747
rect 34944 -11747 35344 -11700
rect 34944 -11764 35034 -11747
rect 34796 -11781 34812 -11764
rect 34560 -11797 34812 -11781
rect 35018 -11781 35034 -11764
rect 35254 -11764 35344 -11747
rect 35402 -11747 35802 -11700
rect 35402 -11764 35492 -11747
rect 35254 -11781 35270 -11764
rect 35018 -11797 35270 -11781
rect 35476 -11781 35492 -11764
rect 35712 -11764 35802 -11747
rect 35860 -11747 36260 -11700
rect 35860 -11764 35950 -11747
rect 35712 -11781 35728 -11764
rect 35476 -11797 35728 -11781
rect 35934 -11781 35950 -11764
rect 36170 -11764 36260 -11747
rect 36318 -11747 36718 -11700
rect 36318 -11764 36408 -11747
rect 36170 -11781 36186 -11764
rect 35934 -11797 36186 -11781
rect 36392 -11781 36408 -11764
rect 36628 -11764 36718 -11747
rect 36628 -11781 36644 -11764
rect 36392 -11797 36644 -11781
rect 9458 -14975 9710 -14959
rect 9458 -14992 9474 -14975
rect 9384 -15009 9474 -14992
rect 9694 -14992 9710 -14975
rect 9916 -14975 10168 -14959
rect 9916 -14992 9932 -14975
rect 9694 -15009 9784 -14992
rect 9384 -15056 9784 -15009
rect 9842 -15009 9932 -14992
rect 10152 -14992 10168 -14975
rect 10374 -14975 10626 -14959
rect 10374 -14992 10390 -14975
rect 10152 -15009 10242 -14992
rect 9842 -15056 10242 -15009
rect 10300 -15009 10390 -14992
rect 10610 -14992 10626 -14975
rect 10832 -14975 11084 -14959
rect 10832 -14992 10848 -14975
rect 10610 -15009 10700 -14992
rect 10300 -15056 10700 -15009
rect 10758 -15009 10848 -14992
rect 11068 -14992 11084 -14975
rect 11290 -14975 11542 -14959
rect 11290 -14992 11306 -14975
rect 11068 -15009 11158 -14992
rect 10758 -15056 11158 -15009
rect 11216 -15009 11306 -14992
rect 11526 -14992 11542 -14975
rect 11748 -14975 12000 -14959
rect 11748 -14992 11764 -14975
rect 11526 -15009 11616 -14992
rect 11216 -15056 11616 -15009
rect 11674 -15009 11764 -14992
rect 11984 -14992 12000 -14975
rect 12206 -14975 12458 -14959
rect 12206 -14992 12222 -14975
rect 11984 -15009 12074 -14992
rect 11674 -15056 12074 -15009
rect 12132 -15009 12222 -14992
rect 12442 -14992 12458 -14975
rect 12664 -14975 12916 -14959
rect 12664 -14992 12680 -14975
rect 12442 -15009 12532 -14992
rect 12132 -15056 12532 -15009
rect 12590 -15009 12680 -14992
rect 12900 -14992 12916 -14975
rect 13122 -14975 13374 -14959
rect 13122 -14992 13138 -14975
rect 12900 -15009 12990 -14992
rect 12590 -15056 12990 -15009
rect 13048 -15009 13138 -14992
rect 13358 -14992 13374 -14975
rect 13580 -14975 13832 -14959
rect 13580 -14992 13596 -14975
rect 13358 -15009 13448 -14992
rect 13048 -15056 13448 -15009
rect 13506 -15009 13596 -14992
rect 13816 -14992 13832 -14975
rect 14038 -14975 14290 -14959
rect 14038 -14992 14054 -14975
rect 13816 -15009 13906 -14992
rect 13506 -15056 13906 -15009
rect 13964 -15009 14054 -14992
rect 14274 -14992 14290 -14975
rect 14496 -14975 14748 -14959
rect 14496 -14992 14512 -14975
rect 14274 -15009 14364 -14992
rect 13964 -15056 14364 -15009
rect 14422 -15009 14512 -14992
rect 14732 -14992 14748 -14975
rect 14954 -14975 15206 -14959
rect 14954 -14992 14970 -14975
rect 14732 -15009 14822 -14992
rect 14422 -15056 14822 -15009
rect 14880 -15009 14970 -14992
rect 15190 -14992 15206 -14975
rect 15412 -14975 15664 -14959
rect 15412 -14992 15428 -14975
rect 15190 -15009 15280 -14992
rect 14880 -15056 15280 -15009
rect 15338 -15009 15428 -14992
rect 15648 -14992 15664 -14975
rect 15870 -14975 16122 -14959
rect 15870 -14992 15886 -14975
rect 15648 -15009 15738 -14992
rect 15338 -15056 15738 -15009
rect 15796 -15009 15886 -14992
rect 16106 -14992 16122 -14975
rect 16328 -14975 16580 -14959
rect 16328 -14992 16344 -14975
rect 16106 -15009 16196 -14992
rect 15796 -15056 16196 -15009
rect 16254 -15009 16344 -14992
rect 16564 -14992 16580 -14975
rect 16786 -14975 17038 -14959
rect 16786 -14992 16802 -14975
rect 16564 -15009 16654 -14992
rect 16254 -15056 16654 -15009
rect 16712 -15009 16802 -14992
rect 17022 -14992 17038 -14975
rect 17244 -14975 17496 -14959
rect 17244 -14992 17260 -14975
rect 17022 -15009 17112 -14992
rect 16712 -15056 17112 -15009
rect 17170 -15009 17260 -14992
rect 17480 -14992 17496 -14975
rect 17480 -15009 17570 -14992
rect 17170 -15056 17570 -15009
rect 9384 -16703 9784 -16656
rect 9384 -16720 9474 -16703
rect 9458 -16737 9474 -16720
rect 9694 -16720 9784 -16703
rect 9842 -16703 10242 -16656
rect 9842 -16720 9932 -16703
rect 9694 -16737 9710 -16720
rect 9458 -16753 9710 -16737
rect 9916 -16737 9932 -16720
rect 10152 -16720 10242 -16703
rect 10300 -16703 10700 -16656
rect 10300 -16720 10390 -16703
rect 10152 -16737 10168 -16720
rect 9916 -16753 10168 -16737
rect 10374 -16737 10390 -16720
rect 10610 -16720 10700 -16703
rect 10758 -16703 11158 -16656
rect 10758 -16720 10848 -16703
rect 10610 -16737 10626 -16720
rect 10374 -16753 10626 -16737
rect 10832 -16737 10848 -16720
rect 11068 -16720 11158 -16703
rect 11216 -16703 11616 -16656
rect 11216 -16720 11306 -16703
rect 11068 -16737 11084 -16720
rect 10832 -16753 11084 -16737
rect 11290 -16737 11306 -16720
rect 11526 -16720 11616 -16703
rect 11674 -16703 12074 -16656
rect 11674 -16720 11764 -16703
rect 11526 -16737 11542 -16720
rect 11290 -16753 11542 -16737
rect 11748 -16737 11764 -16720
rect 11984 -16720 12074 -16703
rect 12132 -16703 12532 -16656
rect 12132 -16720 12222 -16703
rect 11984 -16737 12000 -16720
rect 11748 -16753 12000 -16737
rect 12206 -16737 12222 -16720
rect 12442 -16720 12532 -16703
rect 12590 -16703 12990 -16656
rect 12590 -16720 12680 -16703
rect 12442 -16737 12458 -16720
rect 12206 -16753 12458 -16737
rect 12664 -16737 12680 -16720
rect 12900 -16720 12990 -16703
rect 13048 -16703 13448 -16656
rect 13048 -16720 13138 -16703
rect 12900 -16737 12916 -16720
rect 12664 -16753 12916 -16737
rect 13122 -16737 13138 -16720
rect 13358 -16720 13448 -16703
rect 13506 -16703 13906 -16656
rect 13506 -16720 13596 -16703
rect 13358 -16737 13374 -16720
rect 13122 -16753 13374 -16737
rect 13580 -16737 13596 -16720
rect 13816 -16720 13906 -16703
rect 13964 -16703 14364 -16656
rect 13964 -16720 14054 -16703
rect 13816 -16737 13832 -16720
rect 13580 -16753 13832 -16737
rect 14038 -16737 14054 -16720
rect 14274 -16720 14364 -16703
rect 14422 -16703 14822 -16656
rect 14422 -16720 14512 -16703
rect 14274 -16737 14290 -16720
rect 14038 -16753 14290 -16737
rect 14496 -16737 14512 -16720
rect 14732 -16720 14822 -16703
rect 14880 -16703 15280 -16656
rect 14880 -16720 14970 -16703
rect 14732 -16737 14748 -16720
rect 14496 -16753 14748 -16737
rect 14954 -16737 14970 -16720
rect 15190 -16720 15280 -16703
rect 15338 -16703 15738 -16656
rect 15338 -16720 15428 -16703
rect 15190 -16737 15206 -16720
rect 14954 -16753 15206 -16737
rect 15412 -16737 15428 -16720
rect 15648 -16720 15738 -16703
rect 15796 -16703 16196 -16656
rect 15796 -16720 15886 -16703
rect 15648 -16737 15664 -16720
rect 15412 -16753 15664 -16737
rect 15870 -16737 15886 -16720
rect 16106 -16720 16196 -16703
rect 16254 -16703 16654 -16656
rect 16254 -16720 16344 -16703
rect 16106 -16737 16122 -16720
rect 15870 -16753 16122 -16737
rect 16328 -16737 16344 -16720
rect 16564 -16720 16654 -16703
rect 16712 -16703 17112 -16656
rect 16712 -16720 16802 -16703
rect 16564 -16737 16580 -16720
rect 16328 -16753 16580 -16737
rect 16786 -16737 16802 -16720
rect 17022 -16720 17112 -16703
rect 17170 -16703 17570 -16656
rect 17170 -16720 17260 -16703
rect 17022 -16737 17038 -16720
rect 16786 -16753 17038 -16737
rect 17244 -16737 17260 -16720
rect 17480 -16720 17570 -16703
rect 17480 -16737 17496 -16720
rect 17244 -16753 17496 -16737
rect 8899 -17640 9151 -17624
rect 8899 -17657 8915 -17640
rect 8825 -17674 8915 -17657
rect 9135 -17657 9151 -17640
rect 9357 -17640 9609 -17624
rect 9357 -17657 9373 -17640
rect 9135 -17674 9225 -17657
rect 8825 -17721 9225 -17674
rect 9283 -17674 9373 -17657
rect 9593 -17657 9609 -17640
rect 9815 -17640 10067 -17624
rect 9815 -17657 9831 -17640
rect 9593 -17674 9683 -17657
rect 9283 -17721 9683 -17674
rect 9741 -17674 9831 -17657
rect 10051 -17657 10067 -17640
rect 10273 -17640 10525 -17624
rect 10273 -17657 10289 -17640
rect 10051 -17674 10141 -17657
rect 9741 -17721 10141 -17674
rect 10199 -17674 10289 -17657
rect 10509 -17657 10525 -17640
rect 10731 -17640 10983 -17624
rect 10731 -17657 10747 -17640
rect 10509 -17674 10599 -17657
rect 10199 -17721 10599 -17674
rect 10657 -17674 10747 -17657
rect 10967 -17657 10983 -17640
rect 11189 -17640 11441 -17624
rect 11189 -17657 11205 -17640
rect 10967 -17674 11057 -17657
rect 10657 -17721 11057 -17674
rect 11115 -17674 11205 -17657
rect 11425 -17657 11441 -17640
rect 11647 -17640 11899 -17624
rect 11647 -17657 11663 -17640
rect 11425 -17674 11515 -17657
rect 11115 -17721 11515 -17674
rect 11573 -17674 11663 -17657
rect 11883 -17657 11899 -17640
rect 12105 -17640 12357 -17624
rect 12105 -17657 12121 -17640
rect 11883 -17674 11973 -17657
rect 11573 -17721 11973 -17674
rect 12031 -17674 12121 -17657
rect 12341 -17657 12357 -17640
rect 12563 -17640 12815 -17624
rect 12563 -17657 12579 -17640
rect 12341 -17674 12431 -17657
rect 12031 -17721 12431 -17674
rect 12489 -17674 12579 -17657
rect 12799 -17657 12815 -17640
rect 13021 -17640 13273 -17624
rect 13021 -17657 13037 -17640
rect 12799 -17674 12889 -17657
rect 12489 -17721 12889 -17674
rect 12947 -17674 13037 -17657
rect 13257 -17657 13273 -17640
rect 13899 -17640 14151 -17624
rect 13899 -17657 13915 -17640
rect 13257 -17674 13347 -17657
rect 12947 -17721 13347 -17674
rect 13825 -17674 13915 -17657
rect 14135 -17657 14151 -17640
rect 14357 -17640 14609 -17624
rect 14357 -17657 14373 -17640
rect 14135 -17674 14225 -17657
rect 13825 -17721 14225 -17674
rect 14283 -17674 14373 -17657
rect 14593 -17657 14609 -17640
rect 14815 -17640 15067 -17624
rect 14815 -17657 14831 -17640
rect 14593 -17674 14683 -17657
rect 14283 -17721 14683 -17674
rect 14741 -17674 14831 -17657
rect 15051 -17657 15067 -17640
rect 15273 -17640 15525 -17624
rect 15273 -17657 15289 -17640
rect 15051 -17674 15141 -17657
rect 14741 -17721 15141 -17674
rect 15199 -17674 15289 -17657
rect 15509 -17657 15525 -17640
rect 15731 -17640 15983 -17624
rect 15731 -17657 15747 -17640
rect 15509 -17674 15599 -17657
rect 15199 -17721 15599 -17674
rect 15657 -17674 15747 -17657
rect 15967 -17657 15983 -17640
rect 16189 -17640 16441 -17624
rect 16189 -17657 16205 -17640
rect 15967 -17674 16057 -17657
rect 15657 -17721 16057 -17674
rect 16115 -17674 16205 -17657
rect 16425 -17657 16441 -17640
rect 16647 -17640 16899 -17624
rect 16647 -17657 16663 -17640
rect 16425 -17674 16515 -17657
rect 16115 -17721 16515 -17674
rect 16573 -17674 16663 -17657
rect 16883 -17657 16899 -17640
rect 17105 -17640 17357 -17624
rect 17105 -17657 17121 -17640
rect 16883 -17674 16973 -17657
rect 16573 -17721 16973 -17674
rect 17031 -17674 17121 -17657
rect 17341 -17657 17357 -17640
rect 17563 -17640 17815 -17624
rect 17563 -17657 17579 -17640
rect 17341 -17674 17431 -17657
rect 17031 -17721 17431 -17674
rect 17489 -17674 17579 -17657
rect 17799 -17657 17815 -17640
rect 18021 -17640 18273 -17624
rect 18021 -17657 18037 -17640
rect 17799 -17674 17889 -17657
rect 17489 -17721 17889 -17674
rect 17947 -17674 18037 -17657
rect 18257 -17657 18273 -17640
rect 18257 -17674 18347 -17657
rect 17947 -17721 18347 -17674
rect 8825 -18968 9225 -18921
rect 8825 -18985 8915 -18968
rect 8899 -19002 8915 -18985
rect 9135 -18985 9225 -18968
rect 9283 -18968 9683 -18921
rect 9283 -18985 9373 -18968
rect 9135 -19002 9151 -18985
rect 8899 -19018 9151 -19002
rect 9357 -19002 9373 -18985
rect 9593 -18985 9683 -18968
rect 9741 -18968 10141 -18921
rect 9741 -18985 9831 -18968
rect 9593 -19002 9609 -18985
rect 9357 -19018 9609 -19002
rect 9815 -19002 9831 -18985
rect 10051 -18985 10141 -18968
rect 10199 -18968 10599 -18921
rect 10199 -18985 10289 -18968
rect 10051 -19002 10067 -18985
rect 9815 -19018 10067 -19002
rect 10273 -19002 10289 -18985
rect 10509 -18985 10599 -18968
rect 10657 -18968 11057 -18921
rect 10657 -18985 10747 -18968
rect 10509 -19002 10525 -18985
rect 10273 -19018 10525 -19002
rect 10731 -19002 10747 -18985
rect 10967 -18985 11057 -18968
rect 11115 -18968 11515 -18921
rect 11115 -18985 11205 -18968
rect 10967 -19002 10983 -18985
rect 10731 -19018 10983 -19002
rect 11189 -19002 11205 -18985
rect 11425 -18985 11515 -18968
rect 11573 -18968 11973 -18921
rect 11573 -18985 11663 -18968
rect 11425 -19002 11441 -18985
rect 11189 -19018 11441 -19002
rect 11647 -19002 11663 -18985
rect 11883 -18985 11973 -18968
rect 12031 -18968 12431 -18921
rect 12031 -18985 12121 -18968
rect 11883 -19002 11899 -18985
rect 11647 -19018 11899 -19002
rect 12105 -19002 12121 -18985
rect 12341 -18985 12431 -18968
rect 12489 -18968 12889 -18921
rect 12489 -18985 12579 -18968
rect 12341 -19002 12357 -18985
rect 12105 -19018 12357 -19002
rect 12563 -19002 12579 -18985
rect 12799 -18985 12889 -18968
rect 12947 -18968 13347 -18921
rect 12947 -18985 13037 -18968
rect 12799 -19002 12815 -18985
rect 12563 -19018 12815 -19002
rect 13021 -19002 13037 -18985
rect 13257 -18985 13347 -18968
rect 13825 -18968 14225 -18921
rect 13825 -18985 13915 -18968
rect 13257 -19002 13273 -18985
rect 13021 -19018 13273 -19002
rect 13899 -19002 13915 -18985
rect 14135 -18985 14225 -18968
rect 14283 -18968 14683 -18921
rect 14283 -18985 14373 -18968
rect 14135 -19002 14151 -18985
rect 13899 -19018 14151 -19002
rect 14357 -19002 14373 -18985
rect 14593 -18985 14683 -18968
rect 14741 -18968 15141 -18921
rect 14741 -18985 14831 -18968
rect 14593 -19002 14609 -18985
rect 14357 -19018 14609 -19002
rect 14815 -19002 14831 -18985
rect 15051 -18985 15141 -18968
rect 15199 -18968 15599 -18921
rect 15199 -18985 15289 -18968
rect 15051 -19002 15067 -18985
rect 14815 -19018 15067 -19002
rect 15273 -19002 15289 -18985
rect 15509 -18985 15599 -18968
rect 15657 -18968 16057 -18921
rect 15657 -18985 15747 -18968
rect 15509 -19002 15525 -18985
rect 15273 -19018 15525 -19002
rect 15731 -19002 15747 -18985
rect 15967 -18985 16057 -18968
rect 16115 -18968 16515 -18921
rect 16115 -18985 16205 -18968
rect 15967 -19002 15983 -18985
rect 15731 -19018 15983 -19002
rect 16189 -19002 16205 -18985
rect 16425 -18985 16515 -18968
rect 16573 -18968 16973 -18921
rect 16573 -18985 16663 -18968
rect 16425 -19002 16441 -18985
rect 16189 -19018 16441 -19002
rect 16647 -19002 16663 -18985
rect 16883 -18985 16973 -18968
rect 17031 -18968 17431 -18921
rect 17031 -18985 17121 -18968
rect 16883 -19002 16899 -18985
rect 16647 -19018 16899 -19002
rect 17105 -19002 17121 -18985
rect 17341 -18985 17431 -18968
rect 17489 -18968 17889 -18921
rect 17489 -18985 17579 -18968
rect 17341 -19002 17357 -18985
rect 17105 -19018 17357 -19002
rect 17563 -19002 17579 -18985
rect 17799 -18985 17889 -18968
rect 17947 -18968 18347 -18921
rect 17947 -18985 18037 -18968
rect 17799 -19002 17815 -18985
rect 17563 -19018 17815 -19002
rect 18021 -19002 18037 -18985
rect 18257 -18985 18347 -18968
rect 18257 -19002 18273 -18985
rect 18021 -19018 18273 -19002
rect 24458 -14975 24710 -14959
rect 24458 -14992 24474 -14975
rect 24384 -15009 24474 -14992
rect 24694 -14992 24710 -14975
rect 24916 -14975 25168 -14959
rect 24916 -14992 24932 -14975
rect 24694 -15009 24784 -14992
rect 24384 -15056 24784 -15009
rect 24842 -15009 24932 -14992
rect 25152 -14992 25168 -14975
rect 25374 -14975 25626 -14959
rect 25374 -14992 25390 -14975
rect 25152 -15009 25242 -14992
rect 24842 -15056 25242 -15009
rect 25300 -15009 25390 -14992
rect 25610 -14992 25626 -14975
rect 25832 -14975 26084 -14959
rect 25832 -14992 25848 -14975
rect 25610 -15009 25700 -14992
rect 25300 -15056 25700 -15009
rect 25758 -15009 25848 -14992
rect 26068 -14992 26084 -14975
rect 26290 -14975 26542 -14959
rect 26290 -14992 26306 -14975
rect 26068 -15009 26158 -14992
rect 25758 -15056 26158 -15009
rect 26216 -15009 26306 -14992
rect 26526 -14992 26542 -14975
rect 26748 -14975 27000 -14959
rect 26748 -14992 26764 -14975
rect 26526 -15009 26616 -14992
rect 26216 -15056 26616 -15009
rect 26674 -15009 26764 -14992
rect 26984 -14992 27000 -14975
rect 27206 -14975 27458 -14959
rect 27206 -14992 27222 -14975
rect 26984 -15009 27074 -14992
rect 26674 -15056 27074 -15009
rect 27132 -15009 27222 -14992
rect 27442 -14992 27458 -14975
rect 27664 -14975 27916 -14959
rect 27664 -14992 27680 -14975
rect 27442 -15009 27532 -14992
rect 27132 -15056 27532 -15009
rect 27590 -15009 27680 -14992
rect 27900 -14992 27916 -14975
rect 28122 -14975 28374 -14959
rect 28122 -14992 28138 -14975
rect 27900 -15009 27990 -14992
rect 27590 -15056 27990 -15009
rect 28048 -15009 28138 -14992
rect 28358 -14992 28374 -14975
rect 28580 -14975 28832 -14959
rect 28580 -14992 28596 -14975
rect 28358 -15009 28448 -14992
rect 28048 -15056 28448 -15009
rect 28506 -15009 28596 -14992
rect 28816 -14992 28832 -14975
rect 29038 -14975 29290 -14959
rect 29038 -14992 29054 -14975
rect 28816 -15009 28906 -14992
rect 28506 -15056 28906 -15009
rect 28964 -15009 29054 -14992
rect 29274 -14992 29290 -14975
rect 29496 -14975 29748 -14959
rect 29496 -14992 29512 -14975
rect 29274 -15009 29364 -14992
rect 28964 -15056 29364 -15009
rect 29422 -15009 29512 -14992
rect 29732 -14992 29748 -14975
rect 29954 -14975 30206 -14959
rect 29954 -14992 29970 -14975
rect 29732 -15009 29822 -14992
rect 29422 -15056 29822 -15009
rect 29880 -15009 29970 -14992
rect 30190 -14992 30206 -14975
rect 30412 -14975 30664 -14959
rect 30412 -14992 30428 -14975
rect 30190 -15009 30280 -14992
rect 29880 -15056 30280 -15009
rect 30338 -15009 30428 -14992
rect 30648 -14992 30664 -14975
rect 30870 -14975 31122 -14959
rect 30870 -14992 30886 -14975
rect 30648 -15009 30738 -14992
rect 30338 -15056 30738 -15009
rect 30796 -15009 30886 -14992
rect 31106 -14992 31122 -14975
rect 31328 -14975 31580 -14959
rect 31328 -14992 31344 -14975
rect 31106 -15009 31196 -14992
rect 30796 -15056 31196 -15009
rect 31254 -15009 31344 -14992
rect 31564 -14992 31580 -14975
rect 31786 -14975 32038 -14959
rect 31786 -14992 31802 -14975
rect 31564 -15009 31654 -14992
rect 31254 -15056 31654 -15009
rect 31712 -15009 31802 -14992
rect 32022 -14992 32038 -14975
rect 32244 -14975 32496 -14959
rect 32244 -14992 32260 -14975
rect 32022 -15009 32112 -14992
rect 31712 -15056 32112 -15009
rect 32170 -15009 32260 -14992
rect 32480 -14992 32496 -14975
rect 32480 -15009 32570 -14992
rect 32170 -15056 32570 -15009
rect 24384 -16703 24784 -16656
rect 24384 -16720 24474 -16703
rect 24458 -16737 24474 -16720
rect 24694 -16720 24784 -16703
rect 24842 -16703 25242 -16656
rect 24842 -16720 24932 -16703
rect 24694 -16737 24710 -16720
rect 24458 -16753 24710 -16737
rect 24916 -16737 24932 -16720
rect 25152 -16720 25242 -16703
rect 25300 -16703 25700 -16656
rect 25300 -16720 25390 -16703
rect 25152 -16737 25168 -16720
rect 24916 -16753 25168 -16737
rect 25374 -16737 25390 -16720
rect 25610 -16720 25700 -16703
rect 25758 -16703 26158 -16656
rect 25758 -16720 25848 -16703
rect 25610 -16737 25626 -16720
rect 25374 -16753 25626 -16737
rect 25832 -16737 25848 -16720
rect 26068 -16720 26158 -16703
rect 26216 -16703 26616 -16656
rect 26216 -16720 26306 -16703
rect 26068 -16737 26084 -16720
rect 25832 -16753 26084 -16737
rect 26290 -16737 26306 -16720
rect 26526 -16720 26616 -16703
rect 26674 -16703 27074 -16656
rect 26674 -16720 26764 -16703
rect 26526 -16737 26542 -16720
rect 26290 -16753 26542 -16737
rect 26748 -16737 26764 -16720
rect 26984 -16720 27074 -16703
rect 27132 -16703 27532 -16656
rect 27132 -16720 27222 -16703
rect 26984 -16737 27000 -16720
rect 26748 -16753 27000 -16737
rect 27206 -16737 27222 -16720
rect 27442 -16720 27532 -16703
rect 27590 -16703 27990 -16656
rect 27590 -16720 27680 -16703
rect 27442 -16737 27458 -16720
rect 27206 -16753 27458 -16737
rect 27664 -16737 27680 -16720
rect 27900 -16720 27990 -16703
rect 28048 -16703 28448 -16656
rect 28048 -16720 28138 -16703
rect 27900 -16737 27916 -16720
rect 27664 -16753 27916 -16737
rect 28122 -16737 28138 -16720
rect 28358 -16720 28448 -16703
rect 28506 -16703 28906 -16656
rect 28506 -16720 28596 -16703
rect 28358 -16737 28374 -16720
rect 28122 -16753 28374 -16737
rect 28580 -16737 28596 -16720
rect 28816 -16720 28906 -16703
rect 28964 -16703 29364 -16656
rect 28964 -16720 29054 -16703
rect 28816 -16737 28832 -16720
rect 28580 -16753 28832 -16737
rect 29038 -16737 29054 -16720
rect 29274 -16720 29364 -16703
rect 29422 -16703 29822 -16656
rect 29422 -16720 29512 -16703
rect 29274 -16737 29290 -16720
rect 29038 -16753 29290 -16737
rect 29496 -16737 29512 -16720
rect 29732 -16720 29822 -16703
rect 29880 -16703 30280 -16656
rect 29880 -16720 29970 -16703
rect 29732 -16737 29748 -16720
rect 29496 -16753 29748 -16737
rect 29954 -16737 29970 -16720
rect 30190 -16720 30280 -16703
rect 30338 -16703 30738 -16656
rect 30338 -16720 30428 -16703
rect 30190 -16737 30206 -16720
rect 29954 -16753 30206 -16737
rect 30412 -16737 30428 -16720
rect 30648 -16720 30738 -16703
rect 30796 -16703 31196 -16656
rect 30796 -16720 30886 -16703
rect 30648 -16737 30664 -16720
rect 30412 -16753 30664 -16737
rect 30870 -16737 30886 -16720
rect 31106 -16720 31196 -16703
rect 31254 -16703 31654 -16656
rect 31254 -16720 31344 -16703
rect 31106 -16737 31122 -16720
rect 30870 -16753 31122 -16737
rect 31328 -16737 31344 -16720
rect 31564 -16720 31654 -16703
rect 31712 -16703 32112 -16656
rect 31712 -16720 31802 -16703
rect 31564 -16737 31580 -16720
rect 31328 -16753 31580 -16737
rect 31786 -16737 31802 -16720
rect 32022 -16720 32112 -16703
rect 32170 -16703 32570 -16656
rect 32170 -16720 32260 -16703
rect 32022 -16737 32038 -16720
rect 31786 -16753 32038 -16737
rect 32244 -16737 32260 -16720
rect 32480 -16720 32570 -16703
rect 32480 -16737 32496 -16720
rect 32244 -16753 32496 -16737
rect 23899 -17640 24151 -17624
rect 23899 -17657 23915 -17640
rect 23825 -17674 23915 -17657
rect 24135 -17657 24151 -17640
rect 24357 -17640 24609 -17624
rect 24357 -17657 24373 -17640
rect 24135 -17674 24225 -17657
rect 23825 -17721 24225 -17674
rect 24283 -17674 24373 -17657
rect 24593 -17657 24609 -17640
rect 24815 -17640 25067 -17624
rect 24815 -17657 24831 -17640
rect 24593 -17674 24683 -17657
rect 24283 -17721 24683 -17674
rect 24741 -17674 24831 -17657
rect 25051 -17657 25067 -17640
rect 25273 -17640 25525 -17624
rect 25273 -17657 25289 -17640
rect 25051 -17674 25141 -17657
rect 24741 -17721 25141 -17674
rect 25199 -17674 25289 -17657
rect 25509 -17657 25525 -17640
rect 25731 -17640 25983 -17624
rect 25731 -17657 25747 -17640
rect 25509 -17674 25599 -17657
rect 25199 -17721 25599 -17674
rect 25657 -17674 25747 -17657
rect 25967 -17657 25983 -17640
rect 26189 -17640 26441 -17624
rect 26189 -17657 26205 -17640
rect 25967 -17674 26057 -17657
rect 25657 -17721 26057 -17674
rect 26115 -17674 26205 -17657
rect 26425 -17657 26441 -17640
rect 26647 -17640 26899 -17624
rect 26647 -17657 26663 -17640
rect 26425 -17674 26515 -17657
rect 26115 -17721 26515 -17674
rect 26573 -17674 26663 -17657
rect 26883 -17657 26899 -17640
rect 27105 -17640 27357 -17624
rect 27105 -17657 27121 -17640
rect 26883 -17674 26973 -17657
rect 26573 -17721 26973 -17674
rect 27031 -17674 27121 -17657
rect 27341 -17657 27357 -17640
rect 27563 -17640 27815 -17624
rect 27563 -17657 27579 -17640
rect 27341 -17674 27431 -17657
rect 27031 -17721 27431 -17674
rect 27489 -17674 27579 -17657
rect 27799 -17657 27815 -17640
rect 28021 -17640 28273 -17624
rect 28021 -17657 28037 -17640
rect 27799 -17674 27889 -17657
rect 27489 -17721 27889 -17674
rect 27947 -17674 28037 -17657
rect 28257 -17657 28273 -17640
rect 28899 -17640 29151 -17624
rect 28899 -17657 28915 -17640
rect 28257 -17674 28347 -17657
rect 27947 -17721 28347 -17674
rect 28825 -17674 28915 -17657
rect 29135 -17657 29151 -17640
rect 29357 -17640 29609 -17624
rect 29357 -17657 29373 -17640
rect 29135 -17674 29225 -17657
rect 28825 -17721 29225 -17674
rect 29283 -17674 29373 -17657
rect 29593 -17657 29609 -17640
rect 29815 -17640 30067 -17624
rect 29815 -17657 29831 -17640
rect 29593 -17674 29683 -17657
rect 29283 -17721 29683 -17674
rect 29741 -17674 29831 -17657
rect 30051 -17657 30067 -17640
rect 30273 -17640 30525 -17624
rect 30273 -17657 30289 -17640
rect 30051 -17674 30141 -17657
rect 29741 -17721 30141 -17674
rect 30199 -17674 30289 -17657
rect 30509 -17657 30525 -17640
rect 30731 -17640 30983 -17624
rect 30731 -17657 30747 -17640
rect 30509 -17674 30599 -17657
rect 30199 -17721 30599 -17674
rect 30657 -17674 30747 -17657
rect 30967 -17657 30983 -17640
rect 31189 -17640 31441 -17624
rect 31189 -17657 31205 -17640
rect 30967 -17674 31057 -17657
rect 30657 -17721 31057 -17674
rect 31115 -17674 31205 -17657
rect 31425 -17657 31441 -17640
rect 31647 -17640 31899 -17624
rect 31647 -17657 31663 -17640
rect 31425 -17674 31515 -17657
rect 31115 -17721 31515 -17674
rect 31573 -17674 31663 -17657
rect 31883 -17657 31899 -17640
rect 32105 -17640 32357 -17624
rect 32105 -17657 32121 -17640
rect 31883 -17674 31973 -17657
rect 31573 -17721 31973 -17674
rect 32031 -17674 32121 -17657
rect 32341 -17657 32357 -17640
rect 32563 -17640 32815 -17624
rect 32563 -17657 32579 -17640
rect 32341 -17674 32431 -17657
rect 32031 -17721 32431 -17674
rect 32489 -17674 32579 -17657
rect 32799 -17657 32815 -17640
rect 33021 -17640 33273 -17624
rect 33021 -17657 33037 -17640
rect 32799 -17674 32889 -17657
rect 32489 -17721 32889 -17674
rect 32947 -17674 33037 -17657
rect 33257 -17657 33273 -17640
rect 33257 -17674 33347 -17657
rect 32947 -17721 33347 -17674
rect 23825 -18968 24225 -18921
rect 23825 -18985 23915 -18968
rect 23899 -19002 23915 -18985
rect 24135 -18985 24225 -18968
rect 24283 -18968 24683 -18921
rect 24283 -18985 24373 -18968
rect 24135 -19002 24151 -18985
rect 23899 -19018 24151 -19002
rect 24357 -19002 24373 -18985
rect 24593 -18985 24683 -18968
rect 24741 -18968 25141 -18921
rect 24741 -18985 24831 -18968
rect 24593 -19002 24609 -18985
rect 24357 -19018 24609 -19002
rect 24815 -19002 24831 -18985
rect 25051 -18985 25141 -18968
rect 25199 -18968 25599 -18921
rect 25199 -18985 25289 -18968
rect 25051 -19002 25067 -18985
rect 24815 -19018 25067 -19002
rect 25273 -19002 25289 -18985
rect 25509 -18985 25599 -18968
rect 25657 -18968 26057 -18921
rect 25657 -18985 25747 -18968
rect 25509 -19002 25525 -18985
rect 25273 -19018 25525 -19002
rect 25731 -19002 25747 -18985
rect 25967 -18985 26057 -18968
rect 26115 -18968 26515 -18921
rect 26115 -18985 26205 -18968
rect 25967 -19002 25983 -18985
rect 25731 -19018 25983 -19002
rect 26189 -19002 26205 -18985
rect 26425 -18985 26515 -18968
rect 26573 -18968 26973 -18921
rect 26573 -18985 26663 -18968
rect 26425 -19002 26441 -18985
rect 26189 -19018 26441 -19002
rect 26647 -19002 26663 -18985
rect 26883 -18985 26973 -18968
rect 27031 -18968 27431 -18921
rect 27031 -18985 27121 -18968
rect 26883 -19002 26899 -18985
rect 26647 -19018 26899 -19002
rect 27105 -19002 27121 -18985
rect 27341 -18985 27431 -18968
rect 27489 -18968 27889 -18921
rect 27489 -18985 27579 -18968
rect 27341 -19002 27357 -18985
rect 27105 -19018 27357 -19002
rect 27563 -19002 27579 -18985
rect 27799 -18985 27889 -18968
rect 27947 -18968 28347 -18921
rect 27947 -18985 28037 -18968
rect 27799 -19002 27815 -18985
rect 27563 -19018 27815 -19002
rect 28021 -19002 28037 -18985
rect 28257 -18985 28347 -18968
rect 28825 -18968 29225 -18921
rect 28825 -18985 28915 -18968
rect 28257 -19002 28273 -18985
rect 28021 -19018 28273 -19002
rect 28899 -19002 28915 -18985
rect 29135 -18985 29225 -18968
rect 29283 -18968 29683 -18921
rect 29283 -18985 29373 -18968
rect 29135 -19002 29151 -18985
rect 28899 -19018 29151 -19002
rect 29357 -19002 29373 -18985
rect 29593 -18985 29683 -18968
rect 29741 -18968 30141 -18921
rect 29741 -18985 29831 -18968
rect 29593 -19002 29609 -18985
rect 29357 -19018 29609 -19002
rect 29815 -19002 29831 -18985
rect 30051 -18985 30141 -18968
rect 30199 -18968 30599 -18921
rect 30199 -18985 30289 -18968
rect 30051 -19002 30067 -18985
rect 29815 -19018 30067 -19002
rect 30273 -19002 30289 -18985
rect 30509 -18985 30599 -18968
rect 30657 -18968 31057 -18921
rect 30657 -18985 30747 -18968
rect 30509 -19002 30525 -18985
rect 30273 -19018 30525 -19002
rect 30731 -19002 30747 -18985
rect 30967 -18985 31057 -18968
rect 31115 -18968 31515 -18921
rect 31115 -18985 31205 -18968
rect 30967 -19002 30983 -18985
rect 30731 -19018 30983 -19002
rect 31189 -19002 31205 -18985
rect 31425 -18985 31515 -18968
rect 31573 -18968 31973 -18921
rect 31573 -18985 31663 -18968
rect 31425 -19002 31441 -18985
rect 31189 -19018 31441 -19002
rect 31647 -19002 31663 -18985
rect 31883 -18985 31973 -18968
rect 32031 -18968 32431 -18921
rect 32031 -18985 32121 -18968
rect 31883 -19002 31899 -18985
rect 31647 -19018 31899 -19002
rect 32105 -19002 32121 -18985
rect 32341 -18985 32431 -18968
rect 32489 -18968 32889 -18921
rect 32489 -18985 32579 -18968
rect 32341 -19002 32357 -18985
rect 32105 -19018 32357 -19002
rect 32563 -19002 32579 -18985
rect 32799 -18985 32889 -18968
rect 32947 -18968 33347 -18921
rect 32947 -18985 33037 -18968
rect 32799 -19002 32815 -18985
rect 32563 -19018 32815 -19002
rect 33021 -19002 33037 -18985
rect 33257 -18985 33347 -18968
rect 33257 -19002 33273 -18985
rect 33021 -19018 33273 -19002
rect 8898 -20142 9150 -20126
rect 8898 -20159 8914 -20142
rect 8824 -20176 8914 -20159
rect 9134 -20159 9150 -20142
rect 9356 -20142 9608 -20126
rect 9356 -20159 9372 -20142
rect 9134 -20176 9224 -20159
rect 8824 -20214 9224 -20176
rect 9282 -20176 9372 -20159
rect 9592 -20159 9608 -20142
rect 9814 -20142 10066 -20126
rect 9814 -20159 9830 -20142
rect 9592 -20176 9682 -20159
rect 9282 -20214 9682 -20176
rect 9740 -20176 9830 -20159
rect 10050 -20159 10066 -20142
rect 10272 -20142 10524 -20126
rect 10272 -20159 10288 -20142
rect 10050 -20176 10140 -20159
rect 9740 -20214 10140 -20176
rect 10198 -20176 10288 -20159
rect 10508 -20159 10524 -20142
rect 10730 -20142 10982 -20126
rect 10730 -20159 10746 -20142
rect 10508 -20176 10598 -20159
rect 10198 -20214 10598 -20176
rect 10656 -20176 10746 -20159
rect 10966 -20159 10982 -20142
rect 11188 -20142 11440 -20126
rect 11188 -20159 11204 -20142
rect 10966 -20176 11056 -20159
rect 10656 -20214 11056 -20176
rect 11114 -20176 11204 -20159
rect 11424 -20159 11440 -20142
rect 11646 -20142 11898 -20126
rect 11646 -20159 11662 -20142
rect 11424 -20176 11514 -20159
rect 11114 -20214 11514 -20176
rect 11572 -20176 11662 -20159
rect 11882 -20159 11898 -20142
rect 12104 -20142 12356 -20126
rect 12104 -20159 12120 -20142
rect 11882 -20176 11972 -20159
rect 11572 -20214 11972 -20176
rect 12030 -20176 12120 -20159
rect 12340 -20159 12356 -20142
rect 12562 -20142 12814 -20126
rect 12562 -20159 12578 -20142
rect 12340 -20176 12430 -20159
rect 12030 -20214 12430 -20176
rect 12488 -20176 12578 -20159
rect 12798 -20159 12814 -20142
rect 13020 -20142 13272 -20126
rect 13020 -20159 13036 -20142
rect 12798 -20176 12888 -20159
rect 12488 -20214 12888 -20176
rect 12946 -20176 13036 -20159
rect 13256 -20159 13272 -20142
rect 13898 -20142 14150 -20126
rect 13898 -20159 13914 -20142
rect 13256 -20176 13346 -20159
rect 12946 -20214 13346 -20176
rect 13824 -20176 13914 -20159
rect 14134 -20159 14150 -20142
rect 14356 -20142 14608 -20126
rect 14356 -20159 14372 -20142
rect 14134 -20176 14224 -20159
rect 13824 -20214 14224 -20176
rect 14282 -20176 14372 -20159
rect 14592 -20159 14608 -20142
rect 14814 -20142 15066 -20126
rect 14814 -20159 14830 -20142
rect 14592 -20176 14682 -20159
rect 14282 -20214 14682 -20176
rect 14740 -20176 14830 -20159
rect 15050 -20159 15066 -20142
rect 15272 -20142 15524 -20126
rect 15272 -20159 15288 -20142
rect 15050 -20176 15140 -20159
rect 14740 -20214 15140 -20176
rect 15198 -20176 15288 -20159
rect 15508 -20159 15524 -20142
rect 15730 -20142 15982 -20126
rect 15730 -20159 15746 -20142
rect 15508 -20176 15598 -20159
rect 15198 -20214 15598 -20176
rect 15656 -20176 15746 -20159
rect 15966 -20159 15982 -20142
rect 16188 -20142 16440 -20126
rect 16188 -20159 16204 -20142
rect 15966 -20176 16056 -20159
rect 15656 -20214 16056 -20176
rect 16114 -20176 16204 -20159
rect 16424 -20159 16440 -20142
rect 16646 -20142 16898 -20126
rect 16646 -20159 16662 -20142
rect 16424 -20176 16514 -20159
rect 16114 -20214 16514 -20176
rect 16572 -20176 16662 -20159
rect 16882 -20159 16898 -20142
rect 17104 -20142 17356 -20126
rect 17104 -20159 17120 -20142
rect 16882 -20176 16972 -20159
rect 16572 -20214 16972 -20176
rect 17030 -20176 17120 -20159
rect 17340 -20159 17356 -20142
rect 17562 -20142 17814 -20126
rect 17562 -20159 17578 -20142
rect 17340 -20176 17430 -20159
rect 17030 -20214 17430 -20176
rect 17488 -20176 17578 -20159
rect 17798 -20159 17814 -20142
rect 18020 -20142 18272 -20126
rect 18020 -20159 18036 -20142
rect 17798 -20176 17888 -20159
rect 17488 -20214 17888 -20176
rect 17946 -20176 18036 -20159
rect 18256 -20159 18272 -20142
rect 18256 -20176 18346 -20159
rect 17946 -20214 18346 -20176
rect 8824 -20452 9224 -20414
rect 8824 -20469 8914 -20452
rect 8898 -20486 8914 -20469
rect 9134 -20469 9224 -20452
rect 9282 -20452 9682 -20414
rect 9282 -20469 9372 -20452
rect 9134 -20486 9150 -20469
rect 8898 -20502 9150 -20486
rect 9356 -20486 9372 -20469
rect 9592 -20469 9682 -20452
rect 9740 -20452 10140 -20414
rect 9740 -20469 9830 -20452
rect 9592 -20486 9608 -20469
rect 9356 -20502 9608 -20486
rect 9814 -20486 9830 -20469
rect 10050 -20469 10140 -20452
rect 10198 -20452 10598 -20414
rect 10198 -20469 10288 -20452
rect 10050 -20486 10066 -20469
rect 9814 -20502 10066 -20486
rect 10272 -20486 10288 -20469
rect 10508 -20469 10598 -20452
rect 10656 -20452 11056 -20414
rect 10656 -20469 10746 -20452
rect 10508 -20486 10524 -20469
rect 10272 -20502 10524 -20486
rect 10730 -20486 10746 -20469
rect 10966 -20469 11056 -20452
rect 11114 -20452 11514 -20414
rect 11114 -20469 11204 -20452
rect 10966 -20486 10982 -20469
rect 10730 -20502 10982 -20486
rect 11188 -20486 11204 -20469
rect 11424 -20469 11514 -20452
rect 11572 -20452 11972 -20414
rect 11572 -20469 11662 -20452
rect 11424 -20486 11440 -20469
rect 11188 -20502 11440 -20486
rect 11646 -20486 11662 -20469
rect 11882 -20469 11972 -20452
rect 12030 -20452 12430 -20414
rect 12030 -20469 12120 -20452
rect 11882 -20486 11898 -20469
rect 11646 -20502 11898 -20486
rect 12104 -20486 12120 -20469
rect 12340 -20469 12430 -20452
rect 12488 -20452 12888 -20414
rect 12488 -20469 12578 -20452
rect 12340 -20486 12356 -20469
rect 12104 -20502 12356 -20486
rect 12562 -20486 12578 -20469
rect 12798 -20469 12888 -20452
rect 12946 -20452 13346 -20414
rect 12946 -20469 13036 -20452
rect 12798 -20486 12814 -20469
rect 12562 -20502 12814 -20486
rect 13020 -20486 13036 -20469
rect 13256 -20469 13346 -20452
rect 13824 -20452 14224 -20414
rect 13824 -20469 13914 -20452
rect 13256 -20486 13272 -20469
rect 13020 -20502 13272 -20486
rect 13898 -20486 13914 -20469
rect 14134 -20469 14224 -20452
rect 14282 -20452 14682 -20414
rect 14282 -20469 14372 -20452
rect 14134 -20486 14150 -20469
rect 13898 -20502 14150 -20486
rect 14356 -20486 14372 -20469
rect 14592 -20469 14682 -20452
rect 14740 -20452 15140 -20414
rect 14740 -20469 14830 -20452
rect 14592 -20486 14608 -20469
rect 14356 -20502 14608 -20486
rect 14814 -20486 14830 -20469
rect 15050 -20469 15140 -20452
rect 15198 -20452 15598 -20414
rect 15198 -20469 15288 -20452
rect 15050 -20486 15066 -20469
rect 14814 -20502 15066 -20486
rect 15272 -20486 15288 -20469
rect 15508 -20469 15598 -20452
rect 15656 -20452 16056 -20414
rect 15656 -20469 15746 -20452
rect 15508 -20486 15524 -20469
rect 15272 -20502 15524 -20486
rect 15730 -20486 15746 -20469
rect 15966 -20469 16056 -20452
rect 16114 -20452 16514 -20414
rect 16114 -20469 16204 -20452
rect 15966 -20486 15982 -20469
rect 15730 -20502 15982 -20486
rect 16188 -20486 16204 -20469
rect 16424 -20469 16514 -20452
rect 16572 -20452 16972 -20414
rect 16572 -20469 16662 -20452
rect 16424 -20486 16440 -20469
rect 16188 -20502 16440 -20486
rect 16646 -20486 16662 -20469
rect 16882 -20469 16972 -20452
rect 17030 -20452 17430 -20414
rect 17030 -20469 17120 -20452
rect 16882 -20486 16898 -20469
rect 16646 -20502 16898 -20486
rect 17104 -20486 17120 -20469
rect 17340 -20469 17430 -20452
rect 17488 -20452 17888 -20414
rect 17488 -20469 17578 -20452
rect 17340 -20486 17356 -20469
rect 17104 -20502 17356 -20486
rect 17562 -20486 17578 -20469
rect 17798 -20469 17888 -20452
rect 17946 -20452 18346 -20414
rect 17946 -20469 18036 -20452
rect 17798 -20486 17814 -20469
rect 17562 -20502 17814 -20486
rect 18020 -20486 18036 -20469
rect 18256 -20469 18346 -20452
rect 18256 -20486 18272 -20469
rect 18020 -20502 18272 -20486
rect 8898 -20810 9150 -20794
rect 8898 -20827 8914 -20810
rect 8824 -20844 8914 -20827
rect 9134 -20827 9150 -20810
rect 9356 -20810 9608 -20794
rect 9356 -20827 9372 -20810
rect 9134 -20844 9224 -20827
rect 8824 -20882 9224 -20844
rect 9282 -20844 9372 -20827
rect 9592 -20827 9608 -20810
rect 9814 -20810 10066 -20794
rect 9814 -20827 9830 -20810
rect 9592 -20844 9682 -20827
rect 9282 -20882 9682 -20844
rect 9740 -20844 9830 -20827
rect 10050 -20827 10066 -20810
rect 10272 -20810 10524 -20794
rect 10272 -20827 10288 -20810
rect 10050 -20844 10140 -20827
rect 9740 -20882 10140 -20844
rect 10198 -20844 10288 -20827
rect 10508 -20827 10524 -20810
rect 10730 -20810 10982 -20794
rect 10730 -20827 10746 -20810
rect 10508 -20844 10598 -20827
rect 10198 -20882 10598 -20844
rect 10656 -20844 10746 -20827
rect 10966 -20827 10982 -20810
rect 11188 -20810 11440 -20794
rect 11188 -20827 11204 -20810
rect 10966 -20844 11056 -20827
rect 10656 -20882 11056 -20844
rect 11114 -20844 11204 -20827
rect 11424 -20827 11440 -20810
rect 11646 -20810 11898 -20794
rect 11646 -20827 11662 -20810
rect 11424 -20844 11514 -20827
rect 11114 -20882 11514 -20844
rect 11572 -20844 11662 -20827
rect 11882 -20827 11898 -20810
rect 12104 -20810 12356 -20794
rect 12104 -20827 12120 -20810
rect 11882 -20844 11972 -20827
rect 11572 -20882 11972 -20844
rect 12030 -20844 12120 -20827
rect 12340 -20827 12356 -20810
rect 12562 -20810 12814 -20794
rect 12562 -20827 12578 -20810
rect 12340 -20844 12430 -20827
rect 12030 -20882 12430 -20844
rect 12488 -20844 12578 -20827
rect 12798 -20827 12814 -20810
rect 13020 -20810 13272 -20794
rect 13020 -20827 13036 -20810
rect 12798 -20844 12888 -20827
rect 12488 -20882 12888 -20844
rect 12946 -20844 13036 -20827
rect 13256 -20827 13272 -20810
rect 13256 -20844 13346 -20827
rect 12946 -20882 13346 -20844
rect 8824 -21120 9224 -21082
rect 8824 -21137 8914 -21120
rect 8898 -21154 8914 -21137
rect 9134 -21137 9224 -21120
rect 9282 -21120 9682 -21082
rect 9282 -21137 9372 -21120
rect 9134 -21154 9150 -21137
rect 8898 -21170 9150 -21154
rect 9356 -21154 9372 -21137
rect 9592 -21137 9682 -21120
rect 9740 -21120 10140 -21082
rect 9740 -21137 9830 -21120
rect 9592 -21154 9608 -21137
rect 9356 -21170 9608 -21154
rect 9814 -21154 9830 -21137
rect 10050 -21137 10140 -21120
rect 10198 -21120 10598 -21082
rect 10198 -21137 10288 -21120
rect 10050 -21154 10066 -21137
rect 9814 -21170 10066 -21154
rect 10272 -21154 10288 -21137
rect 10508 -21137 10598 -21120
rect 10656 -21120 11056 -21082
rect 10656 -21137 10746 -21120
rect 10508 -21154 10524 -21137
rect 10272 -21170 10524 -21154
rect 10730 -21154 10746 -21137
rect 10966 -21137 11056 -21120
rect 11114 -21120 11514 -21082
rect 11114 -21137 11204 -21120
rect 10966 -21154 10982 -21137
rect 10730 -21170 10982 -21154
rect 11188 -21154 11204 -21137
rect 11424 -21137 11514 -21120
rect 11572 -21120 11972 -21082
rect 11572 -21137 11662 -21120
rect 11424 -21154 11440 -21137
rect 11188 -21170 11440 -21154
rect 11646 -21154 11662 -21137
rect 11882 -21137 11972 -21120
rect 12030 -21120 12430 -21082
rect 12030 -21137 12120 -21120
rect 11882 -21154 11898 -21137
rect 11646 -21170 11898 -21154
rect 12104 -21154 12120 -21137
rect 12340 -21137 12430 -21120
rect 12488 -21120 12888 -21082
rect 12488 -21137 12578 -21120
rect 12340 -21154 12356 -21137
rect 12104 -21170 12356 -21154
rect 12562 -21154 12578 -21137
rect 12798 -21137 12888 -21120
rect 12946 -21120 13346 -21082
rect 12946 -21137 13036 -21120
rect 12798 -21154 12814 -21137
rect 12562 -21170 12814 -21154
rect 13020 -21154 13036 -21137
rect 13256 -21137 13346 -21120
rect 13256 -21154 13272 -21137
rect 13020 -21170 13272 -21154
rect 23898 -20142 24150 -20126
rect 23898 -20159 23914 -20142
rect 23824 -20176 23914 -20159
rect 24134 -20159 24150 -20142
rect 24356 -20142 24608 -20126
rect 24356 -20159 24372 -20142
rect 24134 -20176 24224 -20159
rect 23824 -20214 24224 -20176
rect 24282 -20176 24372 -20159
rect 24592 -20159 24608 -20142
rect 24814 -20142 25066 -20126
rect 24814 -20159 24830 -20142
rect 24592 -20176 24682 -20159
rect 24282 -20214 24682 -20176
rect 24740 -20176 24830 -20159
rect 25050 -20159 25066 -20142
rect 25272 -20142 25524 -20126
rect 25272 -20159 25288 -20142
rect 25050 -20176 25140 -20159
rect 24740 -20214 25140 -20176
rect 25198 -20176 25288 -20159
rect 25508 -20159 25524 -20142
rect 25730 -20142 25982 -20126
rect 25730 -20159 25746 -20142
rect 25508 -20176 25598 -20159
rect 25198 -20214 25598 -20176
rect 25656 -20176 25746 -20159
rect 25966 -20159 25982 -20142
rect 26188 -20142 26440 -20126
rect 26188 -20159 26204 -20142
rect 25966 -20176 26056 -20159
rect 25656 -20214 26056 -20176
rect 26114 -20176 26204 -20159
rect 26424 -20159 26440 -20142
rect 26646 -20142 26898 -20126
rect 26646 -20159 26662 -20142
rect 26424 -20176 26514 -20159
rect 26114 -20214 26514 -20176
rect 26572 -20176 26662 -20159
rect 26882 -20159 26898 -20142
rect 27104 -20142 27356 -20126
rect 27104 -20159 27120 -20142
rect 26882 -20176 26972 -20159
rect 26572 -20214 26972 -20176
rect 27030 -20176 27120 -20159
rect 27340 -20159 27356 -20142
rect 27562 -20142 27814 -20126
rect 27562 -20159 27578 -20142
rect 27340 -20176 27430 -20159
rect 27030 -20214 27430 -20176
rect 27488 -20176 27578 -20159
rect 27798 -20159 27814 -20142
rect 28020 -20142 28272 -20126
rect 28020 -20159 28036 -20142
rect 27798 -20176 27888 -20159
rect 27488 -20214 27888 -20176
rect 27946 -20176 28036 -20159
rect 28256 -20159 28272 -20142
rect 28898 -20142 29150 -20126
rect 28898 -20159 28914 -20142
rect 28256 -20176 28346 -20159
rect 27946 -20214 28346 -20176
rect 28824 -20176 28914 -20159
rect 29134 -20159 29150 -20142
rect 29356 -20142 29608 -20126
rect 29356 -20159 29372 -20142
rect 29134 -20176 29224 -20159
rect 28824 -20214 29224 -20176
rect 29282 -20176 29372 -20159
rect 29592 -20159 29608 -20142
rect 29814 -20142 30066 -20126
rect 29814 -20159 29830 -20142
rect 29592 -20176 29682 -20159
rect 29282 -20214 29682 -20176
rect 29740 -20176 29830 -20159
rect 30050 -20159 30066 -20142
rect 30272 -20142 30524 -20126
rect 30272 -20159 30288 -20142
rect 30050 -20176 30140 -20159
rect 29740 -20214 30140 -20176
rect 30198 -20176 30288 -20159
rect 30508 -20159 30524 -20142
rect 30730 -20142 30982 -20126
rect 30730 -20159 30746 -20142
rect 30508 -20176 30598 -20159
rect 30198 -20214 30598 -20176
rect 30656 -20176 30746 -20159
rect 30966 -20159 30982 -20142
rect 31188 -20142 31440 -20126
rect 31188 -20159 31204 -20142
rect 30966 -20176 31056 -20159
rect 30656 -20214 31056 -20176
rect 31114 -20176 31204 -20159
rect 31424 -20159 31440 -20142
rect 31646 -20142 31898 -20126
rect 31646 -20159 31662 -20142
rect 31424 -20176 31514 -20159
rect 31114 -20214 31514 -20176
rect 31572 -20176 31662 -20159
rect 31882 -20159 31898 -20142
rect 32104 -20142 32356 -20126
rect 32104 -20159 32120 -20142
rect 31882 -20176 31972 -20159
rect 31572 -20214 31972 -20176
rect 32030 -20176 32120 -20159
rect 32340 -20159 32356 -20142
rect 32562 -20142 32814 -20126
rect 32562 -20159 32578 -20142
rect 32340 -20176 32430 -20159
rect 32030 -20214 32430 -20176
rect 32488 -20176 32578 -20159
rect 32798 -20159 32814 -20142
rect 33020 -20142 33272 -20126
rect 33020 -20159 33036 -20142
rect 32798 -20176 32888 -20159
rect 32488 -20214 32888 -20176
rect 32946 -20176 33036 -20159
rect 33256 -20159 33272 -20142
rect 33256 -20176 33346 -20159
rect 32946 -20214 33346 -20176
rect 23824 -20452 24224 -20414
rect 23824 -20469 23914 -20452
rect 23898 -20486 23914 -20469
rect 24134 -20469 24224 -20452
rect 24282 -20452 24682 -20414
rect 24282 -20469 24372 -20452
rect 24134 -20486 24150 -20469
rect 23898 -20502 24150 -20486
rect 24356 -20486 24372 -20469
rect 24592 -20469 24682 -20452
rect 24740 -20452 25140 -20414
rect 24740 -20469 24830 -20452
rect 24592 -20486 24608 -20469
rect 24356 -20502 24608 -20486
rect 24814 -20486 24830 -20469
rect 25050 -20469 25140 -20452
rect 25198 -20452 25598 -20414
rect 25198 -20469 25288 -20452
rect 25050 -20486 25066 -20469
rect 24814 -20502 25066 -20486
rect 25272 -20486 25288 -20469
rect 25508 -20469 25598 -20452
rect 25656 -20452 26056 -20414
rect 25656 -20469 25746 -20452
rect 25508 -20486 25524 -20469
rect 25272 -20502 25524 -20486
rect 25730 -20486 25746 -20469
rect 25966 -20469 26056 -20452
rect 26114 -20452 26514 -20414
rect 26114 -20469 26204 -20452
rect 25966 -20486 25982 -20469
rect 25730 -20502 25982 -20486
rect 26188 -20486 26204 -20469
rect 26424 -20469 26514 -20452
rect 26572 -20452 26972 -20414
rect 26572 -20469 26662 -20452
rect 26424 -20486 26440 -20469
rect 26188 -20502 26440 -20486
rect 26646 -20486 26662 -20469
rect 26882 -20469 26972 -20452
rect 27030 -20452 27430 -20414
rect 27030 -20469 27120 -20452
rect 26882 -20486 26898 -20469
rect 26646 -20502 26898 -20486
rect 27104 -20486 27120 -20469
rect 27340 -20469 27430 -20452
rect 27488 -20452 27888 -20414
rect 27488 -20469 27578 -20452
rect 27340 -20486 27356 -20469
rect 27104 -20502 27356 -20486
rect 27562 -20486 27578 -20469
rect 27798 -20469 27888 -20452
rect 27946 -20452 28346 -20414
rect 27946 -20469 28036 -20452
rect 27798 -20486 27814 -20469
rect 27562 -20502 27814 -20486
rect 28020 -20486 28036 -20469
rect 28256 -20469 28346 -20452
rect 28824 -20452 29224 -20414
rect 28824 -20469 28914 -20452
rect 28256 -20486 28272 -20469
rect 28020 -20502 28272 -20486
rect 28898 -20486 28914 -20469
rect 29134 -20469 29224 -20452
rect 29282 -20452 29682 -20414
rect 29282 -20469 29372 -20452
rect 29134 -20486 29150 -20469
rect 28898 -20502 29150 -20486
rect 29356 -20486 29372 -20469
rect 29592 -20469 29682 -20452
rect 29740 -20452 30140 -20414
rect 29740 -20469 29830 -20452
rect 29592 -20486 29608 -20469
rect 29356 -20502 29608 -20486
rect 29814 -20486 29830 -20469
rect 30050 -20469 30140 -20452
rect 30198 -20452 30598 -20414
rect 30198 -20469 30288 -20452
rect 30050 -20486 30066 -20469
rect 29814 -20502 30066 -20486
rect 30272 -20486 30288 -20469
rect 30508 -20469 30598 -20452
rect 30656 -20452 31056 -20414
rect 30656 -20469 30746 -20452
rect 30508 -20486 30524 -20469
rect 30272 -20502 30524 -20486
rect 30730 -20486 30746 -20469
rect 30966 -20469 31056 -20452
rect 31114 -20452 31514 -20414
rect 31114 -20469 31204 -20452
rect 30966 -20486 30982 -20469
rect 30730 -20502 30982 -20486
rect 31188 -20486 31204 -20469
rect 31424 -20469 31514 -20452
rect 31572 -20452 31972 -20414
rect 31572 -20469 31662 -20452
rect 31424 -20486 31440 -20469
rect 31188 -20502 31440 -20486
rect 31646 -20486 31662 -20469
rect 31882 -20469 31972 -20452
rect 32030 -20452 32430 -20414
rect 32030 -20469 32120 -20452
rect 31882 -20486 31898 -20469
rect 31646 -20502 31898 -20486
rect 32104 -20486 32120 -20469
rect 32340 -20469 32430 -20452
rect 32488 -20452 32888 -20414
rect 32488 -20469 32578 -20452
rect 32340 -20486 32356 -20469
rect 32104 -20502 32356 -20486
rect 32562 -20486 32578 -20469
rect 32798 -20469 32888 -20452
rect 32946 -20452 33346 -20414
rect 32946 -20469 33036 -20452
rect 32798 -20486 32814 -20469
rect 32562 -20502 32814 -20486
rect 33020 -20486 33036 -20469
rect 33256 -20469 33346 -20452
rect 33256 -20486 33272 -20469
rect 33020 -20502 33272 -20486
rect 23898 -20810 24150 -20794
rect 23898 -20827 23914 -20810
rect 23824 -20844 23914 -20827
rect 24134 -20827 24150 -20810
rect 24356 -20810 24608 -20794
rect 24356 -20827 24372 -20810
rect 24134 -20844 24224 -20827
rect 23824 -20882 24224 -20844
rect 24282 -20844 24372 -20827
rect 24592 -20827 24608 -20810
rect 24814 -20810 25066 -20794
rect 24814 -20827 24830 -20810
rect 24592 -20844 24682 -20827
rect 24282 -20882 24682 -20844
rect 24740 -20844 24830 -20827
rect 25050 -20827 25066 -20810
rect 25272 -20810 25524 -20794
rect 25272 -20827 25288 -20810
rect 25050 -20844 25140 -20827
rect 24740 -20882 25140 -20844
rect 25198 -20844 25288 -20827
rect 25508 -20827 25524 -20810
rect 25730 -20810 25982 -20794
rect 25730 -20827 25746 -20810
rect 25508 -20844 25598 -20827
rect 25198 -20882 25598 -20844
rect 25656 -20844 25746 -20827
rect 25966 -20827 25982 -20810
rect 26188 -20810 26440 -20794
rect 26188 -20827 26204 -20810
rect 25966 -20844 26056 -20827
rect 25656 -20882 26056 -20844
rect 26114 -20844 26204 -20827
rect 26424 -20827 26440 -20810
rect 26646 -20810 26898 -20794
rect 26646 -20827 26662 -20810
rect 26424 -20844 26514 -20827
rect 26114 -20882 26514 -20844
rect 26572 -20844 26662 -20827
rect 26882 -20827 26898 -20810
rect 27104 -20810 27356 -20794
rect 27104 -20827 27120 -20810
rect 26882 -20844 26972 -20827
rect 26572 -20882 26972 -20844
rect 27030 -20844 27120 -20827
rect 27340 -20827 27356 -20810
rect 27562 -20810 27814 -20794
rect 27562 -20827 27578 -20810
rect 27340 -20844 27430 -20827
rect 27030 -20882 27430 -20844
rect 27488 -20844 27578 -20827
rect 27798 -20827 27814 -20810
rect 28020 -20810 28272 -20794
rect 28020 -20827 28036 -20810
rect 27798 -20844 27888 -20827
rect 27488 -20882 27888 -20844
rect 27946 -20844 28036 -20827
rect 28256 -20827 28272 -20810
rect 28256 -20844 28346 -20827
rect 27946 -20882 28346 -20844
rect 23824 -21120 24224 -21082
rect 23824 -21137 23914 -21120
rect 23898 -21154 23914 -21137
rect 24134 -21137 24224 -21120
rect 24282 -21120 24682 -21082
rect 24282 -21137 24372 -21120
rect 24134 -21154 24150 -21137
rect 23898 -21170 24150 -21154
rect 24356 -21154 24372 -21137
rect 24592 -21137 24682 -21120
rect 24740 -21120 25140 -21082
rect 24740 -21137 24830 -21120
rect 24592 -21154 24608 -21137
rect 24356 -21170 24608 -21154
rect 24814 -21154 24830 -21137
rect 25050 -21137 25140 -21120
rect 25198 -21120 25598 -21082
rect 25198 -21137 25288 -21120
rect 25050 -21154 25066 -21137
rect 24814 -21170 25066 -21154
rect 25272 -21154 25288 -21137
rect 25508 -21137 25598 -21120
rect 25656 -21120 26056 -21082
rect 25656 -21137 25746 -21120
rect 25508 -21154 25524 -21137
rect 25272 -21170 25524 -21154
rect 25730 -21154 25746 -21137
rect 25966 -21137 26056 -21120
rect 26114 -21120 26514 -21082
rect 26114 -21137 26204 -21120
rect 25966 -21154 25982 -21137
rect 25730 -21170 25982 -21154
rect 26188 -21154 26204 -21137
rect 26424 -21137 26514 -21120
rect 26572 -21120 26972 -21082
rect 26572 -21137 26662 -21120
rect 26424 -21154 26440 -21137
rect 26188 -21170 26440 -21154
rect 26646 -21154 26662 -21137
rect 26882 -21137 26972 -21120
rect 27030 -21120 27430 -21082
rect 27030 -21137 27120 -21120
rect 26882 -21154 26898 -21137
rect 26646 -21170 26898 -21154
rect 27104 -21154 27120 -21137
rect 27340 -21137 27430 -21120
rect 27488 -21120 27888 -21082
rect 27488 -21137 27578 -21120
rect 27340 -21154 27356 -21137
rect 27104 -21170 27356 -21154
rect 27562 -21154 27578 -21137
rect 27798 -21137 27888 -21120
rect 27946 -21120 28346 -21082
rect 27946 -21137 28036 -21120
rect 27798 -21154 27814 -21137
rect 27562 -21170 27814 -21154
rect 28020 -21154 28036 -21137
rect 28256 -21137 28346 -21120
rect 28256 -21154 28272 -21137
rect 28020 -21170 28272 -21154
<< polycont >>
rect 24030 16481 24414 16515
rect 24888 16481 25272 16515
rect 25746 16481 26130 16515
rect 26604 16481 26988 16515
rect 27462 16481 27846 16515
rect 28320 16481 28704 16515
rect 29178 16481 29562 16515
rect 30036 16481 30420 16515
rect 30894 16481 31278 16515
rect 31752 16481 32136 16515
rect 24030 16153 24414 16187
rect 24888 16153 25272 16187
rect 25746 16153 26130 16187
rect 26604 16153 26988 16187
rect 27462 16153 27846 16187
rect 28320 16153 28704 16187
rect 29178 16153 29562 16187
rect 30036 16153 30420 16187
rect 30894 16153 31278 16187
rect 31752 16153 32136 16187
rect 24030 15881 24414 15915
rect 24888 15881 25272 15915
rect 25746 15881 26130 15915
rect 26604 15881 26988 15915
rect 27462 15881 27846 15915
rect 28320 15881 28704 15915
rect 29178 15881 29562 15915
rect 30036 15881 30420 15915
rect 30894 15881 31278 15915
rect 31752 15881 32136 15915
rect 24030 15553 24414 15587
rect 24888 15553 25272 15587
rect 25746 15553 26130 15587
rect 26604 15553 26988 15587
rect 27462 15553 27846 15587
rect 28320 15553 28704 15587
rect 29178 15553 29562 15587
rect 30036 15553 30420 15587
rect 30894 15553 31278 15587
rect 31752 15553 32136 15587
rect 24259 14841 24359 14875
rect 24517 14841 24617 14875
rect 24775 14841 24875 14875
rect 24259 14313 24359 14347
rect 24517 14313 24617 14347
rect 24775 14313 24875 14347
rect 25381 14841 25481 14875
rect 25639 14841 25739 14875
rect 25897 14841 25997 14875
rect 26155 14841 26255 14875
rect 26413 14841 26513 14875
rect 26671 14841 26771 14875
rect 25381 14313 25481 14347
rect 25639 14313 25739 14347
rect 25897 14313 25997 14347
rect 26155 14313 26255 14347
rect 26413 14313 26513 14347
rect 26671 14313 26771 14347
rect 27292 14129 27326 14163
rect 27394 14144 27428 14178
rect 27782 14245 27816 14279
rect 27601 14190 27635 14224
rect 28031 14219 28065 14253
rect 24259 13945 24359 13979
rect 24517 13945 24617 13979
rect 24775 13945 24875 13979
rect 24259 13635 24359 13669
rect 24517 13635 24617 13669
rect 24775 13635 24875 13669
rect 25381 13945 25481 13979
rect 25639 13945 25739 13979
rect 25897 13945 25997 13979
rect 26155 13945 26255 13979
rect 26413 13945 26513 13979
rect 26671 13945 26771 13979
rect 27760 14083 27794 14117
rect 27862 14077 27896 14111
rect 25381 13635 25481 13669
rect 25639 13635 25739 13669
rect 25897 13635 25997 13669
rect 26155 13635 26255 13669
rect 26413 13635 26513 13669
rect 26671 13635 26771 13669
rect 28117 14083 28151 14117
rect 28213 14131 28247 14165
rect 28496 14245 28530 14279
rect 28361 14071 28395 14105
rect 28457 14119 28491 14153
rect 28774 14229 28808 14263
rect 28601 14093 28635 14127
rect 28697 14121 28731 14155
rect 28897 14129 28931 14163
rect 29237 14129 29271 14163
rect 29456 14129 29490 14163
rect 29688 14129 29722 14163
rect 30772 14229 30806 14263
rect 29856 14129 29890 14163
rect 30090 14129 30124 14163
rect 30309 14129 30343 14163
rect 30649 14129 30683 14163
rect 30849 14121 30883 14155
rect 31050 14245 31084 14279
rect 30945 14093 30979 14127
rect 31089 14119 31123 14153
rect 31333 14131 31367 14165
rect 31515 14219 31549 14253
rect 31185 14071 31219 14105
rect 31429 14083 31463 14117
rect 31764 14245 31798 14279
rect 31945 14190 31979 14224
rect 31684 14077 31718 14111
rect 31786 14083 31820 14117
rect 32152 14144 32186 14178
rect 32254 14129 32288 14163
rect 24466 12892 24926 12926
rect 25324 12892 25784 12926
rect 26182 12892 26642 12926
rect 27040 12892 27500 12926
rect 27898 12892 28358 12926
rect 28756 12892 29216 12926
rect 29614 12892 30074 12926
rect 30472 12892 30932 12926
rect 31330 12892 31790 12926
rect 24466 12582 24926 12616
rect 25324 12582 25784 12616
rect 26182 12582 26642 12616
rect 27040 12582 27500 12616
rect 27898 12582 28358 12616
rect 28756 12582 29216 12616
rect 29614 12582 30074 12616
rect 30472 12582 30932 12616
rect 31330 12582 31790 12616
rect 24466 12310 24926 12344
rect 25324 12310 25784 12344
rect 26182 12310 26642 12344
rect 27040 12310 27500 12344
rect 27898 12310 28358 12344
rect 28756 12310 29216 12344
rect 29614 12310 30074 12344
rect 30472 12310 30932 12344
rect 31330 12310 31790 12344
rect 24466 12000 24926 12034
rect 25324 12000 25784 12034
rect 26182 12000 26642 12034
rect 27040 12000 27500 12034
rect 27898 12000 28358 12034
rect 28756 12000 29216 12034
rect 29614 12000 30074 12034
rect 30472 12000 30932 12034
rect 31330 12000 31790 12034
rect 15304 9706 15524 9740
rect 15762 9706 15982 9740
rect 16220 9706 16440 9740
rect 16678 9706 16898 9740
rect 17136 9706 17356 9740
rect 17594 9706 17814 9740
rect 18052 9706 18272 9740
rect 18510 9706 18730 9740
rect 18968 9706 19188 9740
rect 19426 9706 19646 9740
rect 15304 9396 15524 9430
rect 15762 9396 15982 9430
rect 16220 9396 16440 9430
rect 16678 9396 16898 9430
rect 17136 9396 17356 9430
rect 17594 9396 17814 9430
rect 18052 9396 18272 9430
rect 18510 9396 18730 9430
rect 18968 9396 19188 9430
rect 19426 9396 19646 9430
rect 24066 9706 24286 9740
rect 24524 9706 24744 9740
rect 24982 9706 25202 9740
rect 25440 9706 25660 9740
rect 25898 9706 26118 9740
rect 26356 9706 26576 9740
rect 26814 9706 27034 9740
rect 27272 9706 27492 9740
rect 27730 9706 27950 9740
rect 28188 9706 28408 9740
rect 24066 9396 24286 9430
rect 24524 9396 24744 9430
rect 24982 9396 25202 9430
rect 25440 9396 25660 9430
rect 25898 9396 26118 9430
rect 26356 9396 26576 9430
rect 26814 9396 27034 9430
rect 27272 9396 27492 9430
rect 27730 9396 27950 9430
rect 28188 9396 28408 9430
rect 29156 8665 29190 8699
rect 29389 8665 29423 8699
rect 29481 8665 29515 8699
rect 29565 8665 29599 8699
rect 29649 8665 29683 8699
rect 13472 7864 13692 7898
rect 13930 7864 14150 7898
rect 14388 7864 14608 7898
rect 14846 7864 15066 7898
rect 15304 7864 15524 7898
rect 15762 7864 15982 7898
rect 16220 7864 16440 7898
rect 16678 7864 16898 7898
rect 17136 7864 17356 7898
rect 17594 7864 17814 7898
rect 18052 7864 18272 7898
rect 18510 7864 18730 7898
rect 18968 7864 19188 7898
rect 19426 7864 19646 7898
rect 19884 7864 20104 7898
rect 20342 7864 20562 7898
rect 20800 7864 21020 7898
rect 21258 7864 21478 7898
rect 13472 6136 13692 6170
rect 13930 6136 14150 6170
rect 14388 6136 14608 6170
rect 14846 6136 15066 6170
rect 15304 6136 15524 6170
rect 15762 6136 15982 6170
rect 16220 6136 16440 6170
rect 16678 6136 16898 6170
rect 17136 6136 17356 6170
rect 17594 6136 17814 6170
rect 18052 6136 18272 6170
rect 18510 6136 18730 6170
rect 18968 6136 19188 6170
rect 19426 6136 19646 6170
rect 19884 6136 20104 6170
rect 20342 6136 20562 6170
rect 20800 6136 21020 6170
rect 21258 6136 21478 6170
rect 30584 8631 30618 8665
rect 30848 8699 30882 8733
rect 31100 8747 31134 8781
rect 30686 8646 30720 8680
rect 24067 8284 24287 8318
rect 24525 8284 24745 8318
rect 24983 8284 25203 8318
rect 25441 8284 25661 8318
rect 25899 8284 26119 8318
rect 26357 8284 26577 8318
rect 26815 8284 27035 8318
rect 27273 8284 27493 8318
rect 27731 8284 27951 8318
rect 28189 8284 28409 8318
rect 24067 6956 24287 6990
rect 24525 6956 24745 6990
rect 24983 6956 25203 6990
rect 25441 6956 25661 6990
rect 25899 6956 26119 6990
rect 26357 6956 26577 6990
rect 26815 6956 27035 6990
rect 27273 6956 27493 6990
rect 27731 6956 27951 6990
rect 28189 6956 28409 6990
rect 30991 8669 31025 8703
rect 31011 8573 31045 8607
rect 31512 8747 31546 8781
rect 31648 8747 31682 8781
rect 31274 8681 31308 8715
rect 31410 8681 31444 8715
rect 31210 8585 31244 8619
rect 31453 8573 31487 8607
rect 31722 8631 31756 8665
rect 31906 8631 31940 8665
rect 32167 8631 32201 8665
rect 32380 8631 32414 8665
rect 32613 8631 32647 8665
rect 32705 8631 32739 8665
rect 32789 8631 32823 8665
rect 32873 8631 32907 8665
rect 30584 8167 30618 8201
rect 30686 8152 30720 8186
rect 31011 8225 31045 8259
rect 30848 8099 30882 8133
rect 30991 8129 31025 8163
rect 31210 8213 31244 8247
rect 31100 8051 31134 8085
rect 31453 8225 31487 8259
rect 31274 8117 31308 8151
rect 31410 8117 31444 8151
rect 31722 8167 31756 8201
rect 31906 8167 31940 8201
rect 32167 8167 32201 8201
rect 32380 8167 32414 8201
rect 32613 8167 32647 8201
rect 32705 8167 32739 8201
rect 32789 8167 32823 8201
rect 32873 8167 32907 8201
rect 33282 8167 33316 8201
rect 31512 8051 31546 8085
rect 31648 8051 31682 8085
rect 33384 8152 33418 8186
rect 33709 8225 33743 8259
rect 33546 8099 33580 8133
rect 33689 8129 33723 8163
rect 33908 8213 33942 8247
rect 33798 8051 33832 8085
rect 34151 8225 34185 8259
rect 33972 8117 34006 8151
rect 34108 8117 34142 8151
rect 34420 8167 34454 8201
rect 34604 8167 34638 8201
rect 34865 8167 34899 8201
rect 35078 8167 35112 8201
rect 35311 8167 35345 8201
rect 35403 8167 35437 8201
rect 35487 8167 35521 8201
rect 35571 8167 35605 8201
rect 34210 8051 34244 8085
rect 34346 8051 34380 8085
rect 30584 7543 30618 7577
rect 30848 7611 30882 7645
rect 31100 7659 31134 7693
rect 30686 7558 30720 7592
rect 30991 7581 31025 7615
rect 31011 7485 31045 7519
rect 31512 7659 31546 7693
rect 31648 7659 31682 7693
rect 31274 7593 31308 7627
rect 31410 7593 31444 7627
rect 31210 7497 31244 7531
rect 31453 7485 31487 7519
rect 31722 7543 31756 7577
rect 31906 7543 31940 7577
rect 32167 7543 32201 7577
rect 32380 7543 32414 7577
rect 32613 7543 32647 7577
rect 32705 7543 32739 7577
rect 32789 7543 32823 7577
rect 32873 7543 32907 7577
rect 33282 7543 33316 7577
rect 33546 7611 33580 7645
rect 33798 7659 33832 7693
rect 33384 7558 33418 7592
rect 33689 7581 33723 7615
rect 33709 7485 33743 7519
rect 34210 7659 34244 7693
rect 34346 7659 34380 7693
rect 33972 7593 34006 7627
rect 34108 7593 34142 7627
rect 33908 7497 33942 7531
rect 34151 7485 34185 7519
rect 34420 7543 34454 7577
rect 34604 7543 34638 7577
rect 34865 7543 34899 7577
rect 35078 7543 35112 7577
rect 35311 7543 35345 7577
rect 35403 7543 35437 7577
rect 35487 7543 35521 7577
rect 35571 7543 35605 7577
rect 30584 7079 30618 7113
rect 30686 7064 30720 7098
rect 31011 7137 31045 7171
rect 30848 7011 30882 7045
rect 30991 7041 31025 7075
rect 31210 7125 31244 7159
rect 31100 6963 31134 6997
rect 31453 7137 31487 7171
rect 31274 7029 31308 7063
rect 31410 7029 31444 7063
rect 31722 7079 31756 7113
rect 31906 7079 31940 7113
rect 32167 7079 32201 7113
rect 32380 7079 32414 7113
rect 32613 7079 32647 7113
rect 32705 7079 32739 7113
rect 32789 7079 32823 7113
rect 32873 7079 32907 7113
rect 33282 7079 33316 7113
rect 31512 6963 31546 6997
rect 31648 6963 31682 6997
rect 33384 7064 33418 7098
rect 33709 7137 33743 7171
rect 33546 7011 33580 7045
rect 33689 7041 33723 7075
rect 33908 7125 33942 7159
rect 33798 6963 33832 6997
rect 34151 7137 34185 7171
rect 33972 7029 34006 7063
rect 34108 7029 34142 7063
rect 34420 7079 34454 7113
rect 34604 7079 34638 7113
rect 34865 7079 34899 7113
rect 35078 7079 35112 7113
rect 35311 7079 35345 7113
rect 35403 7079 35437 7113
rect 35487 7079 35521 7113
rect 35571 7079 35605 7113
rect 34210 6963 34244 6997
rect 34346 6963 34380 6997
rect 30584 6455 30618 6489
rect 30848 6523 30882 6557
rect 31100 6571 31134 6605
rect 30686 6470 30720 6504
rect 30991 6493 31025 6527
rect 31011 6397 31045 6431
rect 31512 6571 31546 6605
rect 31648 6571 31682 6605
rect 31274 6505 31308 6539
rect 31410 6505 31444 6539
rect 31210 6409 31244 6443
rect 31453 6397 31487 6431
rect 31722 6455 31756 6489
rect 31906 6455 31940 6489
rect 32167 6455 32201 6489
rect 32380 6455 32414 6489
rect 32613 6455 32647 6489
rect 32705 6455 32739 6489
rect 32789 6455 32823 6489
rect 32873 6455 32907 6489
rect 33282 6455 33316 6489
rect 33546 6523 33580 6557
rect 33798 6571 33832 6605
rect 33384 6470 33418 6504
rect 33689 6493 33723 6527
rect 33709 6397 33743 6431
rect 34210 6571 34244 6605
rect 34346 6571 34380 6605
rect 33972 6505 34006 6539
rect 34108 6505 34142 6539
rect 33908 6409 33942 6443
rect 34151 6397 34185 6431
rect 34420 6455 34454 6489
rect 34604 6455 34638 6489
rect 34865 6455 34899 6489
rect 35078 6455 35112 6489
rect 35311 6455 35345 6489
rect 35403 6455 35437 6489
rect 35487 6455 35521 6489
rect 35571 6455 35605 6489
rect 30584 5991 30618 6025
rect 30686 5976 30720 6010
rect 31011 6049 31045 6083
rect 30848 5923 30882 5957
rect 30991 5953 31025 5987
rect 31210 6037 31244 6071
rect 31100 5875 31134 5909
rect 31453 6049 31487 6083
rect 31274 5941 31308 5975
rect 31410 5941 31444 5975
rect 31722 5991 31756 6025
rect 31906 5991 31940 6025
rect 32167 5991 32201 6025
rect 32380 5991 32414 6025
rect 32613 5991 32647 6025
rect 32705 5991 32739 6025
rect 32789 5991 32823 6025
rect 32873 5991 32907 6025
rect 33282 5991 33316 6025
rect 31512 5875 31546 5909
rect 31648 5875 31682 5909
rect 33384 5976 33418 6010
rect 33709 6049 33743 6083
rect 33546 5923 33580 5957
rect 33689 5953 33723 5987
rect 33908 6037 33942 6071
rect 33798 5875 33832 5909
rect 34151 6049 34185 6083
rect 33972 5941 34006 5975
rect 34108 5941 34142 5975
rect 34420 5991 34454 6025
rect 34604 5991 34638 6025
rect 34865 5991 34899 6025
rect 35078 5991 35112 6025
rect 35311 5991 35345 6025
rect 35403 5991 35437 6025
rect 35487 5991 35521 6025
rect 35571 5991 35605 6025
rect 34210 5875 34244 5909
rect 34346 5875 34380 5909
rect 9474 2991 9694 3025
rect 9932 2991 10152 3025
rect 10390 2991 10610 3025
rect 10848 2991 11068 3025
rect 11306 2991 11526 3025
rect 11764 2991 11984 3025
rect 12222 2991 12442 3025
rect 12680 2991 12900 3025
rect 13138 2991 13358 3025
rect 13596 2991 13816 3025
rect 14054 2991 14274 3025
rect 14512 2991 14732 3025
rect 14970 2991 15190 3025
rect 15428 2991 15648 3025
rect 15886 2991 16106 3025
rect 16344 2991 16564 3025
rect 16802 2991 17022 3025
rect 17260 2991 17480 3025
rect 9474 1263 9694 1297
rect 9932 1263 10152 1297
rect 10390 1263 10610 1297
rect 10848 1263 11068 1297
rect 11306 1263 11526 1297
rect 11764 1263 11984 1297
rect 12222 1263 12442 1297
rect 12680 1263 12900 1297
rect 13138 1263 13358 1297
rect 13596 1263 13816 1297
rect 14054 1263 14274 1297
rect 14512 1263 14732 1297
rect 14970 1263 15190 1297
rect 15428 1263 15648 1297
rect 15886 1263 16106 1297
rect 16344 1263 16564 1297
rect 16802 1263 17022 1297
rect 17260 1263 17480 1297
rect 8915 326 9135 360
rect 9373 326 9593 360
rect 9831 326 10051 360
rect 10289 326 10509 360
rect 10747 326 10967 360
rect 11205 326 11425 360
rect 11663 326 11883 360
rect 12121 326 12341 360
rect 12579 326 12799 360
rect 13037 326 13257 360
rect 13915 326 14135 360
rect 14373 326 14593 360
rect 14831 326 15051 360
rect 15289 326 15509 360
rect 15747 326 15967 360
rect 16205 326 16425 360
rect 16663 326 16883 360
rect 17121 326 17341 360
rect 17579 326 17799 360
rect 18037 326 18257 360
rect 8915 -1002 9135 -968
rect 9373 -1002 9593 -968
rect 9831 -1002 10051 -968
rect 10289 -1002 10509 -968
rect 10747 -1002 10967 -968
rect 11205 -1002 11425 -968
rect 11663 -1002 11883 -968
rect 12121 -1002 12341 -968
rect 12579 -1002 12799 -968
rect 13037 -1002 13257 -968
rect 13915 -1002 14135 -968
rect 14373 -1002 14593 -968
rect 14831 -1002 15051 -968
rect 15289 -1002 15509 -968
rect 15747 -1002 15967 -968
rect 16205 -1002 16425 -968
rect 16663 -1002 16883 -968
rect 17121 -1002 17341 -968
rect 17579 -1002 17799 -968
rect 18037 -1002 18257 -968
rect 24474 2991 24694 3025
rect 24932 2991 25152 3025
rect 25390 2991 25610 3025
rect 25848 2991 26068 3025
rect 26306 2991 26526 3025
rect 26764 2991 26984 3025
rect 27222 2991 27442 3025
rect 27680 2991 27900 3025
rect 28138 2991 28358 3025
rect 28596 2991 28816 3025
rect 29054 2991 29274 3025
rect 29512 2991 29732 3025
rect 29970 2991 30190 3025
rect 30428 2991 30648 3025
rect 30886 2991 31106 3025
rect 31344 2991 31564 3025
rect 31802 2991 32022 3025
rect 32260 2991 32480 3025
rect 24474 1263 24694 1297
rect 24932 1263 25152 1297
rect 25390 1263 25610 1297
rect 25848 1263 26068 1297
rect 26306 1263 26526 1297
rect 26764 1263 26984 1297
rect 27222 1263 27442 1297
rect 27680 1263 27900 1297
rect 28138 1263 28358 1297
rect 28596 1263 28816 1297
rect 29054 1263 29274 1297
rect 29512 1263 29732 1297
rect 29970 1263 30190 1297
rect 30428 1263 30648 1297
rect 30886 1263 31106 1297
rect 31344 1263 31564 1297
rect 31802 1263 32022 1297
rect 32260 1263 32480 1297
rect 23915 326 24135 360
rect 24373 326 24593 360
rect 24831 326 25051 360
rect 25289 326 25509 360
rect 25747 326 25967 360
rect 26205 326 26425 360
rect 26663 326 26883 360
rect 27121 326 27341 360
rect 27579 326 27799 360
rect 28037 326 28257 360
rect 28915 326 29135 360
rect 29373 326 29593 360
rect 29831 326 30051 360
rect 30289 326 30509 360
rect 30747 326 30967 360
rect 31205 326 31425 360
rect 31663 326 31883 360
rect 32121 326 32341 360
rect 32579 326 32799 360
rect 33037 326 33257 360
rect 23915 -1002 24135 -968
rect 24373 -1002 24593 -968
rect 24831 -1002 25051 -968
rect 25289 -1002 25509 -968
rect 25747 -1002 25967 -968
rect 26205 -1002 26425 -968
rect 26663 -1002 26883 -968
rect 27121 -1002 27341 -968
rect 27579 -1002 27799 -968
rect 28037 -1002 28257 -968
rect 28915 -1002 29135 -968
rect 29373 -1002 29593 -968
rect 29831 -1002 30051 -968
rect 30289 -1002 30509 -968
rect 30747 -1002 30967 -968
rect 31205 -1002 31425 -968
rect 31663 -1002 31883 -968
rect 32121 -1002 32341 -968
rect 32579 -1002 32799 -968
rect 33037 -1002 33257 -968
rect 8914 -2176 9134 -2142
rect 9372 -2176 9592 -2142
rect 9830 -2176 10050 -2142
rect 10288 -2176 10508 -2142
rect 10746 -2176 10966 -2142
rect 11204 -2176 11424 -2142
rect 11662 -2176 11882 -2142
rect 12120 -2176 12340 -2142
rect 12578 -2176 12798 -2142
rect 13036 -2176 13256 -2142
rect 13914 -2176 14134 -2142
rect 14372 -2176 14592 -2142
rect 14830 -2176 15050 -2142
rect 15288 -2176 15508 -2142
rect 15746 -2176 15966 -2142
rect 16204 -2176 16424 -2142
rect 16662 -2176 16882 -2142
rect 17120 -2176 17340 -2142
rect 17578 -2176 17798 -2142
rect 18036 -2176 18256 -2142
rect 8914 -2486 9134 -2452
rect 9372 -2486 9592 -2452
rect 9830 -2486 10050 -2452
rect 10288 -2486 10508 -2452
rect 10746 -2486 10966 -2452
rect 11204 -2486 11424 -2452
rect 11662 -2486 11882 -2452
rect 12120 -2486 12340 -2452
rect 12578 -2486 12798 -2452
rect 13036 -2486 13256 -2452
rect 13914 -2486 14134 -2452
rect 14372 -2486 14592 -2452
rect 14830 -2486 15050 -2452
rect 15288 -2486 15508 -2452
rect 15746 -2486 15966 -2452
rect 16204 -2486 16424 -2452
rect 16662 -2486 16882 -2452
rect 17120 -2486 17340 -2452
rect 17578 -2486 17798 -2452
rect 18036 -2486 18256 -2452
rect 8914 -2844 9134 -2810
rect 9372 -2844 9592 -2810
rect 9830 -2844 10050 -2810
rect 10288 -2844 10508 -2810
rect 10746 -2844 10966 -2810
rect 11204 -2844 11424 -2810
rect 11662 -2844 11882 -2810
rect 12120 -2844 12340 -2810
rect 12578 -2844 12798 -2810
rect 13036 -2844 13256 -2810
rect 8914 -3154 9134 -3120
rect 9372 -3154 9592 -3120
rect 9830 -3154 10050 -3120
rect 10288 -3154 10508 -3120
rect 10746 -3154 10966 -3120
rect 11204 -3154 11424 -3120
rect 11662 -3154 11882 -3120
rect 12120 -3154 12340 -3120
rect 12578 -3154 12798 -3120
rect 13036 -3154 13256 -3120
rect 23914 -2176 24134 -2142
rect 24372 -2176 24592 -2142
rect 24830 -2176 25050 -2142
rect 25288 -2176 25508 -2142
rect 25746 -2176 25966 -2142
rect 26204 -2176 26424 -2142
rect 26662 -2176 26882 -2142
rect 27120 -2176 27340 -2142
rect 27578 -2176 27798 -2142
rect 28036 -2176 28256 -2142
rect 28914 -2176 29134 -2142
rect 29372 -2176 29592 -2142
rect 29830 -2176 30050 -2142
rect 30288 -2176 30508 -2142
rect 30746 -2176 30966 -2142
rect 31204 -2176 31424 -2142
rect 31662 -2176 31882 -2142
rect 32120 -2176 32340 -2142
rect 32578 -2176 32798 -2142
rect 33036 -2176 33256 -2142
rect 23914 -2486 24134 -2452
rect 24372 -2486 24592 -2452
rect 24830 -2486 25050 -2452
rect 25288 -2486 25508 -2452
rect 25746 -2486 25966 -2452
rect 26204 -2486 26424 -2452
rect 26662 -2486 26882 -2452
rect 27120 -2486 27340 -2452
rect 27578 -2486 27798 -2452
rect 28036 -2486 28256 -2452
rect 28914 -2486 29134 -2452
rect 29372 -2486 29592 -2452
rect 29830 -2486 30050 -2452
rect 30288 -2486 30508 -2452
rect 30746 -2486 30966 -2452
rect 31204 -2486 31424 -2452
rect 31662 -2486 31882 -2452
rect 32120 -2486 32340 -2452
rect 32578 -2486 32798 -2452
rect 33036 -2486 33256 -2452
rect 23914 -2844 24134 -2810
rect 24372 -2844 24592 -2810
rect 24830 -2844 25050 -2810
rect 25288 -2844 25508 -2810
rect 25746 -2844 25966 -2810
rect 26204 -2844 26424 -2810
rect 26662 -2844 26882 -2810
rect 27120 -2844 27340 -2810
rect 27578 -2844 27798 -2810
rect 28036 -2844 28256 -2810
rect 23914 -3154 24134 -3120
rect 24372 -3154 24592 -3120
rect 24830 -3154 25050 -3120
rect 25288 -3154 25508 -3120
rect 25746 -3154 25966 -3120
rect 26204 -3154 26424 -3120
rect 26662 -3154 26882 -3120
rect 27120 -3154 27340 -3120
rect 27578 -3154 27798 -3120
rect 28036 -3154 28256 -3120
rect 17846 -5636 18066 -5602
rect 18304 -5636 18524 -5602
rect 18762 -5636 18982 -5602
rect 19220 -5636 19440 -5602
rect 19678 -5636 19898 -5602
rect 20136 -5636 20356 -5602
rect 20594 -5636 20814 -5602
rect 21052 -5636 21272 -5602
rect 21510 -5636 21730 -5602
rect 21968 -5636 22188 -5602
rect 17846 -5946 18066 -5912
rect 18304 -5946 18524 -5912
rect 18762 -5946 18982 -5912
rect 19220 -5946 19440 -5912
rect 19678 -5946 19898 -5912
rect 20136 -5946 20356 -5912
rect 20594 -5946 20814 -5912
rect 21052 -5946 21272 -5912
rect 21510 -5946 21730 -5912
rect 21968 -5946 22188 -5912
rect 12846 -6304 13066 -6270
rect 13304 -6304 13524 -6270
rect 13762 -6304 13982 -6270
rect 14220 -6304 14440 -6270
rect 14678 -6304 14898 -6270
rect 15136 -6304 15356 -6270
rect 15594 -6304 15814 -6270
rect 16052 -6304 16272 -6270
rect 16510 -6304 16730 -6270
rect 16968 -6304 17188 -6270
rect 17846 -6304 18066 -6270
rect 18304 -6304 18524 -6270
rect 18762 -6304 18982 -6270
rect 19220 -6304 19440 -6270
rect 19678 -6304 19898 -6270
rect 20136 -6304 20356 -6270
rect 20594 -6304 20814 -6270
rect 21052 -6304 21272 -6270
rect 21510 -6304 21730 -6270
rect 21968 -6304 22188 -6270
rect 12846 -6614 13066 -6580
rect 13304 -6614 13524 -6580
rect 13762 -6614 13982 -6580
rect 14220 -6614 14440 -6580
rect 14678 -6614 14898 -6580
rect 15136 -6614 15356 -6580
rect 15594 -6614 15814 -6580
rect 16052 -6614 16272 -6580
rect 16510 -6614 16730 -6580
rect 16968 -6614 17188 -6580
rect 17846 -6614 18066 -6580
rect 18304 -6614 18524 -6580
rect 18762 -6614 18982 -6580
rect 19220 -6614 19440 -6580
rect 19678 -6614 19898 -6580
rect 20136 -6614 20356 -6580
rect 20594 -6614 20814 -6580
rect 21052 -6614 21272 -6580
rect 21510 -6614 21730 -6580
rect 21968 -6614 22188 -6580
rect 32846 -5636 33066 -5602
rect 33304 -5636 33524 -5602
rect 33762 -5636 33982 -5602
rect 34220 -5636 34440 -5602
rect 34678 -5636 34898 -5602
rect 35136 -5636 35356 -5602
rect 35594 -5636 35814 -5602
rect 36052 -5636 36272 -5602
rect 36510 -5636 36730 -5602
rect 36968 -5636 37188 -5602
rect 32846 -5946 33066 -5912
rect 33304 -5946 33524 -5912
rect 33762 -5946 33982 -5912
rect 34220 -5946 34440 -5912
rect 34678 -5946 34898 -5912
rect 35136 -5946 35356 -5912
rect 35594 -5946 35814 -5912
rect 36052 -5946 36272 -5912
rect 36510 -5946 36730 -5912
rect 36968 -5946 37188 -5912
rect 27846 -6304 28066 -6270
rect 28304 -6304 28524 -6270
rect 28762 -6304 28982 -6270
rect 29220 -6304 29440 -6270
rect 29678 -6304 29898 -6270
rect 30136 -6304 30356 -6270
rect 30594 -6304 30814 -6270
rect 31052 -6304 31272 -6270
rect 31510 -6304 31730 -6270
rect 31968 -6304 32188 -6270
rect 32846 -6304 33066 -6270
rect 33304 -6304 33524 -6270
rect 33762 -6304 33982 -6270
rect 34220 -6304 34440 -6270
rect 34678 -6304 34898 -6270
rect 35136 -6304 35356 -6270
rect 35594 -6304 35814 -6270
rect 36052 -6304 36272 -6270
rect 36510 -6304 36730 -6270
rect 36968 -6304 37188 -6270
rect 27846 -6614 28066 -6580
rect 28304 -6614 28524 -6580
rect 28762 -6614 28982 -6580
rect 29220 -6614 29440 -6580
rect 29678 -6614 29898 -6580
rect 30136 -6614 30356 -6580
rect 30594 -6614 30814 -6580
rect 31052 -6614 31272 -6580
rect 31510 -6614 31730 -6580
rect 31968 -6614 32188 -6580
rect 32846 -6614 33066 -6580
rect 33304 -6614 33524 -6580
rect 33762 -6614 33982 -6580
rect 34220 -6614 34440 -6580
rect 34678 -6614 34898 -6580
rect 35136 -6614 35356 -6580
rect 35594 -6614 35814 -6580
rect 36052 -6614 36272 -6580
rect 36510 -6614 36730 -6580
rect 36968 -6614 37188 -6580
rect 12845 -7788 13065 -7754
rect 13303 -7788 13523 -7754
rect 13761 -7788 13981 -7754
rect 14219 -7788 14439 -7754
rect 14677 -7788 14897 -7754
rect 15135 -7788 15355 -7754
rect 15593 -7788 15813 -7754
rect 16051 -7788 16271 -7754
rect 16509 -7788 16729 -7754
rect 16967 -7788 17187 -7754
rect 17845 -7788 18065 -7754
rect 18303 -7788 18523 -7754
rect 18761 -7788 18981 -7754
rect 19219 -7788 19439 -7754
rect 19677 -7788 19897 -7754
rect 20135 -7788 20355 -7754
rect 20593 -7788 20813 -7754
rect 21051 -7788 21271 -7754
rect 21509 -7788 21729 -7754
rect 21967 -7788 22187 -7754
rect 12845 -9116 13065 -9082
rect 13303 -9116 13523 -9082
rect 13761 -9116 13981 -9082
rect 14219 -9116 14439 -9082
rect 14677 -9116 14897 -9082
rect 15135 -9116 15355 -9082
rect 15593 -9116 15813 -9082
rect 16051 -9116 16271 -9082
rect 16509 -9116 16729 -9082
rect 16967 -9116 17187 -9082
rect 17845 -9116 18065 -9082
rect 18303 -9116 18523 -9082
rect 18761 -9116 18981 -9082
rect 19219 -9116 19439 -9082
rect 19677 -9116 19897 -9082
rect 20135 -9116 20355 -9082
rect 20593 -9116 20813 -9082
rect 21051 -9116 21271 -9082
rect 21509 -9116 21729 -9082
rect 21967 -9116 22187 -9082
rect 13622 -10053 13842 -10019
rect 14080 -10053 14300 -10019
rect 14538 -10053 14758 -10019
rect 14996 -10053 15216 -10019
rect 15454 -10053 15674 -10019
rect 15912 -10053 16132 -10019
rect 16370 -10053 16590 -10019
rect 16828 -10053 17048 -10019
rect 17286 -10053 17506 -10019
rect 17744 -10053 17964 -10019
rect 18202 -10053 18422 -10019
rect 18660 -10053 18880 -10019
rect 19118 -10053 19338 -10019
rect 19576 -10053 19796 -10019
rect 20034 -10053 20254 -10019
rect 20492 -10053 20712 -10019
rect 20950 -10053 21170 -10019
rect 21408 -10053 21628 -10019
rect 13622 -11781 13842 -11747
rect 14080 -11781 14300 -11747
rect 14538 -11781 14758 -11747
rect 14996 -11781 15216 -11747
rect 15454 -11781 15674 -11747
rect 15912 -11781 16132 -11747
rect 16370 -11781 16590 -11747
rect 16828 -11781 17048 -11747
rect 17286 -11781 17506 -11747
rect 17744 -11781 17964 -11747
rect 18202 -11781 18422 -11747
rect 18660 -11781 18880 -11747
rect 19118 -11781 19338 -11747
rect 19576 -11781 19796 -11747
rect 20034 -11781 20254 -11747
rect 20492 -11781 20712 -11747
rect 20950 -11781 21170 -11747
rect 21408 -11781 21628 -11747
rect 27845 -7788 28065 -7754
rect 28303 -7788 28523 -7754
rect 28761 -7788 28981 -7754
rect 29219 -7788 29439 -7754
rect 29677 -7788 29897 -7754
rect 30135 -7788 30355 -7754
rect 30593 -7788 30813 -7754
rect 31051 -7788 31271 -7754
rect 31509 -7788 31729 -7754
rect 31967 -7788 32187 -7754
rect 32845 -7788 33065 -7754
rect 33303 -7788 33523 -7754
rect 33761 -7788 33981 -7754
rect 34219 -7788 34439 -7754
rect 34677 -7788 34897 -7754
rect 35135 -7788 35355 -7754
rect 35593 -7788 35813 -7754
rect 36051 -7788 36271 -7754
rect 36509 -7788 36729 -7754
rect 36967 -7788 37187 -7754
rect 27845 -9116 28065 -9082
rect 28303 -9116 28523 -9082
rect 28761 -9116 28981 -9082
rect 29219 -9116 29439 -9082
rect 29677 -9116 29897 -9082
rect 30135 -9116 30355 -9082
rect 30593 -9116 30813 -9082
rect 31051 -9116 31271 -9082
rect 31509 -9116 31729 -9082
rect 31967 -9116 32187 -9082
rect 32845 -9116 33065 -9082
rect 33303 -9116 33523 -9082
rect 33761 -9116 33981 -9082
rect 34219 -9116 34439 -9082
rect 34677 -9116 34897 -9082
rect 35135 -9116 35355 -9082
rect 35593 -9116 35813 -9082
rect 36051 -9116 36271 -9082
rect 36509 -9116 36729 -9082
rect 36967 -9116 37187 -9082
rect 28622 -10053 28842 -10019
rect 29080 -10053 29300 -10019
rect 29538 -10053 29758 -10019
rect 29996 -10053 30216 -10019
rect 30454 -10053 30674 -10019
rect 30912 -10053 31132 -10019
rect 31370 -10053 31590 -10019
rect 31828 -10053 32048 -10019
rect 32286 -10053 32506 -10019
rect 32744 -10053 32964 -10019
rect 33202 -10053 33422 -10019
rect 33660 -10053 33880 -10019
rect 34118 -10053 34338 -10019
rect 34576 -10053 34796 -10019
rect 35034 -10053 35254 -10019
rect 35492 -10053 35712 -10019
rect 35950 -10053 36170 -10019
rect 36408 -10053 36628 -10019
rect 28622 -11781 28842 -11747
rect 29080 -11781 29300 -11747
rect 29538 -11781 29758 -11747
rect 29996 -11781 30216 -11747
rect 30454 -11781 30674 -11747
rect 30912 -11781 31132 -11747
rect 31370 -11781 31590 -11747
rect 31828 -11781 32048 -11747
rect 32286 -11781 32506 -11747
rect 32744 -11781 32964 -11747
rect 33202 -11781 33422 -11747
rect 33660 -11781 33880 -11747
rect 34118 -11781 34338 -11747
rect 34576 -11781 34796 -11747
rect 35034 -11781 35254 -11747
rect 35492 -11781 35712 -11747
rect 35950 -11781 36170 -11747
rect 36408 -11781 36628 -11747
rect 9474 -15009 9694 -14975
rect 9932 -15009 10152 -14975
rect 10390 -15009 10610 -14975
rect 10848 -15009 11068 -14975
rect 11306 -15009 11526 -14975
rect 11764 -15009 11984 -14975
rect 12222 -15009 12442 -14975
rect 12680 -15009 12900 -14975
rect 13138 -15009 13358 -14975
rect 13596 -15009 13816 -14975
rect 14054 -15009 14274 -14975
rect 14512 -15009 14732 -14975
rect 14970 -15009 15190 -14975
rect 15428 -15009 15648 -14975
rect 15886 -15009 16106 -14975
rect 16344 -15009 16564 -14975
rect 16802 -15009 17022 -14975
rect 17260 -15009 17480 -14975
rect 9474 -16737 9694 -16703
rect 9932 -16737 10152 -16703
rect 10390 -16737 10610 -16703
rect 10848 -16737 11068 -16703
rect 11306 -16737 11526 -16703
rect 11764 -16737 11984 -16703
rect 12222 -16737 12442 -16703
rect 12680 -16737 12900 -16703
rect 13138 -16737 13358 -16703
rect 13596 -16737 13816 -16703
rect 14054 -16737 14274 -16703
rect 14512 -16737 14732 -16703
rect 14970 -16737 15190 -16703
rect 15428 -16737 15648 -16703
rect 15886 -16737 16106 -16703
rect 16344 -16737 16564 -16703
rect 16802 -16737 17022 -16703
rect 17260 -16737 17480 -16703
rect 8915 -17674 9135 -17640
rect 9373 -17674 9593 -17640
rect 9831 -17674 10051 -17640
rect 10289 -17674 10509 -17640
rect 10747 -17674 10967 -17640
rect 11205 -17674 11425 -17640
rect 11663 -17674 11883 -17640
rect 12121 -17674 12341 -17640
rect 12579 -17674 12799 -17640
rect 13037 -17674 13257 -17640
rect 13915 -17674 14135 -17640
rect 14373 -17674 14593 -17640
rect 14831 -17674 15051 -17640
rect 15289 -17674 15509 -17640
rect 15747 -17674 15967 -17640
rect 16205 -17674 16425 -17640
rect 16663 -17674 16883 -17640
rect 17121 -17674 17341 -17640
rect 17579 -17674 17799 -17640
rect 18037 -17674 18257 -17640
rect 8915 -19002 9135 -18968
rect 9373 -19002 9593 -18968
rect 9831 -19002 10051 -18968
rect 10289 -19002 10509 -18968
rect 10747 -19002 10967 -18968
rect 11205 -19002 11425 -18968
rect 11663 -19002 11883 -18968
rect 12121 -19002 12341 -18968
rect 12579 -19002 12799 -18968
rect 13037 -19002 13257 -18968
rect 13915 -19002 14135 -18968
rect 14373 -19002 14593 -18968
rect 14831 -19002 15051 -18968
rect 15289 -19002 15509 -18968
rect 15747 -19002 15967 -18968
rect 16205 -19002 16425 -18968
rect 16663 -19002 16883 -18968
rect 17121 -19002 17341 -18968
rect 17579 -19002 17799 -18968
rect 18037 -19002 18257 -18968
rect 24474 -15009 24694 -14975
rect 24932 -15009 25152 -14975
rect 25390 -15009 25610 -14975
rect 25848 -15009 26068 -14975
rect 26306 -15009 26526 -14975
rect 26764 -15009 26984 -14975
rect 27222 -15009 27442 -14975
rect 27680 -15009 27900 -14975
rect 28138 -15009 28358 -14975
rect 28596 -15009 28816 -14975
rect 29054 -15009 29274 -14975
rect 29512 -15009 29732 -14975
rect 29970 -15009 30190 -14975
rect 30428 -15009 30648 -14975
rect 30886 -15009 31106 -14975
rect 31344 -15009 31564 -14975
rect 31802 -15009 32022 -14975
rect 32260 -15009 32480 -14975
rect 24474 -16737 24694 -16703
rect 24932 -16737 25152 -16703
rect 25390 -16737 25610 -16703
rect 25848 -16737 26068 -16703
rect 26306 -16737 26526 -16703
rect 26764 -16737 26984 -16703
rect 27222 -16737 27442 -16703
rect 27680 -16737 27900 -16703
rect 28138 -16737 28358 -16703
rect 28596 -16737 28816 -16703
rect 29054 -16737 29274 -16703
rect 29512 -16737 29732 -16703
rect 29970 -16737 30190 -16703
rect 30428 -16737 30648 -16703
rect 30886 -16737 31106 -16703
rect 31344 -16737 31564 -16703
rect 31802 -16737 32022 -16703
rect 32260 -16737 32480 -16703
rect 23915 -17674 24135 -17640
rect 24373 -17674 24593 -17640
rect 24831 -17674 25051 -17640
rect 25289 -17674 25509 -17640
rect 25747 -17674 25967 -17640
rect 26205 -17674 26425 -17640
rect 26663 -17674 26883 -17640
rect 27121 -17674 27341 -17640
rect 27579 -17674 27799 -17640
rect 28037 -17674 28257 -17640
rect 28915 -17674 29135 -17640
rect 29373 -17674 29593 -17640
rect 29831 -17674 30051 -17640
rect 30289 -17674 30509 -17640
rect 30747 -17674 30967 -17640
rect 31205 -17674 31425 -17640
rect 31663 -17674 31883 -17640
rect 32121 -17674 32341 -17640
rect 32579 -17674 32799 -17640
rect 33037 -17674 33257 -17640
rect 23915 -19002 24135 -18968
rect 24373 -19002 24593 -18968
rect 24831 -19002 25051 -18968
rect 25289 -19002 25509 -18968
rect 25747 -19002 25967 -18968
rect 26205 -19002 26425 -18968
rect 26663 -19002 26883 -18968
rect 27121 -19002 27341 -18968
rect 27579 -19002 27799 -18968
rect 28037 -19002 28257 -18968
rect 28915 -19002 29135 -18968
rect 29373 -19002 29593 -18968
rect 29831 -19002 30051 -18968
rect 30289 -19002 30509 -18968
rect 30747 -19002 30967 -18968
rect 31205 -19002 31425 -18968
rect 31663 -19002 31883 -18968
rect 32121 -19002 32341 -18968
rect 32579 -19002 32799 -18968
rect 33037 -19002 33257 -18968
rect 8914 -20176 9134 -20142
rect 9372 -20176 9592 -20142
rect 9830 -20176 10050 -20142
rect 10288 -20176 10508 -20142
rect 10746 -20176 10966 -20142
rect 11204 -20176 11424 -20142
rect 11662 -20176 11882 -20142
rect 12120 -20176 12340 -20142
rect 12578 -20176 12798 -20142
rect 13036 -20176 13256 -20142
rect 13914 -20176 14134 -20142
rect 14372 -20176 14592 -20142
rect 14830 -20176 15050 -20142
rect 15288 -20176 15508 -20142
rect 15746 -20176 15966 -20142
rect 16204 -20176 16424 -20142
rect 16662 -20176 16882 -20142
rect 17120 -20176 17340 -20142
rect 17578 -20176 17798 -20142
rect 18036 -20176 18256 -20142
rect 8914 -20486 9134 -20452
rect 9372 -20486 9592 -20452
rect 9830 -20486 10050 -20452
rect 10288 -20486 10508 -20452
rect 10746 -20486 10966 -20452
rect 11204 -20486 11424 -20452
rect 11662 -20486 11882 -20452
rect 12120 -20486 12340 -20452
rect 12578 -20486 12798 -20452
rect 13036 -20486 13256 -20452
rect 13914 -20486 14134 -20452
rect 14372 -20486 14592 -20452
rect 14830 -20486 15050 -20452
rect 15288 -20486 15508 -20452
rect 15746 -20486 15966 -20452
rect 16204 -20486 16424 -20452
rect 16662 -20486 16882 -20452
rect 17120 -20486 17340 -20452
rect 17578 -20486 17798 -20452
rect 18036 -20486 18256 -20452
rect 8914 -20844 9134 -20810
rect 9372 -20844 9592 -20810
rect 9830 -20844 10050 -20810
rect 10288 -20844 10508 -20810
rect 10746 -20844 10966 -20810
rect 11204 -20844 11424 -20810
rect 11662 -20844 11882 -20810
rect 12120 -20844 12340 -20810
rect 12578 -20844 12798 -20810
rect 13036 -20844 13256 -20810
rect 8914 -21154 9134 -21120
rect 9372 -21154 9592 -21120
rect 9830 -21154 10050 -21120
rect 10288 -21154 10508 -21120
rect 10746 -21154 10966 -21120
rect 11204 -21154 11424 -21120
rect 11662 -21154 11882 -21120
rect 12120 -21154 12340 -21120
rect 12578 -21154 12798 -21120
rect 13036 -21154 13256 -21120
rect 23914 -20176 24134 -20142
rect 24372 -20176 24592 -20142
rect 24830 -20176 25050 -20142
rect 25288 -20176 25508 -20142
rect 25746 -20176 25966 -20142
rect 26204 -20176 26424 -20142
rect 26662 -20176 26882 -20142
rect 27120 -20176 27340 -20142
rect 27578 -20176 27798 -20142
rect 28036 -20176 28256 -20142
rect 28914 -20176 29134 -20142
rect 29372 -20176 29592 -20142
rect 29830 -20176 30050 -20142
rect 30288 -20176 30508 -20142
rect 30746 -20176 30966 -20142
rect 31204 -20176 31424 -20142
rect 31662 -20176 31882 -20142
rect 32120 -20176 32340 -20142
rect 32578 -20176 32798 -20142
rect 33036 -20176 33256 -20142
rect 23914 -20486 24134 -20452
rect 24372 -20486 24592 -20452
rect 24830 -20486 25050 -20452
rect 25288 -20486 25508 -20452
rect 25746 -20486 25966 -20452
rect 26204 -20486 26424 -20452
rect 26662 -20486 26882 -20452
rect 27120 -20486 27340 -20452
rect 27578 -20486 27798 -20452
rect 28036 -20486 28256 -20452
rect 28914 -20486 29134 -20452
rect 29372 -20486 29592 -20452
rect 29830 -20486 30050 -20452
rect 30288 -20486 30508 -20452
rect 30746 -20486 30966 -20452
rect 31204 -20486 31424 -20452
rect 31662 -20486 31882 -20452
rect 32120 -20486 32340 -20452
rect 32578 -20486 32798 -20452
rect 33036 -20486 33256 -20452
rect 23914 -20844 24134 -20810
rect 24372 -20844 24592 -20810
rect 24830 -20844 25050 -20810
rect 25288 -20844 25508 -20810
rect 25746 -20844 25966 -20810
rect 26204 -20844 26424 -20810
rect 26662 -20844 26882 -20810
rect 27120 -20844 27340 -20810
rect 27578 -20844 27798 -20810
rect 28036 -20844 28256 -20810
rect 23914 -21154 24134 -21120
rect 24372 -21154 24592 -21120
rect 24830 -21154 25050 -21120
rect 25288 -21154 25508 -21120
rect 25746 -21154 25966 -21120
rect 26204 -21154 26424 -21120
rect 26662 -21154 26882 -21120
rect 27120 -21154 27340 -21120
rect 27578 -21154 27798 -21120
rect 28036 -21154 28256 -21120
<< locali >>
rect 23334 17338 23434 17500
rect 32678 17338 32778 17500
rect 24014 16481 24030 16515
rect 24414 16481 24430 16515
rect 24872 16481 24888 16515
rect 25272 16481 25288 16515
rect 25730 16481 25746 16515
rect 26130 16481 26146 16515
rect 26588 16481 26604 16515
rect 26988 16481 27004 16515
rect 27446 16481 27462 16515
rect 27846 16481 27862 16515
rect 28304 16481 28320 16515
rect 28704 16481 28720 16515
rect 29162 16481 29178 16515
rect 29562 16481 29578 16515
rect 30020 16481 30036 16515
rect 30420 16481 30436 16515
rect 30878 16481 30894 16515
rect 31278 16481 31294 16515
rect 31736 16481 31752 16515
rect 32136 16481 32152 16515
rect 23776 16422 23810 16438
rect 23776 16230 23810 16246
rect 24634 16422 24668 16438
rect 24634 16230 24668 16246
rect 25492 16422 25526 16438
rect 25492 16230 25526 16246
rect 26350 16422 26384 16438
rect 26350 16230 26384 16246
rect 27208 16422 27242 16438
rect 27208 16230 27242 16246
rect 28066 16422 28100 16438
rect 28066 16230 28100 16246
rect 28924 16422 28958 16438
rect 28924 16230 28958 16246
rect 29782 16422 29816 16438
rect 29782 16230 29816 16246
rect 30640 16422 30674 16438
rect 30640 16230 30674 16246
rect 31498 16422 31532 16438
rect 31498 16230 31532 16246
rect 32356 16422 32390 16438
rect 32356 16230 32390 16246
rect 24014 16153 24030 16187
rect 24414 16153 24430 16187
rect 24872 16153 24888 16187
rect 25272 16153 25288 16187
rect 25730 16153 25746 16187
rect 26130 16153 26146 16187
rect 26588 16153 26604 16187
rect 26988 16153 27004 16187
rect 27446 16153 27462 16187
rect 27846 16153 27862 16187
rect 28304 16153 28320 16187
rect 28704 16153 28720 16187
rect 29162 16153 29178 16187
rect 29562 16153 29578 16187
rect 30020 16153 30036 16187
rect 30420 16153 30436 16187
rect 30878 16153 30894 16187
rect 31278 16153 31294 16187
rect 31736 16153 31752 16187
rect 32136 16153 32152 16187
rect 24014 15881 24030 15915
rect 24414 15881 24430 15915
rect 24872 15881 24888 15915
rect 25272 15881 25288 15915
rect 25730 15881 25746 15915
rect 26130 15881 26146 15915
rect 26588 15881 26604 15915
rect 26988 15881 27004 15915
rect 27446 15881 27462 15915
rect 27846 15881 27862 15915
rect 28304 15881 28320 15915
rect 28704 15881 28720 15915
rect 29162 15881 29178 15915
rect 29562 15881 29578 15915
rect 30020 15881 30036 15915
rect 30420 15881 30436 15915
rect 30878 15881 30894 15915
rect 31278 15881 31294 15915
rect 31736 15881 31752 15915
rect 32136 15881 32152 15915
rect 23776 15822 23810 15838
rect 23776 15630 23810 15646
rect 24634 15822 24668 15838
rect 24634 15630 24668 15646
rect 25492 15822 25526 15838
rect 25492 15630 25526 15646
rect 26350 15822 26384 15838
rect 26350 15630 26384 15646
rect 27208 15822 27242 15838
rect 27208 15630 27242 15646
rect 28066 15822 28100 15838
rect 28066 15630 28100 15646
rect 28924 15822 28958 15838
rect 28924 15630 28958 15646
rect 29782 15822 29816 15838
rect 29782 15630 29816 15646
rect 30640 15822 30674 15838
rect 30640 15630 30674 15646
rect 31498 15822 31532 15838
rect 31498 15630 31532 15646
rect 32356 15822 32390 15838
rect 32356 15630 32390 15646
rect 24014 15553 24030 15587
rect 24414 15553 24430 15587
rect 24872 15553 24888 15587
rect 25272 15553 25288 15587
rect 25730 15553 25746 15587
rect 26130 15553 26146 15587
rect 26588 15553 26604 15587
rect 26988 15553 27004 15587
rect 27446 15553 27462 15587
rect 27846 15553 27862 15587
rect 28304 15553 28320 15587
rect 28704 15553 28720 15587
rect 29162 15553 29178 15587
rect 29562 15553 29578 15587
rect 30020 15553 30036 15587
rect 30420 15553 30436 15587
rect 30878 15553 30894 15587
rect 31278 15553 31294 15587
rect 31736 15553 31752 15587
rect 32136 15553 32152 15587
rect 23334 15196 23434 15358
rect 32678 15196 32778 15358
rect 24049 14943 24145 14977
rect 24989 14943 25085 14977
rect 24049 14882 24083 14943
rect 25051 14882 25085 14943
rect 25171 14943 25267 14977
rect 26885 14943 26981 14977
rect 25171 14882 25205 14943
rect 26947 14884 26981 14943
rect 24243 14841 24259 14875
rect 24359 14841 24375 14875
rect 24501 14841 24517 14875
rect 24617 14841 24633 14875
rect 24759 14841 24775 14875
rect 24875 14841 24891 14875
rect 24163 14782 24197 14798
rect 24163 14390 24197 14406
rect 24421 14782 24455 14798
rect 24421 14390 24455 14406
rect 24679 14782 24713 14798
rect 24679 14390 24713 14406
rect 24937 14782 24971 14798
rect 24937 14390 24971 14406
rect 24243 14313 24259 14347
rect 24359 14313 24375 14347
rect 24501 14313 24517 14347
rect 24617 14313 24633 14347
rect 24759 14313 24775 14347
rect 24875 14313 24891 14347
rect 26947 14881 26948 14884
rect 25365 14841 25381 14875
rect 25481 14841 25497 14875
rect 25623 14841 25639 14875
rect 25739 14841 25755 14875
rect 25881 14841 25897 14875
rect 25997 14841 26013 14875
rect 26139 14841 26155 14875
rect 26255 14841 26271 14875
rect 26397 14841 26413 14875
rect 26513 14841 26529 14875
rect 26655 14841 26671 14875
rect 26771 14841 26787 14875
rect 25285 14782 25319 14798
rect 25285 14390 25319 14406
rect 25543 14782 25577 14798
rect 25543 14390 25577 14406
rect 25801 14782 25835 14798
rect 25801 14390 25835 14406
rect 26059 14782 26093 14798
rect 26059 14390 26093 14406
rect 26317 14782 26351 14798
rect 26317 14390 26351 14406
rect 26575 14782 26609 14798
rect 26575 14390 26609 14406
rect 26833 14782 26867 14798
rect 26833 14390 26867 14406
rect 25365 14313 25381 14347
rect 25481 14313 25497 14347
rect 25623 14313 25639 14347
rect 25739 14313 25755 14347
rect 25881 14313 25897 14347
rect 25997 14313 26013 14347
rect 26139 14313 26155 14347
rect 26255 14313 26271 14347
rect 26397 14313 26413 14347
rect 26513 14313 26529 14347
rect 26655 14313 26671 14347
rect 26771 14313 26787 14347
rect 27260 14441 27289 14475
rect 27323 14441 27381 14475
rect 27415 14441 27473 14475
rect 27507 14441 27565 14475
rect 27599 14441 27657 14475
rect 27691 14441 27749 14475
rect 27783 14441 27841 14475
rect 27875 14441 27933 14475
rect 27967 14441 28025 14475
rect 28059 14441 28117 14475
rect 28151 14441 28209 14475
rect 28243 14441 28301 14475
rect 28335 14441 28393 14475
rect 28427 14441 28485 14475
rect 28519 14441 28577 14475
rect 28611 14441 28669 14475
rect 28703 14441 28761 14475
rect 28795 14441 28853 14475
rect 28887 14441 28945 14475
rect 28979 14441 29037 14475
rect 29071 14441 29129 14475
rect 29163 14441 29221 14475
rect 29255 14441 29313 14475
rect 29347 14441 29405 14475
rect 29439 14441 29497 14475
rect 29531 14441 29589 14475
rect 29623 14441 29681 14475
rect 29715 14441 29773 14475
rect 29807 14441 29865 14475
rect 29899 14441 29957 14475
rect 29991 14441 30049 14475
rect 30083 14441 30141 14475
rect 30175 14441 30233 14475
rect 30267 14441 30325 14475
rect 30359 14441 30417 14475
rect 30451 14441 30509 14475
rect 30543 14441 30601 14475
rect 30635 14441 30693 14475
rect 30727 14441 30785 14475
rect 30819 14441 30877 14475
rect 30911 14441 30969 14475
rect 31003 14441 31061 14475
rect 31095 14441 31153 14475
rect 31187 14441 31245 14475
rect 31279 14441 31337 14475
rect 31371 14441 31429 14475
rect 31463 14441 31521 14475
rect 31555 14441 31613 14475
rect 31647 14441 31705 14475
rect 31739 14441 31797 14475
rect 31831 14441 31889 14475
rect 31923 14441 31981 14475
rect 32015 14441 32073 14475
rect 32107 14441 32165 14475
rect 32199 14441 32257 14475
rect 32291 14441 32320 14475
rect 27278 14391 27329 14407
rect 27278 14357 27295 14391
rect 27278 14323 27329 14357
rect 27363 14375 27429 14441
rect 27363 14341 27379 14375
rect 27413 14341 27429 14375
rect 27463 14391 27497 14407
rect 24049 14245 24083 14307
rect 25051 14245 25085 14307
rect 24049 14211 24145 14245
rect 24989 14211 25085 14245
rect 25171 14245 25205 14307
rect 26947 14245 26981 14307
rect 27278 14289 27295 14323
rect 27463 14323 27497 14357
rect 27329 14289 27428 14307
rect 27278 14273 27428 14289
rect 25171 14211 25267 14245
rect 26885 14211 26981 14245
rect 27278 14190 27348 14239
rect 27322 14163 27348 14190
rect 27278 14129 27292 14142
rect 27326 14129 27348 14163
rect 27278 14109 27348 14129
rect 27382 14178 27428 14273
rect 27382 14169 27394 14178
rect 27416 14135 27428 14144
rect 24049 14047 24145 14081
rect 24989 14047 25085 14081
rect 24049 13986 24083 14047
rect 24082 13985 24083 13986
rect 25051 13985 25085 14047
rect 25171 14047 25267 14081
rect 26885 14047 26981 14081
rect 27382 14075 27428 14135
rect 25171 13985 25205 14047
rect 26947 13986 26981 14047
rect 24243 13945 24259 13979
rect 24359 13945 24375 13979
rect 24501 13945 24517 13979
rect 24617 13945 24633 13979
rect 24759 13945 24775 13979
rect 24875 13945 24891 13979
rect 24163 13895 24197 13911
rect 24163 13703 24197 13719
rect 24421 13895 24455 13911
rect 24421 13703 24455 13719
rect 24679 13895 24713 13911
rect 24679 13703 24713 13719
rect 24937 13895 24971 13911
rect 24937 13703 24971 13719
rect 24243 13635 24259 13669
rect 24359 13635 24375 13669
rect 24501 13635 24517 13669
rect 24617 13635 24633 13669
rect 24759 13635 24775 13669
rect 24875 13635 24891 13669
rect 26980 13985 26981 13986
rect 25365 13945 25381 13979
rect 25481 13945 25497 13979
rect 25623 13945 25639 13979
rect 25739 13945 25755 13979
rect 25881 13945 25897 13979
rect 25997 13945 26013 13979
rect 26139 13945 26155 13979
rect 26255 13945 26271 13979
rect 26397 13945 26413 13979
rect 26513 13945 26529 13979
rect 26655 13945 26671 13979
rect 26771 13945 26787 13979
rect 25285 13895 25319 13911
rect 25285 13703 25319 13719
rect 25543 13895 25577 13911
rect 25543 13703 25577 13719
rect 25801 13895 25835 13911
rect 25801 13703 25835 13719
rect 26059 13895 26093 13911
rect 26059 13703 26093 13719
rect 26317 13895 26351 13911
rect 26317 13703 26351 13719
rect 26575 13895 26609 13911
rect 26575 13703 26609 13719
rect 26833 13895 26867 13911
rect 26833 13703 26867 13719
rect 25365 13635 25381 13669
rect 25481 13635 25497 13669
rect 25623 13635 25639 13669
rect 25739 13635 25755 13669
rect 25881 13635 25897 13669
rect 25997 13635 26013 13669
rect 26139 13635 26155 13669
rect 26255 13635 26271 13669
rect 26397 13635 26413 13669
rect 26513 13635 26529 13669
rect 26655 13635 26671 13669
rect 26771 13635 26787 13669
rect 27278 14041 27428 14075
rect 27278 14033 27329 14041
rect 27278 13999 27295 14033
rect 27463 14033 27497 14271
rect 27531 14388 27596 14404
rect 27531 14348 27542 14388
rect 27582 14348 27596 14388
rect 27630 14399 27680 14441
rect 27630 14365 27646 14399
rect 27630 14349 27680 14365
rect 27714 14391 27764 14407
rect 27714 14357 27730 14391
rect 27531 14247 27596 14348
rect 27714 14341 27764 14357
rect 27807 14397 27943 14407
rect 27807 14363 27823 14397
rect 27857 14363 27943 14397
rect 28058 14389 28124 14441
rect 28251 14399 28325 14441
rect 27807 14341 27943 14363
rect 27714 14315 27748 14341
rect 27669 14281 27748 14315
rect 27782 14305 27875 14307
rect 27543 14224 27635 14247
rect 27543 14190 27601 14224
rect 27543 14037 27635 14190
rect 27278 13983 27329 13999
rect 27363 13973 27379 14007
rect 27413 13973 27429 14007
rect 27669 14009 27703 14281
rect 27782 14279 27841 14305
rect 27816 14271 27841 14279
rect 27816 14245 27875 14271
rect 27782 14229 27875 14245
rect 27737 14169 27807 14191
rect 27737 14135 27749 14169
rect 27783 14135 27807 14169
rect 27737 14117 27807 14135
rect 27737 14083 27760 14117
rect 27794 14083 27807 14117
rect 27737 14067 27807 14083
rect 27841 14111 27875 14229
rect 27909 14185 27943 14341
rect 27977 14373 28011 14389
rect 28058 14355 28074 14389
rect 28108 14355 28124 14389
rect 28158 14373 28192 14389
rect 27977 14321 28011 14339
rect 28251 14365 28271 14399
rect 28305 14365 28325 14399
rect 28251 14349 28325 14365
rect 28359 14391 28393 14407
rect 28158 14321 28192 14339
rect 27977 14287 28192 14321
rect 28359 14315 28393 14357
rect 28440 14398 28614 14407
rect 28440 14364 28456 14398
rect 28490 14364 28614 14398
rect 28440 14339 28614 14364
rect 28648 14399 28698 14441
rect 28682 14365 28698 14399
rect 28802 14399 28946 14441
rect 28648 14349 28698 14365
rect 28732 14373 28766 14389
rect 28281 14281 28393 14315
rect 28281 14253 28315 14281
rect 28015 14219 28031 14253
rect 28065 14219 28315 14253
rect 28454 14271 28465 14305
rect 28499 14279 28546 14305
rect 28454 14247 28496 14271
rect 27909 14165 28247 14185
rect 27909 14151 28213 14165
rect 27841 14077 27862 14111
rect 27896 14077 27912 14111
rect 27841 14067 27912 14077
rect 27946 14009 27980 14151
rect 28021 14101 28117 14117
rect 28055 14067 28093 14101
rect 28151 14083 28179 14117
rect 28213 14115 28247 14131
rect 28127 14067 28179 14083
rect 28281 14081 28315 14219
rect 27463 13983 27497 13999
rect 27363 13931 27429 13973
rect 27569 13969 27585 14003
rect 27619 13969 27635 14003
rect 27669 13975 27718 14009
rect 27752 13975 27768 14009
rect 27809 13975 27825 14009
rect 27859 13975 27980 14009
rect 28155 14007 28221 14023
rect 27569 13931 27635 13969
rect 28155 13973 28171 14007
rect 28205 13973 28221 14007
rect 28155 13931 28221 13973
rect 28263 14003 28315 14081
rect 28353 14245 28496 14247
rect 28530 14245 28546 14279
rect 28580 14263 28614 14339
rect 28802 14365 28818 14399
rect 28852 14365 28896 14399
rect 28930 14365 28946 14399
rect 28980 14391 29061 14407
rect 29212 14399 29246 14441
rect 28732 14331 28766 14339
rect 29014 14357 29061 14391
rect 28732 14297 28892 14331
rect 28353 14213 28488 14245
rect 28580 14229 28774 14263
rect 28808 14229 28824 14263
rect 28353 14105 28395 14213
rect 28580 14211 28614 14229
rect 28353 14071 28361 14105
rect 28353 14055 28395 14071
rect 28429 14169 28499 14179
rect 28429 14153 28465 14169
rect 28429 14119 28457 14153
rect 28491 14119 28499 14135
rect 28429 14055 28499 14119
rect 28533 14177 28614 14211
rect 28533 14021 28567 14177
rect 28681 14164 28789 14195
rect 28858 14179 28892 14297
rect 28980 14323 29061 14357
rect 29014 14289 29061 14323
rect 28980 14255 29061 14289
rect 29014 14221 29061 14255
rect 28980 14205 29061 14221
rect 28858 14173 28947 14179
rect 28715 14155 28789 14164
rect 28601 14127 28645 14143
rect 28635 14093 28645 14127
rect 28681 14121 28697 14130
rect 28731 14121 28789 14155
rect 28601 14087 28645 14093
rect 28741 14101 28789 14121
rect 28601 14053 28707 14087
rect 28377 14007 28567 14021
rect 28263 13969 28283 14003
rect 28317 13969 28333 14003
rect 28377 13973 28393 14007
rect 28427 13973 28567 14007
rect 28377 13965 28567 13973
rect 28601 14003 28639 14019
rect 28601 13969 28605 14003
rect 28673 14007 28707 14053
rect 28775 14067 28789 14101
rect 28741 14041 28789 14067
rect 28823 14163 28947 14173
rect 28823 14129 28897 14163
rect 28931 14129 28947 14163
rect 28823 14113 28947 14129
rect 28995 14170 29061 14205
rect 28995 14122 29004 14170
rect 29052 14122 29061 14170
rect 28823 14078 28888 14113
rect 28995 14079 29061 14122
rect 28823 14023 28887 14078
rect 28673 13989 28823 14007
rect 28857 13989 28887 14023
rect 28673 13973 28887 13989
rect 28927 14046 28961 14068
rect 28601 13931 28639 13969
rect 28927 13931 28961 14012
rect 28995 14045 29011 14079
rect 29045 14045 29061 14079
rect 28995 14011 29061 14045
rect 28995 13977 29011 14011
rect 29045 13977 29061 14011
rect 29099 14365 29115 14399
rect 29149 14365 29165 14399
rect 29099 14331 29165 14365
rect 29099 14297 29115 14331
rect 29149 14297 29165 14331
rect 29099 14179 29165 14297
rect 29444 14399 29486 14441
rect 29212 14331 29246 14365
rect 29212 14263 29246 14297
rect 29212 14213 29246 14229
rect 29296 14363 29347 14379
rect 29330 14329 29347 14363
rect 29296 14295 29347 14329
rect 29330 14261 29347 14295
rect 29296 14203 29347 14261
rect 29444 14365 29452 14399
rect 29444 14331 29486 14365
rect 29444 14297 29452 14331
rect 29444 14263 29486 14297
rect 29444 14229 29452 14263
rect 29444 14213 29486 14229
rect 29520 14399 29586 14407
rect 29520 14365 29536 14399
rect 29570 14365 29586 14399
rect 29520 14331 29586 14365
rect 29520 14297 29536 14331
rect 29570 14297 29586 14331
rect 29520 14263 29586 14297
rect 29520 14229 29536 14263
rect 29570 14229 29586 14263
rect 29520 14211 29586 14229
rect 29669 14399 29725 14441
rect 29669 14365 29691 14399
rect 29669 14331 29725 14365
rect 29669 14297 29691 14331
rect 29669 14263 29725 14297
rect 29669 14229 29691 14263
rect 29669 14213 29725 14229
rect 29759 14399 29825 14407
rect 29759 14365 29775 14399
rect 29809 14365 29825 14399
rect 29759 14331 29825 14365
rect 29759 14297 29775 14331
rect 29809 14297 29825 14331
rect 29759 14268 29825 14297
rect 29759 14226 29764 14268
rect 29812 14226 29825 14268
rect 29759 14211 29825 14226
rect 29859 14399 29911 14441
rect 29893 14365 29911 14399
rect 29859 14331 29911 14365
rect 29893 14297 29911 14331
rect 29859 14263 29911 14297
rect 29893 14229 29911 14263
rect 29859 14213 29911 14229
rect 29994 14399 30060 14407
rect 29994 14368 30010 14399
rect 30044 14368 30060 14399
rect 29994 14320 30000 14368
rect 30048 14320 30060 14368
rect 29994 14297 30010 14320
rect 30044 14297 30060 14320
rect 29994 14263 30060 14297
rect 29994 14229 30010 14263
rect 30044 14229 30060 14263
rect 29994 14211 30060 14229
rect 30094 14399 30136 14441
rect 30128 14365 30136 14399
rect 30334 14399 30368 14441
rect 30094 14331 30136 14365
rect 30128 14297 30136 14331
rect 30094 14263 30136 14297
rect 30128 14229 30136 14263
rect 30094 14213 30136 14229
rect 30233 14363 30284 14379
rect 30233 14329 30250 14363
rect 30233 14295 30284 14329
rect 30233 14261 30250 14295
rect 29099 14163 29271 14179
rect 29099 14129 29237 14163
rect 29099 14113 29271 14129
rect 29099 14033 29149 14113
rect 29305 14073 29347 14203
rect 29440 14170 29506 14177
rect 29440 14130 29444 14170
rect 29492 14130 29506 14170
rect 29440 14129 29456 14130
rect 29490 14129 29506 14130
rect 29296 14057 29347 14073
rect 29099 13999 29115 14033
rect 29099 13983 29149 13999
rect 29212 14027 29246 14050
rect 28995 13969 29061 13977
rect 29212 13931 29246 13993
rect 29330 14023 29347 14057
rect 29296 13967 29347 14023
rect 29440 14079 29486 14095
rect 29540 14091 29586 14211
rect 29671 14170 29738 14179
rect 29671 14128 29682 14170
rect 29730 14128 29738 14170
rect 29671 14125 29738 14128
rect 29772 14091 29806 14211
rect 29840 14170 29907 14179
rect 29840 14129 29856 14170
rect 29904 14129 29907 14170
rect 29994 14091 30040 14211
rect 30233 14203 30284 14261
rect 30334 14331 30368 14365
rect 30334 14263 30368 14297
rect 30334 14213 30368 14229
rect 30415 14365 30431 14399
rect 30465 14365 30481 14399
rect 30415 14331 30481 14365
rect 30415 14297 30431 14331
rect 30465 14297 30481 14331
rect 30074 14170 30140 14177
rect 30074 14129 30090 14170
rect 30138 14130 30140 14170
rect 30124 14129 30140 14130
rect 29440 14045 29452 14079
rect 29440 14011 29486 14045
rect 29440 13977 29452 14011
rect 29440 13931 29486 13977
rect 29520 14079 29586 14091
rect 29520 14058 29536 14079
rect 29570 14058 29586 14079
rect 29520 14010 29532 14058
rect 29580 14010 29586 14058
rect 29520 13977 29536 14010
rect 29570 13977 29586 14010
rect 29520 13965 29586 13977
rect 29669 14075 29731 14091
rect 29669 14041 29691 14075
rect 29725 14041 29731 14075
rect 29669 14007 29731 14041
rect 29669 13973 29691 14007
rect 29725 13973 29731 14007
rect 29669 13931 29731 13973
rect 29772 14075 29911 14091
rect 29772 14041 29859 14075
rect 29893 14041 29911 14075
rect 29772 14007 29911 14041
rect 29772 13973 29859 14007
rect 29893 13973 29911 14007
rect 29772 13965 29911 13973
rect 29994 14079 30060 14091
rect 29994 14045 30010 14079
rect 30044 14045 30060 14079
rect 29994 14011 30060 14045
rect 29994 13977 30010 14011
rect 30044 13977 30060 14011
rect 29994 13965 30060 13977
rect 30094 14079 30140 14095
rect 30128 14045 30140 14079
rect 30094 14011 30140 14045
rect 30128 13977 30140 14011
rect 30094 13931 30140 13977
rect 30233 14073 30275 14203
rect 30415 14179 30481 14297
rect 30309 14163 30481 14179
rect 30343 14129 30481 14163
rect 30309 14113 30481 14129
rect 30233 14057 30284 14073
rect 30233 14023 30250 14057
rect 30233 13967 30284 14023
rect 30334 14027 30368 14050
rect 30334 13931 30368 13993
rect 30431 14033 30481 14113
rect 30465 13999 30481 14033
rect 30431 13983 30481 13999
rect 30519 14391 30600 14407
rect 30519 14357 30566 14391
rect 30634 14399 30778 14441
rect 30634 14365 30650 14399
rect 30684 14365 30728 14399
rect 30762 14365 30778 14399
rect 30882 14399 30932 14441
rect 30814 14373 30848 14389
rect 30519 14323 30600 14357
rect 30882 14365 30898 14399
rect 30882 14349 30932 14365
rect 30966 14398 31140 14407
rect 30966 14364 31090 14398
rect 31124 14364 31140 14398
rect 30814 14331 30848 14339
rect 30519 14289 30566 14323
rect 30519 14255 30600 14289
rect 30519 14221 30566 14255
rect 30519 14205 30600 14221
rect 30688 14297 30848 14331
rect 30966 14339 31140 14364
rect 31187 14391 31221 14407
rect 30519 14170 30585 14205
rect 30688 14179 30722 14297
rect 30966 14263 31000 14339
rect 31187 14315 31221 14357
rect 31255 14399 31329 14441
rect 31255 14365 31275 14399
rect 31309 14365 31329 14399
rect 31456 14389 31522 14441
rect 31637 14397 31773 14407
rect 31255 14349 31329 14365
rect 31388 14373 31422 14389
rect 31456 14355 31472 14389
rect 31506 14355 31522 14389
rect 31569 14373 31603 14389
rect 31388 14321 31422 14339
rect 31569 14321 31603 14339
rect 30756 14229 30772 14263
rect 30806 14229 31000 14263
rect 31034 14279 31081 14305
rect 31034 14245 31050 14279
rect 31115 14271 31126 14305
rect 31187 14281 31299 14315
rect 31388 14287 31603 14321
rect 31637 14363 31723 14397
rect 31757 14363 31773 14397
rect 31637 14341 31773 14363
rect 31816 14391 31866 14407
rect 31850 14357 31866 14391
rect 31816 14341 31866 14357
rect 31900 14399 31950 14441
rect 31934 14365 31950 14399
rect 31900 14349 31950 14365
rect 31984 14396 32049 14404
rect 31984 14356 31992 14396
rect 32038 14356 32049 14396
rect 31084 14247 31126 14271
rect 31265 14253 31299 14281
rect 31084 14245 31227 14247
rect 30966 14211 31000 14229
rect 31092 14213 31227 14245
rect 30519 14122 30528 14170
rect 30576 14122 30585 14170
rect 30519 14079 30585 14122
rect 30633 14173 30722 14179
rect 30633 14163 30757 14173
rect 30633 14129 30649 14163
rect 30683 14129 30757 14163
rect 30633 14113 30757 14129
rect 30519 14045 30535 14079
rect 30569 14045 30585 14079
rect 30692 14078 30757 14113
rect 30519 14011 30585 14045
rect 30519 13977 30535 14011
rect 30569 13977 30585 14011
rect 30519 13969 30585 13977
rect 30619 14046 30653 14068
rect 30619 13931 30653 14012
rect 30693 14023 30757 14078
rect 30791 14164 30899 14195
rect 30966 14177 31047 14211
rect 30791 14155 30865 14164
rect 30791 14121 30849 14155
rect 30883 14121 30899 14130
rect 30935 14127 30979 14143
rect 30791 14101 30839 14121
rect 30791 14067 30805 14101
rect 30935 14093 30945 14127
rect 30935 14087 30979 14093
rect 30791 14041 30839 14067
rect 30873 14053 30979 14087
rect 30693 13989 30723 14023
rect 30873 14007 30907 14053
rect 31013 14021 31047 14177
rect 31081 14169 31151 14179
rect 31115 14153 31151 14169
rect 31081 14119 31089 14135
rect 31123 14119 31151 14153
rect 31081 14055 31151 14119
rect 31185 14105 31227 14213
rect 31219 14071 31227 14105
rect 31185 14055 31227 14071
rect 31265 14219 31515 14253
rect 31549 14219 31565 14253
rect 31265 14081 31299 14219
rect 31637 14185 31671 14341
rect 31832 14315 31866 14341
rect 31333 14165 31671 14185
rect 31367 14151 31671 14165
rect 31705 14305 31798 14307
rect 31739 14279 31798 14305
rect 31832 14281 31911 14315
rect 31739 14271 31764 14279
rect 31705 14245 31764 14271
rect 31705 14229 31798 14245
rect 31333 14115 31367 14131
rect 31401 14083 31429 14117
rect 31463 14101 31559 14117
rect 30757 13989 30907 14007
rect 30693 13973 30907 13989
rect 30941 14003 30979 14019
rect 30975 13969 30979 14003
rect 30941 13931 30979 13969
rect 31013 14007 31203 14021
rect 31013 13973 31153 14007
rect 31187 13973 31203 14007
rect 31265 14003 31317 14081
rect 31401 14067 31453 14083
rect 31487 14067 31525 14101
rect 31013 13965 31203 13973
rect 31247 13969 31263 14003
rect 31297 13969 31317 14003
rect 31359 14007 31425 14023
rect 31359 13973 31375 14007
rect 31409 13973 31425 14007
rect 31600 14009 31634 14151
rect 31705 14111 31739 14229
rect 31668 14077 31684 14111
rect 31718 14077 31739 14111
rect 31668 14067 31739 14077
rect 31773 14169 31843 14191
rect 31773 14135 31797 14169
rect 31831 14135 31843 14169
rect 31773 14117 31843 14135
rect 31773 14083 31786 14117
rect 31820 14083 31843 14117
rect 31773 14067 31843 14083
rect 31877 14009 31911 14281
rect 31984 14247 32049 14356
rect 32083 14391 32117 14407
rect 32083 14323 32117 14357
rect 32151 14375 32217 14441
rect 32151 14341 32167 14375
rect 32201 14341 32217 14375
rect 32251 14391 32302 14407
rect 32285 14357 32302 14391
rect 32251 14323 32302 14357
rect 31945 14224 32037 14247
rect 31979 14190 32037 14224
rect 31945 14037 32037 14190
rect 31600 13975 31721 14009
rect 31755 13975 31771 14009
rect 31812 13975 31828 14009
rect 31862 13975 31911 14009
rect 32083 14033 32117 14271
rect 32152 14289 32251 14307
rect 32285 14289 32302 14323
rect 32152 14273 32302 14289
rect 32152 14178 32198 14273
rect 32186 14169 32198 14178
rect 32152 14135 32164 14144
rect 32152 14075 32198 14135
rect 32232 14172 32302 14239
rect 32232 14124 32252 14172
rect 32300 14124 32302 14172
rect 32232 14109 32302 14124
rect 32152 14041 32302 14075
rect 31359 13931 31425 13973
rect 31945 13969 31961 14003
rect 31995 13969 32011 14003
rect 32251 14033 32302 14041
rect 32083 13983 32117 13999
rect 31945 13931 32011 13969
rect 32151 13973 32167 14007
rect 32201 13973 32217 14007
rect 32285 13999 32302 14033
rect 32251 13983 32302 13999
rect 32151 13931 32217 13973
rect 27260 13897 27289 13931
rect 27323 13897 27381 13931
rect 27415 13897 27473 13931
rect 27507 13897 27565 13931
rect 27599 13897 27657 13931
rect 27691 13897 27749 13931
rect 27783 13897 27841 13931
rect 27875 13897 27933 13931
rect 27967 13897 28025 13931
rect 28059 13897 28117 13931
rect 28151 13897 28209 13931
rect 28243 13897 28301 13931
rect 28335 13897 28393 13931
rect 28427 13897 28485 13931
rect 28519 13897 28577 13931
rect 28611 13897 28669 13931
rect 28703 13897 28761 13931
rect 28795 13897 28853 13931
rect 28887 13897 28945 13931
rect 28979 13897 29037 13931
rect 29071 13897 29129 13931
rect 29163 13897 29221 13931
rect 29255 13897 29313 13931
rect 29347 13897 29405 13931
rect 29439 13897 29497 13931
rect 29531 13897 29589 13931
rect 29623 13897 29681 13931
rect 29715 13897 29773 13931
rect 29807 13897 29865 13931
rect 29899 13897 29957 13931
rect 29991 13897 30049 13931
rect 30083 13897 30141 13931
rect 30175 13897 30233 13931
rect 30267 13897 30325 13931
rect 30359 13897 30417 13931
rect 30451 13897 30509 13931
rect 30543 13897 30601 13931
rect 30635 13897 30693 13931
rect 30727 13897 30785 13931
rect 30819 13897 30877 13931
rect 30911 13897 30969 13931
rect 31003 13897 31061 13931
rect 31095 13897 31153 13931
rect 31187 13897 31245 13931
rect 31279 13897 31337 13931
rect 31371 13897 31429 13931
rect 31463 13897 31521 13931
rect 31555 13897 31613 13931
rect 31647 13897 31705 13931
rect 31739 13897 31797 13931
rect 31831 13897 31889 13931
rect 31923 13897 31981 13931
rect 32015 13897 32073 13931
rect 32107 13897 32165 13931
rect 32199 13897 32257 13931
rect 32291 13897 32320 13931
rect 24049 13567 24083 13629
rect 25051 13567 25085 13629
rect 24049 13533 24145 13567
rect 24989 13533 25085 13567
rect 25171 13567 25205 13629
rect 26947 13567 26981 13629
rect 25171 13533 25267 13567
rect 26885 13533 26981 13567
rect 23334 13158 23434 13320
rect 32678 13158 32778 13320
rect 24450 12892 24466 12926
rect 24926 12892 24942 12926
rect 25308 12892 25324 12926
rect 25784 12892 25800 12926
rect 26166 12892 26182 12926
rect 26642 12892 26658 12926
rect 27024 12892 27040 12926
rect 27500 12892 27516 12926
rect 27882 12892 27898 12926
rect 28358 12892 28374 12926
rect 28740 12892 28756 12926
rect 29216 12892 29232 12926
rect 29598 12892 29614 12926
rect 30074 12892 30090 12926
rect 30456 12892 30472 12926
rect 30932 12892 30948 12926
rect 31314 12892 31330 12926
rect 31790 12892 31806 12926
rect 24250 12842 24284 12858
rect 24250 12650 24284 12666
rect 25108 12842 25142 12858
rect 25108 12650 25142 12666
rect 25966 12842 26000 12858
rect 25966 12650 26000 12666
rect 26824 12842 26858 12858
rect 26824 12650 26858 12666
rect 27682 12842 27716 12858
rect 27682 12650 27716 12666
rect 28540 12842 28574 12858
rect 28540 12650 28574 12666
rect 29398 12842 29432 12858
rect 29398 12650 29432 12666
rect 30256 12842 30290 12858
rect 30256 12650 30290 12666
rect 31114 12842 31148 12858
rect 31114 12650 31148 12666
rect 31972 12842 32006 12858
rect 31972 12650 32006 12666
rect 24450 12582 24466 12616
rect 24926 12582 24942 12616
rect 25308 12582 25324 12616
rect 25784 12582 25800 12616
rect 26166 12582 26182 12616
rect 26642 12582 26658 12616
rect 27024 12582 27040 12616
rect 27500 12582 27516 12616
rect 27882 12582 27898 12616
rect 28358 12582 28374 12616
rect 28740 12582 28756 12616
rect 29216 12582 29232 12616
rect 29598 12582 29614 12616
rect 30074 12582 30090 12616
rect 30456 12582 30472 12616
rect 30932 12582 30948 12616
rect 31314 12582 31330 12616
rect 31790 12582 31806 12616
rect 24450 12310 24466 12344
rect 24926 12310 24942 12344
rect 25308 12310 25324 12344
rect 25784 12310 25800 12344
rect 26166 12310 26182 12344
rect 26642 12310 26658 12344
rect 27024 12310 27040 12344
rect 27500 12310 27516 12344
rect 27882 12310 27898 12344
rect 28358 12310 28374 12344
rect 28740 12310 28756 12344
rect 29216 12310 29232 12344
rect 29598 12310 29614 12344
rect 30074 12310 30090 12344
rect 30456 12310 30472 12344
rect 30932 12310 30948 12344
rect 31314 12310 31330 12344
rect 31790 12310 31806 12344
rect 24250 12260 24284 12276
rect 24250 12068 24284 12084
rect 25108 12260 25142 12276
rect 25108 12068 25142 12084
rect 25966 12260 26000 12276
rect 25966 12068 26000 12084
rect 26824 12260 26858 12276
rect 26824 12068 26858 12084
rect 27682 12260 27716 12276
rect 27682 12068 27716 12084
rect 28540 12260 28574 12276
rect 28540 12068 28574 12084
rect 29398 12260 29432 12276
rect 29398 12068 29432 12084
rect 30256 12260 30290 12276
rect 30256 12068 30290 12084
rect 31114 12260 31148 12276
rect 31114 12068 31148 12084
rect 31972 12260 32006 12276
rect 31972 12068 32006 12084
rect 24450 12000 24466 12034
rect 24926 12000 24942 12034
rect 25308 12000 25324 12034
rect 25784 12000 25800 12034
rect 26166 12000 26182 12034
rect 26642 12000 26658 12034
rect 27024 12000 27040 12034
rect 27500 12000 27516 12034
rect 27882 12000 27898 12034
rect 28358 12000 28374 12034
rect 28740 12000 28756 12034
rect 29216 12000 29232 12034
rect 29598 12000 29614 12034
rect 30074 12000 30090 12034
rect 30456 12000 30472 12034
rect 30932 12000 30948 12034
rect 31314 12000 31330 12034
rect 31790 12000 31806 12034
rect 23334 11056 23434 11218
rect 32678 11056 32778 11218
rect 12960 10572 13060 10734
rect 21884 10572 21984 10734
rect 15288 9706 15304 9740
rect 15524 9706 15540 9740
rect 15746 9706 15762 9740
rect 15982 9706 15998 9740
rect 16204 9706 16220 9740
rect 16440 9706 16456 9740
rect 16662 9706 16678 9740
rect 16898 9706 16914 9740
rect 17120 9706 17136 9740
rect 17356 9706 17372 9740
rect 17578 9706 17594 9740
rect 17814 9706 17830 9740
rect 18036 9706 18052 9740
rect 18272 9706 18288 9740
rect 18494 9706 18510 9740
rect 18730 9706 18746 9740
rect 18952 9706 18968 9740
rect 19188 9706 19204 9740
rect 19410 9706 19426 9740
rect 19646 9706 19662 9740
rect 15168 9656 15202 9672
rect 15168 9464 15202 9480
rect 15626 9656 15660 9672
rect 15626 9464 15660 9480
rect 16084 9656 16118 9672
rect 16084 9464 16118 9480
rect 16542 9656 16576 9672
rect 16542 9464 16576 9480
rect 17000 9656 17034 9672
rect 17000 9464 17034 9480
rect 17458 9656 17492 9672
rect 17458 9464 17492 9480
rect 17916 9656 17950 9672
rect 17916 9464 17950 9480
rect 18374 9656 18408 9672
rect 18374 9464 18408 9480
rect 18832 9656 18866 9672
rect 18832 9464 18866 9480
rect 19290 9656 19324 9672
rect 19290 9464 19324 9480
rect 19748 9656 19782 9672
rect 19748 9464 19782 9480
rect 15288 9396 15304 9430
rect 15524 9396 15540 9430
rect 15746 9396 15762 9430
rect 15982 9396 15998 9430
rect 16204 9396 16220 9430
rect 16440 9396 16456 9430
rect 16662 9396 16678 9430
rect 16898 9396 16914 9430
rect 17120 9396 17136 9430
rect 17356 9396 17372 9430
rect 17578 9396 17594 9430
rect 17814 9396 17830 9430
rect 18036 9396 18052 9430
rect 18272 9396 18288 9430
rect 18494 9396 18510 9430
rect 18730 9396 18746 9430
rect 18952 9396 18968 9430
rect 19188 9396 19204 9430
rect 19410 9396 19426 9430
rect 19646 9396 19662 9430
rect 12960 8934 13060 9096
rect 21884 8934 21984 9096
rect 23542 10572 23642 10734
rect 28886 10572 28986 10734
rect 24050 9706 24066 9740
rect 24286 9706 24302 9740
rect 24508 9706 24524 9740
rect 24744 9706 24760 9740
rect 24966 9706 24982 9740
rect 25202 9706 25218 9740
rect 25424 9706 25440 9740
rect 25660 9706 25676 9740
rect 25882 9706 25898 9740
rect 26118 9706 26134 9740
rect 26340 9706 26356 9740
rect 26576 9706 26592 9740
rect 26798 9706 26814 9740
rect 27034 9706 27050 9740
rect 27256 9706 27272 9740
rect 27492 9706 27508 9740
rect 27714 9706 27730 9740
rect 27950 9706 27966 9740
rect 28172 9706 28188 9740
rect 28408 9706 28424 9740
rect 23930 9656 23964 9672
rect 23930 9464 23964 9480
rect 24388 9656 24422 9672
rect 24388 9464 24422 9480
rect 24846 9656 24880 9672
rect 24846 9464 24880 9480
rect 25304 9656 25338 9672
rect 25304 9464 25338 9480
rect 25762 9656 25796 9672
rect 25762 9464 25796 9480
rect 26220 9656 26254 9672
rect 26220 9464 26254 9480
rect 26678 9656 26712 9672
rect 26678 9464 26712 9480
rect 27136 9656 27170 9672
rect 27136 9464 27170 9480
rect 27594 9656 27628 9672
rect 27594 9464 27628 9480
rect 28052 9656 28086 9672
rect 28052 9464 28086 9480
rect 28510 9656 28544 9672
rect 28510 9464 28544 9480
rect 24050 9396 24066 9430
rect 24286 9396 24302 9430
rect 24508 9396 24524 9430
rect 24744 9396 24760 9430
rect 24966 9396 24982 9430
rect 25202 9396 25218 9430
rect 25424 9396 25440 9430
rect 25660 9396 25676 9430
rect 25882 9396 25898 9430
rect 26118 9396 26134 9430
rect 26340 9396 26356 9430
rect 26576 9396 26592 9430
rect 26798 9396 26814 9430
rect 27034 9396 27050 9430
rect 27256 9396 27272 9430
rect 27492 9396 27508 9430
rect 27714 9396 27730 9430
rect 27950 9396 27966 9430
rect 28172 9396 28188 9430
rect 28408 9396 28424 9430
rect 23542 8854 23642 9016
rect 28886 8854 28986 9016
rect 30210 8943 30239 8977
rect 30273 8943 30302 8977
rect 30552 8943 30581 8977
rect 30615 8943 30673 8977
rect 30707 8943 30765 8977
rect 30799 8943 30857 8977
rect 30891 8943 30949 8977
rect 30983 8943 31041 8977
rect 31075 8943 31133 8977
rect 31167 8943 31225 8977
rect 31259 8943 31317 8977
rect 31351 8943 31409 8977
rect 31443 8943 31501 8977
rect 31535 8943 31593 8977
rect 31627 8943 31685 8977
rect 31719 8943 31777 8977
rect 31811 8943 31869 8977
rect 31903 8943 31961 8977
rect 31995 8943 32053 8977
rect 32087 8943 32145 8977
rect 32179 8943 32237 8977
rect 32271 8943 32329 8977
rect 32363 8943 32421 8977
rect 32455 8943 32513 8977
rect 32547 8943 32605 8977
rect 32639 8943 32697 8977
rect 32731 8943 32789 8977
rect 32823 8943 32881 8977
rect 32915 8943 32973 8977
rect 33007 8943 33036 8977
rect 33110 8943 33139 8977
rect 33173 8943 33202 8977
rect 35984 8943 36013 8977
rect 36047 8943 36076 8977
rect 29076 8897 29105 8931
rect 29139 8897 29197 8931
rect 29231 8897 29289 8931
rect 29323 8897 29381 8931
rect 29415 8897 29473 8931
rect 29507 8897 29565 8931
rect 29599 8897 29657 8931
rect 29691 8897 29749 8931
rect 29783 8897 29812 8931
rect 29140 8851 29186 8897
rect 29140 8817 29152 8851
rect 29140 8783 29186 8817
rect 29140 8749 29152 8783
rect 29140 8733 29186 8749
rect 29220 8851 29286 8863
rect 29220 8817 29236 8851
rect 29270 8817 29286 8851
rect 29220 8783 29286 8817
rect 29378 8855 29431 8897
rect 29378 8821 29397 8855
rect 29378 8805 29431 8821
rect 29465 8847 29531 8863
rect 29465 8813 29481 8847
rect 29515 8813 29531 8847
rect 29220 8749 29236 8783
rect 29270 8749 29286 8783
rect 29220 8737 29286 8749
rect 29240 8700 29286 8737
rect 29465 8769 29531 8813
rect 29565 8855 29599 8897
rect 29565 8805 29599 8821
rect 29633 8847 29699 8863
rect 29633 8813 29649 8847
rect 29683 8813 29699 8847
rect 29633 8769 29699 8813
rect 29733 8854 29783 8897
rect 29767 8820 29783 8854
rect 29733 8804 29783 8820
rect 30227 8872 30285 8943
rect 30227 8838 30239 8872
rect 30273 8838 30285 8872
rect 30227 8779 30285 8838
rect 29465 8733 29786 8769
rect 29733 8700 29786 8733
rect 30227 8745 30239 8779
rect 30273 8745 30285 8779
rect 30587 8893 30621 8909
rect 30587 8825 30621 8859
rect 30655 8877 30721 8943
rect 30655 8843 30671 8877
rect 30705 8843 30721 8877
rect 30755 8893 30792 8909
rect 30789 8859 30792 8893
rect 30755 8825 30792 8859
rect 30840 8901 30893 8943
rect 30840 8867 30859 8901
rect 30840 8851 30893 8867
rect 30927 8893 30977 8909
rect 30927 8859 30943 8893
rect 31274 8901 31308 8943
rect 30621 8807 30720 8809
rect 30621 8791 30678 8807
rect 30587 8775 30678 8791
rect 30227 8710 30285 8745
rect 30674 8773 30678 8775
rect 30712 8773 30720 8807
rect 29140 8698 29156 8699
rect 12960 8536 13060 8698
rect 21884 8536 21984 8698
rect 29190 8665 29206 8699
rect 29188 8651 29206 8665
rect 29240 8652 29246 8700
rect 29373 8652 29382 8699
rect 29430 8665 29481 8699
rect 29515 8665 29565 8699
rect 29599 8665 29649 8699
rect 29683 8665 29699 8699
rect 29430 8652 29699 8665
rect 13456 7864 13472 7898
rect 13692 7864 13708 7898
rect 13914 7864 13930 7898
rect 14150 7864 14166 7898
rect 14372 7864 14388 7898
rect 14608 7864 14624 7898
rect 14830 7864 14846 7898
rect 15066 7864 15082 7898
rect 15288 7864 15304 7898
rect 15524 7864 15540 7898
rect 15746 7864 15762 7898
rect 15982 7864 15998 7898
rect 16204 7864 16220 7898
rect 16440 7864 16456 7898
rect 16662 7864 16678 7898
rect 16898 7864 16914 7898
rect 17120 7864 17136 7898
rect 17356 7864 17372 7898
rect 17578 7864 17594 7898
rect 17814 7864 17830 7898
rect 18036 7864 18052 7898
rect 18272 7864 18288 7898
rect 18494 7864 18510 7898
rect 18730 7864 18746 7898
rect 18952 7864 18968 7898
rect 19188 7864 19204 7898
rect 19410 7864 19426 7898
rect 19646 7864 19662 7898
rect 19868 7864 19884 7898
rect 20104 7864 20120 7898
rect 20326 7864 20342 7898
rect 20562 7864 20578 7898
rect 20784 7864 20800 7898
rect 21020 7864 21036 7898
rect 21242 7864 21258 7898
rect 21478 7864 21494 7898
rect 13336 7805 13370 7821
rect 13336 6213 13370 6229
rect 13794 7805 13828 7821
rect 13794 6213 13828 6229
rect 14252 7805 14286 7821
rect 14252 6213 14286 6229
rect 14710 7805 14744 7821
rect 14710 6213 14744 6229
rect 15168 7805 15202 7821
rect 15168 6213 15202 6229
rect 15626 7805 15660 7821
rect 15626 6213 15660 6229
rect 16084 7805 16118 7821
rect 16084 6213 16118 6229
rect 16542 7805 16576 7821
rect 16542 6213 16576 6229
rect 17000 7805 17034 7821
rect 17000 6213 17034 6229
rect 17458 7805 17492 7821
rect 17458 6213 17492 6229
rect 17916 7805 17950 7821
rect 17916 6213 17950 6229
rect 18374 7805 18408 7821
rect 18374 6213 18408 6229
rect 18832 7805 18866 7821
rect 18832 6213 18866 6229
rect 19290 7805 19324 7821
rect 19290 6213 19324 6229
rect 19748 7805 19782 7821
rect 19748 6213 19782 6229
rect 20206 7805 20240 7821
rect 20206 6213 20240 6229
rect 20664 7805 20698 7821
rect 20664 6213 20698 6229
rect 21122 7805 21156 7821
rect 21122 6213 21156 6229
rect 21580 7805 21614 7821
rect 21580 6213 21614 6229
rect 13456 6136 13472 6170
rect 13692 6136 13708 6170
rect 13914 6136 13930 6170
rect 14150 6136 14166 6170
rect 14372 6136 14388 6170
rect 14608 6136 14624 6170
rect 14830 6136 14846 6170
rect 15066 6136 15082 6170
rect 15288 6136 15304 6170
rect 15524 6136 15540 6170
rect 15746 6136 15762 6170
rect 15982 6136 15998 6170
rect 16204 6136 16220 6170
rect 16440 6136 16456 6170
rect 16662 6136 16678 6170
rect 16898 6136 16914 6170
rect 17120 6136 17136 6170
rect 17356 6136 17372 6170
rect 17578 6136 17594 6170
rect 17814 6136 17830 6170
rect 18036 6136 18052 6170
rect 18272 6136 18288 6170
rect 18494 6136 18510 6170
rect 18730 6136 18746 6170
rect 18952 6136 18968 6170
rect 19188 6136 19204 6170
rect 19410 6136 19426 6170
rect 19646 6136 19662 6170
rect 19868 6136 19884 6170
rect 20104 6136 20120 6170
rect 20326 6136 20342 6170
rect 20562 6136 20578 6170
rect 20784 6136 20800 6170
rect 21020 6136 21036 6170
rect 21242 6136 21258 6170
rect 21478 6136 21494 6170
rect 12960 4766 13060 4928
rect 21884 4766 21984 4928
rect 23542 8456 23642 8618
rect 28886 8456 28986 8618
rect 29240 8617 29286 8652
rect 29373 8649 29699 8652
rect 29733 8652 29738 8700
rect 29144 8599 29186 8615
rect 29144 8565 29152 8599
rect 29144 8531 29186 8565
rect 29144 8497 29152 8531
rect 29144 8463 29186 8497
rect 29144 8429 29152 8463
rect 29144 8387 29186 8429
rect 29220 8599 29286 8617
rect 29733 8615 29786 8652
rect 29220 8565 29236 8599
rect 29270 8565 29286 8599
rect 29220 8531 29286 8565
rect 29220 8497 29236 8531
rect 29270 8497 29286 8531
rect 29220 8463 29286 8497
rect 29220 8429 29236 8463
rect 29270 8429 29286 8463
rect 29220 8421 29286 8429
rect 29378 8599 29431 8615
rect 29378 8565 29397 8599
rect 29378 8531 29431 8565
rect 29378 8497 29397 8531
rect 29378 8463 29431 8497
rect 29378 8429 29397 8463
rect 29378 8387 29431 8429
rect 29465 8599 29786 8615
rect 30570 8700 30640 8741
rect 30570 8652 30580 8700
rect 30628 8652 30640 8700
rect 30570 8631 30584 8652
rect 30618 8631 30640 8652
rect 30570 8611 30640 8631
rect 30674 8680 30720 8773
rect 30674 8646 30686 8680
rect 29465 8565 29481 8599
rect 29515 8581 29649 8599
rect 29515 8565 29531 8581
rect 29465 8531 29531 8565
rect 29633 8565 29649 8581
rect 29683 8577 29786 8599
rect 29683 8565 29699 8577
rect 29465 8497 29481 8531
rect 29515 8497 29531 8531
rect 29465 8463 29531 8497
rect 29465 8429 29481 8463
rect 29515 8429 29531 8463
rect 29465 8421 29531 8429
rect 29565 8531 29599 8547
rect 29565 8463 29599 8497
rect 29565 8387 29599 8429
rect 29633 8531 29699 8565
rect 29633 8497 29649 8531
rect 29683 8497 29699 8531
rect 29633 8463 29699 8497
rect 30227 8561 30285 8578
rect 30674 8577 30720 8646
rect 30227 8527 30239 8561
rect 30273 8527 30285 8561
rect 29633 8429 29649 8463
rect 29683 8429 29699 8463
rect 29633 8421 29699 8429
rect 29733 8463 29775 8479
rect 29767 8429 29775 8463
rect 30227 8433 30285 8527
rect 30587 8543 30720 8577
rect 30789 8791 30792 8825
rect 30927 8824 30977 8859
rect 31019 8854 31035 8888
rect 31069 8854 31240 8888
rect 30755 8739 30792 8791
rect 30916 8798 30977 8824
rect 31066 8807 31172 8820
rect 30755 8705 30757 8739
rect 30791 8705 30792 8739
rect 30587 8535 30621 8543
rect 30755 8535 30792 8705
rect 30826 8733 30882 8749
rect 30826 8699 30848 8733
rect 30826 8642 30882 8699
rect 30826 8594 30832 8642
rect 30880 8594 30882 8642
rect 30826 8559 30882 8594
rect 30916 8577 30950 8798
rect 31066 8773 31098 8807
rect 31132 8781 31172 8807
rect 30984 8739 31032 8760
rect 30984 8705 30995 8739
rect 31029 8705 31032 8739
rect 30984 8703 31032 8705
rect 30984 8669 30991 8703
rect 31025 8669 31032 8703
rect 30984 8641 31032 8669
rect 31066 8607 31100 8773
rect 31134 8747 31172 8781
rect 31206 8731 31240 8854
rect 31274 8833 31308 8867
rect 31274 8783 31308 8799
rect 31342 8893 31392 8909
rect 31342 8859 31358 8893
rect 31650 8893 31713 8943
rect 31342 8843 31392 8859
rect 31437 8849 31453 8883
rect 31487 8849 31614 8883
rect 31206 8715 31308 8731
rect 31206 8713 31274 8715
rect 30916 8551 30961 8577
rect 30995 8573 31011 8607
rect 31045 8573 31100 8607
rect 30995 8563 31100 8573
rect 31134 8681 31274 8713
rect 31134 8679 31308 8681
rect 30587 8485 30621 8501
rect 30655 8475 30671 8509
rect 30705 8475 30721 8509
rect 30789 8501 30792 8535
rect 30755 8485 30792 8501
rect 30843 8509 30893 8525
rect 30655 8433 30721 8475
rect 30843 8475 30859 8509
rect 30927 8523 30961 8551
rect 31134 8523 31168 8679
rect 31274 8665 31308 8679
rect 31210 8629 31250 8635
rect 31342 8629 31376 8843
rect 31410 8807 31448 8809
rect 31410 8773 31412 8807
rect 31446 8773 31448 8807
rect 31410 8715 31448 8773
rect 31444 8681 31448 8715
rect 31410 8665 31448 8681
rect 31482 8781 31546 8815
rect 31482 8747 31512 8781
rect 31482 8739 31546 8747
rect 31482 8705 31499 8739
rect 31533 8705 31546 8739
rect 31210 8619 31376 8629
rect 31482 8623 31546 8705
rect 31244 8585 31376 8619
rect 31210 8569 31376 8585
rect 30927 8489 30944 8523
rect 30978 8489 30994 8523
rect 31033 8489 31055 8523
rect 31089 8489 31168 8523
rect 31232 8517 31306 8533
rect 30843 8433 30893 8475
rect 31232 8483 31254 8517
rect 31288 8483 31306 8517
rect 31342 8523 31376 8569
rect 31453 8607 31546 8623
rect 31487 8573 31546 8607
rect 31453 8557 31546 8573
rect 31580 8681 31614 8849
rect 31650 8859 31652 8893
rect 31686 8859 31713 8893
rect 31650 8843 31713 8859
rect 31760 8901 31828 8909
rect 31760 8867 31776 8901
rect 31810 8867 31828 8901
rect 31760 8830 31828 8867
rect 31760 8797 31776 8830
rect 31648 8796 31776 8797
rect 31810 8796 31828 8830
rect 31648 8781 31828 8796
rect 31682 8759 31828 8781
rect 31682 8747 31776 8759
rect 31648 8725 31776 8747
rect 31810 8725 31828 8759
rect 31862 8871 31896 8943
rect 32034 8901 32100 8905
rect 31862 8791 31896 8837
rect 31862 8741 31896 8757
rect 31930 8895 31996 8900
rect 31930 8861 31946 8895
rect 31980 8861 31996 8895
rect 31930 8827 31996 8861
rect 31930 8793 31946 8827
rect 31980 8793 31996 8827
rect 31930 8759 31996 8793
rect 32034 8867 32050 8901
rect 32084 8867 32100 8901
rect 32034 8833 32100 8867
rect 32034 8799 32050 8833
rect 32084 8799 32100 8833
rect 32034 8759 32100 8799
rect 31648 8722 31828 8725
rect 31790 8681 31828 8722
rect 31930 8725 31946 8759
rect 31980 8731 31996 8759
rect 31980 8725 32012 8731
rect 31930 8715 32012 8725
rect 31965 8705 32012 8715
rect 31580 8665 31756 8681
rect 31580 8631 31722 8665
rect 31580 8615 31756 8631
rect 31790 8665 31940 8681
rect 31790 8631 31906 8665
rect 31790 8615 31940 8631
rect 31580 8523 31614 8615
rect 31790 8581 31830 8615
rect 31974 8589 32012 8705
rect 31963 8581 32012 8589
rect 31764 8578 31830 8581
rect 31764 8544 31780 8578
rect 31814 8544 31830 8578
rect 31932 8580 32012 8581
rect 31932 8562 31948 8580
rect 31982 8564 32012 8580
rect 32046 8681 32100 8759
rect 32138 8901 32181 8943
rect 32138 8867 32147 8901
rect 32138 8833 32181 8867
rect 32138 8799 32147 8833
rect 32138 8765 32181 8799
rect 32138 8731 32147 8765
rect 32138 8715 32181 8731
rect 32215 8901 32282 8909
rect 32215 8867 32231 8901
rect 32265 8867 32282 8901
rect 32215 8830 32282 8867
rect 32215 8796 32231 8830
rect 32265 8796 32282 8830
rect 32215 8759 32282 8796
rect 32215 8725 32231 8759
rect 32265 8725 32282 8759
rect 32215 8712 32282 8725
rect 32368 8901 32410 8943
rect 32368 8867 32376 8901
rect 32368 8833 32410 8867
rect 32368 8799 32376 8833
rect 32368 8765 32410 8799
rect 32368 8731 32376 8765
rect 32368 8715 32410 8731
rect 32444 8901 32510 8909
rect 32444 8867 32460 8901
rect 32494 8867 32510 8901
rect 32444 8833 32510 8867
rect 32444 8799 32460 8833
rect 32494 8799 32510 8833
rect 32444 8765 32510 8799
rect 32444 8731 32460 8765
rect 32494 8731 32510 8765
rect 32444 8713 32510 8731
rect 32602 8901 32655 8943
rect 32602 8867 32621 8901
rect 32602 8833 32655 8867
rect 32602 8799 32621 8833
rect 32602 8765 32655 8799
rect 32602 8731 32621 8765
rect 32602 8715 32655 8731
rect 32689 8901 32755 8909
rect 32689 8867 32705 8901
rect 32739 8867 32755 8901
rect 32689 8833 32755 8867
rect 32689 8799 32705 8833
rect 32739 8799 32755 8833
rect 32689 8765 32755 8799
rect 32789 8901 32823 8943
rect 32789 8833 32823 8867
rect 32789 8783 32823 8799
rect 32857 8901 32923 8909
rect 32857 8867 32873 8901
rect 32907 8867 32923 8901
rect 32857 8833 32923 8867
rect 32957 8901 32999 8943
rect 32991 8867 32999 8901
rect 32957 8851 32999 8867
rect 33127 8872 33185 8943
rect 32857 8799 32873 8833
rect 32907 8799 32923 8833
rect 32689 8731 32705 8765
rect 32739 8749 32755 8765
rect 32857 8765 32923 8799
rect 32857 8749 32873 8765
rect 32739 8731 32873 8749
rect 32907 8753 32923 8765
rect 33127 8838 33139 8872
rect 33173 8838 33185 8872
rect 33127 8779 33185 8838
rect 32907 8731 33010 8753
rect 32689 8715 33010 8731
rect 32046 8665 32201 8681
rect 32046 8631 32167 8665
rect 32046 8615 32201 8631
rect 32235 8680 32282 8712
rect 32464 8680 32510 8713
rect 32597 8680 32923 8681
rect 32235 8632 32242 8680
rect 32406 8665 32430 8679
rect 31982 8562 31998 8564
rect 31342 8489 31373 8523
rect 31407 8489 31423 8523
rect 31457 8489 31476 8523
rect 31510 8489 31614 8523
rect 31669 8523 31711 8539
rect 31669 8489 31674 8523
rect 31708 8489 31711 8523
rect 31232 8433 31306 8483
rect 31669 8433 31711 8489
rect 31764 8510 31830 8544
rect 31764 8476 31780 8510
rect 31814 8476 31830 8510
rect 31864 8539 31898 8555
rect 31864 8433 31898 8505
rect 31932 8514 31936 8562
rect 31984 8514 31998 8562
rect 32046 8539 32086 8615
rect 32235 8598 32282 8632
rect 32364 8631 32380 8632
rect 32414 8631 32430 8665
rect 32464 8632 32470 8680
rect 32597 8632 32602 8680
rect 32650 8665 32712 8680
rect 32760 8665 32828 8680
rect 32876 8665 32923 8680
rect 32650 8632 32705 8665
rect 32760 8632 32789 8665
rect 31932 8512 31998 8514
rect 31932 8478 31948 8512
rect 31982 8478 31998 8512
rect 32036 8535 32086 8539
rect 32036 8501 32052 8535
rect 32231 8547 32282 8598
rect 32036 8485 32086 8501
rect 32133 8509 32197 8525
rect 31932 8477 31998 8478
rect 32133 8475 32147 8509
rect 32181 8475 32197 8509
rect 32133 8433 32197 8475
rect 32265 8513 32282 8547
rect 32231 8467 32282 8513
rect 32364 8581 32410 8597
rect 32464 8593 32510 8632
rect 32597 8631 32613 8632
rect 32647 8631 32705 8632
rect 32739 8631 32789 8632
rect 32823 8632 32828 8665
rect 32823 8631 32873 8632
rect 32907 8631 32923 8665
rect 32957 8678 33010 8715
rect 33127 8745 33139 8779
rect 33173 8745 33185 8779
rect 33127 8710 33185 8745
rect 36001 8872 36059 8943
rect 36001 8838 36013 8872
rect 36047 8838 36059 8872
rect 36001 8779 36059 8838
rect 36001 8745 36013 8779
rect 36047 8745 36059 8779
rect 36001 8710 36059 8745
rect 32957 8630 32960 8678
rect 33008 8630 33010 8678
rect 32957 8597 33010 8630
rect 32364 8547 32376 8581
rect 32364 8513 32410 8547
rect 32364 8479 32376 8513
rect 32364 8433 32410 8479
rect 32444 8581 32510 8593
rect 32444 8547 32460 8581
rect 32494 8547 32510 8581
rect 32444 8513 32510 8547
rect 32689 8561 33010 8597
rect 33127 8561 33185 8578
rect 32444 8479 32460 8513
rect 32494 8479 32510 8513
rect 32444 8467 32510 8479
rect 32602 8509 32655 8525
rect 32602 8475 32621 8509
rect 32602 8433 32655 8475
rect 32689 8517 32755 8561
rect 32689 8483 32705 8517
rect 32739 8483 32755 8517
rect 32689 8467 32755 8483
rect 32789 8509 32823 8525
rect 32789 8433 32823 8475
rect 32857 8517 32923 8561
rect 33127 8527 33139 8561
rect 33173 8527 33185 8561
rect 32857 8483 32873 8517
rect 32907 8483 32923 8517
rect 32857 8467 32923 8483
rect 32957 8510 33007 8526
rect 32991 8476 33007 8510
rect 32957 8433 33007 8476
rect 33127 8433 33185 8527
rect 36001 8561 36059 8578
rect 36001 8527 36013 8561
rect 36047 8527 36059 8561
rect 36001 8433 36059 8527
rect 29733 8387 29775 8429
rect 30210 8399 30239 8433
rect 30273 8399 30302 8433
rect 30552 8399 30581 8433
rect 30615 8399 30673 8433
rect 30707 8399 30765 8433
rect 30799 8399 30857 8433
rect 30891 8399 30949 8433
rect 30983 8399 31041 8433
rect 31075 8399 31133 8433
rect 31167 8399 31225 8433
rect 31259 8399 31317 8433
rect 31351 8399 31409 8433
rect 31443 8399 31501 8433
rect 31535 8399 31593 8433
rect 31627 8399 31685 8433
rect 31719 8399 31777 8433
rect 31811 8399 31869 8433
rect 31903 8399 31961 8433
rect 31995 8399 32053 8433
rect 32087 8399 32145 8433
rect 32179 8399 32237 8433
rect 32271 8399 32329 8433
rect 32363 8399 32421 8433
rect 32455 8399 32513 8433
rect 32547 8399 32605 8433
rect 32639 8399 32697 8433
rect 32731 8399 32789 8433
rect 32823 8399 32881 8433
rect 32915 8399 32973 8433
rect 33007 8399 33036 8433
rect 33110 8399 33139 8433
rect 33173 8399 33202 8433
rect 33250 8399 33279 8433
rect 33313 8399 33371 8433
rect 33405 8399 33463 8433
rect 33497 8399 33555 8433
rect 33589 8399 33647 8433
rect 33681 8399 33739 8433
rect 33773 8399 33831 8433
rect 33865 8399 33923 8433
rect 33957 8399 34015 8433
rect 34049 8399 34107 8433
rect 34141 8399 34199 8433
rect 34233 8399 34291 8433
rect 34325 8399 34383 8433
rect 34417 8399 34475 8433
rect 34509 8399 34567 8433
rect 34601 8399 34659 8433
rect 34693 8399 34751 8433
rect 34785 8399 34843 8433
rect 34877 8399 34935 8433
rect 34969 8399 35027 8433
rect 35061 8399 35119 8433
rect 35153 8399 35211 8433
rect 35245 8399 35303 8433
rect 35337 8399 35395 8433
rect 35429 8399 35487 8433
rect 35521 8399 35579 8433
rect 35613 8399 35671 8433
rect 35705 8399 35734 8433
rect 35984 8399 36013 8433
rect 36047 8399 36076 8433
rect 29076 8353 29105 8387
rect 29139 8353 29197 8387
rect 29231 8353 29289 8387
rect 29323 8353 29381 8387
rect 29415 8353 29473 8387
rect 29507 8353 29565 8387
rect 29599 8353 29657 8387
rect 29691 8353 29749 8387
rect 29783 8353 29812 8387
rect 24051 8284 24067 8318
rect 24287 8284 24303 8318
rect 24509 8284 24525 8318
rect 24745 8284 24761 8318
rect 24967 8284 24983 8318
rect 25203 8284 25219 8318
rect 25425 8284 25441 8318
rect 25661 8284 25677 8318
rect 25883 8284 25899 8318
rect 26119 8284 26135 8318
rect 26341 8284 26357 8318
rect 26577 8284 26593 8318
rect 26799 8284 26815 8318
rect 27035 8284 27051 8318
rect 27257 8284 27273 8318
rect 27493 8284 27509 8318
rect 27715 8284 27731 8318
rect 27951 8284 27967 8318
rect 28173 8284 28189 8318
rect 28409 8284 28425 8318
rect 23931 8225 23965 8241
rect 23931 7033 23965 7049
rect 24389 8225 24423 8241
rect 24389 7033 24423 7049
rect 24847 8225 24881 8241
rect 24847 7033 24881 7049
rect 25305 8225 25339 8241
rect 25305 7033 25339 7049
rect 25763 8225 25797 8241
rect 25763 7033 25797 7049
rect 26221 8225 26255 8241
rect 26221 7033 26255 7049
rect 26679 8225 26713 8241
rect 26679 7033 26713 7049
rect 27137 8225 27171 8241
rect 27137 7033 27171 7049
rect 27595 8225 27629 8241
rect 27595 7033 27629 7049
rect 28053 8225 28087 8241
rect 28053 7033 28087 7049
rect 28511 8225 28545 8241
rect 28511 7033 28545 7049
rect 24051 6956 24067 6990
rect 24287 6956 24303 6990
rect 24509 6956 24525 6990
rect 24745 6956 24761 6990
rect 24967 6956 24983 6990
rect 25203 6956 25219 6990
rect 25425 6956 25441 6990
rect 25661 6956 25677 6990
rect 25883 6956 25899 6990
rect 26119 6956 26135 6990
rect 26341 6956 26357 6990
rect 26577 6956 26593 6990
rect 26799 6956 26815 6990
rect 27035 6956 27051 6990
rect 27257 6956 27273 6990
rect 27493 6956 27509 6990
rect 27715 6956 27731 6990
rect 27951 6956 27967 6990
rect 28173 6956 28189 6990
rect 28409 6956 28425 6990
rect 23542 4766 23642 4928
rect 30227 8305 30285 8399
rect 30655 8357 30721 8399
rect 30227 8271 30239 8305
rect 30273 8271 30285 8305
rect 30227 8254 30285 8271
rect 30587 8331 30621 8347
rect 30655 8323 30671 8357
rect 30705 8323 30721 8357
rect 30843 8357 30893 8399
rect 30755 8331 30792 8347
rect 30587 8289 30621 8297
rect 30789 8297 30792 8331
rect 30843 8323 30859 8357
rect 31232 8349 31306 8399
rect 30843 8307 30893 8323
rect 30927 8309 30944 8343
rect 30978 8309 30994 8343
rect 31033 8309 31055 8343
rect 31089 8309 31168 8343
rect 30587 8255 30720 8289
rect 30570 8201 30640 8221
rect 30570 8190 30584 8201
rect 30618 8190 30640 8201
rect 30570 8142 30576 8190
rect 30624 8142 30640 8190
rect 30227 8087 30285 8122
rect 30570 8091 30640 8142
rect 30674 8186 30720 8255
rect 30674 8152 30686 8186
rect 30227 8053 30239 8087
rect 30273 8053 30285 8087
rect 30674 8059 30720 8152
rect 30674 8057 30678 8059
rect 30227 7994 30285 8053
rect 30227 7960 30239 7994
rect 30273 7960 30285 7994
rect 30227 7889 30285 7960
rect 30587 8041 30678 8057
rect 30621 8025 30678 8041
rect 30712 8025 30720 8059
rect 30621 8023 30720 8025
rect 30755 8127 30792 8297
rect 30927 8281 30961 8309
rect 30755 8093 30757 8127
rect 30791 8093 30792 8127
rect 30755 8041 30792 8093
rect 30826 8238 30882 8273
rect 30826 8190 30832 8238
rect 30880 8190 30882 8238
rect 30826 8133 30882 8190
rect 30826 8099 30848 8133
rect 30826 8083 30882 8099
rect 30916 8255 30961 8281
rect 30995 8259 31100 8269
rect 30587 7973 30621 8007
rect 30789 8007 30792 8041
rect 30916 8034 30950 8255
rect 30995 8225 31011 8259
rect 31045 8225 31100 8259
rect 30984 8163 31032 8191
rect 30984 8129 30991 8163
rect 31025 8129 31032 8163
rect 30984 8127 31032 8129
rect 30984 8093 30995 8127
rect 31029 8093 31032 8127
rect 30984 8072 31032 8093
rect 31066 8059 31100 8225
rect 31134 8153 31168 8309
rect 31232 8315 31254 8349
rect 31288 8315 31306 8349
rect 31669 8343 31711 8399
rect 31232 8299 31306 8315
rect 31342 8309 31373 8343
rect 31407 8309 31423 8343
rect 31457 8309 31476 8343
rect 31510 8309 31614 8343
rect 31342 8263 31376 8309
rect 31210 8247 31376 8263
rect 31244 8213 31376 8247
rect 31210 8203 31376 8213
rect 31453 8259 31546 8275
rect 31487 8225 31546 8259
rect 31453 8209 31546 8225
rect 31210 8197 31250 8203
rect 31274 8153 31308 8167
rect 31134 8151 31308 8153
rect 31134 8119 31274 8151
rect 31206 8117 31274 8119
rect 31206 8101 31308 8117
rect 30916 8008 30977 8034
rect 31066 8025 31098 8059
rect 31134 8051 31172 8085
rect 31132 8025 31172 8051
rect 31066 8012 31172 8025
rect 30587 7923 30621 7939
rect 30655 7955 30671 7989
rect 30705 7955 30721 7989
rect 30655 7889 30721 7955
rect 30755 7973 30792 8007
rect 30789 7939 30792 7973
rect 30755 7923 30792 7939
rect 30840 7965 30893 7981
rect 30840 7931 30859 7965
rect 30840 7889 30893 7931
rect 30927 7973 30977 8008
rect 31206 7978 31240 8101
rect 30927 7939 30943 7973
rect 31019 7944 31035 7978
rect 31069 7944 31240 7978
rect 31274 8033 31308 8049
rect 31274 7965 31308 7999
rect 30927 7923 30977 7939
rect 31274 7889 31308 7931
rect 31342 7989 31376 8203
rect 31410 8151 31448 8167
rect 31444 8117 31448 8151
rect 31410 8059 31448 8117
rect 31410 8025 31412 8059
rect 31446 8025 31448 8059
rect 31410 8023 31448 8025
rect 31482 8127 31546 8209
rect 31482 8093 31499 8127
rect 31533 8093 31546 8127
rect 31482 8085 31546 8093
rect 31482 8051 31512 8085
rect 31482 8017 31546 8051
rect 31580 8217 31614 8309
rect 31669 8309 31674 8343
rect 31708 8309 31711 8343
rect 31669 8293 31711 8309
rect 31764 8322 31780 8356
rect 31814 8322 31830 8356
rect 31764 8288 31830 8322
rect 31764 8254 31780 8288
rect 31814 8254 31830 8288
rect 31864 8327 31898 8399
rect 32133 8357 32197 8399
rect 31864 8277 31898 8293
rect 31932 8354 31998 8355
rect 31932 8320 31948 8354
rect 31982 8320 31998 8354
rect 31932 8286 31998 8320
rect 32036 8331 32086 8347
rect 32036 8297 32052 8331
rect 32133 8323 32147 8357
rect 32181 8323 32197 8357
rect 32133 8307 32197 8323
rect 32231 8319 32282 8365
rect 32036 8293 32086 8297
rect 31764 8251 31830 8254
rect 31932 8252 31948 8286
rect 31982 8268 31998 8286
rect 31982 8252 32012 8268
rect 31932 8251 32012 8252
rect 31790 8217 31830 8251
rect 31963 8243 32012 8251
rect 31580 8201 31756 8217
rect 31580 8167 31722 8201
rect 31580 8151 31756 8167
rect 31790 8201 31940 8217
rect 31790 8167 31906 8201
rect 31790 8151 31940 8167
rect 31342 7973 31392 7989
rect 31580 7983 31614 8151
rect 31790 8110 31828 8151
rect 31974 8127 32012 8243
rect 31965 8117 32012 8127
rect 31648 8107 31828 8110
rect 31648 8085 31776 8107
rect 31682 8073 31776 8085
rect 31810 8073 31828 8107
rect 31930 8107 32012 8117
rect 31682 8051 31828 8073
rect 31648 8036 31828 8051
rect 31648 8035 31776 8036
rect 31760 8002 31776 8035
rect 31810 8002 31828 8036
rect 31342 7939 31358 7973
rect 31437 7949 31453 7983
rect 31487 7949 31614 7983
rect 31650 7973 31713 7989
rect 31342 7923 31392 7939
rect 31650 7939 31652 7973
rect 31686 7939 31713 7973
rect 31650 7889 31713 7939
rect 31760 7965 31828 8002
rect 31760 7931 31776 7965
rect 31810 7931 31828 7965
rect 31760 7923 31828 7931
rect 31862 8075 31896 8091
rect 31862 7995 31896 8041
rect 31862 7889 31896 7961
rect 31930 8073 31946 8107
rect 31980 8101 32012 8107
rect 32046 8217 32086 8293
rect 32265 8285 32282 8319
rect 32231 8234 32282 8285
rect 32364 8353 32410 8399
rect 32364 8319 32376 8353
rect 32364 8285 32410 8319
rect 32364 8251 32376 8285
rect 32364 8235 32410 8251
rect 32444 8353 32510 8365
rect 32444 8319 32460 8353
rect 32494 8319 32510 8353
rect 32444 8285 32510 8319
rect 32602 8357 32655 8399
rect 32602 8323 32621 8357
rect 32602 8307 32655 8323
rect 32689 8349 32755 8365
rect 32689 8315 32705 8349
rect 32739 8315 32755 8349
rect 32444 8251 32460 8285
rect 32494 8251 32510 8285
rect 32444 8239 32510 8251
rect 32046 8201 32201 8217
rect 32046 8167 32167 8201
rect 32046 8151 32201 8167
rect 32235 8200 32282 8234
rect 32364 8200 32380 8201
rect 32235 8152 32242 8200
rect 32414 8167 32430 8201
rect 32406 8153 32430 8167
rect 32464 8200 32510 8239
rect 32689 8271 32755 8315
rect 32789 8357 32823 8399
rect 32789 8307 32823 8323
rect 32857 8349 32923 8365
rect 32857 8315 32873 8349
rect 32907 8315 32923 8349
rect 32857 8271 32923 8315
rect 32957 8356 33007 8399
rect 32991 8322 33007 8356
rect 33353 8357 33419 8399
rect 32957 8306 33007 8322
rect 33285 8331 33319 8347
rect 33353 8323 33369 8357
rect 33403 8323 33419 8357
rect 33541 8357 33591 8399
rect 33453 8331 33490 8347
rect 33285 8289 33319 8297
rect 33487 8297 33490 8331
rect 33541 8323 33557 8357
rect 33930 8349 34004 8399
rect 33541 8307 33591 8323
rect 33625 8309 33642 8343
rect 33676 8309 33692 8343
rect 33731 8309 33753 8343
rect 33787 8309 33866 8343
rect 32689 8235 33010 8271
rect 33285 8255 33418 8289
rect 32957 8202 33010 8235
rect 32597 8200 32613 8201
rect 32647 8200 32705 8201
rect 32739 8200 32789 8201
rect 32464 8152 32470 8200
rect 32597 8152 32602 8200
rect 32650 8167 32705 8200
rect 32760 8167 32789 8200
rect 32823 8200 32873 8201
rect 32823 8167 32828 8200
rect 32907 8167 32923 8201
rect 32650 8152 32712 8167
rect 32760 8152 32828 8167
rect 32876 8152 32923 8167
rect 31980 8073 31996 8101
rect 32046 8073 32100 8151
rect 32235 8120 32282 8152
rect 31930 8039 31996 8073
rect 31930 8016 31946 8039
rect 31980 8016 31996 8039
rect 31930 7968 31936 8016
rect 31984 7968 31996 8016
rect 31930 7937 31946 7968
rect 31980 7937 31996 7968
rect 31930 7932 31996 7937
rect 32034 8033 32100 8073
rect 32034 7999 32050 8033
rect 32084 7999 32100 8033
rect 32034 7965 32100 7999
rect 32034 7931 32050 7965
rect 32084 7931 32100 7965
rect 32034 7927 32100 7931
rect 32138 8101 32181 8117
rect 32138 8067 32147 8101
rect 32138 8033 32181 8067
rect 32138 7999 32147 8033
rect 32138 7965 32181 7999
rect 32138 7931 32147 7965
rect 32138 7889 32181 7931
rect 32215 8107 32282 8120
rect 32464 8119 32510 8152
rect 32597 8151 32923 8152
rect 32957 8154 32964 8202
rect 33268 8201 33338 8221
rect 33268 8167 33282 8201
rect 33316 8167 33338 8201
rect 32215 8073 32231 8107
rect 32265 8073 32282 8107
rect 32215 8036 32282 8073
rect 32215 8002 32231 8036
rect 32265 8002 32282 8036
rect 32215 7965 32282 8002
rect 32215 7931 32231 7965
rect 32265 7931 32282 7965
rect 32215 7923 32282 7931
rect 32368 8101 32410 8117
rect 32368 8067 32376 8101
rect 32368 8033 32410 8067
rect 32368 7999 32376 8033
rect 32368 7965 32410 7999
rect 32368 7931 32376 7965
rect 32368 7889 32410 7931
rect 32444 8101 32510 8119
rect 32957 8117 33010 8154
rect 32444 8067 32460 8101
rect 32494 8067 32510 8101
rect 32444 8033 32510 8067
rect 32444 7999 32460 8033
rect 32494 7999 32510 8033
rect 32444 7965 32510 7999
rect 32444 7931 32460 7965
rect 32494 7931 32510 7965
rect 32444 7923 32510 7931
rect 32602 8101 32655 8117
rect 32602 8067 32621 8101
rect 32602 8033 32655 8067
rect 32602 7999 32621 8033
rect 32602 7965 32655 7999
rect 32602 7931 32621 7965
rect 32602 7889 32655 7931
rect 32689 8101 33010 8117
rect 32689 8067 32705 8101
rect 32739 8083 32873 8101
rect 32739 8067 32755 8083
rect 32689 8033 32755 8067
rect 32857 8067 32873 8083
rect 32907 8079 33010 8101
rect 33268 8148 33338 8167
rect 33268 8100 33274 8148
rect 33322 8100 33338 8148
rect 33268 8091 33338 8100
rect 33372 8186 33418 8255
rect 33372 8152 33384 8186
rect 32907 8067 32923 8079
rect 32689 7999 32705 8033
rect 32739 7999 32755 8033
rect 32689 7965 32755 7999
rect 32689 7931 32705 7965
rect 32739 7931 32755 7965
rect 32689 7923 32755 7931
rect 32789 8033 32823 8049
rect 32789 7965 32823 7999
rect 32789 7889 32823 7931
rect 32857 8033 32923 8067
rect 33372 8059 33418 8152
rect 33372 8057 33376 8059
rect 32857 7999 32873 8033
rect 32907 7999 32923 8033
rect 32857 7965 32923 7999
rect 33285 8041 33376 8057
rect 33319 8025 33376 8041
rect 33410 8025 33418 8059
rect 33319 8023 33418 8025
rect 33453 8127 33490 8297
rect 33625 8281 33659 8309
rect 33453 8093 33455 8127
rect 33489 8093 33490 8127
rect 33453 8041 33490 8093
rect 33524 8238 33580 8273
rect 33524 8190 33530 8238
rect 33578 8190 33580 8238
rect 33524 8133 33580 8190
rect 33524 8099 33546 8133
rect 33524 8083 33580 8099
rect 33614 8255 33659 8281
rect 33693 8259 33798 8269
rect 32857 7931 32873 7965
rect 32907 7931 32923 7965
rect 32857 7923 32923 7931
rect 32957 7965 32999 7981
rect 32991 7931 32999 7965
rect 32957 7889 32999 7931
rect 33285 7973 33319 8007
rect 33487 8007 33490 8041
rect 33614 8034 33648 8255
rect 33693 8225 33709 8259
rect 33743 8225 33798 8259
rect 33682 8163 33730 8191
rect 33682 8129 33689 8163
rect 33723 8129 33730 8163
rect 33682 8127 33730 8129
rect 33682 8093 33693 8127
rect 33727 8093 33730 8127
rect 33682 8072 33730 8093
rect 33764 8059 33798 8225
rect 33832 8153 33866 8309
rect 33930 8315 33952 8349
rect 33986 8315 34004 8349
rect 34367 8343 34409 8399
rect 33930 8299 34004 8315
rect 34040 8309 34071 8343
rect 34105 8309 34121 8343
rect 34155 8309 34174 8343
rect 34208 8309 34312 8343
rect 34040 8263 34074 8309
rect 33908 8247 34074 8263
rect 33942 8213 34074 8247
rect 33908 8203 34074 8213
rect 34151 8259 34244 8275
rect 34185 8225 34244 8259
rect 34151 8209 34244 8225
rect 33908 8197 33948 8203
rect 33972 8153 34006 8167
rect 33832 8151 34006 8153
rect 33832 8119 33972 8151
rect 33904 8117 33972 8119
rect 33904 8101 34006 8117
rect 33614 8008 33675 8034
rect 33764 8025 33796 8059
rect 33832 8051 33870 8085
rect 33830 8025 33870 8051
rect 33764 8012 33870 8025
rect 33285 7923 33319 7939
rect 33353 7955 33369 7989
rect 33403 7955 33419 7989
rect 33353 7889 33419 7955
rect 33453 7973 33490 8007
rect 33487 7939 33490 7973
rect 33453 7923 33490 7939
rect 33538 7965 33591 7981
rect 33538 7931 33557 7965
rect 33538 7889 33591 7931
rect 33625 7973 33675 8008
rect 33904 7978 33938 8101
rect 33625 7939 33641 7973
rect 33717 7944 33733 7978
rect 33767 7944 33938 7978
rect 33972 8033 34006 8049
rect 33972 7965 34006 7999
rect 33625 7923 33675 7939
rect 33972 7889 34006 7931
rect 34040 7989 34074 8203
rect 34108 8151 34146 8167
rect 34142 8117 34146 8151
rect 34108 8059 34146 8117
rect 34108 8025 34110 8059
rect 34144 8025 34146 8059
rect 34108 8023 34146 8025
rect 34180 8127 34244 8209
rect 34180 8093 34197 8127
rect 34231 8093 34244 8127
rect 34180 8085 34244 8093
rect 34180 8051 34210 8085
rect 34180 8017 34244 8051
rect 34278 8217 34312 8309
rect 34367 8309 34372 8343
rect 34406 8309 34409 8343
rect 34367 8293 34409 8309
rect 34462 8322 34478 8356
rect 34512 8322 34528 8356
rect 34462 8288 34528 8322
rect 34462 8254 34478 8288
rect 34512 8254 34528 8288
rect 34562 8327 34596 8399
rect 34831 8357 34895 8399
rect 34562 8277 34596 8293
rect 34630 8354 34696 8355
rect 34630 8320 34646 8354
rect 34680 8320 34696 8354
rect 34630 8314 34696 8320
rect 34462 8251 34528 8254
rect 34630 8266 34636 8314
rect 34684 8268 34696 8314
rect 34734 8331 34784 8347
rect 34734 8297 34750 8331
rect 34831 8323 34845 8357
rect 34879 8323 34895 8357
rect 34831 8307 34895 8323
rect 34929 8319 34980 8365
rect 34734 8293 34784 8297
rect 34684 8266 34710 8268
rect 34630 8252 34646 8266
rect 34680 8252 34710 8266
rect 34630 8251 34710 8252
rect 34488 8217 34528 8251
rect 34661 8243 34710 8251
rect 34278 8201 34454 8217
rect 34278 8167 34420 8201
rect 34278 8151 34454 8167
rect 34488 8201 34638 8217
rect 34488 8167 34604 8201
rect 34488 8151 34638 8167
rect 34040 7973 34090 7989
rect 34278 7983 34312 8151
rect 34488 8110 34526 8151
rect 34672 8127 34710 8243
rect 34663 8117 34710 8127
rect 34346 8107 34526 8110
rect 34346 8085 34474 8107
rect 34380 8073 34474 8085
rect 34508 8073 34526 8107
rect 34628 8107 34710 8117
rect 34380 8051 34526 8073
rect 34346 8036 34526 8051
rect 34346 8035 34474 8036
rect 34458 8002 34474 8035
rect 34508 8002 34526 8036
rect 34040 7939 34056 7973
rect 34135 7949 34151 7983
rect 34185 7949 34312 7983
rect 34348 7973 34411 7989
rect 34040 7923 34090 7939
rect 34348 7939 34350 7973
rect 34384 7939 34411 7973
rect 34348 7889 34411 7939
rect 34458 7965 34526 8002
rect 34458 7931 34474 7965
rect 34508 7931 34526 7965
rect 34458 7923 34526 7931
rect 34560 8075 34594 8091
rect 34560 7995 34594 8041
rect 34560 7889 34594 7961
rect 34628 8073 34644 8107
rect 34678 8101 34710 8107
rect 34744 8217 34784 8293
rect 34963 8285 34980 8319
rect 34929 8234 34980 8285
rect 35062 8353 35108 8399
rect 35062 8319 35074 8353
rect 35062 8285 35108 8319
rect 35062 8251 35074 8285
rect 35062 8235 35108 8251
rect 35142 8353 35208 8365
rect 35142 8319 35158 8353
rect 35192 8319 35208 8353
rect 35142 8285 35208 8319
rect 35300 8357 35353 8399
rect 35300 8323 35319 8357
rect 35300 8307 35353 8323
rect 35387 8349 35453 8365
rect 35387 8315 35403 8349
rect 35437 8315 35453 8349
rect 35142 8251 35158 8285
rect 35192 8251 35208 8285
rect 35142 8239 35208 8251
rect 34744 8201 34899 8217
rect 34744 8167 34865 8201
rect 34744 8151 34899 8167
rect 34933 8200 34980 8234
rect 35062 8200 35078 8201
rect 34933 8152 34940 8200
rect 35112 8167 35128 8201
rect 35104 8153 35128 8167
rect 35162 8200 35208 8239
rect 35387 8271 35453 8315
rect 35487 8357 35521 8399
rect 35487 8307 35521 8323
rect 35555 8349 35621 8365
rect 35555 8315 35571 8349
rect 35605 8315 35621 8349
rect 35555 8271 35621 8315
rect 35655 8356 35705 8399
rect 35689 8322 35705 8356
rect 35655 8306 35705 8322
rect 36001 8305 36059 8399
rect 36001 8271 36013 8305
rect 36047 8271 36059 8305
rect 35387 8235 35708 8271
rect 36001 8254 36059 8271
rect 35655 8202 35708 8235
rect 35295 8200 35311 8201
rect 35345 8200 35403 8201
rect 35437 8200 35487 8201
rect 35162 8152 35168 8200
rect 35295 8152 35300 8200
rect 35348 8167 35403 8200
rect 35458 8167 35487 8200
rect 35521 8200 35571 8201
rect 35521 8167 35526 8200
rect 35605 8167 35621 8201
rect 35348 8152 35410 8167
rect 35458 8152 35526 8167
rect 35574 8152 35621 8167
rect 34678 8073 34694 8101
rect 34744 8073 34798 8151
rect 34933 8120 34980 8152
rect 34628 8039 34694 8073
rect 34628 8005 34644 8039
rect 34678 8005 34694 8039
rect 34628 7971 34694 8005
rect 34628 7937 34644 7971
rect 34678 7937 34694 7971
rect 34628 7932 34694 7937
rect 34732 8033 34798 8073
rect 34732 7999 34748 8033
rect 34782 7999 34798 8033
rect 34732 7965 34798 7999
rect 34732 7931 34748 7965
rect 34782 7931 34798 7965
rect 34732 7927 34798 7931
rect 34836 8101 34879 8117
rect 34836 8067 34845 8101
rect 34836 8033 34879 8067
rect 34836 7999 34845 8033
rect 34836 7965 34879 7999
rect 34836 7931 34845 7965
rect 34836 7889 34879 7931
rect 34913 8107 34980 8120
rect 35162 8119 35208 8152
rect 35295 8151 35621 8152
rect 35655 8154 35658 8202
rect 35706 8154 35708 8202
rect 34913 8073 34929 8107
rect 34963 8073 34980 8107
rect 34913 8036 34980 8073
rect 34913 8002 34929 8036
rect 34963 8002 34980 8036
rect 34913 7965 34980 8002
rect 34913 7931 34929 7965
rect 34963 7931 34980 7965
rect 34913 7923 34980 7931
rect 35066 8101 35108 8117
rect 35066 8067 35074 8101
rect 35066 8033 35108 8067
rect 35066 7999 35074 8033
rect 35066 7965 35108 7999
rect 35066 7931 35074 7965
rect 35066 7889 35108 7931
rect 35142 8101 35208 8119
rect 35655 8117 35708 8154
rect 35142 8067 35158 8101
rect 35192 8067 35208 8101
rect 35142 8033 35208 8067
rect 35142 7999 35158 8033
rect 35192 7999 35208 8033
rect 35142 7965 35208 7999
rect 35142 7931 35158 7965
rect 35192 7931 35208 7965
rect 35142 7923 35208 7931
rect 35300 8101 35353 8117
rect 35300 8067 35319 8101
rect 35300 8033 35353 8067
rect 35300 7999 35319 8033
rect 35300 7965 35353 7999
rect 35300 7931 35319 7965
rect 35300 7889 35353 7931
rect 35387 8101 35708 8117
rect 35387 8067 35403 8101
rect 35437 8083 35571 8101
rect 35437 8067 35453 8083
rect 35387 8033 35453 8067
rect 35555 8067 35571 8083
rect 35605 8079 35708 8101
rect 36001 8087 36059 8122
rect 35605 8067 35621 8079
rect 35387 7999 35403 8033
rect 35437 7999 35453 8033
rect 35387 7965 35453 7999
rect 35387 7931 35403 7965
rect 35437 7931 35453 7965
rect 35387 7923 35453 7931
rect 35487 8033 35521 8049
rect 35487 7965 35521 7999
rect 35487 7889 35521 7931
rect 35555 8033 35621 8067
rect 35555 7999 35571 8033
rect 35605 7999 35621 8033
rect 35555 7965 35621 7999
rect 36001 8053 36013 8087
rect 36047 8053 36059 8087
rect 36001 7994 36059 8053
rect 35555 7931 35571 7965
rect 35605 7931 35621 7965
rect 35555 7923 35621 7931
rect 35655 7965 35697 7981
rect 35689 7931 35697 7965
rect 35655 7889 35697 7931
rect 36001 7960 36013 7994
rect 36047 7960 36059 7994
rect 36001 7889 36059 7960
rect 30210 7855 30239 7889
rect 30273 7855 30302 7889
rect 30552 7855 30581 7889
rect 30615 7855 30673 7889
rect 30707 7855 30765 7889
rect 30799 7855 30857 7889
rect 30891 7855 30949 7889
rect 30983 7855 31041 7889
rect 31075 7855 31133 7889
rect 31167 7855 31225 7889
rect 31259 7855 31317 7889
rect 31351 7855 31409 7889
rect 31443 7855 31501 7889
rect 31535 7855 31593 7889
rect 31627 7855 31685 7889
rect 31719 7855 31777 7889
rect 31811 7855 31869 7889
rect 31903 7855 31961 7889
rect 31995 7855 32053 7889
rect 32087 7855 32145 7889
rect 32179 7855 32237 7889
rect 32271 7855 32329 7889
rect 32363 7855 32421 7889
rect 32455 7855 32513 7889
rect 32547 7855 32605 7889
rect 32639 7855 32697 7889
rect 32731 7855 32789 7889
rect 32823 7855 32881 7889
rect 32915 7855 32973 7889
rect 33007 7855 33036 7889
rect 33250 7855 33279 7889
rect 33313 7855 33371 7889
rect 33405 7855 33463 7889
rect 33497 7855 33555 7889
rect 33589 7855 33647 7889
rect 33681 7855 33739 7889
rect 33773 7855 33831 7889
rect 33865 7855 33923 7889
rect 33957 7855 34015 7889
rect 34049 7855 34107 7889
rect 34141 7855 34199 7889
rect 34233 7855 34291 7889
rect 34325 7855 34383 7889
rect 34417 7855 34475 7889
rect 34509 7855 34567 7889
rect 34601 7855 34659 7889
rect 34693 7855 34751 7889
rect 34785 7855 34843 7889
rect 34877 7855 34935 7889
rect 34969 7855 35027 7889
rect 35061 7855 35119 7889
rect 35153 7855 35211 7889
rect 35245 7855 35303 7889
rect 35337 7855 35395 7889
rect 35429 7855 35487 7889
rect 35521 7855 35579 7889
rect 35613 7855 35671 7889
rect 35705 7855 35734 7889
rect 35984 7855 36013 7889
rect 36047 7855 36076 7889
rect 30227 7784 30285 7855
rect 30227 7750 30239 7784
rect 30273 7750 30285 7784
rect 30227 7691 30285 7750
rect 30227 7657 30239 7691
rect 30273 7657 30285 7691
rect 30587 7805 30621 7821
rect 30587 7737 30621 7771
rect 30655 7789 30721 7855
rect 30655 7755 30671 7789
rect 30705 7755 30721 7789
rect 30755 7805 30792 7821
rect 30789 7771 30792 7805
rect 30755 7737 30792 7771
rect 30840 7813 30893 7855
rect 30840 7779 30859 7813
rect 30840 7763 30893 7779
rect 30927 7805 30977 7821
rect 30927 7771 30943 7805
rect 31274 7813 31308 7855
rect 30621 7719 30720 7721
rect 30621 7703 30678 7719
rect 30587 7687 30678 7703
rect 30227 7622 30285 7657
rect 30674 7685 30678 7687
rect 30712 7685 30720 7719
rect 30570 7644 30640 7653
rect 30570 7596 30576 7644
rect 30624 7596 30640 7644
rect 30570 7577 30640 7596
rect 30570 7543 30584 7577
rect 30618 7543 30640 7577
rect 30570 7523 30640 7543
rect 30674 7592 30720 7685
rect 30674 7558 30686 7592
rect 30227 7473 30285 7490
rect 30674 7489 30720 7558
rect 30227 7439 30239 7473
rect 30273 7439 30285 7473
rect 30227 7345 30285 7439
rect 30587 7455 30720 7489
rect 30789 7703 30792 7737
rect 30927 7736 30977 7771
rect 31019 7766 31035 7800
rect 31069 7766 31240 7800
rect 30755 7651 30792 7703
rect 30916 7710 30977 7736
rect 31066 7719 31172 7732
rect 30755 7617 30757 7651
rect 30791 7617 30792 7651
rect 30587 7447 30621 7455
rect 30755 7447 30792 7617
rect 30826 7645 30882 7661
rect 30826 7611 30848 7645
rect 30826 7554 30882 7611
rect 30826 7506 30832 7554
rect 30880 7506 30882 7554
rect 30826 7471 30882 7506
rect 30916 7489 30950 7710
rect 31066 7685 31098 7719
rect 31132 7693 31172 7719
rect 30984 7651 31032 7672
rect 30984 7617 30995 7651
rect 31029 7617 31032 7651
rect 30984 7615 31032 7617
rect 30984 7581 30991 7615
rect 31025 7581 31032 7615
rect 30984 7553 31032 7581
rect 31066 7519 31100 7685
rect 31134 7659 31172 7693
rect 31206 7643 31240 7766
rect 31274 7745 31308 7779
rect 31274 7695 31308 7711
rect 31342 7805 31392 7821
rect 31342 7771 31358 7805
rect 31650 7805 31713 7855
rect 31342 7755 31392 7771
rect 31437 7761 31453 7795
rect 31487 7761 31614 7795
rect 31206 7627 31308 7643
rect 31206 7625 31274 7627
rect 30916 7463 30961 7489
rect 30995 7485 31011 7519
rect 31045 7485 31100 7519
rect 30995 7475 31100 7485
rect 31134 7593 31274 7625
rect 31134 7591 31308 7593
rect 30587 7397 30621 7413
rect 30655 7387 30671 7421
rect 30705 7387 30721 7421
rect 30789 7413 30792 7447
rect 30755 7397 30792 7413
rect 30843 7421 30893 7437
rect 30655 7345 30721 7387
rect 30843 7387 30859 7421
rect 30927 7435 30961 7463
rect 31134 7435 31168 7591
rect 31274 7577 31308 7591
rect 31210 7541 31250 7547
rect 31342 7541 31376 7755
rect 31410 7719 31448 7721
rect 31410 7685 31412 7719
rect 31446 7685 31448 7719
rect 31410 7627 31448 7685
rect 31444 7593 31448 7627
rect 31410 7577 31448 7593
rect 31482 7693 31546 7727
rect 31482 7659 31512 7693
rect 31482 7651 31546 7659
rect 31482 7617 31499 7651
rect 31533 7617 31546 7651
rect 31210 7531 31376 7541
rect 31482 7535 31546 7617
rect 31244 7497 31376 7531
rect 31210 7481 31376 7497
rect 30927 7401 30944 7435
rect 30978 7401 30994 7435
rect 31033 7401 31055 7435
rect 31089 7401 31168 7435
rect 31232 7429 31306 7445
rect 30843 7345 30893 7387
rect 31232 7395 31254 7429
rect 31288 7395 31306 7429
rect 31342 7435 31376 7481
rect 31453 7519 31546 7535
rect 31487 7485 31546 7519
rect 31453 7469 31546 7485
rect 31580 7593 31614 7761
rect 31650 7771 31652 7805
rect 31686 7771 31713 7805
rect 31650 7755 31713 7771
rect 31760 7813 31828 7821
rect 31760 7779 31776 7813
rect 31810 7779 31828 7813
rect 31760 7742 31828 7779
rect 31760 7709 31776 7742
rect 31648 7708 31776 7709
rect 31810 7708 31828 7742
rect 31648 7693 31828 7708
rect 31682 7671 31828 7693
rect 31682 7659 31776 7671
rect 31648 7637 31776 7659
rect 31810 7637 31828 7671
rect 31862 7783 31896 7855
rect 32034 7813 32100 7817
rect 31862 7703 31896 7749
rect 31862 7653 31896 7669
rect 31930 7807 31996 7812
rect 31930 7773 31946 7807
rect 31980 7773 31996 7807
rect 31930 7739 31996 7773
rect 31930 7705 31946 7739
rect 31980 7705 31996 7739
rect 31930 7671 31996 7705
rect 32034 7779 32050 7813
rect 32084 7779 32100 7813
rect 32034 7745 32100 7779
rect 32034 7711 32050 7745
rect 32084 7711 32100 7745
rect 32034 7671 32100 7711
rect 31648 7634 31828 7637
rect 31790 7593 31828 7634
rect 31930 7637 31946 7671
rect 31980 7643 31996 7671
rect 31980 7637 32012 7643
rect 31930 7627 32012 7637
rect 31965 7617 32012 7627
rect 31580 7577 31756 7593
rect 31580 7543 31722 7577
rect 31580 7527 31756 7543
rect 31790 7577 31940 7593
rect 31790 7543 31906 7577
rect 31790 7527 31940 7543
rect 31580 7435 31614 7527
rect 31790 7493 31830 7527
rect 31974 7501 32012 7617
rect 31963 7493 32012 7501
rect 31764 7490 31830 7493
rect 31764 7456 31780 7490
rect 31814 7456 31830 7490
rect 31932 7492 32012 7493
rect 31932 7472 31948 7492
rect 31982 7476 32012 7492
rect 32046 7593 32100 7671
rect 32138 7813 32181 7855
rect 32138 7779 32147 7813
rect 32138 7745 32181 7779
rect 32138 7711 32147 7745
rect 32138 7677 32181 7711
rect 32138 7643 32147 7677
rect 32138 7627 32181 7643
rect 32215 7813 32282 7821
rect 32215 7779 32231 7813
rect 32265 7779 32282 7813
rect 32215 7742 32282 7779
rect 32215 7708 32231 7742
rect 32265 7708 32282 7742
rect 32215 7671 32282 7708
rect 32215 7637 32231 7671
rect 32265 7637 32282 7671
rect 32215 7624 32282 7637
rect 32368 7813 32410 7855
rect 32368 7779 32376 7813
rect 32368 7745 32410 7779
rect 32368 7711 32376 7745
rect 32368 7677 32410 7711
rect 32368 7643 32376 7677
rect 32368 7627 32410 7643
rect 32444 7813 32510 7821
rect 32444 7779 32460 7813
rect 32494 7779 32510 7813
rect 32444 7745 32510 7779
rect 32444 7711 32460 7745
rect 32494 7711 32510 7745
rect 32444 7677 32510 7711
rect 32444 7643 32460 7677
rect 32494 7643 32510 7677
rect 32444 7625 32510 7643
rect 32602 7813 32655 7855
rect 32602 7779 32621 7813
rect 32602 7745 32655 7779
rect 32602 7711 32621 7745
rect 32602 7677 32655 7711
rect 32602 7643 32621 7677
rect 32602 7627 32655 7643
rect 32689 7813 32755 7821
rect 32689 7779 32705 7813
rect 32739 7779 32755 7813
rect 32689 7745 32755 7779
rect 32689 7711 32705 7745
rect 32739 7711 32755 7745
rect 32689 7677 32755 7711
rect 32789 7813 32823 7855
rect 32789 7745 32823 7779
rect 32789 7695 32823 7711
rect 32857 7813 32923 7821
rect 32857 7779 32873 7813
rect 32907 7779 32923 7813
rect 32857 7745 32923 7779
rect 32957 7813 32999 7855
rect 32991 7779 32999 7813
rect 32957 7763 32999 7779
rect 33285 7805 33319 7821
rect 32857 7711 32873 7745
rect 32907 7711 32923 7745
rect 32689 7643 32705 7677
rect 32739 7661 32755 7677
rect 32857 7677 32923 7711
rect 33285 7737 33319 7771
rect 33353 7789 33419 7855
rect 33353 7755 33369 7789
rect 33403 7755 33419 7789
rect 33453 7805 33490 7821
rect 33487 7771 33490 7805
rect 33453 7737 33490 7771
rect 33538 7813 33591 7855
rect 33538 7779 33557 7813
rect 33538 7763 33591 7779
rect 33625 7805 33675 7821
rect 33625 7771 33641 7805
rect 33972 7813 34006 7855
rect 33319 7719 33418 7721
rect 33319 7703 33376 7719
rect 33285 7687 33376 7703
rect 32857 7661 32873 7677
rect 32739 7643 32873 7661
rect 32907 7665 32923 7677
rect 33372 7685 33376 7687
rect 33410 7685 33418 7719
rect 32907 7643 33010 7665
rect 32689 7627 33010 7643
rect 32046 7577 32201 7593
rect 32046 7543 32167 7577
rect 32046 7527 32201 7543
rect 32235 7592 32282 7624
rect 32464 7592 32510 7625
rect 32597 7592 32923 7593
rect 32235 7544 32242 7592
rect 32406 7577 32430 7591
rect 31982 7472 31998 7476
rect 31342 7401 31373 7435
rect 31407 7401 31423 7435
rect 31457 7401 31476 7435
rect 31510 7401 31614 7435
rect 31669 7435 31711 7451
rect 31669 7401 31674 7435
rect 31708 7401 31711 7435
rect 31232 7345 31306 7395
rect 31669 7345 31711 7401
rect 31764 7422 31830 7456
rect 31764 7388 31780 7422
rect 31814 7388 31830 7422
rect 31864 7451 31898 7467
rect 31864 7345 31898 7417
rect 31932 7424 31936 7472
rect 31984 7424 31998 7472
rect 32046 7451 32086 7527
rect 32235 7510 32282 7544
rect 32364 7543 32380 7544
rect 32414 7543 32430 7577
rect 32464 7544 32470 7592
rect 32597 7544 32602 7592
rect 32650 7577 32712 7592
rect 32760 7577 32828 7592
rect 32876 7577 32923 7592
rect 32650 7544 32705 7577
rect 32760 7544 32789 7577
rect 31932 7390 31948 7424
rect 31982 7390 31998 7424
rect 32036 7447 32086 7451
rect 32036 7413 32052 7447
rect 32231 7459 32282 7510
rect 32036 7397 32086 7413
rect 32133 7421 32197 7437
rect 31932 7389 31998 7390
rect 32133 7387 32147 7421
rect 32181 7387 32197 7421
rect 32133 7345 32197 7387
rect 32265 7425 32282 7459
rect 32231 7379 32282 7425
rect 32364 7493 32410 7509
rect 32464 7505 32510 7544
rect 32597 7543 32613 7544
rect 32647 7543 32705 7544
rect 32739 7543 32789 7544
rect 32823 7544 32828 7577
rect 32823 7543 32873 7544
rect 32907 7543 32923 7577
rect 32957 7590 33010 7627
rect 33268 7604 33338 7653
rect 32957 7542 32960 7590
rect 33268 7556 33274 7604
rect 33322 7556 33338 7604
rect 33268 7543 33282 7556
rect 33316 7543 33338 7556
rect 32957 7509 33010 7542
rect 33268 7523 33338 7543
rect 33372 7592 33418 7685
rect 33372 7558 33384 7592
rect 32364 7459 32376 7493
rect 32364 7425 32410 7459
rect 32364 7391 32376 7425
rect 32364 7345 32410 7391
rect 32444 7493 32510 7505
rect 32444 7459 32460 7493
rect 32494 7459 32510 7493
rect 32444 7425 32510 7459
rect 32689 7473 33010 7509
rect 33372 7489 33418 7558
rect 32444 7391 32460 7425
rect 32494 7391 32510 7425
rect 32444 7379 32510 7391
rect 32602 7421 32655 7437
rect 32602 7387 32621 7421
rect 32602 7345 32655 7387
rect 32689 7429 32755 7473
rect 32689 7395 32705 7429
rect 32739 7395 32755 7429
rect 32689 7379 32755 7395
rect 32789 7421 32823 7437
rect 32789 7345 32823 7387
rect 32857 7429 32923 7473
rect 33285 7455 33418 7489
rect 33487 7703 33490 7737
rect 33625 7736 33675 7771
rect 33717 7766 33733 7800
rect 33767 7766 33938 7800
rect 33453 7651 33490 7703
rect 33614 7710 33675 7736
rect 33764 7719 33870 7732
rect 33453 7617 33455 7651
rect 33489 7617 33490 7651
rect 33285 7447 33319 7455
rect 32857 7395 32873 7429
rect 32907 7395 32923 7429
rect 32857 7379 32923 7395
rect 32957 7422 33007 7438
rect 32991 7388 33007 7422
rect 33453 7447 33490 7617
rect 33524 7645 33580 7661
rect 33524 7611 33546 7645
rect 33524 7554 33580 7611
rect 33524 7506 33530 7554
rect 33578 7506 33580 7554
rect 33524 7471 33580 7506
rect 33614 7489 33648 7710
rect 33764 7685 33796 7719
rect 33830 7693 33870 7719
rect 33682 7651 33730 7672
rect 33682 7617 33693 7651
rect 33727 7617 33730 7651
rect 33682 7615 33730 7617
rect 33682 7581 33689 7615
rect 33723 7581 33730 7615
rect 33682 7553 33730 7581
rect 33764 7519 33798 7685
rect 33832 7659 33870 7693
rect 33904 7643 33938 7766
rect 33972 7745 34006 7779
rect 33972 7695 34006 7711
rect 34040 7805 34090 7821
rect 34040 7771 34056 7805
rect 34348 7805 34411 7855
rect 34040 7755 34090 7771
rect 34135 7761 34151 7795
rect 34185 7761 34312 7795
rect 33904 7627 34006 7643
rect 33904 7625 33972 7627
rect 33614 7463 33659 7489
rect 33693 7485 33709 7519
rect 33743 7485 33798 7519
rect 33693 7475 33798 7485
rect 33832 7593 33972 7625
rect 33832 7591 34006 7593
rect 33285 7397 33319 7413
rect 32957 7345 33007 7388
rect 33353 7387 33369 7421
rect 33403 7387 33419 7421
rect 33487 7413 33490 7447
rect 33453 7397 33490 7413
rect 33541 7421 33591 7437
rect 33353 7345 33419 7387
rect 33541 7387 33557 7421
rect 33625 7435 33659 7463
rect 33832 7435 33866 7591
rect 33972 7577 34006 7591
rect 33908 7541 33948 7547
rect 34040 7541 34074 7755
rect 34108 7719 34146 7721
rect 34108 7685 34110 7719
rect 34144 7685 34146 7719
rect 34108 7627 34146 7685
rect 34142 7593 34146 7627
rect 34108 7577 34146 7593
rect 34180 7693 34244 7727
rect 34180 7659 34210 7693
rect 34180 7651 34244 7659
rect 34180 7617 34197 7651
rect 34231 7617 34244 7651
rect 33908 7531 34074 7541
rect 34180 7535 34244 7617
rect 33942 7497 34074 7531
rect 33908 7481 34074 7497
rect 33625 7401 33642 7435
rect 33676 7401 33692 7435
rect 33731 7401 33753 7435
rect 33787 7401 33866 7435
rect 33930 7429 34004 7445
rect 33541 7345 33591 7387
rect 33930 7395 33952 7429
rect 33986 7395 34004 7429
rect 34040 7435 34074 7481
rect 34151 7519 34244 7535
rect 34185 7485 34244 7519
rect 34151 7469 34244 7485
rect 34278 7593 34312 7761
rect 34348 7771 34350 7805
rect 34384 7771 34411 7805
rect 34348 7755 34411 7771
rect 34458 7813 34526 7821
rect 34458 7779 34474 7813
rect 34508 7779 34526 7813
rect 34458 7742 34526 7779
rect 34458 7709 34474 7742
rect 34346 7708 34474 7709
rect 34508 7708 34526 7742
rect 34346 7693 34526 7708
rect 34380 7671 34526 7693
rect 34380 7659 34474 7671
rect 34346 7637 34474 7659
rect 34508 7637 34526 7671
rect 34560 7783 34594 7855
rect 34732 7813 34798 7817
rect 34560 7703 34594 7749
rect 34560 7653 34594 7669
rect 34628 7807 34694 7812
rect 34628 7776 34644 7807
rect 34678 7776 34694 7807
rect 34628 7728 34634 7776
rect 34682 7728 34694 7776
rect 34628 7705 34644 7728
rect 34678 7705 34694 7728
rect 34628 7671 34694 7705
rect 34732 7779 34748 7813
rect 34782 7779 34798 7813
rect 34732 7745 34798 7779
rect 34732 7711 34748 7745
rect 34782 7711 34798 7745
rect 34732 7671 34798 7711
rect 34346 7634 34526 7637
rect 34488 7593 34526 7634
rect 34628 7637 34644 7671
rect 34678 7643 34694 7671
rect 34678 7637 34710 7643
rect 34628 7627 34710 7637
rect 34663 7617 34710 7627
rect 34278 7577 34454 7593
rect 34278 7543 34420 7577
rect 34278 7527 34454 7543
rect 34488 7577 34638 7593
rect 34488 7543 34604 7577
rect 34488 7527 34638 7543
rect 34278 7435 34312 7527
rect 34488 7493 34528 7527
rect 34672 7501 34710 7617
rect 34661 7493 34710 7501
rect 34462 7490 34528 7493
rect 34462 7456 34478 7490
rect 34512 7456 34528 7490
rect 34630 7492 34710 7493
rect 34040 7401 34071 7435
rect 34105 7401 34121 7435
rect 34155 7401 34174 7435
rect 34208 7401 34312 7435
rect 34367 7435 34409 7451
rect 34367 7401 34372 7435
rect 34406 7401 34409 7435
rect 33930 7345 34004 7395
rect 34367 7345 34409 7401
rect 34462 7422 34528 7456
rect 34462 7388 34478 7422
rect 34512 7388 34528 7422
rect 34562 7451 34596 7467
rect 34562 7345 34596 7417
rect 34630 7458 34646 7492
rect 34680 7476 34710 7492
rect 34744 7593 34798 7671
rect 34836 7813 34879 7855
rect 34836 7779 34845 7813
rect 34836 7745 34879 7779
rect 34836 7711 34845 7745
rect 34836 7677 34879 7711
rect 34836 7643 34845 7677
rect 34836 7627 34879 7643
rect 34913 7813 34980 7821
rect 34913 7779 34929 7813
rect 34963 7779 34980 7813
rect 34913 7742 34980 7779
rect 34913 7708 34929 7742
rect 34963 7708 34980 7742
rect 34913 7671 34980 7708
rect 34913 7637 34929 7671
rect 34963 7637 34980 7671
rect 34913 7624 34980 7637
rect 35066 7813 35108 7855
rect 35066 7779 35074 7813
rect 35066 7745 35108 7779
rect 35066 7711 35074 7745
rect 35066 7677 35108 7711
rect 35066 7643 35074 7677
rect 35066 7627 35108 7643
rect 35142 7813 35208 7821
rect 35142 7779 35158 7813
rect 35192 7779 35208 7813
rect 35142 7745 35208 7779
rect 35142 7711 35158 7745
rect 35192 7711 35208 7745
rect 35142 7677 35208 7711
rect 35142 7643 35158 7677
rect 35192 7643 35208 7677
rect 35142 7625 35208 7643
rect 35300 7813 35353 7855
rect 35300 7779 35319 7813
rect 35300 7745 35353 7779
rect 35300 7711 35319 7745
rect 35300 7677 35353 7711
rect 35300 7643 35319 7677
rect 35300 7627 35353 7643
rect 35387 7813 35453 7821
rect 35387 7779 35403 7813
rect 35437 7779 35453 7813
rect 35387 7745 35453 7779
rect 35387 7711 35403 7745
rect 35437 7711 35453 7745
rect 35387 7677 35453 7711
rect 35487 7813 35521 7855
rect 35487 7745 35521 7779
rect 35487 7695 35521 7711
rect 35555 7813 35621 7821
rect 35555 7779 35571 7813
rect 35605 7779 35621 7813
rect 35555 7745 35621 7779
rect 35655 7813 35697 7855
rect 35689 7779 35697 7813
rect 35655 7763 35697 7779
rect 36001 7784 36059 7855
rect 35555 7711 35571 7745
rect 35605 7711 35621 7745
rect 35387 7643 35403 7677
rect 35437 7661 35453 7677
rect 35555 7677 35621 7711
rect 35555 7661 35571 7677
rect 35437 7643 35571 7661
rect 35605 7665 35621 7677
rect 36001 7750 36013 7784
rect 36047 7750 36059 7784
rect 36001 7691 36059 7750
rect 35605 7643 35708 7665
rect 35387 7627 35708 7643
rect 34744 7577 34899 7593
rect 34744 7543 34865 7577
rect 34744 7527 34899 7543
rect 34933 7592 34980 7624
rect 35162 7592 35208 7625
rect 35295 7592 35621 7593
rect 34933 7544 34940 7592
rect 35104 7577 35128 7591
rect 34680 7458 34696 7476
rect 34630 7424 34696 7458
rect 34744 7451 34784 7527
rect 34933 7510 34980 7544
rect 35062 7543 35078 7544
rect 35112 7543 35128 7577
rect 35162 7544 35168 7592
rect 35295 7544 35300 7592
rect 35348 7577 35410 7592
rect 35458 7577 35526 7592
rect 35574 7577 35621 7592
rect 35348 7544 35403 7577
rect 35458 7544 35487 7577
rect 34630 7390 34646 7424
rect 34680 7390 34696 7424
rect 34734 7447 34784 7451
rect 34734 7413 34750 7447
rect 34929 7459 34980 7510
rect 34734 7397 34784 7413
rect 34831 7421 34895 7437
rect 34630 7389 34696 7390
rect 34831 7387 34845 7421
rect 34879 7387 34895 7421
rect 34831 7345 34895 7387
rect 34963 7425 34980 7459
rect 34929 7379 34980 7425
rect 35062 7493 35108 7509
rect 35162 7505 35208 7544
rect 35295 7543 35311 7544
rect 35345 7543 35403 7544
rect 35437 7543 35487 7544
rect 35521 7544 35526 7577
rect 35521 7543 35571 7544
rect 35605 7543 35621 7577
rect 35655 7590 35708 7627
rect 36001 7657 36013 7691
rect 36047 7657 36059 7691
rect 36001 7622 36059 7657
rect 35655 7542 35658 7590
rect 35706 7542 35708 7590
rect 35655 7509 35708 7542
rect 35062 7459 35074 7493
rect 35062 7425 35108 7459
rect 35062 7391 35074 7425
rect 35062 7345 35108 7391
rect 35142 7493 35208 7505
rect 35142 7459 35158 7493
rect 35192 7459 35208 7493
rect 35142 7425 35208 7459
rect 35387 7473 35708 7509
rect 36001 7473 36059 7490
rect 35142 7391 35158 7425
rect 35192 7391 35208 7425
rect 35142 7379 35208 7391
rect 35300 7421 35353 7437
rect 35300 7387 35319 7421
rect 35300 7345 35353 7387
rect 35387 7429 35453 7473
rect 35387 7395 35403 7429
rect 35437 7395 35453 7429
rect 35387 7379 35453 7395
rect 35487 7421 35521 7437
rect 35487 7345 35521 7387
rect 35555 7429 35621 7473
rect 36001 7439 36013 7473
rect 36047 7439 36059 7473
rect 35555 7395 35571 7429
rect 35605 7395 35621 7429
rect 35555 7379 35621 7395
rect 35655 7422 35705 7438
rect 35689 7388 35705 7422
rect 35655 7345 35705 7388
rect 36001 7345 36059 7439
rect 30210 7311 30239 7345
rect 30273 7311 30302 7345
rect 30552 7311 30581 7345
rect 30615 7311 30673 7345
rect 30707 7311 30765 7345
rect 30799 7311 30857 7345
rect 30891 7311 30949 7345
rect 30983 7311 31041 7345
rect 31075 7311 31133 7345
rect 31167 7311 31225 7345
rect 31259 7311 31317 7345
rect 31351 7311 31409 7345
rect 31443 7311 31501 7345
rect 31535 7311 31593 7345
rect 31627 7311 31685 7345
rect 31719 7311 31777 7345
rect 31811 7311 31869 7345
rect 31903 7311 31961 7345
rect 31995 7311 32053 7345
rect 32087 7311 32145 7345
rect 32179 7311 32237 7345
rect 32271 7311 32329 7345
rect 32363 7311 32421 7345
rect 32455 7311 32513 7345
rect 32547 7311 32605 7345
rect 32639 7311 32697 7345
rect 32731 7311 32789 7345
rect 32823 7311 32881 7345
rect 32915 7311 32973 7345
rect 33007 7311 33036 7345
rect 33250 7311 33279 7345
rect 33313 7311 33371 7345
rect 33405 7311 33463 7345
rect 33497 7311 33555 7345
rect 33589 7311 33647 7345
rect 33681 7311 33739 7345
rect 33773 7311 33831 7345
rect 33865 7311 33923 7345
rect 33957 7311 34015 7345
rect 34049 7311 34107 7345
rect 34141 7311 34199 7345
rect 34233 7311 34291 7345
rect 34325 7311 34383 7345
rect 34417 7311 34475 7345
rect 34509 7311 34567 7345
rect 34601 7311 34659 7345
rect 34693 7311 34751 7345
rect 34785 7311 34843 7345
rect 34877 7311 34935 7345
rect 34969 7311 35027 7345
rect 35061 7311 35119 7345
rect 35153 7311 35211 7345
rect 35245 7311 35303 7345
rect 35337 7311 35395 7345
rect 35429 7311 35487 7345
rect 35521 7311 35579 7345
rect 35613 7311 35671 7345
rect 35705 7311 35734 7345
rect 35984 7311 36013 7345
rect 36047 7311 36076 7345
rect 30227 7217 30285 7311
rect 30655 7269 30721 7311
rect 30227 7183 30239 7217
rect 30273 7183 30285 7217
rect 30227 7166 30285 7183
rect 30587 7243 30621 7259
rect 30655 7235 30671 7269
rect 30705 7235 30721 7269
rect 30843 7269 30893 7311
rect 30755 7243 30792 7259
rect 30587 7201 30621 7209
rect 30789 7209 30792 7243
rect 30843 7235 30859 7269
rect 31232 7261 31306 7311
rect 30843 7219 30893 7235
rect 30927 7221 30944 7255
rect 30978 7221 30994 7255
rect 31033 7221 31055 7255
rect 31089 7221 31168 7255
rect 30587 7167 30720 7201
rect 30570 7113 30640 7133
rect 30570 7100 30584 7113
rect 30618 7100 30640 7113
rect 30570 7052 30576 7100
rect 30624 7052 30640 7100
rect 30227 6999 30285 7034
rect 30570 7003 30640 7052
rect 30674 7098 30720 7167
rect 30674 7064 30686 7098
rect 30227 6965 30239 6999
rect 30273 6965 30285 6999
rect 30674 6971 30720 7064
rect 30674 6969 30678 6971
rect 30227 6906 30285 6965
rect 30227 6872 30239 6906
rect 30273 6872 30285 6906
rect 30227 6801 30285 6872
rect 30587 6953 30678 6969
rect 30621 6937 30678 6953
rect 30712 6937 30720 6971
rect 30621 6935 30720 6937
rect 30755 7039 30792 7209
rect 30927 7193 30961 7221
rect 30755 7005 30757 7039
rect 30791 7005 30792 7039
rect 30755 6953 30792 7005
rect 30826 7150 30882 7185
rect 30826 7102 30832 7150
rect 30880 7102 30882 7150
rect 30826 7045 30882 7102
rect 30826 7011 30848 7045
rect 30826 6995 30882 7011
rect 30916 7167 30961 7193
rect 30995 7171 31100 7181
rect 30587 6885 30621 6919
rect 30789 6919 30792 6953
rect 30916 6946 30950 7167
rect 30995 7137 31011 7171
rect 31045 7137 31100 7171
rect 30984 7075 31032 7103
rect 30984 7041 30991 7075
rect 31025 7041 31032 7075
rect 30984 7039 31032 7041
rect 30984 7005 30995 7039
rect 31029 7005 31032 7039
rect 30984 6984 31032 7005
rect 31066 6971 31100 7137
rect 31134 7065 31168 7221
rect 31232 7227 31254 7261
rect 31288 7227 31306 7261
rect 31669 7255 31711 7311
rect 31232 7211 31306 7227
rect 31342 7221 31373 7255
rect 31407 7221 31423 7255
rect 31457 7221 31476 7255
rect 31510 7221 31614 7255
rect 31342 7175 31376 7221
rect 31210 7159 31376 7175
rect 31244 7125 31376 7159
rect 31210 7115 31376 7125
rect 31453 7171 31546 7187
rect 31487 7137 31546 7171
rect 31453 7121 31546 7137
rect 31210 7109 31250 7115
rect 31274 7065 31308 7079
rect 31134 7063 31308 7065
rect 31134 7031 31274 7063
rect 31206 7029 31274 7031
rect 31206 7013 31308 7029
rect 30916 6920 30977 6946
rect 31066 6937 31098 6971
rect 31134 6963 31172 6997
rect 31132 6937 31172 6963
rect 31066 6924 31172 6937
rect 30587 6835 30621 6851
rect 30655 6867 30671 6901
rect 30705 6867 30721 6901
rect 30655 6801 30721 6867
rect 30755 6885 30792 6919
rect 30789 6851 30792 6885
rect 30755 6835 30792 6851
rect 30840 6877 30893 6893
rect 30840 6843 30859 6877
rect 30840 6801 30893 6843
rect 30927 6885 30977 6920
rect 31206 6890 31240 7013
rect 30927 6851 30943 6885
rect 31019 6856 31035 6890
rect 31069 6856 31240 6890
rect 31274 6945 31308 6961
rect 31274 6877 31308 6911
rect 30927 6835 30977 6851
rect 31274 6801 31308 6843
rect 31342 6901 31376 7115
rect 31410 7063 31448 7079
rect 31444 7029 31448 7063
rect 31410 6971 31448 7029
rect 31410 6937 31412 6971
rect 31446 6937 31448 6971
rect 31410 6935 31448 6937
rect 31482 7039 31546 7121
rect 31482 7005 31499 7039
rect 31533 7005 31546 7039
rect 31482 6997 31546 7005
rect 31482 6963 31512 6997
rect 31482 6929 31546 6963
rect 31580 7129 31614 7221
rect 31669 7221 31674 7255
rect 31708 7221 31711 7255
rect 31669 7205 31711 7221
rect 31764 7234 31780 7268
rect 31814 7234 31830 7268
rect 31764 7200 31830 7234
rect 31764 7166 31780 7200
rect 31814 7166 31830 7200
rect 31864 7239 31898 7311
rect 32133 7269 32197 7311
rect 31864 7189 31898 7205
rect 31932 7266 31998 7267
rect 31932 7232 31948 7266
rect 31982 7232 31998 7266
rect 31932 7198 31998 7232
rect 32036 7243 32086 7259
rect 32036 7209 32052 7243
rect 32133 7235 32147 7269
rect 32181 7235 32197 7269
rect 32133 7219 32197 7235
rect 32231 7231 32282 7277
rect 32036 7205 32086 7209
rect 31764 7163 31830 7166
rect 31932 7164 31948 7198
rect 31982 7180 31998 7198
rect 31982 7164 32012 7180
rect 31932 7163 32012 7164
rect 31790 7129 31830 7163
rect 31963 7155 32012 7163
rect 31580 7113 31756 7129
rect 31580 7079 31722 7113
rect 31580 7063 31756 7079
rect 31790 7113 31940 7129
rect 31790 7079 31906 7113
rect 31790 7063 31940 7079
rect 31342 6885 31392 6901
rect 31580 6895 31614 7063
rect 31790 7022 31828 7063
rect 31974 7039 32012 7155
rect 31965 7029 32012 7039
rect 31648 7019 31828 7022
rect 31648 6997 31776 7019
rect 31682 6985 31776 6997
rect 31810 6985 31828 7019
rect 31930 7019 32012 7029
rect 31682 6963 31828 6985
rect 31648 6948 31828 6963
rect 31648 6947 31776 6948
rect 31760 6914 31776 6947
rect 31810 6914 31828 6948
rect 31342 6851 31358 6885
rect 31437 6861 31453 6895
rect 31487 6861 31614 6895
rect 31650 6885 31713 6901
rect 31342 6835 31392 6851
rect 31650 6851 31652 6885
rect 31686 6851 31713 6885
rect 31650 6801 31713 6851
rect 31760 6877 31828 6914
rect 31760 6843 31776 6877
rect 31810 6843 31828 6877
rect 31760 6835 31828 6843
rect 31862 6987 31896 7003
rect 31862 6907 31896 6953
rect 31862 6801 31896 6873
rect 31930 6985 31946 7019
rect 31980 7013 32012 7019
rect 32046 7129 32086 7205
rect 32265 7197 32282 7231
rect 32231 7146 32282 7197
rect 32364 7265 32410 7311
rect 32364 7231 32376 7265
rect 32364 7197 32410 7231
rect 32364 7163 32376 7197
rect 32364 7147 32410 7163
rect 32444 7265 32510 7277
rect 32444 7231 32460 7265
rect 32494 7231 32510 7265
rect 32444 7197 32510 7231
rect 32602 7269 32655 7311
rect 32602 7235 32621 7269
rect 32602 7219 32655 7235
rect 32689 7261 32755 7277
rect 32689 7227 32705 7261
rect 32739 7227 32755 7261
rect 32444 7163 32460 7197
rect 32494 7163 32510 7197
rect 32444 7151 32510 7163
rect 32046 7113 32201 7129
rect 32046 7079 32167 7113
rect 32046 7063 32201 7079
rect 32235 7112 32282 7146
rect 32364 7112 32380 7113
rect 32235 7064 32242 7112
rect 32414 7079 32430 7113
rect 32406 7065 32430 7079
rect 32464 7112 32510 7151
rect 32689 7183 32755 7227
rect 32789 7269 32823 7311
rect 32789 7219 32823 7235
rect 32857 7261 32923 7277
rect 32857 7227 32873 7261
rect 32907 7227 32923 7261
rect 32857 7183 32923 7227
rect 32957 7268 33007 7311
rect 32991 7234 33007 7268
rect 33353 7269 33419 7311
rect 32957 7218 33007 7234
rect 33285 7243 33319 7259
rect 33353 7235 33369 7269
rect 33403 7235 33419 7269
rect 33541 7269 33591 7311
rect 33453 7243 33490 7259
rect 33285 7201 33319 7209
rect 33487 7209 33490 7243
rect 33541 7235 33557 7269
rect 33930 7261 34004 7311
rect 33541 7219 33591 7235
rect 33625 7221 33642 7255
rect 33676 7221 33692 7255
rect 33731 7221 33753 7255
rect 33787 7221 33866 7255
rect 32689 7147 33010 7183
rect 33285 7167 33418 7201
rect 32957 7114 33010 7147
rect 32597 7112 32613 7113
rect 32647 7112 32705 7113
rect 32739 7112 32789 7113
rect 32464 7064 32470 7112
rect 32597 7064 32602 7112
rect 32650 7079 32705 7112
rect 32760 7079 32789 7112
rect 32823 7112 32873 7113
rect 32823 7079 32828 7112
rect 32907 7079 32923 7113
rect 32650 7064 32712 7079
rect 32760 7064 32828 7079
rect 32876 7064 32923 7079
rect 31980 6985 31996 7013
rect 32046 6985 32100 7063
rect 32235 7032 32282 7064
rect 31930 6951 31996 6985
rect 31930 6928 31946 6951
rect 31980 6928 31996 6951
rect 31930 6880 31936 6928
rect 31984 6880 31996 6928
rect 31930 6849 31946 6880
rect 31980 6849 31996 6880
rect 31930 6844 31996 6849
rect 32034 6945 32100 6985
rect 32034 6911 32050 6945
rect 32084 6911 32100 6945
rect 32034 6877 32100 6911
rect 32034 6843 32050 6877
rect 32084 6843 32100 6877
rect 32034 6839 32100 6843
rect 32138 7013 32181 7029
rect 32138 6979 32147 7013
rect 32138 6945 32181 6979
rect 32138 6911 32147 6945
rect 32138 6877 32181 6911
rect 32138 6843 32147 6877
rect 32138 6801 32181 6843
rect 32215 7019 32282 7032
rect 32464 7031 32510 7064
rect 32597 7063 32923 7064
rect 32957 7066 32960 7114
rect 33008 7066 33010 7114
rect 32215 6985 32231 7019
rect 32265 6985 32282 7019
rect 32215 6948 32282 6985
rect 32215 6914 32231 6948
rect 32265 6914 32282 6948
rect 32215 6877 32282 6914
rect 32215 6843 32231 6877
rect 32265 6843 32282 6877
rect 32215 6835 32282 6843
rect 32368 7013 32410 7029
rect 32368 6979 32376 7013
rect 32368 6945 32410 6979
rect 32368 6911 32376 6945
rect 32368 6877 32410 6911
rect 32368 6843 32376 6877
rect 32368 6801 32410 6843
rect 32444 7013 32510 7031
rect 32957 7029 33010 7066
rect 32444 6979 32460 7013
rect 32494 6979 32510 7013
rect 32444 6945 32510 6979
rect 32444 6911 32460 6945
rect 32494 6911 32510 6945
rect 32444 6877 32510 6911
rect 32444 6843 32460 6877
rect 32494 6843 32510 6877
rect 32444 6835 32510 6843
rect 32602 7013 32655 7029
rect 32602 6979 32621 7013
rect 32602 6945 32655 6979
rect 32602 6911 32621 6945
rect 32602 6877 32655 6911
rect 32602 6843 32621 6877
rect 32602 6801 32655 6843
rect 32689 7013 33010 7029
rect 32689 6979 32705 7013
rect 32739 6995 32873 7013
rect 32739 6979 32755 6995
rect 32689 6945 32755 6979
rect 32857 6979 32873 6995
rect 32907 6991 33010 7013
rect 33268 7113 33338 7133
rect 33268 7079 33282 7113
rect 33316 7079 33338 7113
rect 33268 7060 33338 7079
rect 33268 7012 33274 7060
rect 33322 7012 33338 7060
rect 33268 7003 33338 7012
rect 33372 7098 33418 7167
rect 33372 7064 33384 7098
rect 32907 6979 32923 6991
rect 32689 6911 32705 6945
rect 32739 6911 32755 6945
rect 32689 6877 32755 6911
rect 32689 6843 32705 6877
rect 32739 6843 32755 6877
rect 32689 6835 32755 6843
rect 32789 6945 32823 6961
rect 32789 6877 32823 6911
rect 32789 6801 32823 6843
rect 32857 6945 32923 6979
rect 33372 6971 33418 7064
rect 33372 6969 33376 6971
rect 32857 6911 32873 6945
rect 32907 6911 32923 6945
rect 32857 6877 32923 6911
rect 33285 6953 33376 6969
rect 33319 6937 33376 6953
rect 33410 6937 33418 6971
rect 33319 6935 33418 6937
rect 33453 7039 33490 7209
rect 33625 7193 33659 7221
rect 33453 7005 33455 7039
rect 33489 7005 33490 7039
rect 33453 6953 33490 7005
rect 33524 7150 33580 7185
rect 33524 7102 33530 7150
rect 33578 7102 33580 7150
rect 33524 7045 33580 7102
rect 33524 7011 33546 7045
rect 33524 6995 33580 7011
rect 33614 7167 33659 7193
rect 33693 7171 33798 7181
rect 32857 6843 32873 6877
rect 32907 6843 32923 6877
rect 32857 6835 32923 6843
rect 32957 6877 32999 6893
rect 32991 6843 32999 6877
rect 32957 6801 32999 6843
rect 33285 6885 33319 6919
rect 33487 6919 33490 6953
rect 33614 6946 33648 7167
rect 33693 7137 33709 7171
rect 33743 7137 33798 7171
rect 33682 7075 33730 7103
rect 33682 7041 33689 7075
rect 33723 7041 33730 7075
rect 33682 7039 33730 7041
rect 33682 7005 33693 7039
rect 33727 7005 33730 7039
rect 33682 6984 33730 7005
rect 33764 6971 33798 7137
rect 33832 7065 33866 7221
rect 33930 7227 33952 7261
rect 33986 7227 34004 7261
rect 34367 7255 34409 7311
rect 33930 7211 34004 7227
rect 34040 7221 34071 7255
rect 34105 7221 34121 7255
rect 34155 7221 34174 7255
rect 34208 7221 34312 7255
rect 34040 7175 34074 7221
rect 33908 7159 34074 7175
rect 33942 7125 34074 7159
rect 33908 7115 34074 7125
rect 34151 7171 34244 7187
rect 34185 7137 34244 7171
rect 34151 7121 34244 7137
rect 33908 7109 33948 7115
rect 33972 7065 34006 7079
rect 33832 7063 34006 7065
rect 33832 7031 33972 7063
rect 33904 7029 33972 7031
rect 33904 7013 34006 7029
rect 33614 6920 33675 6946
rect 33764 6937 33796 6971
rect 33832 6963 33870 6997
rect 33830 6937 33870 6963
rect 33764 6924 33870 6937
rect 33285 6835 33319 6851
rect 33353 6867 33369 6901
rect 33403 6867 33419 6901
rect 33353 6801 33419 6867
rect 33453 6885 33490 6919
rect 33487 6851 33490 6885
rect 33453 6835 33490 6851
rect 33538 6877 33591 6893
rect 33538 6843 33557 6877
rect 33538 6801 33591 6843
rect 33625 6885 33675 6920
rect 33904 6890 33938 7013
rect 33625 6851 33641 6885
rect 33717 6856 33733 6890
rect 33767 6856 33938 6890
rect 33972 6945 34006 6961
rect 33972 6877 34006 6911
rect 33625 6835 33675 6851
rect 33972 6801 34006 6843
rect 34040 6901 34074 7115
rect 34108 7063 34146 7079
rect 34142 7029 34146 7063
rect 34108 6971 34146 7029
rect 34108 6937 34110 6971
rect 34144 6937 34146 6971
rect 34108 6935 34146 6937
rect 34180 7039 34244 7121
rect 34180 7005 34197 7039
rect 34231 7005 34244 7039
rect 34180 6997 34244 7005
rect 34180 6963 34210 6997
rect 34180 6929 34244 6963
rect 34278 7129 34312 7221
rect 34367 7221 34372 7255
rect 34406 7221 34409 7255
rect 34367 7205 34409 7221
rect 34462 7234 34478 7268
rect 34512 7234 34528 7268
rect 34462 7200 34528 7234
rect 34462 7166 34478 7200
rect 34512 7166 34528 7200
rect 34562 7239 34596 7311
rect 34831 7269 34895 7311
rect 34562 7189 34596 7205
rect 34630 7266 34696 7267
rect 34630 7232 34646 7266
rect 34680 7232 34696 7266
rect 34462 7163 34528 7166
rect 34630 7184 34634 7232
rect 34682 7184 34696 7232
rect 34734 7243 34784 7259
rect 34734 7209 34750 7243
rect 34831 7235 34845 7269
rect 34879 7235 34895 7269
rect 34831 7219 34895 7235
rect 34929 7231 34980 7277
rect 34734 7205 34784 7209
rect 34630 7164 34646 7184
rect 34680 7180 34696 7184
rect 34680 7164 34710 7180
rect 34630 7163 34710 7164
rect 34488 7129 34528 7163
rect 34661 7155 34710 7163
rect 34278 7113 34454 7129
rect 34278 7079 34420 7113
rect 34278 7063 34454 7079
rect 34488 7113 34638 7129
rect 34488 7079 34604 7113
rect 34488 7063 34638 7079
rect 34040 6885 34090 6901
rect 34278 6895 34312 7063
rect 34488 7022 34526 7063
rect 34672 7039 34710 7155
rect 34663 7029 34710 7039
rect 34346 7019 34526 7022
rect 34346 6997 34474 7019
rect 34380 6985 34474 6997
rect 34508 6985 34526 7019
rect 34628 7019 34710 7029
rect 34380 6963 34526 6985
rect 34346 6948 34526 6963
rect 34346 6947 34474 6948
rect 34458 6914 34474 6947
rect 34508 6914 34526 6948
rect 34040 6851 34056 6885
rect 34135 6861 34151 6895
rect 34185 6861 34312 6895
rect 34348 6885 34411 6901
rect 34040 6835 34090 6851
rect 34348 6851 34350 6885
rect 34384 6851 34411 6885
rect 34348 6801 34411 6851
rect 34458 6877 34526 6914
rect 34458 6843 34474 6877
rect 34508 6843 34526 6877
rect 34458 6835 34526 6843
rect 34560 6987 34594 7003
rect 34560 6907 34594 6953
rect 34560 6801 34594 6873
rect 34628 6985 34644 7019
rect 34678 7013 34710 7019
rect 34744 7129 34784 7205
rect 34963 7197 34980 7231
rect 34929 7146 34980 7197
rect 35062 7265 35108 7311
rect 35062 7231 35074 7265
rect 35062 7197 35108 7231
rect 35062 7163 35074 7197
rect 35062 7147 35108 7163
rect 35142 7265 35208 7277
rect 35142 7231 35158 7265
rect 35192 7231 35208 7265
rect 35142 7197 35208 7231
rect 35300 7269 35353 7311
rect 35300 7235 35319 7269
rect 35300 7219 35353 7235
rect 35387 7261 35453 7277
rect 35387 7227 35403 7261
rect 35437 7227 35453 7261
rect 35142 7163 35158 7197
rect 35192 7163 35208 7197
rect 35142 7151 35208 7163
rect 34744 7113 34899 7129
rect 34744 7079 34865 7113
rect 34744 7063 34899 7079
rect 34933 7112 34980 7146
rect 35062 7112 35078 7113
rect 34933 7064 34940 7112
rect 35112 7079 35128 7113
rect 35104 7065 35128 7079
rect 35162 7112 35208 7151
rect 35387 7183 35453 7227
rect 35487 7269 35521 7311
rect 35487 7219 35521 7235
rect 35555 7261 35621 7277
rect 35555 7227 35571 7261
rect 35605 7227 35621 7261
rect 35555 7183 35621 7227
rect 35655 7268 35705 7311
rect 35689 7234 35705 7268
rect 35655 7218 35705 7234
rect 36001 7217 36059 7311
rect 36001 7183 36013 7217
rect 36047 7183 36059 7217
rect 35387 7147 35708 7183
rect 36001 7166 36059 7183
rect 35655 7114 35708 7147
rect 35295 7112 35311 7113
rect 35345 7112 35403 7113
rect 35437 7112 35487 7113
rect 35162 7064 35168 7112
rect 35295 7064 35300 7112
rect 35348 7079 35403 7112
rect 35458 7079 35487 7112
rect 35521 7112 35571 7113
rect 35521 7079 35526 7112
rect 35605 7079 35621 7113
rect 35348 7064 35410 7079
rect 35458 7064 35526 7079
rect 35574 7064 35621 7079
rect 34678 6985 34694 7013
rect 34744 6985 34798 7063
rect 34933 7032 34980 7064
rect 34628 6951 34694 6985
rect 34628 6917 34644 6951
rect 34678 6917 34694 6951
rect 34628 6883 34694 6917
rect 34628 6849 34644 6883
rect 34678 6849 34694 6883
rect 34628 6844 34694 6849
rect 34732 6945 34798 6985
rect 34732 6911 34748 6945
rect 34782 6911 34798 6945
rect 34732 6877 34798 6911
rect 34732 6843 34748 6877
rect 34782 6843 34798 6877
rect 34732 6839 34798 6843
rect 34836 7013 34879 7029
rect 34836 6979 34845 7013
rect 34836 6945 34879 6979
rect 34836 6911 34845 6945
rect 34836 6877 34879 6911
rect 34836 6843 34845 6877
rect 34836 6801 34879 6843
rect 34913 7019 34980 7032
rect 35162 7031 35208 7064
rect 35295 7063 35621 7064
rect 35655 7066 35658 7114
rect 34913 6985 34929 7019
rect 34963 6985 34980 7019
rect 34913 6948 34980 6985
rect 34913 6914 34929 6948
rect 34963 6914 34980 6948
rect 34913 6877 34980 6914
rect 34913 6843 34929 6877
rect 34963 6843 34980 6877
rect 34913 6835 34980 6843
rect 35066 7013 35108 7029
rect 35066 6979 35074 7013
rect 35066 6945 35108 6979
rect 35066 6911 35074 6945
rect 35066 6877 35108 6911
rect 35066 6843 35074 6877
rect 35066 6801 35108 6843
rect 35142 7013 35208 7031
rect 35655 7029 35708 7066
rect 35142 6979 35158 7013
rect 35192 6979 35208 7013
rect 35142 6945 35208 6979
rect 35142 6911 35158 6945
rect 35192 6911 35208 6945
rect 35142 6877 35208 6911
rect 35142 6843 35158 6877
rect 35192 6843 35208 6877
rect 35142 6835 35208 6843
rect 35300 7013 35353 7029
rect 35300 6979 35319 7013
rect 35300 6945 35353 6979
rect 35300 6911 35319 6945
rect 35300 6877 35353 6911
rect 35300 6843 35319 6877
rect 35300 6801 35353 6843
rect 35387 7013 35708 7029
rect 35387 6979 35403 7013
rect 35437 6995 35571 7013
rect 35437 6979 35453 6995
rect 35387 6945 35453 6979
rect 35555 6979 35571 6995
rect 35605 6991 35708 7013
rect 36001 6999 36059 7034
rect 35605 6979 35621 6991
rect 35387 6911 35403 6945
rect 35437 6911 35453 6945
rect 35387 6877 35453 6911
rect 35387 6843 35403 6877
rect 35437 6843 35453 6877
rect 35387 6835 35453 6843
rect 35487 6945 35521 6961
rect 35487 6877 35521 6911
rect 35487 6801 35521 6843
rect 35555 6945 35621 6979
rect 35555 6911 35571 6945
rect 35605 6911 35621 6945
rect 35555 6877 35621 6911
rect 36001 6965 36013 6999
rect 36047 6965 36059 6999
rect 36001 6906 36059 6965
rect 35555 6843 35571 6877
rect 35605 6843 35621 6877
rect 35555 6835 35621 6843
rect 35655 6877 35697 6893
rect 35689 6843 35697 6877
rect 35655 6801 35697 6843
rect 36001 6872 36013 6906
rect 36047 6872 36059 6906
rect 36001 6801 36059 6872
rect 30210 6767 30239 6801
rect 30273 6767 30302 6801
rect 30552 6767 30581 6801
rect 30615 6767 30673 6801
rect 30707 6767 30765 6801
rect 30799 6767 30857 6801
rect 30891 6767 30949 6801
rect 30983 6767 31041 6801
rect 31075 6767 31133 6801
rect 31167 6767 31225 6801
rect 31259 6767 31317 6801
rect 31351 6767 31409 6801
rect 31443 6767 31501 6801
rect 31535 6767 31593 6801
rect 31627 6767 31685 6801
rect 31719 6767 31777 6801
rect 31811 6767 31869 6801
rect 31903 6767 31961 6801
rect 31995 6767 32053 6801
rect 32087 6767 32145 6801
rect 32179 6767 32237 6801
rect 32271 6767 32329 6801
rect 32363 6767 32421 6801
rect 32455 6767 32513 6801
rect 32547 6767 32605 6801
rect 32639 6767 32697 6801
rect 32731 6767 32789 6801
rect 32823 6767 32881 6801
rect 32915 6767 32973 6801
rect 33007 6767 33036 6801
rect 33250 6767 33279 6801
rect 33313 6767 33371 6801
rect 33405 6767 33463 6801
rect 33497 6767 33555 6801
rect 33589 6767 33647 6801
rect 33681 6767 33739 6801
rect 33773 6767 33831 6801
rect 33865 6767 33923 6801
rect 33957 6767 34015 6801
rect 34049 6767 34107 6801
rect 34141 6767 34199 6801
rect 34233 6767 34291 6801
rect 34325 6767 34383 6801
rect 34417 6767 34475 6801
rect 34509 6767 34567 6801
rect 34601 6767 34659 6801
rect 34693 6767 34751 6801
rect 34785 6767 34843 6801
rect 34877 6767 34935 6801
rect 34969 6767 35027 6801
rect 35061 6767 35119 6801
rect 35153 6767 35211 6801
rect 35245 6767 35303 6801
rect 35337 6767 35395 6801
rect 35429 6767 35487 6801
rect 35521 6767 35579 6801
rect 35613 6767 35671 6801
rect 35705 6767 35734 6801
rect 35984 6767 36013 6801
rect 36047 6767 36076 6801
rect 30227 6696 30285 6767
rect 30227 6662 30239 6696
rect 30273 6662 30285 6696
rect 30227 6603 30285 6662
rect 30227 6569 30239 6603
rect 30273 6569 30285 6603
rect 30587 6717 30621 6733
rect 30587 6649 30621 6683
rect 30655 6701 30721 6767
rect 30655 6667 30671 6701
rect 30705 6667 30721 6701
rect 30755 6717 30792 6733
rect 30789 6683 30792 6717
rect 30755 6649 30792 6683
rect 30840 6725 30893 6767
rect 30840 6691 30859 6725
rect 30840 6675 30893 6691
rect 30927 6717 30977 6733
rect 30927 6683 30943 6717
rect 31274 6725 31308 6767
rect 30621 6631 30720 6633
rect 30621 6615 30678 6631
rect 30587 6599 30678 6615
rect 30227 6534 30285 6569
rect 30674 6597 30678 6599
rect 30712 6597 30720 6631
rect 30570 6556 30640 6565
rect 30570 6508 30576 6556
rect 30624 6508 30640 6556
rect 30570 6489 30640 6508
rect 30570 6455 30584 6489
rect 30618 6455 30640 6489
rect 30570 6435 30640 6455
rect 30674 6504 30720 6597
rect 30674 6470 30686 6504
rect 30227 6385 30285 6402
rect 30674 6401 30720 6470
rect 30227 6351 30239 6385
rect 30273 6351 30285 6385
rect 30227 6257 30285 6351
rect 30587 6367 30720 6401
rect 30789 6615 30792 6649
rect 30927 6648 30977 6683
rect 31019 6678 31035 6712
rect 31069 6678 31240 6712
rect 30755 6563 30792 6615
rect 30916 6622 30977 6648
rect 31066 6631 31172 6644
rect 30755 6529 30757 6563
rect 30791 6529 30792 6563
rect 30587 6359 30621 6367
rect 30755 6359 30792 6529
rect 30826 6557 30882 6573
rect 30826 6523 30848 6557
rect 30826 6466 30882 6523
rect 30826 6418 30832 6466
rect 30880 6418 30882 6466
rect 30826 6383 30882 6418
rect 30916 6401 30950 6622
rect 31066 6597 31098 6631
rect 31132 6605 31172 6631
rect 30984 6563 31032 6584
rect 30984 6529 30995 6563
rect 31029 6529 31032 6563
rect 30984 6527 31032 6529
rect 30984 6493 30991 6527
rect 31025 6493 31032 6527
rect 30984 6465 31032 6493
rect 31066 6431 31100 6597
rect 31134 6571 31172 6605
rect 31206 6555 31240 6678
rect 31274 6657 31308 6691
rect 31274 6607 31308 6623
rect 31342 6717 31392 6733
rect 31342 6683 31358 6717
rect 31650 6717 31713 6767
rect 31342 6667 31392 6683
rect 31437 6673 31453 6707
rect 31487 6673 31614 6707
rect 31206 6539 31308 6555
rect 31206 6537 31274 6539
rect 30916 6375 30961 6401
rect 30995 6397 31011 6431
rect 31045 6397 31100 6431
rect 30995 6387 31100 6397
rect 31134 6505 31274 6537
rect 31134 6503 31308 6505
rect 30587 6309 30621 6325
rect 30655 6299 30671 6333
rect 30705 6299 30721 6333
rect 30789 6325 30792 6359
rect 30755 6309 30792 6325
rect 30843 6333 30893 6349
rect 30655 6257 30721 6299
rect 30843 6299 30859 6333
rect 30927 6347 30961 6375
rect 31134 6347 31168 6503
rect 31274 6489 31308 6503
rect 31210 6453 31250 6459
rect 31342 6453 31376 6667
rect 31410 6631 31448 6633
rect 31410 6597 31412 6631
rect 31446 6597 31448 6631
rect 31410 6539 31448 6597
rect 31444 6505 31448 6539
rect 31410 6489 31448 6505
rect 31482 6605 31546 6639
rect 31482 6571 31512 6605
rect 31482 6563 31546 6571
rect 31482 6529 31499 6563
rect 31533 6529 31546 6563
rect 31210 6443 31376 6453
rect 31482 6447 31546 6529
rect 31244 6409 31376 6443
rect 31210 6393 31376 6409
rect 30927 6313 30944 6347
rect 30978 6313 30994 6347
rect 31033 6313 31055 6347
rect 31089 6313 31168 6347
rect 31232 6341 31306 6357
rect 30843 6257 30893 6299
rect 31232 6307 31254 6341
rect 31288 6307 31306 6341
rect 31342 6347 31376 6393
rect 31453 6431 31546 6447
rect 31487 6397 31546 6431
rect 31453 6381 31546 6397
rect 31580 6505 31614 6673
rect 31650 6683 31652 6717
rect 31686 6683 31713 6717
rect 31650 6667 31713 6683
rect 31760 6725 31828 6733
rect 31760 6691 31776 6725
rect 31810 6691 31828 6725
rect 31760 6654 31828 6691
rect 31760 6621 31776 6654
rect 31648 6620 31776 6621
rect 31810 6620 31828 6654
rect 31648 6605 31828 6620
rect 31682 6583 31828 6605
rect 31682 6571 31776 6583
rect 31648 6549 31776 6571
rect 31810 6549 31828 6583
rect 31862 6695 31896 6767
rect 32034 6725 32100 6729
rect 31862 6615 31896 6661
rect 31862 6565 31896 6581
rect 31930 6719 31996 6724
rect 31930 6685 31946 6719
rect 31980 6685 31996 6719
rect 31930 6651 31996 6685
rect 31930 6617 31946 6651
rect 31980 6617 31996 6651
rect 31930 6583 31996 6617
rect 32034 6691 32050 6725
rect 32084 6691 32100 6725
rect 32034 6657 32100 6691
rect 32034 6623 32050 6657
rect 32084 6623 32100 6657
rect 32034 6583 32100 6623
rect 31648 6546 31828 6549
rect 31790 6505 31828 6546
rect 31930 6549 31946 6583
rect 31980 6555 31996 6583
rect 31980 6549 32012 6555
rect 31930 6539 32012 6549
rect 31965 6529 32012 6539
rect 31580 6489 31756 6505
rect 31580 6455 31722 6489
rect 31580 6439 31756 6455
rect 31790 6489 31940 6505
rect 31790 6455 31906 6489
rect 31790 6439 31940 6455
rect 31580 6347 31614 6439
rect 31790 6405 31830 6439
rect 31974 6413 32012 6529
rect 31963 6405 32012 6413
rect 31764 6402 31830 6405
rect 31764 6368 31780 6402
rect 31814 6368 31830 6402
rect 31932 6404 32012 6405
rect 31932 6386 31948 6404
rect 31982 6388 32012 6404
rect 32046 6505 32100 6583
rect 32138 6725 32181 6767
rect 32138 6691 32147 6725
rect 32138 6657 32181 6691
rect 32138 6623 32147 6657
rect 32138 6589 32181 6623
rect 32138 6555 32147 6589
rect 32138 6539 32181 6555
rect 32215 6725 32282 6733
rect 32215 6691 32231 6725
rect 32265 6691 32282 6725
rect 32215 6654 32282 6691
rect 32215 6620 32231 6654
rect 32265 6620 32282 6654
rect 32215 6583 32282 6620
rect 32215 6549 32231 6583
rect 32265 6549 32282 6583
rect 32215 6536 32282 6549
rect 32368 6725 32410 6767
rect 32368 6691 32376 6725
rect 32368 6657 32410 6691
rect 32368 6623 32376 6657
rect 32368 6589 32410 6623
rect 32368 6555 32376 6589
rect 32368 6539 32410 6555
rect 32444 6725 32510 6733
rect 32444 6691 32460 6725
rect 32494 6691 32510 6725
rect 32444 6657 32510 6691
rect 32444 6623 32460 6657
rect 32494 6623 32510 6657
rect 32444 6589 32510 6623
rect 32444 6555 32460 6589
rect 32494 6555 32510 6589
rect 32444 6537 32510 6555
rect 32602 6725 32655 6767
rect 32602 6691 32621 6725
rect 32602 6657 32655 6691
rect 32602 6623 32621 6657
rect 32602 6589 32655 6623
rect 32602 6555 32621 6589
rect 32602 6539 32655 6555
rect 32689 6725 32755 6733
rect 32689 6691 32705 6725
rect 32739 6691 32755 6725
rect 32689 6657 32755 6691
rect 32689 6623 32705 6657
rect 32739 6623 32755 6657
rect 32689 6589 32755 6623
rect 32789 6725 32823 6767
rect 32789 6657 32823 6691
rect 32789 6607 32823 6623
rect 32857 6725 32923 6733
rect 32857 6691 32873 6725
rect 32907 6691 32923 6725
rect 32857 6657 32923 6691
rect 32957 6725 32999 6767
rect 32991 6691 32999 6725
rect 32957 6675 32999 6691
rect 33285 6717 33319 6733
rect 32857 6623 32873 6657
rect 32907 6623 32923 6657
rect 32689 6555 32705 6589
rect 32739 6573 32755 6589
rect 32857 6589 32923 6623
rect 33285 6649 33319 6683
rect 33353 6701 33419 6767
rect 33353 6667 33369 6701
rect 33403 6667 33419 6701
rect 33453 6717 33490 6733
rect 33487 6683 33490 6717
rect 33453 6649 33490 6683
rect 33538 6725 33591 6767
rect 33538 6691 33557 6725
rect 33538 6675 33591 6691
rect 33625 6717 33675 6733
rect 33625 6683 33641 6717
rect 33972 6725 34006 6767
rect 33319 6631 33418 6633
rect 33319 6615 33376 6631
rect 33285 6599 33376 6615
rect 32857 6573 32873 6589
rect 32739 6555 32873 6573
rect 32907 6577 32923 6589
rect 33372 6597 33376 6599
rect 33410 6597 33418 6631
rect 32907 6555 33010 6577
rect 32689 6539 33010 6555
rect 32046 6489 32201 6505
rect 32046 6455 32167 6489
rect 32046 6439 32201 6455
rect 32235 6504 32282 6536
rect 32464 6504 32510 6537
rect 32597 6504 32923 6505
rect 32235 6456 32242 6504
rect 32406 6489 32430 6503
rect 31982 6386 31998 6388
rect 31342 6313 31373 6347
rect 31407 6313 31423 6347
rect 31457 6313 31476 6347
rect 31510 6313 31614 6347
rect 31669 6347 31711 6363
rect 31669 6313 31674 6347
rect 31708 6313 31711 6347
rect 31232 6257 31306 6307
rect 31669 6257 31711 6313
rect 31764 6334 31830 6368
rect 31764 6300 31780 6334
rect 31814 6300 31830 6334
rect 31864 6363 31898 6379
rect 31864 6257 31898 6329
rect 31932 6338 31936 6386
rect 31984 6338 31998 6386
rect 32046 6363 32086 6439
rect 32235 6422 32282 6456
rect 32364 6455 32380 6456
rect 32414 6455 32430 6489
rect 32464 6456 32470 6504
rect 32597 6456 32602 6504
rect 32650 6489 32712 6504
rect 32760 6489 32828 6504
rect 32876 6489 32923 6504
rect 32650 6456 32705 6489
rect 32760 6456 32789 6489
rect 31932 6336 31998 6338
rect 31932 6302 31948 6336
rect 31982 6302 31998 6336
rect 32036 6359 32086 6363
rect 32036 6325 32052 6359
rect 32231 6371 32282 6422
rect 32036 6309 32086 6325
rect 32133 6333 32197 6349
rect 31932 6301 31998 6302
rect 32133 6299 32147 6333
rect 32181 6299 32197 6333
rect 32133 6257 32197 6299
rect 32265 6337 32282 6371
rect 32231 6291 32282 6337
rect 32364 6405 32410 6421
rect 32464 6417 32510 6456
rect 32597 6455 32613 6456
rect 32647 6455 32705 6456
rect 32739 6455 32789 6456
rect 32823 6456 32828 6489
rect 32823 6455 32873 6456
rect 32907 6455 32923 6489
rect 32957 6502 33010 6539
rect 32957 6454 32960 6502
rect 33008 6454 33010 6502
rect 32957 6421 33010 6454
rect 33268 6514 33338 6565
rect 33268 6466 33274 6514
rect 33322 6466 33338 6514
rect 33268 6455 33282 6466
rect 33316 6455 33338 6466
rect 33268 6435 33338 6455
rect 33372 6504 33418 6597
rect 33372 6470 33384 6504
rect 32364 6371 32376 6405
rect 32364 6337 32410 6371
rect 32364 6303 32376 6337
rect 32364 6257 32410 6303
rect 32444 6405 32510 6417
rect 32444 6371 32460 6405
rect 32494 6371 32510 6405
rect 32444 6337 32510 6371
rect 32689 6385 33010 6421
rect 33372 6401 33418 6470
rect 32444 6303 32460 6337
rect 32494 6303 32510 6337
rect 32444 6291 32510 6303
rect 32602 6333 32655 6349
rect 32602 6299 32621 6333
rect 32602 6257 32655 6299
rect 32689 6341 32755 6385
rect 32689 6307 32705 6341
rect 32739 6307 32755 6341
rect 32689 6291 32755 6307
rect 32789 6333 32823 6349
rect 32789 6257 32823 6299
rect 32857 6341 32923 6385
rect 33285 6367 33418 6401
rect 33487 6615 33490 6649
rect 33625 6648 33675 6683
rect 33717 6678 33733 6712
rect 33767 6678 33938 6712
rect 33453 6563 33490 6615
rect 33614 6622 33675 6648
rect 33764 6631 33870 6644
rect 33453 6529 33455 6563
rect 33489 6529 33490 6563
rect 33285 6359 33319 6367
rect 32857 6307 32873 6341
rect 32907 6307 32923 6341
rect 32857 6291 32923 6307
rect 32957 6334 33007 6350
rect 32991 6300 33007 6334
rect 33453 6359 33490 6529
rect 33524 6557 33580 6573
rect 33524 6523 33546 6557
rect 33524 6466 33580 6523
rect 33524 6418 33530 6466
rect 33578 6418 33580 6466
rect 33524 6383 33580 6418
rect 33614 6401 33648 6622
rect 33764 6597 33796 6631
rect 33830 6605 33870 6631
rect 33682 6563 33730 6584
rect 33682 6529 33693 6563
rect 33727 6529 33730 6563
rect 33682 6527 33730 6529
rect 33682 6493 33689 6527
rect 33723 6493 33730 6527
rect 33682 6465 33730 6493
rect 33764 6431 33798 6597
rect 33832 6571 33870 6605
rect 33904 6555 33938 6678
rect 33972 6657 34006 6691
rect 33972 6607 34006 6623
rect 34040 6717 34090 6733
rect 34040 6683 34056 6717
rect 34348 6717 34411 6767
rect 34040 6667 34090 6683
rect 34135 6673 34151 6707
rect 34185 6673 34312 6707
rect 33904 6539 34006 6555
rect 33904 6537 33972 6539
rect 33614 6375 33659 6401
rect 33693 6397 33709 6431
rect 33743 6397 33798 6431
rect 33693 6387 33798 6397
rect 33832 6505 33972 6537
rect 33832 6503 34006 6505
rect 33285 6309 33319 6325
rect 32957 6257 33007 6300
rect 33353 6299 33369 6333
rect 33403 6299 33419 6333
rect 33487 6325 33490 6359
rect 33453 6309 33490 6325
rect 33541 6333 33591 6349
rect 33353 6257 33419 6299
rect 33541 6299 33557 6333
rect 33625 6347 33659 6375
rect 33832 6347 33866 6503
rect 33972 6489 34006 6503
rect 33908 6453 33948 6459
rect 34040 6453 34074 6667
rect 34108 6631 34146 6633
rect 34108 6597 34110 6631
rect 34144 6597 34146 6631
rect 34108 6539 34146 6597
rect 34142 6505 34146 6539
rect 34108 6489 34146 6505
rect 34180 6605 34244 6639
rect 34180 6571 34210 6605
rect 34180 6563 34244 6571
rect 34180 6529 34197 6563
rect 34231 6529 34244 6563
rect 33908 6443 34074 6453
rect 34180 6447 34244 6529
rect 33942 6409 34074 6443
rect 33908 6393 34074 6409
rect 33625 6313 33642 6347
rect 33676 6313 33692 6347
rect 33731 6313 33753 6347
rect 33787 6313 33866 6347
rect 33930 6341 34004 6357
rect 33541 6257 33591 6299
rect 33930 6307 33952 6341
rect 33986 6307 34004 6341
rect 34040 6347 34074 6393
rect 34151 6431 34244 6447
rect 34185 6397 34244 6431
rect 34151 6381 34244 6397
rect 34278 6505 34312 6673
rect 34348 6683 34350 6717
rect 34384 6683 34411 6717
rect 34348 6667 34411 6683
rect 34458 6725 34526 6733
rect 34458 6691 34474 6725
rect 34508 6691 34526 6725
rect 34458 6654 34526 6691
rect 34458 6621 34474 6654
rect 34346 6620 34474 6621
rect 34508 6620 34526 6654
rect 34346 6605 34526 6620
rect 34380 6583 34526 6605
rect 34380 6571 34474 6583
rect 34346 6549 34474 6571
rect 34508 6549 34526 6583
rect 34560 6695 34594 6767
rect 34732 6725 34798 6729
rect 34560 6615 34594 6661
rect 34560 6565 34594 6581
rect 34628 6719 34694 6724
rect 34628 6688 34644 6719
rect 34678 6688 34694 6719
rect 34628 6640 34634 6688
rect 34682 6640 34694 6688
rect 34628 6617 34644 6640
rect 34678 6617 34694 6640
rect 34628 6583 34694 6617
rect 34732 6691 34748 6725
rect 34782 6691 34798 6725
rect 34732 6657 34798 6691
rect 34732 6623 34748 6657
rect 34782 6623 34798 6657
rect 34732 6583 34798 6623
rect 34346 6546 34526 6549
rect 34488 6505 34526 6546
rect 34628 6549 34644 6583
rect 34678 6555 34694 6583
rect 34678 6549 34710 6555
rect 34628 6539 34710 6549
rect 34663 6529 34710 6539
rect 34278 6489 34454 6505
rect 34278 6455 34420 6489
rect 34278 6439 34454 6455
rect 34488 6489 34638 6505
rect 34488 6455 34604 6489
rect 34488 6439 34638 6455
rect 34278 6347 34312 6439
rect 34488 6405 34528 6439
rect 34672 6413 34710 6529
rect 34661 6405 34710 6413
rect 34462 6402 34528 6405
rect 34462 6368 34478 6402
rect 34512 6368 34528 6402
rect 34630 6404 34710 6405
rect 34040 6313 34071 6347
rect 34105 6313 34121 6347
rect 34155 6313 34174 6347
rect 34208 6313 34312 6347
rect 34367 6347 34409 6363
rect 34367 6313 34372 6347
rect 34406 6313 34409 6347
rect 33930 6257 34004 6307
rect 34367 6257 34409 6313
rect 34462 6334 34528 6368
rect 34462 6300 34478 6334
rect 34512 6300 34528 6334
rect 34562 6363 34596 6379
rect 34562 6257 34596 6329
rect 34630 6370 34646 6404
rect 34680 6388 34710 6404
rect 34744 6505 34798 6583
rect 34836 6725 34879 6767
rect 34836 6691 34845 6725
rect 34836 6657 34879 6691
rect 34836 6623 34845 6657
rect 34836 6589 34879 6623
rect 34836 6555 34845 6589
rect 34836 6539 34879 6555
rect 34913 6725 34980 6733
rect 34913 6691 34929 6725
rect 34963 6691 34980 6725
rect 34913 6654 34980 6691
rect 34913 6620 34929 6654
rect 34963 6620 34980 6654
rect 34913 6583 34980 6620
rect 34913 6549 34929 6583
rect 34963 6549 34980 6583
rect 34913 6536 34980 6549
rect 35066 6725 35108 6767
rect 35066 6691 35074 6725
rect 35066 6657 35108 6691
rect 35066 6623 35074 6657
rect 35066 6589 35108 6623
rect 35066 6555 35074 6589
rect 35066 6539 35108 6555
rect 35142 6725 35208 6733
rect 35142 6691 35158 6725
rect 35192 6691 35208 6725
rect 35142 6657 35208 6691
rect 35142 6623 35158 6657
rect 35192 6623 35208 6657
rect 35142 6589 35208 6623
rect 35142 6555 35158 6589
rect 35192 6555 35208 6589
rect 35142 6537 35208 6555
rect 35300 6725 35353 6767
rect 35300 6691 35319 6725
rect 35300 6657 35353 6691
rect 35300 6623 35319 6657
rect 35300 6589 35353 6623
rect 35300 6555 35319 6589
rect 35300 6539 35353 6555
rect 35387 6725 35453 6733
rect 35387 6691 35403 6725
rect 35437 6691 35453 6725
rect 35387 6657 35453 6691
rect 35387 6623 35403 6657
rect 35437 6623 35453 6657
rect 35387 6589 35453 6623
rect 35487 6725 35521 6767
rect 35487 6657 35521 6691
rect 35487 6607 35521 6623
rect 35555 6725 35621 6733
rect 35555 6691 35571 6725
rect 35605 6691 35621 6725
rect 35555 6657 35621 6691
rect 35655 6725 35697 6767
rect 35689 6691 35697 6725
rect 35655 6675 35697 6691
rect 36001 6696 36059 6767
rect 35555 6623 35571 6657
rect 35605 6623 35621 6657
rect 35387 6555 35403 6589
rect 35437 6573 35453 6589
rect 35555 6589 35621 6623
rect 35555 6573 35571 6589
rect 35437 6555 35571 6573
rect 35605 6577 35621 6589
rect 36001 6662 36013 6696
rect 36047 6662 36059 6696
rect 36001 6603 36059 6662
rect 35605 6555 35708 6577
rect 35387 6539 35708 6555
rect 34744 6489 34899 6505
rect 34744 6455 34865 6489
rect 34744 6439 34899 6455
rect 34933 6504 34980 6536
rect 35162 6504 35208 6537
rect 35295 6504 35621 6505
rect 34933 6456 34940 6504
rect 35104 6489 35128 6503
rect 34680 6370 34696 6388
rect 34630 6336 34696 6370
rect 34744 6363 34784 6439
rect 34933 6422 34980 6456
rect 35062 6455 35078 6456
rect 35112 6455 35128 6489
rect 35162 6456 35168 6504
rect 35295 6456 35300 6504
rect 35348 6489 35410 6504
rect 35458 6489 35526 6504
rect 35574 6489 35621 6504
rect 35348 6456 35403 6489
rect 35458 6456 35487 6489
rect 34630 6302 34646 6336
rect 34680 6302 34696 6336
rect 34734 6359 34784 6363
rect 34734 6325 34750 6359
rect 34929 6371 34980 6422
rect 34734 6309 34784 6325
rect 34831 6333 34895 6349
rect 34630 6301 34696 6302
rect 34831 6299 34845 6333
rect 34879 6299 34895 6333
rect 34831 6257 34895 6299
rect 34963 6337 34980 6371
rect 34929 6291 34980 6337
rect 35062 6405 35108 6421
rect 35162 6417 35208 6456
rect 35295 6455 35311 6456
rect 35345 6455 35403 6456
rect 35437 6455 35487 6456
rect 35521 6456 35526 6489
rect 35521 6455 35571 6456
rect 35605 6455 35621 6489
rect 35655 6502 35708 6539
rect 36001 6569 36013 6603
rect 36047 6569 36059 6603
rect 36001 6534 36059 6569
rect 35655 6454 35662 6502
rect 35655 6421 35708 6454
rect 35062 6371 35074 6405
rect 35062 6337 35108 6371
rect 35062 6303 35074 6337
rect 35062 6257 35108 6303
rect 35142 6405 35208 6417
rect 35142 6371 35158 6405
rect 35192 6371 35208 6405
rect 35142 6337 35208 6371
rect 35387 6385 35708 6421
rect 36001 6385 36059 6402
rect 35142 6303 35158 6337
rect 35192 6303 35208 6337
rect 35142 6291 35208 6303
rect 35300 6333 35353 6349
rect 35300 6299 35319 6333
rect 35300 6257 35353 6299
rect 35387 6341 35453 6385
rect 35387 6307 35403 6341
rect 35437 6307 35453 6341
rect 35387 6291 35453 6307
rect 35487 6333 35521 6349
rect 35487 6257 35521 6299
rect 35555 6341 35621 6385
rect 36001 6351 36013 6385
rect 36047 6351 36059 6385
rect 35555 6307 35571 6341
rect 35605 6307 35621 6341
rect 35555 6291 35621 6307
rect 35655 6334 35705 6350
rect 35689 6300 35705 6334
rect 35655 6257 35705 6300
rect 36001 6257 36059 6351
rect 30210 6223 30239 6257
rect 30273 6223 30302 6257
rect 30552 6223 30581 6257
rect 30615 6223 30673 6257
rect 30707 6223 30765 6257
rect 30799 6223 30857 6257
rect 30891 6223 30949 6257
rect 30983 6223 31041 6257
rect 31075 6223 31133 6257
rect 31167 6223 31225 6257
rect 31259 6223 31317 6257
rect 31351 6223 31409 6257
rect 31443 6223 31501 6257
rect 31535 6223 31593 6257
rect 31627 6223 31685 6257
rect 31719 6223 31777 6257
rect 31811 6223 31869 6257
rect 31903 6223 31961 6257
rect 31995 6223 32053 6257
rect 32087 6223 32145 6257
rect 32179 6223 32237 6257
rect 32271 6223 32329 6257
rect 32363 6223 32421 6257
rect 32455 6223 32513 6257
rect 32547 6223 32605 6257
rect 32639 6223 32697 6257
rect 32731 6223 32789 6257
rect 32823 6223 32881 6257
rect 32915 6223 32973 6257
rect 33007 6223 33036 6257
rect 33250 6223 33279 6257
rect 33313 6223 33371 6257
rect 33405 6223 33463 6257
rect 33497 6223 33555 6257
rect 33589 6223 33647 6257
rect 33681 6223 33739 6257
rect 33773 6223 33831 6257
rect 33865 6223 33923 6257
rect 33957 6223 34015 6257
rect 34049 6223 34107 6257
rect 34141 6223 34199 6257
rect 34233 6223 34291 6257
rect 34325 6223 34383 6257
rect 34417 6223 34475 6257
rect 34509 6223 34567 6257
rect 34601 6223 34659 6257
rect 34693 6223 34751 6257
rect 34785 6223 34843 6257
rect 34877 6223 34935 6257
rect 34969 6223 35027 6257
rect 35061 6223 35119 6257
rect 35153 6223 35211 6257
rect 35245 6223 35303 6257
rect 35337 6223 35395 6257
rect 35429 6223 35487 6257
rect 35521 6223 35579 6257
rect 35613 6223 35671 6257
rect 35705 6223 35734 6257
rect 35984 6223 36013 6257
rect 36047 6223 36076 6257
rect 30227 6129 30285 6223
rect 30655 6181 30721 6223
rect 30227 6095 30239 6129
rect 30273 6095 30285 6129
rect 30227 6078 30285 6095
rect 30587 6155 30621 6171
rect 30655 6147 30671 6181
rect 30705 6147 30721 6181
rect 30843 6181 30893 6223
rect 30755 6155 30792 6171
rect 30587 6113 30621 6121
rect 30789 6121 30792 6155
rect 30843 6147 30859 6181
rect 31232 6173 31306 6223
rect 30843 6131 30893 6147
rect 30927 6133 30944 6167
rect 30978 6133 30994 6167
rect 31033 6133 31055 6167
rect 31089 6133 31168 6167
rect 30587 6079 30720 6113
rect 30570 6025 30640 6045
rect 30570 6014 30584 6025
rect 30618 6014 30640 6025
rect 30570 5966 30576 6014
rect 30624 5966 30640 6014
rect 30227 5911 30285 5946
rect 30570 5915 30640 5966
rect 30674 6010 30720 6079
rect 30674 5976 30686 6010
rect 30227 5877 30239 5911
rect 30273 5877 30285 5911
rect 30674 5883 30720 5976
rect 30674 5881 30678 5883
rect 30227 5818 30285 5877
rect 30227 5784 30239 5818
rect 30273 5784 30285 5818
rect 30227 5713 30285 5784
rect 30587 5865 30678 5881
rect 30621 5849 30678 5865
rect 30712 5849 30720 5883
rect 30621 5847 30720 5849
rect 30755 5951 30792 6121
rect 30927 6105 30961 6133
rect 30755 5917 30757 5951
rect 30791 5917 30792 5951
rect 30755 5865 30792 5917
rect 30826 6062 30882 6097
rect 30826 6014 30832 6062
rect 30880 6014 30882 6062
rect 30826 5957 30882 6014
rect 30826 5923 30848 5957
rect 30826 5907 30882 5923
rect 30916 6079 30961 6105
rect 30995 6083 31100 6093
rect 30587 5797 30621 5831
rect 30789 5831 30792 5865
rect 30916 5858 30950 6079
rect 30995 6049 31011 6083
rect 31045 6049 31100 6083
rect 30984 5987 31032 6015
rect 30984 5953 30991 5987
rect 31025 5953 31032 5987
rect 30984 5951 31032 5953
rect 30984 5917 30995 5951
rect 31029 5917 31032 5951
rect 30984 5896 31032 5917
rect 31066 5883 31100 6049
rect 31134 5977 31168 6133
rect 31232 6139 31254 6173
rect 31288 6139 31306 6173
rect 31669 6167 31711 6223
rect 31232 6123 31306 6139
rect 31342 6133 31373 6167
rect 31407 6133 31423 6167
rect 31457 6133 31476 6167
rect 31510 6133 31614 6167
rect 31342 6087 31376 6133
rect 31210 6071 31376 6087
rect 31244 6037 31376 6071
rect 31210 6027 31376 6037
rect 31453 6083 31546 6099
rect 31487 6049 31546 6083
rect 31453 6033 31546 6049
rect 31210 6021 31250 6027
rect 31274 5977 31308 5991
rect 31134 5975 31308 5977
rect 31134 5943 31274 5975
rect 31206 5941 31274 5943
rect 31206 5925 31308 5941
rect 30916 5832 30977 5858
rect 31066 5849 31098 5883
rect 31134 5875 31172 5909
rect 31132 5849 31172 5875
rect 31066 5836 31172 5849
rect 30587 5747 30621 5763
rect 30655 5779 30671 5813
rect 30705 5779 30721 5813
rect 30655 5713 30721 5779
rect 30755 5797 30792 5831
rect 30789 5763 30792 5797
rect 30755 5747 30792 5763
rect 30840 5789 30893 5805
rect 30840 5755 30859 5789
rect 30840 5713 30893 5755
rect 30927 5797 30977 5832
rect 31206 5802 31240 5925
rect 30927 5763 30943 5797
rect 31019 5768 31035 5802
rect 31069 5768 31240 5802
rect 31274 5857 31308 5873
rect 31274 5789 31308 5823
rect 30927 5747 30977 5763
rect 31274 5713 31308 5755
rect 31342 5813 31376 6027
rect 31410 5975 31448 5991
rect 31444 5941 31448 5975
rect 31410 5883 31448 5941
rect 31410 5849 31412 5883
rect 31446 5849 31448 5883
rect 31410 5847 31448 5849
rect 31482 5951 31546 6033
rect 31482 5917 31499 5951
rect 31533 5917 31546 5951
rect 31482 5909 31546 5917
rect 31482 5875 31512 5909
rect 31482 5841 31546 5875
rect 31580 6041 31614 6133
rect 31669 6133 31674 6167
rect 31708 6133 31711 6167
rect 31669 6117 31711 6133
rect 31764 6146 31780 6180
rect 31814 6146 31830 6180
rect 31764 6112 31830 6146
rect 31764 6078 31780 6112
rect 31814 6078 31830 6112
rect 31864 6151 31898 6223
rect 32133 6181 32197 6223
rect 31864 6101 31898 6117
rect 31932 6178 31998 6179
rect 31932 6144 31948 6178
rect 31982 6144 31998 6178
rect 31932 6110 31998 6144
rect 32036 6155 32086 6171
rect 32036 6121 32052 6155
rect 32133 6147 32147 6181
rect 32181 6147 32197 6181
rect 32133 6131 32197 6147
rect 32231 6143 32282 6189
rect 32036 6117 32086 6121
rect 31764 6075 31830 6078
rect 31932 6076 31948 6110
rect 31982 6092 31998 6110
rect 31982 6076 32012 6092
rect 31932 6075 32012 6076
rect 31790 6041 31830 6075
rect 31963 6067 32012 6075
rect 31580 6025 31756 6041
rect 31580 5991 31722 6025
rect 31580 5975 31756 5991
rect 31790 6025 31940 6041
rect 31790 5991 31906 6025
rect 31790 5975 31940 5991
rect 31342 5797 31392 5813
rect 31580 5807 31614 5975
rect 31790 5934 31828 5975
rect 31974 5951 32012 6067
rect 31965 5941 32012 5951
rect 31648 5931 31828 5934
rect 31648 5909 31776 5931
rect 31682 5897 31776 5909
rect 31810 5897 31828 5931
rect 31930 5931 32012 5941
rect 31682 5875 31828 5897
rect 31648 5860 31828 5875
rect 31648 5859 31776 5860
rect 31760 5826 31776 5859
rect 31810 5826 31828 5860
rect 31342 5763 31358 5797
rect 31437 5773 31453 5807
rect 31487 5773 31614 5807
rect 31650 5797 31713 5813
rect 31342 5747 31392 5763
rect 31650 5763 31652 5797
rect 31686 5763 31713 5797
rect 31650 5713 31713 5763
rect 31760 5789 31828 5826
rect 31760 5755 31776 5789
rect 31810 5755 31828 5789
rect 31760 5747 31828 5755
rect 31862 5899 31896 5915
rect 31862 5819 31896 5865
rect 31862 5713 31896 5785
rect 31930 5897 31946 5931
rect 31980 5925 32012 5931
rect 32046 6041 32086 6117
rect 32265 6109 32282 6143
rect 32231 6058 32282 6109
rect 32364 6177 32410 6223
rect 32364 6143 32376 6177
rect 32364 6109 32410 6143
rect 32364 6075 32376 6109
rect 32364 6059 32410 6075
rect 32444 6177 32510 6189
rect 32444 6143 32460 6177
rect 32494 6143 32510 6177
rect 32444 6109 32510 6143
rect 32602 6181 32655 6223
rect 32602 6147 32621 6181
rect 32602 6131 32655 6147
rect 32689 6173 32755 6189
rect 32689 6139 32705 6173
rect 32739 6139 32755 6173
rect 32444 6075 32460 6109
rect 32494 6075 32510 6109
rect 32444 6063 32510 6075
rect 32046 6025 32201 6041
rect 32046 5991 32167 6025
rect 32046 5975 32201 5991
rect 32235 6024 32282 6058
rect 32364 6024 32380 6025
rect 32235 5976 32242 6024
rect 32414 5991 32430 6025
rect 32406 5977 32430 5991
rect 32464 6024 32510 6063
rect 32689 6095 32755 6139
rect 32789 6181 32823 6223
rect 32789 6131 32823 6147
rect 32857 6173 32923 6189
rect 32857 6139 32873 6173
rect 32907 6139 32923 6173
rect 32857 6095 32923 6139
rect 32957 6180 33007 6223
rect 32991 6146 33007 6180
rect 33353 6181 33419 6223
rect 32957 6130 33007 6146
rect 33285 6155 33319 6171
rect 33353 6147 33369 6181
rect 33403 6147 33419 6181
rect 33541 6181 33591 6223
rect 33453 6155 33490 6171
rect 33285 6113 33319 6121
rect 33487 6121 33490 6155
rect 33541 6147 33557 6181
rect 33930 6173 34004 6223
rect 33541 6131 33591 6147
rect 33625 6133 33642 6167
rect 33676 6133 33692 6167
rect 33731 6133 33753 6167
rect 33787 6133 33866 6167
rect 32689 6059 33010 6095
rect 33285 6079 33418 6113
rect 32957 6026 33010 6059
rect 33268 6032 33338 6045
rect 32597 6024 32613 6025
rect 32647 6024 32705 6025
rect 32739 6024 32789 6025
rect 32464 5976 32470 6024
rect 32597 5976 32602 6024
rect 32650 5991 32705 6024
rect 32760 5991 32789 6024
rect 32823 6024 32873 6025
rect 32823 5991 32828 6024
rect 32907 5991 32923 6025
rect 32650 5976 32712 5991
rect 32760 5976 32828 5991
rect 32876 5976 32923 5991
rect 31980 5897 31996 5925
rect 32046 5897 32100 5975
rect 32235 5944 32282 5976
rect 31930 5863 31996 5897
rect 31930 5842 31946 5863
rect 31980 5842 31996 5863
rect 31930 5794 31936 5842
rect 31984 5794 31996 5842
rect 31930 5761 31946 5794
rect 31980 5761 31996 5794
rect 31930 5756 31996 5761
rect 32034 5857 32100 5897
rect 32034 5823 32050 5857
rect 32084 5823 32100 5857
rect 32034 5789 32100 5823
rect 32034 5755 32050 5789
rect 32084 5755 32100 5789
rect 32034 5751 32100 5755
rect 32138 5925 32181 5941
rect 32138 5891 32147 5925
rect 32138 5857 32181 5891
rect 32138 5823 32147 5857
rect 32138 5789 32181 5823
rect 32138 5755 32147 5789
rect 32138 5713 32181 5755
rect 32215 5931 32282 5944
rect 32464 5943 32510 5976
rect 32597 5975 32923 5976
rect 32957 5978 32960 6026
rect 33268 5984 33282 6032
rect 33330 5984 33338 6032
rect 32215 5897 32231 5931
rect 32265 5897 32282 5931
rect 32215 5860 32282 5897
rect 32215 5826 32231 5860
rect 32265 5826 32282 5860
rect 32215 5789 32282 5826
rect 32215 5755 32231 5789
rect 32265 5755 32282 5789
rect 32215 5747 32282 5755
rect 32368 5925 32410 5941
rect 32368 5891 32376 5925
rect 32368 5857 32410 5891
rect 32368 5823 32376 5857
rect 32368 5789 32410 5823
rect 32368 5755 32376 5789
rect 32368 5713 32410 5755
rect 32444 5925 32510 5943
rect 32957 5941 33010 5978
rect 32444 5891 32460 5925
rect 32494 5891 32510 5925
rect 32444 5857 32510 5891
rect 32444 5823 32460 5857
rect 32494 5823 32510 5857
rect 32444 5789 32510 5823
rect 32444 5755 32460 5789
rect 32494 5755 32510 5789
rect 32444 5747 32510 5755
rect 32602 5925 32655 5941
rect 32602 5891 32621 5925
rect 32602 5857 32655 5891
rect 32602 5823 32621 5857
rect 32602 5789 32655 5823
rect 32602 5755 32621 5789
rect 32602 5713 32655 5755
rect 32689 5925 33010 5941
rect 32689 5891 32705 5925
rect 32739 5907 32873 5925
rect 32739 5891 32755 5907
rect 32689 5857 32755 5891
rect 32857 5891 32873 5907
rect 32907 5903 33010 5925
rect 33268 5915 33338 5984
rect 33372 6010 33418 6079
rect 33372 5976 33384 6010
rect 32907 5891 32923 5903
rect 32689 5823 32705 5857
rect 32739 5823 32755 5857
rect 32689 5789 32755 5823
rect 32689 5755 32705 5789
rect 32739 5755 32755 5789
rect 32689 5747 32755 5755
rect 32789 5857 32823 5873
rect 32789 5789 32823 5823
rect 32789 5713 32823 5755
rect 32857 5857 32923 5891
rect 33372 5883 33418 5976
rect 33372 5881 33376 5883
rect 32857 5823 32873 5857
rect 32907 5823 32923 5857
rect 32857 5789 32923 5823
rect 33285 5865 33376 5881
rect 33319 5849 33376 5865
rect 33410 5849 33418 5883
rect 33319 5847 33418 5849
rect 33453 5951 33490 6121
rect 33625 6105 33659 6133
rect 33453 5917 33455 5951
rect 33489 5917 33490 5951
rect 33453 5865 33490 5917
rect 33524 6062 33580 6097
rect 33524 6014 33530 6062
rect 33578 6014 33580 6062
rect 33524 5957 33580 6014
rect 33524 5923 33546 5957
rect 33524 5907 33580 5923
rect 33614 6079 33659 6105
rect 33693 6083 33798 6093
rect 32857 5755 32873 5789
rect 32907 5755 32923 5789
rect 32857 5747 32923 5755
rect 32957 5789 32999 5805
rect 32991 5755 32999 5789
rect 32957 5713 32999 5755
rect 33285 5797 33319 5831
rect 33487 5831 33490 5865
rect 33614 5858 33648 6079
rect 33693 6049 33709 6083
rect 33743 6049 33798 6083
rect 33682 5987 33730 6015
rect 33682 5953 33689 5987
rect 33723 5953 33730 5987
rect 33682 5951 33730 5953
rect 33682 5917 33693 5951
rect 33727 5917 33730 5951
rect 33682 5896 33730 5917
rect 33764 5883 33798 6049
rect 33832 5977 33866 6133
rect 33930 6139 33952 6173
rect 33986 6139 34004 6173
rect 34367 6167 34409 6223
rect 33930 6123 34004 6139
rect 34040 6133 34071 6167
rect 34105 6133 34121 6167
rect 34155 6133 34174 6167
rect 34208 6133 34312 6167
rect 34040 6087 34074 6133
rect 33908 6071 34074 6087
rect 33942 6037 34074 6071
rect 33908 6027 34074 6037
rect 34151 6083 34244 6099
rect 34185 6049 34244 6083
rect 34151 6033 34244 6049
rect 33908 6021 33948 6027
rect 33972 5977 34006 5991
rect 33832 5975 34006 5977
rect 33832 5943 33972 5975
rect 33904 5941 33972 5943
rect 33904 5925 34006 5941
rect 33614 5832 33675 5858
rect 33764 5849 33796 5883
rect 33832 5875 33870 5909
rect 33830 5849 33870 5875
rect 33764 5836 33870 5849
rect 33285 5747 33319 5763
rect 33353 5779 33369 5813
rect 33403 5779 33419 5813
rect 33353 5713 33419 5779
rect 33453 5797 33490 5831
rect 33487 5763 33490 5797
rect 33453 5747 33490 5763
rect 33538 5789 33591 5805
rect 33538 5755 33557 5789
rect 33538 5713 33591 5755
rect 33625 5797 33675 5832
rect 33904 5802 33938 5925
rect 33625 5763 33641 5797
rect 33717 5768 33733 5802
rect 33767 5768 33938 5802
rect 33972 5857 34006 5873
rect 33972 5789 34006 5823
rect 33625 5747 33675 5763
rect 33972 5713 34006 5755
rect 34040 5813 34074 6027
rect 34108 5975 34146 5991
rect 34142 5941 34146 5975
rect 34108 5883 34146 5941
rect 34108 5849 34110 5883
rect 34144 5849 34146 5883
rect 34108 5847 34146 5849
rect 34180 5951 34244 6033
rect 34180 5917 34197 5951
rect 34231 5917 34244 5951
rect 34180 5909 34244 5917
rect 34180 5875 34210 5909
rect 34180 5841 34244 5875
rect 34278 6041 34312 6133
rect 34367 6133 34372 6167
rect 34406 6133 34409 6167
rect 34367 6117 34409 6133
rect 34462 6146 34478 6180
rect 34512 6146 34528 6180
rect 34462 6112 34528 6146
rect 34462 6078 34478 6112
rect 34512 6078 34528 6112
rect 34562 6151 34596 6223
rect 34831 6181 34895 6223
rect 34562 6101 34596 6117
rect 34630 6178 34696 6179
rect 34630 6144 34646 6178
rect 34680 6144 34696 6178
rect 34630 6142 34696 6144
rect 34462 6075 34528 6078
rect 34630 6094 34634 6142
rect 34682 6094 34696 6142
rect 34734 6155 34784 6171
rect 34734 6121 34750 6155
rect 34831 6147 34845 6181
rect 34879 6147 34895 6181
rect 34831 6131 34895 6147
rect 34929 6143 34980 6189
rect 34734 6117 34784 6121
rect 34630 6076 34646 6094
rect 34680 6092 34696 6094
rect 34680 6076 34710 6092
rect 34630 6075 34710 6076
rect 34488 6041 34528 6075
rect 34661 6067 34710 6075
rect 34278 6025 34454 6041
rect 34278 5991 34420 6025
rect 34278 5975 34454 5991
rect 34488 6025 34638 6041
rect 34488 5991 34604 6025
rect 34488 5975 34638 5991
rect 34040 5797 34090 5813
rect 34278 5807 34312 5975
rect 34488 5934 34526 5975
rect 34672 5951 34710 6067
rect 34663 5941 34710 5951
rect 34346 5931 34526 5934
rect 34346 5909 34474 5931
rect 34380 5897 34474 5909
rect 34508 5897 34526 5931
rect 34628 5931 34710 5941
rect 34380 5875 34526 5897
rect 34346 5860 34526 5875
rect 34346 5859 34474 5860
rect 34458 5826 34474 5859
rect 34508 5826 34526 5860
rect 34040 5763 34056 5797
rect 34135 5773 34151 5807
rect 34185 5773 34312 5807
rect 34348 5797 34411 5813
rect 34040 5747 34090 5763
rect 34348 5763 34350 5797
rect 34384 5763 34411 5797
rect 34348 5713 34411 5763
rect 34458 5789 34526 5826
rect 34458 5755 34474 5789
rect 34508 5755 34526 5789
rect 34458 5747 34526 5755
rect 34560 5899 34594 5915
rect 34560 5819 34594 5865
rect 34560 5713 34594 5785
rect 34628 5897 34644 5931
rect 34678 5925 34710 5931
rect 34744 6041 34784 6117
rect 34963 6109 34980 6143
rect 34929 6058 34980 6109
rect 35062 6177 35108 6223
rect 35062 6143 35074 6177
rect 35062 6109 35108 6143
rect 35062 6075 35074 6109
rect 35062 6059 35108 6075
rect 35142 6177 35208 6189
rect 35142 6143 35158 6177
rect 35192 6143 35208 6177
rect 35142 6109 35208 6143
rect 35300 6181 35353 6223
rect 35300 6147 35319 6181
rect 35300 6131 35353 6147
rect 35387 6173 35453 6189
rect 35387 6139 35403 6173
rect 35437 6139 35453 6173
rect 35142 6075 35158 6109
rect 35192 6075 35208 6109
rect 35142 6063 35208 6075
rect 34744 6025 34899 6041
rect 34744 5991 34865 6025
rect 34744 5975 34899 5991
rect 34933 6024 34980 6058
rect 35062 6024 35078 6025
rect 34933 5976 34940 6024
rect 35112 5991 35128 6025
rect 35104 5977 35128 5991
rect 35162 6024 35208 6063
rect 35387 6095 35453 6139
rect 35487 6181 35521 6223
rect 35487 6131 35521 6147
rect 35555 6173 35621 6189
rect 35555 6139 35571 6173
rect 35605 6139 35621 6173
rect 35555 6095 35621 6139
rect 35655 6180 35705 6223
rect 35689 6146 35705 6180
rect 35655 6130 35705 6146
rect 36001 6129 36059 6223
rect 36001 6095 36013 6129
rect 36047 6095 36059 6129
rect 35387 6059 35708 6095
rect 36001 6078 36059 6095
rect 35655 6026 35708 6059
rect 35295 6024 35311 6025
rect 35345 6024 35403 6025
rect 35437 6024 35487 6025
rect 35162 5976 35168 6024
rect 35295 5976 35300 6024
rect 35348 5991 35403 6024
rect 35458 5991 35487 6024
rect 35521 6024 35571 6025
rect 35521 5991 35526 6024
rect 35605 5991 35621 6025
rect 35348 5976 35410 5991
rect 35458 5976 35526 5991
rect 35574 5976 35621 5991
rect 34678 5897 34694 5925
rect 34744 5897 34798 5975
rect 34933 5944 34980 5976
rect 34628 5863 34694 5897
rect 34628 5829 34644 5863
rect 34678 5829 34694 5863
rect 34628 5795 34694 5829
rect 34628 5761 34644 5795
rect 34678 5761 34694 5795
rect 34628 5756 34694 5761
rect 34732 5857 34798 5897
rect 34732 5823 34748 5857
rect 34782 5823 34798 5857
rect 34732 5789 34798 5823
rect 34732 5755 34748 5789
rect 34782 5755 34798 5789
rect 34732 5751 34798 5755
rect 34836 5925 34879 5941
rect 34836 5891 34845 5925
rect 34836 5857 34879 5891
rect 34836 5823 34845 5857
rect 34836 5789 34879 5823
rect 34836 5755 34845 5789
rect 34836 5713 34879 5755
rect 34913 5931 34980 5944
rect 35162 5943 35208 5976
rect 35295 5975 35621 5976
rect 35655 5978 35658 6026
rect 35706 5978 35708 6026
rect 34913 5897 34929 5931
rect 34963 5897 34980 5931
rect 34913 5860 34980 5897
rect 34913 5826 34929 5860
rect 34963 5826 34980 5860
rect 34913 5789 34980 5826
rect 34913 5755 34929 5789
rect 34963 5755 34980 5789
rect 34913 5747 34980 5755
rect 35066 5925 35108 5941
rect 35066 5891 35074 5925
rect 35066 5857 35108 5891
rect 35066 5823 35074 5857
rect 35066 5789 35108 5823
rect 35066 5755 35074 5789
rect 35066 5713 35108 5755
rect 35142 5925 35208 5943
rect 35655 5941 35708 5978
rect 35142 5891 35158 5925
rect 35192 5891 35208 5925
rect 35142 5857 35208 5891
rect 35142 5823 35158 5857
rect 35192 5823 35208 5857
rect 35142 5789 35208 5823
rect 35142 5755 35158 5789
rect 35192 5755 35208 5789
rect 35142 5747 35208 5755
rect 35300 5925 35353 5941
rect 35300 5891 35319 5925
rect 35300 5857 35353 5891
rect 35300 5823 35319 5857
rect 35300 5789 35353 5823
rect 35300 5755 35319 5789
rect 35300 5713 35353 5755
rect 35387 5925 35708 5941
rect 35387 5891 35403 5925
rect 35437 5907 35571 5925
rect 35437 5891 35453 5907
rect 35387 5857 35453 5891
rect 35555 5891 35571 5907
rect 35605 5903 35708 5925
rect 36001 5911 36059 5946
rect 35605 5891 35621 5903
rect 35387 5823 35403 5857
rect 35437 5823 35453 5857
rect 35387 5789 35453 5823
rect 35387 5755 35403 5789
rect 35437 5755 35453 5789
rect 35387 5747 35453 5755
rect 35487 5857 35521 5873
rect 35487 5789 35521 5823
rect 35487 5713 35521 5755
rect 35555 5857 35621 5891
rect 35555 5823 35571 5857
rect 35605 5823 35621 5857
rect 35555 5789 35621 5823
rect 36001 5877 36013 5911
rect 36047 5877 36059 5911
rect 36001 5818 36059 5877
rect 35555 5755 35571 5789
rect 35605 5755 35621 5789
rect 35555 5747 35621 5755
rect 35655 5789 35697 5805
rect 35689 5755 35697 5789
rect 35655 5713 35697 5755
rect 36001 5784 36013 5818
rect 36047 5784 36059 5818
rect 36001 5713 36059 5784
rect 30210 5679 30239 5713
rect 30273 5679 30302 5713
rect 30552 5679 30581 5713
rect 30615 5679 30673 5713
rect 30707 5679 30765 5713
rect 30799 5679 30857 5713
rect 30891 5679 30949 5713
rect 30983 5679 31041 5713
rect 31075 5679 31133 5713
rect 31167 5679 31225 5713
rect 31259 5679 31317 5713
rect 31351 5679 31409 5713
rect 31443 5679 31501 5713
rect 31535 5679 31593 5713
rect 31627 5679 31685 5713
rect 31719 5679 31777 5713
rect 31811 5679 31869 5713
rect 31903 5679 31961 5713
rect 31995 5679 32053 5713
rect 32087 5679 32145 5713
rect 32179 5679 32237 5713
rect 32271 5679 32329 5713
rect 32363 5679 32421 5713
rect 32455 5679 32513 5713
rect 32547 5679 32605 5713
rect 32639 5679 32697 5713
rect 32731 5679 32789 5713
rect 32823 5679 32881 5713
rect 32915 5679 32973 5713
rect 33007 5679 33036 5713
rect 33250 5679 33279 5713
rect 33313 5679 33371 5713
rect 33405 5679 33463 5713
rect 33497 5679 33555 5713
rect 33589 5679 33647 5713
rect 33681 5679 33739 5713
rect 33773 5679 33831 5713
rect 33865 5679 33923 5713
rect 33957 5679 34015 5713
rect 34049 5679 34107 5713
rect 34141 5679 34199 5713
rect 34233 5679 34291 5713
rect 34325 5679 34383 5713
rect 34417 5679 34475 5713
rect 34509 5679 34567 5713
rect 34601 5679 34659 5713
rect 34693 5679 34751 5713
rect 34785 5679 34843 5713
rect 34877 5679 34935 5713
rect 34969 5679 35027 5713
rect 35061 5679 35119 5713
rect 35153 5679 35211 5713
rect 35245 5679 35303 5713
rect 35337 5679 35395 5713
rect 35429 5679 35487 5713
rect 35521 5679 35579 5713
rect 35613 5679 35671 5713
rect 35705 5679 35734 5713
rect 35984 5679 36013 5713
rect 36047 5679 36076 5713
rect 28886 4766 28986 4928
rect 8352 4234 8452 4396
rect 18696 4234 18796 4396
rect 9458 2991 9474 3025
rect 9694 2991 9710 3025
rect 9916 2991 9932 3025
rect 10152 2991 10168 3025
rect 10374 2991 10390 3025
rect 10610 2991 10626 3025
rect 10832 2991 10848 3025
rect 11068 2991 11084 3025
rect 11290 2991 11306 3025
rect 11526 2991 11542 3025
rect 11748 2991 11764 3025
rect 11984 2991 12000 3025
rect 12206 2991 12222 3025
rect 12442 2991 12458 3025
rect 12664 2991 12680 3025
rect 12900 2991 12916 3025
rect 13122 2991 13138 3025
rect 13358 2991 13374 3025
rect 13580 2991 13596 3025
rect 13816 2991 13832 3025
rect 14038 2991 14054 3025
rect 14274 2991 14290 3025
rect 14496 2991 14512 3025
rect 14732 2991 14748 3025
rect 14954 2991 14970 3025
rect 15190 2991 15206 3025
rect 15412 2991 15428 3025
rect 15648 2991 15664 3025
rect 15870 2991 15886 3025
rect 16106 2991 16122 3025
rect 16328 2991 16344 3025
rect 16564 2991 16580 3025
rect 16786 2991 16802 3025
rect 17022 2991 17038 3025
rect 17244 2991 17260 3025
rect 17480 2991 17496 3025
rect 9338 2932 9372 2948
rect 9338 1340 9372 1356
rect 9796 2932 9830 2948
rect 9796 1340 9830 1356
rect 10254 2932 10288 2948
rect 10254 1340 10288 1356
rect 10712 2932 10746 2948
rect 10712 1340 10746 1356
rect 11170 2932 11204 2948
rect 11170 1340 11204 1356
rect 11628 2932 11662 2948
rect 11628 1340 11662 1356
rect 12086 2932 12120 2948
rect 12086 1340 12120 1356
rect 12544 2932 12578 2948
rect 12544 1340 12578 1356
rect 13002 2932 13036 2948
rect 13002 1340 13036 1356
rect 13460 2932 13494 2948
rect 13460 1340 13494 1356
rect 13918 2932 13952 2948
rect 13918 1340 13952 1356
rect 14376 2932 14410 2948
rect 14376 1340 14410 1356
rect 14834 2932 14868 2948
rect 14834 1340 14868 1356
rect 15292 2932 15326 2948
rect 15292 1340 15326 1356
rect 15750 2932 15784 2948
rect 15750 1340 15784 1356
rect 16208 2932 16242 2948
rect 16208 1340 16242 1356
rect 16666 2932 16700 2948
rect 16666 1340 16700 1356
rect 17124 2932 17158 2948
rect 17124 1340 17158 1356
rect 17582 2932 17616 2948
rect 17582 1340 17616 1356
rect 9458 1263 9474 1297
rect 9694 1263 9710 1297
rect 9916 1263 9932 1297
rect 10152 1263 10168 1297
rect 10374 1263 10390 1297
rect 10610 1263 10626 1297
rect 10832 1263 10848 1297
rect 11068 1263 11084 1297
rect 11290 1263 11306 1297
rect 11526 1263 11542 1297
rect 11748 1263 11764 1297
rect 11984 1263 12000 1297
rect 12206 1263 12222 1297
rect 12442 1263 12458 1297
rect 12664 1263 12680 1297
rect 12900 1263 12916 1297
rect 13122 1263 13138 1297
rect 13358 1263 13374 1297
rect 13580 1263 13596 1297
rect 13816 1263 13832 1297
rect 14038 1263 14054 1297
rect 14274 1263 14290 1297
rect 14496 1263 14512 1297
rect 14732 1263 14748 1297
rect 14954 1263 14970 1297
rect 15190 1263 15206 1297
rect 15412 1263 15428 1297
rect 15648 1263 15664 1297
rect 15870 1263 15886 1297
rect 16106 1263 16122 1297
rect 16328 1263 16344 1297
rect 16564 1263 16580 1297
rect 16786 1263 16802 1297
rect 17022 1263 17038 1297
rect 17244 1263 17260 1297
rect 17480 1263 17496 1297
rect 13216 1180 13676 1186
rect 13216 1132 13222 1180
rect 13270 1132 13676 1180
rect 13216 1126 13676 1132
rect 8899 326 8915 360
rect 9135 326 9151 360
rect 9357 326 9373 360
rect 9593 326 9609 360
rect 9815 326 9831 360
rect 10051 326 10067 360
rect 10273 326 10289 360
rect 10509 326 10525 360
rect 10731 326 10747 360
rect 10967 326 10983 360
rect 11189 326 11205 360
rect 11425 326 11441 360
rect 11647 326 11663 360
rect 11883 326 11899 360
rect 12105 326 12121 360
rect 12341 326 12357 360
rect 12563 326 12579 360
rect 12799 326 12815 360
rect 13021 326 13037 360
rect 13257 326 13273 360
rect 13899 326 13915 360
rect 14135 326 14151 360
rect 14357 326 14373 360
rect 14593 326 14609 360
rect 14815 326 14831 360
rect 15051 326 15067 360
rect 15273 326 15289 360
rect 15509 326 15525 360
rect 15731 326 15747 360
rect 15967 326 15983 360
rect 16189 326 16205 360
rect 16425 326 16441 360
rect 16647 326 16663 360
rect 16883 326 16899 360
rect 17105 326 17121 360
rect 17341 326 17357 360
rect 17563 326 17579 360
rect 17799 326 17815 360
rect 18021 326 18037 360
rect 18257 326 18273 360
rect 8779 267 8813 283
rect 8779 -925 8813 -909
rect 9237 267 9271 283
rect 9237 -925 9271 -909
rect 9695 267 9729 283
rect 9695 -925 9729 -909
rect 10153 267 10187 283
rect 10153 -925 10187 -909
rect 10611 267 10645 283
rect 10611 -925 10645 -909
rect 11069 267 11103 283
rect 11069 -925 11103 -909
rect 11527 267 11561 283
rect 11527 -925 11561 -909
rect 11985 267 12019 283
rect 11985 -925 12019 -909
rect 12443 267 12477 283
rect 12443 -925 12477 -909
rect 12901 267 12935 283
rect 12901 -925 12935 -909
rect 13359 267 13393 283
rect 13359 -925 13393 -909
rect 13779 267 13813 283
rect 13779 -925 13813 -909
rect 14237 267 14271 283
rect 14237 -925 14271 -909
rect 14695 267 14729 283
rect 14695 -925 14729 -909
rect 15153 267 15187 283
rect 15153 -925 15187 -909
rect 15611 267 15645 283
rect 15611 -925 15645 -909
rect 16069 267 16103 283
rect 16069 -925 16103 -909
rect 16527 267 16561 283
rect 16527 -925 16561 -909
rect 16985 267 17019 283
rect 16985 -925 17019 -909
rect 17443 267 17477 283
rect 17443 -925 17477 -909
rect 17901 267 17935 283
rect 17901 -925 17935 -909
rect 18359 267 18393 283
rect 18359 -925 18393 -909
rect 8899 -1002 8915 -968
rect 9135 -1002 9151 -968
rect 9357 -1002 9373 -968
rect 9593 -1002 9609 -968
rect 9815 -1002 9831 -968
rect 10051 -1002 10067 -968
rect 10273 -1002 10289 -968
rect 10509 -1002 10525 -968
rect 10731 -1002 10747 -968
rect 10967 -1002 10983 -968
rect 11189 -1002 11205 -968
rect 11425 -1002 11441 -968
rect 11647 -1002 11663 -968
rect 11883 -1002 11899 -968
rect 12105 -1002 12121 -968
rect 12341 -1002 12357 -968
rect 12563 -1002 12579 -968
rect 12799 -1002 12815 -968
rect 13021 -1002 13037 -968
rect 13257 -1002 13273 -968
rect 13899 -1002 13915 -968
rect 14135 -1002 14151 -968
rect 14357 -1002 14373 -968
rect 14593 -1002 14609 -968
rect 14815 -1002 14831 -968
rect 15051 -1002 15067 -968
rect 15273 -1002 15289 -968
rect 15509 -1002 15525 -968
rect 15731 -1002 15747 -968
rect 15967 -1002 15983 -968
rect 16189 -1002 16205 -968
rect 16425 -1002 16441 -968
rect 16647 -1002 16663 -968
rect 16883 -1002 16899 -968
rect 17105 -1002 17121 -968
rect 17341 -1002 17357 -968
rect 17563 -1002 17579 -968
rect 17799 -1002 17815 -968
rect 18021 -1002 18037 -968
rect 18257 -1002 18273 -968
rect 8352 -1448 8452 -1286
rect 18696 -1448 18796 -1286
rect 23352 4234 23452 4396
rect 33696 4234 33796 4396
rect 24458 2991 24474 3025
rect 24694 2991 24710 3025
rect 24916 2991 24932 3025
rect 25152 2991 25168 3025
rect 25374 2991 25390 3025
rect 25610 2991 25626 3025
rect 25832 2991 25848 3025
rect 26068 2991 26084 3025
rect 26290 2991 26306 3025
rect 26526 2991 26542 3025
rect 26748 2991 26764 3025
rect 26984 2991 27000 3025
rect 27206 2991 27222 3025
rect 27442 2991 27458 3025
rect 27664 2991 27680 3025
rect 27900 2991 27916 3025
rect 28122 2991 28138 3025
rect 28358 2991 28374 3025
rect 28580 2991 28596 3025
rect 28816 2991 28832 3025
rect 29038 2991 29054 3025
rect 29274 2991 29290 3025
rect 29496 2991 29512 3025
rect 29732 2991 29748 3025
rect 29954 2991 29970 3025
rect 30190 2991 30206 3025
rect 30412 2991 30428 3025
rect 30648 2991 30664 3025
rect 30870 2991 30886 3025
rect 31106 2991 31122 3025
rect 31328 2991 31344 3025
rect 31564 2991 31580 3025
rect 31786 2991 31802 3025
rect 32022 2991 32038 3025
rect 32244 2991 32260 3025
rect 32480 2991 32496 3025
rect 24338 2932 24372 2948
rect 24338 1340 24372 1356
rect 24796 2932 24830 2948
rect 24796 1340 24830 1356
rect 25254 2932 25288 2948
rect 25254 1340 25288 1356
rect 25712 2932 25746 2948
rect 25712 1340 25746 1356
rect 26170 2932 26204 2948
rect 26170 1340 26204 1356
rect 26628 2932 26662 2948
rect 26628 1340 26662 1356
rect 27086 2932 27120 2948
rect 27086 1340 27120 1356
rect 27544 2932 27578 2948
rect 27544 1340 27578 1356
rect 28002 2932 28036 2948
rect 28002 1340 28036 1356
rect 28460 2932 28494 2948
rect 28460 1340 28494 1356
rect 28918 2932 28952 2948
rect 28918 1340 28952 1356
rect 29376 2932 29410 2948
rect 29376 1340 29410 1356
rect 29834 2932 29868 2948
rect 29834 1340 29868 1356
rect 30292 2932 30326 2948
rect 30292 1340 30326 1356
rect 30750 2932 30784 2948
rect 30750 1340 30784 1356
rect 31208 2932 31242 2948
rect 31208 1340 31242 1356
rect 31666 2932 31700 2948
rect 31666 1340 31700 1356
rect 32124 2932 32158 2948
rect 32124 1340 32158 1356
rect 32582 2932 32616 2948
rect 32582 1340 32616 1356
rect 24458 1263 24474 1297
rect 24694 1263 24710 1297
rect 24916 1263 24932 1297
rect 25152 1263 25168 1297
rect 25374 1263 25390 1297
rect 25610 1263 25626 1297
rect 25832 1263 25848 1297
rect 26068 1263 26084 1297
rect 26290 1263 26306 1297
rect 26526 1263 26542 1297
rect 26748 1263 26764 1297
rect 26984 1263 27000 1297
rect 27206 1263 27222 1297
rect 27442 1263 27458 1297
rect 27664 1263 27680 1297
rect 27900 1263 27916 1297
rect 28122 1263 28138 1297
rect 28358 1263 28374 1297
rect 28580 1263 28596 1297
rect 28816 1263 28832 1297
rect 29038 1263 29054 1297
rect 29274 1263 29290 1297
rect 29496 1263 29512 1297
rect 29732 1263 29748 1297
rect 29954 1263 29970 1297
rect 30190 1263 30206 1297
rect 30412 1263 30428 1297
rect 30648 1263 30664 1297
rect 30870 1263 30886 1297
rect 31106 1263 31122 1297
rect 31328 1263 31344 1297
rect 31564 1263 31580 1297
rect 31786 1263 31802 1297
rect 32022 1263 32038 1297
rect 32244 1263 32260 1297
rect 32480 1263 32496 1297
rect 28216 1180 28676 1186
rect 28216 1132 28222 1180
rect 28270 1132 28676 1180
rect 28216 1126 28676 1132
rect 23899 326 23915 360
rect 24135 326 24151 360
rect 24357 326 24373 360
rect 24593 326 24609 360
rect 24815 326 24831 360
rect 25051 326 25067 360
rect 25273 326 25289 360
rect 25509 326 25525 360
rect 25731 326 25747 360
rect 25967 326 25983 360
rect 26189 326 26205 360
rect 26425 326 26441 360
rect 26647 326 26663 360
rect 26883 326 26899 360
rect 27105 326 27121 360
rect 27341 326 27357 360
rect 27563 326 27579 360
rect 27799 326 27815 360
rect 28021 326 28037 360
rect 28257 326 28273 360
rect 28899 326 28915 360
rect 29135 326 29151 360
rect 29357 326 29373 360
rect 29593 326 29609 360
rect 29815 326 29831 360
rect 30051 326 30067 360
rect 30273 326 30289 360
rect 30509 326 30525 360
rect 30731 326 30747 360
rect 30967 326 30983 360
rect 31189 326 31205 360
rect 31425 326 31441 360
rect 31647 326 31663 360
rect 31883 326 31899 360
rect 32105 326 32121 360
rect 32341 326 32357 360
rect 32563 326 32579 360
rect 32799 326 32815 360
rect 33021 326 33037 360
rect 33257 326 33273 360
rect 23779 267 23813 283
rect 23779 -925 23813 -909
rect 24237 267 24271 283
rect 24237 -925 24271 -909
rect 24695 267 24729 283
rect 24695 -925 24729 -909
rect 25153 267 25187 283
rect 25153 -925 25187 -909
rect 25611 267 25645 283
rect 25611 -925 25645 -909
rect 26069 267 26103 283
rect 26069 -925 26103 -909
rect 26527 267 26561 283
rect 26527 -925 26561 -909
rect 26985 267 27019 283
rect 26985 -925 27019 -909
rect 27443 267 27477 283
rect 27443 -925 27477 -909
rect 27901 267 27935 283
rect 27901 -925 27935 -909
rect 28359 267 28393 283
rect 28359 -925 28393 -909
rect 28779 267 28813 283
rect 28779 -925 28813 -909
rect 29237 267 29271 283
rect 29237 -925 29271 -909
rect 29695 267 29729 283
rect 29695 -925 29729 -909
rect 30153 267 30187 283
rect 30153 -925 30187 -909
rect 30611 267 30645 283
rect 30611 -925 30645 -909
rect 31069 267 31103 283
rect 31069 -925 31103 -909
rect 31527 267 31561 283
rect 31527 -925 31561 -909
rect 31985 267 32019 283
rect 31985 -925 32019 -909
rect 32443 267 32477 283
rect 32443 -925 32477 -909
rect 32901 267 32935 283
rect 32901 -925 32935 -909
rect 33359 267 33393 283
rect 33359 -925 33393 -909
rect 23899 -1002 23915 -968
rect 24135 -1002 24151 -968
rect 24357 -1002 24373 -968
rect 24593 -1002 24609 -968
rect 24815 -1002 24831 -968
rect 25051 -1002 25067 -968
rect 25273 -1002 25289 -968
rect 25509 -1002 25525 -968
rect 25731 -1002 25747 -968
rect 25967 -1002 25983 -968
rect 26189 -1002 26205 -968
rect 26425 -1002 26441 -968
rect 26647 -1002 26663 -968
rect 26883 -1002 26899 -968
rect 27105 -1002 27121 -968
rect 27341 -1002 27357 -968
rect 27563 -1002 27579 -968
rect 27799 -1002 27815 -968
rect 28021 -1002 28037 -968
rect 28257 -1002 28273 -968
rect 28899 -1002 28915 -968
rect 29135 -1002 29151 -968
rect 29357 -1002 29373 -968
rect 29593 -1002 29609 -968
rect 29815 -1002 29831 -968
rect 30051 -1002 30067 -968
rect 30273 -1002 30289 -968
rect 30509 -1002 30525 -968
rect 30731 -1002 30747 -968
rect 30967 -1002 30983 -968
rect 31189 -1002 31205 -968
rect 31425 -1002 31441 -968
rect 31647 -1002 31663 -968
rect 31883 -1002 31899 -968
rect 32105 -1002 32121 -968
rect 32341 -1002 32357 -968
rect 32563 -1002 32579 -968
rect 32799 -1002 32815 -968
rect 33021 -1002 33037 -968
rect 33257 -1002 33273 -968
rect 23352 -1448 23452 -1286
rect 33696 -1448 33796 -1286
rect 8352 -1846 8452 -1684
rect 18696 -1846 18796 -1684
rect 8898 -2176 8914 -2142
rect 9134 -2176 9150 -2142
rect 9356 -2176 9372 -2142
rect 9592 -2176 9608 -2142
rect 9814 -2176 9830 -2142
rect 10050 -2176 10066 -2142
rect 10272 -2176 10288 -2142
rect 10508 -2176 10524 -2142
rect 10730 -2176 10746 -2142
rect 10966 -2176 10982 -2142
rect 11188 -2176 11204 -2142
rect 11424 -2176 11440 -2142
rect 11646 -2176 11662 -2142
rect 11882 -2176 11898 -2142
rect 12104 -2176 12120 -2142
rect 12340 -2176 12356 -2142
rect 12562 -2176 12578 -2142
rect 12798 -2176 12814 -2142
rect 13020 -2176 13036 -2142
rect 13256 -2176 13272 -2142
rect 13898 -2176 13914 -2142
rect 14134 -2176 14150 -2142
rect 14356 -2176 14372 -2142
rect 14592 -2176 14608 -2142
rect 14814 -2176 14830 -2142
rect 15050 -2176 15066 -2142
rect 15272 -2176 15288 -2142
rect 15508 -2176 15524 -2142
rect 15730 -2176 15746 -2142
rect 15966 -2176 15982 -2142
rect 16188 -2176 16204 -2142
rect 16424 -2176 16440 -2142
rect 16646 -2176 16662 -2142
rect 16882 -2176 16898 -2142
rect 17104 -2176 17120 -2142
rect 17340 -2176 17356 -2142
rect 17562 -2176 17578 -2142
rect 17798 -2176 17814 -2142
rect 18020 -2176 18036 -2142
rect 18256 -2176 18272 -2142
rect 8778 -2226 8812 -2210
rect 8778 -2418 8812 -2402
rect 9236 -2226 9270 -2210
rect 9236 -2418 9270 -2402
rect 9694 -2226 9728 -2210
rect 9694 -2418 9728 -2402
rect 10152 -2226 10186 -2210
rect 10152 -2418 10186 -2402
rect 10610 -2226 10644 -2210
rect 10610 -2418 10644 -2402
rect 11068 -2226 11102 -2210
rect 11068 -2418 11102 -2402
rect 11526 -2226 11560 -2210
rect 11526 -2418 11560 -2402
rect 11984 -2226 12018 -2210
rect 11984 -2418 12018 -2402
rect 12442 -2226 12476 -2210
rect 12442 -2418 12476 -2402
rect 12900 -2226 12934 -2210
rect 12900 -2418 12934 -2402
rect 13358 -2226 13392 -2210
rect 13358 -2418 13392 -2402
rect 13778 -2226 13812 -2210
rect 13778 -2418 13812 -2402
rect 14236 -2226 14270 -2210
rect 14236 -2418 14270 -2402
rect 14694 -2226 14728 -2210
rect 14694 -2418 14728 -2402
rect 15152 -2226 15186 -2210
rect 15152 -2418 15186 -2402
rect 15610 -2226 15644 -2210
rect 15610 -2418 15644 -2402
rect 16068 -2226 16102 -2210
rect 16068 -2418 16102 -2402
rect 16526 -2226 16560 -2210
rect 16526 -2418 16560 -2402
rect 16984 -2226 17018 -2210
rect 16984 -2418 17018 -2402
rect 17442 -2226 17476 -2210
rect 17442 -2418 17476 -2402
rect 17900 -2226 17934 -2210
rect 17900 -2418 17934 -2402
rect 18358 -2226 18392 -2210
rect 18358 -2418 18392 -2402
rect 8898 -2486 8914 -2452
rect 9134 -2486 9150 -2452
rect 9356 -2486 9372 -2452
rect 9592 -2486 9608 -2452
rect 9814 -2486 9830 -2452
rect 10050 -2486 10066 -2452
rect 10272 -2486 10288 -2452
rect 10508 -2486 10524 -2452
rect 10730 -2486 10746 -2452
rect 10966 -2486 10982 -2452
rect 11188 -2486 11204 -2452
rect 11424 -2486 11440 -2452
rect 11646 -2486 11662 -2452
rect 11882 -2486 11898 -2452
rect 12104 -2486 12120 -2452
rect 12340 -2486 12356 -2452
rect 12562 -2486 12578 -2452
rect 12798 -2486 12814 -2452
rect 13020 -2486 13036 -2452
rect 13256 -2486 13272 -2452
rect 13898 -2486 13914 -2452
rect 14134 -2486 14150 -2452
rect 14356 -2486 14372 -2452
rect 14592 -2486 14608 -2452
rect 14814 -2486 14830 -2452
rect 15050 -2486 15066 -2452
rect 15272 -2486 15288 -2452
rect 15508 -2486 15524 -2452
rect 15730 -2486 15746 -2452
rect 15966 -2486 15982 -2452
rect 16188 -2486 16204 -2452
rect 16424 -2486 16440 -2452
rect 16646 -2486 16662 -2452
rect 16882 -2486 16898 -2452
rect 17104 -2486 17120 -2452
rect 17340 -2486 17356 -2452
rect 17562 -2486 17578 -2452
rect 17798 -2486 17814 -2452
rect 18020 -2486 18036 -2452
rect 18256 -2486 18272 -2452
rect 8898 -2844 8914 -2810
rect 9134 -2844 9150 -2810
rect 9356 -2844 9372 -2810
rect 9592 -2844 9608 -2810
rect 9814 -2844 9830 -2810
rect 10050 -2844 10066 -2810
rect 10272 -2844 10288 -2810
rect 10508 -2844 10524 -2810
rect 10730 -2844 10746 -2810
rect 10966 -2844 10982 -2810
rect 11188 -2844 11204 -2810
rect 11424 -2844 11440 -2810
rect 11646 -2844 11662 -2810
rect 11882 -2844 11898 -2810
rect 12104 -2844 12120 -2810
rect 12340 -2844 12356 -2810
rect 12562 -2844 12578 -2810
rect 12798 -2844 12814 -2810
rect 13020 -2844 13036 -2810
rect 13256 -2844 13272 -2810
rect 8778 -2894 8812 -2878
rect 8778 -3086 8812 -3070
rect 9236 -2894 9270 -2878
rect 9236 -3086 9270 -3070
rect 9694 -2894 9728 -2878
rect 9694 -3086 9728 -3070
rect 10152 -2894 10186 -2878
rect 10152 -3086 10186 -3070
rect 10610 -2894 10644 -2878
rect 10610 -3086 10644 -3070
rect 11068 -2894 11102 -2878
rect 11068 -3086 11102 -3070
rect 11526 -2894 11560 -2878
rect 11526 -3086 11560 -3070
rect 11984 -2894 12018 -2878
rect 11984 -3086 12018 -3070
rect 12442 -2894 12476 -2878
rect 12442 -3086 12476 -3070
rect 12900 -2894 12934 -2878
rect 12900 -3086 12934 -3070
rect 13358 -2894 13392 -2878
rect 13358 -3086 13392 -3070
rect 8898 -3154 8914 -3120
rect 9134 -3154 9150 -3120
rect 9356 -3154 9372 -3120
rect 9592 -3154 9608 -3120
rect 9814 -3154 9830 -3120
rect 10050 -3154 10066 -3120
rect 10272 -3154 10288 -3120
rect 10508 -3154 10524 -3120
rect 10730 -3154 10746 -3120
rect 10966 -3154 10982 -3120
rect 11188 -3154 11204 -3120
rect 11424 -3154 11440 -3120
rect 11646 -3154 11662 -3120
rect 11882 -3154 11898 -3120
rect 12104 -3154 12120 -3120
rect 12340 -3154 12356 -3120
rect 12562 -3154 12578 -3120
rect 12798 -3154 12814 -3120
rect 13020 -3154 13036 -3120
rect 13256 -3154 13272 -3120
rect 8352 -4148 8452 -3986
rect 18696 -4148 18796 -3986
rect 23352 -1846 23452 -1684
rect 33696 -1846 33796 -1684
rect 23898 -2176 23914 -2142
rect 24134 -2176 24150 -2142
rect 24356 -2176 24372 -2142
rect 24592 -2176 24608 -2142
rect 24814 -2176 24830 -2142
rect 25050 -2176 25066 -2142
rect 25272 -2176 25288 -2142
rect 25508 -2176 25524 -2142
rect 25730 -2176 25746 -2142
rect 25966 -2176 25982 -2142
rect 26188 -2176 26204 -2142
rect 26424 -2176 26440 -2142
rect 26646 -2176 26662 -2142
rect 26882 -2176 26898 -2142
rect 27104 -2176 27120 -2142
rect 27340 -2176 27356 -2142
rect 27562 -2176 27578 -2142
rect 27798 -2176 27814 -2142
rect 28020 -2176 28036 -2142
rect 28256 -2176 28272 -2142
rect 28898 -2176 28914 -2142
rect 29134 -2176 29150 -2142
rect 29356 -2176 29372 -2142
rect 29592 -2176 29608 -2142
rect 29814 -2176 29830 -2142
rect 30050 -2176 30066 -2142
rect 30272 -2176 30288 -2142
rect 30508 -2176 30524 -2142
rect 30730 -2176 30746 -2142
rect 30966 -2176 30982 -2142
rect 31188 -2176 31204 -2142
rect 31424 -2176 31440 -2142
rect 31646 -2176 31662 -2142
rect 31882 -2176 31898 -2142
rect 32104 -2176 32120 -2142
rect 32340 -2176 32356 -2142
rect 32562 -2176 32578 -2142
rect 32798 -2176 32814 -2142
rect 33020 -2176 33036 -2142
rect 33256 -2176 33272 -2142
rect 23778 -2226 23812 -2210
rect 23778 -2418 23812 -2402
rect 24236 -2226 24270 -2210
rect 24236 -2418 24270 -2402
rect 24694 -2226 24728 -2210
rect 24694 -2418 24728 -2402
rect 25152 -2226 25186 -2210
rect 25152 -2418 25186 -2402
rect 25610 -2226 25644 -2210
rect 25610 -2418 25644 -2402
rect 26068 -2226 26102 -2210
rect 26068 -2418 26102 -2402
rect 26526 -2226 26560 -2210
rect 26526 -2418 26560 -2402
rect 26984 -2226 27018 -2210
rect 26984 -2418 27018 -2402
rect 27442 -2226 27476 -2210
rect 27442 -2418 27476 -2402
rect 27900 -2226 27934 -2210
rect 27900 -2418 27934 -2402
rect 28358 -2226 28392 -2210
rect 28358 -2418 28392 -2402
rect 28778 -2226 28812 -2210
rect 28778 -2418 28812 -2402
rect 29236 -2226 29270 -2210
rect 29236 -2418 29270 -2402
rect 29694 -2226 29728 -2210
rect 29694 -2418 29728 -2402
rect 30152 -2226 30186 -2210
rect 30152 -2418 30186 -2402
rect 30610 -2226 30644 -2210
rect 30610 -2418 30644 -2402
rect 31068 -2226 31102 -2210
rect 31068 -2418 31102 -2402
rect 31526 -2226 31560 -2210
rect 31526 -2418 31560 -2402
rect 31984 -2226 32018 -2210
rect 31984 -2418 32018 -2402
rect 32442 -2226 32476 -2210
rect 32442 -2418 32476 -2402
rect 32900 -2226 32934 -2210
rect 32900 -2418 32934 -2402
rect 33358 -2226 33392 -2210
rect 33358 -2418 33392 -2402
rect 23898 -2486 23914 -2452
rect 24134 -2486 24150 -2452
rect 24356 -2486 24372 -2452
rect 24592 -2486 24608 -2452
rect 24814 -2486 24830 -2452
rect 25050 -2486 25066 -2452
rect 25272 -2486 25288 -2452
rect 25508 -2486 25524 -2452
rect 25730 -2486 25746 -2452
rect 25966 -2486 25982 -2452
rect 26188 -2486 26204 -2452
rect 26424 -2486 26440 -2452
rect 26646 -2486 26662 -2452
rect 26882 -2486 26898 -2452
rect 27104 -2486 27120 -2452
rect 27340 -2486 27356 -2452
rect 27562 -2486 27578 -2452
rect 27798 -2486 27814 -2452
rect 28020 -2486 28036 -2452
rect 28256 -2486 28272 -2452
rect 28898 -2486 28914 -2452
rect 29134 -2486 29150 -2452
rect 29356 -2486 29372 -2452
rect 29592 -2486 29608 -2452
rect 29814 -2486 29830 -2452
rect 30050 -2486 30066 -2452
rect 30272 -2486 30288 -2452
rect 30508 -2486 30524 -2452
rect 30730 -2486 30746 -2452
rect 30966 -2486 30982 -2452
rect 31188 -2486 31204 -2452
rect 31424 -2486 31440 -2452
rect 31646 -2486 31662 -2452
rect 31882 -2486 31898 -2452
rect 32104 -2486 32120 -2452
rect 32340 -2486 32356 -2452
rect 32562 -2486 32578 -2452
rect 32798 -2486 32814 -2452
rect 33020 -2486 33036 -2452
rect 33256 -2486 33272 -2452
rect 23898 -2844 23914 -2810
rect 24134 -2844 24150 -2810
rect 24356 -2844 24372 -2810
rect 24592 -2844 24608 -2810
rect 24814 -2844 24830 -2810
rect 25050 -2844 25066 -2810
rect 25272 -2844 25288 -2810
rect 25508 -2844 25524 -2810
rect 25730 -2844 25746 -2810
rect 25966 -2844 25982 -2810
rect 26188 -2844 26204 -2810
rect 26424 -2844 26440 -2810
rect 26646 -2844 26662 -2810
rect 26882 -2844 26898 -2810
rect 27104 -2844 27120 -2810
rect 27340 -2844 27356 -2810
rect 27562 -2844 27578 -2810
rect 27798 -2844 27814 -2810
rect 28020 -2844 28036 -2810
rect 28256 -2844 28272 -2810
rect 23778 -2894 23812 -2878
rect 23778 -3086 23812 -3070
rect 24236 -2894 24270 -2878
rect 24236 -3086 24270 -3070
rect 24694 -2894 24728 -2878
rect 24694 -3086 24728 -3070
rect 25152 -2894 25186 -2878
rect 25152 -3086 25186 -3070
rect 25610 -2894 25644 -2878
rect 25610 -3086 25644 -3070
rect 26068 -2894 26102 -2878
rect 26068 -3086 26102 -3070
rect 26526 -2894 26560 -2878
rect 26526 -3086 26560 -3070
rect 26984 -2894 27018 -2878
rect 26984 -3086 27018 -3070
rect 27442 -2894 27476 -2878
rect 27442 -3086 27476 -3070
rect 27900 -2894 27934 -2878
rect 27900 -3086 27934 -3070
rect 28358 -2894 28392 -2878
rect 28358 -3086 28392 -3070
rect 23898 -3154 23914 -3120
rect 24134 -3154 24150 -3120
rect 24356 -3154 24372 -3120
rect 24592 -3154 24608 -3120
rect 24814 -3154 24830 -3120
rect 25050 -3154 25066 -3120
rect 25272 -3154 25288 -3120
rect 25508 -3154 25524 -3120
rect 25730 -3154 25746 -3120
rect 25966 -3154 25982 -3120
rect 26188 -3154 26204 -3120
rect 26424 -3154 26440 -3120
rect 26646 -3154 26662 -3120
rect 26882 -3154 26898 -3120
rect 27104 -3154 27120 -3120
rect 27340 -3154 27356 -3120
rect 27562 -3154 27578 -3120
rect 27798 -3154 27814 -3120
rect 28020 -3154 28036 -3120
rect 28256 -3154 28272 -3120
rect 23352 -4148 23452 -3986
rect 33696 -4148 33796 -3986
rect 12306 -4770 12406 -4608
rect 22650 -4770 22750 -4608
rect 17830 -5636 17846 -5602
rect 18066 -5636 18082 -5602
rect 18288 -5636 18304 -5602
rect 18524 -5636 18540 -5602
rect 18746 -5636 18762 -5602
rect 18982 -5636 18998 -5602
rect 19204 -5636 19220 -5602
rect 19440 -5636 19456 -5602
rect 19662 -5636 19678 -5602
rect 19898 -5636 19914 -5602
rect 20120 -5636 20136 -5602
rect 20356 -5636 20372 -5602
rect 20578 -5636 20594 -5602
rect 20814 -5636 20830 -5602
rect 21036 -5636 21052 -5602
rect 21272 -5636 21288 -5602
rect 21494 -5636 21510 -5602
rect 21730 -5636 21746 -5602
rect 21952 -5636 21968 -5602
rect 22188 -5636 22204 -5602
rect 17710 -5686 17744 -5670
rect 17710 -5878 17744 -5862
rect 18168 -5686 18202 -5670
rect 18168 -5878 18202 -5862
rect 18626 -5686 18660 -5670
rect 18626 -5878 18660 -5862
rect 19084 -5686 19118 -5670
rect 19084 -5878 19118 -5862
rect 19542 -5686 19576 -5670
rect 19542 -5878 19576 -5862
rect 20000 -5686 20034 -5670
rect 20000 -5878 20034 -5862
rect 20458 -5686 20492 -5670
rect 20458 -5878 20492 -5862
rect 20916 -5686 20950 -5670
rect 20916 -5878 20950 -5862
rect 21374 -5686 21408 -5670
rect 21374 -5878 21408 -5862
rect 21832 -5686 21866 -5670
rect 21832 -5878 21866 -5862
rect 22290 -5686 22324 -5670
rect 22290 -5878 22324 -5862
rect 17830 -5946 17846 -5912
rect 18066 -5946 18082 -5912
rect 18288 -5946 18304 -5912
rect 18524 -5946 18540 -5912
rect 18746 -5946 18762 -5912
rect 18982 -5946 18998 -5912
rect 19204 -5946 19220 -5912
rect 19440 -5946 19456 -5912
rect 19662 -5946 19678 -5912
rect 19898 -5946 19914 -5912
rect 20120 -5946 20136 -5912
rect 20356 -5946 20372 -5912
rect 20578 -5946 20594 -5912
rect 20814 -5946 20830 -5912
rect 21036 -5946 21052 -5912
rect 21272 -5946 21288 -5912
rect 21494 -5946 21510 -5912
rect 21730 -5946 21746 -5912
rect 21952 -5946 21968 -5912
rect 22188 -5946 22204 -5912
rect 12830 -6304 12846 -6270
rect 13066 -6304 13082 -6270
rect 13288 -6304 13304 -6270
rect 13524 -6304 13540 -6270
rect 13746 -6304 13762 -6270
rect 13982 -6304 13998 -6270
rect 14204 -6304 14220 -6270
rect 14440 -6304 14456 -6270
rect 14662 -6304 14678 -6270
rect 14898 -6304 14914 -6270
rect 15120 -6304 15136 -6270
rect 15356 -6304 15372 -6270
rect 15578 -6304 15594 -6270
rect 15814 -6304 15830 -6270
rect 16036 -6304 16052 -6270
rect 16272 -6304 16288 -6270
rect 16494 -6304 16510 -6270
rect 16730 -6304 16746 -6270
rect 16952 -6304 16968 -6270
rect 17188 -6304 17204 -6270
rect 17830 -6304 17846 -6270
rect 18066 -6304 18082 -6270
rect 18288 -6304 18304 -6270
rect 18524 -6304 18540 -6270
rect 18746 -6304 18762 -6270
rect 18982 -6304 18998 -6270
rect 19204 -6304 19220 -6270
rect 19440 -6304 19456 -6270
rect 19662 -6304 19678 -6270
rect 19898 -6304 19914 -6270
rect 20120 -6304 20136 -6270
rect 20356 -6304 20372 -6270
rect 20578 -6304 20594 -6270
rect 20814 -6304 20830 -6270
rect 21036 -6304 21052 -6270
rect 21272 -6304 21288 -6270
rect 21494 -6304 21510 -6270
rect 21730 -6304 21746 -6270
rect 21952 -6304 21968 -6270
rect 22188 -6304 22204 -6270
rect 12710 -6354 12744 -6338
rect 12710 -6546 12744 -6530
rect 13168 -6354 13202 -6338
rect 13168 -6546 13202 -6530
rect 13626 -6354 13660 -6338
rect 13626 -6546 13660 -6530
rect 14084 -6354 14118 -6338
rect 14084 -6546 14118 -6530
rect 14542 -6354 14576 -6338
rect 14542 -6546 14576 -6530
rect 15000 -6354 15034 -6338
rect 15000 -6546 15034 -6530
rect 15458 -6354 15492 -6338
rect 15458 -6546 15492 -6530
rect 15916 -6354 15950 -6338
rect 15916 -6546 15950 -6530
rect 16374 -6354 16408 -6338
rect 16374 -6546 16408 -6530
rect 16832 -6354 16866 -6338
rect 16832 -6546 16866 -6530
rect 17290 -6354 17324 -6338
rect 17290 -6546 17324 -6530
rect 17710 -6354 17744 -6338
rect 17710 -6546 17744 -6530
rect 18168 -6354 18202 -6338
rect 18168 -6546 18202 -6530
rect 18626 -6354 18660 -6338
rect 18626 -6546 18660 -6530
rect 19084 -6354 19118 -6338
rect 19084 -6546 19118 -6530
rect 19542 -6354 19576 -6338
rect 19542 -6546 19576 -6530
rect 20000 -6354 20034 -6338
rect 20000 -6546 20034 -6530
rect 20458 -6354 20492 -6338
rect 20458 -6546 20492 -6530
rect 20916 -6354 20950 -6338
rect 20916 -6546 20950 -6530
rect 21374 -6354 21408 -6338
rect 21374 -6546 21408 -6530
rect 21832 -6354 21866 -6338
rect 21832 -6546 21866 -6530
rect 22290 -6354 22324 -6338
rect 22290 -6546 22324 -6530
rect 12830 -6614 12846 -6580
rect 13066 -6614 13082 -6580
rect 13288 -6614 13304 -6580
rect 13524 -6614 13540 -6580
rect 13746 -6614 13762 -6580
rect 13982 -6614 13998 -6580
rect 14204 -6614 14220 -6580
rect 14440 -6614 14456 -6580
rect 14662 -6614 14678 -6580
rect 14898 -6614 14914 -6580
rect 15120 -6614 15136 -6580
rect 15356 -6614 15372 -6580
rect 15578 -6614 15594 -6580
rect 15814 -6614 15830 -6580
rect 16036 -6614 16052 -6580
rect 16272 -6614 16288 -6580
rect 16494 -6614 16510 -6580
rect 16730 -6614 16746 -6580
rect 16952 -6614 16968 -6580
rect 17188 -6614 17204 -6580
rect 17830 -6614 17846 -6580
rect 18066 -6614 18082 -6580
rect 18288 -6614 18304 -6580
rect 18524 -6614 18540 -6580
rect 18746 -6614 18762 -6580
rect 18982 -6614 18998 -6580
rect 19204 -6614 19220 -6580
rect 19440 -6614 19456 -6580
rect 19662 -6614 19678 -6580
rect 19898 -6614 19914 -6580
rect 20120 -6614 20136 -6580
rect 20356 -6614 20372 -6580
rect 20578 -6614 20594 -6580
rect 20814 -6614 20830 -6580
rect 21036 -6614 21052 -6580
rect 21272 -6614 21288 -6580
rect 21494 -6614 21510 -6580
rect 21730 -6614 21746 -6580
rect 21952 -6614 21968 -6580
rect 22188 -6614 22204 -6580
rect 12306 -7072 12406 -6910
rect 22650 -7072 22750 -6910
rect 27306 -4770 27406 -4608
rect 37650 -4770 37750 -4608
rect 32830 -5636 32846 -5602
rect 33066 -5636 33082 -5602
rect 33288 -5636 33304 -5602
rect 33524 -5636 33540 -5602
rect 33746 -5636 33762 -5602
rect 33982 -5636 33998 -5602
rect 34204 -5636 34220 -5602
rect 34440 -5636 34456 -5602
rect 34662 -5636 34678 -5602
rect 34898 -5636 34914 -5602
rect 35120 -5636 35136 -5602
rect 35356 -5636 35372 -5602
rect 35578 -5636 35594 -5602
rect 35814 -5636 35830 -5602
rect 36036 -5636 36052 -5602
rect 36272 -5636 36288 -5602
rect 36494 -5636 36510 -5602
rect 36730 -5636 36746 -5602
rect 36952 -5636 36968 -5602
rect 37188 -5636 37204 -5602
rect 32710 -5686 32744 -5670
rect 32710 -5878 32744 -5862
rect 33168 -5686 33202 -5670
rect 33168 -5878 33202 -5862
rect 33626 -5686 33660 -5670
rect 33626 -5878 33660 -5862
rect 34084 -5686 34118 -5670
rect 34084 -5878 34118 -5862
rect 34542 -5686 34576 -5670
rect 34542 -5878 34576 -5862
rect 35000 -5686 35034 -5670
rect 35000 -5878 35034 -5862
rect 35458 -5686 35492 -5670
rect 35458 -5878 35492 -5862
rect 35916 -5686 35950 -5670
rect 35916 -5878 35950 -5862
rect 36374 -5686 36408 -5670
rect 36374 -5878 36408 -5862
rect 36832 -5686 36866 -5670
rect 36832 -5878 36866 -5862
rect 37290 -5686 37324 -5670
rect 37290 -5878 37324 -5862
rect 32830 -5946 32846 -5912
rect 33066 -5946 33082 -5912
rect 33288 -5946 33304 -5912
rect 33524 -5946 33540 -5912
rect 33746 -5946 33762 -5912
rect 33982 -5946 33998 -5912
rect 34204 -5946 34220 -5912
rect 34440 -5946 34456 -5912
rect 34662 -5946 34678 -5912
rect 34898 -5946 34914 -5912
rect 35120 -5946 35136 -5912
rect 35356 -5946 35372 -5912
rect 35578 -5946 35594 -5912
rect 35814 -5946 35830 -5912
rect 36036 -5946 36052 -5912
rect 36272 -5946 36288 -5912
rect 36494 -5946 36510 -5912
rect 36730 -5946 36746 -5912
rect 36952 -5946 36968 -5912
rect 37188 -5946 37204 -5912
rect 27830 -6304 27846 -6270
rect 28066 -6304 28082 -6270
rect 28288 -6304 28304 -6270
rect 28524 -6304 28540 -6270
rect 28746 -6304 28762 -6270
rect 28982 -6304 28998 -6270
rect 29204 -6304 29220 -6270
rect 29440 -6304 29456 -6270
rect 29662 -6304 29678 -6270
rect 29898 -6304 29914 -6270
rect 30120 -6304 30136 -6270
rect 30356 -6304 30372 -6270
rect 30578 -6304 30594 -6270
rect 30814 -6304 30830 -6270
rect 31036 -6304 31052 -6270
rect 31272 -6304 31288 -6270
rect 31494 -6304 31510 -6270
rect 31730 -6304 31746 -6270
rect 31952 -6304 31968 -6270
rect 32188 -6304 32204 -6270
rect 32830 -6304 32846 -6270
rect 33066 -6304 33082 -6270
rect 33288 -6304 33304 -6270
rect 33524 -6304 33540 -6270
rect 33746 -6304 33762 -6270
rect 33982 -6304 33998 -6270
rect 34204 -6304 34220 -6270
rect 34440 -6304 34456 -6270
rect 34662 -6304 34678 -6270
rect 34898 -6304 34914 -6270
rect 35120 -6304 35136 -6270
rect 35356 -6304 35372 -6270
rect 35578 -6304 35594 -6270
rect 35814 -6304 35830 -6270
rect 36036 -6304 36052 -6270
rect 36272 -6304 36288 -6270
rect 36494 -6304 36510 -6270
rect 36730 -6304 36746 -6270
rect 36952 -6304 36968 -6270
rect 37188 -6304 37204 -6270
rect 27710 -6354 27744 -6338
rect 27710 -6546 27744 -6530
rect 28168 -6354 28202 -6338
rect 28168 -6546 28202 -6530
rect 28626 -6354 28660 -6338
rect 28626 -6546 28660 -6530
rect 29084 -6354 29118 -6338
rect 29084 -6546 29118 -6530
rect 29542 -6354 29576 -6338
rect 29542 -6546 29576 -6530
rect 30000 -6354 30034 -6338
rect 30000 -6546 30034 -6530
rect 30458 -6354 30492 -6338
rect 30458 -6546 30492 -6530
rect 30916 -6354 30950 -6338
rect 30916 -6546 30950 -6530
rect 31374 -6354 31408 -6338
rect 31374 -6546 31408 -6530
rect 31832 -6354 31866 -6338
rect 31832 -6546 31866 -6530
rect 32290 -6354 32324 -6338
rect 32290 -6546 32324 -6530
rect 32710 -6354 32744 -6338
rect 32710 -6546 32744 -6530
rect 33168 -6354 33202 -6338
rect 33168 -6546 33202 -6530
rect 33626 -6354 33660 -6338
rect 33626 -6546 33660 -6530
rect 34084 -6354 34118 -6338
rect 34084 -6546 34118 -6530
rect 34542 -6354 34576 -6338
rect 34542 -6546 34576 -6530
rect 35000 -6354 35034 -6338
rect 35000 -6546 35034 -6530
rect 35458 -6354 35492 -6338
rect 35458 -6546 35492 -6530
rect 35916 -6354 35950 -6338
rect 35916 -6546 35950 -6530
rect 36374 -6354 36408 -6338
rect 36374 -6546 36408 -6530
rect 36832 -6354 36866 -6338
rect 36832 -6546 36866 -6530
rect 37290 -6354 37324 -6338
rect 37290 -6546 37324 -6530
rect 27830 -6614 27846 -6580
rect 28066 -6614 28082 -6580
rect 28288 -6614 28304 -6580
rect 28524 -6614 28540 -6580
rect 28746 -6614 28762 -6580
rect 28982 -6614 28998 -6580
rect 29204 -6614 29220 -6580
rect 29440 -6614 29456 -6580
rect 29662 -6614 29678 -6580
rect 29898 -6614 29914 -6580
rect 30120 -6614 30136 -6580
rect 30356 -6614 30372 -6580
rect 30578 -6614 30594 -6580
rect 30814 -6614 30830 -6580
rect 31036 -6614 31052 -6580
rect 31272 -6614 31288 -6580
rect 31494 -6614 31510 -6580
rect 31730 -6614 31746 -6580
rect 31952 -6614 31968 -6580
rect 32188 -6614 32204 -6580
rect 32830 -6614 32846 -6580
rect 33066 -6614 33082 -6580
rect 33288 -6614 33304 -6580
rect 33524 -6614 33540 -6580
rect 33746 -6614 33762 -6580
rect 33982 -6614 33998 -6580
rect 34204 -6614 34220 -6580
rect 34440 -6614 34456 -6580
rect 34662 -6614 34678 -6580
rect 34898 -6614 34914 -6580
rect 35120 -6614 35136 -6580
rect 35356 -6614 35372 -6580
rect 35578 -6614 35594 -6580
rect 35814 -6614 35830 -6580
rect 36036 -6614 36052 -6580
rect 36272 -6614 36288 -6580
rect 36494 -6614 36510 -6580
rect 36730 -6614 36746 -6580
rect 36952 -6614 36968 -6580
rect 37188 -6614 37204 -6580
rect 27306 -7072 27406 -6910
rect 37650 -7072 37750 -6910
rect 12306 -7470 12406 -7308
rect 22650 -7470 22750 -7308
rect 12829 -7788 12845 -7754
rect 13065 -7788 13081 -7754
rect 13287 -7788 13303 -7754
rect 13523 -7788 13539 -7754
rect 13745 -7788 13761 -7754
rect 13981 -7788 13997 -7754
rect 14203 -7788 14219 -7754
rect 14439 -7788 14455 -7754
rect 14661 -7788 14677 -7754
rect 14897 -7788 14913 -7754
rect 15119 -7788 15135 -7754
rect 15355 -7788 15371 -7754
rect 15577 -7788 15593 -7754
rect 15813 -7788 15829 -7754
rect 16035 -7788 16051 -7754
rect 16271 -7788 16287 -7754
rect 16493 -7788 16509 -7754
rect 16729 -7788 16745 -7754
rect 16951 -7788 16967 -7754
rect 17187 -7788 17203 -7754
rect 17829 -7788 17845 -7754
rect 18065 -7788 18081 -7754
rect 18287 -7788 18303 -7754
rect 18523 -7788 18539 -7754
rect 18745 -7788 18761 -7754
rect 18981 -7788 18997 -7754
rect 19203 -7788 19219 -7754
rect 19439 -7788 19455 -7754
rect 19661 -7788 19677 -7754
rect 19897 -7788 19913 -7754
rect 20119 -7788 20135 -7754
rect 20355 -7788 20371 -7754
rect 20577 -7788 20593 -7754
rect 20813 -7788 20829 -7754
rect 21035 -7788 21051 -7754
rect 21271 -7788 21287 -7754
rect 21493 -7788 21509 -7754
rect 21729 -7788 21745 -7754
rect 21951 -7788 21967 -7754
rect 22187 -7788 22203 -7754
rect 12709 -7847 12743 -7831
rect 12709 -9039 12743 -9023
rect 13167 -7847 13201 -7831
rect 13167 -9039 13201 -9023
rect 13625 -7847 13659 -7831
rect 13625 -9039 13659 -9023
rect 14083 -7847 14117 -7831
rect 14083 -9039 14117 -9023
rect 14541 -7847 14575 -7831
rect 14541 -9039 14575 -9023
rect 14999 -7847 15033 -7831
rect 14999 -9039 15033 -9023
rect 15457 -7847 15491 -7831
rect 15457 -9039 15491 -9023
rect 15915 -7847 15949 -7831
rect 15915 -9039 15949 -9023
rect 16373 -7847 16407 -7831
rect 16373 -9039 16407 -9023
rect 16831 -7847 16865 -7831
rect 16831 -9039 16865 -9023
rect 17289 -7847 17323 -7831
rect 17289 -9039 17323 -9023
rect 17709 -7847 17743 -7831
rect 17709 -9039 17743 -9023
rect 18167 -7847 18201 -7831
rect 18167 -9039 18201 -9023
rect 18625 -7847 18659 -7831
rect 18625 -9039 18659 -9023
rect 19083 -7847 19117 -7831
rect 19083 -9039 19117 -9023
rect 19541 -7847 19575 -7831
rect 19541 -9039 19575 -9023
rect 19999 -7847 20033 -7831
rect 19999 -9039 20033 -9023
rect 20457 -7847 20491 -7831
rect 20457 -9039 20491 -9023
rect 20915 -7847 20949 -7831
rect 20915 -9039 20949 -9023
rect 21373 -7847 21407 -7831
rect 21373 -9039 21407 -9023
rect 21831 -7847 21865 -7831
rect 21831 -9039 21865 -9023
rect 22289 -7847 22323 -7831
rect 22289 -9039 22323 -9023
rect 12829 -9116 12845 -9082
rect 13065 -9116 13081 -9082
rect 13287 -9116 13303 -9082
rect 13523 -9116 13539 -9082
rect 13745 -9116 13761 -9082
rect 13981 -9116 13997 -9082
rect 14203 -9116 14219 -9082
rect 14439 -9116 14455 -9082
rect 14661 -9116 14677 -9082
rect 14897 -9116 14913 -9082
rect 15119 -9116 15135 -9082
rect 15355 -9116 15371 -9082
rect 15577 -9116 15593 -9082
rect 15813 -9116 15829 -9082
rect 16035 -9116 16051 -9082
rect 16271 -9116 16287 -9082
rect 16493 -9116 16509 -9082
rect 16729 -9116 16745 -9082
rect 16951 -9116 16967 -9082
rect 17187 -9116 17203 -9082
rect 17829 -9116 17845 -9082
rect 18065 -9116 18081 -9082
rect 18287 -9116 18303 -9082
rect 18523 -9116 18539 -9082
rect 18745 -9116 18761 -9082
rect 18981 -9116 18997 -9082
rect 19203 -9116 19219 -9082
rect 19439 -9116 19455 -9082
rect 19661 -9116 19677 -9082
rect 19897 -9116 19913 -9082
rect 20119 -9116 20135 -9082
rect 20355 -9116 20371 -9082
rect 20577 -9116 20593 -9082
rect 20813 -9116 20829 -9082
rect 21035 -9116 21051 -9082
rect 21271 -9116 21287 -9082
rect 21493 -9116 21509 -9082
rect 21729 -9116 21745 -9082
rect 21951 -9116 21967 -9082
rect 22187 -9116 22203 -9082
rect 17426 -9888 17886 -9882
rect 17426 -9936 17832 -9888
rect 17880 -9936 17886 -9888
rect 17426 -9942 17886 -9936
rect 13606 -10053 13622 -10019
rect 13842 -10053 13858 -10019
rect 14064 -10053 14080 -10019
rect 14300 -10053 14316 -10019
rect 14522 -10053 14538 -10019
rect 14758 -10053 14774 -10019
rect 14980 -10053 14996 -10019
rect 15216 -10053 15232 -10019
rect 15438 -10053 15454 -10019
rect 15674 -10053 15690 -10019
rect 15896 -10053 15912 -10019
rect 16132 -10053 16148 -10019
rect 16354 -10053 16370 -10019
rect 16590 -10053 16606 -10019
rect 16812 -10053 16828 -10019
rect 17048 -10053 17064 -10019
rect 17270 -10053 17286 -10019
rect 17506 -10053 17522 -10019
rect 17728 -10053 17744 -10019
rect 17964 -10053 17980 -10019
rect 18186 -10053 18202 -10019
rect 18422 -10053 18438 -10019
rect 18644 -10053 18660 -10019
rect 18880 -10053 18896 -10019
rect 19102 -10053 19118 -10019
rect 19338 -10053 19354 -10019
rect 19560 -10053 19576 -10019
rect 19796 -10053 19812 -10019
rect 20018 -10053 20034 -10019
rect 20254 -10053 20270 -10019
rect 20476 -10053 20492 -10019
rect 20712 -10053 20728 -10019
rect 20934 -10053 20950 -10019
rect 21170 -10053 21186 -10019
rect 21392 -10053 21408 -10019
rect 21628 -10053 21644 -10019
rect 13486 -10112 13520 -10096
rect 13486 -11704 13520 -11688
rect 13944 -10112 13978 -10096
rect 13944 -11704 13978 -11688
rect 14402 -10112 14436 -10096
rect 14402 -11704 14436 -11688
rect 14860 -10112 14894 -10096
rect 14860 -11704 14894 -11688
rect 15318 -10112 15352 -10096
rect 15318 -11704 15352 -11688
rect 15776 -10112 15810 -10096
rect 15776 -11704 15810 -11688
rect 16234 -10112 16268 -10096
rect 16234 -11704 16268 -11688
rect 16692 -10112 16726 -10096
rect 16692 -11704 16726 -11688
rect 17150 -10112 17184 -10096
rect 17150 -11704 17184 -11688
rect 17608 -10112 17642 -10096
rect 17608 -11704 17642 -11688
rect 18066 -10112 18100 -10096
rect 18066 -11704 18100 -11688
rect 18524 -10112 18558 -10096
rect 18524 -11704 18558 -11688
rect 18982 -10112 19016 -10096
rect 18982 -11704 19016 -11688
rect 19440 -10112 19474 -10096
rect 19440 -11704 19474 -11688
rect 19898 -10112 19932 -10096
rect 19898 -11704 19932 -11688
rect 20356 -10112 20390 -10096
rect 20356 -11704 20390 -11688
rect 20814 -10112 20848 -10096
rect 20814 -11704 20848 -11688
rect 21272 -10112 21306 -10096
rect 21272 -11704 21306 -11688
rect 21730 -10112 21764 -10096
rect 21730 -11704 21764 -11688
rect 13606 -11781 13622 -11747
rect 13842 -11781 13858 -11747
rect 14064 -11781 14080 -11747
rect 14300 -11781 14316 -11747
rect 14522 -11781 14538 -11747
rect 14758 -11781 14774 -11747
rect 14980 -11781 14996 -11747
rect 15216 -11781 15232 -11747
rect 15438 -11781 15454 -11747
rect 15674 -11781 15690 -11747
rect 15896 -11781 15912 -11747
rect 16132 -11781 16148 -11747
rect 16354 -11781 16370 -11747
rect 16590 -11781 16606 -11747
rect 16812 -11781 16828 -11747
rect 17048 -11781 17064 -11747
rect 17270 -11781 17286 -11747
rect 17506 -11781 17522 -11747
rect 17728 -11781 17744 -11747
rect 17964 -11781 17980 -11747
rect 18186 -11781 18202 -11747
rect 18422 -11781 18438 -11747
rect 18644 -11781 18660 -11747
rect 18880 -11781 18896 -11747
rect 19102 -11781 19118 -11747
rect 19338 -11781 19354 -11747
rect 19560 -11781 19576 -11747
rect 19796 -11781 19812 -11747
rect 20018 -11781 20034 -11747
rect 20254 -11781 20270 -11747
rect 20476 -11781 20492 -11747
rect 20712 -11781 20728 -11747
rect 20934 -11781 20950 -11747
rect 21170 -11781 21186 -11747
rect 21392 -11781 21408 -11747
rect 21628 -11781 21644 -11747
rect 12306 -13152 12406 -12990
rect 22650 -13152 22750 -12990
rect 27306 -7470 27406 -7308
rect 37650 -7470 37750 -7308
rect 27829 -7788 27845 -7754
rect 28065 -7788 28081 -7754
rect 28287 -7788 28303 -7754
rect 28523 -7788 28539 -7754
rect 28745 -7788 28761 -7754
rect 28981 -7788 28997 -7754
rect 29203 -7788 29219 -7754
rect 29439 -7788 29455 -7754
rect 29661 -7788 29677 -7754
rect 29897 -7788 29913 -7754
rect 30119 -7788 30135 -7754
rect 30355 -7788 30371 -7754
rect 30577 -7788 30593 -7754
rect 30813 -7788 30829 -7754
rect 31035 -7788 31051 -7754
rect 31271 -7788 31287 -7754
rect 31493 -7788 31509 -7754
rect 31729 -7788 31745 -7754
rect 31951 -7788 31967 -7754
rect 32187 -7788 32203 -7754
rect 32829 -7788 32845 -7754
rect 33065 -7788 33081 -7754
rect 33287 -7788 33303 -7754
rect 33523 -7788 33539 -7754
rect 33745 -7788 33761 -7754
rect 33981 -7788 33997 -7754
rect 34203 -7788 34219 -7754
rect 34439 -7788 34455 -7754
rect 34661 -7788 34677 -7754
rect 34897 -7788 34913 -7754
rect 35119 -7788 35135 -7754
rect 35355 -7788 35371 -7754
rect 35577 -7788 35593 -7754
rect 35813 -7788 35829 -7754
rect 36035 -7788 36051 -7754
rect 36271 -7788 36287 -7754
rect 36493 -7788 36509 -7754
rect 36729 -7788 36745 -7754
rect 36951 -7788 36967 -7754
rect 37187 -7788 37203 -7754
rect 27709 -7847 27743 -7831
rect 27709 -9039 27743 -9023
rect 28167 -7847 28201 -7831
rect 28167 -9039 28201 -9023
rect 28625 -7847 28659 -7831
rect 28625 -9039 28659 -9023
rect 29083 -7847 29117 -7831
rect 29083 -9039 29117 -9023
rect 29541 -7847 29575 -7831
rect 29541 -9039 29575 -9023
rect 29999 -7847 30033 -7831
rect 29999 -9039 30033 -9023
rect 30457 -7847 30491 -7831
rect 30457 -9039 30491 -9023
rect 30915 -7847 30949 -7831
rect 30915 -9039 30949 -9023
rect 31373 -7847 31407 -7831
rect 31373 -9039 31407 -9023
rect 31831 -7847 31865 -7831
rect 31831 -9039 31865 -9023
rect 32289 -7847 32323 -7831
rect 32289 -9039 32323 -9023
rect 32709 -7847 32743 -7831
rect 32709 -9039 32743 -9023
rect 33167 -7847 33201 -7831
rect 33167 -9039 33201 -9023
rect 33625 -7847 33659 -7831
rect 33625 -9039 33659 -9023
rect 34083 -7847 34117 -7831
rect 34083 -9039 34117 -9023
rect 34541 -7847 34575 -7831
rect 34541 -9039 34575 -9023
rect 34999 -7847 35033 -7831
rect 34999 -9039 35033 -9023
rect 35457 -7847 35491 -7831
rect 35457 -9039 35491 -9023
rect 35915 -7847 35949 -7831
rect 35915 -9039 35949 -9023
rect 36373 -7847 36407 -7831
rect 36373 -9039 36407 -9023
rect 36831 -7847 36865 -7831
rect 36831 -9039 36865 -9023
rect 37289 -7847 37323 -7831
rect 37289 -9039 37323 -9023
rect 27829 -9116 27845 -9082
rect 28065 -9116 28081 -9082
rect 28287 -9116 28303 -9082
rect 28523 -9116 28539 -9082
rect 28745 -9116 28761 -9082
rect 28981 -9116 28997 -9082
rect 29203 -9116 29219 -9082
rect 29439 -9116 29455 -9082
rect 29661 -9116 29677 -9082
rect 29897 -9116 29913 -9082
rect 30119 -9116 30135 -9082
rect 30355 -9116 30371 -9082
rect 30577 -9116 30593 -9082
rect 30813 -9116 30829 -9082
rect 31035 -9116 31051 -9082
rect 31271 -9116 31287 -9082
rect 31493 -9116 31509 -9082
rect 31729 -9116 31745 -9082
rect 31951 -9116 31967 -9082
rect 32187 -9116 32203 -9082
rect 32829 -9116 32845 -9082
rect 33065 -9116 33081 -9082
rect 33287 -9116 33303 -9082
rect 33523 -9116 33539 -9082
rect 33745 -9116 33761 -9082
rect 33981 -9116 33997 -9082
rect 34203 -9116 34219 -9082
rect 34439 -9116 34455 -9082
rect 34661 -9116 34677 -9082
rect 34897 -9116 34913 -9082
rect 35119 -9116 35135 -9082
rect 35355 -9116 35371 -9082
rect 35577 -9116 35593 -9082
rect 35813 -9116 35829 -9082
rect 36035 -9116 36051 -9082
rect 36271 -9116 36287 -9082
rect 36493 -9116 36509 -9082
rect 36729 -9116 36745 -9082
rect 36951 -9116 36967 -9082
rect 37187 -9116 37203 -9082
rect 32426 -9888 32886 -9882
rect 32426 -9936 32832 -9888
rect 32880 -9936 32886 -9888
rect 32426 -9942 32886 -9936
rect 28606 -10053 28622 -10019
rect 28842 -10053 28858 -10019
rect 29064 -10053 29080 -10019
rect 29300 -10053 29316 -10019
rect 29522 -10053 29538 -10019
rect 29758 -10053 29774 -10019
rect 29980 -10053 29996 -10019
rect 30216 -10053 30232 -10019
rect 30438 -10053 30454 -10019
rect 30674 -10053 30690 -10019
rect 30896 -10053 30912 -10019
rect 31132 -10053 31148 -10019
rect 31354 -10053 31370 -10019
rect 31590 -10053 31606 -10019
rect 31812 -10053 31828 -10019
rect 32048 -10053 32064 -10019
rect 32270 -10053 32286 -10019
rect 32506 -10053 32522 -10019
rect 32728 -10053 32744 -10019
rect 32964 -10053 32980 -10019
rect 33186 -10053 33202 -10019
rect 33422 -10053 33438 -10019
rect 33644 -10053 33660 -10019
rect 33880 -10053 33896 -10019
rect 34102 -10053 34118 -10019
rect 34338 -10053 34354 -10019
rect 34560 -10053 34576 -10019
rect 34796 -10053 34812 -10019
rect 35018 -10053 35034 -10019
rect 35254 -10053 35270 -10019
rect 35476 -10053 35492 -10019
rect 35712 -10053 35728 -10019
rect 35934 -10053 35950 -10019
rect 36170 -10053 36186 -10019
rect 36392 -10053 36408 -10019
rect 36628 -10053 36644 -10019
rect 28486 -10112 28520 -10096
rect 28486 -11704 28520 -11688
rect 28944 -10112 28978 -10096
rect 28944 -11704 28978 -11688
rect 29402 -10112 29436 -10096
rect 29402 -11704 29436 -11688
rect 29860 -10112 29894 -10096
rect 29860 -11704 29894 -11688
rect 30318 -10112 30352 -10096
rect 30318 -11704 30352 -11688
rect 30776 -10112 30810 -10096
rect 30776 -11704 30810 -11688
rect 31234 -10112 31268 -10096
rect 31234 -11704 31268 -11688
rect 31692 -10112 31726 -10096
rect 31692 -11704 31726 -11688
rect 32150 -10112 32184 -10096
rect 32150 -11704 32184 -11688
rect 32608 -10112 32642 -10096
rect 32608 -11704 32642 -11688
rect 33066 -10112 33100 -10096
rect 33066 -11704 33100 -11688
rect 33524 -10112 33558 -10096
rect 33524 -11704 33558 -11688
rect 33982 -10112 34016 -10096
rect 33982 -11704 34016 -11688
rect 34440 -10112 34474 -10096
rect 34440 -11704 34474 -11688
rect 34898 -10112 34932 -10096
rect 34898 -11704 34932 -11688
rect 35356 -10112 35390 -10096
rect 35356 -11704 35390 -11688
rect 35814 -10112 35848 -10096
rect 35814 -11704 35848 -11688
rect 36272 -10112 36306 -10096
rect 36272 -11704 36306 -11688
rect 36730 -10112 36764 -10096
rect 36730 -11704 36764 -11688
rect 28606 -11781 28622 -11747
rect 28842 -11781 28858 -11747
rect 29064 -11781 29080 -11747
rect 29300 -11781 29316 -11747
rect 29522 -11781 29538 -11747
rect 29758 -11781 29774 -11747
rect 29980 -11781 29996 -11747
rect 30216 -11781 30232 -11747
rect 30438 -11781 30454 -11747
rect 30674 -11781 30690 -11747
rect 30896 -11781 30912 -11747
rect 31132 -11781 31148 -11747
rect 31354 -11781 31370 -11747
rect 31590 -11781 31606 -11747
rect 31812 -11781 31828 -11747
rect 32048 -11781 32064 -11747
rect 32270 -11781 32286 -11747
rect 32506 -11781 32522 -11747
rect 32728 -11781 32744 -11747
rect 32964 -11781 32980 -11747
rect 33186 -11781 33202 -11747
rect 33422 -11781 33438 -11747
rect 33644 -11781 33660 -11747
rect 33880 -11781 33896 -11747
rect 34102 -11781 34118 -11747
rect 34338 -11781 34354 -11747
rect 34560 -11781 34576 -11747
rect 34796 -11781 34812 -11747
rect 35018 -11781 35034 -11747
rect 35254 -11781 35270 -11747
rect 35476 -11781 35492 -11747
rect 35712 -11781 35728 -11747
rect 35934 -11781 35950 -11747
rect 36170 -11781 36186 -11747
rect 36392 -11781 36408 -11747
rect 36628 -11781 36644 -11747
rect 27306 -13152 27406 -12990
rect 37650 -13152 37750 -12990
rect 8352 -13766 8452 -13604
rect 18696 -13766 18796 -13604
rect 9458 -15009 9474 -14975
rect 9694 -15009 9710 -14975
rect 9916 -15009 9932 -14975
rect 10152 -15009 10168 -14975
rect 10374 -15009 10390 -14975
rect 10610 -15009 10626 -14975
rect 10832 -15009 10848 -14975
rect 11068 -15009 11084 -14975
rect 11290 -15009 11306 -14975
rect 11526 -15009 11542 -14975
rect 11748 -15009 11764 -14975
rect 11984 -15009 12000 -14975
rect 12206 -15009 12222 -14975
rect 12442 -15009 12458 -14975
rect 12664 -15009 12680 -14975
rect 12900 -15009 12916 -14975
rect 13122 -15009 13138 -14975
rect 13358 -15009 13374 -14975
rect 13580 -15009 13596 -14975
rect 13816 -15009 13832 -14975
rect 14038 -15009 14054 -14975
rect 14274 -15009 14290 -14975
rect 14496 -15009 14512 -14975
rect 14732 -15009 14748 -14975
rect 14954 -15009 14970 -14975
rect 15190 -15009 15206 -14975
rect 15412 -15009 15428 -14975
rect 15648 -15009 15664 -14975
rect 15870 -15009 15886 -14975
rect 16106 -15009 16122 -14975
rect 16328 -15009 16344 -14975
rect 16564 -15009 16580 -14975
rect 16786 -15009 16802 -14975
rect 17022 -15009 17038 -14975
rect 17244 -15009 17260 -14975
rect 17480 -15009 17496 -14975
rect 9338 -15068 9372 -15052
rect 9338 -16660 9372 -16644
rect 9796 -15068 9830 -15052
rect 9796 -16660 9830 -16644
rect 10254 -15068 10288 -15052
rect 10254 -16660 10288 -16644
rect 10712 -15068 10746 -15052
rect 10712 -16660 10746 -16644
rect 11170 -15068 11204 -15052
rect 11170 -16660 11204 -16644
rect 11628 -15068 11662 -15052
rect 11628 -16660 11662 -16644
rect 12086 -15068 12120 -15052
rect 12086 -16660 12120 -16644
rect 12544 -15068 12578 -15052
rect 12544 -16660 12578 -16644
rect 13002 -15068 13036 -15052
rect 13002 -16660 13036 -16644
rect 13460 -15068 13494 -15052
rect 13460 -16660 13494 -16644
rect 13918 -15068 13952 -15052
rect 13918 -16660 13952 -16644
rect 14376 -15068 14410 -15052
rect 14376 -16660 14410 -16644
rect 14834 -15068 14868 -15052
rect 14834 -16660 14868 -16644
rect 15292 -15068 15326 -15052
rect 15292 -16660 15326 -16644
rect 15750 -15068 15784 -15052
rect 15750 -16660 15784 -16644
rect 16208 -15068 16242 -15052
rect 16208 -16660 16242 -16644
rect 16666 -15068 16700 -15052
rect 16666 -16660 16700 -16644
rect 17124 -15068 17158 -15052
rect 17124 -16660 17158 -16644
rect 17582 -15068 17616 -15052
rect 17582 -16660 17616 -16644
rect 9458 -16737 9474 -16703
rect 9694 -16737 9710 -16703
rect 9916 -16737 9932 -16703
rect 10152 -16737 10168 -16703
rect 10374 -16737 10390 -16703
rect 10610 -16737 10626 -16703
rect 10832 -16737 10848 -16703
rect 11068 -16737 11084 -16703
rect 11290 -16737 11306 -16703
rect 11526 -16737 11542 -16703
rect 11748 -16737 11764 -16703
rect 11984 -16737 12000 -16703
rect 12206 -16737 12222 -16703
rect 12442 -16737 12458 -16703
rect 12664 -16737 12680 -16703
rect 12900 -16737 12916 -16703
rect 13122 -16737 13138 -16703
rect 13358 -16737 13374 -16703
rect 13580 -16737 13596 -16703
rect 13816 -16737 13832 -16703
rect 14038 -16737 14054 -16703
rect 14274 -16737 14290 -16703
rect 14496 -16737 14512 -16703
rect 14732 -16737 14748 -16703
rect 14954 -16737 14970 -16703
rect 15190 -16737 15206 -16703
rect 15412 -16737 15428 -16703
rect 15648 -16737 15664 -16703
rect 15870 -16737 15886 -16703
rect 16106 -16737 16122 -16703
rect 16328 -16737 16344 -16703
rect 16564 -16737 16580 -16703
rect 16786 -16737 16802 -16703
rect 17022 -16737 17038 -16703
rect 17244 -16737 17260 -16703
rect 17480 -16737 17496 -16703
rect 13216 -16820 13676 -16814
rect 13216 -16868 13222 -16820
rect 13270 -16868 13676 -16820
rect 13216 -16874 13676 -16868
rect 8899 -17674 8915 -17640
rect 9135 -17674 9151 -17640
rect 9357 -17674 9373 -17640
rect 9593 -17674 9609 -17640
rect 9815 -17674 9831 -17640
rect 10051 -17674 10067 -17640
rect 10273 -17674 10289 -17640
rect 10509 -17674 10525 -17640
rect 10731 -17674 10747 -17640
rect 10967 -17674 10983 -17640
rect 11189 -17674 11205 -17640
rect 11425 -17674 11441 -17640
rect 11647 -17674 11663 -17640
rect 11883 -17674 11899 -17640
rect 12105 -17674 12121 -17640
rect 12341 -17674 12357 -17640
rect 12563 -17674 12579 -17640
rect 12799 -17674 12815 -17640
rect 13021 -17674 13037 -17640
rect 13257 -17674 13273 -17640
rect 13899 -17674 13915 -17640
rect 14135 -17674 14151 -17640
rect 14357 -17674 14373 -17640
rect 14593 -17674 14609 -17640
rect 14815 -17674 14831 -17640
rect 15051 -17674 15067 -17640
rect 15273 -17674 15289 -17640
rect 15509 -17674 15525 -17640
rect 15731 -17674 15747 -17640
rect 15967 -17674 15983 -17640
rect 16189 -17674 16205 -17640
rect 16425 -17674 16441 -17640
rect 16647 -17674 16663 -17640
rect 16883 -17674 16899 -17640
rect 17105 -17674 17121 -17640
rect 17341 -17674 17357 -17640
rect 17563 -17674 17579 -17640
rect 17799 -17674 17815 -17640
rect 18021 -17674 18037 -17640
rect 18257 -17674 18273 -17640
rect 8779 -17733 8813 -17717
rect 8779 -18925 8813 -18909
rect 9237 -17733 9271 -17717
rect 9237 -18925 9271 -18909
rect 9695 -17733 9729 -17717
rect 9695 -18925 9729 -18909
rect 10153 -17733 10187 -17717
rect 10153 -18925 10187 -18909
rect 10611 -17733 10645 -17717
rect 10611 -18925 10645 -18909
rect 11069 -17733 11103 -17717
rect 11069 -18925 11103 -18909
rect 11527 -17733 11561 -17717
rect 11527 -18925 11561 -18909
rect 11985 -17733 12019 -17717
rect 11985 -18925 12019 -18909
rect 12443 -17733 12477 -17717
rect 12443 -18925 12477 -18909
rect 12901 -17733 12935 -17717
rect 12901 -18925 12935 -18909
rect 13359 -17733 13393 -17717
rect 13359 -18925 13393 -18909
rect 13779 -17733 13813 -17717
rect 13779 -18925 13813 -18909
rect 14237 -17733 14271 -17717
rect 14237 -18925 14271 -18909
rect 14695 -17733 14729 -17717
rect 14695 -18925 14729 -18909
rect 15153 -17733 15187 -17717
rect 15153 -18925 15187 -18909
rect 15611 -17733 15645 -17717
rect 15611 -18925 15645 -18909
rect 16069 -17733 16103 -17717
rect 16069 -18925 16103 -18909
rect 16527 -17733 16561 -17717
rect 16527 -18925 16561 -18909
rect 16985 -17733 17019 -17717
rect 16985 -18925 17019 -18909
rect 17443 -17733 17477 -17717
rect 17443 -18925 17477 -18909
rect 17901 -17733 17935 -17717
rect 17901 -18925 17935 -18909
rect 18359 -17733 18393 -17717
rect 18359 -18925 18393 -18909
rect 8899 -19002 8915 -18968
rect 9135 -19002 9151 -18968
rect 9357 -19002 9373 -18968
rect 9593 -19002 9609 -18968
rect 9815 -19002 9831 -18968
rect 10051 -19002 10067 -18968
rect 10273 -19002 10289 -18968
rect 10509 -19002 10525 -18968
rect 10731 -19002 10747 -18968
rect 10967 -19002 10983 -18968
rect 11189 -19002 11205 -18968
rect 11425 -19002 11441 -18968
rect 11647 -19002 11663 -18968
rect 11883 -19002 11899 -18968
rect 12105 -19002 12121 -18968
rect 12341 -19002 12357 -18968
rect 12563 -19002 12579 -18968
rect 12799 -19002 12815 -18968
rect 13021 -19002 13037 -18968
rect 13257 -19002 13273 -18968
rect 13899 -19002 13915 -18968
rect 14135 -19002 14151 -18968
rect 14357 -19002 14373 -18968
rect 14593 -19002 14609 -18968
rect 14815 -19002 14831 -18968
rect 15051 -19002 15067 -18968
rect 15273 -19002 15289 -18968
rect 15509 -19002 15525 -18968
rect 15731 -19002 15747 -18968
rect 15967 -19002 15983 -18968
rect 16189 -19002 16205 -18968
rect 16425 -19002 16441 -18968
rect 16647 -19002 16663 -18968
rect 16883 -19002 16899 -18968
rect 17105 -19002 17121 -18968
rect 17341 -19002 17357 -18968
rect 17563 -19002 17579 -18968
rect 17799 -19002 17815 -18968
rect 18021 -19002 18037 -18968
rect 18257 -19002 18273 -18968
rect 8352 -19448 8452 -19286
rect 18696 -19448 18796 -19286
rect 23352 -13766 23452 -13604
rect 33696 -13766 33796 -13604
rect 24458 -15009 24474 -14975
rect 24694 -15009 24710 -14975
rect 24916 -15009 24932 -14975
rect 25152 -15009 25168 -14975
rect 25374 -15009 25390 -14975
rect 25610 -15009 25626 -14975
rect 25832 -15009 25848 -14975
rect 26068 -15009 26084 -14975
rect 26290 -15009 26306 -14975
rect 26526 -15009 26542 -14975
rect 26748 -15009 26764 -14975
rect 26984 -15009 27000 -14975
rect 27206 -15009 27222 -14975
rect 27442 -15009 27458 -14975
rect 27664 -15009 27680 -14975
rect 27900 -15009 27916 -14975
rect 28122 -15009 28138 -14975
rect 28358 -15009 28374 -14975
rect 28580 -15009 28596 -14975
rect 28816 -15009 28832 -14975
rect 29038 -15009 29054 -14975
rect 29274 -15009 29290 -14975
rect 29496 -15009 29512 -14975
rect 29732 -15009 29748 -14975
rect 29954 -15009 29970 -14975
rect 30190 -15009 30206 -14975
rect 30412 -15009 30428 -14975
rect 30648 -15009 30664 -14975
rect 30870 -15009 30886 -14975
rect 31106 -15009 31122 -14975
rect 31328 -15009 31344 -14975
rect 31564 -15009 31580 -14975
rect 31786 -15009 31802 -14975
rect 32022 -15009 32038 -14975
rect 32244 -15009 32260 -14975
rect 32480 -15009 32496 -14975
rect 24338 -15068 24372 -15052
rect 24338 -16660 24372 -16644
rect 24796 -15068 24830 -15052
rect 24796 -16660 24830 -16644
rect 25254 -15068 25288 -15052
rect 25254 -16660 25288 -16644
rect 25712 -15068 25746 -15052
rect 25712 -16660 25746 -16644
rect 26170 -15068 26204 -15052
rect 26170 -16660 26204 -16644
rect 26628 -15068 26662 -15052
rect 26628 -16660 26662 -16644
rect 27086 -15068 27120 -15052
rect 27086 -16660 27120 -16644
rect 27544 -15068 27578 -15052
rect 27544 -16660 27578 -16644
rect 28002 -15068 28036 -15052
rect 28002 -16660 28036 -16644
rect 28460 -15068 28494 -15052
rect 28460 -16660 28494 -16644
rect 28918 -15068 28952 -15052
rect 28918 -16660 28952 -16644
rect 29376 -15068 29410 -15052
rect 29376 -16660 29410 -16644
rect 29834 -15068 29868 -15052
rect 29834 -16660 29868 -16644
rect 30292 -15068 30326 -15052
rect 30292 -16660 30326 -16644
rect 30750 -15068 30784 -15052
rect 30750 -16660 30784 -16644
rect 31208 -15068 31242 -15052
rect 31208 -16660 31242 -16644
rect 31666 -15068 31700 -15052
rect 31666 -16660 31700 -16644
rect 32124 -15068 32158 -15052
rect 32124 -16660 32158 -16644
rect 32582 -15068 32616 -15052
rect 32582 -16660 32616 -16644
rect 24458 -16737 24474 -16703
rect 24694 -16737 24710 -16703
rect 24916 -16737 24932 -16703
rect 25152 -16737 25168 -16703
rect 25374 -16737 25390 -16703
rect 25610 -16737 25626 -16703
rect 25832 -16737 25848 -16703
rect 26068 -16737 26084 -16703
rect 26290 -16737 26306 -16703
rect 26526 -16737 26542 -16703
rect 26748 -16737 26764 -16703
rect 26984 -16737 27000 -16703
rect 27206 -16737 27222 -16703
rect 27442 -16737 27458 -16703
rect 27664 -16737 27680 -16703
rect 27900 -16737 27916 -16703
rect 28122 -16737 28138 -16703
rect 28358 -16737 28374 -16703
rect 28580 -16737 28596 -16703
rect 28816 -16737 28832 -16703
rect 29038 -16737 29054 -16703
rect 29274 -16737 29290 -16703
rect 29496 -16737 29512 -16703
rect 29732 -16737 29748 -16703
rect 29954 -16737 29970 -16703
rect 30190 -16737 30206 -16703
rect 30412 -16737 30428 -16703
rect 30648 -16737 30664 -16703
rect 30870 -16737 30886 -16703
rect 31106 -16737 31122 -16703
rect 31328 -16737 31344 -16703
rect 31564 -16737 31580 -16703
rect 31786 -16737 31802 -16703
rect 32022 -16737 32038 -16703
rect 32244 -16737 32260 -16703
rect 32480 -16737 32496 -16703
rect 28216 -16820 28676 -16814
rect 28216 -16868 28222 -16820
rect 28270 -16868 28676 -16820
rect 28216 -16874 28676 -16868
rect 23899 -17674 23915 -17640
rect 24135 -17674 24151 -17640
rect 24357 -17674 24373 -17640
rect 24593 -17674 24609 -17640
rect 24815 -17674 24831 -17640
rect 25051 -17674 25067 -17640
rect 25273 -17674 25289 -17640
rect 25509 -17674 25525 -17640
rect 25731 -17674 25747 -17640
rect 25967 -17674 25983 -17640
rect 26189 -17674 26205 -17640
rect 26425 -17674 26441 -17640
rect 26647 -17674 26663 -17640
rect 26883 -17674 26899 -17640
rect 27105 -17674 27121 -17640
rect 27341 -17674 27357 -17640
rect 27563 -17674 27579 -17640
rect 27799 -17674 27815 -17640
rect 28021 -17674 28037 -17640
rect 28257 -17674 28273 -17640
rect 28899 -17674 28915 -17640
rect 29135 -17674 29151 -17640
rect 29357 -17674 29373 -17640
rect 29593 -17674 29609 -17640
rect 29815 -17674 29831 -17640
rect 30051 -17674 30067 -17640
rect 30273 -17674 30289 -17640
rect 30509 -17674 30525 -17640
rect 30731 -17674 30747 -17640
rect 30967 -17674 30983 -17640
rect 31189 -17674 31205 -17640
rect 31425 -17674 31441 -17640
rect 31647 -17674 31663 -17640
rect 31883 -17674 31899 -17640
rect 32105 -17674 32121 -17640
rect 32341 -17674 32357 -17640
rect 32563 -17674 32579 -17640
rect 32799 -17674 32815 -17640
rect 33021 -17674 33037 -17640
rect 33257 -17674 33273 -17640
rect 23779 -17733 23813 -17717
rect 23779 -18925 23813 -18909
rect 24237 -17733 24271 -17717
rect 24237 -18925 24271 -18909
rect 24695 -17733 24729 -17717
rect 24695 -18925 24729 -18909
rect 25153 -17733 25187 -17717
rect 25153 -18925 25187 -18909
rect 25611 -17733 25645 -17717
rect 25611 -18925 25645 -18909
rect 26069 -17733 26103 -17717
rect 26069 -18925 26103 -18909
rect 26527 -17733 26561 -17717
rect 26527 -18925 26561 -18909
rect 26985 -17733 27019 -17717
rect 26985 -18925 27019 -18909
rect 27443 -17733 27477 -17717
rect 27443 -18925 27477 -18909
rect 27901 -17733 27935 -17717
rect 27901 -18925 27935 -18909
rect 28359 -17733 28393 -17717
rect 28359 -18925 28393 -18909
rect 28779 -17733 28813 -17717
rect 28779 -18925 28813 -18909
rect 29237 -17733 29271 -17717
rect 29237 -18925 29271 -18909
rect 29695 -17733 29729 -17717
rect 29695 -18925 29729 -18909
rect 30153 -17733 30187 -17717
rect 30153 -18925 30187 -18909
rect 30611 -17733 30645 -17717
rect 30611 -18925 30645 -18909
rect 31069 -17733 31103 -17717
rect 31069 -18925 31103 -18909
rect 31527 -17733 31561 -17717
rect 31527 -18925 31561 -18909
rect 31985 -17733 32019 -17717
rect 31985 -18925 32019 -18909
rect 32443 -17733 32477 -17717
rect 32443 -18925 32477 -18909
rect 32901 -17733 32935 -17717
rect 32901 -18925 32935 -18909
rect 33359 -17733 33393 -17717
rect 33359 -18925 33393 -18909
rect 23899 -19002 23915 -18968
rect 24135 -19002 24151 -18968
rect 24357 -19002 24373 -18968
rect 24593 -19002 24609 -18968
rect 24815 -19002 24831 -18968
rect 25051 -19002 25067 -18968
rect 25273 -19002 25289 -18968
rect 25509 -19002 25525 -18968
rect 25731 -19002 25747 -18968
rect 25967 -19002 25983 -18968
rect 26189 -19002 26205 -18968
rect 26425 -19002 26441 -18968
rect 26647 -19002 26663 -18968
rect 26883 -19002 26899 -18968
rect 27105 -19002 27121 -18968
rect 27341 -19002 27357 -18968
rect 27563 -19002 27579 -18968
rect 27799 -19002 27815 -18968
rect 28021 -19002 28037 -18968
rect 28257 -19002 28273 -18968
rect 28899 -19002 28915 -18968
rect 29135 -19002 29151 -18968
rect 29357 -19002 29373 -18968
rect 29593 -19002 29609 -18968
rect 29815 -19002 29831 -18968
rect 30051 -19002 30067 -18968
rect 30273 -19002 30289 -18968
rect 30509 -19002 30525 -18968
rect 30731 -19002 30747 -18968
rect 30967 -19002 30983 -18968
rect 31189 -19002 31205 -18968
rect 31425 -19002 31441 -18968
rect 31647 -19002 31663 -18968
rect 31883 -19002 31899 -18968
rect 32105 -19002 32121 -18968
rect 32341 -19002 32357 -18968
rect 32563 -19002 32579 -18968
rect 32799 -19002 32815 -18968
rect 33021 -19002 33037 -18968
rect 33257 -19002 33273 -18968
rect 23352 -19448 23452 -19286
rect 33696 -19448 33796 -19286
rect 8352 -19846 8452 -19684
rect 18696 -19846 18796 -19684
rect 8898 -20176 8914 -20142
rect 9134 -20176 9150 -20142
rect 9356 -20176 9372 -20142
rect 9592 -20176 9608 -20142
rect 9814 -20176 9830 -20142
rect 10050 -20176 10066 -20142
rect 10272 -20176 10288 -20142
rect 10508 -20176 10524 -20142
rect 10730 -20176 10746 -20142
rect 10966 -20176 10982 -20142
rect 11188 -20176 11204 -20142
rect 11424 -20176 11440 -20142
rect 11646 -20176 11662 -20142
rect 11882 -20176 11898 -20142
rect 12104 -20176 12120 -20142
rect 12340 -20176 12356 -20142
rect 12562 -20176 12578 -20142
rect 12798 -20176 12814 -20142
rect 13020 -20176 13036 -20142
rect 13256 -20176 13272 -20142
rect 13898 -20176 13914 -20142
rect 14134 -20176 14150 -20142
rect 14356 -20176 14372 -20142
rect 14592 -20176 14608 -20142
rect 14814 -20176 14830 -20142
rect 15050 -20176 15066 -20142
rect 15272 -20176 15288 -20142
rect 15508 -20176 15524 -20142
rect 15730 -20176 15746 -20142
rect 15966 -20176 15982 -20142
rect 16188 -20176 16204 -20142
rect 16424 -20176 16440 -20142
rect 16646 -20176 16662 -20142
rect 16882 -20176 16898 -20142
rect 17104 -20176 17120 -20142
rect 17340 -20176 17356 -20142
rect 17562 -20176 17578 -20142
rect 17798 -20176 17814 -20142
rect 18020 -20176 18036 -20142
rect 18256 -20176 18272 -20142
rect 8778 -20226 8812 -20210
rect 8778 -20418 8812 -20402
rect 9236 -20226 9270 -20210
rect 9236 -20418 9270 -20402
rect 9694 -20226 9728 -20210
rect 9694 -20418 9728 -20402
rect 10152 -20226 10186 -20210
rect 10152 -20418 10186 -20402
rect 10610 -20226 10644 -20210
rect 10610 -20418 10644 -20402
rect 11068 -20226 11102 -20210
rect 11068 -20418 11102 -20402
rect 11526 -20226 11560 -20210
rect 11526 -20418 11560 -20402
rect 11984 -20226 12018 -20210
rect 11984 -20418 12018 -20402
rect 12442 -20226 12476 -20210
rect 12442 -20418 12476 -20402
rect 12900 -20226 12934 -20210
rect 12900 -20418 12934 -20402
rect 13358 -20226 13392 -20210
rect 13358 -20418 13392 -20402
rect 13778 -20226 13812 -20210
rect 13778 -20418 13812 -20402
rect 14236 -20226 14270 -20210
rect 14236 -20418 14270 -20402
rect 14694 -20226 14728 -20210
rect 14694 -20418 14728 -20402
rect 15152 -20226 15186 -20210
rect 15152 -20418 15186 -20402
rect 15610 -20226 15644 -20210
rect 15610 -20418 15644 -20402
rect 16068 -20226 16102 -20210
rect 16068 -20418 16102 -20402
rect 16526 -20226 16560 -20210
rect 16526 -20418 16560 -20402
rect 16984 -20226 17018 -20210
rect 16984 -20418 17018 -20402
rect 17442 -20226 17476 -20210
rect 17442 -20418 17476 -20402
rect 17900 -20226 17934 -20210
rect 17900 -20418 17934 -20402
rect 18358 -20226 18392 -20210
rect 18358 -20418 18392 -20402
rect 8898 -20486 8914 -20452
rect 9134 -20486 9150 -20452
rect 9356 -20486 9372 -20452
rect 9592 -20486 9608 -20452
rect 9814 -20486 9830 -20452
rect 10050 -20486 10066 -20452
rect 10272 -20486 10288 -20452
rect 10508 -20486 10524 -20452
rect 10730 -20486 10746 -20452
rect 10966 -20486 10982 -20452
rect 11188 -20486 11204 -20452
rect 11424 -20486 11440 -20452
rect 11646 -20486 11662 -20452
rect 11882 -20486 11898 -20452
rect 12104 -20486 12120 -20452
rect 12340 -20486 12356 -20452
rect 12562 -20486 12578 -20452
rect 12798 -20486 12814 -20452
rect 13020 -20486 13036 -20452
rect 13256 -20486 13272 -20452
rect 13898 -20486 13914 -20452
rect 14134 -20486 14150 -20452
rect 14356 -20486 14372 -20452
rect 14592 -20486 14608 -20452
rect 14814 -20486 14830 -20452
rect 15050 -20486 15066 -20452
rect 15272 -20486 15288 -20452
rect 15508 -20486 15524 -20452
rect 15730 -20486 15746 -20452
rect 15966 -20486 15982 -20452
rect 16188 -20486 16204 -20452
rect 16424 -20486 16440 -20452
rect 16646 -20486 16662 -20452
rect 16882 -20486 16898 -20452
rect 17104 -20486 17120 -20452
rect 17340 -20486 17356 -20452
rect 17562 -20486 17578 -20452
rect 17798 -20486 17814 -20452
rect 18020 -20486 18036 -20452
rect 18256 -20486 18272 -20452
rect 8898 -20844 8914 -20810
rect 9134 -20844 9150 -20810
rect 9356 -20844 9372 -20810
rect 9592 -20844 9608 -20810
rect 9814 -20844 9830 -20810
rect 10050 -20844 10066 -20810
rect 10272 -20844 10288 -20810
rect 10508 -20844 10524 -20810
rect 10730 -20844 10746 -20810
rect 10966 -20844 10982 -20810
rect 11188 -20844 11204 -20810
rect 11424 -20844 11440 -20810
rect 11646 -20844 11662 -20810
rect 11882 -20844 11898 -20810
rect 12104 -20844 12120 -20810
rect 12340 -20844 12356 -20810
rect 12562 -20844 12578 -20810
rect 12798 -20844 12814 -20810
rect 13020 -20844 13036 -20810
rect 13256 -20844 13272 -20810
rect 8778 -20894 8812 -20878
rect 8778 -21086 8812 -21070
rect 9236 -20894 9270 -20878
rect 9236 -21086 9270 -21070
rect 9694 -20894 9728 -20878
rect 9694 -21086 9728 -21070
rect 10152 -20894 10186 -20878
rect 10152 -21086 10186 -21070
rect 10610 -20894 10644 -20878
rect 10610 -21086 10644 -21070
rect 11068 -20894 11102 -20878
rect 11068 -21086 11102 -21070
rect 11526 -20894 11560 -20878
rect 11526 -21086 11560 -21070
rect 11984 -20894 12018 -20878
rect 11984 -21086 12018 -21070
rect 12442 -20894 12476 -20878
rect 12442 -21086 12476 -21070
rect 12900 -20894 12934 -20878
rect 12900 -21086 12934 -21070
rect 13358 -20894 13392 -20878
rect 13358 -21086 13392 -21070
rect 8898 -21154 8914 -21120
rect 9134 -21154 9150 -21120
rect 9356 -21154 9372 -21120
rect 9592 -21154 9608 -21120
rect 9814 -21154 9830 -21120
rect 10050 -21154 10066 -21120
rect 10272 -21154 10288 -21120
rect 10508 -21154 10524 -21120
rect 10730 -21154 10746 -21120
rect 10966 -21154 10982 -21120
rect 11188 -21154 11204 -21120
rect 11424 -21154 11440 -21120
rect 11646 -21154 11662 -21120
rect 11882 -21154 11898 -21120
rect 12104 -21154 12120 -21120
rect 12340 -21154 12356 -21120
rect 12562 -21154 12578 -21120
rect 12798 -21154 12814 -21120
rect 13020 -21154 13036 -21120
rect 13256 -21154 13272 -21120
rect 8352 -22148 8452 -21986
rect 18696 -22148 18796 -21986
rect 23352 -19846 23452 -19684
rect 33696 -19846 33796 -19684
rect 23898 -20176 23914 -20142
rect 24134 -20176 24150 -20142
rect 24356 -20176 24372 -20142
rect 24592 -20176 24608 -20142
rect 24814 -20176 24830 -20142
rect 25050 -20176 25066 -20142
rect 25272 -20176 25288 -20142
rect 25508 -20176 25524 -20142
rect 25730 -20176 25746 -20142
rect 25966 -20176 25982 -20142
rect 26188 -20176 26204 -20142
rect 26424 -20176 26440 -20142
rect 26646 -20176 26662 -20142
rect 26882 -20176 26898 -20142
rect 27104 -20176 27120 -20142
rect 27340 -20176 27356 -20142
rect 27562 -20176 27578 -20142
rect 27798 -20176 27814 -20142
rect 28020 -20176 28036 -20142
rect 28256 -20176 28272 -20142
rect 28898 -20176 28914 -20142
rect 29134 -20176 29150 -20142
rect 29356 -20176 29372 -20142
rect 29592 -20176 29608 -20142
rect 29814 -20176 29830 -20142
rect 30050 -20176 30066 -20142
rect 30272 -20176 30288 -20142
rect 30508 -20176 30524 -20142
rect 30730 -20176 30746 -20142
rect 30966 -20176 30982 -20142
rect 31188 -20176 31204 -20142
rect 31424 -20176 31440 -20142
rect 31646 -20176 31662 -20142
rect 31882 -20176 31898 -20142
rect 32104 -20176 32120 -20142
rect 32340 -20176 32356 -20142
rect 32562 -20176 32578 -20142
rect 32798 -20176 32814 -20142
rect 33020 -20176 33036 -20142
rect 33256 -20176 33272 -20142
rect 23778 -20226 23812 -20210
rect 23778 -20418 23812 -20402
rect 24236 -20226 24270 -20210
rect 24236 -20418 24270 -20402
rect 24694 -20226 24728 -20210
rect 24694 -20418 24728 -20402
rect 25152 -20226 25186 -20210
rect 25152 -20418 25186 -20402
rect 25610 -20226 25644 -20210
rect 25610 -20418 25644 -20402
rect 26068 -20226 26102 -20210
rect 26068 -20418 26102 -20402
rect 26526 -20226 26560 -20210
rect 26526 -20418 26560 -20402
rect 26984 -20226 27018 -20210
rect 26984 -20418 27018 -20402
rect 27442 -20226 27476 -20210
rect 27442 -20418 27476 -20402
rect 27900 -20226 27934 -20210
rect 27900 -20418 27934 -20402
rect 28358 -20226 28392 -20210
rect 28358 -20418 28392 -20402
rect 28778 -20226 28812 -20210
rect 28778 -20418 28812 -20402
rect 29236 -20226 29270 -20210
rect 29236 -20418 29270 -20402
rect 29694 -20226 29728 -20210
rect 29694 -20418 29728 -20402
rect 30152 -20226 30186 -20210
rect 30152 -20418 30186 -20402
rect 30610 -20226 30644 -20210
rect 30610 -20418 30644 -20402
rect 31068 -20226 31102 -20210
rect 31068 -20418 31102 -20402
rect 31526 -20226 31560 -20210
rect 31526 -20418 31560 -20402
rect 31984 -20226 32018 -20210
rect 31984 -20418 32018 -20402
rect 32442 -20226 32476 -20210
rect 32442 -20418 32476 -20402
rect 32900 -20226 32934 -20210
rect 32900 -20418 32934 -20402
rect 33358 -20226 33392 -20210
rect 33358 -20418 33392 -20402
rect 23898 -20486 23914 -20452
rect 24134 -20486 24150 -20452
rect 24356 -20486 24372 -20452
rect 24592 -20486 24608 -20452
rect 24814 -20486 24830 -20452
rect 25050 -20486 25066 -20452
rect 25272 -20486 25288 -20452
rect 25508 -20486 25524 -20452
rect 25730 -20486 25746 -20452
rect 25966 -20486 25982 -20452
rect 26188 -20486 26204 -20452
rect 26424 -20486 26440 -20452
rect 26646 -20486 26662 -20452
rect 26882 -20486 26898 -20452
rect 27104 -20486 27120 -20452
rect 27340 -20486 27356 -20452
rect 27562 -20486 27578 -20452
rect 27798 -20486 27814 -20452
rect 28020 -20486 28036 -20452
rect 28256 -20486 28272 -20452
rect 28898 -20486 28914 -20452
rect 29134 -20486 29150 -20452
rect 29356 -20486 29372 -20452
rect 29592 -20486 29608 -20452
rect 29814 -20486 29830 -20452
rect 30050 -20486 30066 -20452
rect 30272 -20486 30288 -20452
rect 30508 -20486 30524 -20452
rect 30730 -20486 30746 -20452
rect 30966 -20486 30982 -20452
rect 31188 -20486 31204 -20452
rect 31424 -20486 31440 -20452
rect 31646 -20486 31662 -20452
rect 31882 -20486 31898 -20452
rect 32104 -20486 32120 -20452
rect 32340 -20486 32356 -20452
rect 32562 -20486 32578 -20452
rect 32798 -20486 32814 -20452
rect 33020 -20486 33036 -20452
rect 33256 -20486 33272 -20452
rect 23898 -20844 23914 -20810
rect 24134 -20844 24150 -20810
rect 24356 -20844 24372 -20810
rect 24592 -20844 24608 -20810
rect 24814 -20844 24830 -20810
rect 25050 -20844 25066 -20810
rect 25272 -20844 25288 -20810
rect 25508 -20844 25524 -20810
rect 25730 -20844 25746 -20810
rect 25966 -20844 25982 -20810
rect 26188 -20844 26204 -20810
rect 26424 -20844 26440 -20810
rect 26646 -20844 26662 -20810
rect 26882 -20844 26898 -20810
rect 27104 -20844 27120 -20810
rect 27340 -20844 27356 -20810
rect 27562 -20844 27578 -20810
rect 27798 -20844 27814 -20810
rect 28020 -20844 28036 -20810
rect 28256 -20844 28272 -20810
rect 23778 -20894 23812 -20878
rect 23778 -21086 23812 -21070
rect 24236 -20894 24270 -20878
rect 24236 -21086 24270 -21070
rect 24694 -20894 24728 -20878
rect 24694 -21086 24728 -21070
rect 25152 -20894 25186 -20878
rect 25152 -21086 25186 -21070
rect 25610 -20894 25644 -20878
rect 25610 -21086 25644 -21070
rect 26068 -20894 26102 -20878
rect 26068 -21086 26102 -21070
rect 26526 -20894 26560 -20878
rect 26526 -21086 26560 -21070
rect 26984 -20894 27018 -20878
rect 26984 -21086 27018 -21070
rect 27442 -20894 27476 -20878
rect 27442 -21086 27476 -21070
rect 27900 -20894 27934 -20878
rect 27900 -21086 27934 -21070
rect 28358 -20894 28392 -20878
rect 28358 -21086 28392 -21070
rect 23898 -21154 23914 -21120
rect 24134 -21154 24150 -21120
rect 24356 -21154 24372 -21120
rect 24592 -21154 24608 -21120
rect 24814 -21154 24830 -21120
rect 25050 -21154 25066 -21120
rect 25272 -21154 25288 -21120
rect 25508 -21154 25524 -21120
rect 25730 -21154 25746 -21120
rect 25966 -21154 25982 -21120
rect 26188 -21154 26204 -21120
rect 26424 -21154 26440 -21120
rect 26646 -21154 26662 -21120
rect 26882 -21154 26898 -21120
rect 27104 -21154 27120 -21120
rect 27340 -21154 27356 -21120
rect 27562 -21154 27578 -21120
rect 27798 -21154 27814 -21120
rect 28020 -21154 28036 -21120
rect 28256 -21154 28272 -21120
rect 23352 -22148 23452 -21986
rect 33696 -22148 33796 -21986
<< viali >>
rect 23434 17400 23496 17500
rect 23496 17400 32616 17500
rect 32616 17400 32678 17500
rect 23334 15401 23434 17295
rect 24030 16481 24414 16515
rect 24888 16481 25272 16515
rect 25746 16481 26130 16515
rect 26604 16481 26988 16515
rect 27462 16481 27846 16515
rect 28320 16481 28704 16515
rect 29178 16481 29562 16515
rect 30036 16481 30420 16515
rect 30894 16481 31278 16515
rect 31752 16481 32136 16515
rect 23776 16246 23810 16422
rect 24634 16246 24668 16422
rect 25492 16246 25526 16422
rect 26350 16246 26384 16422
rect 27208 16246 27242 16422
rect 28066 16246 28100 16422
rect 28924 16246 28958 16422
rect 29782 16246 29816 16422
rect 30640 16246 30674 16422
rect 31498 16246 31532 16422
rect 32356 16246 32390 16422
rect 24030 16153 24414 16187
rect 24888 16153 25272 16187
rect 25746 16153 26130 16187
rect 26604 16153 26988 16187
rect 27462 16153 27846 16187
rect 28320 16153 28704 16187
rect 29178 16153 29562 16187
rect 30036 16153 30420 16187
rect 30894 16153 31278 16187
rect 31752 16153 32136 16187
rect 24030 15881 24414 15915
rect 24888 15881 25272 15915
rect 25746 15881 26130 15915
rect 26604 15881 26988 15915
rect 27462 15881 27846 15915
rect 28320 15881 28704 15915
rect 29178 15881 29562 15915
rect 30036 15881 30420 15915
rect 30894 15881 31278 15915
rect 31752 15881 32136 15915
rect 23776 15646 23810 15822
rect 24634 15646 24668 15822
rect 25492 15646 25526 15822
rect 26350 15646 26384 15822
rect 27208 15646 27242 15822
rect 28066 15646 28100 15822
rect 28924 15646 28958 15822
rect 29782 15646 29816 15822
rect 30640 15646 30674 15822
rect 31498 15646 31532 15822
rect 32356 15646 32390 15822
rect 24030 15553 24414 15587
rect 24888 15553 25272 15587
rect 25746 15553 26130 15587
rect 26604 15553 26988 15587
rect 27462 15553 27846 15587
rect 28320 15553 28704 15587
rect 29178 15553 29562 15587
rect 30036 15553 30420 15587
rect 30894 15553 31278 15587
rect 31752 15553 32136 15587
rect 32678 15401 32778 17295
rect 23434 15196 23496 15296
rect 23496 15196 32616 15296
rect 32616 15196 32678 15296
rect 24048 14881 24084 14882
rect 24048 14308 24049 14881
rect 24049 14308 24083 14881
rect 24083 14308 24084 14881
rect 25050 14881 25086 14882
rect 24267 14841 24351 14875
rect 24525 14841 24609 14875
rect 24783 14841 24867 14875
rect 24163 14406 24197 14782
rect 24421 14406 24455 14782
rect 24679 14406 24713 14782
rect 24937 14406 24971 14782
rect 24267 14313 24351 14347
rect 24525 14313 24609 14347
rect 24783 14313 24867 14347
rect 25050 14308 25051 14881
rect 25051 14308 25085 14881
rect 25085 14308 25086 14881
rect 25170 14881 25206 14882
rect 25170 14308 25171 14881
rect 25171 14308 25205 14881
rect 25205 14308 25206 14881
rect 26948 14881 26982 14884
rect 25389 14841 25473 14875
rect 25647 14841 25731 14875
rect 25905 14841 25989 14875
rect 26163 14841 26247 14875
rect 26421 14841 26505 14875
rect 26679 14841 26763 14875
rect 25285 14406 25319 14782
rect 25543 14406 25577 14782
rect 25801 14406 25835 14782
rect 26059 14406 26093 14782
rect 26317 14406 26351 14782
rect 26575 14406 26609 14782
rect 26833 14406 26867 14782
rect 25389 14313 25473 14347
rect 25647 14313 25731 14347
rect 25905 14313 25989 14347
rect 26163 14313 26247 14347
rect 26421 14313 26505 14347
rect 26679 14313 26763 14347
rect 26948 14308 26981 14881
rect 26981 14308 26982 14881
rect 27289 14441 27323 14475
rect 27381 14441 27415 14475
rect 27473 14441 27507 14475
rect 27565 14441 27599 14475
rect 27657 14441 27691 14475
rect 27749 14441 27783 14475
rect 27841 14441 27875 14475
rect 27933 14441 27967 14475
rect 28025 14441 28059 14475
rect 28117 14441 28151 14475
rect 28209 14441 28243 14475
rect 28301 14441 28335 14475
rect 28393 14441 28427 14475
rect 28485 14441 28519 14475
rect 28577 14441 28611 14475
rect 28669 14441 28703 14475
rect 28761 14441 28795 14475
rect 28853 14441 28887 14475
rect 28945 14441 28979 14475
rect 29037 14441 29071 14475
rect 29129 14441 29163 14475
rect 29221 14441 29255 14475
rect 29313 14441 29347 14475
rect 29405 14441 29439 14475
rect 29497 14441 29531 14475
rect 29589 14441 29623 14475
rect 29681 14441 29715 14475
rect 29773 14441 29807 14475
rect 29865 14441 29899 14475
rect 29957 14441 29991 14475
rect 30049 14441 30083 14475
rect 30141 14441 30175 14475
rect 30233 14441 30267 14475
rect 30325 14441 30359 14475
rect 30417 14441 30451 14475
rect 30509 14441 30543 14475
rect 30601 14441 30635 14475
rect 30693 14441 30727 14475
rect 30785 14441 30819 14475
rect 30877 14441 30911 14475
rect 30969 14441 31003 14475
rect 31061 14441 31095 14475
rect 31153 14441 31187 14475
rect 31245 14441 31279 14475
rect 31337 14441 31371 14475
rect 31429 14441 31463 14475
rect 31521 14441 31555 14475
rect 31613 14441 31647 14475
rect 31705 14441 31739 14475
rect 31797 14441 31831 14475
rect 31889 14441 31923 14475
rect 31981 14441 32015 14475
rect 32073 14441 32107 14475
rect 32165 14441 32199 14475
rect 32257 14441 32291 14475
rect 27274 14163 27322 14190
rect 27274 14142 27292 14163
rect 27292 14142 27322 14163
rect 27382 14144 27394 14169
rect 27394 14144 27416 14169
rect 27382 14135 27416 14144
rect 24048 13985 24082 13986
rect 24048 13630 24049 13985
rect 24049 13630 24082 13985
rect 24267 13945 24351 13979
rect 24525 13945 24609 13979
rect 24783 13945 24867 13979
rect 24163 13719 24197 13895
rect 24421 13719 24455 13895
rect 24679 13719 24713 13895
rect 24937 13719 24971 13895
rect 24267 13635 24351 13669
rect 24525 13635 24609 13669
rect 24783 13635 24867 13669
rect 25050 13630 25051 13984
rect 25051 13630 25084 13984
rect 25170 13630 25171 13984
rect 25171 13630 25204 13984
rect 26946 13985 26980 13986
rect 25389 13945 25473 13979
rect 25647 13945 25731 13979
rect 25905 13945 25989 13979
rect 26163 13945 26247 13979
rect 26421 13945 26505 13979
rect 26679 13945 26763 13979
rect 25285 13719 25319 13895
rect 25543 13719 25577 13895
rect 25801 13719 25835 13895
rect 26059 13719 26093 13895
rect 26317 13719 26351 13895
rect 26575 13719 26609 13895
rect 26833 13719 26867 13895
rect 25389 13635 25473 13669
rect 25647 13635 25731 13669
rect 25905 13635 25989 13669
rect 26163 13635 26247 13669
rect 26421 13635 26505 13669
rect 26679 13635 26763 13669
rect 26946 13630 26947 13985
rect 26947 13630 26980 13985
rect 27463 14289 27497 14305
rect 27463 14271 27497 14289
rect 27542 14348 27582 14388
rect 27841 14271 27875 14305
rect 27749 14135 27783 14169
rect 28465 14279 28499 14305
rect 28465 14271 28496 14279
rect 28496 14271 28499 14279
rect 28021 14067 28055 14101
rect 28093 14083 28117 14101
rect 28117 14083 28127 14101
rect 28093 14067 28127 14083
rect 28465 14153 28499 14169
rect 28465 14135 28491 14153
rect 28491 14135 28499 14153
rect 28681 14155 28715 14164
rect 28681 14130 28697 14155
rect 28697 14130 28715 14155
rect 28741 14067 28775 14101
rect 29004 14122 29052 14170
rect 29764 14263 29812 14268
rect 29764 14229 29775 14263
rect 29775 14229 29809 14263
rect 29809 14229 29812 14263
rect 29764 14226 29812 14229
rect 30000 14365 30010 14368
rect 30010 14365 30044 14368
rect 30044 14365 30048 14368
rect 30000 14331 30048 14365
rect 30000 14320 30010 14331
rect 30010 14320 30044 14331
rect 30044 14320 30048 14331
rect 29444 14163 29492 14170
rect 29444 14130 29456 14163
rect 29456 14130 29490 14163
rect 29490 14130 29492 14163
rect 29682 14163 29730 14170
rect 29682 14129 29688 14163
rect 29688 14129 29722 14163
rect 29722 14129 29730 14163
rect 29682 14128 29730 14129
rect 29856 14163 29904 14170
rect 29856 14129 29890 14163
rect 29890 14129 29904 14163
rect 29856 14128 29904 14129
rect 30090 14163 30138 14170
rect 30090 14130 30124 14163
rect 30124 14130 30138 14163
rect 29532 14045 29536 14058
rect 29536 14045 29570 14058
rect 29570 14045 29580 14058
rect 29532 14011 29580 14045
rect 29532 14010 29536 14011
rect 29536 14010 29570 14011
rect 29570 14010 29580 14011
rect 31081 14279 31115 14305
rect 31081 14271 31084 14279
rect 31084 14271 31115 14279
rect 31992 14356 32038 14396
rect 30528 14122 30576 14170
rect 30865 14155 30899 14164
rect 30865 14130 30883 14155
rect 30883 14130 30899 14155
rect 30805 14067 30839 14101
rect 31081 14153 31115 14169
rect 31081 14135 31089 14153
rect 31089 14135 31115 14153
rect 31705 14271 31739 14305
rect 31453 14083 31463 14101
rect 31463 14083 31487 14101
rect 31453 14067 31487 14083
rect 31525 14067 31559 14101
rect 31797 14135 31831 14169
rect 32083 14289 32117 14305
rect 32083 14271 32117 14289
rect 32164 14144 32186 14169
rect 32186 14144 32198 14169
rect 32164 14135 32198 14144
rect 32252 14163 32300 14172
rect 32252 14129 32254 14163
rect 32254 14129 32288 14163
rect 32288 14129 32300 14163
rect 32252 14124 32300 14129
rect 27289 13897 27323 13931
rect 27381 13897 27415 13931
rect 27473 13897 27507 13931
rect 27565 13897 27599 13931
rect 27657 13897 27691 13931
rect 27749 13897 27783 13931
rect 27841 13897 27875 13931
rect 27933 13897 27967 13931
rect 28025 13897 28059 13931
rect 28117 13897 28151 13931
rect 28209 13897 28243 13931
rect 28301 13897 28335 13931
rect 28393 13897 28427 13931
rect 28485 13897 28519 13931
rect 28577 13897 28611 13931
rect 28669 13897 28703 13931
rect 28761 13897 28795 13931
rect 28853 13897 28887 13931
rect 28945 13897 28979 13931
rect 29037 13897 29071 13931
rect 29129 13897 29163 13931
rect 29221 13897 29255 13931
rect 29313 13897 29347 13931
rect 29405 13897 29439 13931
rect 29497 13897 29531 13931
rect 29589 13897 29623 13931
rect 29681 13897 29715 13931
rect 29773 13897 29807 13931
rect 29865 13897 29899 13931
rect 29957 13897 29991 13931
rect 30049 13897 30083 13931
rect 30141 13897 30175 13931
rect 30233 13897 30267 13931
rect 30325 13897 30359 13931
rect 30417 13897 30451 13931
rect 30509 13897 30543 13931
rect 30601 13897 30635 13931
rect 30693 13897 30727 13931
rect 30785 13897 30819 13931
rect 30877 13897 30911 13931
rect 30969 13897 31003 13931
rect 31061 13897 31095 13931
rect 31153 13897 31187 13931
rect 31245 13897 31279 13931
rect 31337 13897 31371 13931
rect 31429 13897 31463 13931
rect 31521 13897 31555 13931
rect 31613 13897 31647 13931
rect 31705 13897 31739 13931
rect 31797 13897 31831 13931
rect 31889 13897 31923 13931
rect 31981 13897 32015 13931
rect 32073 13897 32107 13931
rect 32165 13897 32199 13931
rect 32257 13897 32291 13931
rect 23434 13220 23496 13320
rect 23496 13220 32616 13320
rect 32616 13220 32678 13320
rect 23334 11254 23434 13122
rect 24504 12892 24888 12926
rect 25362 12892 25746 12926
rect 26220 12892 26604 12926
rect 27078 12892 27462 12926
rect 27936 12892 28320 12926
rect 28794 12892 29178 12926
rect 29652 12892 30036 12926
rect 30510 12892 30894 12926
rect 31368 12892 31752 12926
rect 24250 12666 24284 12842
rect 25108 12666 25142 12842
rect 25966 12666 26000 12842
rect 26824 12666 26858 12842
rect 27682 12666 27716 12842
rect 28540 12666 28574 12842
rect 29398 12666 29432 12842
rect 30256 12666 30290 12842
rect 31114 12666 31148 12842
rect 31972 12666 32006 12842
rect 24504 12582 24888 12616
rect 25362 12582 25746 12616
rect 26220 12582 26604 12616
rect 27078 12582 27462 12616
rect 27936 12582 28320 12616
rect 28794 12582 29178 12616
rect 29652 12582 30036 12616
rect 30510 12582 30894 12616
rect 31368 12582 31752 12616
rect 24504 12310 24888 12344
rect 25362 12310 25746 12344
rect 26220 12310 26604 12344
rect 27078 12310 27462 12344
rect 27936 12310 28320 12344
rect 28794 12310 29178 12344
rect 29652 12310 30036 12344
rect 30510 12310 30894 12344
rect 31368 12310 31752 12344
rect 24250 12084 24284 12260
rect 25108 12084 25142 12260
rect 25966 12084 26000 12260
rect 26824 12084 26858 12260
rect 27682 12084 27716 12260
rect 28540 12084 28574 12260
rect 29398 12084 29432 12260
rect 30256 12084 30290 12260
rect 31114 12084 31148 12260
rect 31972 12084 32006 12260
rect 24504 12000 24888 12034
rect 25362 12000 25746 12034
rect 26220 12000 26604 12034
rect 27078 12000 27462 12034
rect 27936 12000 28320 12034
rect 28794 12000 29178 12034
rect 29652 12000 30036 12034
rect 30510 12000 30894 12034
rect 31368 12000 31752 12034
rect 32678 11254 32778 13122
rect 23434 11056 23496 11156
rect 23496 11056 32616 11156
rect 32616 11056 32678 11156
rect 13060 10634 13122 10734
rect 13122 10634 21822 10734
rect 21822 10634 21884 10734
rect 12960 9122 13060 10546
rect 15322 9706 15506 9740
rect 15780 9706 15964 9740
rect 16238 9706 16422 9740
rect 16696 9706 16880 9740
rect 17154 9706 17338 9740
rect 17612 9706 17796 9740
rect 18070 9706 18254 9740
rect 18528 9706 18712 9740
rect 18986 9706 19170 9740
rect 19444 9706 19628 9740
rect 15168 9480 15202 9656
rect 15626 9480 15660 9656
rect 16084 9480 16118 9656
rect 16542 9480 16576 9656
rect 17000 9480 17034 9656
rect 17458 9480 17492 9656
rect 17916 9480 17950 9656
rect 18374 9480 18408 9656
rect 18832 9480 18866 9656
rect 19290 9480 19324 9656
rect 19748 9480 19782 9656
rect 15322 9396 15506 9430
rect 15780 9396 15964 9430
rect 16238 9396 16422 9430
rect 16696 9396 16880 9430
rect 17154 9396 17338 9430
rect 17612 9396 17796 9430
rect 18070 9396 18254 9430
rect 18528 9396 18712 9430
rect 18986 9396 19170 9430
rect 19444 9396 19628 9430
rect 21884 9122 21984 10546
rect 13060 8934 13122 9034
rect 13122 8934 21822 9034
rect 21822 8934 21884 9034
rect 23642 10634 23704 10734
rect 23704 10634 28824 10734
rect 28824 10634 28886 10734
rect 23542 9038 23642 10550
rect 24084 9706 24268 9740
rect 24542 9706 24726 9740
rect 25000 9706 25184 9740
rect 25458 9706 25642 9740
rect 25916 9706 26100 9740
rect 26374 9706 26558 9740
rect 26832 9706 27016 9740
rect 27290 9706 27474 9740
rect 27748 9706 27932 9740
rect 28206 9706 28390 9740
rect 23930 9480 23964 9656
rect 24388 9480 24422 9656
rect 24846 9480 24880 9656
rect 25304 9480 25338 9656
rect 25762 9480 25796 9656
rect 26220 9480 26254 9656
rect 26678 9480 26712 9656
rect 27136 9480 27170 9656
rect 27594 9480 27628 9656
rect 28052 9480 28086 9656
rect 28510 9480 28544 9656
rect 24084 9396 24268 9430
rect 24542 9396 24726 9430
rect 25000 9396 25184 9430
rect 25458 9396 25642 9430
rect 25916 9396 26100 9430
rect 26374 9396 26558 9430
rect 26832 9396 27016 9430
rect 27290 9396 27474 9430
rect 27748 9396 27932 9430
rect 28206 9396 28390 9430
rect 28886 9038 28986 10550
rect 23642 8854 23704 8954
rect 23704 8854 28824 8954
rect 28824 8854 28886 8954
rect 30239 8943 30273 8977
rect 30581 8943 30615 8977
rect 30673 8943 30707 8977
rect 30765 8943 30799 8977
rect 30857 8943 30891 8977
rect 30949 8943 30983 8977
rect 31041 8943 31075 8977
rect 31133 8943 31167 8977
rect 31225 8943 31259 8977
rect 31317 8943 31351 8977
rect 31409 8943 31443 8977
rect 31501 8943 31535 8977
rect 31593 8943 31627 8977
rect 31685 8943 31719 8977
rect 31777 8943 31811 8977
rect 31869 8943 31903 8977
rect 31961 8943 31995 8977
rect 32053 8943 32087 8977
rect 32145 8943 32179 8977
rect 32237 8943 32271 8977
rect 32329 8943 32363 8977
rect 32421 8943 32455 8977
rect 32513 8943 32547 8977
rect 32605 8943 32639 8977
rect 32697 8943 32731 8977
rect 32789 8943 32823 8977
rect 32881 8943 32915 8977
rect 32973 8943 33007 8977
rect 33139 8943 33173 8977
rect 36013 8943 36047 8977
rect 29105 8897 29139 8931
rect 29197 8897 29231 8931
rect 29289 8897 29323 8931
rect 29381 8897 29415 8931
rect 29473 8897 29507 8931
rect 29565 8897 29599 8931
rect 29657 8897 29691 8931
rect 29749 8897 29783 8931
rect 30678 8773 30712 8807
rect 13060 8598 13122 8698
rect 13122 8598 21822 8698
rect 21822 8598 21884 8698
rect 12960 5064 13060 8400
rect 29140 8665 29156 8698
rect 29156 8665 29188 8698
rect 29140 8650 29188 8665
rect 29246 8652 29294 8700
rect 29382 8699 29430 8700
rect 29382 8665 29389 8699
rect 29389 8665 29423 8699
rect 29423 8665 29430 8699
rect 29382 8652 29430 8665
rect 13490 7864 13674 7898
rect 13948 7864 14132 7898
rect 14406 7864 14590 7898
rect 14864 7864 15048 7898
rect 15322 7864 15506 7898
rect 15780 7864 15964 7898
rect 16238 7864 16422 7898
rect 16696 7864 16880 7898
rect 17154 7864 17338 7898
rect 17612 7864 17796 7898
rect 18070 7864 18254 7898
rect 18528 7864 18712 7898
rect 18986 7864 19170 7898
rect 19444 7864 19628 7898
rect 19902 7864 20086 7898
rect 20360 7864 20544 7898
rect 20818 7864 21002 7898
rect 21276 7864 21460 7898
rect 13336 6229 13370 7805
rect 13794 6229 13828 7805
rect 14252 6229 14286 7805
rect 14710 6229 14744 7805
rect 15168 6229 15202 7805
rect 15626 6229 15660 7805
rect 16084 6229 16118 7805
rect 16542 6229 16576 7805
rect 17000 6229 17034 7805
rect 17458 6229 17492 7805
rect 17916 6229 17950 7805
rect 18374 6229 18408 7805
rect 18832 6229 18866 7805
rect 19290 6229 19324 7805
rect 19748 6229 19782 7805
rect 20206 6229 20240 7805
rect 20664 6229 20698 7805
rect 21122 6229 21156 7805
rect 21580 6229 21614 7805
rect 13490 6136 13674 6170
rect 13948 6136 14132 6170
rect 14406 6136 14590 6170
rect 14864 6136 15048 6170
rect 15322 6136 15506 6170
rect 15780 6136 15964 6170
rect 16238 6136 16422 6170
rect 16696 6136 16880 6170
rect 17154 6136 17338 6170
rect 17612 6136 17796 6170
rect 18070 6136 18254 6170
rect 18528 6136 18712 6170
rect 18986 6136 19170 6170
rect 19444 6136 19628 6170
rect 19902 6136 20086 6170
rect 20360 6136 20544 6170
rect 20818 6136 21002 6170
rect 21276 6136 21460 6170
rect 21884 5064 21984 8400
rect 13060 4766 13122 4866
rect 13122 4766 21822 4866
rect 21822 4766 21884 4866
rect 23642 8518 23704 8618
rect 23704 8518 28824 8618
rect 28824 8518 28886 8618
rect 23542 5049 23642 8335
rect 29738 8652 29786 8700
rect 30580 8665 30628 8700
rect 30580 8652 30584 8665
rect 30584 8652 30618 8665
rect 30618 8652 30628 8665
rect 30757 8705 30791 8739
rect 30832 8594 30880 8642
rect 31098 8781 31132 8807
rect 31098 8773 31100 8781
rect 31100 8773 31132 8781
rect 30995 8705 31029 8739
rect 31412 8773 31446 8807
rect 31499 8705 31533 8739
rect 32242 8632 32290 8680
rect 32358 8665 32406 8680
rect 32358 8632 32380 8665
rect 32380 8632 32406 8665
rect 31936 8546 31948 8562
rect 31948 8546 31982 8562
rect 31982 8546 31984 8562
rect 31936 8514 31984 8546
rect 32470 8632 32518 8680
rect 32602 8665 32650 8680
rect 32712 8665 32760 8680
rect 32828 8665 32876 8680
rect 32602 8632 32613 8665
rect 32613 8632 32647 8665
rect 32647 8632 32650 8665
rect 32712 8632 32739 8665
rect 32739 8632 32760 8665
rect 32828 8632 32873 8665
rect 32873 8632 32876 8665
rect 32960 8630 33008 8678
rect 30239 8399 30273 8433
rect 30581 8399 30615 8433
rect 30673 8399 30707 8433
rect 30765 8399 30799 8433
rect 30857 8399 30891 8433
rect 30949 8399 30983 8433
rect 31041 8399 31075 8433
rect 31133 8399 31167 8433
rect 31225 8399 31259 8433
rect 31317 8399 31351 8433
rect 31409 8399 31443 8433
rect 31501 8399 31535 8433
rect 31593 8399 31627 8433
rect 31685 8399 31719 8433
rect 31777 8399 31811 8433
rect 31869 8399 31903 8433
rect 31961 8399 31995 8433
rect 32053 8399 32087 8433
rect 32145 8399 32179 8433
rect 32237 8399 32271 8433
rect 32329 8399 32363 8433
rect 32421 8399 32455 8433
rect 32513 8399 32547 8433
rect 32605 8399 32639 8433
rect 32697 8399 32731 8433
rect 32789 8399 32823 8433
rect 32881 8399 32915 8433
rect 32973 8399 33007 8433
rect 33139 8399 33173 8433
rect 33279 8399 33313 8433
rect 33371 8399 33405 8433
rect 33463 8399 33497 8433
rect 33555 8399 33589 8433
rect 33647 8399 33681 8433
rect 33739 8399 33773 8433
rect 33831 8399 33865 8433
rect 33923 8399 33957 8433
rect 34015 8399 34049 8433
rect 34107 8399 34141 8433
rect 34199 8399 34233 8433
rect 34291 8399 34325 8433
rect 34383 8399 34417 8433
rect 34475 8399 34509 8433
rect 34567 8399 34601 8433
rect 34659 8399 34693 8433
rect 34751 8399 34785 8433
rect 34843 8399 34877 8433
rect 34935 8399 34969 8433
rect 35027 8399 35061 8433
rect 35119 8399 35153 8433
rect 35211 8399 35245 8433
rect 35303 8399 35337 8433
rect 35395 8399 35429 8433
rect 35487 8399 35521 8433
rect 35579 8399 35613 8433
rect 35671 8399 35705 8433
rect 36013 8399 36047 8433
rect 29105 8353 29139 8387
rect 29197 8353 29231 8387
rect 29289 8353 29323 8387
rect 29381 8353 29415 8387
rect 29473 8353 29507 8387
rect 29565 8353 29599 8387
rect 29657 8353 29691 8387
rect 29749 8353 29783 8387
rect 24085 8284 24269 8318
rect 24543 8284 24727 8318
rect 25001 8284 25185 8318
rect 25459 8284 25643 8318
rect 25917 8284 26101 8318
rect 26375 8284 26559 8318
rect 26833 8284 27017 8318
rect 27291 8284 27475 8318
rect 27749 8284 27933 8318
rect 28207 8284 28391 8318
rect 23931 7049 23965 8225
rect 24389 7049 24423 8225
rect 24847 7049 24881 8225
rect 25305 7049 25339 8225
rect 25763 7049 25797 8225
rect 26221 7049 26255 8225
rect 26679 7049 26713 8225
rect 27137 7049 27171 8225
rect 27595 7049 27629 8225
rect 28053 7049 28087 8225
rect 28511 7049 28545 8225
rect 24085 6956 24269 6990
rect 24543 6956 24727 6990
rect 25001 6956 25185 6990
rect 25459 6956 25643 6990
rect 25917 6956 26101 6990
rect 26375 6956 26559 6990
rect 26833 6956 27017 6990
rect 27291 6956 27475 6990
rect 27749 6956 27933 6990
rect 28207 6956 28391 6990
rect 28886 5049 28986 8335
rect 30576 8167 30584 8190
rect 30584 8167 30618 8190
rect 30618 8167 30624 8190
rect 30576 8142 30624 8167
rect 30678 8025 30712 8059
rect 30757 8093 30791 8127
rect 30832 8190 30880 8238
rect 30995 8093 31029 8127
rect 31098 8051 31100 8059
rect 31100 8051 31132 8059
rect 31098 8025 31132 8051
rect 31412 8025 31446 8059
rect 31499 8093 31533 8127
rect 32242 8152 32290 8200
rect 32358 8167 32380 8200
rect 32380 8167 32406 8200
rect 32358 8152 32406 8167
rect 32470 8152 32518 8200
rect 32602 8167 32613 8200
rect 32613 8167 32647 8200
rect 32647 8167 32650 8200
rect 32712 8167 32739 8200
rect 32739 8167 32760 8200
rect 32828 8167 32873 8200
rect 32873 8167 32876 8200
rect 32602 8152 32650 8167
rect 32712 8152 32760 8167
rect 32828 8152 32876 8167
rect 31936 8005 31946 8016
rect 31946 8005 31980 8016
rect 31980 8005 31984 8016
rect 31936 7971 31984 8005
rect 31936 7968 31946 7971
rect 31946 7968 31980 7971
rect 31980 7968 31984 7971
rect 32964 8154 33012 8202
rect 33274 8100 33322 8148
rect 33376 8025 33410 8059
rect 33455 8093 33489 8127
rect 33530 8190 33578 8238
rect 33693 8093 33727 8127
rect 33796 8051 33798 8059
rect 33798 8051 33830 8059
rect 33796 8025 33830 8051
rect 34110 8025 34144 8059
rect 34197 8093 34231 8127
rect 34636 8286 34684 8314
rect 34636 8266 34646 8286
rect 34646 8266 34680 8286
rect 34680 8266 34684 8286
rect 34940 8152 34988 8200
rect 35056 8167 35078 8200
rect 35078 8167 35104 8200
rect 35056 8152 35104 8167
rect 35168 8152 35216 8200
rect 35300 8167 35311 8200
rect 35311 8167 35345 8200
rect 35345 8167 35348 8200
rect 35410 8167 35437 8200
rect 35437 8167 35458 8200
rect 35526 8167 35571 8200
rect 35571 8167 35574 8200
rect 35300 8152 35348 8167
rect 35410 8152 35458 8167
rect 35526 8152 35574 8167
rect 35658 8154 35706 8202
rect 30239 7855 30273 7889
rect 30581 7855 30615 7889
rect 30673 7855 30707 7889
rect 30765 7855 30799 7889
rect 30857 7855 30891 7889
rect 30949 7855 30983 7889
rect 31041 7855 31075 7889
rect 31133 7855 31167 7889
rect 31225 7855 31259 7889
rect 31317 7855 31351 7889
rect 31409 7855 31443 7889
rect 31501 7855 31535 7889
rect 31593 7855 31627 7889
rect 31685 7855 31719 7889
rect 31777 7855 31811 7889
rect 31869 7855 31903 7889
rect 31961 7855 31995 7889
rect 32053 7855 32087 7889
rect 32145 7855 32179 7889
rect 32237 7855 32271 7889
rect 32329 7855 32363 7889
rect 32421 7855 32455 7889
rect 32513 7855 32547 7889
rect 32605 7855 32639 7889
rect 32697 7855 32731 7889
rect 32789 7855 32823 7889
rect 32881 7855 32915 7889
rect 32973 7855 33007 7889
rect 33279 7855 33313 7889
rect 33371 7855 33405 7889
rect 33463 7855 33497 7889
rect 33555 7855 33589 7889
rect 33647 7855 33681 7889
rect 33739 7855 33773 7889
rect 33831 7855 33865 7889
rect 33923 7855 33957 7889
rect 34015 7855 34049 7889
rect 34107 7855 34141 7889
rect 34199 7855 34233 7889
rect 34291 7855 34325 7889
rect 34383 7855 34417 7889
rect 34475 7855 34509 7889
rect 34567 7855 34601 7889
rect 34659 7855 34693 7889
rect 34751 7855 34785 7889
rect 34843 7855 34877 7889
rect 34935 7855 34969 7889
rect 35027 7855 35061 7889
rect 35119 7855 35153 7889
rect 35211 7855 35245 7889
rect 35303 7855 35337 7889
rect 35395 7855 35429 7889
rect 35487 7855 35521 7889
rect 35579 7855 35613 7889
rect 35671 7855 35705 7889
rect 36013 7855 36047 7889
rect 30678 7685 30712 7719
rect 30576 7596 30624 7644
rect 30757 7617 30791 7651
rect 30832 7506 30880 7554
rect 31098 7693 31132 7719
rect 31098 7685 31100 7693
rect 31100 7685 31132 7693
rect 30995 7617 31029 7651
rect 31412 7685 31446 7719
rect 31499 7617 31533 7651
rect 33376 7685 33410 7719
rect 32242 7544 32290 7592
rect 32358 7577 32406 7592
rect 32358 7544 32380 7577
rect 32380 7544 32406 7577
rect 31936 7458 31948 7472
rect 31948 7458 31982 7472
rect 31982 7458 31984 7472
rect 31936 7424 31984 7458
rect 32470 7544 32518 7592
rect 32602 7577 32650 7592
rect 32712 7577 32760 7592
rect 32828 7577 32876 7592
rect 32602 7544 32613 7577
rect 32613 7544 32647 7577
rect 32647 7544 32650 7577
rect 32712 7544 32739 7577
rect 32739 7544 32760 7577
rect 32828 7544 32873 7577
rect 32873 7544 32876 7577
rect 32960 7542 33012 7590
rect 33274 7577 33322 7604
rect 33274 7556 33282 7577
rect 33282 7556 33316 7577
rect 33316 7556 33322 7577
rect 33455 7617 33489 7651
rect 33530 7506 33578 7554
rect 33796 7693 33830 7719
rect 33796 7685 33798 7693
rect 33798 7685 33830 7693
rect 33693 7617 33727 7651
rect 34110 7685 34144 7719
rect 34197 7617 34231 7651
rect 34634 7773 34644 7776
rect 34644 7773 34678 7776
rect 34678 7773 34682 7776
rect 34634 7739 34682 7773
rect 34634 7728 34644 7739
rect 34644 7728 34678 7739
rect 34678 7728 34682 7739
rect 34940 7544 34988 7592
rect 35056 7577 35104 7592
rect 35056 7544 35078 7577
rect 35078 7544 35104 7577
rect 35168 7544 35216 7592
rect 35300 7577 35348 7592
rect 35410 7577 35458 7592
rect 35526 7577 35574 7592
rect 35300 7544 35311 7577
rect 35311 7544 35345 7577
rect 35345 7544 35348 7577
rect 35410 7544 35437 7577
rect 35437 7544 35458 7577
rect 35526 7544 35571 7577
rect 35571 7544 35574 7577
rect 35658 7542 35706 7590
rect 30239 7311 30273 7345
rect 30581 7311 30615 7345
rect 30673 7311 30707 7345
rect 30765 7311 30799 7345
rect 30857 7311 30891 7345
rect 30949 7311 30983 7345
rect 31041 7311 31075 7345
rect 31133 7311 31167 7345
rect 31225 7311 31259 7345
rect 31317 7311 31351 7345
rect 31409 7311 31443 7345
rect 31501 7311 31535 7345
rect 31593 7311 31627 7345
rect 31685 7311 31719 7345
rect 31777 7311 31811 7345
rect 31869 7311 31903 7345
rect 31961 7311 31995 7345
rect 32053 7311 32087 7345
rect 32145 7311 32179 7345
rect 32237 7311 32271 7345
rect 32329 7311 32363 7345
rect 32421 7311 32455 7345
rect 32513 7311 32547 7345
rect 32605 7311 32639 7345
rect 32697 7311 32731 7345
rect 32789 7311 32823 7345
rect 32881 7311 32915 7345
rect 32973 7311 33007 7345
rect 33279 7311 33313 7345
rect 33371 7311 33405 7345
rect 33463 7311 33497 7345
rect 33555 7311 33589 7345
rect 33647 7311 33681 7345
rect 33739 7311 33773 7345
rect 33831 7311 33865 7345
rect 33923 7311 33957 7345
rect 34015 7311 34049 7345
rect 34107 7311 34141 7345
rect 34199 7311 34233 7345
rect 34291 7311 34325 7345
rect 34383 7311 34417 7345
rect 34475 7311 34509 7345
rect 34567 7311 34601 7345
rect 34659 7311 34693 7345
rect 34751 7311 34785 7345
rect 34843 7311 34877 7345
rect 34935 7311 34969 7345
rect 35027 7311 35061 7345
rect 35119 7311 35153 7345
rect 35211 7311 35245 7345
rect 35303 7311 35337 7345
rect 35395 7311 35429 7345
rect 35487 7311 35521 7345
rect 35579 7311 35613 7345
rect 35671 7311 35705 7345
rect 36013 7311 36047 7345
rect 30576 7079 30584 7100
rect 30584 7079 30618 7100
rect 30618 7079 30624 7100
rect 30576 7052 30624 7079
rect 30678 6937 30712 6971
rect 30757 7005 30791 7039
rect 30832 7102 30880 7150
rect 30995 7005 31029 7039
rect 31098 6963 31100 6971
rect 31100 6963 31132 6971
rect 31098 6937 31132 6963
rect 31412 6937 31446 6971
rect 31499 7005 31533 7039
rect 32242 7064 32290 7112
rect 32358 7079 32380 7112
rect 32380 7079 32406 7112
rect 32358 7064 32406 7079
rect 32470 7064 32518 7112
rect 32602 7079 32613 7112
rect 32613 7079 32647 7112
rect 32647 7079 32650 7112
rect 32712 7079 32739 7112
rect 32739 7079 32760 7112
rect 32828 7079 32873 7112
rect 32873 7079 32876 7112
rect 32602 7064 32650 7079
rect 32712 7064 32760 7079
rect 32828 7064 32876 7079
rect 31936 6917 31946 6928
rect 31946 6917 31980 6928
rect 31980 6917 31984 6928
rect 31936 6883 31984 6917
rect 31936 6880 31946 6883
rect 31946 6880 31980 6883
rect 31980 6880 31984 6883
rect 32960 7066 33008 7114
rect 33274 7012 33322 7060
rect 33376 6937 33410 6971
rect 33455 7005 33489 7039
rect 33530 7102 33578 7150
rect 33693 7005 33727 7039
rect 33796 6963 33798 6971
rect 33798 6963 33830 6971
rect 33796 6937 33830 6963
rect 34110 6937 34144 6971
rect 34197 7005 34231 7039
rect 34634 7198 34682 7232
rect 34634 7184 34646 7198
rect 34646 7184 34680 7198
rect 34680 7184 34682 7198
rect 34940 7064 34988 7112
rect 35056 7079 35078 7112
rect 35078 7079 35104 7112
rect 35056 7064 35104 7079
rect 35168 7064 35216 7112
rect 35300 7079 35311 7112
rect 35311 7079 35345 7112
rect 35345 7079 35348 7112
rect 35410 7079 35437 7112
rect 35437 7079 35458 7112
rect 35526 7079 35571 7112
rect 35571 7079 35574 7112
rect 35300 7064 35348 7079
rect 35410 7064 35458 7079
rect 35526 7064 35574 7079
rect 35658 7066 35710 7114
rect 30239 6767 30273 6801
rect 30581 6767 30615 6801
rect 30673 6767 30707 6801
rect 30765 6767 30799 6801
rect 30857 6767 30891 6801
rect 30949 6767 30983 6801
rect 31041 6767 31075 6801
rect 31133 6767 31167 6801
rect 31225 6767 31259 6801
rect 31317 6767 31351 6801
rect 31409 6767 31443 6801
rect 31501 6767 31535 6801
rect 31593 6767 31627 6801
rect 31685 6767 31719 6801
rect 31777 6767 31811 6801
rect 31869 6767 31903 6801
rect 31961 6767 31995 6801
rect 32053 6767 32087 6801
rect 32145 6767 32179 6801
rect 32237 6767 32271 6801
rect 32329 6767 32363 6801
rect 32421 6767 32455 6801
rect 32513 6767 32547 6801
rect 32605 6767 32639 6801
rect 32697 6767 32731 6801
rect 32789 6767 32823 6801
rect 32881 6767 32915 6801
rect 32973 6767 33007 6801
rect 33279 6767 33313 6801
rect 33371 6767 33405 6801
rect 33463 6767 33497 6801
rect 33555 6767 33589 6801
rect 33647 6767 33681 6801
rect 33739 6767 33773 6801
rect 33831 6767 33865 6801
rect 33923 6767 33957 6801
rect 34015 6767 34049 6801
rect 34107 6767 34141 6801
rect 34199 6767 34233 6801
rect 34291 6767 34325 6801
rect 34383 6767 34417 6801
rect 34475 6767 34509 6801
rect 34567 6767 34601 6801
rect 34659 6767 34693 6801
rect 34751 6767 34785 6801
rect 34843 6767 34877 6801
rect 34935 6767 34969 6801
rect 35027 6767 35061 6801
rect 35119 6767 35153 6801
rect 35211 6767 35245 6801
rect 35303 6767 35337 6801
rect 35395 6767 35429 6801
rect 35487 6767 35521 6801
rect 35579 6767 35613 6801
rect 35671 6767 35705 6801
rect 36013 6767 36047 6801
rect 30678 6597 30712 6631
rect 30576 6508 30624 6556
rect 30757 6529 30791 6563
rect 30832 6418 30880 6466
rect 31098 6605 31132 6631
rect 31098 6597 31100 6605
rect 31100 6597 31132 6605
rect 30995 6529 31029 6563
rect 31412 6597 31446 6631
rect 31499 6529 31533 6563
rect 33376 6597 33410 6631
rect 32242 6456 32290 6504
rect 32358 6489 32406 6504
rect 32358 6456 32380 6489
rect 32380 6456 32406 6489
rect 31936 6370 31948 6386
rect 31948 6370 31982 6386
rect 31982 6370 31984 6386
rect 31936 6338 31984 6370
rect 32470 6456 32518 6504
rect 32602 6489 32650 6504
rect 32712 6489 32760 6504
rect 32828 6489 32876 6504
rect 32602 6456 32613 6489
rect 32613 6456 32647 6489
rect 32647 6456 32650 6489
rect 32712 6456 32739 6489
rect 32739 6456 32760 6489
rect 32828 6456 32873 6489
rect 32873 6456 32876 6489
rect 32960 6454 33008 6502
rect 33274 6489 33322 6514
rect 33274 6466 33282 6489
rect 33282 6466 33316 6489
rect 33316 6466 33322 6489
rect 33455 6529 33489 6563
rect 33530 6418 33578 6466
rect 33796 6605 33830 6631
rect 33796 6597 33798 6605
rect 33798 6597 33830 6605
rect 33693 6529 33727 6563
rect 34110 6597 34144 6631
rect 34197 6529 34231 6563
rect 34634 6685 34644 6688
rect 34644 6685 34678 6688
rect 34678 6685 34682 6688
rect 34634 6651 34682 6685
rect 34634 6640 34644 6651
rect 34644 6640 34678 6651
rect 34678 6640 34682 6651
rect 34940 6456 34988 6504
rect 35056 6489 35104 6504
rect 35056 6456 35078 6489
rect 35078 6456 35104 6489
rect 35168 6456 35216 6504
rect 35300 6489 35348 6504
rect 35410 6489 35458 6504
rect 35526 6489 35574 6504
rect 35300 6456 35311 6489
rect 35311 6456 35345 6489
rect 35345 6456 35348 6489
rect 35410 6456 35437 6489
rect 35437 6456 35458 6489
rect 35526 6456 35571 6489
rect 35571 6456 35574 6489
rect 35662 6454 35710 6502
rect 30239 6223 30273 6257
rect 30581 6223 30615 6257
rect 30673 6223 30707 6257
rect 30765 6223 30799 6257
rect 30857 6223 30891 6257
rect 30949 6223 30983 6257
rect 31041 6223 31075 6257
rect 31133 6223 31167 6257
rect 31225 6223 31259 6257
rect 31317 6223 31351 6257
rect 31409 6223 31443 6257
rect 31501 6223 31535 6257
rect 31593 6223 31627 6257
rect 31685 6223 31719 6257
rect 31777 6223 31811 6257
rect 31869 6223 31903 6257
rect 31961 6223 31995 6257
rect 32053 6223 32087 6257
rect 32145 6223 32179 6257
rect 32237 6223 32271 6257
rect 32329 6223 32363 6257
rect 32421 6223 32455 6257
rect 32513 6223 32547 6257
rect 32605 6223 32639 6257
rect 32697 6223 32731 6257
rect 32789 6223 32823 6257
rect 32881 6223 32915 6257
rect 32973 6223 33007 6257
rect 33279 6223 33313 6257
rect 33371 6223 33405 6257
rect 33463 6223 33497 6257
rect 33555 6223 33589 6257
rect 33647 6223 33681 6257
rect 33739 6223 33773 6257
rect 33831 6223 33865 6257
rect 33923 6223 33957 6257
rect 34015 6223 34049 6257
rect 34107 6223 34141 6257
rect 34199 6223 34233 6257
rect 34291 6223 34325 6257
rect 34383 6223 34417 6257
rect 34475 6223 34509 6257
rect 34567 6223 34601 6257
rect 34659 6223 34693 6257
rect 34751 6223 34785 6257
rect 34843 6223 34877 6257
rect 34935 6223 34969 6257
rect 35027 6223 35061 6257
rect 35119 6223 35153 6257
rect 35211 6223 35245 6257
rect 35303 6223 35337 6257
rect 35395 6223 35429 6257
rect 35487 6223 35521 6257
rect 35579 6223 35613 6257
rect 35671 6223 35705 6257
rect 36013 6223 36047 6257
rect 30576 5991 30584 6014
rect 30584 5991 30618 6014
rect 30618 5991 30624 6014
rect 30576 5966 30624 5991
rect 30678 5849 30712 5883
rect 30757 5917 30791 5951
rect 30832 6014 30880 6062
rect 30995 5917 31029 5951
rect 31098 5875 31100 5883
rect 31100 5875 31132 5883
rect 31098 5849 31132 5875
rect 31412 5849 31446 5883
rect 31499 5917 31533 5951
rect 32242 5976 32290 6024
rect 32358 5991 32380 6024
rect 32380 5991 32406 6024
rect 32358 5976 32406 5991
rect 32470 5976 32518 6024
rect 32602 5991 32613 6024
rect 32613 5991 32647 6024
rect 32647 5991 32650 6024
rect 32712 5991 32739 6024
rect 32739 5991 32760 6024
rect 32828 5991 32873 6024
rect 32873 5991 32876 6024
rect 32602 5976 32650 5991
rect 32712 5976 32760 5991
rect 32828 5976 32876 5991
rect 31936 5829 31946 5842
rect 31946 5829 31980 5842
rect 31980 5829 31984 5842
rect 31936 5795 31984 5829
rect 31936 5794 31946 5795
rect 31946 5794 31980 5795
rect 31980 5794 31984 5795
rect 32960 5978 33012 6026
rect 33282 6025 33330 6032
rect 33282 5991 33316 6025
rect 33316 5991 33330 6025
rect 33282 5984 33330 5991
rect 33376 5849 33410 5883
rect 33455 5917 33489 5951
rect 33530 6014 33578 6062
rect 33693 5917 33727 5951
rect 33796 5875 33798 5883
rect 33798 5875 33830 5883
rect 33796 5849 33830 5875
rect 34110 5849 34144 5883
rect 34197 5917 34231 5951
rect 34634 6110 34682 6142
rect 34634 6094 34646 6110
rect 34646 6094 34680 6110
rect 34680 6094 34682 6110
rect 34940 5976 34988 6024
rect 35056 5991 35078 6024
rect 35078 5991 35104 6024
rect 35056 5976 35104 5991
rect 35168 5976 35216 6024
rect 35300 5991 35311 6024
rect 35311 5991 35345 6024
rect 35345 5991 35348 6024
rect 35410 5991 35437 6024
rect 35437 5991 35458 6024
rect 35526 5991 35571 6024
rect 35571 5991 35574 6024
rect 35300 5976 35348 5991
rect 35410 5976 35458 5991
rect 35526 5976 35574 5991
rect 35658 5978 35706 6026
rect 30239 5679 30273 5713
rect 30581 5679 30615 5713
rect 30673 5679 30707 5713
rect 30765 5679 30799 5713
rect 30857 5679 30891 5713
rect 30949 5679 30983 5713
rect 31041 5679 31075 5713
rect 31133 5679 31167 5713
rect 31225 5679 31259 5713
rect 31317 5679 31351 5713
rect 31409 5679 31443 5713
rect 31501 5679 31535 5713
rect 31593 5679 31627 5713
rect 31685 5679 31719 5713
rect 31777 5679 31811 5713
rect 31869 5679 31903 5713
rect 31961 5679 31995 5713
rect 32053 5679 32087 5713
rect 32145 5679 32179 5713
rect 32237 5679 32271 5713
rect 32329 5679 32363 5713
rect 32421 5679 32455 5713
rect 32513 5679 32547 5713
rect 32605 5679 32639 5713
rect 32697 5679 32731 5713
rect 32789 5679 32823 5713
rect 32881 5679 32915 5713
rect 32973 5679 33007 5713
rect 33279 5679 33313 5713
rect 33371 5679 33405 5713
rect 33463 5679 33497 5713
rect 33555 5679 33589 5713
rect 33647 5679 33681 5713
rect 33739 5679 33773 5713
rect 33831 5679 33865 5713
rect 33923 5679 33957 5713
rect 34015 5679 34049 5713
rect 34107 5679 34141 5713
rect 34199 5679 34233 5713
rect 34291 5679 34325 5713
rect 34383 5679 34417 5713
rect 34475 5679 34509 5713
rect 34567 5679 34601 5713
rect 34659 5679 34693 5713
rect 34751 5679 34785 5713
rect 34843 5679 34877 5713
rect 34935 5679 34969 5713
rect 35027 5679 35061 5713
rect 35119 5679 35153 5713
rect 35211 5679 35245 5713
rect 35303 5679 35337 5713
rect 35395 5679 35429 5713
rect 35487 5679 35521 5713
rect 35579 5679 35613 5713
rect 35671 5679 35705 5713
rect 36013 5679 36047 5713
rect 23642 4766 23704 4866
rect 23704 4766 28824 4866
rect 28824 4766 28886 4866
rect 8452 4296 8514 4396
rect 8514 4296 18634 4396
rect 18634 4296 18696 4396
rect 8352 -1166 8452 4006
rect 9492 2991 9676 3025
rect 9950 2991 10134 3025
rect 10408 2991 10592 3025
rect 10866 2991 11050 3025
rect 11324 2991 11508 3025
rect 11782 2991 11966 3025
rect 12240 2991 12424 3025
rect 12698 2991 12882 3025
rect 13156 2991 13340 3025
rect 13614 2991 13798 3025
rect 14072 2991 14256 3025
rect 14530 2991 14714 3025
rect 14988 2991 15172 3025
rect 15446 2991 15630 3025
rect 15904 2991 16088 3025
rect 16362 2991 16546 3025
rect 16820 2991 17004 3025
rect 17278 2991 17462 3025
rect 9338 1356 9372 2932
rect 9796 1356 9830 2932
rect 10254 1356 10288 2932
rect 10712 1356 10746 2932
rect 11170 1356 11204 2932
rect 11628 1356 11662 2932
rect 12086 1356 12120 2932
rect 12544 1356 12578 2932
rect 13002 1356 13036 2932
rect 13460 1356 13494 2932
rect 13918 1356 13952 2932
rect 14376 1356 14410 2932
rect 14834 1356 14868 2932
rect 15292 1356 15326 2932
rect 15750 1356 15784 2932
rect 16208 1356 16242 2932
rect 16666 1356 16700 2932
rect 17124 1356 17158 2932
rect 17582 1356 17616 2932
rect 9492 1263 9676 1297
rect 9950 1263 10134 1297
rect 10408 1263 10592 1297
rect 10866 1263 11050 1297
rect 11324 1263 11508 1297
rect 11782 1263 11966 1297
rect 12240 1263 12424 1297
rect 12698 1263 12882 1297
rect 13156 1263 13340 1297
rect 13614 1263 13798 1297
rect 14072 1263 14256 1297
rect 14530 1263 14714 1297
rect 14988 1263 15172 1297
rect 15446 1263 15630 1297
rect 15904 1263 16088 1297
rect 16362 1263 16546 1297
rect 16820 1263 17004 1297
rect 17278 1263 17462 1297
rect 13222 1132 13270 1180
rect 13676 1126 13736 1186
rect 8933 326 9117 360
rect 9391 326 9575 360
rect 9849 326 10033 360
rect 10307 326 10491 360
rect 10765 326 10949 360
rect 11223 326 11407 360
rect 11681 326 11865 360
rect 12139 326 12323 360
rect 12597 326 12781 360
rect 13055 326 13239 360
rect 13933 326 14117 360
rect 14391 326 14575 360
rect 14849 326 15033 360
rect 15307 326 15491 360
rect 15765 326 15949 360
rect 16223 326 16407 360
rect 16681 326 16865 360
rect 17139 326 17323 360
rect 17597 326 17781 360
rect 18055 326 18239 360
rect 8779 -909 8813 267
rect 9237 -909 9271 267
rect 9695 -909 9729 267
rect 10153 -909 10187 267
rect 10611 -909 10645 267
rect 11069 -909 11103 267
rect 11527 -909 11561 267
rect 11985 -909 12019 267
rect 12443 -909 12477 267
rect 12901 -909 12935 267
rect 13359 -909 13393 267
rect 13779 -909 13813 267
rect 14237 -909 14271 267
rect 14695 -909 14729 267
rect 15153 -909 15187 267
rect 15611 -909 15645 267
rect 16069 -909 16103 267
rect 16527 -909 16561 267
rect 16985 -909 17019 267
rect 17443 -909 17477 267
rect 17901 -909 17935 267
rect 18359 -909 18393 267
rect 8933 -1002 9117 -968
rect 9391 -1002 9575 -968
rect 9849 -1002 10033 -968
rect 10307 -1002 10491 -968
rect 10765 -1002 10949 -968
rect 11223 -1002 11407 -968
rect 11681 -1002 11865 -968
rect 12139 -1002 12323 -968
rect 12597 -1002 12781 -968
rect 13055 -1002 13239 -968
rect 13933 -1002 14117 -968
rect 14391 -1002 14575 -968
rect 14849 -1002 15033 -968
rect 15307 -1002 15491 -968
rect 15765 -1002 15949 -968
rect 16223 -1002 16407 -968
rect 16681 -1002 16865 -968
rect 17139 -1002 17323 -968
rect 17597 -1002 17781 -968
rect 18055 -1002 18239 -968
rect 18696 -1166 18796 4006
rect 8452 -1448 8514 -1348
rect 8514 -1448 18634 -1348
rect 18634 -1448 18696 -1348
rect 23452 4296 23514 4396
rect 23514 4296 33634 4396
rect 33634 4296 33696 4396
rect 23352 -1166 23452 4006
rect 24492 2991 24676 3025
rect 24950 2991 25134 3025
rect 25408 2991 25592 3025
rect 25866 2991 26050 3025
rect 26324 2991 26508 3025
rect 26782 2991 26966 3025
rect 27240 2991 27424 3025
rect 27698 2991 27882 3025
rect 28156 2991 28340 3025
rect 28614 2991 28798 3025
rect 29072 2991 29256 3025
rect 29530 2991 29714 3025
rect 29988 2991 30172 3025
rect 30446 2991 30630 3025
rect 30904 2991 31088 3025
rect 31362 2991 31546 3025
rect 31820 2991 32004 3025
rect 32278 2991 32462 3025
rect 24338 1356 24372 2932
rect 24796 1356 24830 2932
rect 25254 1356 25288 2932
rect 25712 1356 25746 2932
rect 26170 1356 26204 2932
rect 26628 1356 26662 2932
rect 27086 1356 27120 2932
rect 27544 1356 27578 2932
rect 28002 1356 28036 2932
rect 28460 1356 28494 2932
rect 28918 1356 28952 2932
rect 29376 1356 29410 2932
rect 29834 1356 29868 2932
rect 30292 1356 30326 2932
rect 30750 1356 30784 2932
rect 31208 1356 31242 2932
rect 31666 1356 31700 2932
rect 32124 1356 32158 2932
rect 32582 1356 32616 2932
rect 24492 1263 24676 1297
rect 24950 1263 25134 1297
rect 25408 1263 25592 1297
rect 25866 1263 26050 1297
rect 26324 1263 26508 1297
rect 26782 1263 26966 1297
rect 27240 1263 27424 1297
rect 27698 1263 27882 1297
rect 28156 1263 28340 1297
rect 28614 1263 28798 1297
rect 29072 1263 29256 1297
rect 29530 1263 29714 1297
rect 29988 1263 30172 1297
rect 30446 1263 30630 1297
rect 30904 1263 31088 1297
rect 31362 1263 31546 1297
rect 31820 1263 32004 1297
rect 32278 1263 32462 1297
rect 28222 1132 28270 1180
rect 28676 1126 28736 1186
rect 23933 326 24117 360
rect 24391 326 24575 360
rect 24849 326 25033 360
rect 25307 326 25491 360
rect 25765 326 25949 360
rect 26223 326 26407 360
rect 26681 326 26865 360
rect 27139 326 27323 360
rect 27597 326 27781 360
rect 28055 326 28239 360
rect 28933 326 29117 360
rect 29391 326 29575 360
rect 29849 326 30033 360
rect 30307 326 30491 360
rect 30765 326 30949 360
rect 31223 326 31407 360
rect 31681 326 31865 360
rect 32139 326 32323 360
rect 32597 326 32781 360
rect 33055 326 33239 360
rect 23779 -909 23813 267
rect 24237 -909 24271 267
rect 24695 -909 24729 267
rect 25153 -909 25187 267
rect 25611 -909 25645 267
rect 26069 -909 26103 267
rect 26527 -909 26561 267
rect 26985 -909 27019 267
rect 27443 -909 27477 267
rect 27901 -909 27935 267
rect 28359 -909 28393 267
rect 28779 -909 28813 267
rect 29237 -909 29271 267
rect 29695 -909 29729 267
rect 30153 -909 30187 267
rect 30611 -909 30645 267
rect 31069 -909 31103 267
rect 31527 -909 31561 267
rect 31985 -909 32019 267
rect 32443 -909 32477 267
rect 32901 -909 32935 267
rect 33359 -909 33393 267
rect 23933 -1002 24117 -968
rect 24391 -1002 24575 -968
rect 24849 -1002 25033 -968
rect 25307 -1002 25491 -968
rect 25765 -1002 25949 -968
rect 26223 -1002 26407 -968
rect 26681 -1002 26865 -968
rect 27139 -1002 27323 -968
rect 27597 -1002 27781 -968
rect 28055 -1002 28239 -968
rect 28933 -1002 29117 -968
rect 29391 -1002 29575 -968
rect 29849 -1002 30033 -968
rect 30307 -1002 30491 -968
rect 30765 -1002 30949 -968
rect 31223 -1002 31407 -968
rect 31681 -1002 31865 -968
rect 32139 -1002 32323 -968
rect 32597 -1002 32781 -968
rect 33055 -1002 33239 -968
rect 33696 -1166 33796 4006
rect 23452 -1448 23514 -1348
rect 23514 -1448 33634 -1348
rect 33634 -1448 33696 -1348
rect 8452 -1784 8514 -1684
rect 8514 -1784 18634 -1684
rect 18634 -1784 18696 -1684
rect 8352 -3918 8452 -1914
rect 8932 -2176 9116 -2142
rect 9390 -2176 9574 -2142
rect 9848 -2176 10032 -2142
rect 10306 -2176 10490 -2142
rect 10764 -2176 10948 -2142
rect 11222 -2176 11406 -2142
rect 11680 -2176 11864 -2142
rect 12138 -2176 12322 -2142
rect 12596 -2176 12780 -2142
rect 13054 -2176 13238 -2142
rect 13932 -2176 14116 -2142
rect 14390 -2176 14574 -2142
rect 14848 -2176 15032 -2142
rect 15306 -2176 15490 -2142
rect 15764 -2176 15948 -2142
rect 16222 -2176 16406 -2142
rect 16680 -2176 16864 -2142
rect 17138 -2176 17322 -2142
rect 17596 -2176 17780 -2142
rect 18054 -2176 18238 -2142
rect 8778 -2402 8812 -2226
rect 9236 -2402 9270 -2226
rect 9694 -2402 9728 -2226
rect 10152 -2402 10186 -2226
rect 10610 -2402 10644 -2226
rect 11068 -2402 11102 -2226
rect 11526 -2402 11560 -2226
rect 11984 -2402 12018 -2226
rect 12442 -2402 12476 -2226
rect 12900 -2402 12934 -2226
rect 13358 -2402 13392 -2226
rect 13778 -2402 13812 -2226
rect 14236 -2402 14270 -2226
rect 14694 -2402 14728 -2226
rect 15152 -2402 15186 -2226
rect 15610 -2402 15644 -2226
rect 16068 -2402 16102 -2226
rect 16526 -2402 16560 -2226
rect 16984 -2402 17018 -2226
rect 17442 -2402 17476 -2226
rect 17900 -2402 17934 -2226
rect 18358 -2402 18392 -2226
rect 8932 -2486 9116 -2452
rect 9390 -2486 9574 -2452
rect 9848 -2486 10032 -2452
rect 10306 -2486 10490 -2452
rect 10764 -2486 10948 -2452
rect 11222 -2486 11406 -2452
rect 11680 -2486 11864 -2452
rect 12138 -2486 12322 -2452
rect 12596 -2486 12780 -2452
rect 13054 -2486 13238 -2452
rect 13932 -2486 14116 -2452
rect 14390 -2486 14574 -2452
rect 14848 -2486 15032 -2452
rect 15306 -2486 15490 -2452
rect 15764 -2486 15948 -2452
rect 16222 -2486 16406 -2452
rect 16680 -2486 16864 -2452
rect 17138 -2486 17322 -2452
rect 17596 -2486 17780 -2452
rect 18054 -2486 18238 -2452
rect 8932 -2844 9116 -2810
rect 9390 -2844 9574 -2810
rect 9848 -2844 10032 -2810
rect 10306 -2844 10490 -2810
rect 10764 -2844 10948 -2810
rect 11222 -2844 11406 -2810
rect 11680 -2844 11864 -2810
rect 12138 -2844 12322 -2810
rect 12596 -2844 12780 -2810
rect 13054 -2844 13238 -2810
rect 8778 -3070 8812 -2894
rect 9236 -3070 9270 -2894
rect 9694 -3070 9728 -2894
rect 10152 -3070 10186 -2894
rect 10610 -3070 10644 -2894
rect 11068 -3070 11102 -2894
rect 11526 -3070 11560 -2894
rect 11984 -3070 12018 -2894
rect 12442 -3070 12476 -2894
rect 12900 -3070 12934 -2894
rect 13358 -3070 13392 -2894
rect 8932 -3154 9116 -3120
rect 9390 -3154 9574 -3120
rect 9848 -3154 10032 -3120
rect 10306 -3154 10490 -3120
rect 10764 -3154 10948 -3120
rect 11222 -3154 11406 -3120
rect 11680 -3154 11864 -3120
rect 12138 -3154 12322 -3120
rect 12596 -3154 12780 -3120
rect 13054 -3154 13238 -3120
rect 18696 -3918 18796 -1914
rect 8452 -4148 8514 -4048
rect 8514 -4148 18634 -4048
rect 18634 -4148 18696 -4048
rect 23452 -1784 23514 -1684
rect 23514 -1784 33634 -1684
rect 33634 -1784 33696 -1684
rect 23352 -3918 23452 -1914
rect 23932 -2176 24116 -2142
rect 24390 -2176 24574 -2142
rect 24848 -2176 25032 -2142
rect 25306 -2176 25490 -2142
rect 25764 -2176 25948 -2142
rect 26222 -2176 26406 -2142
rect 26680 -2176 26864 -2142
rect 27138 -2176 27322 -2142
rect 27596 -2176 27780 -2142
rect 28054 -2176 28238 -2142
rect 28932 -2176 29116 -2142
rect 29390 -2176 29574 -2142
rect 29848 -2176 30032 -2142
rect 30306 -2176 30490 -2142
rect 30764 -2176 30948 -2142
rect 31222 -2176 31406 -2142
rect 31680 -2176 31864 -2142
rect 32138 -2176 32322 -2142
rect 32596 -2176 32780 -2142
rect 33054 -2176 33238 -2142
rect 23778 -2402 23812 -2226
rect 24236 -2402 24270 -2226
rect 24694 -2402 24728 -2226
rect 25152 -2402 25186 -2226
rect 25610 -2402 25644 -2226
rect 26068 -2402 26102 -2226
rect 26526 -2402 26560 -2226
rect 26984 -2402 27018 -2226
rect 27442 -2402 27476 -2226
rect 27900 -2402 27934 -2226
rect 28358 -2402 28392 -2226
rect 28778 -2402 28812 -2226
rect 29236 -2402 29270 -2226
rect 29694 -2402 29728 -2226
rect 30152 -2402 30186 -2226
rect 30610 -2402 30644 -2226
rect 31068 -2402 31102 -2226
rect 31526 -2402 31560 -2226
rect 31984 -2402 32018 -2226
rect 32442 -2402 32476 -2226
rect 32900 -2402 32934 -2226
rect 33358 -2402 33392 -2226
rect 23932 -2486 24116 -2452
rect 24390 -2486 24574 -2452
rect 24848 -2486 25032 -2452
rect 25306 -2486 25490 -2452
rect 25764 -2486 25948 -2452
rect 26222 -2486 26406 -2452
rect 26680 -2486 26864 -2452
rect 27138 -2486 27322 -2452
rect 27596 -2486 27780 -2452
rect 28054 -2486 28238 -2452
rect 28932 -2486 29116 -2452
rect 29390 -2486 29574 -2452
rect 29848 -2486 30032 -2452
rect 30306 -2486 30490 -2452
rect 30764 -2486 30948 -2452
rect 31222 -2486 31406 -2452
rect 31680 -2486 31864 -2452
rect 32138 -2486 32322 -2452
rect 32596 -2486 32780 -2452
rect 33054 -2486 33238 -2452
rect 23932 -2844 24116 -2810
rect 24390 -2844 24574 -2810
rect 24848 -2844 25032 -2810
rect 25306 -2844 25490 -2810
rect 25764 -2844 25948 -2810
rect 26222 -2844 26406 -2810
rect 26680 -2844 26864 -2810
rect 27138 -2844 27322 -2810
rect 27596 -2844 27780 -2810
rect 28054 -2844 28238 -2810
rect 23778 -3070 23812 -2894
rect 24236 -3070 24270 -2894
rect 24694 -3070 24728 -2894
rect 25152 -3070 25186 -2894
rect 25610 -3070 25644 -2894
rect 26068 -3070 26102 -2894
rect 26526 -3070 26560 -2894
rect 26984 -3070 27018 -2894
rect 27442 -3070 27476 -2894
rect 27900 -3070 27934 -2894
rect 28358 -3070 28392 -2894
rect 23932 -3154 24116 -3120
rect 24390 -3154 24574 -3120
rect 24848 -3154 25032 -3120
rect 25306 -3154 25490 -3120
rect 25764 -3154 25948 -3120
rect 26222 -3154 26406 -3120
rect 26680 -3154 26864 -3120
rect 27138 -3154 27322 -3120
rect 27596 -3154 27780 -3120
rect 28054 -3154 28238 -3120
rect 33696 -3918 33796 -1914
rect 23452 -4148 23514 -4048
rect 23514 -4148 33634 -4048
rect 33634 -4148 33696 -4048
rect 12406 -4708 12468 -4608
rect 12468 -4708 22588 -4608
rect 22588 -4708 22650 -4608
rect 12306 -6842 12406 -4838
rect 17864 -5636 18048 -5602
rect 18322 -5636 18506 -5602
rect 18780 -5636 18964 -5602
rect 19238 -5636 19422 -5602
rect 19696 -5636 19880 -5602
rect 20154 -5636 20338 -5602
rect 20612 -5636 20796 -5602
rect 21070 -5636 21254 -5602
rect 21528 -5636 21712 -5602
rect 21986 -5636 22170 -5602
rect 17710 -5862 17744 -5686
rect 18168 -5862 18202 -5686
rect 18626 -5862 18660 -5686
rect 19084 -5862 19118 -5686
rect 19542 -5862 19576 -5686
rect 20000 -5862 20034 -5686
rect 20458 -5862 20492 -5686
rect 20916 -5862 20950 -5686
rect 21374 -5862 21408 -5686
rect 21832 -5862 21866 -5686
rect 22290 -5862 22324 -5686
rect 17864 -5946 18048 -5912
rect 18322 -5946 18506 -5912
rect 18780 -5946 18964 -5912
rect 19238 -5946 19422 -5912
rect 19696 -5946 19880 -5912
rect 20154 -5946 20338 -5912
rect 20612 -5946 20796 -5912
rect 21070 -5946 21254 -5912
rect 21528 -5946 21712 -5912
rect 21986 -5946 22170 -5912
rect 12864 -6304 13048 -6270
rect 13322 -6304 13506 -6270
rect 13780 -6304 13964 -6270
rect 14238 -6304 14422 -6270
rect 14696 -6304 14880 -6270
rect 15154 -6304 15338 -6270
rect 15612 -6304 15796 -6270
rect 16070 -6304 16254 -6270
rect 16528 -6304 16712 -6270
rect 16986 -6304 17170 -6270
rect 17864 -6304 18048 -6270
rect 18322 -6304 18506 -6270
rect 18780 -6304 18964 -6270
rect 19238 -6304 19422 -6270
rect 19696 -6304 19880 -6270
rect 20154 -6304 20338 -6270
rect 20612 -6304 20796 -6270
rect 21070 -6304 21254 -6270
rect 21528 -6304 21712 -6270
rect 21986 -6304 22170 -6270
rect 12710 -6530 12744 -6354
rect 13168 -6530 13202 -6354
rect 13626 -6530 13660 -6354
rect 14084 -6530 14118 -6354
rect 14542 -6530 14576 -6354
rect 15000 -6530 15034 -6354
rect 15458 -6530 15492 -6354
rect 15916 -6530 15950 -6354
rect 16374 -6530 16408 -6354
rect 16832 -6530 16866 -6354
rect 17290 -6530 17324 -6354
rect 17710 -6530 17744 -6354
rect 18168 -6530 18202 -6354
rect 18626 -6530 18660 -6354
rect 19084 -6530 19118 -6354
rect 19542 -6530 19576 -6354
rect 20000 -6530 20034 -6354
rect 20458 -6530 20492 -6354
rect 20916 -6530 20950 -6354
rect 21374 -6530 21408 -6354
rect 21832 -6530 21866 -6354
rect 22290 -6530 22324 -6354
rect 12864 -6614 13048 -6580
rect 13322 -6614 13506 -6580
rect 13780 -6614 13964 -6580
rect 14238 -6614 14422 -6580
rect 14696 -6614 14880 -6580
rect 15154 -6614 15338 -6580
rect 15612 -6614 15796 -6580
rect 16070 -6614 16254 -6580
rect 16528 -6614 16712 -6580
rect 16986 -6614 17170 -6580
rect 17864 -6614 18048 -6580
rect 18322 -6614 18506 -6580
rect 18780 -6614 18964 -6580
rect 19238 -6614 19422 -6580
rect 19696 -6614 19880 -6580
rect 20154 -6614 20338 -6580
rect 20612 -6614 20796 -6580
rect 21070 -6614 21254 -6580
rect 21528 -6614 21712 -6580
rect 21986 -6614 22170 -6580
rect 22650 -6842 22750 -4838
rect 12406 -7072 12468 -6972
rect 12468 -7072 22588 -6972
rect 22588 -7072 22650 -6972
rect 27406 -4708 27468 -4608
rect 27468 -4708 37588 -4608
rect 37588 -4708 37650 -4608
rect 27306 -6842 27406 -4838
rect 32864 -5636 33048 -5602
rect 33322 -5636 33506 -5602
rect 33780 -5636 33964 -5602
rect 34238 -5636 34422 -5602
rect 34696 -5636 34880 -5602
rect 35154 -5636 35338 -5602
rect 35612 -5636 35796 -5602
rect 36070 -5636 36254 -5602
rect 36528 -5636 36712 -5602
rect 36986 -5636 37170 -5602
rect 32710 -5862 32744 -5686
rect 33168 -5862 33202 -5686
rect 33626 -5862 33660 -5686
rect 34084 -5862 34118 -5686
rect 34542 -5862 34576 -5686
rect 35000 -5862 35034 -5686
rect 35458 -5862 35492 -5686
rect 35916 -5862 35950 -5686
rect 36374 -5862 36408 -5686
rect 36832 -5862 36866 -5686
rect 37290 -5862 37324 -5686
rect 32864 -5946 33048 -5912
rect 33322 -5946 33506 -5912
rect 33780 -5946 33964 -5912
rect 34238 -5946 34422 -5912
rect 34696 -5946 34880 -5912
rect 35154 -5946 35338 -5912
rect 35612 -5946 35796 -5912
rect 36070 -5946 36254 -5912
rect 36528 -5946 36712 -5912
rect 36986 -5946 37170 -5912
rect 27864 -6304 28048 -6270
rect 28322 -6304 28506 -6270
rect 28780 -6304 28964 -6270
rect 29238 -6304 29422 -6270
rect 29696 -6304 29880 -6270
rect 30154 -6304 30338 -6270
rect 30612 -6304 30796 -6270
rect 31070 -6304 31254 -6270
rect 31528 -6304 31712 -6270
rect 31986 -6304 32170 -6270
rect 32864 -6304 33048 -6270
rect 33322 -6304 33506 -6270
rect 33780 -6304 33964 -6270
rect 34238 -6304 34422 -6270
rect 34696 -6304 34880 -6270
rect 35154 -6304 35338 -6270
rect 35612 -6304 35796 -6270
rect 36070 -6304 36254 -6270
rect 36528 -6304 36712 -6270
rect 36986 -6304 37170 -6270
rect 27710 -6530 27744 -6354
rect 28168 -6530 28202 -6354
rect 28626 -6530 28660 -6354
rect 29084 -6530 29118 -6354
rect 29542 -6530 29576 -6354
rect 30000 -6530 30034 -6354
rect 30458 -6530 30492 -6354
rect 30916 -6530 30950 -6354
rect 31374 -6530 31408 -6354
rect 31832 -6530 31866 -6354
rect 32290 -6530 32324 -6354
rect 32710 -6530 32744 -6354
rect 33168 -6530 33202 -6354
rect 33626 -6530 33660 -6354
rect 34084 -6530 34118 -6354
rect 34542 -6530 34576 -6354
rect 35000 -6530 35034 -6354
rect 35458 -6530 35492 -6354
rect 35916 -6530 35950 -6354
rect 36374 -6530 36408 -6354
rect 36832 -6530 36866 -6354
rect 37290 -6530 37324 -6354
rect 27864 -6614 28048 -6580
rect 28322 -6614 28506 -6580
rect 28780 -6614 28964 -6580
rect 29238 -6614 29422 -6580
rect 29696 -6614 29880 -6580
rect 30154 -6614 30338 -6580
rect 30612 -6614 30796 -6580
rect 31070 -6614 31254 -6580
rect 31528 -6614 31712 -6580
rect 31986 -6614 32170 -6580
rect 32864 -6614 33048 -6580
rect 33322 -6614 33506 -6580
rect 33780 -6614 33964 -6580
rect 34238 -6614 34422 -6580
rect 34696 -6614 34880 -6580
rect 35154 -6614 35338 -6580
rect 35612 -6614 35796 -6580
rect 36070 -6614 36254 -6580
rect 36528 -6614 36712 -6580
rect 36986 -6614 37170 -6580
rect 37650 -6842 37750 -4838
rect 27406 -7072 27468 -6972
rect 27468 -7072 37588 -6972
rect 37588 -7072 37650 -6972
rect 12406 -7408 12468 -7308
rect 12468 -7408 22588 -7308
rect 22588 -7408 22650 -7308
rect 12306 -12762 12406 -7590
rect 12863 -7788 13047 -7754
rect 13321 -7788 13505 -7754
rect 13779 -7788 13963 -7754
rect 14237 -7788 14421 -7754
rect 14695 -7788 14879 -7754
rect 15153 -7788 15337 -7754
rect 15611 -7788 15795 -7754
rect 16069 -7788 16253 -7754
rect 16527 -7788 16711 -7754
rect 16985 -7788 17169 -7754
rect 17863 -7788 18047 -7754
rect 18321 -7788 18505 -7754
rect 18779 -7788 18963 -7754
rect 19237 -7788 19421 -7754
rect 19695 -7788 19879 -7754
rect 20153 -7788 20337 -7754
rect 20611 -7788 20795 -7754
rect 21069 -7788 21253 -7754
rect 21527 -7788 21711 -7754
rect 21985 -7788 22169 -7754
rect 12709 -9023 12743 -7847
rect 13167 -9023 13201 -7847
rect 13625 -9023 13659 -7847
rect 14083 -9023 14117 -7847
rect 14541 -9023 14575 -7847
rect 14999 -9023 15033 -7847
rect 15457 -9023 15491 -7847
rect 15915 -9023 15949 -7847
rect 16373 -9023 16407 -7847
rect 16831 -9023 16865 -7847
rect 17289 -9023 17323 -7847
rect 17709 -9023 17743 -7847
rect 18167 -9023 18201 -7847
rect 18625 -9023 18659 -7847
rect 19083 -9023 19117 -7847
rect 19541 -9023 19575 -7847
rect 19999 -9023 20033 -7847
rect 20457 -9023 20491 -7847
rect 20915 -9023 20949 -7847
rect 21373 -9023 21407 -7847
rect 21831 -9023 21865 -7847
rect 22289 -9023 22323 -7847
rect 12863 -9116 13047 -9082
rect 13321 -9116 13505 -9082
rect 13779 -9116 13963 -9082
rect 14237 -9116 14421 -9082
rect 14695 -9116 14879 -9082
rect 15153 -9116 15337 -9082
rect 15611 -9116 15795 -9082
rect 16069 -9116 16253 -9082
rect 16527 -9116 16711 -9082
rect 16985 -9116 17169 -9082
rect 17863 -9116 18047 -9082
rect 18321 -9116 18505 -9082
rect 18779 -9116 18963 -9082
rect 19237 -9116 19421 -9082
rect 19695 -9116 19879 -9082
rect 20153 -9116 20337 -9082
rect 20611 -9116 20795 -9082
rect 21069 -9116 21253 -9082
rect 21527 -9116 21711 -9082
rect 21985 -9116 22169 -9082
rect 17366 -9942 17426 -9882
rect 17832 -9936 17880 -9888
rect 13640 -10053 13824 -10019
rect 14098 -10053 14282 -10019
rect 14556 -10053 14740 -10019
rect 15014 -10053 15198 -10019
rect 15472 -10053 15656 -10019
rect 15930 -10053 16114 -10019
rect 16388 -10053 16572 -10019
rect 16846 -10053 17030 -10019
rect 17304 -10053 17488 -10019
rect 17762 -10053 17946 -10019
rect 18220 -10053 18404 -10019
rect 18678 -10053 18862 -10019
rect 19136 -10053 19320 -10019
rect 19594 -10053 19778 -10019
rect 20052 -10053 20236 -10019
rect 20510 -10053 20694 -10019
rect 20968 -10053 21152 -10019
rect 21426 -10053 21610 -10019
rect 13486 -11688 13520 -10112
rect 13944 -11688 13978 -10112
rect 14402 -11688 14436 -10112
rect 14860 -11688 14894 -10112
rect 15318 -11688 15352 -10112
rect 15776 -11688 15810 -10112
rect 16234 -11688 16268 -10112
rect 16692 -11688 16726 -10112
rect 17150 -11688 17184 -10112
rect 17608 -11688 17642 -10112
rect 18066 -11688 18100 -10112
rect 18524 -11688 18558 -10112
rect 18982 -11688 19016 -10112
rect 19440 -11688 19474 -10112
rect 19898 -11688 19932 -10112
rect 20356 -11688 20390 -10112
rect 20814 -11688 20848 -10112
rect 21272 -11688 21306 -10112
rect 21730 -11688 21764 -10112
rect 13640 -11781 13824 -11747
rect 14098 -11781 14282 -11747
rect 14556 -11781 14740 -11747
rect 15014 -11781 15198 -11747
rect 15472 -11781 15656 -11747
rect 15930 -11781 16114 -11747
rect 16388 -11781 16572 -11747
rect 16846 -11781 17030 -11747
rect 17304 -11781 17488 -11747
rect 17762 -11781 17946 -11747
rect 18220 -11781 18404 -11747
rect 18678 -11781 18862 -11747
rect 19136 -11781 19320 -11747
rect 19594 -11781 19778 -11747
rect 20052 -11781 20236 -11747
rect 20510 -11781 20694 -11747
rect 20968 -11781 21152 -11747
rect 21426 -11781 21610 -11747
rect 22650 -12762 22750 -7590
rect 12406 -13152 12468 -13052
rect 12468 -13152 22588 -13052
rect 22588 -13152 22650 -13052
rect 27406 -7408 27468 -7308
rect 27468 -7408 37588 -7308
rect 37588 -7408 37650 -7308
rect 27306 -12762 27406 -7590
rect 27863 -7788 28047 -7754
rect 28321 -7788 28505 -7754
rect 28779 -7788 28963 -7754
rect 29237 -7788 29421 -7754
rect 29695 -7788 29879 -7754
rect 30153 -7788 30337 -7754
rect 30611 -7788 30795 -7754
rect 31069 -7788 31253 -7754
rect 31527 -7788 31711 -7754
rect 31985 -7788 32169 -7754
rect 32863 -7788 33047 -7754
rect 33321 -7788 33505 -7754
rect 33779 -7788 33963 -7754
rect 34237 -7788 34421 -7754
rect 34695 -7788 34879 -7754
rect 35153 -7788 35337 -7754
rect 35611 -7788 35795 -7754
rect 36069 -7788 36253 -7754
rect 36527 -7788 36711 -7754
rect 36985 -7788 37169 -7754
rect 27709 -9023 27743 -7847
rect 28167 -9023 28201 -7847
rect 28625 -9023 28659 -7847
rect 29083 -9023 29117 -7847
rect 29541 -9023 29575 -7847
rect 29999 -9023 30033 -7847
rect 30457 -9023 30491 -7847
rect 30915 -9023 30949 -7847
rect 31373 -9023 31407 -7847
rect 31831 -9023 31865 -7847
rect 32289 -9023 32323 -7847
rect 32709 -9023 32743 -7847
rect 33167 -9023 33201 -7847
rect 33625 -9023 33659 -7847
rect 34083 -9023 34117 -7847
rect 34541 -9023 34575 -7847
rect 34999 -9023 35033 -7847
rect 35457 -9023 35491 -7847
rect 35915 -9023 35949 -7847
rect 36373 -9023 36407 -7847
rect 36831 -9023 36865 -7847
rect 37289 -9023 37323 -7847
rect 27863 -9116 28047 -9082
rect 28321 -9116 28505 -9082
rect 28779 -9116 28963 -9082
rect 29237 -9116 29421 -9082
rect 29695 -9116 29879 -9082
rect 30153 -9116 30337 -9082
rect 30611 -9116 30795 -9082
rect 31069 -9116 31253 -9082
rect 31527 -9116 31711 -9082
rect 31985 -9116 32169 -9082
rect 32863 -9116 33047 -9082
rect 33321 -9116 33505 -9082
rect 33779 -9116 33963 -9082
rect 34237 -9116 34421 -9082
rect 34695 -9116 34879 -9082
rect 35153 -9116 35337 -9082
rect 35611 -9116 35795 -9082
rect 36069 -9116 36253 -9082
rect 36527 -9116 36711 -9082
rect 36985 -9116 37169 -9082
rect 32366 -9942 32426 -9882
rect 32832 -9936 32880 -9888
rect 28640 -10053 28824 -10019
rect 29098 -10053 29282 -10019
rect 29556 -10053 29740 -10019
rect 30014 -10053 30198 -10019
rect 30472 -10053 30656 -10019
rect 30930 -10053 31114 -10019
rect 31388 -10053 31572 -10019
rect 31846 -10053 32030 -10019
rect 32304 -10053 32488 -10019
rect 32762 -10053 32946 -10019
rect 33220 -10053 33404 -10019
rect 33678 -10053 33862 -10019
rect 34136 -10053 34320 -10019
rect 34594 -10053 34778 -10019
rect 35052 -10053 35236 -10019
rect 35510 -10053 35694 -10019
rect 35968 -10053 36152 -10019
rect 36426 -10053 36610 -10019
rect 28486 -11688 28520 -10112
rect 28944 -11688 28978 -10112
rect 29402 -11688 29436 -10112
rect 29860 -11688 29894 -10112
rect 30318 -11688 30352 -10112
rect 30776 -11688 30810 -10112
rect 31234 -11688 31268 -10112
rect 31692 -11688 31726 -10112
rect 32150 -11688 32184 -10112
rect 32608 -11688 32642 -10112
rect 33066 -11688 33100 -10112
rect 33524 -11688 33558 -10112
rect 33982 -11688 34016 -10112
rect 34440 -11688 34474 -10112
rect 34898 -11688 34932 -10112
rect 35356 -11688 35390 -10112
rect 35814 -11688 35848 -10112
rect 36272 -11688 36306 -10112
rect 36730 -11688 36764 -10112
rect 28640 -11781 28824 -11747
rect 29098 -11781 29282 -11747
rect 29556 -11781 29740 -11747
rect 30014 -11781 30198 -11747
rect 30472 -11781 30656 -11747
rect 30930 -11781 31114 -11747
rect 31388 -11781 31572 -11747
rect 31846 -11781 32030 -11747
rect 32304 -11781 32488 -11747
rect 32762 -11781 32946 -11747
rect 33220 -11781 33404 -11747
rect 33678 -11781 33862 -11747
rect 34136 -11781 34320 -11747
rect 34594 -11781 34778 -11747
rect 35052 -11781 35236 -11747
rect 35510 -11781 35694 -11747
rect 35968 -11781 36152 -11747
rect 36426 -11781 36610 -11747
rect 37650 -12762 37750 -7590
rect 27406 -13152 27468 -13052
rect 27468 -13152 37588 -13052
rect 37588 -13152 37650 -13052
rect 8452 -13704 8514 -13604
rect 8514 -13704 18634 -13604
rect 18634 -13704 18696 -13604
rect 8352 -19166 8452 -13994
rect 9492 -15009 9676 -14975
rect 9950 -15009 10134 -14975
rect 10408 -15009 10592 -14975
rect 10866 -15009 11050 -14975
rect 11324 -15009 11508 -14975
rect 11782 -15009 11966 -14975
rect 12240 -15009 12424 -14975
rect 12698 -15009 12882 -14975
rect 13156 -15009 13340 -14975
rect 13614 -15009 13798 -14975
rect 14072 -15009 14256 -14975
rect 14530 -15009 14714 -14975
rect 14988 -15009 15172 -14975
rect 15446 -15009 15630 -14975
rect 15904 -15009 16088 -14975
rect 16362 -15009 16546 -14975
rect 16820 -15009 17004 -14975
rect 17278 -15009 17462 -14975
rect 9338 -16644 9372 -15068
rect 9796 -16644 9830 -15068
rect 10254 -16644 10288 -15068
rect 10712 -16644 10746 -15068
rect 11170 -16644 11204 -15068
rect 11628 -16644 11662 -15068
rect 12086 -16644 12120 -15068
rect 12544 -16644 12578 -15068
rect 13002 -16644 13036 -15068
rect 13460 -16644 13494 -15068
rect 13918 -16644 13952 -15068
rect 14376 -16644 14410 -15068
rect 14834 -16644 14868 -15068
rect 15292 -16644 15326 -15068
rect 15750 -16644 15784 -15068
rect 16208 -16644 16242 -15068
rect 16666 -16644 16700 -15068
rect 17124 -16644 17158 -15068
rect 17582 -16644 17616 -15068
rect 9492 -16737 9676 -16703
rect 9950 -16737 10134 -16703
rect 10408 -16737 10592 -16703
rect 10866 -16737 11050 -16703
rect 11324 -16737 11508 -16703
rect 11782 -16737 11966 -16703
rect 12240 -16737 12424 -16703
rect 12698 -16737 12882 -16703
rect 13156 -16737 13340 -16703
rect 13614 -16737 13798 -16703
rect 14072 -16737 14256 -16703
rect 14530 -16737 14714 -16703
rect 14988 -16737 15172 -16703
rect 15446 -16737 15630 -16703
rect 15904 -16737 16088 -16703
rect 16362 -16737 16546 -16703
rect 16820 -16737 17004 -16703
rect 17278 -16737 17462 -16703
rect 13222 -16868 13270 -16820
rect 13676 -16874 13736 -16814
rect 8933 -17674 9117 -17640
rect 9391 -17674 9575 -17640
rect 9849 -17674 10033 -17640
rect 10307 -17674 10491 -17640
rect 10765 -17674 10949 -17640
rect 11223 -17674 11407 -17640
rect 11681 -17674 11865 -17640
rect 12139 -17674 12323 -17640
rect 12597 -17674 12781 -17640
rect 13055 -17674 13239 -17640
rect 13933 -17674 14117 -17640
rect 14391 -17674 14575 -17640
rect 14849 -17674 15033 -17640
rect 15307 -17674 15491 -17640
rect 15765 -17674 15949 -17640
rect 16223 -17674 16407 -17640
rect 16681 -17674 16865 -17640
rect 17139 -17674 17323 -17640
rect 17597 -17674 17781 -17640
rect 18055 -17674 18239 -17640
rect 8779 -18909 8813 -17733
rect 9237 -18909 9271 -17733
rect 9695 -18909 9729 -17733
rect 10153 -18909 10187 -17733
rect 10611 -18909 10645 -17733
rect 11069 -18909 11103 -17733
rect 11527 -18909 11561 -17733
rect 11985 -18909 12019 -17733
rect 12443 -18909 12477 -17733
rect 12901 -18909 12935 -17733
rect 13359 -18909 13393 -17733
rect 13779 -18909 13813 -17733
rect 14237 -18909 14271 -17733
rect 14695 -18909 14729 -17733
rect 15153 -18909 15187 -17733
rect 15611 -18909 15645 -17733
rect 16069 -18909 16103 -17733
rect 16527 -18909 16561 -17733
rect 16985 -18909 17019 -17733
rect 17443 -18909 17477 -17733
rect 17901 -18909 17935 -17733
rect 18359 -18909 18393 -17733
rect 8933 -19002 9117 -18968
rect 9391 -19002 9575 -18968
rect 9849 -19002 10033 -18968
rect 10307 -19002 10491 -18968
rect 10765 -19002 10949 -18968
rect 11223 -19002 11407 -18968
rect 11681 -19002 11865 -18968
rect 12139 -19002 12323 -18968
rect 12597 -19002 12781 -18968
rect 13055 -19002 13239 -18968
rect 13933 -19002 14117 -18968
rect 14391 -19002 14575 -18968
rect 14849 -19002 15033 -18968
rect 15307 -19002 15491 -18968
rect 15765 -19002 15949 -18968
rect 16223 -19002 16407 -18968
rect 16681 -19002 16865 -18968
rect 17139 -19002 17323 -18968
rect 17597 -19002 17781 -18968
rect 18055 -19002 18239 -18968
rect 18696 -19166 18796 -13994
rect 8452 -19448 8514 -19348
rect 8514 -19448 18634 -19348
rect 18634 -19448 18696 -19348
rect 23452 -13704 23514 -13604
rect 23514 -13704 33634 -13604
rect 33634 -13704 33696 -13604
rect 23352 -19166 23452 -13994
rect 24492 -15009 24676 -14975
rect 24950 -15009 25134 -14975
rect 25408 -15009 25592 -14975
rect 25866 -15009 26050 -14975
rect 26324 -15009 26508 -14975
rect 26782 -15009 26966 -14975
rect 27240 -15009 27424 -14975
rect 27698 -15009 27882 -14975
rect 28156 -15009 28340 -14975
rect 28614 -15009 28798 -14975
rect 29072 -15009 29256 -14975
rect 29530 -15009 29714 -14975
rect 29988 -15009 30172 -14975
rect 30446 -15009 30630 -14975
rect 30904 -15009 31088 -14975
rect 31362 -15009 31546 -14975
rect 31820 -15009 32004 -14975
rect 32278 -15009 32462 -14975
rect 24338 -16644 24372 -15068
rect 24796 -16644 24830 -15068
rect 25254 -16644 25288 -15068
rect 25712 -16644 25746 -15068
rect 26170 -16644 26204 -15068
rect 26628 -16644 26662 -15068
rect 27086 -16644 27120 -15068
rect 27544 -16644 27578 -15068
rect 28002 -16644 28036 -15068
rect 28460 -16644 28494 -15068
rect 28918 -16644 28952 -15068
rect 29376 -16644 29410 -15068
rect 29834 -16644 29868 -15068
rect 30292 -16644 30326 -15068
rect 30750 -16644 30784 -15068
rect 31208 -16644 31242 -15068
rect 31666 -16644 31700 -15068
rect 32124 -16644 32158 -15068
rect 32582 -16644 32616 -15068
rect 24492 -16737 24676 -16703
rect 24950 -16737 25134 -16703
rect 25408 -16737 25592 -16703
rect 25866 -16737 26050 -16703
rect 26324 -16737 26508 -16703
rect 26782 -16737 26966 -16703
rect 27240 -16737 27424 -16703
rect 27698 -16737 27882 -16703
rect 28156 -16737 28340 -16703
rect 28614 -16737 28798 -16703
rect 29072 -16737 29256 -16703
rect 29530 -16737 29714 -16703
rect 29988 -16737 30172 -16703
rect 30446 -16737 30630 -16703
rect 30904 -16737 31088 -16703
rect 31362 -16737 31546 -16703
rect 31820 -16737 32004 -16703
rect 32278 -16737 32462 -16703
rect 28222 -16868 28270 -16820
rect 28676 -16874 28736 -16814
rect 23933 -17674 24117 -17640
rect 24391 -17674 24575 -17640
rect 24849 -17674 25033 -17640
rect 25307 -17674 25491 -17640
rect 25765 -17674 25949 -17640
rect 26223 -17674 26407 -17640
rect 26681 -17674 26865 -17640
rect 27139 -17674 27323 -17640
rect 27597 -17674 27781 -17640
rect 28055 -17674 28239 -17640
rect 28933 -17674 29117 -17640
rect 29391 -17674 29575 -17640
rect 29849 -17674 30033 -17640
rect 30307 -17674 30491 -17640
rect 30765 -17674 30949 -17640
rect 31223 -17674 31407 -17640
rect 31681 -17674 31865 -17640
rect 32139 -17674 32323 -17640
rect 32597 -17674 32781 -17640
rect 33055 -17674 33239 -17640
rect 23779 -18909 23813 -17733
rect 24237 -18909 24271 -17733
rect 24695 -18909 24729 -17733
rect 25153 -18909 25187 -17733
rect 25611 -18909 25645 -17733
rect 26069 -18909 26103 -17733
rect 26527 -18909 26561 -17733
rect 26985 -18909 27019 -17733
rect 27443 -18909 27477 -17733
rect 27901 -18909 27935 -17733
rect 28359 -18909 28393 -17733
rect 28779 -18909 28813 -17733
rect 29237 -18909 29271 -17733
rect 29695 -18909 29729 -17733
rect 30153 -18909 30187 -17733
rect 30611 -18909 30645 -17733
rect 31069 -18909 31103 -17733
rect 31527 -18909 31561 -17733
rect 31985 -18909 32019 -17733
rect 32443 -18909 32477 -17733
rect 32901 -18909 32935 -17733
rect 33359 -18909 33393 -17733
rect 23933 -19002 24117 -18968
rect 24391 -19002 24575 -18968
rect 24849 -19002 25033 -18968
rect 25307 -19002 25491 -18968
rect 25765 -19002 25949 -18968
rect 26223 -19002 26407 -18968
rect 26681 -19002 26865 -18968
rect 27139 -19002 27323 -18968
rect 27597 -19002 27781 -18968
rect 28055 -19002 28239 -18968
rect 28933 -19002 29117 -18968
rect 29391 -19002 29575 -18968
rect 29849 -19002 30033 -18968
rect 30307 -19002 30491 -18968
rect 30765 -19002 30949 -18968
rect 31223 -19002 31407 -18968
rect 31681 -19002 31865 -18968
rect 32139 -19002 32323 -18968
rect 32597 -19002 32781 -18968
rect 33055 -19002 33239 -18968
rect 33696 -19166 33796 -13994
rect 23452 -19448 23514 -19348
rect 23514 -19448 33634 -19348
rect 33634 -19448 33696 -19348
rect 8452 -19784 8514 -19684
rect 8514 -19784 18634 -19684
rect 18634 -19784 18696 -19684
rect 8352 -21918 8452 -19914
rect 8932 -20176 9116 -20142
rect 9390 -20176 9574 -20142
rect 9848 -20176 10032 -20142
rect 10306 -20176 10490 -20142
rect 10764 -20176 10948 -20142
rect 11222 -20176 11406 -20142
rect 11680 -20176 11864 -20142
rect 12138 -20176 12322 -20142
rect 12596 -20176 12780 -20142
rect 13054 -20176 13238 -20142
rect 13932 -20176 14116 -20142
rect 14390 -20176 14574 -20142
rect 14848 -20176 15032 -20142
rect 15306 -20176 15490 -20142
rect 15764 -20176 15948 -20142
rect 16222 -20176 16406 -20142
rect 16680 -20176 16864 -20142
rect 17138 -20176 17322 -20142
rect 17596 -20176 17780 -20142
rect 18054 -20176 18238 -20142
rect 8778 -20402 8812 -20226
rect 9236 -20402 9270 -20226
rect 9694 -20402 9728 -20226
rect 10152 -20402 10186 -20226
rect 10610 -20402 10644 -20226
rect 11068 -20402 11102 -20226
rect 11526 -20402 11560 -20226
rect 11984 -20402 12018 -20226
rect 12442 -20402 12476 -20226
rect 12900 -20402 12934 -20226
rect 13358 -20402 13392 -20226
rect 13778 -20402 13812 -20226
rect 14236 -20402 14270 -20226
rect 14694 -20402 14728 -20226
rect 15152 -20402 15186 -20226
rect 15610 -20402 15644 -20226
rect 16068 -20402 16102 -20226
rect 16526 -20402 16560 -20226
rect 16984 -20402 17018 -20226
rect 17442 -20402 17476 -20226
rect 17900 -20402 17934 -20226
rect 18358 -20402 18392 -20226
rect 8932 -20486 9116 -20452
rect 9390 -20486 9574 -20452
rect 9848 -20486 10032 -20452
rect 10306 -20486 10490 -20452
rect 10764 -20486 10948 -20452
rect 11222 -20486 11406 -20452
rect 11680 -20486 11864 -20452
rect 12138 -20486 12322 -20452
rect 12596 -20486 12780 -20452
rect 13054 -20486 13238 -20452
rect 13932 -20486 14116 -20452
rect 14390 -20486 14574 -20452
rect 14848 -20486 15032 -20452
rect 15306 -20486 15490 -20452
rect 15764 -20486 15948 -20452
rect 16222 -20486 16406 -20452
rect 16680 -20486 16864 -20452
rect 17138 -20486 17322 -20452
rect 17596 -20486 17780 -20452
rect 18054 -20486 18238 -20452
rect 8932 -20844 9116 -20810
rect 9390 -20844 9574 -20810
rect 9848 -20844 10032 -20810
rect 10306 -20844 10490 -20810
rect 10764 -20844 10948 -20810
rect 11222 -20844 11406 -20810
rect 11680 -20844 11864 -20810
rect 12138 -20844 12322 -20810
rect 12596 -20844 12780 -20810
rect 13054 -20844 13238 -20810
rect 8778 -21070 8812 -20894
rect 9236 -21070 9270 -20894
rect 9694 -21070 9728 -20894
rect 10152 -21070 10186 -20894
rect 10610 -21070 10644 -20894
rect 11068 -21070 11102 -20894
rect 11526 -21070 11560 -20894
rect 11984 -21070 12018 -20894
rect 12442 -21070 12476 -20894
rect 12900 -21070 12934 -20894
rect 13358 -21070 13392 -20894
rect 8932 -21154 9116 -21120
rect 9390 -21154 9574 -21120
rect 9848 -21154 10032 -21120
rect 10306 -21154 10490 -21120
rect 10764 -21154 10948 -21120
rect 11222 -21154 11406 -21120
rect 11680 -21154 11864 -21120
rect 12138 -21154 12322 -21120
rect 12596 -21154 12780 -21120
rect 13054 -21154 13238 -21120
rect 18696 -21918 18796 -19914
rect 8452 -22148 8514 -22048
rect 8514 -22148 18634 -22048
rect 18634 -22148 18696 -22048
rect 23452 -19784 23514 -19684
rect 23514 -19784 33634 -19684
rect 33634 -19784 33696 -19684
rect 23352 -21918 23452 -19914
rect 23932 -20176 24116 -20142
rect 24390 -20176 24574 -20142
rect 24848 -20176 25032 -20142
rect 25306 -20176 25490 -20142
rect 25764 -20176 25948 -20142
rect 26222 -20176 26406 -20142
rect 26680 -20176 26864 -20142
rect 27138 -20176 27322 -20142
rect 27596 -20176 27780 -20142
rect 28054 -20176 28238 -20142
rect 28932 -20176 29116 -20142
rect 29390 -20176 29574 -20142
rect 29848 -20176 30032 -20142
rect 30306 -20176 30490 -20142
rect 30764 -20176 30948 -20142
rect 31222 -20176 31406 -20142
rect 31680 -20176 31864 -20142
rect 32138 -20176 32322 -20142
rect 32596 -20176 32780 -20142
rect 33054 -20176 33238 -20142
rect 23778 -20402 23812 -20226
rect 24236 -20402 24270 -20226
rect 24694 -20402 24728 -20226
rect 25152 -20402 25186 -20226
rect 25610 -20402 25644 -20226
rect 26068 -20402 26102 -20226
rect 26526 -20402 26560 -20226
rect 26984 -20402 27018 -20226
rect 27442 -20402 27476 -20226
rect 27900 -20402 27934 -20226
rect 28358 -20402 28392 -20226
rect 28778 -20402 28812 -20226
rect 29236 -20402 29270 -20226
rect 29694 -20402 29728 -20226
rect 30152 -20402 30186 -20226
rect 30610 -20402 30644 -20226
rect 31068 -20402 31102 -20226
rect 31526 -20402 31560 -20226
rect 31984 -20402 32018 -20226
rect 32442 -20402 32476 -20226
rect 32900 -20402 32934 -20226
rect 33358 -20402 33392 -20226
rect 23932 -20486 24116 -20452
rect 24390 -20486 24574 -20452
rect 24848 -20486 25032 -20452
rect 25306 -20486 25490 -20452
rect 25764 -20486 25948 -20452
rect 26222 -20486 26406 -20452
rect 26680 -20486 26864 -20452
rect 27138 -20486 27322 -20452
rect 27596 -20486 27780 -20452
rect 28054 -20486 28238 -20452
rect 28932 -20486 29116 -20452
rect 29390 -20486 29574 -20452
rect 29848 -20486 30032 -20452
rect 30306 -20486 30490 -20452
rect 30764 -20486 30948 -20452
rect 31222 -20486 31406 -20452
rect 31680 -20486 31864 -20452
rect 32138 -20486 32322 -20452
rect 32596 -20486 32780 -20452
rect 33054 -20486 33238 -20452
rect 23932 -20844 24116 -20810
rect 24390 -20844 24574 -20810
rect 24848 -20844 25032 -20810
rect 25306 -20844 25490 -20810
rect 25764 -20844 25948 -20810
rect 26222 -20844 26406 -20810
rect 26680 -20844 26864 -20810
rect 27138 -20844 27322 -20810
rect 27596 -20844 27780 -20810
rect 28054 -20844 28238 -20810
rect 23778 -21070 23812 -20894
rect 24236 -21070 24270 -20894
rect 24694 -21070 24728 -20894
rect 25152 -21070 25186 -20894
rect 25610 -21070 25644 -20894
rect 26068 -21070 26102 -20894
rect 26526 -21070 26560 -20894
rect 26984 -21070 27018 -20894
rect 27442 -21070 27476 -20894
rect 27900 -21070 27934 -20894
rect 28358 -21070 28392 -20894
rect 23932 -21154 24116 -21120
rect 24390 -21154 24574 -21120
rect 24848 -21154 25032 -21120
rect 25306 -21154 25490 -21120
rect 25764 -21154 25948 -21120
rect 26222 -21154 26406 -21120
rect 26680 -21154 26864 -21120
rect 27138 -21154 27322 -21120
rect 27596 -21154 27780 -21120
rect 28054 -21154 28238 -21120
rect 33696 -21918 33796 -19914
rect 23452 -22148 23514 -22048
rect 23514 -22148 33634 -22048
rect 33634 -22148 33696 -22048
<< metal1 >>
rect 23328 17500 32784 17506
rect 23328 17400 23434 17500
rect 32678 17400 32784 17500
rect 23328 17394 32784 17400
rect 23328 17295 23440 17394
rect 23328 15401 23334 17295
rect 23434 15401 23440 17295
rect 24040 17094 24050 17394
rect 32062 17094 32072 17394
rect 32672 17295 32784 17394
rect 23526 16978 32596 17012
rect 23526 16868 23562 16978
rect 32558 16868 32596 16978
rect 23526 16830 32596 16868
rect 23596 16606 23602 16666
rect 23662 16606 23668 16666
rect 23764 16658 23824 16830
rect 24196 16658 24256 16830
rect 25480 16670 25540 16830
rect 27194 16670 27254 16830
rect 23602 15474 23662 16606
rect 23764 16598 24256 16658
rect 24616 16606 24622 16666
rect 24682 16606 24688 16666
rect 25480 16610 27254 16670
rect 28910 16666 28970 16830
rect 30628 16666 30688 16830
rect 23764 16422 23824 16598
rect 24196 16521 24256 16598
rect 24018 16515 24426 16521
rect 24018 16481 24030 16515
rect 24414 16481 24426 16515
rect 24018 16475 24426 16481
rect 23764 16246 23776 16422
rect 23810 16246 23824 16422
rect 24622 16422 24682 16606
rect 24876 16515 25284 16521
rect 24876 16481 24888 16515
rect 25272 16481 25284 16515
rect 24876 16475 25284 16481
rect 24622 16392 24634 16422
rect 23764 16064 23824 16246
rect 24628 16246 24634 16392
rect 24668 16392 24682 16422
rect 25480 16422 25540 16610
rect 25734 16515 26142 16521
rect 25734 16481 25746 16515
rect 26130 16481 26142 16515
rect 25734 16475 26142 16481
rect 26592 16515 27000 16521
rect 26592 16481 26604 16515
rect 26988 16481 27000 16515
rect 26592 16475 27000 16481
rect 24668 16246 24674 16392
rect 24628 16234 24674 16246
rect 25480 16246 25492 16422
rect 25526 16246 25540 16422
rect 26344 16422 26390 16434
rect 26344 16308 26350 16422
rect 24018 16187 24426 16193
rect 24018 16153 24030 16187
rect 24414 16153 24426 16187
rect 24018 16147 24426 16153
rect 24876 16187 25284 16193
rect 24876 16153 24888 16187
rect 25272 16153 25284 16187
rect 24876 16147 25284 16153
rect 24196 16064 24256 16147
rect 25060 16066 25120 16147
rect 23764 16004 24256 16064
rect 24614 16006 24620 16066
rect 24680 16006 24686 16066
rect 25054 16006 25060 16066
rect 25120 16006 25126 16066
rect 23764 15822 23824 16004
rect 24196 15921 24256 16004
rect 24018 15915 24426 15921
rect 24018 15881 24030 15915
rect 24414 15881 24426 15915
rect 24018 15875 24426 15881
rect 23764 15646 23776 15822
rect 23810 15646 23824 15822
rect 24620 15822 24680 16006
rect 25060 15921 25120 16006
rect 24876 15915 25284 15921
rect 24876 15881 24888 15915
rect 25272 15881 25284 15915
rect 24876 15875 25284 15881
rect 24620 15776 24634 15822
rect 23764 15482 23824 15646
rect 24628 15646 24634 15776
rect 24668 15776 24680 15822
rect 25480 15822 25540 16246
rect 26336 16246 26350 16308
rect 26384 16308 26390 16422
rect 27194 16422 27254 16610
rect 28050 16606 28056 16666
rect 28116 16606 28122 16666
rect 28910 16606 30688 16666
rect 31480 16612 31486 16672
rect 31546 16612 31552 16672
rect 31920 16644 31980 16830
rect 32342 16644 32402 16830
rect 27450 16515 27858 16521
rect 27450 16481 27462 16515
rect 27846 16481 27858 16515
rect 27450 16475 27858 16481
rect 26384 16246 26396 16308
rect 25734 16187 26142 16193
rect 25734 16153 25746 16187
rect 26130 16153 26142 16187
rect 25734 16147 26142 16153
rect 25900 16066 25960 16147
rect 26336 16066 26396 16246
rect 27194 16246 27208 16422
rect 27242 16246 27254 16422
rect 28056 16422 28116 16606
rect 28308 16515 28716 16521
rect 28308 16481 28320 16515
rect 28704 16481 28716 16515
rect 28308 16475 28716 16481
rect 28056 16368 28066 16422
rect 26592 16187 27000 16193
rect 26592 16153 26604 16187
rect 26988 16153 27000 16187
rect 26592 16147 27000 16153
rect 26770 16066 26830 16147
rect 25894 16006 25900 16066
rect 25960 16006 25966 16066
rect 26330 16006 26336 16066
rect 26396 16006 26402 16066
rect 26764 16006 26770 16066
rect 26830 16006 26836 16066
rect 25900 15921 25960 16006
rect 26770 15921 26830 16006
rect 25734 15915 26142 15921
rect 25734 15881 25746 15915
rect 26130 15881 26142 15915
rect 25734 15875 26142 15881
rect 26592 15915 27000 15921
rect 26592 15881 26604 15915
rect 26988 15881 27000 15915
rect 26592 15875 27000 15881
rect 25480 15778 25492 15822
rect 24668 15646 24674 15776
rect 24628 15634 24674 15646
rect 25486 15646 25492 15778
rect 25526 15778 25540 15822
rect 26344 15822 26390 15834
rect 25526 15646 25532 15778
rect 26344 15696 26350 15822
rect 25486 15634 25532 15646
rect 26340 15646 26350 15696
rect 26384 15696 26390 15822
rect 27194 15822 27254 16246
rect 28060 16246 28066 16368
rect 28100 16368 28116 16422
rect 28910 16422 28970 16606
rect 29166 16515 29574 16521
rect 29166 16481 29178 16515
rect 29562 16481 29574 16515
rect 29166 16475 29574 16481
rect 30024 16515 30432 16521
rect 30024 16481 30036 16515
rect 30420 16481 30432 16515
rect 30024 16475 30432 16481
rect 28100 16246 28106 16368
rect 28060 16234 28106 16246
rect 28910 16246 28924 16422
rect 28958 16246 28970 16422
rect 29776 16422 29822 16434
rect 29776 16308 29782 16422
rect 27450 16187 27858 16193
rect 27450 16153 27462 16187
rect 27846 16153 27858 16187
rect 27450 16147 27858 16153
rect 28308 16187 28716 16193
rect 28308 16153 28320 16187
rect 28704 16153 28716 16187
rect 28308 16147 28716 16153
rect 27632 16066 27692 16147
rect 28484 16066 28544 16147
rect 27626 16006 27632 16066
rect 27692 16006 27698 16066
rect 28046 16006 28052 16066
rect 28112 16006 28118 16066
rect 28478 16006 28484 16066
rect 28544 16006 28550 16066
rect 27632 15921 27692 16006
rect 27450 15915 27858 15921
rect 27450 15881 27462 15915
rect 27846 15881 27858 15915
rect 27450 15875 27858 15881
rect 27194 15772 27208 15822
rect 26384 15646 26400 15696
rect 24018 15587 24426 15593
rect 24018 15553 24030 15587
rect 24414 15553 24426 15587
rect 24018 15547 24426 15553
rect 24876 15587 25284 15593
rect 24876 15553 24888 15587
rect 25272 15553 25284 15587
rect 24876 15547 25284 15553
rect 25734 15587 26142 15593
rect 25734 15553 25746 15587
rect 26130 15553 26142 15587
rect 25734 15547 26142 15553
rect 24200 15482 24260 15547
rect 23596 15414 23602 15474
rect 23662 15414 23668 15474
rect 23762 15422 24260 15482
rect 26340 15474 26400 15646
rect 27202 15646 27208 15772
rect 27242 15772 27254 15822
rect 28052 15822 28112 16006
rect 28484 15921 28544 16006
rect 28308 15915 28716 15921
rect 28308 15881 28320 15915
rect 28704 15881 28716 15915
rect 28308 15875 28716 15881
rect 28052 15776 28066 15822
rect 27242 15646 27248 15772
rect 27202 15634 27248 15646
rect 28060 15646 28066 15776
rect 28100 15776 28112 15822
rect 28910 15822 28970 16246
rect 29770 16246 29782 16308
rect 29816 16308 29822 16422
rect 30628 16422 30688 16606
rect 30882 16515 31290 16521
rect 30882 16481 30894 16515
rect 31278 16481 31290 16515
rect 30882 16475 31290 16481
rect 29816 16246 29830 16308
rect 29166 16187 29574 16193
rect 29166 16153 29178 16187
rect 29562 16153 29574 16187
rect 29166 16147 29574 16153
rect 29340 16066 29400 16147
rect 29770 16066 29830 16246
rect 30628 16246 30640 16422
rect 30674 16246 30688 16422
rect 31486 16422 31546 16612
rect 31920 16584 32402 16644
rect 32488 16612 32494 16672
rect 32554 16612 32560 16672
rect 31920 16521 31980 16584
rect 31740 16515 32148 16521
rect 31740 16481 31752 16515
rect 32136 16481 32148 16515
rect 31740 16475 32148 16481
rect 31486 16374 31498 16422
rect 30024 16187 30432 16193
rect 30024 16153 30036 16187
rect 30420 16153 30432 16187
rect 30024 16147 30432 16153
rect 30202 16066 30262 16147
rect 29334 16006 29340 16066
rect 29400 16006 29406 16066
rect 29764 16006 29770 16066
rect 29830 16006 29836 16066
rect 30196 16006 30202 16066
rect 30262 16006 30268 16066
rect 29340 15921 29400 16006
rect 30202 15921 30262 16006
rect 29166 15915 29574 15921
rect 29166 15881 29178 15915
rect 29562 15881 29574 15915
rect 29166 15875 29574 15881
rect 30024 15915 30432 15921
rect 30024 15881 30036 15915
rect 30420 15881 30432 15915
rect 30024 15875 30432 15881
rect 28100 15646 28106 15776
rect 28910 15768 28924 15822
rect 28060 15634 28106 15646
rect 28918 15646 28924 15768
rect 28958 15768 28970 15822
rect 29776 15822 29822 15834
rect 28958 15646 28964 15768
rect 29776 15692 29782 15822
rect 28918 15634 28964 15646
rect 29770 15646 29782 15692
rect 29816 15692 29822 15822
rect 30628 15822 30688 16246
rect 31492 16246 31498 16374
rect 31532 16374 31546 16422
rect 32342 16422 32402 16584
rect 31532 16246 31538 16374
rect 31492 16234 31538 16246
rect 32342 16246 32356 16422
rect 32390 16246 32402 16422
rect 30882 16187 31290 16193
rect 30882 16153 30894 16187
rect 31278 16153 31290 16187
rect 30882 16147 31290 16153
rect 31740 16187 32148 16193
rect 31740 16153 31752 16187
rect 32136 16153 32148 16187
rect 31740 16147 32148 16153
rect 31052 16066 31112 16147
rect 31918 16066 31978 16147
rect 32342 16066 32402 16246
rect 31046 16006 31052 16066
rect 31112 16006 31118 16066
rect 31480 16006 31486 16066
rect 31546 16006 31552 16066
rect 31918 16006 32402 16066
rect 31052 15921 31112 16006
rect 30882 15915 31290 15921
rect 30882 15881 30894 15915
rect 31278 15881 31290 15915
rect 30882 15875 31290 15881
rect 30628 15784 30640 15822
rect 29816 15646 29830 15692
rect 26592 15587 27000 15593
rect 26592 15553 26604 15587
rect 26988 15553 27000 15587
rect 26592 15547 27000 15553
rect 27450 15587 27858 15593
rect 27450 15553 27462 15587
rect 27846 15553 27858 15587
rect 27450 15547 27858 15553
rect 28308 15587 28716 15593
rect 28308 15553 28320 15587
rect 28704 15553 28716 15587
rect 28308 15547 28716 15553
rect 29166 15587 29574 15593
rect 29166 15553 29178 15587
rect 29562 15553 29574 15587
rect 29166 15547 29574 15553
rect 29770 15474 29830 15646
rect 30634 15646 30640 15784
rect 30674 15784 30688 15822
rect 31486 15822 31546 16006
rect 31918 15921 31978 16006
rect 31740 15915 32148 15921
rect 31740 15881 31752 15915
rect 32136 15881 32148 15915
rect 31740 15875 32148 15881
rect 30674 15646 30680 15784
rect 31486 15780 31498 15822
rect 30634 15634 30680 15646
rect 31492 15646 31498 15780
rect 31532 15780 31546 15822
rect 32342 15822 32402 16006
rect 31532 15646 31538 15780
rect 31492 15634 31538 15646
rect 32342 15646 32356 15822
rect 32390 15646 32402 15822
rect 30024 15587 30432 15593
rect 30024 15553 30036 15587
rect 30420 15553 30432 15587
rect 30024 15547 30432 15553
rect 30882 15587 31290 15593
rect 30882 15553 30894 15587
rect 31278 15553 31290 15587
rect 30882 15547 31290 15553
rect 31740 15587 32148 15593
rect 31740 15553 31752 15587
rect 32136 15553 32148 15587
rect 31740 15547 32148 15553
rect 31922 15486 31982 15547
rect 32342 15486 32402 15646
rect 23328 15302 23440 15401
rect 23764 15302 23824 15422
rect 24200 15302 24260 15422
rect 26334 15414 26340 15474
rect 26400 15414 26406 15474
rect 29764 15414 29770 15474
rect 29830 15414 29836 15474
rect 31922 15426 32402 15486
rect 32494 15474 32554 16612
rect 31922 15302 31982 15426
rect 32342 15302 32402 15426
rect 32488 15414 32494 15474
rect 32554 15414 32560 15474
rect 32672 15401 32678 17295
rect 32778 15401 32784 17295
rect 32672 15302 32784 15401
rect 23328 15296 32784 15302
rect 23328 15196 23434 15296
rect 32678 15196 32784 15296
rect 23328 15190 32784 15196
rect 24034 15002 24098 15190
rect 24152 15002 24212 15190
rect 24276 15002 24336 15190
rect 24528 15078 24534 15138
rect 24594 15078 24600 15138
rect 24034 14942 24336 15002
rect 24034 14882 24098 14942
rect 24034 14308 24048 14882
rect 24084 14308 24098 14882
rect 24152 14782 24212 14942
rect 24276 14881 24336 14942
rect 24534 14881 24594 15078
rect 24792 14997 24852 15190
rect 24922 14997 24982 15190
rect 25032 14997 25222 15190
rect 24658 14934 24664 14994
rect 24724 14934 24730 14994
rect 24792 14937 25222 14997
rect 24255 14875 24363 14881
rect 24255 14841 24267 14875
rect 24351 14841 24363 14875
rect 24255 14835 24363 14841
rect 24513 14875 24621 14881
rect 24513 14841 24525 14875
rect 24609 14841 24621 14875
rect 24513 14835 24621 14841
rect 24152 14754 24163 14782
rect 24157 14406 24163 14754
rect 24197 14754 24212 14782
rect 24415 14782 24461 14794
rect 24197 14406 24203 14754
rect 24415 14432 24421 14782
rect 24157 14394 24203 14406
rect 24408 14406 24421 14432
rect 24455 14432 24461 14782
rect 24664 14782 24724 14934
rect 24792 14881 24852 14937
rect 24771 14875 24879 14881
rect 24771 14841 24783 14875
rect 24867 14841 24879 14875
rect 24771 14835 24879 14841
rect 24664 14746 24679 14782
rect 24455 14406 24468 14432
rect 24034 14296 24098 14308
rect 24255 14347 24363 14353
rect 24255 14313 24267 14347
rect 24351 14313 24363 14347
rect 24255 14307 24363 14313
rect 23080 14160 23140 14166
rect 24408 14160 24468 14406
rect 24673 14406 24679 14746
rect 24713 14746 24724 14782
rect 24922 14782 24982 14937
rect 24713 14406 24719 14746
rect 24922 14740 24937 14782
rect 24673 14394 24719 14406
rect 24931 14406 24937 14740
rect 24971 14740 24982 14782
rect 25032 14882 25222 14937
rect 24971 14406 24977 14740
rect 24931 14394 24977 14406
rect 24513 14347 24621 14353
rect 24513 14313 24525 14347
rect 24609 14313 24621 14347
rect 24513 14307 24621 14313
rect 24771 14347 24879 14353
rect 24771 14313 24783 14347
rect 24867 14313 24879 14347
rect 24771 14307 24879 14313
rect 25032 14308 25050 14882
rect 25086 14308 25170 14882
rect 25206 14308 25222 14882
rect 25268 15002 25328 15190
rect 25398 15002 25458 15190
rect 25268 14942 25458 15002
rect 25268 14782 25328 14942
rect 25398 14881 25458 14942
rect 25522 14934 25528 14994
rect 25588 14934 25594 14994
rect 25650 14936 25656 14996
rect 25716 14936 25722 14996
rect 25916 14994 25976 15190
rect 26044 14994 26104 15190
rect 26174 14994 26234 15190
rect 25377 14875 25485 14881
rect 25377 14841 25389 14875
rect 25473 14841 25485 14875
rect 25377 14835 25485 14841
rect 25268 14731 25285 14782
rect 25279 14406 25285 14731
rect 25319 14731 25328 14782
rect 25528 14782 25588 14934
rect 25656 14881 25716 14936
rect 25916 14934 26234 14994
rect 25916 14881 25976 14934
rect 25635 14875 25743 14881
rect 25635 14841 25647 14875
rect 25731 14841 25743 14875
rect 25635 14835 25743 14841
rect 25893 14875 26001 14881
rect 25893 14841 25905 14875
rect 25989 14841 26001 14875
rect 25893 14835 26001 14841
rect 25528 14742 25543 14782
rect 25319 14406 25325 14731
rect 25279 14394 25325 14406
rect 25537 14406 25543 14742
rect 25577 14742 25588 14782
rect 25795 14782 25841 14794
rect 25577 14406 25583 14742
rect 25795 14440 25801 14782
rect 25537 14394 25583 14406
rect 25786 14406 25801 14440
rect 25835 14440 25841 14782
rect 26044 14782 26104 14934
rect 26174 14881 26234 14934
rect 26562 14994 26622 15190
rect 26686 14994 26746 15190
rect 26820 14994 26880 15190
rect 26932 14994 26996 15190
rect 26562 14934 26996 14994
rect 26151 14875 26259 14881
rect 26151 14841 26163 14875
rect 26247 14841 26259 14875
rect 26151 14835 26259 14841
rect 26409 14875 26517 14881
rect 26409 14841 26421 14875
rect 26505 14841 26517 14875
rect 26409 14835 26517 14841
rect 26044 14754 26059 14782
rect 25835 14406 25846 14440
rect 25032 14294 25222 14308
rect 25377 14347 25485 14353
rect 25377 14313 25389 14347
rect 25473 14313 25485 14347
rect 25377 14307 25485 14313
rect 25635 14347 25743 14353
rect 25635 14313 25647 14347
rect 25731 14313 25743 14347
rect 25635 14307 25743 14313
rect 23140 14100 24468 14160
rect 23080 14094 23140 14100
rect 24030 13986 24098 14004
rect 24030 13630 24048 13986
rect 24082 13630 24098 13986
rect 24255 13979 24363 13985
rect 24255 13945 24267 13979
rect 24351 13945 24363 13979
rect 24255 13939 24363 13945
rect 24157 13895 24203 13907
rect 24157 13744 24163 13895
rect 24030 13562 24098 13630
rect 24148 13719 24163 13744
rect 24197 13744 24203 13895
rect 24408 13895 24468 14100
rect 25786 14094 25846 14406
rect 26053 14406 26059 14754
rect 26093 14754 26104 14782
rect 26311 14782 26357 14794
rect 26093 14406 26099 14754
rect 26311 14454 26317 14782
rect 26053 14394 26099 14406
rect 26304 14406 26317 14454
rect 26351 14454 26357 14782
rect 26562 14782 26622 14934
rect 26686 14881 26746 14934
rect 26667 14875 26775 14881
rect 26667 14841 26679 14875
rect 26763 14841 26775 14875
rect 26667 14835 26775 14841
rect 26562 14744 26575 14782
rect 26351 14406 26364 14454
rect 25893 14347 26001 14353
rect 25893 14313 25905 14347
rect 25989 14313 26001 14347
rect 25893 14307 26001 14313
rect 26151 14347 26259 14353
rect 26151 14313 26163 14347
rect 26247 14313 26259 14347
rect 26151 14307 26259 14313
rect 26304 14264 26364 14406
rect 26569 14406 26575 14744
rect 26609 14744 26622 14782
rect 26820 14782 26880 14934
rect 26820 14766 26833 14782
rect 26609 14406 26615 14744
rect 26569 14394 26615 14406
rect 26827 14406 26833 14766
rect 26867 14766 26880 14782
rect 26932 14884 26996 14934
rect 26867 14406 26873 14766
rect 26827 14394 26873 14406
rect 26409 14347 26517 14353
rect 26409 14313 26421 14347
rect 26505 14313 26517 14347
rect 26409 14307 26517 14313
rect 26667 14347 26775 14353
rect 26667 14313 26679 14347
rect 26763 14313 26775 14347
rect 26667 14307 26775 14313
rect 26932 14308 26948 14884
rect 26982 14308 26996 14884
rect 27262 14506 27506 15190
rect 28078 14506 28322 15190
rect 29078 14506 29322 15190
rect 30078 14506 30322 15190
rect 31078 14506 31322 15190
rect 32078 14506 32322 15190
rect 27260 14475 32322 14506
rect 27260 14441 27289 14475
rect 27323 14441 27381 14475
rect 27415 14441 27473 14475
rect 27507 14441 27565 14475
rect 27599 14441 27657 14475
rect 27691 14441 27749 14475
rect 27783 14441 27841 14475
rect 27875 14441 27933 14475
rect 27967 14441 28025 14475
rect 28059 14441 28117 14475
rect 28151 14441 28209 14475
rect 28243 14441 28301 14475
rect 28335 14441 28393 14475
rect 28427 14441 28485 14475
rect 28519 14441 28577 14475
rect 28611 14441 28669 14475
rect 28703 14441 28761 14475
rect 28795 14441 28853 14475
rect 28887 14441 28945 14475
rect 28979 14441 29037 14475
rect 29071 14441 29129 14475
rect 29163 14441 29221 14475
rect 29255 14441 29313 14475
rect 29347 14441 29405 14475
rect 29439 14441 29497 14475
rect 29531 14441 29589 14475
rect 29623 14441 29681 14475
rect 29715 14441 29773 14475
rect 29807 14441 29865 14475
rect 29899 14441 29957 14475
rect 29991 14441 30049 14475
rect 30083 14441 30141 14475
rect 30175 14441 30233 14475
rect 30267 14441 30325 14475
rect 30359 14441 30417 14475
rect 30451 14441 30509 14475
rect 30543 14441 30601 14475
rect 30635 14441 30693 14475
rect 30727 14441 30785 14475
rect 30819 14441 30877 14475
rect 30911 14441 30969 14475
rect 31003 14441 31061 14475
rect 31095 14441 31153 14475
rect 31187 14441 31245 14475
rect 31279 14441 31337 14475
rect 31371 14441 31429 14475
rect 31463 14441 31521 14475
rect 31555 14441 31613 14475
rect 31647 14441 31705 14475
rect 31739 14441 31797 14475
rect 31831 14441 31889 14475
rect 31923 14441 31981 14475
rect 32015 14441 32073 14475
rect 32107 14441 32165 14475
rect 32199 14441 32257 14475
rect 32291 14441 32322 14475
rect 27260 14410 32322 14441
rect 27530 14388 27596 14410
rect 27530 14348 27542 14388
rect 27582 14348 27596 14388
rect 31984 14396 32050 14410
rect 29994 14374 30054 14380
rect 27530 14336 27596 14348
rect 29988 14314 29994 14374
rect 30054 14314 30060 14374
rect 31984 14356 31992 14396
rect 32038 14356 32050 14396
rect 31984 14342 32050 14356
rect 26432 14264 26492 14307
rect 26932 14298 26996 14308
rect 27451 14305 27509 14311
rect 27451 14271 27463 14305
rect 27497 14302 27509 14305
rect 27829 14305 27887 14311
rect 27829 14302 27841 14305
rect 27497 14274 27841 14302
rect 27497 14271 27509 14274
rect 27451 14265 27509 14271
rect 27829 14271 27841 14274
rect 27875 14302 27887 14305
rect 28453 14305 28511 14311
rect 29994 14308 30054 14314
rect 28453 14302 28465 14305
rect 27875 14274 28465 14302
rect 27875 14271 27887 14274
rect 27829 14265 27887 14271
rect 28453 14271 28465 14274
rect 28499 14271 28511 14305
rect 31069 14305 31127 14311
rect 28453 14265 28511 14271
rect 28670 14268 30916 14274
rect 26304 14204 26624 14264
rect 25658 14034 25846 14094
rect 24513 13979 24621 13985
rect 24513 13945 24525 13979
rect 24609 13945 24621 13979
rect 24513 13939 24621 13945
rect 24771 13979 24879 13985
rect 24771 13945 24783 13979
rect 24867 13945 24879 13979
rect 24771 13939 24879 13945
rect 25030 13984 25224 14006
rect 25658 13985 25718 14034
rect 24408 13868 24421 13895
rect 24197 13719 24208 13744
rect 24148 13562 24208 13719
rect 24415 13719 24421 13868
rect 24455 13868 24468 13895
rect 24673 13895 24719 13907
rect 24455 13719 24461 13868
rect 24673 13750 24679 13895
rect 24415 13707 24461 13719
rect 24666 13719 24679 13750
rect 24713 13750 24719 13895
rect 24931 13895 24977 13907
rect 24931 13756 24937 13895
rect 24713 13719 24726 13750
rect 24255 13669 24363 13675
rect 24255 13635 24267 13669
rect 24351 13635 24363 13669
rect 24255 13629 24363 13635
rect 24513 13669 24621 13675
rect 24513 13635 24525 13669
rect 24609 13635 24621 13669
rect 24666 13656 24726 13719
rect 24922 13719 24937 13756
rect 24971 13756 24977 13895
rect 24971 13719 24982 13756
rect 24513 13629 24621 13635
rect 24280 13562 24340 13629
rect 24530 13564 24590 13629
rect 24664 13590 24726 13656
rect 24771 13669 24879 13675
rect 24771 13635 24783 13669
rect 24867 13635 24879 13669
rect 24771 13629 24879 13635
rect 24030 13502 24340 13562
rect 24524 13504 24530 13564
rect 24590 13504 24596 13564
rect 24030 13326 24098 13502
rect 24148 13326 24208 13502
rect 24280 13326 24340 13502
rect 24664 13446 24724 13590
rect 24794 13568 24854 13629
rect 24922 13568 24982 13719
rect 25030 13630 25050 13984
rect 25084 13630 25170 13984
rect 25204 13630 25224 13984
rect 25377 13979 25485 13985
rect 25377 13945 25389 13979
rect 25473 13945 25485 13979
rect 25377 13939 25485 13945
rect 25635 13979 25743 13985
rect 25635 13945 25647 13979
rect 25731 13945 25743 13979
rect 25635 13939 25743 13945
rect 25279 13895 25325 13907
rect 25279 13758 25285 13895
rect 25030 13568 25224 13630
rect 24794 13566 25224 13568
rect 25274 13719 25285 13758
rect 25319 13758 25325 13895
rect 25537 13895 25583 13907
rect 25537 13758 25543 13895
rect 25319 13719 25334 13758
rect 25274 13566 25334 13719
rect 25530 13719 25543 13758
rect 25577 13758 25583 13895
rect 25786 13895 25846 14034
rect 25893 13979 26001 13985
rect 25893 13945 25905 13979
rect 25989 13945 26001 13979
rect 25893 13939 26001 13945
rect 26151 13979 26259 13985
rect 26151 13945 26163 13979
rect 26247 13945 26259 13979
rect 26151 13939 26259 13945
rect 26409 13979 26517 13985
rect 26409 13945 26421 13979
rect 26505 13945 26517 13979
rect 26409 13939 26517 13945
rect 25786 13856 25801 13895
rect 25577 13719 25590 13758
rect 25377 13669 25485 13675
rect 25377 13635 25389 13669
rect 25473 13635 25485 13669
rect 25377 13629 25485 13635
rect 25402 13566 25462 13629
rect 25530 13566 25590 13719
rect 25795 13719 25801 13856
rect 25835 13856 25846 13895
rect 26053 13895 26099 13907
rect 25835 13719 25841 13856
rect 26053 13756 26059 13895
rect 25795 13707 25841 13719
rect 26046 13719 26059 13756
rect 26093 13756 26099 13895
rect 26311 13895 26357 13907
rect 26093 13719 26106 13756
rect 26311 13752 26317 13895
rect 25635 13669 25743 13675
rect 25635 13635 25647 13669
rect 25731 13635 25743 13669
rect 25635 13629 25743 13635
rect 25893 13669 26001 13675
rect 25893 13635 25905 13669
rect 25989 13635 26001 13669
rect 25893 13629 26001 13635
rect 24794 13508 25590 13566
rect 24664 13380 24724 13386
rect 25030 13506 25590 13508
rect 25916 13578 25976 13629
rect 26046 13578 26106 13719
rect 26304 13719 26317 13752
rect 26351 13752 26357 13895
rect 26564 13895 26624 14204
rect 28670 14226 29764 14268
rect 29812 14226 30916 14268
rect 31069 14271 31081 14305
rect 31115 14302 31127 14305
rect 31693 14305 31751 14311
rect 31693 14302 31705 14305
rect 31115 14274 31705 14302
rect 31115 14271 31127 14274
rect 31069 14265 31127 14271
rect 31693 14271 31705 14274
rect 31739 14302 31751 14305
rect 32071 14305 32129 14311
rect 32071 14302 32083 14305
rect 31739 14274 32083 14302
rect 31739 14271 31751 14274
rect 31693 14265 31751 14271
rect 32071 14271 32083 14274
rect 32117 14271 32129 14305
rect 32071 14265 32129 14271
rect 28670 14214 30916 14226
rect 27146 14096 27152 14196
rect 27252 14190 27334 14196
rect 27252 14142 27274 14190
rect 27322 14142 27334 14190
rect 27252 14136 27334 14142
rect 27370 14169 27428 14175
rect 27252 14096 27258 14136
rect 27370 14135 27382 14169
rect 27416 14166 27428 14169
rect 27737 14169 27795 14175
rect 27737 14166 27749 14169
rect 27416 14138 27749 14166
rect 27416 14135 27428 14138
rect 27370 14129 27428 14135
rect 27737 14135 27749 14138
rect 27783 14166 27795 14169
rect 28453 14169 28511 14175
rect 28670 14170 28730 14214
rect 29760 14212 29820 14214
rect 29356 14176 29416 14182
rect 29848 14176 29908 14182
rect 28453 14166 28465 14169
rect 27783 14138 28465 14166
rect 27783 14135 27795 14138
rect 27737 14129 27795 14135
rect 28453 14135 28465 14138
rect 28499 14135 28511 14169
rect 28453 14129 28511 14135
rect 28669 14164 28730 14170
rect 28669 14130 28681 14164
rect 28715 14130 28730 14164
rect 28669 14107 28730 14130
rect 28992 14170 29356 14176
rect 28992 14122 29004 14170
rect 29052 14122 29356 14170
rect 28992 14116 29356 14122
rect 29416 14170 29742 14176
rect 29416 14130 29444 14170
rect 29492 14130 29682 14170
rect 29416 14128 29682 14130
rect 29730 14128 29742 14170
rect 29416 14116 29742 14128
rect 29844 14116 29848 14176
rect 29908 14170 30588 14176
rect 30856 14170 30916 14214
rect 29908 14130 30090 14170
rect 30138 14130 30528 14170
rect 29908 14122 30528 14130
rect 30576 14122 30588 14170
rect 29908 14116 30588 14122
rect 30853 14164 30916 14170
rect 30853 14130 30865 14164
rect 30899 14130 30916 14164
rect 29356 14110 29416 14116
rect 29848 14110 29908 14116
rect 30853 14107 30916 14130
rect 31069 14169 31127 14175
rect 31069 14135 31081 14169
rect 31115 14166 31127 14169
rect 31785 14169 31843 14175
rect 31785 14166 31797 14169
rect 31115 14138 31797 14166
rect 31115 14135 31127 14138
rect 31069 14129 31127 14135
rect 31785 14135 31797 14138
rect 31831 14166 31843 14169
rect 32152 14169 32210 14175
rect 32152 14166 32164 14169
rect 31831 14138 32164 14166
rect 31831 14135 31843 14138
rect 31785 14129 31843 14135
rect 32152 14135 32164 14138
rect 32198 14135 32210 14169
rect 32152 14129 32210 14135
rect 32240 14172 32930 14178
rect 32240 14124 32252 14172
rect 32300 14124 32930 14172
rect 32240 14118 32930 14124
rect 28009 14101 28139 14107
rect 28009 14067 28021 14101
rect 28055 14067 28093 14101
rect 28127 14098 28139 14101
rect 28669 14101 28787 14107
rect 28669 14098 28741 14101
rect 28127 14070 28741 14098
rect 28127 14067 28139 14070
rect 28009 14061 28139 14067
rect 28729 14067 28741 14070
rect 28775 14067 28787 14101
rect 30793 14101 30916 14107
rect 28729 14061 28787 14067
rect 29526 14064 29586 14070
rect 30793 14067 30805 14101
rect 30839 14098 30916 14101
rect 31441 14101 31571 14107
rect 31441 14098 31453 14101
rect 30839 14070 31453 14098
rect 30839 14067 30851 14070
rect 29520 14004 29526 14064
rect 29586 14004 29592 14064
rect 30793 14061 30851 14067
rect 31441 14067 31453 14070
rect 31487 14067 31525 14101
rect 31559 14067 31571 14101
rect 31441 14061 31571 14067
rect 29526 13998 29586 14004
rect 26930 13986 26994 13998
rect 26667 13979 26775 13985
rect 26667 13945 26679 13979
rect 26763 13945 26775 13979
rect 26667 13939 26775 13945
rect 26564 13856 26575 13895
rect 26351 13719 26364 13752
rect 26151 13669 26259 13675
rect 26151 13635 26163 13669
rect 26247 13635 26259 13669
rect 26151 13629 26259 13635
rect 26174 13578 26234 13629
rect 25916 13518 26234 13578
rect 25030 13326 25224 13506
rect 25916 13326 25976 13518
rect 26046 13326 26106 13518
rect 26174 13326 26234 13518
rect 26304 13442 26364 13719
rect 26569 13719 26575 13856
rect 26609 13856 26624 13895
rect 26827 13895 26873 13907
rect 26609 13719 26615 13856
rect 26827 13766 26833 13895
rect 26569 13707 26615 13719
rect 26820 13719 26833 13766
rect 26867 13766 26873 13895
rect 26867 13719 26880 13766
rect 26409 13669 26517 13675
rect 26409 13635 26421 13669
rect 26505 13635 26517 13669
rect 26409 13629 26517 13635
rect 26667 13669 26775 13675
rect 26667 13635 26679 13669
rect 26763 13635 26775 13669
rect 26667 13629 26775 13635
rect 26442 13444 26502 13629
rect 26686 13580 26746 13629
rect 26820 13580 26880 13719
rect 26930 13630 26946 13986
rect 26980 13630 26994 13986
rect 26930 13580 26994 13630
rect 26686 13520 26994 13580
rect 26298 13382 26304 13442
rect 26364 13382 26370 13442
rect 26436 13384 26442 13444
rect 26502 13384 26508 13444
rect 26686 13326 26746 13520
rect 26820 13326 26880 13520
rect 26930 13326 26994 13520
rect 27260 13931 32320 13962
rect 27260 13897 27289 13931
rect 27323 13897 27381 13931
rect 27415 13897 27473 13931
rect 27507 13897 27565 13931
rect 27599 13897 27657 13931
rect 27691 13897 27749 13931
rect 27783 13897 27841 13931
rect 27875 13897 27933 13931
rect 27967 13897 28025 13931
rect 28059 13897 28117 13931
rect 28151 13897 28209 13931
rect 28243 13897 28301 13931
rect 28335 13897 28393 13931
rect 28427 13897 28485 13931
rect 28519 13897 28577 13931
rect 28611 13897 28669 13931
rect 28703 13897 28761 13931
rect 28795 13897 28853 13931
rect 28887 13897 28945 13931
rect 28979 13897 29037 13931
rect 29071 13897 29129 13931
rect 29163 13897 29221 13931
rect 29255 13897 29313 13931
rect 29347 13897 29405 13931
rect 29439 13897 29497 13931
rect 29531 13897 29589 13931
rect 29623 13897 29681 13931
rect 29715 13897 29773 13931
rect 29807 13897 29865 13931
rect 29899 13897 29957 13931
rect 29991 13897 30049 13931
rect 30083 13897 30141 13931
rect 30175 13897 30233 13931
rect 30267 13897 30325 13931
rect 30359 13897 30417 13931
rect 30451 13897 30509 13931
rect 30543 13897 30601 13931
rect 30635 13897 30693 13931
rect 30727 13897 30785 13931
rect 30819 13897 30877 13931
rect 30911 13897 30969 13931
rect 31003 13897 31061 13931
rect 31095 13897 31153 13931
rect 31187 13897 31245 13931
rect 31279 13897 31337 13931
rect 31371 13897 31429 13931
rect 31463 13897 31521 13931
rect 31555 13897 31613 13931
rect 31647 13897 31705 13931
rect 31739 13897 31797 13931
rect 31831 13897 31889 13931
rect 31923 13897 31981 13931
rect 32015 13897 32073 13931
rect 32107 13897 32165 13931
rect 32199 13897 32257 13931
rect 32291 13897 32320 13931
rect 27260 13896 32320 13897
rect 27260 13866 32322 13896
rect 27260 13326 27504 13866
rect 28078 13326 28322 13866
rect 29078 13326 29322 13866
rect 30078 13326 30322 13866
rect 31078 13326 31322 13866
rect 32078 13326 32322 13866
rect 23328 13320 32784 13326
rect 23328 13220 23434 13320
rect 32678 13220 32784 13320
rect 23328 13214 32784 13220
rect 23328 13122 23440 13214
rect 23328 11254 23334 13122
rect 23434 11254 23440 13122
rect 24664 13164 24724 13170
rect 26304 13164 26364 13168
rect 24724 13162 26364 13164
rect 24724 13104 26304 13162
rect 24664 13098 24724 13104
rect 26364 13102 27730 13162
rect 26304 13096 26364 13102
rect 24238 12990 25098 13050
rect 25158 12990 25164 13050
rect 26802 12990 26808 13050
rect 26868 12990 26874 13050
rect 27240 12990 27246 13050
rect 27306 12990 27312 13050
rect 24238 12842 24298 12990
rect 24678 12932 24738 12990
rect 24492 12926 24900 12932
rect 24492 12892 24504 12926
rect 24888 12892 24900 12926
rect 24492 12886 24900 12892
rect 24238 12666 24250 12842
rect 24284 12666 24298 12842
rect 25098 12842 25158 12990
rect 25350 12926 25758 12932
rect 25350 12892 25362 12926
rect 25746 12892 25758 12926
rect 25350 12886 25758 12892
rect 26208 12926 26616 12932
rect 26208 12892 26220 12926
rect 26604 12892 26616 12926
rect 26208 12886 26616 12892
rect 25098 12792 25108 12842
rect 24238 12502 24298 12666
rect 25102 12666 25108 12792
rect 25142 12792 25158 12842
rect 25960 12842 26006 12854
rect 25142 12666 25148 12792
rect 25960 12716 25966 12842
rect 25102 12654 25148 12666
rect 25952 12666 25966 12716
rect 26000 12716 26006 12842
rect 26808 12842 26868 12990
rect 27246 12932 27306 12990
rect 27066 12926 27474 12932
rect 27066 12892 27078 12926
rect 27462 12892 27474 12926
rect 27066 12886 27474 12892
rect 26808 12802 26824 12842
rect 26000 12666 26012 12716
rect 24492 12616 24900 12622
rect 24492 12582 24504 12616
rect 24888 12582 24900 12616
rect 24492 12576 24900 12582
rect 25350 12616 25758 12622
rect 25350 12582 25362 12616
rect 25746 12582 25758 12616
rect 25350 12576 25758 12582
rect 24680 12502 24740 12576
rect 24238 12442 24740 12502
rect 25530 12498 25590 12576
rect 25952 12498 26012 12666
rect 26818 12666 26824 12802
rect 26858 12802 26868 12842
rect 27670 12842 27730 13102
rect 32672 13122 32784 13214
rect 28520 12990 28526 13050
rect 28586 12990 28592 13050
rect 30238 12990 30244 13050
rect 30304 12990 32020 13050
rect 27924 12926 28332 12932
rect 27924 12892 27936 12926
rect 28320 12892 28332 12926
rect 27924 12886 28332 12892
rect 27670 12812 27682 12842
rect 26858 12666 26864 12802
rect 26818 12654 26864 12666
rect 27676 12666 27682 12812
rect 27716 12812 27730 12842
rect 28526 12842 28586 12990
rect 28782 12926 29190 12932
rect 28782 12892 28794 12926
rect 29178 12892 29190 12926
rect 28782 12886 29190 12892
rect 29640 12926 30048 12932
rect 29640 12892 29652 12926
rect 30036 12892 30048 12926
rect 29640 12886 30048 12892
rect 27716 12666 27722 12812
rect 28526 12806 28540 12842
rect 27676 12654 27722 12666
rect 28534 12666 28540 12806
rect 28574 12806 28586 12842
rect 29392 12842 29438 12854
rect 28574 12666 28580 12806
rect 29392 12704 29398 12842
rect 28534 12654 28580 12666
rect 29386 12666 29398 12704
rect 29432 12704 29438 12842
rect 30244 12842 30304 12990
rect 31536 12932 31596 12990
rect 30498 12926 30906 12932
rect 30498 12892 30510 12926
rect 30894 12892 30906 12926
rect 30498 12886 30906 12892
rect 31356 12926 31764 12932
rect 31356 12892 31368 12926
rect 31752 12892 31764 12926
rect 31356 12886 31764 12892
rect 30244 12796 30256 12842
rect 29432 12666 29446 12704
rect 26208 12616 26616 12622
rect 26208 12582 26220 12616
rect 26604 12582 26616 12616
rect 26208 12576 26616 12582
rect 27066 12616 27474 12622
rect 27066 12582 27078 12616
rect 27462 12582 27474 12616
rect 27066 12576 27474 12582
rect 27924 12616 28332 12622
rect 27924 12582 27936 12616
rect 28320 12582 28332 12616
rect 27924 12576 28332 12582
rect 28782 12616 29190 12622
rect 28782 12582 28794 12616
rect 29178 12582 29190 12616
rect 28782 12576 29190 12582
rect 26378 12498 26438 12576
rect 28102 12498 28162 12576
rect 28966 12498 29026 12576
rect 29386 12498 29446 12666
rect 30250 12666 30256 12796
rect 30290 12796 30304 12842
rect 31108 12842 31154 12854
rect 30290 12666 30296 12796
rect 31108 12714 31114 12842
rect 30250 12654 30296 12666
rect 31104 12666 31114 12714
rect 31148 12714 31154 12842
rect 31960 12842 32020 12990
rect 31148 12666 31164 12714
rect 29640 12616 30048 12622
rect 29640 12582 29652 12616
rect 30036 12582 30048 12616
rect 29640 12576 30048 12582
rect 30498 12616 30906 12622
rect 30498 12582 30510 12616
rect 30894 12582 30906 12616
rect 30498 12576 30906 12582
rect 29818 12498 29878 12576
rect 30672 12498 30732 12576
rect 31104 12498 31164 12666
rect 31960 12666 31972 12842
rect 32006 12666 32020 12842
rect 31356 12616 31764 12622
rect 31356 12582 31368 12616
rect 31752 12582 31764 12616
rect 31356 12576 31764 12582
rect 24238 12260 24298 12442
rect 24680 12350 24740 12442
rect 25090 12438 25096 12498
rect 25156 12438 25162 12498
rect 25524 12438 25530 12498
rect 25590 12438 25596 12498
rect 25946 12438 25952 12498
rect 26012 12438 26018 12498
rect 26372 12438 26378 12498
rect 26438 12438 26444 12498
rect 26806 12438 26812 12498
rect 26872 12438 26878 12498
rect 27240 12438 27246 12498
rect 27306 12438 27312 12498
rect 28096 12438 28102 12498
rect 28162 12438 28168 12498
rect 28960 12438 28966 12498
rect 29026 12438 29032 12498
rect 29380 12438 29386 12498
rect 29446 12438 29452 12498
rect 29812 12438 29818 12498
rect 29878 12438 29884 12498
rect 30242 12438 30248 12498
rect 30308 12438 30314 12498
rect 30666 12438 30672 12498
rect 30732 12438 30738 12498
rect 31098 12438 31104 12498
rect 31164 12438 31170 12498
rect 31544 12494 31604 12576
rect 31960 12494 32020 12666
rect 24492 12344 24900 12350
rect 24492 12310 24504 12344
rect 24888 12310 24900 12344
rect 24492 12304 24900 12310
rect 24238 12084 24250 12260
rect 24284 12084 24298 12260
rect 25096 12260 25156 12438
rect 25530 12350 25590 12438
rect 26378 12350 26438 12438
rect 25350 12344 25758 12350
rect 25350 12310 25362 12344
rect 25746 12310 25758 12344
rect 25350 12304 25758 12310
rect 26208 12344 26616 12350
rect 26208 12310 26220 12344
rect 26604 12310 26616 12344
rect 26208 12304 26616 12310
rect 25096 12220 25108 12260
rect 24238 11934 24298 12084
rect 25102 12084 25108 12220
rect 25142 12220 25156 12260
rect 25960 12260 26006 12272
rect 25142 12084 25148 12220
rect 25960 12138 25966 12260
rect 25102 12072 25148 12084
rect 25954 12084 25966 12138
rect 26000 12138 26006 12260
rect 26812 12260 26872 12438
rect 27246 12350 27306 12438
rect 28102 12350 28162 12438
rect 29818 12350 29878 12438
rect 27066 12344 27474 12350
rect 27066 12310 27078 12344
rect 27462 12310 27474 12344
rect 27066 12304 27474 12310
rect 27924 12344 28332 12350
rect 27924 12310 27936 12344
rect 28320 12310 28332 12344
rect 27924 12304 28332 12310
rect 28782 12344 29190 12350
rect 28782 12310 28794 12344
rect 29178 12310 29190 12344
rect 28782 12304 29190 12310
rect 29640 12344 30048 12350
rect 29640 12310 29652 12344
rect 30036 12310 30048 12344
rect 29640 12304 30048 12310
rect 26812 12202 26824 12260
rect 26000 12084 26014 12138
rect 24492 12034 24900 12040
rect 24492 12000 24504 12034
rect 24888 12000 24900 12034
rect 24492 11994 24900 12000
rect 25350 12034 25758 12040
rect 25350 12000 25362 12034
rect 25746 12000 25758 12034
rect 25350 11994 25758 12000
rect 24680 11934 24740 11994
rect 24238 11874 24740 11934
rect 24238 11756 24298 11874
rect 24680 11756 24740 11874
rect 25954 11756 26014 12084
rect 26818 12084 26824 12202
rect 26858 12202 26872 12260
rect 27676 12260 27722 12272
rect 26858 12084 26864 12202
rect 27676 12102 27682 12260
rect 26818 12072 26864 12084
rect 27670 12084 27682 12102
rect 27716 12102 27722 12260
rect 28534 12260 28580 12272
rect 28534 12142 28540 12260
rect 27716 12084 27730 12102
rect 26208 12034 26616 12040
rect 26208 12000 26220 12034
rect 26604 12000 26616 12034
rect 26208 11994 26616 12000
rect 27066 12034 27474 12040
rect 27066 12000 27078 12034
rect 27462 12000 27474 12034
rect 27066 11994 27474 12000
rect 27670 11756 27730 12084
rect 28526 12084 28540 12142
rect 28574 12142 28580 12260
rect 29392 12260 29438 12272
rect 28574 12084 28586 12142
rect 29392 12138 29398 12260
rect 27924 12034 28332 12040
rect 27924 12000 27936 12034
rect 28320 12000 28332 12034
rect 27924 11994 28332 12000
rect 28526 11934 28586 12084
rect 29388 12084 29398 12138
rect 29432 12138 29438 12260
rect 30248 12260 30308 12438
rect 30672 12350 30732 12438
rect 31104 12432 31164 12438
rect 31544 12434 32020 12494
rect 31544 12350 31604 12434
rect 30498 12344 30906 12350
rect 30498 12310 30510 12344
rect 30894 12310 30906 12344
rect 30498 12304 30906 12310
rect 31356 12344 31764 12350
rect 31356 12310 31368 12344
rect 31752 12310 31764 12344
rect 31356 12304 31764 12310
rect 30248 12212 30256 12260
rect 29432 12084 29448 12138
rect 28782 12034 29190 12040
rect 28782 12000 28794 12034
rect 29178 12000 29190 12034
rect 28782 11994 29190 12000
rect 28520 11874 28526 11934
rect 28586 11874 28592 11934
rect 28962 11932 29022 11994
rect 29388 11932 29448 12084
rect 30250 12084 30256 12212
rect 30290 12212 30308 12260
rect 31108 12260 31154 12272
rect 30290 12084 30296 12212
rect 31108 12116 31114 12260
rect 30250 12072 30296 12084
rect 31102 12084 31114 12116
rect 31148 12116 31154 12260
rect 31960 12260 32020 12434
rect 31148 12084 31162 12116
rect 29640 12034 30048 12040
rect 29640 12000 29652 12034
rect 30036 12000 30048 12034
rect 29640 11994 30048 12000
rect 30498 12034 30906 12040
rect 30498 12000 30510 12034
rect 30894 12000 30906 12034
rect 30498 11994 30906 12000
rect 28962 11872 29448 11932
rect 28962 11756 29022 11872
rect 29388 11756 29448 11872
rect 31102 11946 31162 12084
rect 31960 12084 31972 12260
rect 32006 12084 32020 12260
rect 31356 12034 31764 12040
rect 31356 12000 31368 12034
rect 31752 12000 31764 12034
rect 31356 11994 31764 12000
rect 31536 11946 31596 11994
rect 31960 11946 32020 12084
rect 31102 11886 32020 11946
rect 31102 11756 31162 11886
rect 31536 11756 31596 11886
rect 31960 11756 32020 11886
rect 24136 11716 32076 11756
rect 24136 11572 24176 11716
rect 32038 11572 32076 11716
rect 24136 11542 32076 11572
rect 23328 11162 23440 11254
rect 24040 11162 24050 11462
rect 32062 11162 32072 11462
rect 32672 11254 32678 13122
rect 32778 11254 32784 13122
rect 32672 11162 32784 11254
rect 23328 11156 32784 11162
rect 23328 11056 23434 11156
rect 32678 11056 32784 11156
rect 23328 11050 32784 11056
rect 12954 10734 21990 10740
rect 12954 10634 13060 10734
rect 21884 10634 21990 10734
rect 12954 10628 21990 10634
rect 12954 10546 13066 10628
rect 12954 9122 12960 10546
rect 13060 9122 13066 10546
rect 13448 10328 13458 10628
rect 21190 10328 21200 10628
rect 21878 10546 21990 10628
rect 15084 10150 20056 10180
rect 15084 10064 15134 10150
rect 15230 10064 15714 10150
rect 15810 10064 16314 10150
rect 16410 10064 16914 10150
rect 17010 10064 17514 10150
rect 17610 10064 18114 10150
rect 18210 10064 18714 10150
rect 18810 10064 19314 10150
rect 19410 10064 19914 10150
rect 20010 10064 20056 10150
rect 15084 10036 20056 10064
rect 15148 9656 15208 10036
rect 15388 9746 15448 10036
rect 15838 9812 19048 9872
rect 19108 9812 19114 9872
rect 15838 9746 15898 9812
rect 16300 9746 16360 9812
rect 16754 9746 16814 9812
rect 17216 9746 17276 9812
rect 17670 9746 17730 9812
rect 18120 9746 18180 9812
rect 18586 9746 18646 9812
rect 19042 9746 19102 9812
rect 15310 9740 15518 9746
rect 15310 9706 15322 9740
rect 15506 9706 15518 9740
rect 15310 9700 15518 9706
rect 15768 9740 15976 9746
rect 15768 9706 15780 9740
rect 15964 9706 15976 9740
rect 15768 9700 15976 9706
rect 16226 9740 16434 9746
rect 16226 9706 16238 9740
rect 16422 9706 16434 9740
rect 16226 9700 16434 9706
rect 16684 9740 16892 9746
rect 16684 9706 16696 9740
rect 16880 9706 16892 9740
rect 16684 9700 16892 9706
rect 17142 9740 17350 9746
rect 17142 9706 17154 9740
rect 17338 9706 17350 9740
rect 17142 9700 17350 9706
rect 17600 9740 17808 9746
rect 17600 9706 17612 9740
rect 17796 9706 17808 9740
rect 17600 9700 17808 9706
rect 18058 9740 18266 9746
rect 18058 9706 18070 9740
rect 18254 9706 18266 9740
rect 18058 9700 18266 9706
rect 18516 9740 18724 9746
rect 18516 9706 18528 9740
rect 18712 9706 18724 9740
rect 18516 9700 18724 9706
rect 18974 9740 19182 9746
rect 18974 9706 18986 9740
rect 19170 9706 19182 9740
rect 18974 9700 19182 9706
rect 15148 9626 15168 9656
rect 15162 9500 15168 9626
rect 12954 9040 13066 9122
rect 15156 9480 15168 9500
rect 15202 9500 15208 9656
rect 15620 9656 15666 9668
rect 15620 9508 15626 9656
rect 15202 9480 15216 9500
rect 15156 9040 15216 9480
rect 15612 9480 15626 9508
rect 15660 9508 15666 9656
rect 16078 9656 16124 9668
rect 15660 9480 15672 9508
rect 15310 9430 15518 9436
rect 15310 9396 15322 9430
rect 15506 9396 15518 9430
rect 15310 9390 15518 9396
rect 15384 9040 15444 9390
rect 15612 9192 15672 9480
rect 16078 9480 16084 9656
rect 16118 9480 16124 9656
rect 16078 9468 16124 9480
rect 16536 9656 16582 9668
rect 16536 9480 16542 9656
rect 16576 9480 16582 9656
rect 16536 9468 16582 9480
rect 16994 9656 17040 9668
rect 16994 9480 17000 9656
rect 17034 9480 17040 9656
rect 16994 9468 17040 9480
rect 17452 9656 17498 9668
rect 17452 9480 17458 9656
rect 17492 9480 17498 9656
rect 17452 9468 17498 9480
rect 17910 9656 17956 9668
rect 17910 9480 17916 9656
rect 17950 9480 17956 9656
rect 17910 9468 17956 9480
rect 18368 9656 18414 9668
rect 18368 9480 18374 9656
rect 18408 9480 18414 9656
rect 18368 9468 18414 9480
rect 18826 9656 18872 9668
rect 18826 9480 18832 9656
rect 18866 9480 18872 9656
rect 19276 9656 19336 10036
rect 19502 9746 19562 10036
rect 19432 9740 19640 9746
rect 19432 9706 19444 9740
rect 19628 9706 19640 9740
rect 19432 9700 19640 9706
rect 19276 9628 19290 9656
rect 19284 9500 19290 9628
rect 18826 9468 18872 9480
rect 19282 9480 19290 9500
rect 19324 9628 19336 9656
rect 19742 9656 19802 10036
rect 19324 9500 19330 9628
rect 19324 9480 19342 9500
rect 15768 9430 15976 9436
rect 15768 9396 15780 9430
rect 15964 9396 15976 9430
rect 15768 9390 15976 9396
rect 16226 9430 16434 9436
rect 16226 9396 16238 9430
rect 16422 9396 16434 9430
rect 16226 9390 16434 9396
rect 16684 9430 16892 9436
rect 16684 9396 16696 9430
rect 16880 9396 16892 9430
rect 16684 9390 16892 9396
rect 17142 9430 17350 9436
rect 17142 9396 17154 9430
rect 17338 9396 17350 9430
rect 17142 9390 17350 9396
rect 17600 9430 17808 9436
rect 17600 9396 17612 9430
rect 17796 9396 17808 9430
rect 17600 9390 17808 9396
rect 18058 9430 18266 9436
rect 18058 9396 18070 9430
rect 18254 9396 18266 9430
rect 18058 9390 18266 9396
rect 18516 9430 18724 9436
rect 18516 9396 18528 9430
rect 18712 9396 18724 9430
rect 18516 9390 18724 9396
rect 18974 9430 19182 9436
rect 18974 9396 18986 9430
rect 19170 9396 19182 9430
rect 18974 9390 19182 9396
rect 15844 9318 15910 9390
rect 16306 9318 16372 9390
rect 16760 9318 16826 9390
rect 17222 9318 17288 9390
rect 17676 9318 17742 9390
rect 18126 9318 18192 9390
rect 18592 9318 18658 9390
rect 19048 9318 19114 9390
rect 15844 9252 19114 9318
rect 15612 9126 15672 9132
rect 19282 9040 19342 9480
rect 19742 9480 19748 9656
rect 19782 9480 19802 9656
rect 19432 9430 19640 9436
rect 19432 9396 19444 9430
rect 19628 9396 19640 9430
rect 19432 9390 19640 9396
rect 19510 9040 19570 9390
rect 19742 9040 19802 9480
rect 21878 9122 21884 10546
rect 21984 9122 21990 10546
rect 21878 9040 21990 9122
rect 12954 9034 21990 9040
rect 12954 8934 13060 9034
rect 21884 8934 21990 9034
rect 12954 8928 21990 8934
rect 23536 10734 28992 10740
rect 23536 10634 23642 10734
rect 28886 10634 28992 10734
rect 23536 10628 28992 10634
rect 23536 10550 23648 10628
rect 23536 9038 23542 10550
rect 23642 9038 23648 10550
rect 24248 10328 24258 10628
rect 28270 10328 28280 10628
rect 28880 10550 28992 10628
rect 23846 10150 28818 10180
rect 23846 10064 23896 10150
rect 23992 10064 24476 10150
rect 24572 10064 25076 10150
rect 25172 10064 25676 10150
rect 25772 10064 26276 10150
rect 26372 10064 26876 10150
rect 26972 10064 27476 10150
rect 27572 10064 28076 10150
rect 28172 10064 28676 10150
rect 28772 10064 28818 10150
rect 23846 10036 28818 10064
rect 23910 9656 23970 10036
rect 24150 9746 24210 10036
rect 24072 9740 24280 9746
rect 24072 9706 24084 9740
rect 24268 9706 24280 9740
rect 24072 9700 24280 9706
rect 23910 9626 23930 9656
rect 23924 9500 23930 9626
rect 23536 8960 23648 9038
rect 23918 9480 23930 9500
rect 23964 9500 23970 9656
rect 24374 9656 24434 10036
rect 24600 9812 27864 9872
rect 24600 9746 24660 9812
rect 25062 9746 25122 9812
rect 25516 9746 25576 9812
rect 25978 9746 26038 9812
rect 26432 9746 26492 9812
rect 26882 9746 26942 9812
rect 27348 9746 27408 9812
rect 27804 9746 27864 9812
rect 28264 9746 28324 10036
rect 24530 9740 24738 9746
rect 24530 9706 24542 9740
rect 24726 9706 24738 9740
rect 24530 9700 24738 9706
rect 24988 9740 25196 9746
rect 24988 9706 25000 9740
rect 25184 9706 25196 9740
rect 24988 9700 25196 9706
rect 25446 9740 25654 9746
rect 25446 9706 25458 9740
rect 25642 9706 25654 9740
rect 25446 9700 25654 9706
rect 25904 9740 26112 9746
rect 25904 9706 25916 9740
rect 26100 9706 26112 9740
rect 25904 9700 26112 9706
rect 26362 9740 26570 9746
rect 26362 9706 26374 9740
rect 26558 9706 26570 9740
rect 26362 9700 26570 9706
rect 26820 9740 27028 9746
rect 26820 9706 26832 9740
rect 27016 9706 27028 9740
rect 26820 9700 27028 9706
rect 27278 9740 27486 9746
rect 27278 9706 27290 9740
rect 27474 9706 27486 9740
rect 27278 9700 27486 9706
rect 27736 9740 27944 9746
rect 27736 9706 27748 9740
rect 27932 9706 27944 9740
rect 27736 9700 27944 9706
rect 28194 9740 28402 9746
rect 28194 9706 28206 9740
rect 28390 9706 28402 9740
rect 28194 9700 28402 9706
rect 23964 9480 23978 9500
rect 23918 8960 23978 9480
rect 24374 9480 24388 9656
rect 24422 9480 24434 9656
rect 24072 9430 24280 9436
rect 24072 9396 24084 9430
rect 24268 9396 24280 9430
rect 24072 9390 24280 9396
rect 24146 8960 24206 9390
rect 24374 8960 24434 9480
rect 24840 9656 24886 9668
rect 24840 9480 24846 9656
rect 24880 9480 24886 9656
rect 24840 9468 24886 9480
rect 25298 9656 25344 9668
rect 25298 9480 25304 9656
rect 25338 9480 25344 9656
rect 25298 9468 25344 9480
rect 25756 9656 25802 9668
rect 25756 9480 25762 9656
rect 25796 9480 25802 9656
rect 25756 9468 25802 9480
rect 26214 9656 26260 9668
rect 26214 9480 26220 9656
rect 26254 9480 26260 9656
rect 26214 9468 26260 9480
rect 26672 9656 26718 9668
rect 26672 9480 26678 9656
rect 26712 9480 26718 9656
rect 26672 9468 26718 9480
rect 27130 9656 27176 9668
rect 27130 9480 27136 9656
rect 27170 9480 27176 9656
rect 27130 9468 27176 9480
rect 27588 9656 27634 9668
rect 27588 9480 27594 9656
rect 27628 9480 27634 9656
rect 28046 9656 28092 9668
rect 28046 9534 28052 9656
rect 27588 9468 27634 9480
rect 28038 9480 28052 9534
rect 28086 9534 28092 9656
rect 28504 9656 28564 10036
rect 28086 9480 28098 9534
rect 24530 9430 24738 9436
rect 24530 9396 24542 9430
rect 24726 9396 24738 9430
rect 24530 9390 24738 9396
rect 24988 9430 25196 9436
rect 24988 9396 25000 9430
rect 25184 9396 25196 9430
rect 24988 9390 25196 9396
rect 25446 9430 25654 9436
rect 25446 9396 25458 9430
rect 25642 9396 25654 9430
rect 25446 9390 25654 9396
rect 25904 9430 26112 9436
rect 25904 9396 25916 9430
rect 26100 9396 26112 9430
rect 25904 9390 26112 9396
rect 26362 9430 26570 9436
rect 26362 9396 26374 9430
rect 26558 9396 26570 9430
rect 26362 9390 26570 9396
rect 26820 9430 27028 9436
rect 26820 9396 26832 9430
rect 27016 9396 27028 9430
rect 26820 9390 27028 9396
rect 27278 9430 27486 9436
rect 27278 9396 27290 9430
rect 27474 9396 27486 9430
rect 27278 9390 27486 9396
rect 27736 9430 27944 9436
rect 27736 9396 27748 9430
rect 27932 9396 27944 9430
rect 27736 9390 27944 9396
rect 24600 9318 24660 9390
rect 25062 9318 25122 9390
rect 25516 9320 25576 9390
rect 25510 9318 25516 9320
rect 24593 9258 24600 9318
rect 24660 9258 25062 9318
rect 25122 9260 25516 9318
rect 25576 9318 25582 9320
rect 25978 9318 26038 9390
rect 26432 9318 26492 9390
rect 26882 9318 26942 9390
rect 27348 9318 27408 9390
rect 27804 9318 27864 9390
rect 25576 9260 25978 9318
rect 25122 9258 25978 9260
rect 26038 9258 26432 9318
rect 26492 9258 26882 9318
rect 26942 9258 27348 9318
rect 27408 9258 27804 9318
rect 27864 9258 27871 9318
rect 24593 9252 27871 9258
rect 28038 9110 28098 9480
rect 28504 9480 28510 9656
rect 28544 9480 28564 9656
rect 28194 9430 28402 9436
rect 28194 9396 28206 9430
rect 28390 9396 28402 9430
rect 28194 9390 28402 9396
rect 28032 9050 28038 9110
rect 28098 9050 28104 9110
rect 28272 8960 28332 9390
rect 28504 8960 28564 9480
rect 28880 9038 28886 10550
rect 28986 9038 28992 10550
rect 28880 8962 28992 9038
rect 30210 8996 36076 9008
rect 30210 8977 33086 8996
rect 33182 8977 36076 8996
rect 28880 8960 29812 8962
rect 23536 8954 29812 8960
rect 23536 8854 23642 8954
rect 28886 8931 29812 8954
rect 28886 8897 29105 8931
rect 29139 8897 29197 8931
rect 29231 8897 29289 8931
rect 29323 8897 29381 8931
rect 29415 8897 29473 8931
rect 29507 8897 29565 8931
rect 29599 8897 29657 8931
rect 29691 8897 29749 8931
rect 29783 8897 29812 8931
rect 30210 8943 30239 8977
rect 30273 8943 30581 8977
rect 30615 8943 30673 8977
rect 30707 8943 30765 8977
rect 30799 8943 30857 8977
rect 30891 8943 30949 8977
rect 30983 8943 31041 8977
rect 31075 8943 31133 8977
rect 31167 8943 31225 8977
rect 31259 8943 31317 8977
rect 31351 8943 31409 8977
rect 31443 8943 31501 8977
rect 31535 8943 31593 8977
rect 31627 8943 31685 8977
rect 31719 8943 31777 8977
rect 31811 8943 31869 8977
rect 31903 8943 31961 8977
rect 31995 8943 32053 8977
rect 32087 8943 32145 8977
rect 32179 8943 32237 8977
rect 32271 8943 32329 8977
rect 32363 8943 32421 8977
rect 32455 8943 32513 8977
rect 32547 8943 32605 8977
rect 32639 8943 32697 8977
rect 32731 8943 32789 8977
rect 32823 8943 32881 8977
rect 32915 8943 32973 8977
rect 33007 8943 33086 8977
rect 33182 8943 36013 8977
rect 36047 8943 36076 8977
rect 30210 8924 33086 8943
rect 33182 8924 36076 8943
rect 30210 8912 36076 8924
rect 28886 8866 29812 8897
rect 28886 8854 28992 8866
rect 23536 8848 28992 8854
rect 30666 8807 30724 8813
rect 28038 8768 28098 8774
rect 30666 8773 30678 8807
rect 30712 8804 30724 8807
rect 31086 8807 31144 8813
rect 31086 8804 31098 8807
rect 30712 8776 31098 8804
rect 30712 8773 30724 8776
rect 22768 8708 28038 8768
rect 28098 8708 29100 8768
rect 30666 8767 30724 8773
rect 31086 8773 31098 8776
rect 31132 8804 31144 8807
rect 31400 8807 31458 8813
rect 31400 8804 31412 8807
rect 31132 8776 31412 8804
rect 31132 8773 31144 8776
rect 31086 8767 31144 8773
rect 31400 8773 31412 8776
rect 31446 8773 31458 8807
rect 31400 8767 31458 8773
rect 12954 8698 21990 8704
rect 12954 8598 13060 8698
rect 21884 8598 21990 8698
rect 12954 8592 21990 8598
rect 12954 8400 13066 8592
rect 12954 5064 12960 8400
rect 13060 8038 13066 8400
rect 13324 8038 13384 8592
rect 13552 8038 13612 8592
rect 13778 8038 13838 8592
rect 14236 8450 20712 8510
rect 13060 7978 13838 8038
rect 14002 7978 14008 8038
rect 14068 7978 14074 8038
rect 13060 5064 13066 7978
rect 13324 7805 13384 7978
rect 13552 7904 13612 7978
rect 13478 7898 13686 7904
rect 13478 7864 13490 7898
rect 13674 7864 13686 7898
rect 13478 7858 13686 7864
rect 13324 7746 13336 7805
rect 13330 6262 13336 7746
rect 13322 6229 13336 6262
rect 13370 7746 13384 7805
rect 13778 7805 13838 7978
rect 14008 7904 14068 7978
rect 13936 7898 14144 7904
rect 13936 7864 13948 7898
rect 14132 7864 14144 7898
rect 13936 7858 14144 7864
rect 13778 7762 13794 7805
rect 13370 6262 13376 7746
rect 13788 6294 13794 7762
rect 13370 6229 13382 6262
rect 13322 5442 13382 6229
rect 13780 6229 13794 6294
rect 13828 7762 13838 7805
rect 14236 7805 14296 8450
rect 15154 8326 19798 8386
rect 14458 7978 14464 8038
rect 14524 7978 14530 8038
rect 14918 7978 14924 8038
rect 14984 7978 14990 8038
rect 14464 7904 14524 7978
rect 14924 7904 14984 7978
rect 14394 7898 14602 7904
rect 14394 7864 14406 7898
rect 14590 7864 14602 7898
rect 14394 7858 14602 7864
rect 14852 7898 15060 7904
rect 14852 7864 14864 7898
rect 15048 7864 15060 7898
rect 14852 7858 15060 7864
rect 13828 6294 13834 7762
rect 14236 7722 14252 7805
rect 13828 6229 13840 6294
rect 13478 6170 13686 6176
rect 13478 6136 13490 6170
rect 13674 6136 13686 6170
rect 13478 6130 13686 6136
rect 13554 5442 13614 6130
rect 13780 5442 13840 6229
rect 14246 6229 14252 7722
rect 14286 7722 14296 7805
rect 14704 7805 14750 7817
rect 14286 6229 14292 7722
rect 14704 6288 14710 7805
rect 14246 6217 14292 6229
rect 14696 6229 14710 6288
rect 14744 6288 14750 7805
rect 15154 7805 15214 8326
rect 16062 8202 18878 8262
rect 15374 7978 15380 8038
rect 15440 7978 15446 8038
rect 15832 7978 15838 8038
rect 15898 7978 15904 8038
rect 15380 7904 15440 7978
rect 15838 7904 15898 7978
rect 15310 7898 15518 7904
rect 15310 7864 15322 7898
rect 15506 7864 15518 7898
rect 15310 7858 15518 7864
rect 15768 7898 15976 7904
rect 15768 7864 15780 7898
rect 15964 7864 15976 7898
rect 15768 7858 15976 7864
rect 16062 7817 16122 8202
rect 16986 8086 17964 8146
rect 16296 7978 16302 8038
rect 16362 7978 16368 8038
rect 16750 7978 16756 8038
rect 16816 7978 16822 8038
rect 16302 7904 16362 7978
rect 16756 7904 16816 7978
rect 16226 7898 16434 7904
rect 16226 7864 16238 7898
rect 16422 7864 16434 7898
rect 16226 7858 16434 7864
rect 16684 7898 16892 7904
rect 16684 7864 16696 7898
rect 16880 7864 16892 7898
rect 16684 7858 16892 7864
rect 15154 7728 15168 7805
rect 14744 6229 14756 6288
rect 13936 6170 14144 6176
rect 13936 6136 13948 6170
rect 14132 6136 14144 6170
rect 13936 6130 14144 6136
rect 14394 6170 14602 6176
rect 14394 6136 14406 6170
rect 14590 6136 14602 6170
rect 14394 6130 14602 6136
rect 14012 6064 14072 6130
rect 14468 6064 14528 6130
rect 14006 6004 14012 6064
rect 14072 6004 14078 6064
rect 14462 6004 14468 6064
rect 14528 6004 14534 6064
rect 14696 5696 14756 6229
rect 15162 6229 15168 7728
rect 15202 7728 15214 7805
rect 15620 7805 15666 7817
rect 15202 6229 15208 7728
rect 15620 6290 15626 7805
rect 15162 6217 15208 6229
rect 15612 6229 15626 6290
rect 15660 6290 15666 7805
rect 16062 7805 16124 7817
rect 16062 7734 16084 7805
rect 15660 6229 15672 6290
rect 14852 6170 15060 6176
rect 14852 6136 14864 6170
rect 15048 6136 15060 6170
rect 14852 6130 15060 6136
rect 15310 6170 15518 6176
rect 15310 6136 15322 6170
rect 15506 6136 15518 6170
rect 15310 6130 15518 6136
rect 14928 6064 14988 6130
rect 15384 6064 15444 6130
rect 14922 6004 14928 6064
rect 14988 6004 14994 6064
rect 15378 6004 15384 6064
rect 15444 6004 15450 6064
rect 15612 5830 15672 6229
rect 16078 6229 16084 7734
rect 16118 6229 16124 7805
rect 16536 7805 16582 7817
rect 16536 6308 16542 7805
rect 16078 6217 16124 6229
rect 16528 6229 16542 6308
rect 16576 6308 16582 7805
rect 16986 7805 17046 8086
rect 17210 7978 17216 8038
rect 17276 7978 17282 8038
rect 17440 7978 17446 8038
rect 17506 7978 17512 8038
rect 17668 7978 17674 8038
rect 17734 7978 17740 8038
rect 17216 7904 17276 7978
rect 17142 7898 17350 7904
rect 17142 7864 17154 7898
rect 17338 7864 17350 7898
rect 17142 7858 17350 7864
rect 16986 7726 17000 7805
rect 16576 6229 16588 6308
rect 15768 6170 15976 6176
rect 15768 6136 15780 6170
rect 15964 6136 15976 6170
rect 15768 6130 15976 6136
rect 16226 6170 16434 6176
rect 16226 6136 16238 6170
rect 16422 6136 16434 6170
rect 16226 6130 16434 6136
rect 15842 6064 15902 6130
rect 16306 6064 16366 6130
rect 15836 6004 15842 6064
rect 15902 6004 15908 6064
rect 16300 6004 16306 6064
rect 16366 6004 16372 6064
rect 16528 5954 16588 6229
rect 16994 6229 17000 7726
rect 17034 7726 17046 7805
rect 17446 7805 17506 7978
rect 17674 7904 17734 7978
rect 17600 7898 17808 7904
rect 17600 7864 17612 7898
rect 17796 7864 17808 7898
rect 17600 7858 17808 7864
rect 17446 7756 17458 7805
rect 17034 6229 17040 7726
rect 16994 6217 17040 6229
rect 17452 6229 17458 7756
rect 17492 7756 17506 7805
rect 17904 7805 17964 8086
rect 18124 7978 18130 8038
rect 18190 7978 18196 8038
rect 18584 7978 18590 8038
rect 18650 7978 18656 8038
rect 18130 7904 18190 7978
rect 18590 7904 18650 7978
rect 18058 7898 18266 7904
rect 18058 7864 18070 7898
rect 18254 7864 18266 7898
rect 18058 7858 18266 7864
rect 18516 7898 18724 7904
rect 18516 7864 18528 7898
rect 18712 7864 18724 7898
rect 18516 7858 18724 7864
rect 17904 7778 17916 7805
rect 17492 6229 17498 7756
rect 17452 6217 17498 6229
rect 17910 6229 17916 7778
rect 17950 7778 17964 7805
rect 18368 7805 18414 7817
rect 17950 6229 17956 7778
rect 18368 6274 18374 7805
rect 17910 6217 17956 6229
rect 18358 6229 18374 6274
rect 18408 6274 18414 7805
rect 18818 7805 18878 8202
rect 19040 7978 19046 8038
rect 19106 7978 19112 8038
rect 19496 7978 19502 8038
rect 19562 7978 19568 8038
rect 19046 7904 19106 7978
rect 19502 7904 19562 7978
rect 18974 7898 19182 7904
rect 18974 7864 18986 7898
rect 19170 7864 19182 7898
rect 18974 7858 19182 7864
rect 19432 7898 19640 7904
rect 19432 7864 19444 7898
rect 19628 7864 19640 7898
rect 19432 7858 19640 7864
rect 18818 7774 18832 7805
rect 18408 6229 18418 6274
rect 16684 6170 16892 6176
rect 16684 6136 16696 6170
rect 16880 6136 16892 6170
rect 16684 6130 16892 6136
rect 17142 6170 17350 6176
rect 17142 6136 17154 6170
rect 17338 6136 17350 6170
rect 17142 6130 17350 6136
rect 17600 6170 17808 6176
rect 17600 6136 17612 6170
rect 17796 6136 17808 6170
rect 17600 6130 17808 6136
rect 18058 6170 18266 6176
rect 18058 6136 18070 6170
rect 18254 6136 18266 6170
rect 18058 6130 18266 6136
rect 16756 6064 16816 6130
rect 17212 6064 17272 6130
rect 17680 6064 17740 6130
rect 18138 6064 18198 6130
rect 16750 6004 16756 6064
rect 16816 6004 16822 6064
rect 17206 6004 17212 6064
rect 17272 6004 17278 6064
rect 17674 6004 17680 6064
rect 17740 6004 17746 6064
rect 18132 6004 18138 6064
rect 18198 6004 18204 6064
rect 18358 5954 18418 6229
rect 18826 6229 18832 7774
rect 18866 7774 18878 7805
rect 19284 7805 19330 7817
rect 18866 6229 18872 7774
rect 19284 6288 19290 7805
rect 18826 6217 18872 6229
rect 19274 6229 19290 6288
rect 19324 6288 19330 7805
rect 19738 7805 19798 8326
rect 19952 7978 19958 8038
rect 20018 7978 20024 8038
rect 20410 7978 20416 8038
rect 20476 7978 20482 8038
rect 19958 7904 20018 7978
rect 20416 7904 20476 7978
rect 19890 7898 20098 7904
rect 19890 7864 19902 7898
rect 20086 7864 20098 7898
rect 19890 7858 20098 7864
rect 20348 7898 20556 7904
rect 20348 7864 20360 7898
rect 20544 7864 20556 7898
rect 20348 7858 20556 7864
rect 19738 7738 19748 7805
rect 19324 6229 19334 6288
rect 18516 6170 18724 6176
rect 18516 6136 18528 6170
rect 18712 6136 18724 6170
rect 18516 6130 18724 6136
rect 18974 6170 19182 6176
rect 18974 6136 18986 6170
rect 19170 6136 19182 6170
rect 18974 6130 19182 6136
rect 18594 6064 18654 6130
rect 19050 6064 19110 6130
rect 18588 6004 18594 6064
rect 18654 6004 18660 6064
rect 19044 6004 19050 6064
rect 19110 6004 19116 6064
rect 16528 5894 18418 5954
rect 19274 5830 19334 6229
rect 19742 6229 19748 7738
rect 19782 7738 19798 7805
rect 20200 7805 20246 7817
rect 19782 6229 19788 7738
rect 20200 6286 20206 7805
rect 19742 6217 19788 6229
rect 20194 6229 20206 6286
rect 20240 6286 20246 7805
rect 20652 7805 20712 8450
rect 21106 8038 21166 8592
rect 21338 8038 21398 8592
rect 21564 8038 21624 8592
rect 21878 8400 21990 8592
rect 21878 8038 21884 8400
rect 20870 7978 20876 8038
rect 20936 7978 20942 8038
rect 21106 7978 21884 8038
rect 20876 7904 20936 7978
rect 20806 7898 21014 7904
rect 20806 7864 20818 7898
rect 21002 7864 21014 7898
rect 20806 7858 21014 7864
rect 20652 7746 20664 7805
rect 20240 6229 20254 6286
rect 19432 6170 19640 6176
rect 19432 6136 19444 6170
rect 19628 6136 19640 6170
rect 19432 6130 19640 6136
rect 19890 6170 20098 6176
rect 19890 6136 19902 6170
rect 20086 6136 20098 6170
rect 19890 6130 20098 6136
rect 19506 6064 19566 6130
rect 19962 6064 20022 6130
rect 19500 6004 19506 6064
rect 19566 6004 19572 6064
rect 19956 6004 19962 6064
rect 20022 6004 20028 6064
rect 15612 5770 19334 5830
rect 20194 5696 20254 6229
rect 20658 6229 20664 7746
rect 20698 7746 20712 7805
rect 21106 7805 21166 7978
rect 21338 7904 21398 7978
rect 21264 7898 21472 7904
rect 21264 7864 21276 7898
rect 21460 7864 21472 7898
rect 21264 7858 21472 7864
rect 20698 6229 20704 7746
rect 21106 7744 21122 7805
rect 21116 6306 21122 7744
rect 20658 6217 20704 6229
rect 21110 6229 21122 6306
rect 21156 7744 21166 7805
rect 21564 7805 21624 7978
rect 21564 7762 21580 7805
rect 21156 6306 21162 7744
rect 21156 6229 21170 6306
rect 21574 6300 21580 7762
rect 20348 6170 20556 6176
rect 20348 6136 20360 6170
rect 20544 6136 20556 6170
rect 20348 6130 20556 6136
rect 20806 6170 21014 6176
rect 20806 6136 20818 6170
rect 21002 6136 21014 6170
rect 20806 6130 21014 6136
rect 20420 6064 20480 6130
rect 20880 6064 20940 6130
rect 20414 6004 20420 6064
rect 20480 6004 20486 6064
rect 20874 6004 20880 6064
rect 20940 6004 20946 6064
rect 14696 5636 20254 5696
rect 21110 5442 21170 6229
rect 21568 6229 21580 6300
rect 21614 7762 21624 7805
rect 21614 6300 21620 7762
rect 21614 6229 21628 6300
rect 21264 6170 21472 6176
rect 21264 6136 21276 6170
rect 21460 6136 21472 6170
rect 21264 6130 21472 6136
rect 21340 5442 21400 6130
rect 21568 5442 21628 6229
rect 21878 5442 21884 7978
rect 13294 5432 21884 5442
rect 13294 5346 13308 5432
rect 13404 5346 13908 5432
rect 14004 5346 14508 5432
rect 14604 5346 15108 5432
rect 15204 5346 15708 5432
rect 15804 5346 16308 5432
rect 16404 5346 16908 5432
rect 17004 5346 17508 5432
rect 17604 5346 18108 5432
rect 18204 5346 18708 5432
rect 18804 5346 19308 5432
rect 19404 5346 19908 5432
rect 20004 5346 20508 5432
rect 20604 5346 21108 5432
rect 21204 5346 21528 5432
rect 21624 5346 21884 5432
rect 13294 5332 21884 5346
rect 12954 4872 13066 5064
rect 13448 4872 13458 5172
rect 21190 4872 21200 5172
rect 21878 5064 21884 5332
rect 21984 5442 21990 8400
rect 21984 5332 21992 5442
rect 21984 5064 21990 5332
rect 21878 4872 21990 5064
rect 12954 4866 21990 4872
rect 12954 4766 13060 4866
rect 21884 4766 21990 4866
rect 12954 4760 21990 4766
rect 8346 4396 18802 4402
rect 8346 4296 8452 4396
rect 18696 4296 18802 4396
rect 8346 4290 18802 4296
rect 8346 4006 8458 4290
rect 8346 -1166 8352 4006
rect 8452 1184 8458 4006
rect 9058 3990 9068 4290
rect 18080 3990 18090 4290
rect 18690 4006 18802 4290
rect 9296 3816 17652 3830
rect 9296 3730 9310 3816
rect 9406 3730 9910 3816
rect 10006 3730 10510 3816
rect 10606 3730 11110 3816
rect 11206 3730 11710 3816
rect 11806 3730 12310 3816
rect 12406 3730 12910 3816
rect 13006 3730 13510 3816
rect 13606 3730 14110 3816
rect 14206 3730 14710 3816
rect 14806 3730 15310 3816
rect 15406 3730 15910 3816
rect 16006 3730 16510 3816
rect 16606 3730 17110 3816
rect 17206 3730 17530 3816
rect 17626 3730 17652 3816
rect 9296 3720 17652 3730
rect 9324 2932 9384 3720
rect 9556 3031 9616 3720
rect 9480 3025 9688 3031
rect 9480 2991 9492 3025
rect 9676 2991 9688 3025
rect 9480 2985 9688 2991
rect 9324 2900 9338 2932
rect 9332 1416 9338 2900
rect 9326 1356 9338 1416
rect 9372 2900 9384 2932
rect 9782 2932 9842 3720
rect 10698 3466 16256 3526
rect 10008 3098 10014 3158
rect 10074 3098 10080 3158
rect 10464 3098 10470 3158
rect 10530 3098 10536 3158
rect 10014 3031 10074 3098
rect 10470 3031 10530 3098
rect 9938 3025 10146 3031
rect 9938 2991 9950 3025
rect 10134 2991 10146 3025
rect 9938 2985 10146 2991
rect 10396 3025 10604 3031
rect 10396 2991 10408 3025
rect 10592 2991 10604 3025
rect 10396 2985 10604 2991
rect 9372 1416 9378 2900
rect 9782 2868 9796 2932
rect 9372 1356 9386 1416
rect 9790 1400 9796 2868
rect 9326 1184 9386 1356
rect 9780 1356 9796 1400
rect 9830 2868 9842 2932
rect 10248 2932 10294 2944
rect 9830 1400 9836 2868
rect 10248 1440 10254 2932
rect 9830 1356 9840 1400
rect 9480 1297 9688 1303
rect 9480 1263 9492 1297
rect 9676 1263 9688 1297
rect 9480 1257 9688 1263
rect 9554 1184 9614 1257
rect 9780 1184 9840 1356
rect 10238 1356 10254 1440
rect 10288 1440 10294 2932
rect 10698 2932 10758 3466
rect 11614 3332 15336 3392
rect 10924 3098 10930 3158
rect 10990 3098 10996 3158
rect 11380 3098 11386 3158
rect 11446 3098 11452 3158
rect 10930 3031 10990 3098
rect 11386 3031 11446 3098
rect 10854 3025 11062 3031
rect 10854 2991 10866 3025
rect 11050 2991 11062 3025
rect 10854 2985 11062 2991
rect 11312 3025 11520 3031
rect 11312 2991 11324 3025
rect 11508 2991 11520 3025
rect 11312 2985 11520 2991
rect 10698 2874 10712 2932
rect 10288 1356 10298 1440
rect 9938 1297 10146 1303
rect 9938 1263 9950 1297
rect 10134 1263 10146 1297
rect 9938 1257 10146 1263
rect 10010 1184 10070 1257
rect 8452 1124 9840 1184
rect 10004 1124 10010 1184
rect 10070 1124 10076 1184
rect 8452 752 8458 1124
rect 9326 752 9386 1124
rect 8452 692 9386 752
rect 10238 704 10298 1356
rect 10706 1356 10712 2874
rect 10746 2874 10758 2932
rect 11164 2932 11210 2944
rect 10746 1356 10752 2874
rect 11164 1434 11170 2932
rect 10706 1344 10752 1356
rect 11156 1356 11170 1434
rect 11204 1434 11210 2932
rect 11614 2932 11674 3332
rect 12530 3208 14420 3268
rect 11838 3098 11844 3158
rect 11904 3098 11910 3158
rect 12302 3098 12308 3158
rect 12368 3098 12374 3158
rect 11844 3031 11904 3098
rect 12308 3031 12368 3098
rect 11770 3025 11978 3031
rect 11770 2991 11782 3025
rect 11966 2991 11978 3025
rect 11770 2985 11978 2991
rect 12228 3025 12436 3031
rect 12228 2991 12240 3025
rect 12424 2991 12436 3025
rect 12228 2985 12436 2991
rect 11614 2872 11628 2932
rect 11204 1356 11216 1434
rect 10396 1297 10604 1303
rect 10396 1263 10408 1297
rect 10592 1263 10604 1297
rect 10396 1257 10604 1263
rect 10854 1297 11062 1303
rect 10854 1263 10866 1297
rect 11050 1263 11062 1297
rect 10854 1257 11062 1263
rect 10466 1184 10526 1257
rect 10926 1184 10986 1257
rect 10460 1124 10466 1184
rect 10526 1124 10532 1184
rect 10920 1124 10926 1184
rect 10986 1124 10992 1184
rect 11156 834 11216 1356
rect 11622 1356 11628 2872
rect 11662 2872 11674 2932
rect 12080 2932 12126 2944
rect 11662 1356 11668 2872
rect 12080 1428 12086 2932
rect 11622 1344 11668 1356
rect 12064 1356 12086 1428
rect 12120 1356 12126 2932
rect 12530 2932 12590 3208
rect 12752 3098 12758 3158
rect 12818 3098 12824 3158
rect 13208 3098 13214 3158
rect 13274 3098 13280 3158
rect 13676 3098 13682 3158
rect 13742 3098 13748 3158
rect 14134 3098 14140 3158
rect 14200 3098 14206 3158
rect 12758 3031 12818 3098
rect 13214 3031 13274 3098
rect 13682 3031 13742 3098
rect 14140 3031 14200 3098
rect 12686 3025 12894 3031
rect 12686 2991 12698 3025
rect 12882 2991 12894 3025
rect 12686 2985 12894 2991
rect 13144 3025 13352 3031
rect 13144 2991 13156 3025
rect 13340 2991 13352 3025
rect 13144 2985 13352 2991
rect 13602 3025 13810 3031
rect 13602 2991 13614 3025
rect 13798 2991 13810 3025
rect 13602 2985 13810 2991
rect 14060 3025 14268 3031
rect 14060 2991 14072 3025
rect 14256 2991 14268 3025
rect 14060 2985 14268 2991
rect 12530 2854 12544 2932
rect 12064 1344 12126 1356
rect 12538 1356 12544 2854
rect 12578 2854 12590 2932
rect 12996 2932 13042 2944
rect 12578 1356 12584 2854
rect 12996 1436 13002 2932
rect 12538 1344 12584 1356
rect 12988 1356 13002 1436
rect 13036 1436 13042 2932
rect 13454 2932 13500 2944
rect 13036 1356 13048 1436
rect 13454 1378 13460 2932
rect 11312 1297 11520 1303
rect 11312 1263 11324 1297
rect 11508 1263 11520 1297
rect 11312 1257 11520 1263
rect 11770 1297 11978 1303
rect 11770 1263 11782 1297
rect 11966 1263 11978 1297
rect 11770 1257 11978 1263
rect 11382 1184 11442 1257
rect 11840 1184 11900 1257
rect 11376 1124 11382 1184
rect 11442 1124 11448 1184
rect 11834 1124 11840 1184
rect 11900 1124 11906 1184
rect 12064 960 12124 1344
rect 12228 1297 12436 1303
rect 12228 1263 12240 1297
rect 12424 1263 12436 1297
rect 12228 1257 12436 1263
rect 12686 1297 12894 1303
rect 12686 1263 12698 1297
rect 12882 1263 12894 1297
rect 12686 1257 12894 1263
rect 12304 1184 12364 1257
rect 12758 1184 12818 1257
rect 12298 1124 12304 1184
rect 12364 1124 12370 1184
rect 12752 1124 12758 1184
rect 12818 1124 12824 1184
rect 12988 1076 13048 1356
rect 13450 1356 13460 1378
rect 13494 1378 13500 2932
rect 13912 2932 13958 2944
rect 13912 1384 13918 2932
rect 13494 1356 13510 1378
rect 13144 1297 13352 1303
rect 13144 1263 13156 1297
rect 13340 1263 13352 1297
rect 13144 1257 13352 1263
rect 13216 1186 13276 1257
rect 13450 1196 13510 1356
rect 13906 1356 13918 1384
rect 13952 1384 13958 2932
rect 14360 2932 14420 3208
rect 14590 3098 14596 3158
rect 14656 3098 14662 3158
rect 15046 3098 15052 3158
rect 15112 3098 15118 3158
rect 14596 3031 14656 3098
rect 15052 3031 15112 3098
rect 14518 3025 14726 3031
rect 14518 2991 14530 3025
rect 14714 2991 14726 3025
rect 14518 2985 14726 2991
rect 14976 3025 15184 3031
rect 14976 2991 14988 3025
rect 15172 2991 15184 3025
rect 14976 2985 15184 2991
rect 14360 2888 14376 2932
rect 13952 1356 13966 1384
rect 13602 1297 13810 1303
rect 13602 1263 13614 1297
rect 13798 1263 13810 1297
rect 13602 1257 13810 1263
rect 13210 1184 13282 1186
rect 13210 1124 13216 1184
rect 13276 1124 13282 1184
rect 13676 1192 13736 1257
rect 13450 1130 13510 1136
rect 13664 1186 13748 1192
rect 13664 1124 13676 1186
rect 13736 1124 13748 1186
rect 13664 1120 13748 1124
rect 13906 1076 13966 1356
rect 14370 1356 14376 2888
rect 14410 2888 14420 2932
rect 14828 2932 14874 2944
rect 14410 1356 14416 2888
rect 14828 1388 14834 2932
rect 14370 1344 14416 1356
rect 14820 1356 14834 1388
rect 14868 1388 14874 2932
rect 15276 2932 15336 3332
rect 15502 3098 15508 3158
rect 15568 3098 15574 3158
rect 15958 3098 15964 3158
rect 16024 3098 16030 3158
rect 15508 3031 15568 3098
rect 15964 3031 16024 3098
rect 15434 3025 15642 3031
rect 15434 2991 15446 3025
rect 15630 2991 15642 3025
rect 15434 2985 15642 2991
rect 15892 3025 16100 3031
rect 15892 2991 15904 3025
rect 16088 2991 16100 3025
rect 15892 2985 16100 2991
rect 15276 2874 15292 2932
rect 14868 1356 14880 1388
rect 14060 1297 14268 1303
rect 14060 1263 14072 1297
rect 14256 1263 14268 1297
rect 14060 1257 14268 1263
rect 14518 1297 14726 1303
rect 14518 1263 14530 1297
rect 14714 1263 14726 1297
rect 14518 1257 14726 1263
rect 14132 1184 14192 1257
rect 14592 1184 14652 1257
rect 14126 1124 14132 1184
rect 14192 1124 14198 1184
rect 14586 1124 14592 1184
rect 14652 1124 14658 1184
rect 12988 1016 13966 1076
rect 14820 960 14880 1356
rect 15286 1356 15292 2874
rect 15326 2874 15336 2932
rect 15744 2932 15790 2944
rect 15326 1356 15332 2874
rect 15744 1424 15750 2932
rect 15286 1344 15332 1356
rect 15740 1356 15750 1424
rect 15784 1424 15790 2932
rect 16196 2932 16256 3466
rect 16416 3098 16422 3158
rect 16482 3098 16488 3158
rect 16876 3098 16882 3158
rect 16942 3098 16948 3158
rect 16422 3031 16482 3098
rect 16882 3031 16942 3098
rect 16350 3025 16558 3031
rect 16350 2991 16362 3025
rect 16546 2991 16558 3025
rect 16350 2985 16558 2991
rect 16808 3025 17016 3031
rect 16808 2991 16820 3025
rect 17004 2991 17016 3025
rect 16808 2985 17016 2991
rect 16196 2876 16208 2932
rect 15784 1356 15800 1424
rect 14976 1297 15184 1303
rect 14976 1263 14988 1297
rect 15172 1263 15184 1297
rect 14976 1257 15184 1263
rect 15434 1297 15642 1303
rect 15434 1263 15446 1297
rect 15630 1263 15642 1297
rect 15434 1257 15642 1263
rect 15048 1184 15108 1257
rect 15504 1184 15564 1257
rect 15042 1124 15048 1184
rect 15108 1124 15114 1184
rect 15498 1124 15504 1184
rect 15564 1124 15570 1184
rect 12064 900 14880 960
rect 15740 834 15800 1356
rect 16202 1356 16208 2876
rect 16242 2876 16256 2932
rect 16660 2932 16706 2944
rect 16242 1356 16248 2876
rect 16660 1416 16666 2932
rect 16202 1344 16248 1356
rect 16654 1356 16666 1416
rect 16700 1416 16706 2932
rect 17112 2932 17172 3720
rect 17342 3031 17402 3720
rect 17266 3025 17474 3031
rect 17266 2991 17278 3025
rect 17462 2991 17474 3025
rect 17266 2985 17474 2991
rect 17112 2856 17124 2932
rect 17118 1418 17124 2856
rect 16700 1356 16714 1416
rect 15892 1297 16100 1303
rect 15892 1263 15904 1297
rect 16088 1263 16100 1297
rect 15892 1257 16100 1263
rect 16350 1297 16558 1303
rect 16350 1263 16362 1297
rect 16546 1263 16558 1297
rect 16350 1257 16558 1263
rect 15960 1184 16020 1257
rect 16418 1184 16478 1257
rect 15954 1124 15960 1184
rect 16020 1124 16026 1184
rect 16412 1124 16418 1184
rect 16478 1124 16484 1184
rect 11156 774 15800 834
rect 16654 704 16714 1356
rect 17108 1356 17124 1418
rect 17158 2856 17172 2932
rect 17570 2932 17630 3720
rect 17570 2862 17582 2932
rect 17158 1418 17164 2856
rect 17158 1356 17168 1418
rect 17576 1400 17582 2862
rect 16808 1297 17016 1303
rect 16808 1263 16820 1297
rect 17004 1263 17016 1297
rect 16808 1257 17016 1263
rect 16878 1184 16938 1257
rect 16872 1124 16878 1184
rect 16938 1124 16944 1184
rect 17108 1182 17168 1356
rect 17566 1356 17582 1400
rect 17616 2862 17630 2932
rect 17616 1400 17622 2862
rect 17616 1356 17626 1400
rect 17266 1297 17474 1303
rect 17266 1263 17278 1297
rect 17462 1263 17474 1297
rect 17266 1257 17474 1263
rect 17340 1182 17400 1257
rect 17566 1182 17626 1356
rect 18690 1182 18696 4006
rect 17108 1122 18696 1182
rect 8452 -1166 8458 692
rect 8766 267 8826 692
rect 8994 366 9054 692
rect 10238 644 16714 704
rect 17566 688 17626 1122
rect 18690 688 18696 1122
rect 17566 628 18696 688
rect 9218 538 9224 598
rect 9284 538 9290 598
rect 8921 360 9129 366
rect 8921 326 8933 360
rect 9117 326 9129 360
rect 8921 320 9129 326
rect 8766 220 8779 267
rect 8773 -888 8779 220
rect 8346 -1342 8458 -1166
rect 8766 -909 8779 -888
rect 8813 220 8826 267
rect 9224 267 9284 538
rect 9456 436 12658 496
rect 12718 436 12724 496
rect 9456 366 9516 436
rect 9918 366 9978 436
rect 10372 366 10432 436
rect 10834 366 10894 436
rect 11288 366 11348 436
rect 11738 366 11798 436
rect 12204 366 12264 436
rect 12660 366 12720 436
rect 13116 418 14284 478
rect 13116 366 13176 418
rect 9379 360 9587 366
rect 9379 326 9391 360
rect 9575 326 9587 360
rect 9379 320 9587 326
rect 9837 360 10045 366
rect 9837 326 9849 360
rect 10033 326 10045 360
rect 9837 320 10045 326
rect 10295 360 10503 366
rect 10295 326 10307 360
rect 10491 326 10503 360
rect 10295 320 10503 326
rect 10753 360 10961 366
rect 10753 326 10765 360
rect 10949 326 10961 360
rect 10753 320 10961 326
rect 11211 360 11419 366
rect 11211 326 11223 360
rect 11407 326 11419 360
rect 11211 320 11419 326
rect 11669 360 11877 366
rect 11669 326 11681 360
rect 11865 326 11877 360
rect 11669 320 11877 326
rect 12127 360 12335 366
rect 12127 326 12139 360
rect 12323 326 12335 360
rect 12127 320 12335 326
rect 12585 360 12793 366
rect 12585 326 12597 360
rect 12781 326 12793 360
rect 12585 320 12793 326
rect 13043 360 13251 366
rect 13043 326 13055 360
rect 13239 326 13251 360
rect 13043 320 13251 326
rect 8813 -888 8819 220
rect 9224 200 9237 267
rect 8813 -909 8826 -888
rect 8766 -1342 8826 -909
rect 9231 -909 9237 200
rect 9271 200 9284 267
rect 9689 267 9735 279
rect 9271 -909 9277 200
rect 9231 -921 9277 -909
rect 9689 -909 9695 267
rect 9729 -909 9735 267
rect 9689 -921 9735 -909
rect 10147 267 10193 279
rect 10147 -909 10153 267
rect 10187 -909 10193 267
rect 10147 -921 10193 -909
rect 10605 267 10651 279
rect 10605 -909 10611 267
rect 10645 -909 10651 267
rect 10605 -921 10651 -909
rect 11063 267 11109 279
rect 11063 -909 11069 267
rect 11103 -909 11109 267
rect 11063 -921 11109 -909
rect 11521 267 11567 279
rect 11521 -909 11527 267
rect 11561 -909 11567 267
rect 11521 -921 11567 -909
rect 11979 267 12025 279
rect 11979 -909 11985 267
rect 12019 -909 12025 267
rect 11979 -921 12025 -909
rect 12437 267 12483 279
rect 12437 -909 12443 267
rect 12477 -909 12483 267
rect 12895 267 12941 279
rect 12895 -842 12901 267
rect 12437 -921 12483 -909
rect 12886 -909 12901 -842
rect 12935 -842 12941 267
rect 13346 267 13406 418
rect 13346 252 13359 267
rect 12935 -909 12946 -842
rect 13353 -874 13359 252
rect 8921 -968 9129 -962
rect 8921 -1002 8933 -968
rect 9117 -1002 9129 -968
rect 8921 -1008 9129 -1002
rect 9379 -968 9587 -962
rect 9379 -1002 9391 -968
rect 9575 -1002 9587 -968
rect 9379 -1008 9587 -1002
rect 9837 -968 10045 -962
rect 9837 -1002 9849 -968
rect 10033 -1002 10045 -968
rect 9837 -1008 10045 -1002
rect 10295 -968 10503 -962
rect 10295 -1002 10307 -968
rect 10491 -1002 10503 -968
rect 10295 -1008 10503 -1002
rect 10753 -968 10961 -962
rect 10753 -1002 10765 -968
rect 10949 -1002 10961 -968
rect 10753 -1008 10961 -1002
rect 11211 -968 11419 -962
rect 11211 -1002 11223 -968
rect 11407 -1002 11419 -968
rect 11211 -1008 11419 -1002
rect 11669 -968 11877 -962
rect 11669 -1002 11681 -968
rect 11865 -1002 11877 -968
rect 11669 -1008 11877 -1002
rect 12127 -968 12335 -962
rect 12127 -1002 12139 -968
rect 12323 -1002 12335 -968
rect 12127 -1008 12335 -1002
rect 12585 -968 12793 -962
rect 12585 -1002 12597 -968
rect 12781 -1002 12793 -968
rect 12585 -1008 12793 -1002
rect 8994 -1342 9054 -1008
rect 9448 -1076 9508 -1008
rect 9910 -1076 9970 -1008
rect 10364 -1076 10424 -1008
rect 10826 -1076 10886 -1008
rect 11280 -1076 11340 -1008
rect 11730 -1076 11790 -1008
rect 12196 -1076 12256 -1008
rect 12652 -1076 12712 -1008
rect 9448 -1080 10364 -1076
rect 9508 -1136 9910 -1080
rect 9448 -1146 9508 -1140
rect 9970 -1136 10364 -1080
rect 10424 -1136 10826 -1076
rect 10886 -1082 11730 -1076
rect 10886 -1136 11280 -1082
rect 9910 -1146 9970 -1140
rect 10364 -1142 10424 -1136
rect 10826 -1142 10886 -1136
rect 11340 -1136 11730 -1082
rect 11790 -1136 12196 -1076
rect 12256 -1080 12712 -1076
rect 12256 -1136 12652 -1080
rect 11730 -1142 11790 -1136
rect 12196 -1142 12256 -1136
rect 11280 -1148 11340 -1142
rect 12652 -1146 12712 -1140
rect 12886 -1202 12946 -909
rect 13344 -909 13359 -874
rect 13393 252 13406 267
rect 13766 267 13826 418
rect 13998 366 14058 418
rect 13921 360 14129 366
rect 13921 326 13933 360
rect 14117 326 14129 360
rect 13921 320 14129 326
rect 13393 -874 13399 252
rect 13766 246 13779 267
rect 13773 -874 13779 246
rect 13393 -909 13404 -874
rect 13043 -968 13251 -962
rect 13043 -1002 13055 -968
rect 13239 -1002 13251 -968
rect 13043 -1008 13251 -1002
rect 12880 -1262 12886 -1202
rect 12946 -1262 12952 -1202
rect 13116 -1342 13176 -1008
rect 13344 -1342 13404 -909
rect 13764 -909 13779 -874
rect 13813 246 13826 267
rect 14224 267 14284 418
rect 14450 436 17714 496
rect 14450 366 14510 436
rect 14912 366 14972 436
rect 15366 366 15426 436
rect 15828 366 15888 436
rect 16282 366 16342 436
rect 16732 366 16792 436
rect 17198 366 17258 436
rect 17654 366 17714 436
rect 18116 366 18176 628
rect 14379 360 14587 366
rect 14379 326 14391 360
rect 14575 326 14587 360
rect 14379 320 14587 326
rect 14837 360 15045 366
rect 14837 326 14849 360
rect 15033 326 15045 360
rect 14837 320 15045 326
rect 15295 360 15503 366
rect 15295 326 15307 360
rect 15491 326 15503 360
rect 15295 320 15503 326
rect 15753 360 15961 366
rect 15753 326 15765 360
rect 15949 326 15961 360
rect 15753 320 15961 326
rect 16211 360 16419 366
rect 16211 326 16223 360
rect 16407 326 16419 360
rect 16211 320 16419 326
rect 16669 360 16877 366
rect 16669 326 16681 360
rect 16865 326 16877 360
rect 16669 320 16877 326
rect 17127 360 17335 366
rect 17127 326 17139 360
rect 17323 326 17335 360
rect 17127 320 17335 326
rect 17585 360 17793 366
rect 17585 326 17597 360
rect 17781 326 17793 360
rect 17585 320 17793 326
rect 18043 360 18251 366
rect 18043 326 18055 360
rect 18239 326 18251 360
rect 18043 320 18251 326
rect 13813 -874 13819 246
rect 14224 224 14237 267
rect 14231 -868 14237 224
rect 13813 -909 13824 -874
rect 13764 -1342 13824 -909
rect 14222 -909 14237 -868
rect 14271 224 14284 267
rect 14689 267 14735 279
rect 14271 -868 14277 224
rect 14271 -909 14282 -868
rect 13921 -968 14129 -962
rect 13921 -1002 13933 -968
rect 14117 -1002 14129 -968
rect 13921 -1008 14129 -1002
rect 13992 -1342 14052 -1008
rect 14222 -1342 14282 -909
rect 14689 -909 14695 267
rect 14729 -909 14735 267
rect 14689 -921 14735 -909
rect 15147 267 15193 279
rect 15147 -909 15153 267
rect 15187 -909 15193 267
rect 15147 -921 15193 -909
rect 15605 267 15651 279
rect 15605 -909 15611 267
rect 15645 -909 15651 267
rect 15605 -921 15651 -909
rect 16063 267 16109 279
rect 16063 -909 16069 267
rect 16103 -909 16109 267
rect 16063 -921 16109 -909
rect 16521 267 16567 279
rect 16521 -909 16527 267
rect 16561 -909 16567 267
rect 16521 -921 16567 -909
rect 16979 267 17025 279
rect 16979 -909 16985 267
rect 17019 -909 17025 267
rect 16979 -921 17025 -909
rect 17437 267 17483 279
rect 17437 -909 17443 267
rect 17477 -909 17483 267
rect 17895 267 17941 279
rect 17895 -902 17901 267
rect 17437 -921 17483 -909
rect 17886 -909 17901 -902
rect 17935 -902 17941 267
rect 18342 267 18402 628
rect 18342 214 18359 267
rect 18353 -876 18359 214
rect 17935 -909 17946 -902
rect 14379 -968 14587 -962
rect 14379 -1002 14391 -968
rect 14575 -1002 14587 -968
rect 14379 -1008 14587 -1002
rect 14837 -968 15045 -962
rect 14837 -1002 14849 -968
rect 15033 -1002 15045 -968
rect 14837 -1008 15045 -1002
rect 15295 -968 15503 -962
rect 15295 -1002 15307 -968
rect 15491 -1002 15503 -968
rect 15295 -1008 15503 -1002
rect 15753 -968 15961 -962
rect 15753 -1002 15765 -968
rect 15949 -1002 15961 -968
rect 15753 -1008 15961 -1002
rect 16211 -968 16419 -962
rect 16211 -1002 16223 -968
rect 16407 -1002 16419 -968
rect 16211 -1008 16419 -1002
rect 16669 -968 16877 -962
rect 16669 -1002 16681 -968
rect 16865 -1002 16877 -968
rect 16669 -1008 16877 -1002
rect 17127 -968 17335 -962
rect 17127 -1002 17139 -968
rect 17323 -1002 17335 -968
rect 17127 -1008 17335 -1002
rect 17585 -968 17793 -962
rect 17585 -1002 17597 -968
rect 17781 -1002 17793 -968
rect 17585 -1008 17793 -1002
rect 14450 -1076 14510 -1008
rect 14912 -1072 14972 -1008
rect 14450 -1080 14912 -1076
rect 14510 -1132 14912 -1080
rect 15366 -1076 15426 -1008
rect 15828 -1076 15888 -1008
rect 16282 -1076 16342 -1008
rect 16732 -1072 16792 -1008
rect 14972 -1078 16732 -1076
rect 14972 -1132 15366 -1078
rect 14510 -1136 15366 -1132
rect 14912 -1138 14972 -1136
rect 15426 -1136 15828 -1078
rect 14450 -1146 14510 -1140
rect 15366 -1144 15426 -1138
rect 15888 -1136 16282 -1078
rect 15828 -1144 15888 -1138
rect 16342 -1132 16732 -1078
rect 17198 -1076 17258 -1008
rect 17654 -1076 17714 -1008
rect 16792 -1078 17714 -1076
rect 16792 -1132 17198 -1078
rect 16342 -1136 17198 -1132
rect 16732 -1138 16792 -1136
rect 17258 -1136 17654 -1078
rect 16282 -1144 16342 -1138
rect 17198 -1144 17258 -1138
rect 17654 -1144 17714 -1138
rect 17886 -1208 17946 -909
rect 18344 -909 18359 -876
rect 18393 214 18402 267
rect 18393 -876 18399 214
rect 18393 -909 18404 -876
rect 18043 -968 18251 -962
rect 18043 -1002 18055 -968
rect 18239 -1002 18251 -968
rect 18043 -1008 18251 -1002
rect 17886 -1274 17946 -1268
rect 18116 -1342 18176 -1008
rect 18344 -1342 18404 -909
rect 18690 -1166 18696 628
rect 18796 -1166 18802 4006
rect 22768 760 22828 8708
rect 28038 8702 28098 8708
rect 29040 8704 29100 8708
rect 30745 8739 30803 8745
rect 29040 8698 29200 8704
rect 29040 8650 29140 8698
rect 29188 8650 29200 8698
rect 29040 8644 29200 8650
rect 29234 8700 29442 8706
rect 29234 8652 29246 8700
rect 29294 8652 29382 8700
rect 29430 8652 29442 8700
rect 29234 8646 29442 8652
rect 29726 8700 30640 8706
rect 29726 8652 29738 8700
rect 29786 8652 30580 8700
rect 30628 8652 30640 8700
rect 30745 8705 30757 8739
rect 30791 8736 30803 8739
rect 30983 8739 31041 8745
rect 30983 8736 30995 8739
rect 30791 8708 30995 8736
rect 30791 8705 30803 8708
rect 30745 8699 30803 8705
rect 30983 8705 30995 8708
rect 31029 8736 31041 8739
rect 31487 8739 31545 8745
rect 31487 8736 31499 8739
rect 31029 8708 31499 8736
rect 31029 8705 31041 8708
rect 30983 8699 31041 8705
rect 31487 8705 31499 8708
rect 31533 8705 31545 8739
rect 31487 8699 31545 8705
rect 32230 8680 32418 8686
rect 29726 8646 30640 8652
rect 30826 8648 30886 8654
rect 23080 8624 23140 8630
rect 22934 6004 22940 6064
rect 23000 6004 23006 6064
rect 22940 3164 23000 6004
rect 22940 3158 23002 3164
rect 22940 3098 22942 3158
rect 22940 3092 23002 3098
rect 22762 700 22768 760
rect 22828 700 22834 760
rect 18690 -1342 18802 -1166
rect 8346 -1348 18802 -1342
rect 8346 -1448 8452 -1348
rect 18696 -1448 18802 -1348
rect 8346 -1454 18802 -1448
rect 8346 -1684 18802 -1678
rect 8346 -1784 8452 -1684
rect 18696 -1784 18802 -1684
rect 8346 -1790 18802 -1784
rect 8346 -1914 8458 -1790
rect 8346 -3918 8352 -1914
rect 8452 -3918 8458 -1914
rect 8766 -2226 8826 -1790
rect 8996 -2136 9056 -1790
rect 12886 -1882 12946 -1876
rect 9454 -2016 9910 -2010
rect 9442 -2076 9448 -2016
rect 9508 -2070 9910 -2016
rect 9970 -2016 10826 -2010
rect 9970 -2070 10364 -2016
rect 9508 -2076 9514 -2070
rect 9448 -2136 9514 -2076
rect 9910 -2136 9976 -2070
rect 10358 -2076 10364 -2070
rect 10424 -2070 10826 -2016
rect 10886 -2070 11280 -2010
rect 11340 -2070 11730 -2010
rect 11790 -2016 12652 -2010
rect 11790 -2070 12196 -2016
rect 10424 -2076 10430 -2070
rect 10364 -2136 10430 -2076
rect 10826 -2136 10892 -2070
rect 11280 -2136 11346 -2070
rect 11730 -2136 11796 -2070
rect 12190 -2076 12196 -2070
rect 12256 -2070 12652 -2016
rect 12712 -2070 12718 -2010
rect 12256 -2076 12262 -2070
rect 12196 -2136 12262 -2076
rect 12652 -2136 12718 -2070
rect 8920 -2142 9128 -2136
rect 8920 -2176 8932 -2142
rect 9116 -2176 9128 -2142
rect 8920 -2182 9128 -2176
rect 9378 -2142 9586 -2136
rect 9378 -2176 9390 -2142
rect 9574 -2176 9586 -2142
rect 9378 -2182 9586 -2176
rect 9836 -2142 10044 -2136
rect 9836 -2176 9848 -2142
rect 10032 -2176 10044 -2142
rect 9836 -2182 10044 -2176
rect 10294 -2142 10502 -2136
rect 10294 -2176 10306 -2142
rect 10490 -2176 10502 -2142
rect 10294 -2182 10502 -2176
rect 10752 -2142 10960 -2136
rect 10752 -2176 10764 -2142
rect 10948 -2176 10960 -2142
rect 10752 -2182 10960 -2176
rect 11210 -2142 11418 -2136
rect 11210 -2176 11222 -2142
rect 11406 -2176 11418 -2142
rect 11210 -2182 11418 -2176
rect 11668 -2142 11876 -2136
rect 11668 -2176 11680 -2142
rect 11864 -2176 11876 -2142
rect 11668 -2182 11876 -2176
rect 12126 -2142 12334 -2136
rect 12126 -2176 12138 -2142
rect 12322 -2176 12334 -2142
rect 12126 -2182 12334 -2176
rect 12584 -2142 12792 -2136
rect 12584 -2176 12596 -2142
rect 12780 -2176 12792 -2142
rect 12584 -2182 12792 -2176
rect 8766 -2266 8778 -2226
rect 8772 -2362 8778 -2266
rect 8766 -2402 8778 -2362
rect 8812 -2266 8826 -2226
rect 9230 -2226 9276 -2214
rect 8812 -2362 8818 -2266
rect 9230 -2360 9236 -2226
rect 8812 -2402 8826 -2362
rect 8766 -2618 8826 -2402
rect 9222 -2402 9236 -2360
rect 9270 -2360 9276 -2226
rect 9688 -2226 9734 -2214
rect 9270 -2402 9282 -2360
rect 8920 -2452 9128 -2446
rect 8920 -2486 8932 -2452
rect 9116 -2486 9128 -2452
rect 8920 -2492 9128 -2486
rect 8994 -2618 9054 -2492
rect 8766 -2678 9054 -2618
rect 8766 -2894 8826 -2678
rect 8994 -2804 9054 -2678
rect 8920 -2810 9128 -2804
rect 8920 -2844 8932 -2810
rect 9116 -2844 9128 -2810
rect 8920 -2850 9128 -2844
rect 8766 -2914 8778 -2894
rect 8772 -3040 8778 -2914
rect 8758 -3070 8778 -3040
rect 8812 -2914 8826 -2894
rect 9222 -2894 9282 -2402
rect 9688 -2402 9694 -2226
rect 9728 -2402 9734 -2226
rect 9688 -2414 9734 -2402
rect 10146 -2226 10192 -2214
rect 10146 -2402 10152 -2226
rect 10186 -2402 10192 -2226
rect 10146 -2414 10192 -2402
rect 10604 -2226 10650 -2214
rect 10604 -2402 10610 -2226
rect 10644 -2402 10650 -2226
rect 10604 -2414 10650 -2402
rect 11062 -2226 11108 -2214
rect 11062 -2402 11068 -2226
rect 11102 -2402 11108 -2226
rect 11062 -2414 11108 -2402
rect 11520 -2226 11566 -2214
rect 11520 -2402 11526 -2226
rect 11560 -2402 11566 -2226
rect 11520 -2414 11566 -2402
rect 11978 -2226 12024 -2214
rect 11978 -2402 11984 -2226
rect 12018 -2402 12024 -2226
rect 11978 -2414 12024 -2402
rect 12436 -2226 12482 -2214
rect 12436 -2402 12442 -2226
rect 12476 -2402 12482 -2226
rect 12886 -2226 12946 -1942
rect 13114 -2136 13174 -1790
rect 13042 -2142 13250 -2136
rect 13042 -2176 13054 -2142
rect 13238 -2176 13250 -2142
rect 13042 -2182 13250 -2176
rect 12886 -2256 12900 -2226
rect 12436 -2414 12482 -2402
rect 12894 -2402 12900 -2256
rect 12934 -2256 12946 -2226
rect 13346 -2226 13406 -1790
rect 13346 -2254 13358 -2226
rect 12934 -2402 12940 -2256
rect 13352 -2346 13358 -2254
rect 12894 -2414 12940 -2402
rect 13346 -2402 13358 -2346
rect 13392 -2254 13406 -2226
rect 13766 -2226 13826 -1790
rect 14000 -2136 14060 -1790
rect 13920 -2142 14128 -2136
rect 13920 -2176 13932 -2142
rect 14116 -2176 14128 -2142
rect 13920 -2182 14128 -2176
rect 13392 -2346 13398 -2254
rect 13766 -2262 13778 -2226
rect 13392 -2402 13406 -2346
rect 13772 -2366 13778 -2262
rect 9378 -2452 9586 -2446
rect 9378 -2486 9390 -2452
rect 9574 -2486 9586 -2452
rect 9378 -2492 9586 -2486
rect 9836 -2452 10044 -2446
rect 9836 -2486 9848 -2452
rect 10032 -2486 10044 -2452
rect 9836 -2492 10044 -2486
rect 10294 -2452 10502 -2446
rect 10294 -2486 10306 -2452
rect 10490 -2486 10502 -2452
rect 10294 -2492 10502 -2486
rect 10752 -2452 10960 -2446
rect 10752 -2486 10764 -2452
rect 10948 -2486 10960 -2452
rect 10752 -2492 10960 -2486
rect 11210 -2452 11418 -2446
rect 11210 -2486 11222 -2452
rect 11406 -2486 11418 -2452
rect 11210 -2492 11418 -2486
rect 11668 -2452 11876 -2446
rect 11668 -2486 11680 -2452
rect 11864 -2486 11876 -2452
rect 11668 -2492 11876 -2486
rect 12126 -2452 12334 -2446
rect 12126 -2486 12138 -2452
rect 12322 -2486 12334 -2452
rect 12126 -2492 12334 -2486
rect 12584 -2452 12792 -2446
rect 12584 -2486 12596 -2452
rect 12780 -2486 12792 -2452
rect 12584 -2492 12792 -2486
rect 13042 -2452 13250 -2446
rect 13042 -2486 13054 -2452
rect 13238 -2486 13250 -2452
rect 13042 -2492 13250 -2486
rect 9448 -2558 9508 -2492
rect 9910 -2558 9970 -2492
rect 10364 -2558 10424 -2492
rect 10826 -2558 10886 -2492
rect 11280 -2558 11340 -2492
rect 11730 -2558 11790 -2492
rect 12196 -2558 12256 -2492
rect 12652 -2558 12712 -2492
rect 9448 -2618 12712 -2558
rect 9454 -2738 12718 -2678
rect 9454 -2804 9514 -2738
rect 9916 -2804 9976 -2738
rect 10370 -2804 10430 -2738
rect 10832 -2804 10892 -2738
rect 11286 -2804 11346 -2738
rect 11736 -2804 11796 -2738
rect 12202 -2804 12262 -2738
rect 12658 -2804 12718 -2738
rect 13114 -2804 13174 -2492
rect 9378 -2810 9586 -2804
rect 9378 -2844 9390 -2810
rect 9574 -2844 9586 -2810
rect 9378 -2850 9586 -2844
rect 9836 -2810 10044 -2804
rect 9836 -2844 9848 -2810
rect 10032 -2844 10044 -2810
rect 9836 -2850 10044 -2844
rect 10294 -2810 10502 -2804
rect 10294 -2844 10306 -2810
rect 10490 -2844 10502 -2810
rect 10294 -2850 10502 -2844
rect 10752 -2810 10960 -2804
rect 10752 -2844 10764 -2810
rect 10948 -2844 10960 -2810
rect 10752 -2850 10960 -2844
rect 11210 -2810 11418 -2804
rect 11210 -2844 11222 -2810
rect 11406 -2844 11418 -2810
rect 11210 -2850 11418 -2844
rect 11668 -2810 11876 -2804
rect 11668 -2844 11680 -2810
rect 11864 -2844 11876 -2810
rect 11668 -2850 11876 -2844
rect 12126 -2810 12334 -2804
rect 12126 -2844 12138 -2810
rect 12322 -2844 12334 -2810
rect 12126 -2850 12334 -2844
rect 12584 -2810 12792 -2804
rect 12584 -2844 12596 -2810
rect 12780 -2844 12792 -2810
rect 12584 -2850 12792 -2844
rect 13042 -2810 13250 -2804
rect 13042 -2844 13054 -2810
rect 13238 -2844 13250 -2810
rect 13042 -2850 13250 -2844
rect 8812 -3070 8818 -2914
rect 9222 -2922 9236 -2894
rect 8758 -3450 8818 -3070
rect 9230 -3070 9236 -2922
rect 9270 -2922 9282 -2894
rect 9688 -2894 9734 -2882
rect 9270 -3070 9276 -2922
rect 9230 -3082 9276 -3070
rect 9688 -3070 9694 -2894
rect 9728 -3070 9734 -2894
rect 9688 -3082 9734 -3070
rect 10146 -2894 10192 -2882
rect 10146 -3070 10152 -2894
rect 10186 -3070 10192 -2894
rect 10146 -3082 10192 -3070
rect 10604 -2894 10650 -2882
rect 10604 -3070 10610 -2894
rect 10644 -3070 10650 -2894
rect 10604 -3082 10650 -3070
rect 11062 -2894 11108 -2882
rect 11062 -3070 11068 -2894
rect 11102 -3070 11108 -2894
rect 11062 -3082 11108 -3070
rect 11520 -2894 11566 -2882
rect 11520 -3070 11526 -2894
rect 11560 -3070 11566 -2894
rect 11520 -3082 11566 -3070
rect 11978 -2894 12024 -2882
rect 11978 -3070 11984 -2894
rect 12018 -3070 12024 -2894
rect 11978 -3082 12024 -3070
rect 12436 -2894 12482 -2882
rect 12436 -3070 12442 -2894
rect 12476 -3070 12482 -2894
rect 12894 -2894 12940 -2882
rect 12894 -3042 12900 -2894
rect 12436 -3082 12482 -3070
rect 12886 -3070 12900 -3042
rect 12934 -3042 12940 -2894
rect 13346 -2894 13406 -2402
rect 12934 -3070 12946 -3042
rect 8920 -3120 9128 -3114
rect 8920 -3154 8932 -3120
rect 9116 -3154 9128 -3120
rect 8920 -3160 9128 -3154
rect 9378 -3120 9586 -3114
rect 9378 -3154 9390 -3120
rect 9574 -3154 9586 -3120
rect 9378 -3160 9586 -3154
rect 9836 -3120 10044 -3114
rect 9836 -3154 9848 -3120
rect 10032 -3154 10044 -3120
rect 9836 -3160 10044 -3154
rect 10294 -3120 10502 -3114
rect 10294 -3154 10306 -3120
rect 10490 -3154 10502 -3120
rect 10294 -3160 10502 -3154
rect 10752 -3120 10960 -3114
rect 10752 -3154 10764 -3120
rect 10948 -3154 10960 -3120
rect 10752 -3160 10960 -3154
rect 11210 -3120 11418 -3114
rect 11210 -3154 11222 -3120
rect 11406 -3154 11418 -3120
rect 11210 -3160 11418 -3154
rect 11668 -3120 11876 -3114
rect 11668 -3154 11680 -3120
rect 11864 -3154 11876 -3120
rect 11668 -3160 11876 -3154
rect 12126 -3120 12334 -3114
rect 12126 -3154 12138 -3120
rect 12322 -3154 12334 -3120
rect 12126 -3160 12334 -3154
rect 12584 -3120 12792 -3114
rect 12584 -3154 12596 -3120
rect 12780 -3154 12792 -3120
rect 12584 -3160 12792 -3154
rect 8998 -3450 9058 -3160
rect 9448 -3226 9508 -3160
rect 9910 -3226 9970 -3160
rect 10364 -3226 10424 -3160
rect 10826 -3226 10886 -3160
rect 11280 -3226 11340 -3160
rect 11730 -3226 11790 -3160
rect 12196 -3226 12256 -3160
rect 12652 -3226 12712 -3160
rect 9448 -3286 12650 -3226
rect 12710 -3286 12716 -3226
rect 12886 -3450 12946 -3070
rect 13346 -3070 13358 -2894
rect 13392 -3070 13406 -2894
rect 13042 -3120 13250 -3114
rect 13042 -3154 13054 -3120
rect 13238 -3154 13250 -3120
rect 13042 -3160 13250 -3154
rect 13112 -3450 13172 -3160
rect 13346 -3450 13406 -3070
rect 13762 -2402 13778 -2366
rect 13812 -2262 13826 -2226
rect 14222 -2226 14282 -1790
rect 17880 -1930 17886 -1870
rect 17946 -1930 17952 -1870
rect 16726 -2010 16732 -2006
rect 14444 -2070 14450 -2010
rect 14510 -2012 16732 -2010
rect 14510 -2070 14912 -2012
rect 14450 -2136 14514 -2070
rect 14906 -2072 14912 -2070
rect 14972 -2070 15366 -2012
rect 14972 -2072 14978 -2070
rect 15360 -2072 15366 -2070
rect 15426 -2070 15828 -2012
rect 15426 -2072 15432 -2070
rect 15822 -2072 15828 -2070
rect 15888 -2070 16282 -2012
rect 15888 -2072 15894 -2070
rect 16276 -2072 16282 -2070
rect 16342 -2066 16732 -2012
rect 16792 -2010 16798 -2006
rect 16792 -2066 17198 -2010
rect 16342 -2070 17198 -2066
rect 17258 -2070 17654 -2010
rect 17714 -2070 17720 -2010
rect 16342 -2072 16348 -2070
rect 14912 -2136 14976 -2072
rect 15366 -2136 15430 -2072
rect 15828 -2136 15892 -2072
rect 16282 -2136 16346 -2072
rect 16732 -2136 16796 -2070
rect 17198 -2136 17262 -2070
rect 17654 -2136 17718 -2070
rect 14378 -2142 14586 -2136
rect 14378 -2176 14390 -2142
rect 14574 -2176 14586 -2142
rect 14378 -2182 14586 -2176
rect 14836 -2142 15044 -2136
rect 14836 -2176 14848 -2142
rect 15032 -2176 15044 -2142
rect 14836 -2182 15044 -2176
rect 15294 -2142 15502 -2136
rect 15294 -2176 15306 -2142
rect 15490 -2176 15502 -2142
rect 15294 -2182 15502 -2176
rect 15752 -2142 15960 -2136
rect 15752 -2176 15764 -2142
rect 15948 -2176 15960 -2142
rect 15752 -2182 15960 -2176
rect 16210 -2142 16418 -2136
rect 16210 -2176 16222 -2142
rect 16406 -2176 16418 -2142
rect 16210 -2182 16418 -2176
rect 16668 -2142 16876 -2136
rect 16668 -2176 16680 -2142
rect 16864 -2176 16876 -2142
rect 16668 -2182 16876 -2176
rect 17126 -2142 17334 -2136
rect 17126 -2176 17138 -2142
rect 17322 -2176 17334 -2142
rect 17126 -2182 17334 -2176
rect 17584 -2142 17792 -2136
rect 17584 -2176 17596 -2142
rect 17780 -2176 17792 -2142
rect 17584 -2182 17792 -2176
rect 13812 -2366 13818 -2262
rect 14222 -2290 14236 -2226
rect 14230 -2358 14236 -2290
rect 13812 -2402 13822 -2366
rect 13762 -2556 13822 -2402
rect 14222 -2402 14236 -2358
rect 14270 -2290 14282 -2226
rect 14688 -2226 14734 -2214
rect 14270 -2358 14276 -2290
rect 14270 -2402 14282 -2358
rect 13920 -2452 14128 -2446
rect 13920 -2486 13932 -2452
rect 14116 -2486 14128 -2452
rect 13920 -2492 14128 -2486
rect 13990 -2556 14050 -2492
rect 14222 -2556 14282 -2402
rect 14688 -2402 14694 -2226
rect 14728 -2402 14734 -2226
rect 14688 -2414 14734 -2402
rect 15146 -2226 15192 -2214
rect 15146 -2402 15152 -2226
rect 15186 -2402 15192 -2226
rect 15146 -2414 15192 -2402
rect 15604 -2226 15650 -2214
rect 15604 -2402 15610 -2226
rect 15644 -2402 15650 -2226
rect 15604 -2414 15650 -2402
rect 16062 -2226 16108 -2214
rect 16062 -2402 16068 -2226
rect 16102 -2402 16108 -2226
rect 16062 -2414 16108 -2402
rect 16520 -2226 16566 -2214
rect 16520 -2402 16526 -2226
rect 16560 -2402 16566 -2226
rect 16520 -2414 16566 -2402
rect 16978 -2226 17024 -2214
rect 16978 -2402 16984 -2226
rect 17018 -2402 17024 -2226
rect 16978 -2414 17024 -2402
rect 17436 -2226 17482 -2214
rect 17436 -2402 17442 -2226
rect 17476 -2402 17482 -2226
rect 17886 -2226 17946 -1930
rect 18126 -2136 18186 -1790
rect 18042 -2142 18250 -2136
rect 18042 -2176 18054 -2142
rect 18238 -2176 18250 -2142
rect 18042 -2182 18250 -2176
rect 17886 -2268 17900 -2226
rect 17436 -2414 17482 -2402
rect 17894 -2402 17900 -2268
rect 17934 -2268 17946 -2226
rect 18344 -2226 18404 -1790
rect 18344 -2266 18358 -2226
rect 17934 -2402 17940 -2268
rect 18352 -2356 18358 -2266
rect 17894 -2414 17940 -2402
rect 18342 -2402 18358 -2356
rect 18392 -2266 18404 -2226
rect 18690 -1914 18802 -1790
rect 18392 -2356 18398 -2266
rect 18392 -2402 18402 -2356
rect 14378 -2452 14586 -2446
rect 14378 -2486 14390 -2452
rect 14574 -2486 14586 -2452
rect 14378 -2492 14586 -2486
rect 14836 -2452 15044 -2446
rect 14836 -2486 14848 -2452
rect 15032 -2486 15044 -2452
rect 14836 -2492 15044 -2486
rect 15294 -2452 15502 -2446
rect 15294 -2486 15306 -2452
rect 15490 -2486 15502 -2452
rect 15294 -2492 15502 -2486
rect 15752 -2452 15960 -2446
rect 15752 -2486 15764 -2452
rect 15948 -2486 15960 -2452
rect 15752 -2492 15960 -2486
rect 16210 -2452 16418 -2446
rect 16210 -2486 16222 -2452
rect 16406 -2486 16418 -2452
rect 16210 -2492 16418 -2486
rect 16668 -2452 16876 -2446
rect 16668 -2486 16680 -2452
rect 16864 -2486 16876 -2452
rect 16668 -2492 16876 -2486
rect 17126 -2452 17334 -2446
rect 17126 -2486 17138 -2452
rect 17322 -2486 17334 -2452
rect 17126 -2492 17334 -2486
rect 17584 -2452 17792 -2446
rect 17584 -2486 17596 -2452
rect 17780 -2486 17792 -2452
rect 17584 -2492 17792 -2486
rect 18042 -2452 18250 -2446
rect 18042 -2486 18054 -2452
rect 18238 -2486 18250 -2452
rect 18042 -2492 18250 -2486
rect 13762 -2616 14282 -2556
rect 13762 -3450 13822 -2616
rect 13990 -3450 14050 -2616
rect 14222 -3450 14282 -2616
rect 14448 -2558 14508 -2492
rect 14910 -2558 14970 -2492
rect 15364 -2558 15424 -2492
rect 15826 -2558 15886 -2492
rect 16280 -2558 16340 -2492
rect 16730 -2558 16790 -2492
rect 17196 -2558 17256 -2492
rect 17652 -2558 17712 -2492
rect 14448 -2618 17712 -2558
rect 18116 -3450 18176 -2492
rect 18342 -3450 18402 -2402
rect 8694 -3478 18464 -3450
rect 8694 -3564 8744 -3478
rect 8840 -3564 9324 -3478
rect 9420 -3564 9924 -3478
rect 10020 -3564 10524 -3478
rect 10620 -3564 11124 -3478
rect 11220 -3564 11724 -3478
rect 11820 -3564 12324 -3478
rect 12420 -3564 12924 -3478
rect 13020 -3564 13524 -3478
rect 13620 -3564 14124 -3478
rect 14220 -3564 14724 -3478
rect 14820 -3564 15324 -3478
rect 15420 -3564 15924 -3478
rect 16020 -3564 16524 -3478
rect 16620 -3564 17124 -3478
rect 17220 -3564 17724 -3478
rect 17820 -3564 18324 -3478
rect 18420 -3564 18464 -3478
rect 8694 -3594 18464 -3564
rect 8346 -4042 8458 -3918
rect 9058 -4042 9068 -3742
rect 18080 -4042 18090 -3742
rect 18690 -3918 18696 -1914
rect 18796 -3918 18802 -1914
rect 18690 -4042 18802 -3918
rect 8346 -4048 18802 -4042
rect 8346 -4148 8452 -4048
rect 18696 -4148 18802 -4048
rect 8346 -4154 18802 -4148
rect 12300 -4608 22756 -4602
rect 12300 -4708 12406 -4608
rect 22650 -4708 22756 -4608
rect 12300 -4714 22756 -4708
rect 12300 -4838 12412 -4714
rect 12300 -6842 12306 -4838
rect 12406 -6842 12412 -4838
rect 13012 -5014 13022 -4714
rect 22034 -5014 22044 -4714
rect 22644 -4838 22756 -4714
rect 12638 -5192 22408 -5162
rect 12638 -5278 12682 -5192
rect 12778 -5278 13282 -5192
rect 13378 -5278 13882 -5192
rect 13978 -5278 14482 -5192
rect 14578 -5278 15082 -5192
rect 15178 -5278 15682 -5192
rect 15778 -5278 16282 -5192
rect 16378 -5278 16882 -5192
rect 16978 -5278 17482 -5192
rect 17578 -5278 18082 -5192
rect 18178 -5278 18682 -5192
rect 18778 -5278 19282 -5192
rect 19378 -5278 19882 -5192
rect 19978 -5278 20482 -5192
rect 20578 -5278 21082 -5192
rect 21178 -5278 21682 -5192
rect 21778 -5278 22262 -5192
rect 22358 -5278 22408 -5192
rect 12638 -5306 22408 -5278
rect 12700 -6354 12760 -5306
rect 12926 -6264 12986 -5306
rect 13390 -6198 16654 -6138
rect 13390 -6264 13450 -6198
rect 13846 -6264 13906 -6198
rect 14312 -6264 14372 -6198
rect 14762 -6264 14822 -6198
rect 15216 -6264 15276 -6198
rect 15678 -6264 15738 -6198
rect 16132 -6264 16192 -6198
rect 16594 -6264 16654 -6198
rect 16820 -6140 16880 -5306
rect 17052 -6140 17112 -5306
rect 17280 -6140 17340 -5306
rect 16820 -6200 17340 -6140
rect 12852 -6270 13060 -6264
rect 12852 -6304 12864 -6270
rect 13048 -6304 13060 -6270
rect 12852 -6310 13060 -6304
rect 13310 -6270 13518 -6264
rect 13310 -6304 13322 -6270
rect 13506 -6304 13518 -6270
rect 13310 -6310 13518 -6304
rect 13768 -6270 13976 -6264
rect 13768 -6304 13780 -6270
rect 13964 -6304 13976 -6270
rect 13768 -6310 13976 -6304
rect 14226 -6270 14434 -6264
rect 14226 -6304 14238 -6270
rect 14422 -6304 14434 -6270
rect 14226 -6310 14434 -6304
rect 14684 -6270 14892 -6264
rect 14684 -6304 14696 -6270
rect 14880 -6304 14892 -6270
rect 14684 -6310 14892 -6304
rect 15142 -6270 15350 -6264
rect 15142 -6304 15154 -6270
rect 15338 -6304 15350 -6270
rect 15142 -6310 15350 -6304
rect 15600 -6270 15808 -6264
rect 15600 -6304 15612 -6270
rect 15796 -6304 15808 -6270
rect 15600 -6310 15808 -6304
rect 16058 -6270 16266 -6264
rect 16058 -6304 16070 -6270
rect 16254 -6304 16266 -6270
rect 16058 -6310 16266 -6304
rect 16516 -6270 16724 -6264
rect 16516 -6304 16528 -6270
rect 16712 -6304 16724 -6270
rect 16516 -6310 16724 -6304
rect 12700 -6400 12710 -6354
rect 12704 -6490 12710 -6400
rect 12300 -6966 12412 -6842
rect 12698 -6530 12710 -6490
rect 12744 -6400 12760 -6354
rect 13162 -6354 13208 -6342
rect 12744 -6490 12750 -6400
rect 13162 -6488 13168 -6354
rect 12744 -6530 12758 -6490
rect 12698 -6966 12758 -6530
rect 13156 -6530 13168 -6488
rect 13202 -6488 13208 -6354
rect 13620 -6354 13666 -6342
rect 13202 -6530 13216 -6488
rect 12852 -6580 13060 -6574
rect 12852 -6614 12864 -6580
rect 13048 -6614 13060 -6580
rect 12852 -6620 13060 -6614
rect 12916 -6966 12976 -6620
rect 13156 -6826 13216 -6530
rect 13620 -6530 13626 -6354
rect 13660 -6530 13666 -6354
rect 13620 -6542 13666 -6530
rect 14078 -6354 14124 -6342
rect 14078 -6530 14084 -6354
rect 14118 -6530 14124 -6354
rect 14078 -6542 14124 -6530
rect 14536 -6354 14582 -6342
rect 14536 -6530 14542 -6354
rect 14576 -6530 14582 -6354
rect 14536 -6542 14582 -6530
rect 14994 -6354 15040 -6342
rect 14994 -6530 15000 -6354
rect 15034 -6530 15040 -6354
rect 14994 -6542 15040 -6530
rect 15452 -6354 15498 -6342
rect 15452 -6530 15458 -6354
rect 15492 -6530 15498 -6354
rect 15452 -6542 15498 -6530
rect 15910 -6354 15956 -6342
rect 15910 -6530 15916 -6354
rect 15950 -6530 15956 -6354
rect 15910 -6542 15956 -6530
rect 16368 -6354 16414 -6342
rect 16368 -6530 16374 -6354
rect 16408 -6530 16414 -6354
rect 16820 -6354 16880 -6200
rect 17052 -6264 17112 -6200
rect 16974 -6270 17182 -6264
rect 16974 -6304 16986 -6270
rect 17170 -6304 17182 -6270
rect 16974 -6310 17182 -6304
rect 16820 -6398 16832 -6354
rect 16826 -6466 16832 -6398
rect 16368 -6542 16414 -6530
rect 16820 -6530 16832 -6466
rect 16866 -6398 16880 -6354
rect 17280 -6354 17340 -6200
rect 17280 -6390 17290 -6354
rect 16866 -6466 16872 -6398
rect 16866 -6530 16880 -6466
rect 17284 -6494 17290 -6390
rect 13310 -6580 13518 -6574
rect 13310 -6614 13322 -6580
rect 13506 -6614 13518 -6580
rect 13310 -6620 13518 -6614
rect 13768 -6580 13976 -6574
rect 13768 -6614 13780 -6580
rect 13964 -6614 13976 -6580
rect 13768 -6620 13976 -6614
rect 14226 -6580 14434 -6574
rect 14226 -6614 14238 -6580
rect 14422 -6614 14434 -6580
rect 14226 -6620 14434 -6614
rect 14684 -6580 14892 -6574
rect 14684 -6614 14696 -6580
rect 14880 -6614 14892 -6580
rect 14684 -6620 14892 -6614
rect 15142 -6580 15350 -6574
rect 15142 -6614 15154 -6580
rect 15338 -6614 15350 -6580
rect 15142 -6620 15350 -6614
rect 15600 -6580 15808 -6574
rect 15600 -6614 15612 -6580
rect 15796 -6614 15808 -6580
rect 15600 -6620 15808 -6614
rect 16058 -6580 16266 -6574
rect 16058 -6614 16070 -6580
rect 16254 -6614 16266 -6580
rect 16058 -6620 16266 -6614
rect 16516 -6580 16724 -6574
rect 16516 -6614 16528 -6580
rect 16712 -6614 16724 -6580
rect 16516 -6620 16724 -6614
rect 13384 -6686 13448 -6620
rect 13840 -6686 13904 -6620
rect 14306 -6686 14370 -6620
rect 14756 -6684 14820 -6620
rect 15210 -6684 15274 -6620
rect 15672 -6684 15736 -6620
rect 16126 -6684 16190 -6620
rect 14754 -6686 14760 -6684
rect 13382 -6746 13388 -6686
rect 13448 -6746 13844 -6686
rect 13904 -6690 14760 -6686
rect 13904 -6746 14310 -6690
rect 14304 -6750 14310 -6746
rect 14370 -6744 14760 -6690
rect 14820 -6686 14826 -6684
rect 15208 -6686 15214 -6684
rect 14820 -6744 15214 -6686
rect 15274 -6686 15280 -6684
rect 15670 -6686 15676 -6684
rect 15274 -6744 15676 -6686
rect 15736 -6686 15742 -6684
rect 16124 -6686 16130 -6684
rect 15736 -6744 16130 -6686
rect 16190 -6686 16196 -6684
rect 16588 -6686 16652 -6620
rect 16190 -6744 16592 -6686
rect 14370 -6746 16592 -6744
rect 16652 -6746 16658 -6686
rect 14370 -6750 14376 -6746
rect 13150 -6886 13156 -6826
rect 13216 -6886 13222 -6826
rect 16820 -6966 16880 -6530
rect 17276 -6530 17290 -6494
rect 17324 -6390 17340 -6354
rect 17696 -5686 17756 -5306
rect 17930 -5596 17990 -5306
rect 17852 -5602 18060 -5596
rect 17852 -5636 17864 -5602
rect 18048 -5636 18060 -5602
rect 17852 -5642 18060 -5636
rect 17696 -5862 17710 -5686
rect 17744 -5862 17756 -5686
rect 18156 -5686 18216 -5306
rect 18390 -5530 21596 -5470
rect 21656 -5530 21662 -5470
rect 18390 -5596 18450 -5530
rect 18846 -5596 18906 -5530
rect 19312 -5596 19372 -5530
rect 19762 -5596 19822 -5530
rect 20216 -5596 20276 -5530
rect 20678 -5596 20738 -5530
rect 21132 -5596 21192 -5530
rect 21594 -5596 21654 -5530
rect 22044 -5596 22104 -5306
rect 18310 -5602 18518 -5596
rect 18310 -5636 18322 -5602
rect 18506 -5636 18518 -5602
rect 18310 -5642 18518 -5636
rect 18768 -5602 18976 -5596
rect 18768 -5636 18780 -5602
rect 18964 -5636 18976 -5602
rect 18768 -5642 18976 -5636
rect 19226 -5602 19434 -5596
rect 19226 -5636 19238 -5602
rect 19422 -5636 19434 -5602
rect 19226 -5642 19434 -5636
rect 19684 -5602 19892 -5596
rect 19684 -5636 19696 -5602
rect 19880 -5636 19892 -5602
rect 19684 -5642 19892 -5636
rect 20142 -5602 20350 -5596
rect 20142 -5636 20154 -5602
rect 20338 -5636 20350 -5602
rect 20142 -5642 20350 -5636
rect 20600 -5602 20808 -5596
rect 20600 -5636 20612 -5602
rect 20796 -5636 20808 -5602
rect 20600 -5642 20808 -5636
rect 21058 -5602 21266 -5596
rect 21058 -5636 21070 -5602
rect 21254 -5636 21266 -5602
rect 21058 -5642 21266 -5636
rect 21516 -5602 21724 -5596
rect 21516 -5636 21528 -5602
rect 21712 -5636 21724 -5602
rect 21516 -5642 21724 -5636
rect 21974 -5602 22182 -5596
rect 21974 -5636 21986 -5602
rect 22170 -5636 22182 -5602
rect 21974 -5642 22182 -5636
rect 18156 -5714 18168 -5686
rect 17696 -6354 17756 -5862
rect 18162 -5862 18168 -5714
rect 18202 -5714 18216 -5686
rect 18620 -5686 18666 -5674
rect 18202 -5862 18208 -5714
rect 18162 -5874 18208 -5862
rect 18620 -5862 18626 -5686
rect 18660 -5862 18666 -5686
rect 18620 -5874 18666 -5862
rect 19078 -5686 19124 -5674
rect 19078 -5862 19084 -5686
rect 19118 -5862 19124 -5686
rect 19078 -5874 19124 -5862
rect 19536 -5686 19582 -5674
rect 19536 -5862 19542 -5686
rect 19576 -5862 19582 -5686
rect 19536 -5874 19582 -5862
rect 19994 -5686 20040 -5674
rect 19994 -5862 20000 -5686
rect 20034 -5862 20040 -5686
rect 19994 -5874 20040 -5862
rect 20452 -5686 20498 -5674
rect 20452 -5862 20458 -5686
rect 20492 -5862 20498 -5686
rect 20452 -5874 20498 -5862
rect 20910 -5686 20956 -5674
rect 20910 -5862 20916 -5686
rect 20950 -5862 20956 -5686
rect 20910 -5874 20956 -5862
rect 21368 -5686 21414 -5674
rect 21368 -5862 21374 -5686
rect 21408 -5862 21414 -5686
rect 21826 -5686 21872 -5674
rect 21826 -5834 21832 -5686
rect 21368 -5874 21414 -5862
rect 21820 -5862 21832 -5834
rect 21866 -5834 21872 -5686
rect 22284 -5686 22344 -5306
rect 21866 -5862 21880 -5834
rect 22284 -5842 22290 -5686
rect 17852 -5912 18060 -5906
rect 17852 -5946 17864 -5912
rect 18048 -5946 18060 -5912
rect 17852 -5952 18060 -5946
rect 18310 -5912 18518 -5906
rect 18310 -5946 18322 -5912
rect 18506 -5946 18518 -5912
rect 18310 -5952 18518 -5946
rect 18768 -5912 18976 -5906
rect 18768 -5946 18780 -5912
rect 18964 -5946 18976 -5912
rect 18768 -5952 18976 -5946
rect 19226 -5912 19434 -5906
rect 19226 -5946 19238 -5912
rect 19422 -5946 19434 -5912
rect 19226 -5952 19434 -5946
rect 19684 -5912 19892 -5906
rect 19684 -5946 19696 -5912
rect 19880 -5946 19892 -5912
rect 19684 -5952 19892 -5946
rect 20142 -5912 20350 -5906
rect 20142 -5946 20154 -5912
rect 20338 -5946 20350 -5912
rect 20142 -5952 20350 -5946
rect 20600 -5912 20808 -5906
rect 20600 -5946 20612 -5912
rect 20796 -5946 20808 -5912
rect 20600 -5952 20808 -5946
rect 21058 -5912 21266 -5906
rect 21058 -5946 21070 -5912
rect 21254 -5946 21266 -5912
rect 21058 -5952 21266 -5946
rect 21516 -5912 21724 -5906
rect 21516 -5946 21528 -5912
rect 21712 -5946 21724 -5912
rect 21516 -5952 21724 -5946
rect 17928 -6264 17988 -5952
rect 18384 -6018 18444 -5952
rect 18840 -6018 18900 -5952
rect 19306 -6018 19366 -5952
rect 19756 -6018 19816 -5952
rect 20210 -6018 20270 -5952
rect 20672 -6018 20732 -5952
rect 21126 -6018 21186 -5952
rect 21588 -6018 21648 -5952
rect 18384 -6078 21648 -6018
rect 18390 -6198 21654 -6138
rect 18390 -6264 18450 -6198
rect 18846 -6264 18906 -6198
rect 19312 -6264 19372 -6198
rect 19762 -6264 19822 -6198
rect 20216 -6264 20276 -6198
rect 20678 -6264 20738 -6198
rect 21132 -6264 21192 -6198
rect 21594 -6264 21654 -6198
rect 17852 -6270 18060 -6264
rect 17852 -6304 17864 -6270
rect 18048 -6304 18060 -6270
rect 17852 -6310 18060 -6304
rect 18310 -6270 18518 -6264
rect 18310 -6304 18322 -6270
rect 18506 -6304 18518 -6270
rect 18310 -6310 18518 -6304
rect 18768 -6270 18976 -6264
rect 18768 -6304 18780 -6270
rect 18964 -6304 18976 -6270
rect 18768 -6310 18976 -6304
rect 19226 -6270 19434 -6264
rect 19226 -6304 19238 -6270
rect 19422 -6304 19434 -6270
rect 19226 -6310 19434 -6304
rect 19684 -6270 19892 -6264
rect 19684 -6304 19696 -6270
rect 19880 -6304 19892 -6270
rect 19684 -6310 19892 -6304
rect 20142 -6270 20350 -6264
rect 20142 -6304 20154 -6270
rect 20338 -6304 20350 -6270
rect 20142 -6310 20350 -6304
rect 20600 -6270 20808 -6264
rect 20600 -6304 20612 -6270
rect 20796 -6304 20808 -6270
rect 20600 -6310 20808 -6304
rect 21058 -6270 21266 -6264
rect 21058 -6304 21070 -6270
rect 21254 -6304 21266 -6270
rect 21058 -6310 21266 -6304
rect 21516 -6270 21724 -6264
rect 21516 -6304 21528 -6270
rect 21712 -6304 21724 -6270
rect 21516 -6310 21724 -6304
rect 17324 -6494 17330 -6390
rect 17696 -6410 17710 -6354
rect 17324 -6530 17336 -6494
rect 17704 -6502 17710 -6410
rect 16974 -6580 17182 -6574
rect 16974 -6614 16986 -6580
rect 17170 -6614 17182 -6580
rect 16974 -6620 17182 -6614
rect 17042 -6966 17102 -6620
rect 17276 -6966 17336 -6530
rect 17696 -6530 17710 -6502
rect 17744 -6410 17756 -6354
rect 18162 -6354 18208 -6342
rect 17744 -6502 17750 -6410
rect 18162 -6500 18168 -6354
rect 17744 -6530 17756 -6502
rect 17696 -6966 17756 -6530
rect 18156 -6530 18168 -6500
rect 18202 -6500 18208 -6354
rect 18620 -6354 18666 -6342
rect 18202 -6530 18216 -6500
rect 17852 -6580 18060 -6574
rect 17852 -6614 17864 -6580
rect 18048 -6614 18060 -6580
rect 17852 -6620 18060 -6614
rect 17928 -6966 17988 -6620
rect 18156 -6814 18216 -6530
rect 18620 -6530 18626 -6354
rect 18660 -6530 18666 -6354
rect 18620 -6542 18666 -6530
rect 19078 -6354 19124 -6342
rect 19078 -6530 19084 -6354
rect 19118 -6530 19124 -6354
rect 19078 -6542 19124 -6530
rect 19536 -6354 19582 -6342
rect 19536 -6530 19542 -6354
rect 19576 -6530 19582 -6354
rect 19536 -6542 19582 -6530
rect 19994 -6354 20040 -6342
rect 19994 -6530 20000 -6354
rect 20034 -6530 20040 -6354
rect 19994 -6542 20040 -6530
rect 20452 -6354 20498 -6342
rect 20452 -6530 20458 -6354
rect 20492 -6530 20498 -6354
rect 20452 -6542 20498 -6530
rect 20910 -6354 20956 -6342
rect 20910 -6530 20916 -6354
rect 20950 -6530 20956 -6354
rect 20910 -6542 20956 -6530
rect 21368 -6354 21414 -6342
rect 21368 -6530 21374 -6354
rect 21408 -6530 21414 -6354
rect 21820 -6354 21880 -5862
rect 22276 -5862 22290 -5842
rect 22324 -5716 22344 -5686
rect 22324 -5842 22330 -5716
rect 22324 -5862 22336 -5842
rect 21974 -5912 22182 -5906
rect 21974 -5946 21986 -5912
rect 22170 -5946 22182 -5912
rect 21974 -5952 22182 -5946
rect 22048 -6078 22108 -5952
rect 22276 -6078 22336 -5862
rect 22048 -6138 22336 -6078
rect 22048 -6264 22108 -6138
rect 21974 -6270 22182 -6264
rect 21974 -6304 21986 -6270
rect 22170 -6304 22182 -6270
rect 21974 -6310 22182 -6304
rect 21820 -6396 21832 -6354
rect 21368 -6542 21414 -6530
rect 21826 -6530 21832 -6396
rect 21866 -6396 21880 -6354
rect 22276 -6354 22336 -6138
rect 22276 -6394 22290 -6354
rect 21866 -6530 21872 -6396
rect 22284 -6490 22290 -6394
rect 21826 -6542 21872 -6530
rect 22276 -6530 22290 -6490
rect 22324 -6394 22336 -6354
rect 22324 -6490 22330 -6394
rect 22324 -6530 22336 -6490
rect 18310 -6580 18518 -6574
rect 18310 -6614 18322 -6580
rect 18506 -6614 18518 -6580
rect 18310 -6620 18518 -6614
rect 18768 -6580 18976 -6574
rect 18768 -6614 18780 -6580
rect 18964 -6614 18976 -6580
rect 18768 -6620 18976 -6614
rect 19226 -6580 19434 -6574
rect 19226 -6614 19238 -6580
rect 19422 -6614 19434 -6580
rect 19226 -6620 19434 -6614
rect 19684 -6580 19892 -6574
rect 19684 -6614 19696 -6580
rect 19880 -6614 19892 -6580
rect 19684 -6620 19892 -6614
rect 20142 -6580 20350 -6574
rect 20142 -6614 20154 -6580
rect 20338 -6614 20350 -6580
rect 20142 -6620 20350 -6614
rect 20600 -6580 20808 -6574
rect 20600 -6614 20612 -6580
rect 20796 -6614 20808 -6580
rect 20600 -6620 20808 -6614
rect 21058 -6580 21266 -6574
rect 21058 -6614 21070 -6580
rect 21254 -6614 21266 -6580
rect 21058 -6620 21266 -6614
rect 21516 -6580 21724 -6574
rect 21516 -6614 21528 -6580
rect 21712 -6614 21724 -6580
rect 21516 -6620 21724 -6614
rect 21974 -6580 22182 -6574
rect 21974 -6614 21986 -6580
rect 22170 -6614 22182 -6580
rect 21974 -6620 22182 -6614
rect 18384 -6686 18450 -6620
rect 18840 -6680 18906 -6620
rect 18840 -6686 18846 -6680
rect 18384 -6746 18390 -6686
rect 18450 -6740 18846 -6686
rect 18906 -6686 18912 -6680
rect 19306 -6686 19372 -6620
rect 19756 -6686 19822 -6620
rect 20210 -6686 20276 -6620
rect 20672 -6680 20738 -6620
rect 20672 -6686 20678 -6680
rect 18906 -6740 19312 -6686
rect 18450 -6746 19312 -6740
rect 19372 -6746 19762 -6686
rect 19822 -6746 20216 -6686
rect 20276 -6740 20678 -6686
rect 20738 -6686 20744 -6680
rect 21126 -6686 21192 -6620
rect 21588 -6680 21654 -6620
rect 21588 -6686 21594 -6680
rect 20738 -6740 21132 -6686
rect 20276 -6746 21132 -6740
rect 21192 -6740 21594 -6686
rect 21654 -6740 21660 -6680
rect 21192 -6746 21648 -6740
rect 18156 -6880 18216 -6874
rect 22046 -6966 22106 -6620
rect 22276 -6966 22336 -6530
rect 22644 -6842 22650 -4838
rect 22750 -6842 22756 -4838
rect 22644 -6966 22756 -6842
rect 12300 -6972 22756 -6966
rect 12300 -7072 12406 -6972
rect 22650 -7072 22756 -6972
rect 12300 -7078 22756 -7072
rect 12300 -7308 22756 -7302
rect 12300 -7408 12406 -7308
rect 22650 -7408 22756 -7308
rect 12300 -7414 22756 -7408
rect 12300 -7590 12412 -7414
rect 12300 -12762 12306 -7590
rect 12406 -9384 12412 -7590
rect 12698 -7847 12758 -7414
rect 12926 -7748 12986 -7414
rect 13156 -7488 13216 -7482
rect 12851 -7754 13059 -7748
rect 12851 -7788 12863 -7754
rect 13047 -7788 13059 -7754
rect 12851 -7794 13059 -7788
rect 12698 -7880 12709 -7847
rect 12703 -8970 12709 -7880
rect 12700 -9023 12709 -8970
rect 12743 -7880 12758 -7847
rect 13156 -7847 13216 -7548
rect 13388 -7618 13448 -7612
rect 13844 -7618 13904 -7612
rect 14760 -7618 14820 -7612
rect 13448 -7678 13844 -7620
rect 14310 -7620 14370 -7618
rect 13904 -7624 14760 -7620
rect 13904 -7678 14310 -7624
rect 13388 -7680 14310 -7678
rect 13388 -7748 13448 -7680
rect 13844 -7748 13904 -7680
rect 14370 -7678 14760 -7624
rect 15214 -7618 15274 -7612
rect 14820 -7678 15214 -7620
rect 15676 -7618 15736 -7612
rect 16592 -7616 16652 -7610
rect 15274 -7678 15676 -7620
rect 16130 -7620 16190 -7618
rect 15736 -7624 16592 -7620
rect 15736 -7678 16130 -7624
rect 14370 -7680 16130 -7678
rect 14310 -7748 14370 -7684
rect 14760 -7748 14820 -7680
rect 15214 -7748 15274 -7680
rect 15676 -7748 15736 -7680
rect 16190 -7676 16592 -7624
rect 16190 -7680 16652 -7676
rect 16130 -7748 16190 -7684
rect 16592 -7748 16652 -7680
rect 13309 -7754 13517 -7748
rect 13309 -7788 13321 -7754
rect 13505 -7788 13517 -7754
rect 13309 -7794 13517 -7788
rect 13767 -7754 13975 -7748
rect 13767 -7788 13779 -7754
rect 13963 -7788 13975 -7754
rect 13767 -7794 13975 -7788
rect 14225 -7754 14433 -7748
rect 14225 -7788 14237 -7754
rect 14421 -7788 14433 -7754
rect 14225 -7794 14433 -7788
rect 14683 -7754 14891 -7748
rect 14683 -7788 14695 -7754
rect 14879 -7788 14891 -7754
rect 14683 -7794 14891 -7788
rect 15141 -7754 15349 -7748
rect 15141 -7788 15153 -7754
rect 15337 -7788 15349 -7754
rect 15141 -7794 15349 -7788
rect 15599 -7754 15807 -7748
rect 15599 -7788 15611 -7754
rect 15795 -7788 15807 -7754
rect 15599 -7794 15807 -7788
rect 16057 -7754 16265 -7748
rect 16057 -7788 16069 -7754
rect 16253 -7788 16265 -7754
rect 16057 -7794 16265 -7788
rect 16515 -7754 16723 -7748
rect 16515 -7788 16527 -7754
rect 16711 -7788 16723 -7754
rect 16515 -7794 16723 -7788
rect 13156 -7854 13167 -7847
rect 12743 -8970 12749 -7880
rect 12743 -9023 12760 -8970
rect 12700 -9384 12760 -9023
rect 13161 -9023 13167 -7854
rect 13201 -7854 13216 -7847
rect 13619 -7847 13665 -7835
rect 13201 -9023 13207 -7854
rect 13161 -9035 13207 -9023
rect 13619 -9023 13625 -7847
rect 13659 -9023 13665 -7847
rect 13619 -9035 13665 -9023
rect 14077 -7847 14123 -7835
rect 14077 -9023 14083 -7847
rect 14117 -9023 14123 -7847
rect 14077 -9035 14123 -9023
rect 14535 -7847 14581 -7835
rect 14535 -9023 14541 -7847
rect 14575 -9023 14581 -7847
rect 14535 -9035 14581 -9023
rect 14993 -7847 15039 -7835
rect 14993 -9023 14999 -7847
rect 15033 -9023 15039 -7847
rect 14993 -9035 15039 -9023
rect 15451 -7847 15497 -7835
rect 15451 -9023 15457 -7847
rect 15491 -9023 15497 -7847
rect 15451 -9035 15497 -9023
rect 15909 -7847 15955 -7835
rect 15909 -9023 15915 -7847
rect 15949 -9023 15955 -7847
rect 15909 -9035 15955 -9023
rect 16367 -7847 16413 -7835
rect 16367 -9023 16373 -7847
rect 16407 -9023 16413 -7847
rect 16820 -7847 16880 -7414
rect 17050 -7748 17110 -7414
rect 16973 -7754 17181 -7748
rect 16973 -7788 16985 -7754
rect 17169 -7788 17181 -7754
rect 16973 -7794 17181 -7788
rect 16820 -7888 16831 -7847
rect 16825 -8980 16831 -7888
rect 16367 -9035 16413 -9023
rect 16818 -9023 16831 -8980
rect 16865 -7888 16880 -7847
rect 17278 -7847 17338 -7414
rect 17278 -7882 17289 -7847
rect 16865 -8980 16871 -7888
rect 16865 -9023 16878 -8980
rect 17283 -9002 17289 -7882
rect 12851 -9082 13059 -9076
rect 12851 -9116 12863 -9082
rect 13047 -9116 13059 -9082
rect 12851 -9122 13059 -9116
rect 13309 -9082 13517 -9076
rect 13309 -9116 13321 -9082
rect 13505 -9116 13517 -9082
rect 13309 -9122 13517 -9116
rect 13767 -9082 13975 -9076
rect 13767 -9116 13779 -9082
rect 13963 -9116 13975 -9082
rect 13767 -9122 13975 -9116
rect 14225 -9082 14433 -9076
rect 14225 -9116 14237 -9082
rect 14421 -9116 14433 -9082
rect 14225 -9122 14433 -9116
rect 14683 -9082 14891 -9076
rect 14683 -9116 14695 -9082
rect 14879 -9116 14891 -9082
rect 14683 -9122 14891 -9116
rect 15141 -9082 15349 -9076
rect 15141 -9116 15153 -9082
rect 15337 -9116 15349 -9082
rect 15141 -9122 15349 -9116
rect 15599 -9082 15807 -9076
rect 15599 -9116 15611 -9082
rect 15795 -9116 15807 -9082
rect 15599 -9122 15807 -9116
rect 16057 -9082 16265 -9076
rect 16057 -9116 16069 -9082
rect 16253 -9116 16265 -9082
rect 16057 -9122 16265 -9116
rect 16515 -9082 16723 -9076
rect 16515 -9116 16527 -9082
rect 16711 -9116 16723 -9082
rect 16515 -9122 16723 -9116
rect 12926 -9384 12986 -9122
rect 13388 -9192 13448 -9122
rect 13844 -9192 13904 -9122
rect 14310 -9192 14370 -9122
rect 14760 -9192 14820 -9122
rect 15214 -9192 15274 -9122
rect 15676 -9192 15736 -9122
rect 16130 -9192 16190 -9122
rect 16592 -9192 16652 -9122
rect 13388 -9252 16652 -9192
rect 16818 -9174 16878 -9023
rect 17276 -9023 17289 -9002
rect 17323 -7882 17338 -7847
rect 17698 -7847 17758 -7414
rect 17926 -7748 17986 -7414
rect 18150 -7554 18156 -7494
rect 18216 -7554 18222 -7494
rect 17851 -7754 18059 -7748
rect 17851 -7788 17863 -7754
rect 18047 -7788 18059 -7754
rect 17851 -7794 18059 -7788
rect 17698 -7882 17709 -7847
rect 17323 -9002 17329 -7882
rect 17323 -9023 17336 -9002
rect 17703 -9008 17709 -7882
rect 16973 -9082 17181 -9076
rect 16973 -9116 16985 -9082
rect 17169 -9116 17181 -9082
rect 16973 -9122 17181 -9116
rect 17044 -9174 17104 -9122
rect 17276 -9174 17336 -9023
rect 17696 -9023 17709 -9008
rect 17743 -7882 17758 -7847
rect 18156 -7847 18216 -7554
rect 18390 -7616 18450 -7610
rect 19762 -7614 19822 -7608
rect 18846 -7620 18906 -7614
rect 19312 -7620 19372 -7614
rect 18450 -7676 18846 -7620
rect 18390 -7680 18846 -7676
rect 18906 -7680 19312 -7620
rect 19372 -7674 19762 -7620
rect 20216 -7620 20276 -7614
rect 20678 -7620 20738 -7614
rect 21132 -7616 21192 -7610
rect 19822 -7674 20216 -7620
rect 19372 -7680 20216 -7674
rect 20276 -7680 20678 -7620
rect 20738 -7676 21132 -7620
rect 21594 -7616 21654 -7610
rect 21192 -7676 21594 -7620
rect 20738 -7680 21654 -7676
rect 18390 -7748 18450 -7680
rect 18846 -7748 18906 -7680
rect 19312 -7748 19372 -7680
rect 19762 -7748 19822 -7680
rect 20216 -7748 20276 -7680
rect 20678 -7748 20738 -7680
rect 21132 -7748 21192 -7680
rect 21594 -7748 21654 -7680
rect 22048 -7748 22108 -7414
rect 18309 -7754 18517 -7748
rect 18309 -7788 18321 -7754
rect 18505 -7788 18517 -7754
rect 18309 -7794 18517 -7788
rect 18767 -7754 18975 -7748
rect 18767 -7788 18779 -7754
rect 18963 -7788 18975 -7754
rect 18767 -7794 18975 -7788
rect 19225 -7754 19433 -7748
rect 19225 -7788 19237 -7754
rect 19421 -7788 19433 -7754
rect 19225 -7794 19433 -7788
rect 19683 -7754 19891 -7748
rect 19683 -7788 19695 -7754
rect 19879 -7788 19891 -7754
rect 19683 -7794 19891 -7788
rect 20141 -7754 20349 -7748
rect 20141 -7788 20153 -7754
rect 20337 -7788 20349 -7754
rect 20141 -7794 20349 -7788
rect 20599 -7754 20807 -7748
rect 20599 -7788 20611 -7754
rect 20795 -7788 20807 -7754
rect 20599 -7794 20807 -7788
rect 21057 -7754 21265 -7748
rect 21057 -7788 21069 -7754
rect 21253 -7788 21265 -7754
rect 21057 -7794 21265 -7788
rect 21515 -7754 21723 -7748
rect 21515 -7788 21527 -7754
rect 21711 -7788 21723 -7754
rect 21515 -7794 21723 -7788
rect 21973 -7754 22181 -7748
rect 21973 -7788 21985 -7754
rect 22169 -7788 22181 -7754
rect 21973 -7794 22181 -7788
rect 17743 -9008 17749 -7882
rect 18156 -7914 18167 -7847
rect 17743 -9023 17756 -9008
rect 17696 -9174 17756 -9023
rect 18161 -9023 18167 -7914
rect 18201 -7914 18216 -7847
rect 18619 -7847 18665 -7835
rect 18201 -9023 18207 -7914
rect 18161 -9035 18207 -9023
rect 18619 -9023 18625 -7847
rect 18659 -9023 18665 -7847
rect 18619 -9035 18665 -9023
rect 19077 -7847 19123 -7835
rect 19077 -9023 19083 -7847
rect 19117 -9023 19123 -7847
rect 19077 -9035 19123 -9023
rect 19535 -7847 19581 -7835
rect 19535 -9023 19541 -7847
rect 19575 -9023 19581 -7847
rect 19535 -9035 19581 -9023
rect 19993 -7847 20039 -7835
rect 19993 -9023 19999 -7847
rect 20033 -9023 20039 -7847
rect 19993 -9035 20039 -9023
rect 20451 -7847 20497 -7835
rect 20451 -9023 20457 -7847
rect 20491 -9023 20497 -7847
rect 20451 -9035 20497 -9023
rect 20909 -7847 20955 -7835
rect 20909 -9023 20915 -7847
rect 20949 -9023 20955 -7847
rect 20909 -9035 20955 -9023
rect 21367 -7847 21413 -7835
rect 21367 -9023 21373 -7847
rect 21407 -9023 21413 -7847
rect 21825 -7847 21871 -7835
rect 21825 -8956 21831 -7847
rect 21367 -9035 21413 -9023
rect 21818 -9023 21831 -8956
rect 21865 -8956 21871 -7847
rect 22276 -7847 22336 -7414
rect 22276 -7868 22289 -7847
rect 21865 -9023 21878 -8956
rect 22283 -8976 22289 -7868
rect 17851 -9082 18059 -9076
rect 17851 -9116 17863 -9082
rect 18047 -9116 18059 -9082
rect 17851 -9122 18059 -9116
rect 18309 -9082 18517 -9076
rect 18309 -9116 18321 -9082
rect 18505 -9116 18517 -9082
rect 18309 -9122 18517 -9116
rect 18767 -9082 18975 -9076
rect 18767 -9116 18779 -9082
rect 18963 -9116 18975 -9082
rect 18767 -9122 18975 -9116
rect 19225 -9082 19433 -9076
rect 19225 -9116 19237 -9082
rect 19421 -9116 19433 -9082
rect 19225 -9122 19433 -9116
rect 19683 -9082 19891 -9076
rect 19683 -9116 19695 -9082
rect 19879 -9116 19891 -9082
rect 19683 -9122 19891 -9116
rect 20141 -9082 20349 -9076
rect 20141 -9116 20153 -9082
rect 20337 -9116 20349 -9082
rect 20141 -9122 20349 -9116
rect 20599 -9082 20807 -9076
rect 20599 -9116 20611 -9082
rect 20795 -9116 20807 -9082
rect 20599 -9122 20807 -9116
rect 21057 -9082 21265 -9076
rect 21057 -9116 21069 -9082
rect 21253 -9116 21265 -9082
rect 21057 -9122 21265 -9116
rect 21515 -9082 21723 -9076
rect 21515 -9116 21527 -9082
rect 21711 -9116 21723 -9082
rect 21515 -9122 21723 -9116
rect 17926 -9174 17986 -9122
rect 16818 -9234 17986 -9174
rect 18382 -9192 18442 -9122
rect 18838 -9192 18898 -9122
rect 19304 -9192 19364 -9122
rect 19754 -9192 19814 -9122
rect 20208 -9192 20268 -9122
rect 20670 -9192 20730 -9122
rect 21124 -9192 21184 -9122
rect 21586 -9192 21646 -9122
rect 18382 -9252 21646 -9192
rect 21818 -9294 21878 -9023
rect 22276 -9023 22289 -8976
rect 22323 -7868 22336 -7847
rect 22644 -7590 22756 -7414
rect 22323 -8976 22329 -7868
rect 22323 -9023 22336 -8976
rect 21973 -9082 22181 -9076
rect 21973 -9116 21985 -9082
rect 22169 -9116 22181 -9082
rect 21973 -9122 22181 -9116
rect 21812 -9354 21818 -9294
rect 21878 -9354 21884 -9294
rect 12406 -9444 13536 -9384
rect 12406 -9878 12412 -9444
rect 13476 -9878 13536 -9444
rect 14388 -9460 20864 -9400
rect 22048 -9448 22108 -9122
rect 22276 -9448 22336 -9023
rect 22644 -9448 22650 -7590
rect 12406 -9938 13994 -9878
rect 12406 -12762 12412 -9938
rect 13476 -10112 13536 -9938
rect 13702 -10013 13762 -9938
rect 13628 -10019 13836 -10013
rect 13628 -10053 13640 -10019
rect 13824 -10053 13836 -10019
rect 13628 -10059 13836 -10053
rect 13476 -10156 13486 -10112
rect 13480 -11618 13486 -10156
rect 13472 -11688 13486 -11618
rect 13520 -10156 13536 -10112
rect 13934 -10112 13994 -9938
rect 14158 -9940 14164 -9880
rect 14224 -9940 14230 -9880
rect 14164 -10013 14224 -9940
rect 14086 -10019 14294 -10013
rect 14086 -10053 14098 -10019
rect 14282 -10053 14294 -10019
rect 14086 -10059 14294 -10053
rect 13520 -11618 13526 -10156
rect 13934 -10174 13944 -10112
rect 13938 -11612 13944 -10174
rect 13520 -11688 13532 -11618
rect 13472 -12476 13532 -11688
rect 13930 -11688 13944 -11612
rect 13978 -10174 13994 -10112
rect 14388 -10112 14448 -9460
rect 15302 -9590 19946 -9530
rect 14618 -9940 14624 -9880
rect 14684 -9940 14690 -9880
rect 15076 -9940 15082 -9880
rect 15142 -9940 15148 -9880
rect 14624 -10013 14684 -9940
rect 15082 -10013 15142 -9940
rect 14544 -10019 14752 -10013
rect 14544 -10053 14556 -10019
rect 14740 -10053 14752 -10019
rect 14544 -10059 14752 -10053
rect 15002 -10019 15210 -10013
rect 15002 -10053 15014 -10019
rect 15198 -10053 15210 -10019
rect 15002 -10059 15210 -10053
rect 14388 -10172 14402 -10112
rect 13978 -11612 13984 -10174
rect 13978 -11688 13990 -11612
rect 13628 -11747 13836 -11741
rect 13628 -11781 13640 -11747
rect 13824 -11781 13836 -11747
rect 13628 -11787 13836 -11781
rect 13700 -12476 13760 -11787
rect 13930 -12476 13990 -11688
rect 14396 -11688 14402 -10172
rect 14436 -10172 14448 -10112
rect 14854 -10112 14900 -10100
rect 14436 -11688 14442 -10172
rect 14854 -11632 14860 -10112
rect 14396 -11700 14442 -11688
rect 14846 -11688 14860 -11632
rect 14894 -11632 14900 -10112
rect 15302 -10112 15362 -9590
rect 16222 -9716 19038 -9656
rect 15532 -9940 15538 -9880
rect 15598 -9940 15604 -9880
rect 15988 -9940 15994 -9880
rect 16054 -9940 16060 -9880
rect 15538 -10013 15598 -9940
rect 15994 -10013 16054 -9940
rect 15460 -10019 15668 -10013
rect 15460 -10053 15472 -10019
rect 15656 -10053 15668 -10019
rect 15460 -10059 15668 -10053
rect 15918 -10019 16126 -10013
rect 15918 -10053 15930 -10019
rect 16114 -10053 16126 -10019
rect 15918 -10059 16126 -10053
rect 15302 -10180 15318 -10112
rect 14894 -11688 14906 -11632
rect 14086 -11747 14294 -11741
rect 14086 -11781 14098 -11747
rect 14282 -11781 14294 -11747
rect 14086 -11787 14294 -11781
rect 14544 -11747 14752 -11741
rect 14544 -11781 14556 -11747
rect 14740 -11781 14752 -11747
rect 14544 -11787 14752 -11781
rect 14160 -11854 14220 -11787
rect 14620 -11854 14680 -11787
rect 14154 -11914 14160 -11854
rect 14220 -11914 14226 -11854
rect 14614 -11914 14620 -11854
rect 14680 -11914 14686 -11854
rect 14846 -12222 14906 -11688
rect 15312 -11688 15318 -10180
rect 15352 -10180 15362 -10112
rect 15770 -10112 15816 -10100
rect 15352 -11688 15358 -10180
rect 15770 -11630 15776 -10112
rect 15312 -11700 15358 -11688
rect 15766 -11688 15776 -11630
rect 15810 -11630 15816 -10112
rect 16222 -10112 16282 -9716
rect 17136 -9832 18114 -9772
rect 16444 -9940 16450 -9880
rect 16510 -9940 16516 -9880
rect 16904 -9940 16910 -9880
rect 16970 -9940 16976 -9880
rect 16450 -10013 16510 -9940
rect 16910 -10013 16970 -9940
rect 16376 -10019 16584 -10013
rect 16376 -10053 16388 -10019
rect 16572 -10053 16584 -10019
rect 16376 -10059 16584 -10053
rect 16834 -10019 17042 -10013
rect 16834 -10053 16846 -10019
rect 17030 -10053 17042 -10019
rect 16834 -10059 17042 -10053
rect 16222 -10144 16234 -10112
rect 15810 -11688 15826 -11630
rect 15002 -11747 15210 -11741
rect 15002 -11781 15014 -11747
rect 15198 -11781 15210 -11747
rect 15002 -11787 15210 -11781
rect 15460 -11747 15668 -11741
rect 15460 -11781 15472 -11747
rect 15656 -11781 15668 -11747
rect 15460 -11787 15668 -11781
rect 15078 -11854 15138 -11787
rect 15534 -11854 15594 -11787
rect 15072 -11914 15078 -11854
rect 15138 -11914 15144 -11854
rect 15528 -11914 15534 -11854
rect 15594 -11914 15600 -11854
rect 15766 -12088 15826 -11688
rect 16228 -11688 16234 -10144
rect 16268 -10144 16282 -10112
rect 16686 -10112 16732 -10100
rect 16268 -11688 16274 -10144
rect 16686 -11644 16692 -10112
rect 16228 -11700 16274 -11688
rect 16682 -11688 16692 -11644
rect 16726 -11644 16732 -10112
rect 17136 -10112 17196 -9832
rect 17354 -9880 17438 -9876
rect 17354 -9942 17366 -9880
rect 17426 -9942 17438 -9880
rect 17354 -9948 17438 -9942
rect 17592 -9892 17652 -9886
rect 17366 -10013 17426 -9948
rect 17820 -9940 17826 -9880
rect 17886 -9940 17892 -9880
rect 17820 -9942 17892 -9940
rect 17292 -10019 17500 -10013
rect 17292 -10053 17304 -10019
rect 17488 -10053 17500 -10019
rect 17292 -10059 17500 -10053
rect 17136 -10140 17150 -10112
rect 16726 -11688 16742 -11644
rect 15918 -11747 16126 -11741
rect 15918 -11781 15930 -11747
rect 16114 -11781 16126 -11747
rect 15918 -11787 16126 -11781
rect 16376 -11747 16584 -11741
rect 16376 -11781 16388 -11747
rect 16572 -11781 16584 -11747
rect 16376 -11787 16584 -11781
rect 15990 -11854 16050 -11787
rect 16446 -11854 16506 -11787
rect 15984 -11914 15990 -11854
rect 16050 -11914 16056 -11854
rect 16440 -11914 16446 -11854
rect 16506 -11914 16512 -11854
rect 16682 -11964 16742 -11688
rect 17144 -11688 17150 -10140
rect 17184 -10140 17196 -10112
rect 17592 -10112 17652 -9952
rect 17826 -10013 17886 -9942
rect 17750 -10019 17958 -10013
rect 17750 -10053 17762 -10019
rect 17946 -10053 17958 -10019
rect 17750 -10059 17958 -10053
rect 17592 -10134 17608 -10112
rect 17184 -11688 17190 -10140
rect 17144 -11700 17190 -11688
rect 17602 -11688 17608 -10134
rect 17642 -10134 17652 -10112
rect 18054 -10112 18114 -9832
rect 18278 -9940 18284 -9880
rect 18344 -9940 18350 -9880
rect 18732 -9940 18738 -9880
rect 18798 -9940 18804 -9880
rect 18284 -10013 18344 -9940
rect 18738 -10013 18798 -9940
rect 18208 -10019 18416 -10013
rect 18208 -10053 18220 -10019
rect 18404 -10053 18416 -10019
rect 18208 -10059 18416 -10053
rect 18666 -10019 18874 -10013
rect 18666 -10053 18678 -10019
rect 18862 -10053 18874 -10019
rect 18666 -10059 18874 -10053
rect 18978 -10100 19038 -9716
rect 19196 -9940 19202 -9880
rect 19262 -9940 19268 -9880
rect 19654 -9940 19660 -9880
rect 19720 -9940 19726 -9880
rect 19202 -10013 19262 -9940
rect 19660 -10013 19720 -9940
rect 19124 -10019 19332 -10013
rect 19124 -10053 19136 -10019
rect 19320 -10053 19332 -10019
rect 19124 -10059 19332 -10053
rect 19582 -10019 19790 -10013
rect 19582 -10053 19594 -10019
rect 19778 -10053 19790 -10019
rect 19582 -10059 19790 -10053
rect 17642 -11688 17648 -10134
rect 18054 -10192 18066 -10112
rect 17602 -11700 17648 -11688
rect 18060 -11688 18066 -10192
rect 18100 -10192 18114 -10112
rect 18518 -10112 18564 -10100
rect 18100 -11688 18106 -10192
rect 18518 -11610 18524 -10112
rect 18060 -11700 18106 -11688
rect 18512 -11688 18524 -11610
rect 18558 -11610 18564 -10112
rect 18976 -10112 19038 -10100
rect 18558 -11688 18572 -11610
rect 16834 -11747 17042 -11741
rect 16834 -11781 16846 -11747
rect 17030 -11781 17042 -11747
rect 16834 -11787 17042 -11781
rect 17292 -11747 17500 -11741
rect 17292 -11781 17304 -11747
rect 17488 -11781 17500 -11747
rect 17292 -11787 17500 -11781
rect 17750 -11747 17958 -11741
rect 17750 -11781 17762 -11747
rect 17946 -11781 17958 -11747
rect 17750 -11787 17958 -11781
rect 18208 -11747 18416 -11741
rect 18208 -11781 18220 -11747
rect 18404 -11781 18416 -11747
rect 18208 -11787 18416 -11781
rect 16902 -11854 16962 -11787
rect 17360 -11854 17420 -11787
rect 17828 -11854 17888 -11787
rect 18284 -11854 18344 -11787
rect 16896 -11914 16902 -11854
rect 16962 -11914 16968 -11854
rect 17354 -11914 17360 -11854
rect 17420 -11914 17426 -11854
rect 17822 -11914 17828 -11854
rect 17888 -11914 17894 -11854
rect 18278 -11914 18284 -11854
rect 18344 -11914 18350 -11854
rect 18512 -11964 18572 -11688
rect 18976 -11688 18982 -10112
rect 19016 -10184 19038 -10112
rect 19434 -10112 19480 -10100
rect 19016 -11688 19022 -10184
rect 19434 -11628 19440 -10112
rect 18976 -11700 19022 -11688
rect 19428 -11688 19440 -11628
rect 19474 -11628 19480 -10112
rect 19886 -10112 19946 -9590
rect 20110 -9940 20116 -9880
rect 20176 -9940 20182 -9880
rect 20570 -9940 20576 -9880
rect 20636 -9940 20642 -9880
rect 20116 -10013 20176 -9940
rect 20576 -10013 20636 -9940
rect 20040 -10019 20248 -10013
rect 20040 -10053 20052 -10019
rect 20236 -10053 20248 -10019
rect 20040 -10059 20248 -10053
rect 20498 -10019 20706 -10013
rect 20498 -10053 20510 -10019
rect 20694 -10053 20706 -10019
rect 20498 -10059 20706 -10053
rect 19886 -10190 19898 -10112
rect 19474 -11688 19488 -11628
rect 18666 -11747 18874 -11741
rect 18666 -11781 18678 -11747
rect 18862 -11781 18874 -11747
rect 18666 -11787 18874 -11781
rect 19124 -11747 19332 -11741
rect 19124 -11781 19136 -11747
rect 19320 -11781 19332 -11747
rect 19124 -11787 19332 -11781
rect 18734 -11854 18794 -11787
rect 19198 -11854 19258 -11787
rect 18728 -11914 18734 -11854
rect 18794 -11914 18800 -11854
rect 19192 -11914 19198 -11854
rect 19258 -11914 19264 -11854
rect 16682 -12024 18572 -11964
rect 19428 -12088 19488 -11688
rect 19892 -11688 19898 -10190
rect 19932 -10190 19946 -10112
rect 20350 -10112 20396 -10100
rect 19932 -11688 19938 -10190
rect 20350 -11630 20356 -10112
rect 19892 -11700 19938 -11688
rect 20344 -11688 20356 -11630
rect 20390 -11630 20396 -10112
rect 20804 -10112 20864 -9460
rect 21716 -9508 22650 -9448
rect 21716 -9880 21776 -9508
rect 22644 -9880 22650 -9508
rect 21026 -9940 21032 -9880
rect 21092 -9940 21098 -9880
rect 21262 -9940 22650 -9880
rect 21032 -10013 21092 -9940
rect 20956 -10019 21164 -10013
rect 20956 -10053 20968 -10019
rect 21152 -10053 21164 -10019
rect 20956 -10059 21164 -10053
rect 20804 -10196 20814 -10112
rect 20390 -11688 20404 -11630
rect 19582 -11747 19790 -11741
rect 19582 -11781 19594 -11747
rect 19778 -11781 19790 -11747
rect 19582 -11787 19790 -11781
rect 20040 -11747 20248 -11741
rect 20040 -11781 20052 -11747
rect 20236 -11781 20248 -11747
rect 20040 -11787 20248 -11781
rect 19656 -11854 19716 -11787
rect 20112 -11854 20172 -11787
rect 19650 -11914 19656 -11854
rect 19716 -11914 19722 -11854
rect 20106 -11914 20112 -11854
rect 20172 -11914 20178 -11854
rect 15766 -12148 19488 -12088
rect 20344 -12222 20404 -11688
rect 20808 -11688 20814 -10196
rect 20848 -10196 20864 -10112
rect 21262 -10112 21322 -9940
rect 21488 -10013 21548 -9940
rect 21414 -10019 21622 -10013
rect 21414 -10053 21426 -10019
rect 21610 -10053 21622 -10019
rect 21414 -10059 21622 -10053
rect 21262 -10156 21272 -10112
rect 20848 -11688 20854 -10196
rect 21266 -11624 21272 -10156
rect 20808 -11700 20854 -11688
rect 21260 -11688 21272 -11624
rect 21306 -10156 21322 -10112
rect 21716 -10112 21776 -9940
rect 21306 -11624 21312 -10156
rect 21716 -10172 21730 -10112
rect 21306 -11688 21320 -11624
rect 21724 -11656 21730 -10172
rect 20498 -11747 20706 -11741
rect 20498 -11781 20510 -11747
rect 20694 -11781 20706 -11747
rect 20498 -11787 20706 -11781
rect 20956 -11747 21164 -11741
rect 20956 -11781 20968 -11747
rect 21152 -11781 21164 -11747
rect 20956 -11787 21164 -11781
rect 20572 -11854 20632 -11787
rect 21028 -11854 21088 -11787
rect 20566 -11914 20572 -11854
rect 20632 -11914 20638 -11854
rect 21022 -11914 21028 -11854
rect 21088 -11914 21094 -11854
rect 14846 -12282 20404 -12222
rect 21260 -12476 21320 -11688
rect 21718 -11688 21730 -11656
rect 21764 -10172 21776 -10112
rect 21764 -11656 21770 -10172
rect 21764 -11688 21778 -11656
rect 21414 -11747 21622 -11741
rect 21414 -11781 21426 -11747
rect 21610 -11781 21622 -11747
rect 21414 -11787 21622 -11781
rect 21486 -12476 21546 -11787
rect 21718 -12476 21778 -11688
rect 13450 -12486 21806 -12476
rect 13450 -12572 13476 -12486
rect 13572 -12572 13896 -12486
rect 13992 -12572 14496 -12486
rect 14592 -12572 15096 -12486
rect 15192 -12572 15696 -12486
rect 15792 -12572 16296 -12486
rect 16392 -12572 16896 -12486
rect 16992 -12572 17496 -12486
rect 17592 -12572 18096 -12486
rect 18192 -12572 18696 -12486
rect 18792 -12572 19296 -12486
rect 19392 -12572 19896 -12486
rect 19992 -12572 20496 -12486
rect 20592 -12572 21096 -12486
rect 21192 -12572 21696 -12486
rect 21792 -12572 21806 -12486
rect 13450 -12586 21806 -12572
rect 12300 -13046 12412 -12762
rect 13012 -13046 13022 -12746
rect 22034 -13046 22044 -12746
rect 22644 -12762 22650 -9940
rect 22750 -12762 22756 -7590
rect 22644 -13046 22756 -12762
rect 12300 -13052 22756 -13046
rect 12300 -13152 12406 -13052
rect 22650 -13152 22756 -13052
rect 12300 -13158 22756 -13152
rect 22940 -9880 23000 3092
rect 23080 -3226 23140 8564
rect 23536 8618 28992 8624
rect 23536 8518 23642 8618
rect 28886 8518 28992 8618
rect 30820 8588 30826 8648
rect 30886 8588 30892 8648
rect 32230 8632 32242 8680
rect 32290 8632 32358 8680
rect 32406 8632 32418 8680
rect 32230 8626 32418 8632
rect 32458 8680 32888 8686
rect 32954 8684 33014 8690
rect 32458 8632 32470 8680
rect 32518 8632 32602 8680
rect 32650 8632 32712 8680
rect 32760 8632 32828 8680
rect 32876 8632 32888 8680
rect 32458 8626 32888 8632
rect 32948 8624 32954 8684
rect 33014 8624 33020 8684
rect 32954 8618 33014 8624
rect 30826 8582 30886 8588
rect 31930 8568 31990 8574
rect 23536 8512 28992 8518
rect 23536 8335 23648 8512
rect 23536 5442 23542 8335
rect 23534 5332 23542 5442
rect 23536 5049 23542 5332
rect 23642 6844 23648 8335
rect 23918 8225 23978 8512
rect 24146 8324 24206 8512
rect 24073 8318 24281 8324
rect 24073 8284 24085 8318
rect 24269 8284 24281 8318
rect 24073 8278 24281 8284
rect 23918 8202 23931 8225
rect 23925 7094 23931 8202
rect 23918 7049 23931 7094
rect 23965 8202 23978 8225
rect 24376 8225 24436 8512
rect 28038 8456 28098 8462
rect 24600 8450 24660 8456
rect 25062 8450 25122 8456
rect 25516 8450 25576 8456
rect 25978 8450 26038 8456
rect 26432 8450 26492 8456
rect 26882 8450 26942 8456
rect 27348 8450 27408 8456
rect 27804 8450 27864 8456
rect 24594 8390 24600 8450
rect 24660 8390 25062 8450
rect 25122 8390 25516 8450
rect 25576 8390 25978 8450
rect 26038 8390 26432 8450
rect 26492 8390 26882 8450
rect 26942 8390 27348 8450
rect 27408 8390 27804 8450
rect 27864 8390 27870 8450
rect 24600 8324 24660 8390
rect 25062 8324 25122 8390
rect 25516 8324 25576 8390
rect 25978 8324 26038 8390
rect 26432 8324 26492 8390
rect 26882 8324 26942 8390
rect 27348 8324 27408 8390
rect 27804 8324 27864 8390
rect 24531 8318 24739 8324
rect 24531 8284 24543 8318
rect 24727 8284 24739 8318
rect 24531 8278 24739 8284
rect 24989 8318 25197 8324
rect 24989 8284 25001 8318
rect 25185 8284 25197 8318
rect 24989 8278 25197 8284
rect 25447 8318 25655 8324
rect 25447 8284 25459 8318
rect 25643 8284 25655 8318
rect 25447 8278 25655 8284
rect 25905 8318 26113 8324
rect 25905 8284 25917 8318
rect 26101 8284 26113 8318
rect 25905 8278 26113 8284
rect 26363 8318 26571 8324
rect 26363 8284 26375 8318
rect 26559 8284 26571 8318
rect 26363 8278 26571 8284
rect 26821 8318 27029 8324
rect 26821 8284 26833 8318
rect 27017 8284 27029 8318
rect 26821 8278 27029 8284
rect 27279 8318 27487 8324
rect 27279 8284 27291 8318
rect 27475 8284 27487 8318
rect 27279 8278 27487 8284
rect 27737 8318 27945 8324
rect 27737 8284 27749 8318
rect 27933 8284 27945 8318
rect 27737 8278 27945 8284
rect 23965 7094 23971 8202
rect 23965 7049 23978 7094
rect 23918 6844 23978 7049
rect 24376 7049 24389 8225
rect 24423 7049 24436 8225
rect 24073 6990 24281 6996
rect 24073 6956 24085 6990
rect 24269 6956 24281 6990
rect 24073 6950 24281 6956
rect 24146 6844 24206 6950
rect 24376 6844 24436 7049
rect 24841 8225 24887 8237
rect 24841 7049 24847 8225
rect 24881 7049 24887 8225
rect 24841 7037 24887 7049
rect 25299 8225 25345 8237
rect 25299 7049 25305 8225
rect 25339 7049 25345 8225
rect 25299 7037 25345 7049
rect 25757 8225 25803 8237
rect 25757 7049 25763 8225
rect 25797 7049 25803 8225
rect 25757 7037 25803 7049
rect 26215 8225 26261 8237
rect 26215 7049 26221 8225
rect 26255 7049 26261 8225
rect 26215 7037 26261 7049
rect 26673 8225 26719 8237
rect 26673 7049 26679 8225
rect 26713 7049 26719 8225
rect 26673 7037 26719 7049
rect 27131 8225 27177 8237
rect 27131 7049 27137 8225
rect 27171 7049 27177 8225
rect 27131 7037 27177 7049
rect 27589 8225 27635 8237
rect 27589 7049 27595 8225
rect 27629 7049 27635 8225
rect 28038 8225 28098 8396
rect 28268 8324 28328 8512
rect 28195 8318 28403 8324
rect 28195 8284 28207 8318
rect 28391 8284 28403 8318
rect 28195 8278 28403 8284
rect 28038 8156 28053 8225
rect 27589 7037 27635 7049
rect 28047 7049 28053 8156
rect 28087 8156 28098 8225
rect 28496 8225 28556 8512
rect 28496 8188 28511 8225
rect 28087 7049 28093 8156
rect 28505 7062 28511 8188
rect 28047 7037 28093 7049
rect 28498 7049 28511 7062
rect 28545 8188 28556 8225
rect 28880 8418 28992 8512
rect 31924 8508 31930 8568
rect 31990 8508 31996 8568
rect 31930 8502 31990 8508
rect 30210 8452 36076 8464
rect 30210 8433 30406 8452
rect 28880 8387 29812 8418
rect 28880 8353 29105 8387
rect 29139 8353 29197 8387
rect 29231 8353 29289 8387
rect 29323 8353 29381 8387
rect 29415 8353 29473 8387
rect 29507 8353 29565 8387
rect 29599 8353 29657 8387
rect 29691 8353 29749 8387
rect 29783 8353 29812 8387
rect 30210 8399 30239 8433
rect 30273 8399 30406 8433
rect 30210 8380 30406 8399
rect 30502 8433 35784 8452
rect 30502 8399 30581 8433
rect 30615 8399 30673 8433
rect 30707 8399 30765 8433
rect 30799 8399 30857 8433
rect 30891 8399 30949 8433
rect 30983 8399 31041 8433
rect 31075 8399 31133 8433
rect 31167 8399 31225 8433
rect 31259 8399 31317 8433
rect 31351 8399 31409 8433
rect 31443 8399 31501 8433
rect 31535 8399 31593 8433
rect 31627 8399 31685 8433
rect 31719 8399 31777 8433
rect 31811 8399 31869 8433
rect 31903 8399 31961 8433
rect 31995 8399 32053 8433
rect 32087 8399 32145 8433
rect 32179 8399 32237 8433
rect 32271 8399 32329 8433
rect 32363 8399 32421 8433
rect 32455 8399 32513 8433
rect 32547 8399 32605 8433
rect 32639 8399 32697 8433
rect 32731 8399 32789 8433
rect 32823 8399 32881 8433
rect 32915 8399 32973 8433
rect 33007 8399 33139 8433
rect 33173 8399 33279 8433
rect 33313 8399 33371 8433
rect 33405 8399 33463 8433
rect 33497 8399 33555 8433
rect 33589 8399 33647 8433
rect 33681 8399 33739 8433
rect 33773 8399 33831 8433
rect 33865 8399 33923 8433
rect 33957 8399 34015 8433
rect 34049 8399 34107 8433
rect 34141 8399 34199 8433
rect 34233 8399 34291 8433
rect 34325 8399 34383 8433
rect 34417 8399 34475 8433
rect 34509 8399 34567 8433
rect 34601 8399 34659 8433
rect 34693 8399 34751 8433
rect 34785 8399 34843 8433
rect 34877 8399 34935 8433
rect 34969 8399 35027 8433
rect 35061 8399 35119 8433
rect 35153 8399 35211 8433
rect 35245 8399 35303 8433
rect 35337 8399 35395 8433
rect 35429 8399 35487 8433
rect 35521 8399 35579 8433
rect 35613 8399 35671 8433
rect 35705 8399 35784 8433
rect 30502 8380 35784 8399
rect 35880 8433 36076 8452
rect 35880 8399 36013 8433
rect 36047 8399 36076 8433
rect 35880 8380 36076 8399
rect 30210 8368 36076 8380
rect 28880 8335 29812 8353
rect 28545 7062 28551 8188
rect 28545 7049 28558 7062
rect 24531 6990 24739 6996
rect 24531 6956 24543 6990
rect 24727 6956 24739 6990
rect 24531 6950 24739 6956
rect 24989 6990 25197 6996
rect 24989 6956 25001 6990
rect 25185 6956 25197 6990
rect 24989 6950 25197 6956
rect 25447 6990 25655 6996
rect 25447 6956 25459 6990
rect 25643 6956 25655 6990
rect 25447 6950 25655 6956
rect 25905 6990 26113 6996
rect 25905 6956 25917 6990
rect 26101 6956 26113 6990
rect 25905 6950 26113 6956
rect 26363 6990 26571 6996
rect 26363 6956 26375 6990
rect 26559 6956 26571 6990
rect 26363 6950 26571 6956
rect 26821 6990 27029 6996
rect 26821 6956 26833 6990
rect 27017 6956 27029 6990
rect 26821 6950 27029 6956
rect 27279 6990 27487 6996
rect 27279 6956 27291 6990
rect 27475 6956 27487 6990
rect 27279 6950 27487 6956
rect 27737 6990 27945 6996
rect 27737 6956 27749 6990
rect 27933 6956 27945 6990
rect 27737 6950 27945 6956
rect 28195 6990 28403 6996
rect 28195 6956 28207 6990
rect 28391 6956 28403 6990
rect 28195 6950 28403 6956
rect 23642 6784 24436 6844
rect 24608 6878 24668 6950
rect 25070 6878 25130 6950
rect 25524 6878 25584 6950
rect 25986 6878 26046 6950
rect 26440 6878 26500 6950
rect 26890 6878 26950 6950
rect 27356 6878 27416 6950
rect 27812 6878 27872 6950
rect 28268 6896 28328 6950
rect 28498 6896 28558 7049
rect 28880 6896 28886 8335
rect 24608 6818 27812 6878
rect 27872 6818 27878 6878
rect 28268 6836 28886 6896
rect 23642 5442 23648 6784
rect 23918 5442 23978 6784
rect 24146 5442 24206 6784
rect 24376 5442 24436 6784
rect 28268 5442 28328 6836
rect 28498 5442 28558 6836
rect 23642 5432 28808 5442
rect 23642 5346 23824 5432
rect 23920 5346 24424 5432
rect 24520 5346 25024 5432
rect 25120 5346 25624 5432
rect 25720 5346 26224 5432
rect 26320 5346 26824 5432
rect 26920 5346 27424 5432
rect 27520 5346 28024 5432
rect 28120 5346 28624 5432
rect 28720 5346 28808 5432
rect 23642 5332 28808 5346
rect 23642 5049 23648 5332
rect 23536 4872 23648 5049
rect 24248 4872 24258 5172
rect 28270 4872 28280 5172
rect 28880 5049 28886 6836
rect 28986 8322 29812 8335
rect 28986 5049 28992 8322
rect 34630 8320 34690 8326
rect 34624 8260 34630 8320
rect 34690 8260 34696 8320
rect 34630 8254 34690 8260
rect 30826 8244 30886 8250
rect 33524 8244 33584 8250
rect 30570 8196 30630 8202
rect 30564 8136 30570 8196
rect 30630 8136 30636 8196
rect 30820 8184 30826 8244
rect 30886 8184 30892 8244
rect 32230 8200 32418 8206
rect 30826 8178 30886 8184
rect 32230 8152 32242 8200
rect 32290 8152 32358 8200
rect 32406 8152 32418 8200
rect 32230 8146 32418 8152
rect 32458 8200 32888 8206
rect 32458 8152 32470 8200
rect 32518 8152 32602 8200
rect 32650 8152 32712 8200
rect 32760 8152 32828 8200
rect 32876 8152 32888 8200
rect 32458 8146 32888 8152
rect 32946 8148 32952 8208
rect 33012 8148 33024 8208
rect 33518 8184 33524 8244
rect 33584 8184 33590 8244
rect 35652 8208 35712 8214
rect 34928 8200 35116 8206
rect 33524 8178 33584 8184
rect 33268 8154 33328 8160
rect 30570 8130 30630 8136
rect 30745 8127 30803 8133
rect 30745 8093 30757 8127
rect 30791 8124 30803 8127
rect 30983 8127 31041 8133
rect 30983 8124 30995 8127
rect 30791 8096 30995 8124
rect 30791 8093 30803 8096
rect 30745 8087 30803 8093
rect 30983 8093 30995 8096
rect 31029 8124 31041 8127
rect 31487 8127 31545 8133
rect 31487 8124 31499 8127
rect 31029 8096 31499 8124
rect 31029 8093 31041 8096
rect 30983 8087 31041 8093
rect 31487 8093 31499 8096
rect 31533 8093 31545 8127
rect 33262 8094 33268 8154
rect 33328 8094 33334 8154
rect 34928 8152 34940 8200
rect 34988 8152 35056 8200
rect 35104 8152 35116 8200
rect 34928 8146 35116 8152
rect 35156 8200 35586 8206
rect 35156 8152 35168 8200
rect 35216 8152 35300 8200
rect 35348 8152 35410 8200
rect 35458 8152 35526 8200
rect 35574 8152 35586 8200
rect 35156 8146 35586 8152
rect 35646 8148 35652 8208
rect 35712 8148 35718 8208
rect 35652 8142 35712 8148
rect 33443 8127 33501 8133
rect 31487 8087 31545 8093
rect 33268 8088 33328 8094
rect 33443 8093 33455 8127
rect 33489 8124 33501 8127
rect 33681 8127 33739 8133
rect 33681 8124 33693 8127
rect 33489 8096 33693 8124
rect 33489 8093 33501 8096
rect 33443 8087 33501 8093
rect 33681 8093 33693 8096
rect 33727 8124 33739 8127
rect 34185 8127 34243 8133
rect 34185 8124 34197 8127
rect 33727 8096 34197 8124
rect 33727 8093 33739 8096
rect 33681 8087 33739 8093
rect 34185 8093 34197 8096
rect 34231 8093 34243 8127
rect 34185 8087 34243 8093
rect 30666 8059 30724 8065
rect 30666 8025 30678 8059
rect 30712 8056 30724 8059
rect 31086 8059 31144 8065
rect 31086 8056 31098 8059
rect 30712 8028 31098 8056
rect 30712 8025 30724 8028
rect 30666 8019 30724 8025
rect 31086 8025 31098 8028
rect 31132 8056 31144 8059
rect 31400 8059 31458 8065
rect 31400 8056 31412 8059
rect 31132 8028 31412 8056
rect 31132 8025 31144 8028
rect 31086 8019 31144 8025
rect 31400 8025 31412 8028
rect 31446 8025 31458 8059
rect 33364 8059 33422 8065
rect 31400 8019 31458 8025
rect 31930 8022 31990 8028
rect 33364 8025 33376 8059
rect 33410 8056 33422 8059
rect 33784 8059 33842 8065
rect 33784 8056 33796 8059
rect 33410 8028 33796 8056
rect 33410 8025 33422 8028
rect 31924 7962 31930 8022
rect 31990 7962 31996 8022
rect 33364 8019 33422 8025
rect 33784 8025 33796 8028
rect 33830 8056 33842 8059
rect 34098 8059 34156 8065
rect 34098 8056 34110 8059
rect 33830 8028 34110 8056
rect 33830 8025 33842 8028
rect 33784 8019 33842 8025
rect 34098 8025 34110 8028
rect 34144 8025 34156 8059
rect 34098 8019 34156 8025
rect 31930 7956 31990 7962
rect 30210 7908 36076 7920
rect 30210 7889 33086 7908
rect 30210 7855 30239 7889
rect 30273 7855 30581 7889
rect 30615 7855 30673 7889
rect 30707 7855 30765 7889
rect 30799 7855 30857 7889
rect 30891 7855 30949 7889
rect 30983 7855 31041 7889
rect 31075 7855 31133 7889
rect 31167 7855 31225 7889
rect 31259 7855 31317 7889
rect 31351 7855 31409 7889
rect 31443 7855 31501 7889
rect 31535 7855 31593 7889
rect 31627 7855 31685 7889
rect 31719 7855 31777 7889
rect 31811 7855 31869 7889
rect 31903 7855 31961 7889
rect 31995 7855 32053 7889
rect 32087 7855 32145 7889
rect 32179 7855 32237 7889
rect 32271 7855 32329 7889
rect 32363 7855 32421 7889
rect 32455 7855 32513 7889
rect 32547 7855 32605 7889
rect 32639 7855 32697 7889
rect 32731 7855 32789 7889
rect 32823 7855 32881 7889
rect 32915 7855 32973 7889
rect 33007 7855 33086 7889
rect 30210 7836 33086 7855
rect 33182 7889 36076 7908
rect 33182 7855 33279 7889
rect 33313 7855 33371 7889
rect 33405 7855 33463 7889
rect 33497 7855 33555 7889
rect 33589 7855 33647 7889
rect 33681 7855 33739 7889
rect 33773 7855 33831 7889
rect 33865 7855 33923 7889
rect 33957 7855 34015 7889
rect 34049 7855 34107 7889
rect 34141 7855 34199 7889
rect 34233 7855 34291 7889
rect 34325 7855 34383 7889
rect 34417 7855 34475 7889
rect 34509 7855 34567 7889
rect 34601 7855 34659 7889
rect 34693 7855 34751 7889
rect 34785 7855 34843 7889
rect 34877 7855 34935 7889
rect 34969 7855 35027 7889
rect 35061 7855 35119 7889
rect 35153 7855 35211 7889
rect 35245 7855 35303 7889
rect 35337 7855 35395 7889
rect 35429 7855 35487 7889
rect 35521 7855 35579 7889
rect 35613 7855 35671 7889
rect 35705 7855 36013 7889
rect 36047 7855 36076 7889
rect 33182 7836 36076 7855
rect 30210 7824 36076 7836
rect 34628 7782 34688 7788
rect 30666 7719 30724 7725
rect 30666 7685 30678 7719
rect 30712 7716 30724 7719
rect 31086 7719 31144 7725
rect 31086 7716 31098 7719
rect 30712 7688 31098 7716
rect 30712 7685 30724 7688
rect 30666 7679 30724 7685
rect 31086 7685 31098 7688
rect 31132 7716 31144 7719
rect 31400 7719 31458 7725
rect 31400 7716 31412 7719
rect 31132 7688 31412 7716
rect 31132 7685 31144 7688
rect 31086 7679 31144 7685
rect 31400 7685 31412 7688
rect 31446 7685 31458 7719
rect 31400 7679 31458 7685
rect 33364 7719 33422 7725
rect 33364 7685 33376 7719
rect 33410 7716 33422 7719
rect 33784 7719 33842 7725
rect 33784 7716 33796 7719
rect 33410 7688 33796 7716
rect 33410 7685 33422 7688
rect 33364 7679 33422 7685
rect 33784 7685 33796 7688
rect 33830 7716 33842 7719
rect 34098 7719 34156 7725
rect 34622 7722 34628 7782
rect 34688 7722 34694 7782
rect 34098 7716 34110 7719
rect 33830 7688 34110 7716
rect 33830 7685 33842 7688
rect 33784 7679 33842 7685
rect 34098 7685 34110 7688
rect 34144 7685 34156 7719
rect 34628 7716 34688 7722
rect 34098 7679 34156 7685
rect 30570 7650 30630 7656
rect 30745 7651 30803 7657
rect 30564 7590 30570 7650
rect 30630 7590 30636 7650
rect 30745 7617 30757 7651
rect 30791 7648 30803 7651
rect 30983 7651 31041 7657
rect 30983 7648 30995 7651
rect 30791 7620 30995 7648
rect 30791 7617 30803 7620
rect 30745 7611 30803 7617
rect 30983 7617 30995 7620
rect 31029 7648 31041 7651
rect 31487 7651 31545 7657
rect 31487 7648 31499 7651
rect 31029 7620 31499 7648
rect 31029 7617 31041 7620
rect 30983 7611 31041 7617
rect 31487 7617 31499 7620
rect 31533 7617 31545 7651
rect 31487 7611 31545 7617
rect 33443 7651 33501 7657
rect 33443 7617 33455 7651
rect 33489 7648 33501 7651
rect 33681 7651 33739 7657
rect 33681 7648 33693 7651
rect 33489 7620 33693 7648
rect 33489 7617 33501 7620
rect 33268 7610 33328 7616
rect 33443 7611 33501 7617
rect 33681 7617 33693 7620
rect 33727 7648 33739 7651
rect 34185 7651 34243 7657
rect 34185 7648 34197 7651
rect 33727 7620 34197 7648
rect 33727 7617 33739 7620
rect 33681 7611 33739 7617
rect 34185 7617 34197 7620
rect 34231 7617 34243 7651
rect 34185 7611 34243 7617
rect 32230 7592 32418 7598
rect 30570 7584 30630 7590
rect 30826 7560 30886 7566
rect 30820 7500 30826 7560
rect 30886 7500 30892 7560
rect 32230 7544 32242 7592
rect 32290 7544 32358 7592
rect 32406 7544 32418 7592
rect 32230 7538 32418 7544
rect 32458 7592 32888 7598
rect 32954 7596 33014 7602
rect 32458 7544 32470 7592
rect 32518 7544 32602 7592
rect 32650 7544 32712 7592
rect 32760 7544 32828 7592
rect 32876 7544 32888 7592
rect 32458 7538 32888 7544
rect 32948 7536 32954 7596
rect 33014 7536 33020 7596
rect 33262 7550 33268 7610
rect 33328 7550 33334 7610
rect 34928 7592 35116 7598
rect 33524 7560 33584 7566
rect 33268 7544 33328 7550
rect 32954 7530 33014 7536
rect 33518 7500 33524 7560
rect 33584 7500 33590 7560
rect 34928 7544 34940 7592
rect 34988 7544 35056 7592
rect 35104 7544 35116 7592
rect 34928 7538 35116 7544
rect 35156 7592 35586 7598
rect 35652 7596 35712 7602
rect 35156 7544 35168 7592
rect 35216 7544 35300 7592
rect 35348 7544 35410 7592
rect 35458 7544 35526 7592
rect 35574 7544 35586 7592
rect 35156 7538 35586 7544
rect 35646 7536 35652 7596
rect 35712 7536 35718 7596
rect 35652 7530 35712 7536
rect 30826 7494 30886 7500
rect 33524 7494 33584 7500
rect 31930 7478 31990 7484
rect 31924 7418 31930 7478
rect 31990 7418 31996 7478
rect 31930 7412 31990 7418
rect 30210 7364 36076 7376
rect 30210 7345 30406 7364
rect 30210 7311 30239 7345
rect 30273 7311 30406 7345
rect 30210 7292 30406 7311
rect 30502 7345 35784 7364
rect 30502 7311 30581 7345
rect 30615 7311 30673 7345
rect 30707 7311 30765 7345
rect 30799 7311 30857 7345
rect 30891 7311 30949 7345
rect 30983 7311 31041 7345
rect 31075 7311 31133 7345
rect 31167 7311 31225 7345
rect 31259 7311 31317 7345
rect 31351 7311 31409 7345
rect 31443 7311 31501 7345
rect 31535 7311 31593 7345
rect 31627 7311 31685 7345
rect 31719 7311 31777 7345
rect 31811 7311 31869 7345
rect 31903 7311 31961 7345
rect 31995 7311 32053 7345
rect 32087 7311 32145 7345
rect 32179 7311 32237 7345
rect 32271 7311 32329 7345
rect 32363 7311 32421 7345
rect 32455 7311 32513 7345
rect 32547 7311 32605 7345
rect 32639 7311 32697 7345
rect 32731 7311 32789 7345
rect 32823 7311 32881 7345
rect 32915 7311 32973 7345
rect 33007 7311 33279 7345
rect 33313 7311 33371 7345
rect 33405 7311 33463 7345
rect 33497 7311 33555 7345
rect 33589 7311 33647 7345
rect 33681 7311 33739 7345
rect 33773 7311 33831 7345
rect 33865 7311 33923 7345
rect 33957 7311 34015 7345
rect 34049 7311 34107 7345
rect 34141 7311 34199 7345
rect 34233 7311 34291 7345
rect 34325 7311 34383 7345
rect 34417 7311 34475 7345
rect 34509 7311 34567 7345
rect 34601 7311 34659 7345
rect 34693 7311 34751 7345
rect 34785 7311 34843 7345
rect 34877 7311 34935 7345
rect 34969 7311 35027 7345
rect 35061 7311 35119 7345
rect 35153 7311 35211 7345
rect 35245 7311 35303 7345
rect 35337 7311 35395 7345
rect 35429 7311 35487 7345
rect 35521 7311 35579 7345
rect 35613 7311 35671 7345
rect 35705 7311 35784 7345
rect 30502 7292 35784 7311
rect 35880 7345 36076 7364
rect 35880 7311 36013 7345
rect 36047 7311 36076 7345
rect 35880 7292 36076 7311
rect 30210 7280 36076 7292
rect 34628 7238 34688 7244
rect 34622 7178 34628 7238
rect 34688 7178 34694 7238
rect 34628 7172 34688 7178
rect 30826 7156 30886 7162
rect 33524 7156 33584 7162
rect 30570 7106 30630 7112
rect 30564 7046 30570 7106
rect 30630 7046 30636 7106
rect 30820 7096 30826 7156
rect 30886 7096 30892 7156
rect 32954 7120 33014 7126
rect 32230 7112 32418 7118
rect 30826 7090 30886 7096
rect 32230 7064 32242 7112
rect 32290 7064 32358 7112
rect 32406 7064 32418 7112
rect 32230 7058 32418 7064
rect 32458 7112 32888 7118
rect 32458 7064 32470 7112
rect 32518 7064 32602 7112
rect 32650 7064 32712 7112
rect 32760 7064 32828 7112
rect 32876 7064 32888 7112
rect 32458 7058 32888 7064
rect 32948 7060 32954 7120
rect 33014 7060 33020 7120
rect 33518 7096 33524 7156
rect 33584 7096 33590 7156
rect 35652 7120 35712 7126
rect 34928 7112 35116 7118
rect 33524 7090 33584 7096
rect 33268 7066 33328 7072
rect 32954 7054 33014 7060
rect 30570 7040 30630 7046
rect 30745 7039 30803 7045
rect 30745 7005 30757 7039
rect 30791 7036 30803 7039
rect 30983 7039 31041 7045
rect 30983 7036 30995 7039
rect 30791 7008 30995 7036
rect 30791 7005 30803 7008
rect 30745 6999 30803 7005
rect 30983 7005 30995 7008
rect 31029 7036 31041 7039
rect 31487 7039 31545 7045
rect 31487 7036 31499 7039
rect 31029 7008 31499 7036
rect 31029 7005 31041 7008
rect 30983 6999 31041 7005
rect 31487 7005 31499 7008
rect 31533 7005 31545 7039
rect 33262 7006 33268 7066
rect 33328 7006 33334 7066
rect 34928 7064 34940 7112
rect 34988 7064 35056 7112
rect 35104 7064 35116 7112
rect 34928 7058 35116 7064
rect 35156 7112 35586 7118
rect 35156 7064 35168 7112
rect 35216 7064 35300 7112
rect 35348 7064 35410 7112
rect 35458 7064 35526 7112
rect 35574 7064 35586 7112
rect 35156 7058 35586 7064
rect 35646 7060 35652 7120
rect 35712 7060 35718 7120
rect 35652 7054 35712 7060
rect 33443 7039 33501 7045
rect 31487 6999 31545 7005
rect 33268 7000 33328 7006
rect 33443 7005 33455 7039
rect 33489 7036 33501 7039
rect 33681 7039 33739 7045
rect 33681 7036 33693 7039
rect 33489 7008 33693 7036
rect 33489 7005 33501 7008
rect 33443 6999 33501 7005
rect 33681 7005 33693 7008
rect 33727 7036 33739 7039
rect 34185 7039 34243 7045
rect 34185 7036 34197 7039
rect 33727 7008 34197 7036
rect 33727 7005 33739 7008
rect 33681 6999 33739 7005
rect 34185 7005 34197 7008
rect 34231 7005 34243 7039
rect 34185 6999 34243 7005
rect 30666 6971 30724 6977
rect 30666 6937 30678 6971
rect 30712 6968 30724 6971
rect 31086 6971 31144 6977
rect 31086 6968 31098 6971
rect 30712 6940 31098 6968
rect 30712 6937 30724 6940
rect 30666 6931 30724 6937
rect 31086 6937 31098 6940
rect 31132 6968 31144 6971
rect 31400 6971 31458 6977
rect 31400 6968 31412 6971
rect 31132 6940 31412 6968
rect 31132 6937 31144 6940
rect 31086 6931 31144 6937
rect 31400 6937 31412 6940
rect 31446 6937 31458 6971
rect 33364 6971 33422 6977
rect 31400 6931 31458 6937
rect 31930 6934 31990 6940
rect 33364 6937 33376 6971
rect 33410 6968 33422 6971
rect 33784 6971 33842 6977
rect 33784 6968 33796 6971
rect 33410 6940 33796 6968
rect 33410 6937 33422 6940
rect 31924 6874 31930 6934
rect 31990 6874 31996 6934
rect 33364 6931 33422 6937
rect 33784 6937 33796 6940
rect 33830 6968 33842 6971
rect 34098 6971 34156 6977
rect 34098 6968 34110 6971
rect 33830 6940 34110 6968
rect 33830 6937 33842 6940
rect 33784 6931 33842 6937
rect 34098 6937 34110 6940
rect 34144 6937 34156 6971
rect 34098 6931 34156 6937
rect 31930 6868 31990 6874
rect 30210 6820 36076 6832
rect 30210 6801 33086 6820
rect 30210 6767 30239 6801
rect 30273 6767 30581 6801
rect 30615 6767 30673 6801
rect 30707 6767 30765 6801
rect 30799 6767 30857 6801
rect 30891 6767 30949 6801
rect 30983 6767 31041 6801
rect 31075 6767 31133 6801
rect 31167 6767 31225 6801
rect 31259 6767 31317 6801
rect 31351 6767 31409 6801
rect 31443 6767 31501 6801
rect 31535 6767 31593 6801
rect 31627 6767 31685 6801
rect 31719 6767 31777 6801
rect 31811 6767 31869 6801
rect 31903 6767 31961 6801
rect 31995 6767 32053 6801
rect 32087 6767 32145 6801
rect 32179 6767 32237 6801
rect 32271 6767 32329 6801
rect 32363 6767 32421 6801
rect 32455 6767 32513 6801
rect 32547 6767 32605 6801
rect 32639 6767 32697 6801
rect 32731 6767 32789 6801
rect 32823 6767 32881 6801
rect 32915 6767 32973 6801
rect 33007 6767 33086 6801
rect 30210 6748 33086 6767
rect 33182 6801 36076 6820
rect 33182 6767 33279 6801
rect 33313 6767 33371 6801
rect 33405 6767 33463 6801
rect 33497 6767 33555 6801
rect 33589 6767 33647 6801
rect 33681 6767 33739 6801
rect 33773 6767 33831 6801
rect 33865 6767 33923 6801
rect 33957 6767 34015 6801
rect 34049 6767 34107 6801
rect 34141 6767 34199 6801
rect 34233 6767 34291 6801
rect 34325 6767 34383 6801
rect 34417 6767 34475 6801
rect 34509 6767 34567 6801
rect 34601 6767 34659 6801
rect 34693 6767 34751 6801
rect 34785 6767 34843 6801
rect 34877 6767 34935 6801
rect 34969 6767 35027 6801
rect 35061 6767 35119 6801
rect 35153 6767 35211 6801
rect 35245 6767 35303 6801
rect 35337 6767 35395 6801
rect 35429 6767 35487 6801
rect 35521 6767 35579 6801
rect 35613 6767 35671 6801
rect 35705 6767 36013 6801
rect 36047 6767 36076 6801
rect 33182 6748 36076 6767
rect 30210 6736 36076 6748
rect 34628 6694 34688 6700
rect 30666 6631 30724 6637
rect 30666 6597 30678 6631
rect 30712 6628 30724 6631
rect 31086 6631 31144 6637
rect 31086 6628 31098 6631
rect 30712 6600 31098 6628
rect 30712 6597 30724 6600
rect 30666 6591 30724 6597
rect 31086 6597 31098 6600
rect 31132 6628 31144 6631
rect 31400 6631 31458 6637
rect 31400 6628 31412 6631
rect 31132 6600 31412 6628
rect 31132 6597 31144 6600
rect 31086 6591 31144 6597
rect 31400 6597 31412 6600
rect 31446 6597 31458 6631
rect 31400 6591 31458 6597
rect 33364 6631 33422 6637
rect 33364 6597 33376 6631
rect 33410 6628 33422 6631
rect 33784 6631 33842 6637
rect 33784 6628 33796 6631
rect 33410 6600 33796 6628
rect 33410 6597 33422 6600
rect 33364 6591 33422 6597
rect 33784 6597 33796 6600
rect 33830 6628 33842 6631
rect 34098 6631 34156 6637
rect 34622 6634 34628 6694
rect 34688 6634 34694 6694
rect 34098 6628 34110 6631
rect 33830 6600 34110 6628
rect 33830 6597 33842 6600
rect 33784 6591 33842 6597
rect 34098 6597 34110 6600
rect 34144 6597 34156 6631
rect 34628 6628 34688 6634
rect 34098 6591 34156 6597
rect 30570 6562 30630 6568
rect 30745 6563 30803 6569
rect 30564 6502 30570 6562
rect 30630 6502 30636 6562
rect 30745 6529 30757 6563
rect 30791 6560 30803 6563
rect 30983 6563 31041 6569
rect 30983 6560 30995 6563
rect 30791 6532 30995 6560
rect 30791 6529 30803 6532
rect 30745 6523 30803 6529
rect 30983 6529 30995 6532
rect 31029 6560 31041 6563
rect 31487 6563 31545 6569
rect 31487 6560 31499 6563
rect 31029 6532 31499 6560
rect 31029 6529 31041 6532
rect 30983 6523 31041 6529
rect 31487 6529 31499 6532
rect 31533 6529 31545 6563
rect 31487 6523 31545 6529
rect 33443 6563 33501 6569
rect 33443 6529 33455 6563
rect 33489 6560 33501 6563
rect 33681 6563 33739 6569
rect 33681 6560 33693 6563
rect 33489 6532 33693 6560
rect 33489 6529 33501 6532
rect 33268 6520 33328 6526
rect 33443 6523 33501 6529
rect 33681 6529 33693 6532
rect 33727 6560 33739 6563
rect 34185 6563 34243 6569
rect 34185 6560 34197 6563
rect 33727 6532 34197 6560
rect 33727 6529 33739 6532
rect 33681 6523 33739 6529
rect 34185 6529 34197 6532
rect 34231 6529 34243 6563
rect 34185 6523 34243 6529
rect 32230 6504 32418 6510
rect 30570 6496 30630 6502
rect 30826 6472 30886 6478
rect 30820 6412 30826 6472
rect 30886 6412 30892 6472
rect 32230 6456 32242 6504
rect 32290 6456 32358 6504
rect 32406 6456 32418 6504
rect 32230 6450 32418 6456
rect 32458 6504 32888 6510
rect 32954 6508 33014 6514
rect 32458 6456 32470 6504
rect 32518 6456 32602 6504
rect 32650 6456 32712 6504
rect 32760 6456 32828 6504
rect 32876 6456 32888 6504
rect 32458 6450 32888 6456
rect 32948 6448 32954 6508
rect 33014 6448 33020 6508
rect 33262 6460 33268 6520
rect 33328 6460 33334 6520
rect 34928 6504 35116 6510
rect 33524 6472 33584 6478
rect 33268 6454 33328 6460
rect 32954 6442 33014 6448
rect 33518 6412 33524 6472
rect 33584 6412 33590 6472
rect 34928 6456 34940 6504
rect 34988 6456 35056 6504
rect 35104 6456 35116 6504
rect 34928 6450 35116 6456
rect 35156 6504 35586 6510
rect 35156 6456 35168 6504
rect 35216 6456 35300 6504
rect 35348 6456 35410 6504
rect 35458 6456 35526 6504
rect 35574 6456 35586 6504
rect 35156 6450 35586 6456
rect 35644 6448 35650 6508
rect 35710 6448 35722 6508
rect 30826 6406 30886 6412
rect 33524 6406 33584 6412
rect 31930 6392 31990 6398
rect 31924 6332 31930 6392
rect 31990 6332 31996 6392
rect 31930 6326 31990 6332
rect 30210 6276 36076 6288
rect 30210 6257 30406 6276
rect 30210 6223 30239 6257
rect 30273 6223 30406 6257
rect 30210 6204 30406 6223
rect 30502 6257 35784 6276
rect 30502 6223 30581 6257
rect 30615 6223 30673 6257
rect 30707 6223 30765 6257
rect 30799 6223 30857 6257
rect 30891 6223 30949 6257
rect 30983 6223 31041 6257
rect 31075 6223 31133 6257
rect 31167 6223 31225 6257
rect 31259 6223 31317 6257
rect 31351 6223 31409 6257
rect 31443 6223 31501 6257
rect 31535 6223 31593 6257
rect 31627 6223 31685 6257
rect 31719 6223 31777 6257
rect 31811 6223 31869 6257
rect 31903 6223 31961 6257
rect 31995 6223 32053 6257
rect 32087 6223 32145 6257
rect 32179 6223 32237 6257
rect 32271 6223 32329 6257
rect 32363 6223 32421 6257
rect 32455 6223 32513 6257
rect 32547 6223 32605 6257
rect 32639 6223 32697 6257
rect 32731 6223 32789 6257
rect 32823 6223 32881 6257
rect 32915 6223 32973 6257
rect 33007 6223 33279 6257
rect 33313 6223 33371 6257
rect 33405 6223 33463 6257
rect 33497 6223 33555 6257
rect 33589 6223 33647 6257
rect 33681 6223 33739 6257
rect 33773 6223 33831 6257
rect 33865 6223 33923 6257
rect 33957 6223 34015 6257
rect 34049 6223 34107 6257
rect 34141 6223 34199 6257
rect 34233 6223 34291 6257
rect 34325 6223 34383 6257
rect 34417 6223 34475 6257
rect 34509 6223 34567 6257
rect 34601 6223 34659 6257
rect 34693 6223 34751 6257
rect 34785 6223 34843 6257
rect 34877 6223 34935 6257
rect 34969 6223 35027 6257
rect 35061 6223 35119 6257
rect 35153 6223 35211 6257
rect 35245 6223 35303 6257
rect 35337 6223 35395 6257
rect 35429 6223 35487 6257
rect 35521 6223 35579 6257
rect 35613 6223 35671 6257
rect 35705 6223 35784 6257
rect 30502 6204 35784 6223
rect 35880 6257 36076 6276
rect 35880 6223 36013 6257
rect 36047 6223 36076 6257
rect 35880 6204 36076 6223
rect 30210 6192 36076 6204
rect 34628 6148 34688 6154
rect 34622 6088 34628 6148
rect 34688 6088 34694 6148
rect 34628 6082 34688 6088
rect 30826 6068 30886 6074
rect 33524 6068 33584 6074
rect 30570 6020 30630 6026
rect 30564 5960 30570 6020
rect 30630 5960 30636 6020
rect 30820 6008 30826 6068
rect 30886 6008 30892 6068
rect 33276 6038 33336 6044
rect 32954 6032 33014 6038
rect 32230 6024 32418 6030
rect 30826 6002 30886 6008
rect 32230 5976 32242 6024
rect 32290 5976 32358 6024
rect 32406 5976 32418 6024
rect 32230 5970 32418 5976
rect 32458 6024 32888 6030
rect 32458 5976 32470 6024
rect 32518 5976 32602 6024
rect 32650 5976 32712 6024
rect 32760 5976 32828 6024
rect 32876 5976 32888 6024
rect 32458 5970 32888 5976
rect 32948 5972 32954 6032
rect 33014 5972 33020 6032
rect 33270 5978 33276 6038
rect 33336 5978 33342 6038
rect 33518 6008 33524 6068
rect 33584 6008 33590 6068
rect 35652 6032 35712 6038
rect 34928 6024 35116 6030
rect 33524 6002 33584 6008
rect 33276 5972 33336 5978
rect 34928 5976 34940 6024
rect 34988 5976 35056 6024
rect 35104 5976 35116 6024
rect 32954 5966 33014 5972
rect 34928 5970 35116 5976
rect 35156 6024 35586 6030
rect 35156 5976 35168 6024
rect 35216 5976 35300 6024
rect 35348 5976 35410 6024
rect 35458 5976 35526 6024
rect 35574 5976 35586 6024
rect 35156 5970 35586 5976
rect 35646 5972 35652 6032
rect 35712 5972 35718 6032
rect 35652 5966 35712 5972
rect 30570 5954 30630 5960
rect 30745 5951 30803 5957
rect 30745 5917 30757 5951
rect 30791 5948 30803 5951
rect 30983 5951 31041 5957
rect 30983 5948 30995 5951
rect 30791 5920 30995 5948
rect 30791 5917 30803 5920
rect 30745 5911 30803 5917
rect 30983 5917 30995 5920
rect 31029 5948 31041 5951
rect 31487 5951 31545 5957
rect 31487 5948 31499 5951
rect 31029 5920 31499 5948
rect 31029 5917 31041 5920
rect 30983 5911 31041 5917
rect 31487 5917 31499 5920
rect 31533 5917 31545 5951
rect 31487 5911 31545 5917
rect 33443 5951 33501 5957
rect 33443 5917 33455 5951
rect 33489 5948 33501 5951
rect 33681 5951 33739 5957
rect 33681 5948 33693 5951
rect 33489 5920 33693 5948
rect 33489 5917 33501 5920
rect 33443 5911 33501 5917
rect 33681 5917 33693 5920
rect 33727 5948 33739 5951
rect 34185 5951 34243 5957
rect 34185 5948 34197 5951
rect 33727 5920 34197 5948
rect 33727 5917 33739 5920
rect 33681 5911 33739 5917
rect 34185 5917 34197 5920
rect 34231 5917 34243 5951
rect 34185 5911 34243 5917
rect 30666 5883 30724 5889
rect 30666 5849 30678 5883
rect 30712 5880 30724 5883
rect 31086 5883 31144 5889
rect 31086 5880 31098 5883
rect 30712 5852 31098 5880
rect 30712 5849 30724 5852
rect 30666 5843 30724 5849
rect 31086 5849 31098 5852
rect 31132 5880 31144 5883
rect 31400 5883 31458 5889
rect 31400 5880 31412 5883
rect 31132 5852 31412 5880
rect 31132 5849 31144 5852
rect 31086 5843 31144 5849
rect 31400 5849 31412 5852
rect 31446 5849 31458 5883
rect 33364 5883 33422 5889
rect 31400 5843 31458 5849
rect 31930 5848 31990 5854
rect 33364 5849 33376 5883
rect 33410 5880 33422 5883
rect 33784 5883 33842 5889
rect 33784 5880 33796 5883
rect 33410 5852 33796 5880
rect 33410 5849 33422 5852
rect 31924 5788 31930 5848
rect 31990 5788 31996 5848
rect 33364 5843 33422 5849
rect 33784 5849 33796 5852
rect 33830 5880 33842 5883
rect 34098 5883 34156 5889
rect 34098 5880 34110 5883
rect 33830 5852 34110 5880
rect 33830 5849 33842 5852
rect 33784 5843 33842 5849
rect 34098 5849 34110 5852
rect 34144 5849 34156 5883
rect 34098 5843 34156 5849
rect 31930 5782 31990 5788
rect 30210 5732 36076 5744
rect 30210 5713 33086 5732
rect 30210 5679 30239 5713
rect 30273 5679 30581 5713
rect 30615 5679 30673 5713
rect 30707 5679 30765 5713
rect 30799 5679 30857 5713
rect 30891 5679 30949 5713
rect 30983 5679 31041 5713
rect 31075 5679 31133 5713
rect 31167 5679 31225 5713
rect 31259 5679 31317 5713
rect 31351 5679 31409 5713
rect 31443 5679 31501 5713
rect 31535 5679 31593 5713
rect 31627 5679 31685 5713
rect 31719 5679 31777 5713
rect 31811 5679 31869 5713
rect 31903 5679 31961 5713
rect 31995 5679 32053 5713
rect 32087 5679 32145 5713
rect 32179 5679 32237 5713
rect 32271 5679 32329 5713
rect 32363 5679 32421 5713
rect 32455 5679 32513 5713
rect 32547 5679 32605 5713
rect 32639 5679 32697 5713
rect 32731 5679 32789 5713
rect 32823 5679 32881 5713
rect 32915 5679 32973 5713
rect 33007 5679 33086 5713
rect 30210 5660 33086 5679
rect 33182 5713 36076 5732
rect 33182 5679 33279 5713
rect 33313 5679 33371 5713
rect 33405 5679 33463 5713
rect 33497 5679 33555 5713
rect 33589 5679 33647 5713
rect 33681 5679 33739 5713
rect 33773 5679 33831 5713
rect 33865 5679 33923 5713
rect 33957 5679 34015 5713
rect 34049 5679 34107 5713
rect 34141 5679 34199 5713
rect 34233 5679 34291 5713
rect 34325 5679 34383 5713
rect 34417 5679 34475 5713
rect 34509 5679 34567 5713
rect 34601 5679 34659 5713
rect 34693 5679 34751 5713
rect 34785 5679 34843 5713
rect 34877 5679 34935 5713
rect 34969 5679 35027 5713
rect 35061 5679 35119 5713
rect 35153 5679 35211 5713
rect 35245 5679 35303 5713
rect 35337 5679 35395 5713
rect 35429 5679 35487 5713
rect 35521 5679 35579 5713
rect 35613 5679 35671 5713
rect 35705 5679 36013 5713
rect 36047 5679 36076 5713
rect 33182 5660 36076 5679
rect 30210 5648 36076 5660
rect 28880 4872 28992 5049
rect 23536 4866 28992 4872
rect 23536 4766 23642 4866
rect 28886 4766 28992 4866
rect 23536 4760 28992 4766
rect 23346 4396 33802 4402
rect 23346 4296 23452 4396
rect 33696 4296 33802 4396
rect 23346 4290 33802 4296
rect 23346 4006 23458 4290
rect 23346 -1166 23352 4006
rect 23452 1184 23458 4006
rect 24058 3990 24068 4290
rect 33080 3990 33090 4290
rect 33690 4006 33802 4290
rect 24296 3816 32652 3830
rect 24296 3730 24310 3816
rect 24406 3730 24910 3816
rect 25006 3730 25510 3816
rect 25606 3730 26110 3816
rect 26206 3730 26710 3816
rect 26806 3730 27310 3816
rect 27406 3730 27910 3816
rect 28006 3730 28510 3816
rect 28606 3730 29110 3816
rect 29206 3730 29710 3816
rect 29806 3730 30310 3816
rect 30406 3730 30910 3816
rect 31006 3730 31510 3816
rect 31606 3730 32110 3816
rect 32206 3730 32530 3816
rect 32626 3730 32652 3816
rect 24296 3720 32652 3730
rect 24324 2932 24384 3720
rect 24556 3031 24616 3720
rect 24480 3025 24688 3031
rect 24480 2991 24492 3025
rect 24676 2991 24688 3025
rect 24480 2985 24688 2991
rect 24324 2900 24338 2932
rect 24332 1416 24338 2900
rect 24326 1356 24338 1416
rect 24372 2900 24384 2932
rect 24782 2932 24842 3720
rect 25698 3466 31256 3526
rect 25008 3098 25014 3158
rect 25074 3098 25080 3158
rect 25464 3098 25470 3158
rect 25530 3098 25536 3158
rect 25014 3031 25074 3098
rect 25470 3031 25530 3098
rect 24938 3025 25146 3031
rect 24938 2991 24950 3025
rect 25134 2991 25146 3025
rect 24938 2985 25146 2991
rect 25396 3025 25604 3031
rect 25396 2991 25408 3025
rect 25592 2991 25604 3025
rect 25396 2985 25604 2991
rect 24372 1416 24378 2900
rect 24782 2868 24796 2932
rect 24372 1356 24386 1416
rect 24790 1400 24796 2868
rect 24326 1184 24386 1356
rect 24780 1356 24796 1400
rect 24830 2868 24842 2932
rect 25248 2932 25294 2944
rect 24830 1400 24836 2868
rect 25248 1440 25254 2932
rect 24830 1356 24840 1400
rect 24480 1297 24688 1303
rect 24480 1263 24492 1297
rect 24676 1263 24688 1297
rect 24480 1257 24688 1263
rect 24554 1184 24614 1257
rect 24780 1184 24840 1356
rect 25238 1356 25254 1440
rect 25288 1440 25294 2932
rect 25698 2932 25758 3466
rect 26614 3332 30336 3392
rect 25924 3098 25930 3158
rect 25990 3098 25996 3158
rect 26380 3098 26386 3158
rect 26446 3098 26452 3158
rect 25930 3031 25990 3098
rect 26386 3031 26446 3098
rect 25854 3025 26062 3031
rect 25854 2991 25866 3025
rect 26050 2991 26062 3025
rect 25854 2985 26062 2991
rect 26312 3025 26520 3031
rect 26312 2991 26324 3025
rect 26508 2991 26520 3025
rect 26312 2985 26520 2991
rect 25698 2874 25712 2932
rect 25288 1356 25298 1440
rect 24938 1297 25146 1303
rect 24938 1263 24950 1297
rect 25134 1263 25146 1297
rect 24938 1257 25146 1263
rect 25010 1184 25070 1257
rect 23452 1124 24840 1184
rect 25004 1124 25010 1184
rect 25070 1124 25076 1184
rect 23452 752 23458 1124
rect 24326 752 24386 1124
rect 23452 692 24386 752
rect 25238 704 25298 1356
rect 25706 1356 25712 2874
rect 25746 2874 25758 2932
rect 26164 2932 26210 2944
rect 25746 1356 25752 2874
rect 26164 1434 26170 2932
rect 25706 1344 25752 1356
rect 26156 1356 26170 1434
rect 26204 1434 26210 2932
rect 26614 2932 26674 3332
rect 27530 3208 29420 3268
rect 26838 3098 26844 3158
rect 26904 3098 26910 3158
rect 27302 3098 27308 3158
rect 27368 3098 27374 3158
rect 26844 3031 26904 3098
rect 27308 3031 27368 3098
rect 26770 3025 26978 3031
rect 26770 2991 26782 3025
rect 26966 2991 26978 3025
rect 26770 2985 26978 2991
rect 27228 3025 27436 3031
rect 27228 2991 27240 3025
rect 27424 2991 27436 3025
rect 27228 2985 27436 2991
rect 26614 2872 26628 2932
rect 26204 1356 26216 1434
rect 25396 1297 25604 1303
rect 25396 1263 25408 1297
rect 25592 1263 25604 1297
rect 25396 1257 25604 1263
rect 25854 1297 26062 1303
rect 25854 1263 25866 1297
rect 26050 1263 26062 1297
rect 25854 1257 26062 1263
rect 25466 1184 25526 1257
rect 25926 1184 25986 1257
rect 25460 1124 25466 1184
rect 25526 1124 25532 1184
rect 25920 1124 25926 1184
rect 25986 1124 25992 1184
rect 26156 834 26216 1356
rect 26622 1356 26628 2872
rect 26662 2872 26674 2932
rect 27080 2932 27126 2944
rect 26662 1356 26668 2872
rect 27080 1428 27086 2932
rect 26622 1344 26668 1356
rect 27064 1356 27086 1428
rect 27120 1356 27126 2932
rect 27530 2932 27590 3208
rect 27752 3098 27758 3158
rect 27818 3098 27824 3158
rect 28208 3098 28214 3158
rect 28274 3098 28280 3158
rect 28676 3098 28682 3158
rect 28742 3098 28748 3158
rect 29134 3098 29140 3158
rect 29200 3098 29206 3158
rect 27758 3031 27818 3098
rect 28214 3031 28274 3098
rect 28682 3031 28742 3098
rect 29140 3031 29200 3098
rect 27686 3025 27894 3031
rect 27686 2991 27698 3025
rect 27882 2991 27894 3025
rect 27686 2985 27894 2991
rect 28144 3025 28352 3031
rect 28144 2991 28156 3025
rect 28340 2991 28352 3025
rect 28144 2985 28352 2991
rect 28602 3025 28810 3031
rect 28602 2991 28614 3025
rect 28798 2991 28810 3025
rect 28602 2985 28810 2991
rect 29060 3025 29268 3031
rect 29060 2991 29072 3025
rect 29256 2991 29268 3025
rect 29060 2985 29268 2991
rect 27530 2854 27544 2932
rect 27064 1344 27126 1356
rect 27538 1356 27544 2854
rect 27578 2854 27590 2932
rect 27996 2932 28042 2944
rect 27578 1356 27584 2854
rect 27996 1436 28002 2932
rect 27538 1344 27584 1356
rect 27988 1356 28002 1436
rect 28036 1436 28042 2932
rect 28454 2932 28500 2944
rect 28036 1356 28048 1436
rect 28454 1378 28460 2932
rect 26312 1297 26520 1303
rect 26312 1263 26324 1297
rect 26508 1263 26520 1297
rect 26312 1257 26520 1263
rect 26770 1297 26978 1303
rect 26770 1263 26782 1297
rect 26966 1263 26978 1297
rect 26770 1257 26978 1263
rect 26382 1184 26442 1257
rect 26840 1184 26900 1257
rect 26376 1124 26382 1184
rect 26442 1124 26448 1184
rect 26834 1124 26840 1184
rect 26900 1124 26906 1184
rect 27064 960 27124 1344
rect 27228 1297 27436 1303
rect 27228 1263 27240 1297
rect 27424 1263 27436 1297
rect 27228 1257 27436 1263
rect 27686 1297 27894 1303
rect 27686 1263 27698 1297
rect 27882 1263 27894 1297
rect 27686 1257 27894 1263
rect 27304 1184 27364 1257
rect 27758 1184 27818 1257
rect 27298 1124 27304 1184
rect 27364 1124 27370 1184
rect 27752 1124 27758 1184
rect 27818 1124 27824 1184
rect 27988 1076 28048 1356
rect 28450 1356 28460 1378
rect 28494 1378 28500 2932
rect 28912 2932 28958 2944
rect 28912 1384 28918 2932
rect 28494 1356 28510 1378
rect 28144 1297 28352 1303
rect 28144 1263 28156 1297
rect 28340 1263 28352 1297
rect 28144 1257 28352 1263
rect 28216 1186 28276 1257
rect 28450 1196 28510 1356
rect 28906 1356 28918 1384
rect 28952 1384 28958 2932
rect 29360 2932 29420 3208
rect 29590 3098 29596 3158
rect 29656 3098 29662 3158
rect 30046 3098 30052 3158
rect 30112 3098 30118 3158
rect 29596 3031 29656 3098
rect 30052 3031 30112 3098
rect 29518 3025 29726 3031
rect 29518 2991 29530 3025
rect 29714 2991 29726 3025
rect 29518 2985 29726 2991
rect 29976 3025 30184 3031
rect 29976 2991 29988 3025
rect 30172 2991 30184 3025
rect 29976 2985 30184 2991
rect 29360 2888 29376 2932
rect 28952 1356 28966 1384
rect 28602 1297 28810 1303
rect 28602 1263 28614 1297
rect 28798 1263 28810 1297
rect 28602 1257 28810 1263
rect 28210 1184 28282 1186
rect 28210 1124 28216 1184
rect 28276 1124 28282 1184
rect 28676 1192 28736 1257
rect 28450 1130 28510 1136
rect 28664 1186 28748 1192
rect 28664 1124 28676 1186
rect 28736 1124 28748 1186
rect 28664 1120 28748 1124
rect 28906 1076 28966 1356
rect 29370 1356 29376 2888
rect 29410 2888 29420 2932
rect 29828 2932 29874 2944
rect 29410 1356 29416 2888
rect 29828 1388 29834 2932
rect 29370 1344 29416 1356
rect 29820 1356 29834 1388
rect 29868 1388 29874 2932
rect 30276 2932 30336 3332
rect 30502 3098 30508 3158
rect 30568 3098 30574 3158
rect 30958 3098 30964 3158
rect 31024 3098 31030 3158
rect 30508 3031 30568 3098
rect 30964 3031 31024 3098
rect 30434 3025 30642 3031
rect 30434 2991 30446 3025
rect 30630 2991 30642 3025
rect 30434 2985 30642 2991
rect 30892 3025 31100 3031
rect 30892 2991 30904 3025
rect 31088 2991 31100 3025
rect 30892 2985 31100 2991
rect 30276 2874 30292 2932
rect 29868 1356 29880 1388
rect 29060 1297 29268 1303
rect 29060 1263 29072 1297
rect 29256 1263 29268 1297
rect 29060 1257 29268 1263
rect 29518 1297 29726 1303
rect 29518 1263 29530 1297
rect 29714 1263 29726 1297
rect 29518 1257 29726 1263
rect 29132 1184 29192 1257
rect 29592 1184 29652 1257
rect 29126 1124 29132 1184
rect 29192 1124 29198 1184
rect 29586 1124 29592 1184
rect 29652 1124 29658 1184
rect 27988 1016 28966 1076
rect 29820 960 29880 1356
rect 30286 1356 30292 2874
rect 30326 2874 30336 2932
rect 30744 2932 30790 2944
rect 30326 1356 30332 2874
rect 30744 1424 30750 2932
rect 30286 1344 30332 1356
rect 30740 1356 30750 1424
rect 30784 1424 30790 2932
rect 31196 2932 31256 3466
rect 31416 3098 31422 3158
rect 31482 3098 31488 3158
rect 31876 3098 31882 3158
rect 31942 3098 31948 3158
rect 31422 3031 31482 3098
rect 31882 3031 31942 3098
rect 31350 3025 31558 3031
rect 31350 2991 31362 3025
rect 31546 2991 31558 3025
rect 31350 2985 31558 2991
rect 31808 3025 32016 3031
rect 31808 2991 31820 3025
rect 32004 2991 32016 3025
rect 31808 2985 32016 2991
rect 31196 2876 31208 2932
rect 30784 1356 30800 1424
rect 29976 1297 30184 1303
rect 29976 1263 29988 1297
rect 30172 1263 30184 1297
rect 29976 1257 30184 1263
rect 30434 1297 30642 1303
rect 30434 1263 30446 1297
rect 30630 1263 30642 1297
rect 30434 1257 30642 1263
rect 30048 1184 30108 1257
rect 30504 1184 30564 1257
rect 30042 1124 30048 1184
rect 30108 1124 30114 1184
rect 30498 1124 30504 1184
rect 30564 1124 30570 1184
rect 27064 900 29880 960
rect 30740 834 30800 1356
rect 31202 1356 31208 2876
rect 31242 2876 31256 2932
rect 31660 2932 31706 2944
rect 31242 1356 31248 2876
rect 31660 1416 31666 2932
rect 31202 1344 31248 1356
rect 31654 1356 31666 1416
rect 31700 1416 31706 2932
rect 32112 2932 32172 3720
rect 32342 3031 32402 3720
rect 32266 3025 32474 3031
rect 32266 2991 32278 3025
rect 32462 2991 32474 3025
rect 32266 2985 32474 2991
rect 32112 2856 32124 2932
rect 32118 1418 32124 2856
rect 31700 1356 31714 1416
rect 30892 1297 31100 1303
rect 30892 1263 30904 1297
rect 31088 1263 31100 1297
rect 30892 1257 31100 1263
rect 31350 1297 31558 1303
rect 31350 1263 31362 1297
rect 31546 1263 31558 1297
rect 31350 1257 31558 1263
rect 30960 1184 31020 1257
rect 31418 1184 31478 1257
rect 30954 1124 30960 1184
rect 31020 1124 31026 1184
rect 31412 1124 31418 1184
rect 31478 1124 31484 1184
rect 26156 774 30800 834
rect 31654 704 31714 1356
rect 32108 1356 32124 1418
rect 32158 2856 32172 2932
rect 32570 2932 32630 3720
rect 32570 2862 32582 2932
rect 32158 1418 32164 2856
rect 32158 1356 32168 1418
rect 32576 1400 32582 2862
rect 31808 1297 32016 1303
rect 31808 1263 31820 1297
rect 32004 1263 32016 1297
rect 31808 1257 32016 1263
rect 31878 1184 31938 1257
rect 31872 1124 31878 1184
rect 31938 1124 31944 1184
rect 32108 1182 32168 1356
rect 32566 1356 32582 1400
rect 32616 2862 32630 2932
rect 32616 1400 32622 2862
rect 32616 1356 32626 1400
rect 32266 1297 32474 1303
rect 32266 1263 32278 1297
rect 32462 1263 32474 1297
rect 32266 1257 32474 1263
rect 32340 1182 32400 1257
rect 32566 1182 32626 1356
rect 33690 1182 33696 4006
rect 32108 1122 33696 1182
rect 23452 -1166 23458 692
rect 23766 267 23826 692
rect 23994 366 24054 692
rect 25238 644 31714 704
rect 32566 688 32626 1122
rect 33690 688 33696 1122
rect 32566 628 33696 688
rect 24218 538 24224 598
rect 24284 538 24290 598
rect 23921 360 24129 366
rect 23921 326 23933 360
rect 24117 326 24129 360
rect 23921 320 24129 326
rect 23766 220 23779 267
rect 23773 -888 23779 220
rect 23346 -1342 23458 -1166
rect 23766 -909 23779 -888
rect 23813 220 23826 267
rect 24224 267 24284 538
rect 24456 436 27720 496
rect 24456 366 24516 436
rect 24918 366 24978 436
rect 25372 366 25432 436
rect 25834 366 25894 436
rect 26288 366 26348 436
rect 26738 366 26798 436
rect 27204 366 27264 436
rect 27660 366 27720 436
rect 28116 418 29284 478
rect 28116 366 28176 418
rect 24379 360 24587 366
rect 24379 326 24391 360
rect 24575 326 24587 360
rect 24379 320 24587 326
rect 24837 360 25045 366
rect 24837 326 24849 360
rect 25033 326 25045 360
rect 24837 320 25045 326
rect 25295 360 25503 366
rect 25295 326 25307 360
rect 25491 326 25503 360
rect 25295 320 25503 326
rect 25753 360 25961 366
rect 25753 326 25765 360
rect 25949 326 25961 360
rect 25753 320 25961 326
rect 26211 360 26419 366
rect 26211 326 26223 360
rect 26407 326 26419 360
rect 26211 320 26419 326
rect 26669 360 26877 366
rect 26669 326 26681 360
rect 26865 326 26877 360
rect 26669 320 26877 326
rect 27127 360 27335 366
rect 27127 326 27139 360
rect 27323 326 27335 360
rect 27127 320 27335 326
rect 27585 360 27793 366
rect 27585 326 27597 360
rect 27781 326 27793 360
rect 27585 320 27793 326
rect 28043 360 28251 366
rect 28043 326 28055 360
rect 28239 326 28251 360
rect 28043 320 28251 326
rect 23813 -888 23819 220
rect 24224 200 24237 267
rect 23813 -909 23826 -888
rect 23766 -1342 23826 -909
rect 24231 -909 24237 200
rect 24271 200 24284 267
rect 24689 267 24735 279
rect 24271 -909 24277 200
rect 24231 -921 24277 -909
rect 24689 -909 24695 267
rect 24729 -909 24735 267
rect 24689 -921 24735 -909
rect 25147 267 25193 279
rect 25147 -909 25153 267
rect 25187 -909 25193 267
rect 25147 -921 25193 -909
rect 25605 267 25651 279
rect 25605 -909 25611 267
rect 25645 -909 25651 267
rect 25605 -921 25651 -909
rect 26063 267 26109 279
rect 26063 -909 26069 267
rect 26103 -909 26109 267
rect 26063 -921 26109 -909
rect 26521 267 26567 279
rect 26521 -909 26527 267
rect 26561 -909 26567 267
rect 26521 -921 26567 -909
rect 26979 267 27025 279
rect 26979 -909 26985 267
rect 27019 -909 27025 267
rect 26979 -921 27025 -909
rect 27437 267 27483 279
rect 27437 -909 27443 267
rect 27477 -909 27483 267
rect 27895 267 27941 279
rect 27895 -842 27901 267
rect 27437 -921 27483 -909
rect 27886 -909 27901 -842
rect 27935 -842 27941 267
rect 28346 267 28406 418
rect 28346 252 28359 267
rect 27935 -909 27946 -842
rect 28353 -874 28359 252
rect 23921 -968 24129 -962
rect 23921 -1002 23933 -968
rect 24117 -1002 24129 -968
rect 23921 -1008 24129 -1002
rect 24379 -968 24587 -962
rect 24379 -1002 24391 -968
rect 24575 -1002 24587 -968
rect 24379 -1008 24587 -1002
rect 24837 -968 25045 -962
rect 24837 -1002 24849 -968
rect 25033 -1002 25045 -968
rect 24837 -1008 25045 -1002
rect 25295 -968 25503 -962
rect 25295 -1002 25307 -968
rect 25491 -1002 25503 -968
rect 25295 -1008 25503 -1002
rect 25753 -968 25961 -962
rect 25753 -1002 25765 -968
rect 25949 -1002 25961 -968
rect 25753 -1008 25961 -1002
rect 26211 -968 26419 -962
rect 26211 -1002 26223 -968
rect 26407 -1002 26419 -968
rect 26211 -1008 26419 -1002
rect 26669 -968 26877 -962
rect 26669 -1002 26681 -968
rect 26865 -1002 26877 -968
rect 26669 -1008 26877 -1002
rect 27127 -968 27335 -962
rect 27127 -1002 27139 -968
rect 27323 -1002 27335 -968
rect 27127 -1008 27335 -1002
rect 27585 -968 27793 -962
rect 27585 -1002 27597 -968
rect 27781 -1002 27793 -968
rect 27585 -1008 27793 -1002
rect 23994 -1342 24054 -1008
rect 24448 -1076 24508 -1008
rect 24910 -1076 24970 -1008
rect 25364 -1076 25424 -1008
rect 25826 -1076 25886 -1008
rect 26280 -1076 26340 -1008
rect 26730 -1076 26790 -1008
rect 27196 -1076 27256 -1008
rect 27652 -1076 27712 -1008
rect 24448 -1080 25364 -1076
rect 24508 -1136 24910 -1080
rect 24448 -1146 24508 -1140
rect 24970 -1136 25364 -1080
rect 25424 -1136 25826 -1076
rect 25886 -1082 26730 -1076
rect 25886 -1136 26280 -1082
rect 24910 -1146 24970 -1140
rect 25364 -1142 25424 -1136
rect 25826 -1142 25886 -1136
rect 26340 -1136 26730 -1082
rect 26790 -1136 27196 -1076
rect 27256 -1080 27712 -1076
rect 27256 -1136 27652 -1080
rect 26730 -1142 26790 -1136
rect 27196 -1142 27256 -1136
rect 26280 -1148 26340 -1142
rect 27652 -1146 27712 -1140
rect 27886 -1202 27946 -909
rect 28344 -909 28359 -874
rect 28393 252 28406 267
rect 28766 267 28826 418
rect 28998 366 29058 418
rect 28921 360 29129 366
rect 28921 326 28933 360
rect 29117 326 29129 360
rect 28921 320 29129 326
rect 28393 -874 28399 252
rect 28766 246 28779 267
rect 28773 -874 28779 246
rect 28393 -909 28404 -874
rect 28043 -968 28251 -962
rect 28043 -1002 28055 -968
rect 28239 -1002 28251 -968
rect 28043 -1008 28251 -1002
rect 27880 -1262 27886 -1202
rect 27946 -1262 27952 -1202
rect 28116 -1342 28176 -1008
rect 28344 -1342 28404 -909
rect 28764 -909 28779 -874
rect 28813 246 28826 267
rect 29224 267 29284 418
rect 29450 436 32714 496
rect 29450 366 29510 436
rect 29912 366 29972 436
rect 30366 366 30426 436
rect 30828 366 30888 436
rect 31282 366 31342 436
rect 31732 366 31792 436
rect 32198 366 32258 436
rect 32654 366 32714 436
rect 33116 366 33176 628
rect 29379 360 29587 366
rect 29379 326 29391 360
rect 29575 326 29587 360
rect 29379 320 29587 326
rect 29837 360 30045 366
rect 29837 326 29849 360
rect 30033 326 30045 360
rect 29837 320 30045 326
rect 30295 360 30503 366
rect 30295 326 30307 360
rect 30491 326 30503 360
rect 30295 320 30503 326
rect 30753 360 30961 366
rect 30753 326 30765 360
rect 30949 326 30961 360
rect 30753 320 30961 326
rect 31211 360 31419 366
rect 31211 326 31223 360
rect 31407 326 31419 360
rect 31211 320 31419 326
rect 31669 360 31877 366
rect 31669 326 31681 360
rect 31865 326 31877 360
rect 31669 320 31877 326
rect 32127 360 32335 366
rect 32127 326 32139 360
rect 32323 326 32335 360
rect 32127 320 32335 326
rect 32585 360 32793 366
rect 32585 326 32597 360
rect 32781 326 32793 360
rect 32585 320 32793 326
rect 33043 360 33251 366
rect 33043 326 33055 360
rect 33239 326 33251 360
rect 33043 320 33251 326
rect 28813 -874 28819 246
rect 29224 224 29237 267
rect 29231 -868 29237 224
rect 28813 -909 28824 -874
rect 28764 -1342 28824 -909
rect 29222 -909 29237 -868
rect 29271 224 29284 267
rect 29689 267 29735 279
rect 29271 -868 29277 224
rect 29271 -909 29282 -868
rect 28921 -968 29129 -962
rect 28921 -1002 28933 -968
rect 29117 -1002 29129 -968
rect 28921 -1008 29129 -1002
rect 28992 -1342 29052 -1008
rect 29222 -1342 29282 -909
rect 29689 -909 29695 267
rect 29729 -909 29735 267
rect 29689 -921 29735 -909
rect 30147 267 30193 279
rect 30147 -909 30153 267
rect 30187 -909 30193 267
rect 30147 -921 30193 -909
rect 30605 267 30651 279
rect 30605 -909 30611 267
rect 30645 -909 30651 267
rect 30605 -921 30651 -909
rect 31063 267 31109 279
rect 31063 -909 31069 267
rect 31103 -909 31109 267
rect 31063 -921 31109 -909
rect 31521 267 31567 279
rect 31521 -909 31527 267
rect 31561 -909 31567 267
rect 31521 -921 31567 -909
rect 31979 267 32025 279
rect 31979 -909 31985 267
rect 32019 -909 32025 267
rect 31979 -921 32025 -909
rect 32437 267 32483 279
rect 32437 -909 32443 267
rect 32477 -909 32483 267
rect 32895 267 32941 279
rect 32895 -902 32901 267
rect 32437 -921 32483 -909
rect 32886 -909 32901 -902
rect 32935 -902 32941 267
rect 33342 267 33402 628
rect 33342 214 33359 267
rect 33353 -876 33359 214
rect 32935 -909 32946 -902
rect 29379 -968 29587 -962
rect 29379 -1002 29391 -968
rect 29575 -1002 29587 -968
rect 29379 -1008 29587 -1002
rect 29837 -968 30045 -962
rect 29837 -1002 29849 -968
rect 30033 -1002 30045 -968
rect 29837 -1008 30045 -1002
rect 30295 -968 30503 -962
rect 30295 -1002 30307 -968
rect 30491 -1002 30503 -968
rect 30295 -1008 30503 -1002
rect 30753 -968 30961 -962
rect 30753 -1002 30765 -968
rect 30949 -1002 30961 -968
rect 30753 -1008 30961 -1002
rect 31211 -968 31419 -962
rect 31211 -1002 31223 -968
rect 31407 -1002 31419 -968
rect 31211 -1008 31419 -1002
rect 31669 -968 31877 -962
rect 31669 -1002 31681 -968
rect 31865 -1002 31877 -968
rect 31669 -1008 31877 -1002
rect 32127 -968 32335 -962
rect 32127 -1002 32139 -968
rect 32323 -1002 32335 -968
rect 32127 -1008 32335 -1002
rect 32585 -968 32793 -962
rect 32585 -1002 32597 -968
rect 32781 -1002 32793 -968
rect 32585 -1008 32793 -1002
rect 29450 -1076 29510 -1008
rect 29912 -1072 29972 -1008
rect 29450 -1080 29912 -1076
rect 29510 -1132 29912 -1080
rect 30366 -1076 30426 -1008
rect 30828 -1076 30888 -1008
rect 31282 -1076 31342 -1008
rect 31732 -1072 31792 -1008
rect 29972 -1078 31732 -1076
rect 29972 -1132 30366 -1078
rect 29510 -1136 30366 -1132
rect 29912 -1138 29972 -1136
rect 30426 -1136 30828 -1078
rect 29450 -1146 29510 -1140
rect 30366 -1144 30426 -1138
rect 30888 -1136 31282 -1078
rect 30828 -1144 30888 -1138
rect 31342 -1132 31732 -1078
rect 32198 -1076 32258 -1008
rect 32654 -1076 32714 -1008
rect 31792 -1078 32714 -1076
rect 31792 -1132 32198 -1078
rect 31342 -1136 32198 -1132
rect 31732 -1138 31792 -1136
rect 32258 -1136 32654 -1078
rect 31282 -1144 31342 -1138
rect 32198 -1144 32258 -1138
rect 32654 -1144 32714 -1138
rect 32886 -1208 32946 -909
rect 33344 -909 33359 -876
rect 33393 214 33402 267
rect 33393 -876 33399 214
rect 33393 -909 33404 -876
rect 33043 -968 33251 -962
rect 33043 -1002 33055 -968
rect 33239 -1002 33251 -968
rect 33043 -1008 33251 -1002
rect 32886 -1274 32946 -1268
rect 33116 -1342 33176 -1008
rect 33344 -1342 33404 -909
rect 33690 -1166 33696 628
rect 33796 -1166 33802 4006
rect 33690 -1342 33802 -1166
rect 23346 -1348 33802 -1342
rect 23346 -1448 23452 -1348
rect 33696 -1448 33802 -1348
rect 23346 -1454 33802 -1448
rect 23346 -1684 33802 -1678
rect 23346 -1784 23452 -1684
rect 33696 -1784 33802 -1684
rect 23346 -1790 33802 -1784
rect 23346 -1914 23458 -1790
rect 23074 -3286 23080 -3226
rect 23140 -3286 23146 -3226
rect 8346 -13604 18802 -13598
rect 8346 -13704 8452 -13604
rect 18696 -13704 18802 -13604
rect 8346 -13710 18802 -13704
rect 8346 -13994 8458 -13710
rect 8346 -19166 8352 -13994
rect 8452 -16816 8458 -13994
rect 9058 -14010 9068 -13710
rect 18080 -14010 18090 -13710
rect 18690 -13994 18802 -13710
rect 9296 -14184 17652 -14170
rect 9296 -14270 9310 -14184
rect 9406 -14270 9910 -14184
rect 10006 -14270 10510 -14184
rect 10606 -14270 11110 -14184
rect 11206 -14270 11710 -14184
rect 11806 -14270 12310 -14184
rect 12406 -14270 12910 -14184
rect 13006 -14270 13510 -14184
rect 13606 -14270 14110 -14184
rect 14206 -14270 14710 -14184
rect 14806 -14270 15310 -14184
rect 15406 -14270 15910 -14184
rect 16006 -14270 16510 -14184
rect 16606 -14270 17110 -14184
rect 17206 -14270 17530 -14184
rect 17626 -14270 17652 -14184
rect 9296 -14280 17652 -14270
rect 9324 -15068 9384 -14280
rect 9556 -14969 9616 -14280
rect 9480 -14975 9688 -14969
rect 9480 -15009 9492 -14975
rect 9676 -15009 9688 -14975
rect 9480 -15015 9688 -15009
rect 9324 -15100 9338 -15068
rect 9332 -16584 9338 -15100
rect 9326 -16644 9338 -16584
rect 9372 -15100 9384 -15068
rect 9782 -15068 9842 -14280
rect 10698 -14534 16256 -14474
rect 10008 -14902 10014 -14842
rect 10074 -14902 10080 -14842
rect 10464 -14902 10470 -14842
rect 10530 -14902 10536 -14842
rect 10014 -14969 10074 -14902
rect 10470 -14969 10530 -14902
rect 9938 -14975 10146 -14969
rect 9938 -15009 9950 -14975
rect 10134 -15009 10146 -14975
rect 9938 -15015 10146 -15009
rect 10396 -14975 10604 -14969
rect 10396 -15009 10408 -14975
rect 10592 -15009 10604 -14975
rect 10396 -15015 10604 -15009
rect 9372 -16584 9378 -15100
rect 9782 -15132 9796 -15068
rect 9372 -16644 9386 -16584
rect 9790 -16600 9796 -15132
rect 9326 -16816 9386 -16644
rect 9780 -16644 9796 -16600
rect 9830 -15132 9842 -15068
rect 10248 -15068 10294 -15056
rect 9830 -16600 9836 -15132
rect 10248 -16560 10254 -15068
rect 9830 -16644 9840 -16600
rect 9480 -16703 9688 -16697
rect 9480 -16737 9492 -16703
rect 9676 -16737 9688 -16703
rect 9480 -16743 9688 -16737
rect 9554 -16816 9614 -16743
rect 9780 -16816 9840 -16644
rect 10238 -16644 10254 -16560
rect 10288 -16560 10294 -15068
rect 10698 -15068 10758 -14534
rect 11614 -14668 15336 -14608
rect 10924 -14902 10930 -14842
rect 10990 -14902 10996 -14842
rect 11380 -14902 11386 -14842
rect 11446 -14902 11452 -14842
rect 10930 -14969 10990 -14902
rect 11386 -14969 11446 -14902
rect 10854 -14975 11062 -14969
rect 10854 -15009 10866 -14975
rect 11050 -15009 11062 -14975
rect 10854 -15015 11062 -15009
rect 11312 -14975 11520 -14969
rect 11312 -15009 11324 -14975
rect 11508 -15009 11520 -14975
rect 11312 -15015 11520 -15009
rect 10698 -15126 10712 -15068
rect 10288 -16644 10298 -16560
rect 9938 -16703 10146 -16697
rect 9938 -16737 9950 -16703
rect 10134 -16737 10146 -16703
rect 9938 -16743 10146 -16737
rect 10010 -16816 10070 -16743
rect 8452 -16876 9840 -16816
rect 10004 -16876 10010 -16816
rect 10070 -16876 10076 -16816
rect 8452 -17248 8458 -16876
rect 9326 -17248 9386 -16876
rect 8452 -17308 9386 -17248
rect 10238 -17296 10298 -16644
rect 10706 -16644 10712 -15126
rect 10746 -15126 10758 -15068
rect 11164 -15068 11210 -15056
rect 10746 -16644 10752 -15126
rect 11164 -16566 11170 -15068
rect 10706 -16656 10752 -16644
rect 11156 -16644 11170 -16566
rect 11204 -16566 11210 -15068
rect 11614 -15068 11674 -14668
rect 12530 -14792 14420 -14732
rect 11838 -14902 11844 -14842
rect 11904 -14902 11910 -14842
rect 12302 -14902 12308 -14842
rect 12368 -14902 12374 -14842
rect 11844 -14969 11904 -14902
rect 12308 -14969 12368 -14902
rect 11770 -14975 11978 -14969
rect 11770 -15009 11782 -14975
rect 11966 -15009 11978 -14975
rect 11770 -15015 11978 -15009
rect 12228 -14975 12436 -14969
rect 12228 -15009 12240 -14975
rect 12424 -15009 12436 -14975
rect 12228 -15015 12436 -15009
rect 11614 -15128 11628 -15068
rect 11204 -16644 11216 -16566
rect 10396 -16703 10604 -16697
rect 10396 -16737 10408 -16703
rect 10592 -16737 10604 -16703
rect 10396 -16743 10604 -16737
rect 10854 -16703 11062 -16697
rect 10854 -16737 10866 -16703
rect 11050 -16737 11062 -16703
rect 10854 -16743 11062 -16737
rect 10466 -16816 10526 -16743
rect 10926 -16816 10986 -16743
rect 10460 -16876 10466 -16816
rect 10526 -16876 10532 -16816
rect 10920 -16876 10926 -16816
rect 10986 -16876 10992 -16816
rect 11156 -17166 11216 -16644
rect 11622 -16644 11628 -15128
rect 11662 -15128 11674 -15068
rect 12080 -15068 12126 -15056
rect 11662 -16644 11668 -15128
rect 12080 -16572 12086 -15068
rect 11622 -16656 11668 -16644
rect 12064 -16644 12086 -16572
rect 12120 -16644 12126 -15068
rect 12530 -15068 12590 -14792
rect 12752 -14902 12758 -14842
rect 12818 -14902 12824 -14842
rect 13208 -14902 13214 -14842
rect 13274 -14902 13280 -14842
rect 13676 -14902 13682 -14842
rect 13742 -14902 13748 -14842
rect 14134 -14902 14140 -14842
rect 14200 -14902 14206 -14842
rect 12758 -14969 12818 -14902
rect 13214 -14969 13274 -14902
rect 13682 -14969 13742 -14902
rect 14140 -14969 14200 -14902
rect 12686 -14975 12894 -14969
rect 12686 -15009 12698 -14975
rect 12882 -15009 12894 -14975
rect 12686 -15015 12894 -15009
rect 13144 -14975 13352 -14969
rect 13144 -15009 13156 -14975
rect 13340 -15009 13352 -14975
rect 13144 -15015 13352 -15009
rect 13602 -14975 13810 -14969
rect 13602 -15009 13614 -14975
rect 13798 -15009 13810 -14975
rect 13602 -15015 13810 -15009
rect 14060 -14975 14268 -14969
rect 14060 -15009 14072 -14975
rect 14256 -15009 14268 -14975
rect 14060 -15015 14268 -15009
rect 12530 -15146 12544 -15068
rect 12064 -16656 12126 -16644
rect 12538 -16644 12544 -15146
rect 12578 -15146 12590 -15068
rect 12996 -15068 13042 -15056
rect 12578 -16644 12584 -15146
rect 12996 -16564 13002 -15068
rect 12538 -16656 12584 -16644
rect 12988 -16644 13002 -16564
rect 13036 -16564 13042 -15068
rect 13454 -15068 13500 -15056
rect 13036 -16644 13048 -16564
rect 13454 -16622 13460 -15068
rect 11312 -16703 11520 -16697
rect 11312 -16737 11324 -16703
rect 11508 -16737 11520 -16703
rect 11312 -16743 11520 -16737
rect 11770 -16703 11978 -16697
rect 11770 -16737 11782 -16703
rect 11966 -16737 11978 -16703
rect 11770 -16743 11978 -16737
rect 11382 -16816 11442 -16743
rect 11840 -16816 11900 -16743
rect 11376 -16876 11382 -16816
rect 11442 -16876 11448 -16816
rect 11834 -16876 11840 -16816
rect 11900 -16876 11906 -16816
rect 12064 -17040 12124 -16656
rect 12228 -16703 12436 -16697
rect 12228 -16737 12240 -16703
rect 12424 -16737 12436 -16703
rect 12228 -16743 12436 -16737
rect 12686 -16703 12894 -16697
rect 12686 -16737 12698 -16703
rect 12882 -16737 12894 -16703
rect 12686 -16743 12894 -16737
rect 12304 -16816 12364 -16743
rect 12758 -16816 12818 -16743
rect 12298 -16876 12304 -16816
rect 12364 -16876 12370 -16816
rect 12752 -16876 12758 -16816
rect 12818 -16876 12824 -16816
rect 12988 -16924 13048 -16644
rect 13450 -16644 13460 -16622
rect 13494 -16622 13500 -15068
rect 13912 -15068 13958 -15056
rect 13912 -16616 13918 -15068
rect 13494 -16644 13510 -16622
rect 13144 -16703 13352 -16697
rect 13144 -16737 13156 -16703
rect 13340 -16737 13352 -16703
rect 13144 -16743 13352 -16737
rect 13216 -16814 13276 -16743
rect 13450 -16804 13510 -16644
rect 13906 -16644 13918 -16616
rect 13952 -16616 13958 -15068
rect 14360 -15068 14420 -14792
rect 14590 -14902 14596 -14842
rect 14656 -14902 14662 -14842
rect 15046 -14902 15052 -14842
rect 15112 -14902 15118 -14842
rect 14596 -14969 14656 -14902
rect 15052 -14969 15112 -14902
rect 14518 -14975 14726 -14969
rect 14518 -15009 14530 -14975
rect 14714 -15009 14726 -14975
rect 14518 -15015 14726 -15009
rect 14976 -14975 15184 -14969
rect 14976 -15009 14988 -14975
rect 15172 -15009 15184 -14975
rect 14976 -15015 15184 -15009
rect 14360 -15112 14376 -15068
rect 13952 -16644 13966 -16616
rect 13602 -16703 13810 -16697
rect 13602 -16737 13614 -16703
rect 13798 -16737 13810 -16703
rect 13602 -16743 13810 -16737
rect 13210 -16816 13282 -16814
rect 13210 -16876 13216 -16816
rect 13276 -16876 13282 -16816
rect 13676 -16808 13736 -16743
rect 13450 -16870 13510 -16864
rect 13664 -16814 13748 -16808
rect 13664 -16876 13676 -16814
rect 13736 -16876 13748 -16814
rect 13664 -16880 13748 -16876
rect 13906 -16924 13966 -16644
rect 14370 -16644 14376 -15112
rect 14410 -15112 14420 -15068
rect 14828 -15068 14874 -15056
rect 14410 -16644 14416 -15112
rect 14828 -16612 14834 -15068
rect 14370 -16656 14416 -16644
rect 14820 -16644 14834 -16612
rect 14868 -16612 14874 -15068
rect 15276 -15068 15336 -14668
rect 15502 -14902 15508 -14842
rect 15568 -14902 15574 -14842
rect 15958 -14902 15964 -14842
rect 16024 -14902 16030 -14842
rect 15508 -14969 15568 -14902
rect 15964 -14969 16024 -14902
rect 15434 -14975 15642 -14969
rect 15434 -15009 15446 -14975
rect 15630 -15009 15642 -14975
rect 15434 -15015 15642 -15009
rect 15892 -14975 16100 -14969
rect 15892 -15009 15904 -14975
rect 16088 -15009 16100 -14975
rect 15892 -15015 16100 -15009
rect 15276 -15126 15292 -15068
rect 14868 -16644 14880 -16612
rect 14060 -16703 14268 -16697
rect 14060 -16737 14072 -16703
rect 14256 -16737 14268 -16703
rect 14060 -16743 14268 -16737
rect 14518 -16703 14726 -16697
rect 14518 -16737 14530 -16703
rect 14714 -16737 14726 -16703
rect 14518 -16743 14726 -16737
rect 14132 -16816 14192 -16743
rect 14592 -16816 14652 -16743
rect 14126 -16876 14132 -16816
rect 14192 -16876 14198 -16816
rect 14586 -16876 14592 -16816
rect 14652 -16876 14658 -16816
rect 12988 -16984 13966 -16924
rect 14820 -17040 14880 -16644
rect 15286 -16644 15292 -15126
rect 15326 -15126 15336 -15068
rect 15744 -15068 15790 -15056
rect 15326 -16644 15332 -15126
rect 15744 -16576 15750 -15068
rect 15286 -16656 15332 -16644
rect 15740 -16644 15750 -16576
rect 15784 -16576 15790 -15068
rect 16196 -15068 16256 -14534
rect 16416 -14902 16422 -14842
rect 16482 -14902 16488 -14842
rect 16876 -14902 16882 -14842
rect 16942 -14902 16948 -14842
rect 16422 -14969 16482 -14902
rect 16882 -14969 16942 -14902
rect 16350 -14975 16558 -14969
rect 16350 -15009 16362 -14975
rect 16546 -15009 16558 -14975
rect 16350 -15015 16558 -15009
rect 16808 -14975 17016 -14969
rect 16808 -15009 16820 -14975
rect 17004 -15009 17016 -14975
rect 16808 -15015 17016 -15009
rect 16196 -15124 16208 -15068
rect 15784 -16644 15800 -16576
rect 14976 -16703 15184 -16697
rect 14976 -16737 14988 -16703
rect 15172 -16737 15184 -16703
rect 14976 -16743 15184 -16737
rect 15434 -16703 15642 -16697
rect 15434 -16737 15446 -16703
rect 15630 -16737 15642 -16703
rect 15434 -16743 15642 -16737
rect 15048 -16816 15108 -16743
rect 15504 -16816 15564 -16743
rect 15042 -16876 15048 -16816
rect 15108 -16876 15114 -16816
rect 15498 -16876 15504 -16816
rect 15564 -16876 15570 -16816
rect 12064 -17100 14880 -17040
rect 15740 -17166 15800 -16644
rect 16202 -16644 16208 -15124
rect 16242 -15124 16256 -15068
rect 16660 -15068 16706 -15056
rect 16242 -16644 16248 -15124
rect 16660 -16584 16666 -15068
rect 16202 -16656 16248 -16644
rect 16654 -16644 16666 -16584
rect 16700 -16584 16706 -15068
rect 17112 -15068 17172 -14280
rect 17342 -14969 17402 -14280
rect 17266 -14975 17474 -14969
rect 17266 -15009 17278 -14975
rect 17462 -15009 17474 -14975
rect 17266 -15015 17474 -15009
rect 17112 -15144 17124 -15068
rect 17118 -16582 17124 -15144
rect 16700 -16644 16714 -16584
rect 15892 -16703 16100 -16697
rect 15892 -16737 15904 -16703
rect 16088 -16737 16100 -16703
rect 15892 -16743 16100 -16737
rect 16350 -16703 16558 -16697
rect 16350 -16737 16362 -16703
rect 16546 -16737 16558 -16703
rect 16350 -16743 16558 -16737
rect 15960 -16816 16020 -16743
rect 16418 -16816 16478 -16743
rect 15954 -16876 15960 -16816
rect 16020 -16876 16026 -16816
rect 16412 -16876 16418 -16816
rect 16478 -16876 16484 -16816
rect 11156 -17226 15800 -17166
rect 16654 -17296 16714 -16644
rect 17108 -16644 17124 -16582
rect 17158 -15144 17172 -15068
rect 17570 -15068 17630 -14280
rect 17570 -15138 17582 -15068
rect 17158 -16582 17164 -15144
rect 17158 -16644 17168 -16582
rect 17576 -16600 17582 -15138
rect 16808 -16703 17016 -16697
rect 16808 -16737 16820 -16703
rect 17004 -16737 17016 -16703
rect 16808 -16743 17016 -16737
rect 16878 -16816 16938 -16743
rect 16872 -16876 16878 -16816
rect 16938 -16876 16944 -16816
rect 17108 -16818 17168 -16644
rect 17566 -16644 17582 -16600
rect 17616 -15138 17630 -15068
rect 17616 -16600 17622 -15138
rect 17616 -16644 17626 -16600
rect 17266 -16703 17474 -16697
rect 17266 -16737 17278 -16703
rect 17462 -16737 17474 -16703
rect 17266 -16743 17474 -16737
rect 17340 -16818 17400 -16743
rect 17566 -16818 17626 -16644
rect 18690 -16818 18696 -13994
rect 17108 -16878 18696 -16818
rect 8452 -19166 8458 -17308
rect 8766 -17733 8826 -17308
rect 8994 -17634 9054 -17308
rect 10238 -17356 16714 -17296
rect 17566 -17312 17626 -16878
rect 18690 -17312 18696 -16878
rect 17566 -17372 18696 -17312
rect 9218 -17462 9224 -17402
rect 9284 -17462 9290 -17402
rect 8921 -17640 9129 -17634
rect 8921 -17674 8933 -17640
rect 9117 -17674 9129 -17640
rect 8921 -17680 9129 -17674
rect 8766 -17780 8779 -17733
rect 8773 -18888 8779 -17780
rect 8346 -19342 8458 -19166
rect 8766 -18909 8779 -18888
rect 8813 -17780 8826 -17733
rect 9224 -17733 9284 -17462
rect 9456 -17564 12720 -17504
rect 9456 -17634 9516 -17564
rect 9918 -17634 9978 -17564
rect 10372 -17634 10432 -17564
rect 10834 -17634 10894 -17564
rect 11288 -17634 11348 -17564
rect 11738 -17634 11798 -17564
rect 12204 -17634 12264 -17564
rect 12660 -17634 12720 -17564
rect 13116 -17582 14284 -17522
rect 13116 -17634 13176 -17582
rect 9379 -17640 9587 -17634
rect 9379 -17674 9391 -17640
rect 9575 -17674 9587 -17640
rect 9379 -17680 9587 -17674
rect 9837 -17640 10045 -17634
rect 9837 -17674 9849 -17640
rect 10033 -17674 10045 -17640
rect 9837 -17680 10045 -17674
rect 10295 -17640 10503 -17634
rect 10295 -17674 10307 -17640
rect 10491 -17674 10503 -17640
rect 10295 -17680 10503 -17674
rect 10753 -17640 10961 -17634
rect 10753 -17674 10765 -17640
rect 10949 -17674 10961 -17640
rect 10753 -17680 10961 -17674
rect 11211 -17640 11419 -17634
rect 11211 -17674 11223 -17640
rect 11407 -17674 11419 -17640
rect 11211 -17680 11419 -17674
rect 11669 -17640 11877 -17634
rect 11669 -17674 11681 -17640
rect 11865 -17674 11877 -17640
rect 11669 -17680 11877 -17674
rect 12127 -17640 12335 -17634
rect 12127 -17674 12139 -17640
rect 12323 -17674 12335 -17640
rect 12127 -17680 12335 -17674
rect 12585 -17640 12793 -17634
rect 12585 -17674 12597 -17640
rect 12781 -17674 12793 -17640
rect 12585 -17680 12793 -17674
rect 13043 -17640 13251 -17634
rect 13043 -17674 13055 -17640
rect 13239 -17674 13251 -17640
rect 13043 -17680 13251 -17674
rect 8813 -18888 8819 -17780
rect 9224 -17800 9237 -17733
rect 8813 -18909 8826 -18888
rect 8766 -19342 8826 -18909
rect 9231 -18909 9237 -17800
rect 9271 -17800 9284 -17733
rect 9689 -17733 9735 -17721
rect 9271 -18909 9277 -17800
rect 9231 -18921 9277 -18909
rect 9689 -18909 9695 -17733
rect 9729 -18909 9735 -17733
rect 9689 -18921 9735 -18909
rect 10147 -17733 10193 -17721
rect 10147 -18909 10153 -17733
rect 10187 -18909 10193 -17733
rect 10147 -18921 10193 -18909
rect 10605 -17733 10651 -17721
rect 10605 -18909 10611 -17733
rect 10645 -18909 10651 -17733
rect 10605 -18921 10651 -18909
rect 11063 -17733 11109 -17721
rect 11063 -18909 11069 -17733
rect 11103 -18909 11109 -17733
rect 11063 -18921 11109 -18909
rect 11521 -17733 11567 -17721
rect 11521 -18909 11527 -17733
rect 11561 -18909 11567 -17733
rect 11521 -18921 11567 -18909
rect 11979 -17733 12025 -17721
rect 11979 -18909 11985 -17733
rect 12019 -18909 12025 -17733
rect 11979 -18921 12025 -18909
rect 12437 -17733 12483 -17721
rect 12437 -18909 12443 -17733
rect 12477 -18909 12483 -17733
rect 12895 -17733 12941 -17721
rect 12895 -18842 12901 -17733
rect 12437 -18921 12483 -18909
rect 12886 -18909 12901 -18842
rect 12935 -18842 12941 -17733
rect 13346 -17733 13406 -17582
rect 13346 -17748 13359 -17733
rect 12935 -18909 12946 -18842
rect 13353 -18874 13359 -17748
rect 8921 -18968 9129 -18962
rect 8921 -19002 8933 -18968
rect 9117 -19002 9129 -18968
rect 8921 -19008 9129 -19002
rect 9379 -18968 9587 -18962
rect 9379 -19002 9391 -18968
rect 9575 -19002 9587 -18968
rect 9379 -19008 9587 -19002
rect 9837 -18968 10045 -18962
rect 9837 -19002 9849 -18968
rect 10033 -19002 10045 -18968
rect 9837 -19008 10045 -19002
rect 10295 -18968 10503 -18962
rect 10295 -19002 10307 -18968
rect 10491 -19002 10503 -18968
rect 10295 -19008 10503 -19002
rect 10753 -18968 10961 -18962
rect 10753 -19002 10765 -18968
rect 10949 -19002 10961 -18968
rect 10753 -19008 10961 -19002
rect 11211 -18968 11419 -18962
rect 11211 -19002 11223 -18968
rect 11407 -19002 11419 -18968
rect 11211 -19008 11419 -19002
rect 11669 -18968 11877 -18962
rect 11669 -19002 11681 -18968
rect 11865 -19002 11877 -18968
rect 11669 -19008 11877 -19002
rect 12127 -18968 12335 -18962
rect 12127 -19002 12139 -18968
rect 12323 -19002 12335 -18968
rect 12127 -19008 12335 -19002
rect 12585 -18968 12793 -18962
rect 12585 -19002 12597 -18968
rect 12781 -19002 12793 -18968
rect 12585 -19008 12793 -19002
rect 8994 -19342 9054 -19008
rect 9448 -19076 9508 -19008
rect 9910 -19076 9970 -19008
rect 10364 -19076 10424 -19008
rect 10826 -19076 10886 -19008
rect 11280 -19076 11340 -19008
rect 11730 -19076 11790 -19008
rect 12196 -19076 12256 -19008
rect 12652 -19076 12712 -19008
rect 9448 -19080 10364 -19076
rect 9508 -19136 9910 -19080
rect 9448 -19146 9508 -19140
rect 9970 -19136 10364 -19080
rect 10424 -19136 10826 -19076
rect 10886 -19082 11730 -19076
rect 10886 -19136 11280 -19082
rect 9910 -19146 9970 -19140
rect 10364 -19142 10424 -19136
rect 10826 -19142 10886 -19136
rect 11340 -19136 11730 -19082
rect 11790 -19136 12196 -19076
rect 12256 -19080 12712 -19076
rect 12256 -19136 12652 -19080
rect 11730 -19142 11790 -19136
rect 12196 -19142 12256 -19136
rect 11280 -19148 11340 -19142
rect 12652 -19146 12712 -19140
rect 12886 -19202 12946 -18909
rect 13344 -18909 13359 -18874
rect 13393 -17748 13406 -17733
rect 13766 -17733 13826 -17582
rect 13998 -17634 14058 -17582
rect 13921 -17640 14129 -17634
rect 13921 -17674 13933 -17640
rect 14117 -17674 14129 -17640
rect 13921 -17680 14129 -17674
rect 13393 -18874 13399 -17748
rect 13766 -17754 13779 -17733
rect 13773 -18874 13779 -17754
rect 13393 -18909 13404 -18874
rect 13043 -18968 13251 -18962
rect 13043 -19002 13055 -18968
rect 13239 -19002 13251 -18968
rect 13043 -19008 13251 -19002
rect 12880 -19262 12886 -19202
rect 12946 -19262 12952 -19202
rect 13116 -19342 13176 -19008
rect 13344 -19342 13404 -18909
rect 13764 -18909 13779 -18874
rect 13813 -17754 13826 -17733
rect 14224 -17733 14284 -17582
rect 14450 -17564 17714 -17504
rect 14450 -17634 14510 -17564
rect 14912 -17634 14972 -17564
rect 15366 -17634 15426 -17564
rect 15828 -17634 15888 -17564
rect 16282 -17634 16342 -17564
rect 16732 -17634 16792 -17564
rect 17198 -17634 17258 -17564
rect 17654 -17634 17714 -17564
rect 18116 -17634 18176 -17372
rect 14379 -17640 14587 -17634
rect 14379 -17674 14391 -17640
rect 14575 -17674 14587 -17640
rect 14379 -17680 14587 -17674
rect 14837 -17640 15045 -17634
rect 14837 -17674 14849 -17640
rect 15033 -17674 15045 -17640
rect 14837 -17680 15045 -17674
rect 15295 -17640 15503 -17634
rect 15295 -17674 15307 -17640
rect 15491 -17674 15503 -17640
rect 15295 -17680 15503 -17674
rect 15753 -17640 15961 -17634
rect 15753 -17674 15765 -17640
rect 15949 -17674 15961 -17640
rect 15753 -17680 15961 -17674
rect 16211 -17640 16419 -17634
rect 16211 -17674 16223 -17640
rect 16407 -17674 16419 -17640
rect 16211 -17680 16419 -17674
rect 16669 -17640 16877 -17634
rect 16669 -17674 16681 -17640
rect 16865 -17674 16877 -17640
rect 16669 -17680 16877 -17674
rect 17127 -17640 17335 -17634
rect 17127 -17674 17139 -17640
rect 17323 -17674 17335 -17640
rect 17127 -17680 17335 -17674
rect 17585 -17640 17793 -17634
rect 17585 -17674 17597 -17640
rect 17781 -17674 17793 -17640
rect 17585 -17680 17793 -17674
rect 18043 -17640 18251 -17634
rect 18043 -17674 18055 -17640
rect 18239 -17674 18251 -17640
rect 18043 -17680 18251 -17674
rect 13813 -18874 13819 -17754
rect 14224 -17776 14237 -17733
rect 14231 -18868 14237 -17776
rect 13813 -18909 13824 -18874
rect 13764 -19342 13824 -18909
rect 14222 -18909 14237 -18868
rect 14271 -17776 14284 -17733
rect 14689 -17733 14735 -17721
rect 14271 -18868 14277 -17776
rect 14271 -18909 14282 -18868
rect 13921 -18968 14129 -18962
rect 13921 -19002 13933 -18968
rect 14117 -19002 14129 -18968
rect 13921 -19008 14129 -19002
rect 13992 -19342 14052 -19008
rect 14222 -19342 14282 -18909
rect 14689 -18909 14695 -17733
rect 14729 -18909 14735 -17733
rect 14689 -18921 14735 -18909
rect 15147 -17733 15193 -17721
rect 15147 -18909 15153 -17733
rect 15187 -18909 15193 -17733
rect 15147 -18921 15193 -18909
rect 15605 -17733 15651 -17721
rect 15605 -18909 15611 -17733
rect 15645 -18909 15651 -17733
rect 15605 -18921 15651 -18909
rect 16063 -17733 16109 -17721
rect 16063 -18909 16069 -17733
rect 16103 -18909 16109 -17733
rect 16063 -18921 16109 -18909
rect 16521 -17733 16567 -17721
rect 16521 -18909 16527 -17733
rect 16561 -18909 16567 -17733
rect 16521 -18921 16567 -18909
rect 16979 -17733 17025 -17721
rect 16979 -18909 16985 -17733
rect 17019 -18909 17025 -17733
rect 16979 -18921 17025 -18909
rect 17437 -17733 17483 -17721
rect 17437 -18909 17443 -17733
rect 17477 -18909 17483 -17733
rect 17895 -17733 17941 -17721
rect 17895 -18902 17901 -17733
rect 17437 -18921 17483 -18909
rect 17886 -18909 17901 -18902
rect 17935 -18902 17941 -17733
rect 18342 -17733 18402 -17372
rect 18342 -17786 18359 -17733
rect 18353 -18876 18359 -17786
rect 17935 -18909 17946 -18902
rect 14379 -18968 14587 -18962
rect 14379 -19002 14391 -18968
rect 14575 -19002 14587 -18968
rect 14379 -19008 14587 -19002
rect 14837 -18968 15045 -18962
rect 14837 -19002 14849 -18968
rect 15033 -19002 15045 -18968
rect 14837 -19008 15045 -19002
rect 15295 -18968 15503 -18962
rect 15295 -19002 15307 -18968
rect 15491 -19002 15503 -18968
rect 15295 -19008 15503 -19002
rect 15753 -18968 15961 -18962
rect 15753 -19002 15765 -18968
rect 15949 -19002 15961 -18968
rect 15753 -19008 15961 -19002
rect 16211 -18968 16419 -18962
rect 16211 -19002 16223 -18968
rect 16407 -19002 16419 -18968
rect 16211 -19008 16419 -19002
rect 16669 -18968 16877 -18962
rect 16669 -19002 16681 -18968
rect 16865 -19002 16877 -18968
rect 16669 -19008 16877 -19002
rect 17127 -18968 17335 -18962
rect 17127 -19002 17139 -18968
rect 17323 -19002 17335 -18968
rect 17127 -19008 17335 -19002
rect 17585 -18968 17793 -18962
rect 17585 -19002 17597 -18968
rect 17781 -19002 17793 -18968
rect 17585 -19008 17793 -19002
rect 14450 -19076 14510 -19008
rect 14912 -19072 14972 -19008
rect 14450 -19080 14912 -19076
rect 14510 -19132 14912 -19080
rect 15366 -19076 15426 -19008
rect 15828 -19076 15888 -19008
rect 16282 -19076 16342 -19008
rect 16732 -19072 16792 -19008
rect 14972 -19078 16732 -19076
rect 14972 -19132 15366 -19078
rect 14510 -19136 15366 -19132
rect 14912 -19138 14972 -19136
rect 15426 -19136 15828 -19078
rect 14450 -19146 14510 -19140
rect 15366 -19144 15426 -19138
rect 15888 -19136 16282 -19078
rect 15828 -19144 15888 -19138
rect 16342 -19132 16732 -19078
rect 17198 -19076 17258 -19008
rect 17654 -19076 17714 -19008
rect 16792 -19078 17714 -19076
rect 16792 -19132 17198 -19078
rect 16342 -19136 17198 -19132
rect 16732 -19138 16792 -19136
rect 17258 -19136 17654 -19078
rect 16282 -19144 16342 -19138
rect 17198 -19144 17258 -19138
rect 17654 -19144 17714 -19138
rect 17886 -19208 17946 -18909
rect 18344 -18909 18359 -18876
rect 18393 -17786 18402 -17733
rect 18393 -18876 18399 -17786
rect 18393 -18909 18404 -18876
rect 18043 -18968 18251 -18962
rect 18043 -19002 18055 -18968
rect 18239 -19002 18251 -18968
rect 18043 -19008 18251 -19002
rect 17886 -19274 17946 -19268
rect 18116 -19342 18176 -19008
rect 18344 -19342 18404 -18909
rect 18690 -19166 18696 -17372
rect 18796 -19166 18802 -13994
rect 22940 -16816 23000 -9940
rect 23080 -5470 23140 -3286
rect 23346 -3918 23352 -1914
rect 23452 -3918 23458 -1914
rect 23766 -2226 23826 -1790
rect 23996 -2136 24056 -1790
rect 27886 -1882 27946 -1876
rect 24454 -2016 24910 -2010
rect 24442 -2076 24448 -2016
rect 24508 -2070 24910 -2016
rect 24970 -2016 25826 -2010
rect 24970 -2070 25364 -2016
rect 24508 -2076 24514 -2070
rect 24448 -2136 24514 -2076
rect 24910 -2136 24976 -2070
rect 25358 -2076 25364 -2070
rect 25424 -2070 25826 -2016
rect 25886 -2070 26280 -2010
rect 26340 -2070 26730 -2010
rect 26790 -2016 27652 -2010
rect 26790 -2070 27196 -2016
rect 25424 -2076 25430 -2070
rect 25364 -2136 25430 -2076
rect 25826 -2136 25892 -2070
rect 26280 -2136 26346 -2070
rect 26730 -2136 26796 -2070
rect 27190 -2076 27196 -2070
rect 27256 -2070 27652 -2016
rect 27712 -2070 27718 -2010
rect 27256 -2076 27262 -2070
rect 27196 -2136 27262 -2076
rect 27652 -2136 27718 -2070
rect 23920 -2142 24128 -2136
rect 23920 -2176 23932 -2142
rect 24116 -2176 24128 -2142
rect 23920 -2182 24128 -2176
rect 24378 -2142 24586 -2136
rect 24378 -2176 24390 -2142
rect 24574 -2176 24586 -2142
rect 24378 -2182 24586 -2176
rect 24836 -2142 25044 -2136
rect 24836 -2176 24848 -2142
rect 25032 -2176 25044 -2142
rect 24836 -2182 25044 -2176
rect 25294 -2142 25502 -2136
rect 25294 -2176 25306 -2142
rect 25490 -2176 25502 -2142
rect 25294 -2182 25502 -2176
rect 25752 -2142 25960 -2136
rect 25752 -2176 25764 -2142
rect 25948 -2176 25960 -2142
rect 25752 -2182 25960 -2176
rect 26210 -2142 26418 -2136
rect 26210 -2176 26222 -2142
rect 26406 -2176 26418 -2142
rect 26210 -2182 26418 -2176
rect 26668 -2142 26876 -2136
rect 26668 -2176 26680 -2142
rect 26864 -2176 26876 -2142
rect 26668 -2182 26876 -2176
rect 27126 -2142 27334 -2136
rect 27126 -2176 27138 -2142
rect 27322 -2176 27334 -2142
rect 27126 -2182 27334 -2176
rect 27584 -2142 27792 -2136
rect 27584 -2176 27596 -2142
rect 27780 -2176 27792 -2142
rect 27584 -2182 27792 -2176
rect 23766 -2266 23778 -2226
rect 23772 -2362 23778 -2266
rect 23766 -2402 23778 -2362
rect 23812 -2266 23826 -2226
rect 24230 -2226 24276 -2214
rect 23812 -2362 23818 -2266
rect 24230 -2360 24236 -2226
rect 23812 -2402 23826 -2362
rect 23766 -2618 23826 -2402
rect 24222 -2402 24236 -2360
rect 24270 -2360 24276 -2226
rect 24688 -2226 24734 -2214
rect 24270 -2402 24282 -2360
rect 23920 -2452 24128 -2446
rect 23920 -2486 23932 -2452
rect 24116 -2486 24128 -2452
rect 23920 -2492 24128 -2486
rect 23994 -2618 24054 -2492
rect 23766 -2678 24054 -2618
rect 23766 -2894 23826 -2678
rect 23994 -2804 24054 -2678
rect 23920 -2810 24128 -2804
rect 23920 -2844 23932 -2810
rect 24116 -2844 24128 -2810
rect 23920 -2850 24128 -2844
rect 23766 -2914 23778 -2894
rect 23772 -3040 23778 -2914
rect 23758 -3070 23778 -3040
rect 23812 -2914 23826 -2894
rect 24222 -2894 24282 -2402
rect 24688 -2402 24694 -2226
rect 24728 -2402 24734 -2226
rect 24688 -2414 24734 -2402
rect 25146 -2226 25192 -2214
rect 25146 -2402 25152 -2226
rect 25186 -2402 25192 -2226
rect 25146 -2414 25192 -2402
rect 25604 -2226 25650 -2214
rect 25604 -2402 25610 -2226
rect 25644 -2402 25650 -2226
rect 25604 -2414 25650 -2402
rect 26062 -2226 26108 -2214
rect 26062 -2402 26068 -2226
rect 26102 -2402 26108 -2226
rect 26062 -2414 26108 -2402
rect 26520 -2226 26566 -2214
rect 26520 -2402 26526 -2226
rect 26560 -2402 26566 -2226
rect 26520 -2414 26566 -2402
rect 26978 -2226 27024 -2214
rect 26978 -2402 26984 -2226
rect 27018 -2402 27024 -2226
rect 26978 -2414 27024 -2402
rect 27436 -2226 27482 -2214
rect 27436 -2402 27442 -2226
rect 27476 -2402 27482 -2226
rect 27886 -2226 27946 -1942
rect 28114 -2136 28174 -1790
rect 28042 -2142 28250 -2136
rect 28042 -2176 28054 -2142
rect 28238 -2176 28250 -2142
rect 28042 -2182 28250 -2176
rect 27886 -2256 27900 -2226
rect 27436 -2414 27482 -2402
rect 27894 -2402 27900 -2256
rect 27934 -2256 27946 -2226
rect 28346 -2226 28406 -1790
rect 28346 -2254 28358 -2226
rect 27934 -2402 27940 -2256
rect 28352 -2346 28358 -2254
rect 27894 -2414 27940 -2402
rect 28346 -2402 28358 -2346
rect 28392 -2254 28406 -2226
rect 28766 -2226 28826 -1790
rect 29000 -2136 29060 -1790
rect 28920 -2142 29128 -2136
rect 28920 -2176 28932 -2142
rect 29116 -2176 29128 -2142
rect 28920 -2182 29128 -2176
rect 28392 -2346 28398 -2254
rect 28766 -2262 28778 -2226
rect 28392 -2402 28406 -2346
rect 28772 -2366 28778 -2262
rect 24378 -2452 24586 -2446
rect 24378 -2486 24390 -2452
rect 24574 -2486 24586 -2452
rect 24378 -2492 24586 -2486
rect 24836 -2452 25044 -2446
rect 24836 -2486 24848 -2452
rect 25032 -2486 25044 -2452
rect 24836 -2492 25044 -2486
rect 25294 -2452 25502 -2446
rect 25294 -2486 25306 -2452
rect 25490 -2486 25502 -2452
rect 25294 -2492 25502 -2486
rect 25752 -2452 25960 -2446
rect 25752 -2486 25764 -2452
rect 25948 -2486 25960 -2452
rect 25752 -2492 25960 -2486
rect 26210 -2452 26418 -2446
rect 26210 -2486 26222 -2452
rect 26406 -2486 26418 -2452
rect 26210 -2492 26418 -2486
rect 26668 -2452 26876 -2446
rect 26668 -2486 26680 -2452
rect 26864 -2486 26876 -2452
rect 26668 -2492 26876 -2486
rect 27126 -2452 27334 -2446
rect 27126 -2486 27138 -2452
rect 27322 -2486 27334 -2452
rect 27126 -2492 27334 -2486
rect 27584 -2452 27792 -2446
rect 27584 -2486 27596 -2452
rect 27780 -2486 27792 -2452
rect 27584 -2492 27792 -2486
rect 28042 -2452 28250 -2446
rect 28042 -2486 28054 -2452
rect 28238 -2486 28250 -2452
rect 28042 -2492 28250 -2486
rect 24448 -2558 24508 -2492
rect 24910 -2558 24970 -2492
rect 25364 -2558 25424 -2492
rect 25826 -2558 25886 -2492
rect 26280 -2558 26340 -2492
rect 26730 -2558 26790 -2492
rect 27196 -2558 27256 -2492
rect 27652 -2558 27712 -2492
rect 24448 -2618 27712 -2558
rect 24454 -2738 27718 -2678
rect 24454 -2804 24514 -2738
rect 24916 -2804 24976 -2738
rect 25370 -2804 25430 -2738
rect 25832 -2804 25892 -2738
rect 26286 -2804 26346 -2738
rect 26736 -2804 26796 -2738
rect 27202 -2804 27262 -2738
rect 27658 -2804 27718 -2738
rect 28114 -2804 28174 -2492
rect 24378 -2810 24586 -2804
rect 24378 -2844 24390 -2810
rect 24574 -2844 24586 -2810
rect 24378 -2850 24586 -2844
rect 24836 -2810 25044 -2804
rect 24836 -2844 24848 -2810
rect 25032 -2844 25044 -2810
rect 24836 -2850 25044 -2844
rect 25294 -2810 25502 -2804
rect 25294 -2844 25306 -2810
rect 25490 -2844 25502 -2810
rect 25294 -2850 25502 -2844
rect 25752 -2810 25960 -2804
rect 25752 -2844 25764 -2810
rect 25948 -2844 25960 -2810
rect 25752 -2850 25960 -2844
rect 26210 -2810 26418 -2804
rect 26210 -2844 26222 -2810
rect 26406 -2844 26418 -2810
rect 26210 -2850 26418 -2844
rect 26668 -2810 26876 -2804
rect 26668 -2844 26680 -2810
rect 26864 -2844 26876 -2810
rect 26668 -2850 26876 -2844
rect 27126 -2810 27334 -2804
rect 27126 -2844 27138 -2810
rect 27322 -2844 27334 -2810
rect 27126 -2850 27334 -2844
rect 27584 -2810 27792 -2804
rect 27584 -2844 27596 -2810
rect 27780 -2844 27792 -2810
rect 27584 -2850 27792 -2844
rect 28042 -2810 28250 -2804
rect 28042 -2844 28054 -2810
rect 28238 -2844 28250 -2810
rect 28042 -2850 28250 -2844
rect 23812 -3070 23818 -2914
rect 24222 -2922 24236 -2894
rect 23758 -3450 23818 -3070
rect 24230 -3070 24236 -2922
rect 24270 -2922 24282 -2894
rect 24688 -2894 24734 -2882
rect 24270 -3070 24276 -2922
rect 24230 -3082 24276 -3070
rect 24688 -3070 24694 -2894
rect 24728 -3070 24734 -2894
rect 24688 -3082 24734 -3070
rect 25146 -2894 25192 -2882
rect 25146 -3070 25152 -2894
rect 25186 -3070 25192 -2894
rect 25146 -3082 25192 -3070
rect 25604 -2894 25650 -2882
rect 25604 -3070 25610 -2894
rect 25644 -3070 25650 -2894
rect 25604 -3082 25650 -3070
rect 26062 -2894 26108 -2882
rect 26062 -3070 26068 -2894
rect 26102 -3070 26108 -2894
rect 26062 -3082 26108 -3070
rect 26520 -2894 26566 -2882
rect 26520 -3070 26526 -2894
rect 26560 -3070 26566 -2894
rect 26520 -3082 26566 -3070
rect 26978 -2894 27024 -2882
rect 26978 -3070 26984 -2894
rect 27018 -3070 27024 -2894
rect 26978 -3082 27024 -3070
rect 27436 -2894 27482 -2882
rect 27436 -3070 27442 -2894
rect 27476 -3070 27482 -2894
rect 27894 -2894 27940 -2882
rect 27894 -3042 27900 -2894
rect 27436 -3082 27482 -3070
rect 27886 -3070 27900 -3042
rect 27934 -3042 27940 -2894
rect 28346 -2894 28406 -2402
rect 27934 -3070 27946 -3042
rect 23920 -3120 24128 -3114
rect 23920 -3154 23932 -3120
rect 24116 -3154 24128 -3120
rect 23920 -3160 24128 -3154
rect 24378 -3120 24586 -3114
rect 24378 -3154 24390 -3120
rect 24574 -3154 24586 -3120
rect 24378 -3160 24586 -3154
rect 24836 -3120 25044 -3114
rect 24836 -3154 24848 -3120
rect 25032 -3154 25044 -3120
rect 24836 -3160 25044 -3154
rect 25294 -3120 25502 -3114
rect 25294 -3154 25306 -3120
rect 25490 -3154 25502 -3120
rect 25294 -3160 25502 -3154
rect 25752 -3120 25960 -3114
rect 25752 -3154 25764 -3120
rect 25948 -3154 25960 -3120
rect 25752 -3160 25960 -3154
rect 26210 -3120 26418 -3114
rect 26210 -3154 26222 -3120
rect 26406 -3154 26418 -3120
rect 26210 -3160 26418 -3154
rect 26668 -3120 26876 -3114
rect 26668 -3154 26680 -3120
rect 26864 -3154 26876 -3120
rect 26668 -3160 26876 -3154
rect 27126 -3120 27334 -3114
rect 27126 -3154 27138 -3120
rect 27322 -3154 27334 -3120
rect 27126 -3160 27334 -3154
rect 27584 -3120 27792 -3114
rect 27584 -3154 27596 -3120
rect 27780 -3154 27792 -3120
rect 27584 -3160 27792 -3154
rect 23998 -3450 24058 -3160
rect 24448 -3226 24508 -3160
rect 24910 -3226 24970 -3160
rect 25364 -3226 25424 -3160
rect 25826 -3226 25886 -3160
rect 26280 -3226 26340 -3160
rect 26730 -3226 26790 -3160
rect 27196 -3226 27256 -3160
rect 27652 -3226 27712 -3160
rect 24508 -3286 27712 -3226
rect 24448 -3292 24508 -3286
rect 27886 -3450 27946 -3070
rect 28346 -3070 28358 -2894
rect 28392 -3070 28406 -2894
rect 28042 -3120 28250 -3114
rect 28042 -3154 28054 -3120
rect 28238 -3154 28250 -3120
rect 28042 -3160 28250 -3154
rect 28112 -3450 28172 -3160
rect 28346 -3450 28406 -3070
rect 28762 -2402 28778 -2366
rect 28812 -2262 28826 -2226
rect 29222 -2226 29282 -1790
rect 32880 -1930 32886 -1870
rect 32946 -1930 32952 -1870
rect 31726 -2010 31732 -2006
rect 29444 -2070 29450 -2010
rect 29510 -2012 31732 -2010
rect 29510 -2070 29912 -2012
rect 29450 -2136 29514 -2070
rect 29906 -2072 29912 -2070
rect 29972 -2070 30366 -2012
rect 29972 -2072 29978 -2070
rect 30360 -2072 30366 -2070
rect 30426 -2070 30828 -2012
rect 30426 -2072 30432 -2070
rect 30822 -2072 30828 -2070
rect 30888 -2070 31282 -2012
rect 30888 -2072 30894 -2070
rect 31276 -2072 31282 -2070
rect 31342 -2066 31732 -2012
rect 31792 -2010 31798 -2006
rect 31792 -2066 32198 -2010
rect 31342 -2070 32198 -2066
rect 32258 -2070 32654 -2010
rect 32714 -2070 32720 -2010
rect 31342 -2072 31348 -2070
rect 29912 -2136 29976 -2072
rect 30366 -2136 30430 -2072
rect 30828 -2136 30892 -2072
rect 31282 -2136 31346 -2072
rect 31732 -2136 31796 -2070
rect 32198 -2136 32262 -2070
rect 32654 -2136 32718 -2070
rect 29378 -2142 29586 -2136
rect 29378 -2176 29390 -2142
rect 29574 -2176 29586 -2142
rect 29378 -2182 29586 -2176
rect 29836 -2142 30044 -2136
rect 29836 -2176 29848 -2142
rect 30032 -2176 30044 -2142
rect 29836 -2182 30044 -2176
rect 30294 -2142 30502 -2136
rect 30294 -2176 30306 -2142
rect 30490 -2176 30502 -2142
rect 30294 -2182 30502 -2176
rect 30752 -2142 30960 -2136
rect 30752 -2176 30764 -2142
rect 30948 -2176 30960 -2142
rect 30752 -2182 30960 -2176
rect 31210 -2142 31418 -2136
rect 31210 -2176 31222 -2142
rect 31406 -2176 31418 -2142
rect 31210 -2182 31418 -2176
rect 31668 -2142 31876 -2136
rect 31668 -2176 31680 -2142
rect 31864 -2176 31876 -2142
rect 31668 -2182 31876 -2176
rect 32126 -2142 32334 -2136
rect 32126 -2176 32138 -2142
rect 32322 -2176 32334 -2142
rect 32126 -2182 32334 -2176
rect 32584 -2142 32792 -2136
rect 32584 -2176 32596 -2142
rect 32780 -2176 32792 -2142
rect 32584 -2182 32792 -2176
rect 28812 -2366 28818 -2262
rect 29222 -2290 29236 -2226
rect 29230 -2358 29236 -2290
rect 28812 -2402 28822 -2366
rect 28762 -2556 28822 -2402
rect 29222 -2402 29236 -2358
rect 29270 -2290 29282 -2226
rect 29688 -2226 29734 -2214
rect 29270 -2358 29276 -2290
rect 29270 -2402 29282 -2358
rect 28920 -2452 29128 -2446
rect 28920 -2486 28932 -2452
rect 29116 -2486 29128 -2452
rect 28920 -2492 29128 -2486
rect 28990 -2556 29050 -2492
rect 29222 -2556 29282 -2402
rect 29688 -2402 29694 -2226
rect 29728 -2402 29734 -2226
rect 29688 -2414 29734 -2402
rect 30146 -2226 30192 -2214
rect 30146 -2402 30152 -2226
rect 30186 -2402 30192 -2226
rect 30146 -2414 30192 -2402
rect 30604 -2226 30650 -2214
rect 30604 -2402 30610 -2226
rect 30644 -2402 30650 -2226
rect 30604 -2414 30650 -2402
rect 31062 -2226 31108 -2214
rect 31062 -2402 31068 -2226
rect 31102 -2402 31108 -2226
rect 31062 -2414 31108 -2402
rect 31520 -2226 31566 -2214
rect 31520 -2402 31526 -2226
rect 31560 -2402 31566 -2226
rect 31520 -2414 31566 -2402
rect 31978 -2226 32024 -2214
rect 31978 -2402 31984 -2226
rect 32018 -2402 32024 -2226
rect 31978 -2414 32024 -2402
rect 32436 -2226 32482 -2214
rect 32436 -2402 32442 -2226
rect 32476 -2402 32482 -2226
rect 32886 -2226 32946 -1930
rect 33126 -2136 33186 -1790
rect 33042 -2142 33250 -2136
rect 33042 -2176 33054 -2142
rect 33238 -2176 33250 -2142
rect 33042 -2182 33250 -2176
rect 32886 -2268 32900 -2226
rect 32436 -2414 32482 -2402
rect 32894 -2402 32900 -2268
rect 32934 -2268 32946 -2226
rect 33344 -2226 33404 -1790
rect 33344 -2266 33358 -2226
rect 32934 -2402 32940 -2268
rect 33352 -2356 33358 -2266
rect 32894 -2414 32940 -2402
rect 33342 -2402 33358 -2356
rect 33392 -2266 33404 -2226
rect 33690 -1914 33802 -1790
rect 33392 -2356 33398 -2266
rect 33392 -2402 33402 -2356
rect 29378 -2452 29586 -2446
rect 29378 -2486 29390 -2452
rect 29574 -2486 29586 -2452
rect 29378 -2492 29586 -2486
rect 29836 -2452 30044 -2446
rect 29836 -2486 29848 -2452
rect 30032 -2486 30044 -2452
rect 29836 -2492 30044 -2486
rect 30294 -2452 30502 -2446
rect 30294 -2486 30306 -2452
rect 30490 -2486 30502 -2452
rect 30294 -2492 30502 -2486
rect 30752 -2452 30960 -2446
rect 30752 -2486 30764 -2452
rect 30948 -2486 30960 -2452
rect 30752 -2492 30960 -2486
rect 31210 -2452 31418 -2446
rect 31210 -2486 31222 -2452
rect 31406 -2486 31418 -2452
rect 31210 -2492 31418 -2486
rect 31668 -2452 31876 -2446
rect 31668 -2486 31680 -2452
rect 31864 -2486 31876 -2452
rect 31668 -2492 31876 -2486
rect 32126 -2452 32334 -2446
rect 32126 -2486 32138 -2452
rect 32322 -2486 32334 -2452
rect 32126 -2492 32334 -2486
rect 32584 -2452 32792 -2446
rect 32584 -2486 32596 -2452
rect 32780 -2486 32792 -2452
rect 32584 -2492 32792 -2486
rect 33042 -2452 33250 -2446
rect 33042 -2486 33054 -2452
rect 33238 -2486 33250 -2452
rect 33042 -2492 33250 -2486
rect 28762 -2616 29282 -2556
rect 28762 -3450 28822 -2616
rect 28990 -3450 29050 -2616
rect 29222 -3450 29282 -2616
rect 29448 -2558 29508 -2492
rect 29910 -2558 29970 -2492
rect 30364 -2558 30424 -2492
rect 30826 -2558 30886 -2492
rect 31280 -2558 31340 -2492
rect 31730 -2558 31790 -2492
rect 32196 -2558 32256 -2492
rect 32652 -2558 32712 -2492
rect 29448 -2618 32712 -2558
rect 33116 -3450 33176 -2492
rect 33342 -3450 33402 -2402
rect 23694 -3478 33464 -3450
rect 23694 -3564 23744 -3478
rect 23840 -3564 24324 -3478
rect 24420 -3564 24924 -3478
rect 25020 -3564 25524 -3478
rect 25620 -3564 26124 -3478
rect 26220 -3564 26724 -3478
rect 26820 -3564 27324 -3478
rect 27420 -3564 27924 -3478
rect 28020 -3564 28524 -3478
rect 28620 -3564 29124 -3478
rect 29220 -3564 29724 -3478
rect 29820 -3564 30324 -3478
rect 30420 -3564 30924 -3478
rect 31020 -3564 31524 -3478
rect 31620 -3564 32124 -3478
rect 32220 -3564 32724 -3478
rect 32820 -3564 33324 -3478
rect 33420 -3564 33464 -3478
rect 23694 -3594 33464 -3564
rect 23346 -4042 23458 -3918
rect 24058 -4042 24068 -3742
rect 33080 -4042 33090 -3742
rect 33690 -3918 33696 -1914
rect 33796 -3918 33802 -1914
rect 33690 -4042 33802 -3918
rect 23346 -4048 33802 -4042
rect 23346 -4148 23452 -4048
rect 33696 -4148 33802 -4048
rect 23346 -4154 33802 -4148
rect 22934 -16876 22940 -16816
rect 23000 -16876 23006 -16816
rect 18690 -19342 18802 -19166
rect 8346 -19348 18802 -19342
rect 8346 -19448 8452 -19348
rect 18696 -19448 18802 -19348
rect 8346 -19454 18802 -19448
rect 8346 -19684 18802 -19678
rect 8346 -19784 8452 -19684
rect 18696 -19784 18802 -19684
rect 8346 -19790 18802 -19784
rect 8346 -19914 8458 -19790
rect 8346 -21918 8352 -19914
rect 8452 -21918 8458 -19914
rect 8766 -20226 8826 -19790
rect 8996 -20136 9056 -19790
rect 12886 -19882 12946 -19876
rect 9454 -20016 9910 -20010
rect 9442 -20076 9448 -20016
rect 9508 -20070 9910 -20016
rect 9970 -20016 10826 -20010
rect 9970 -20070 10364 -20016
rect 9508 -20076 9514 -20070
rect 9448 -20136 9514 -20076
rect 9910 -20136 9976 -20070
rect 10358 -20076 10364 -20070
rect 10424 -20070 10826 -20016
rect 10886 -20070 11280 -20010
rect 11340 -20070 11730 -20010
rect 11790 -20016 12652 -20010
rect 11790 -20070 12196 -20016
rect 10424 -20076 10430 -20070
rect 10364 -20136 10430 -20076
rect 10826 -20136 10892 -20070
rect 11280 -20136 11346 -20070
rect 11730 -20136 11796 -20070
rect 12190 -20076 12196 -20070
rect 12256 -20070 12652 -20016
rect 12712 -20070 12718 -20010
rect 12256 -20076 12262 -20070
rect 12196 -20136 12262 -20076
rect 12652 -20136 12718 -20070
rect 8920 -20142 9128 -20136
rect 8920 -20176 8932 -20142
rect 9116 -20176 9128 -20142
rect 8920 -20182 9128 -20176
rect 9378 -20142 9586 -20136
rect 9378 -20176 9390 -20142
rect 9574 -20176 9586 -20142
rect 9378 -20182 9586 -20176
rect 9836 -20142 10044 -20136
rect 9836 -20176 9848 -20142
rect 10032 -20176 10044 -20142
rect 9836 -20182 10044 -20176
rect 10294 -20142 10502 -20136
rect 10294 -20176 10306 -20142
rect 10490 -20176 10502 -20142
rect 10294 -20182 10502 -20176
rect 10752 -20142 10960 -20136
rect 10752 -20176 10764 -20142
rect 10948 -20176 10960 -20142
rect 10752 -20182 10960 -20176
rect 11210 -20142 11418 -20136
rect 11210 -20176 11222 -20142
rect 11406 -20176 11418 -20142
rect 11210 -20182 11418 -20176
rect 11668 -20142 11876 -20136
rect 11668 -20176 11680 -20142
rect 11864 -20176 11876 -20142
rect 11668 -20182 11876 -20176
rect 12126 -20142 12334 -20136
rect 12126 -20176 12138 -20142
rect 12322 -20176 12334 -20142
rect 12126 -20182 12334 -20176
rect 12584 -20142 12792 -20136
rect 12584 -20176 12596 -20142
rect 12780 -20176 12792 -20142
rect 12584 -20182 12792 -20176
rect 8766 -20266 8778 -20226
rect 8772 -20362 8778 -20266
rect 8766 -20402 8778 -20362
rect 8812 -20266 8826 -20226
rect 9230 -20226 9276 -20214
rect 8812 -20362 8818 -20266
rect 9230 -20360 9236 -20226
rect 8812 -20402 8826 -20362
rect 8766 -20618 8826 -20402
rect 9222 -20402 9236 -20360
rect 9270 -20360 9276 -20226
rect 9688 -20226 9734 -20214
rect 9270 -20402 9282 -20360
rect 8920 -20452 9128 -20446
rect 8920 -20486 8932 -20452
rect 9116 -20486 9128 -20452
rect 8920 -20492 9128 -20486
rect 8994 -20618 9054 -20492
rect 8766 -20678 9054 -20618
rect 8766 -20894 8826 -20678
rect 8994 -20804 9054 -20678
rect 8920 -20810 9128 -20804
rect 8920 -20844 8932 -20810
rect 9116 -20844 9128 -20810
rect 8920 -20850 9128 -20844
rect 8766 -20914 8778 -20894
rect 8772 -21040 8778 -20914
rect 8758 -21070 8778 -21040
rect 8812 -20914 8826 -20894
rect 9222 -20894 9282 -20402
rect 9688 -20402 9694 -20226
rect 9728 -20402 9734 -20226
rect 9688 -20414 9734 -20402
rect 10146 -20226 10192 -20214
rect 10146 -20402 10152 -20226
rect 10186 -20402 10192 -20226
rect 10146 -20414 10192 -20402
rect 10604 -20226 10650 -20214
rect 10604 -20402 10610 -20226
rect 10644 -20402 10650 -20226
rect 10604 -20414 10650 -20402
rect 11062 -20226 11108 -20214
rect 11062 -20402 11068 -20226
rect 11102 -20402 11108 -20226
rect 11062 -20414 11108 -20402
rect 11520 -20226 11566 -20214
rect 11520 -20402 11526 -20226
rect 11560 -20402 11566 -20226
rect 11520 -20414 11566 -20402
rect 11978 -20226 12024 -20214
rect 11978 -20402 11984 -20226
rect 12018 -20402 12024 -20226
rect 11978 -20414 12024 -20402
rect 12436 -20226 12482 -20214
rect 12436 -20402 12442 -20226
rect 12476 -20402 12482 -20226
rect 12886 -20226 12946 -19942
rect 13114 -20136 13174 -19790
rect 13042 -20142 13250 -20136
rect 13042 -20176 13054 -20142
rect 13238 -20176 13250 -20142
rect 13042 -20182 13250 -20176
rect 12886 -20256 12900 -20226
rect 12436 -20414 12482 -20402
rect 12894 -20402 12900 -20256
rect 12934 -20256 12946 -20226
rect 13346 -20226 13406 -19790
rect 13346 -20254 13358 -20226
rect 12934 -20402 12940 -20256
rect 13352 -20346 13358 -20254
rect 12894 -20414 12940 -20402
rect 13346 -20402 13358 -20346
rect 13392 -20254 13406 -20226
rect 13766 -20226 13826 -19790
rect 14000 -20136 14060 -19790
rect 13920 -20142 14128 -20136
rect 13920 -20176 13932 -20142
rect 14116 -20176 14128 -20142
rect 13920 -20182 14128 -20176
rect 13392 -20346 13398 -20254
rect 13766 -20262 13778 -20226
rect 13392 -20402 13406 -20346
rect 13772 -20366 13778 -20262
rect 9378 -20452 9586 -20446
rect 9378 -20486 9390 -20452
rect 9574 -20486 9586 -20452
rect 9378 -20492 9586 -20486
rect 9836 -20452 10044 -20446
rect 9836 -20486 9848 -20452
rect 10032 -20486 10044 -20452
rect 9836 -20492 10044 -20486
rect 10294 -20452 10502 -20446
rect 10294 -20486 10306 -20452
rect 10490 -20486 10502 -20452
rect 10294 -20492 10502 -20486
rect 10752 -20452 10960 -20446
rect 10752 -20486 10764 -20452
rect 10948 -20486 10960 -20452
rect 10752 -20492 10960 -20486
rect 11210 -20452 11418 -20446
rect 11210 -20486 11222 -20452
rect 11406 -20486 11418 -20452
rect 11210 -20492 11418 -20486
rect 11668 -20452 11876 -20446
rect 11668 -20486 11680 -20452
rect 11864 -20486 11876 -20452
rect 11668 -20492 11876 -20486
rect 12126 -20452 12334 -20446
rect 12126 -20486 12138 -20452
rect 12322 -20486 12334 -20452
rect 12126 -20492 12334 -20486
rect 12584 -20452 12792 -20446
rect 12584 -20486 12596 -20452
rect 12780 -20486 12792 -20452
rect 12584 -20492 12792 -20486
rect 13042 -20452 13250 -20446
rect 13042 -20486 13054 -20452
rect 13238 -20486 13250 -20452
rect 13042 -20492 13250 -20486
rect 9448 -20558 9508 -20492
rect 9910 -20558 9970 -20492
rect 10364 -20558 10424 -20492
rect 10826 -20558 10886 -20492
rect 11280 -20558 11340 -20492
rect 11730 -20558 11790 -20492
rect 12196 -20558 12256 -20492
rect 12652 -20558 12712 -20492
rect 9448 -20618 12712 -20558
rect 9454 -20738 12718 -20678
rect 9454 -20804 9514 -20738
rect 9916 -20804 9976 -20738
rect 10370 -20804 10430 -20738
rect 10832 -20804 10892 -20738
rect 11286 -20804 11346 -20738
rect 11736 -20804 11796 -20738
rect 12202 -20804 12262 -20738
rect 12658 -20804 12718 -20738
rect 13114 -20804 13174 -20492
rect 9378 -20810 9586 -20804
rect 9378 -20844 9390 -20810
rect 9574 -20844 9586 -20810
rect 9378 -20850 9586 -20844
rect 9836 -20810 10044 -20804
rect 9836 -20844 9848 -20810
rect 10032 -20844 10044 -20810
rect 9836 -20850 10044 -20844
rect 10294 -20810 10502 -20804
rect 10294 -20844 10306 -20810
rect 10490 -20844 10502 -20810
rect 10294 -20850 10502 -20844
rect 10752 -20810 10960 -20804
rect 10752 -20844 10764 -20810
rect 10948 -20844 10960 -20810
rect 10752 -20850 10960 -20844
rect 11210 -20810 11418 -20804
rect 11210 -20844 11222 -20810
rect 11406 -20844 11418 -20810
rect 11210 -20850 11418 -20844
rect 11668 -20810 11876 -20804
rect 11668 -20844 11680 -20810
rect 11864 -20844 11876 -20810
rect 11668 -20850 11876 -20844
rect 12126 -20810 12334 -20804
rect 12126 -20844 12138 -20810
rect 12322 -20844 12334 -20810
rect 12126 -20850 12334 -20844
rect 12584 -20810 12792 -20804
rect 12584 -20844 12596 -20810
rect 12780 -20844 12792 -20810
rect 12584 -20850 12792 -20844
rect 13042 -20810 13250 -20804
rect 13042 -20844 13054 -20810
rect 13238 -20844 13250 -20810
rect 13042 -20850 13250 -20844
rect 8812 -21070 8818 -20914
rect 9222 -20922 9236 -20894
rect 8758 -21450 8818 -21070
rect 9230 -21070 9236 -20922
rect 9270 -20922 9282 -20894
rect 9688 -20894 9734 -20882
rect 9270 -21070 9276 -20922
rect 9230 -21082 9276 -21070
rect 9688 -21070 9694 -20894
rect 9728 -21070 9734 -20894
rect 9688 -21082 9734 -21070
rect 10146 -20894 10192 -20882
rect 10146 -21070 10152 -20894
rect 10186 -21070 10192 -20894
rect 10146 -21082 10192 -21070
rect 10604 -20894 10650 -20882
rect 10604 -21070 10610 -20894
rect 10644 -21070 10650 -20894
rect 10604 -21082 10650 -21070
rect 11062 -20894 11108 -20882
rect 11062 -21070 11068 -20894
rect 11102 -21070 11108 -20894
rect 11062 -21082 11108 -21070
rect 11520 -20894 11566 -20882
rect 11520 -21070 11526 -20894
rect 11560 -21070 11566 -20894
rect 11520 -21082 11566 -21070
rect 11978 -20894 12024 -20882
rect 11978 -21070 11984 -20894
rect 12018 -21070 12024 -20894
rect 11978 -21082 12024 -21070
rect 12436 -20894 12482 -20882
rect 12436 -21070 12442 -20894
rect 12476 -21070 12482 -20894
rect 12894 -20894 12940 -20882
rect 12894 -21042 12900 -20894
rect 12436 -21082 12482 -21070
rect 12886 -21070 12900 -21042
rect 12934 -21042 12940 -20894
rect 13346 -20894 13406 -20402
rect 12934 -21070 12946 -21042
rect 8920 -21120 9128 -21114
rect 8920 -21154 8932 -21120
rect 9116 -21154 9128 -21120
rect 8920 -21160 9128 -21154
rect 9378 -21120 9586 -21114
rect 9378 -21154 9390 -21120
rect 9574 -21154 9586 -21120
rect 9378 -21160 9586 -21154
rect 9836 -21120 10044 -21114
rect 9836 -21154 9848 -21120
rect 10032 -21154 10044 -21120
rect 9836 -21160 10044 -21154
rect 10294 -21120 10502 -21114
rect 10294 -21154 10306 -21120
rect 10490 -21154 10502 -21120
rect 10294 -21160 10502 -21154
rect 10752 -21120 10960 -21114
rect 10752 -21154 10764 -21120
rect 10948 -21154 10960 -21120
rect 10752 -21160 10960 -21154
rect 11210 -21120 11418 -21114
rect 11210 -21154 11222 -21120
rect 11406 -21154 11418 -21120
rect 11210 -21160 11418 -21154
rect 11668 -21120 11876 -21114
rect 11668 -21154 11680 -21120
rect 11864 -21154 11876 -21120
rect 11668 -21160 11876 -21154
rect 12126 -21120 12334 -21114
rect 12126 -21154 12138 -21120
rect 12322 -21154 12334 -21120
rect 12126 -21160 12334 -21154
rect 12584 -21120 12792 -21114
rect 12584 -21154 12596 -21120
rect 12780 -21154 12792 -21120
rect 12584 -21160 12792 -21154
rect 8998 -21450 9058 -21160
rect 9448 -21226 9508 -21160
rect 9910 -21226 9970 -21160
rect 10364 -21226 10424 -21160
rect 10826 -21226 10886 -21160
rect 11280 -21226 11340 -21160
rect 11730 -21226 11790 -21160
rect 12196 -21226 12256 -21160
rect 12652 -21226 12712 -21160
rect 9448 -21286 12652 -21226
rect 12652 -21292 12712 -21286
rect 12886 -21450 12946 -21070
rect 13346 -21070 13358 -20894
rect 13392 -21070 13406 -20894
rect 13042 -21120 13250 -21114
rect 13042 -21154 13054 -21120
rect 13238 -21154 13250 -21120
rect 13042 -21160 13250 -21154
rect 13112 -21450 13172 -21160
rect 13346 -21450 13406 -21070
rect 13762 -20402 13778 -20366
rect 13812 -20262 13826 -20226
rect 14222 -20226 14282 -19790
rect 17880 -19930 17886 -19870
rect 17946 -19930 17952 -19870
rect 16726 -20010 16732 -20006
rect 14444 -20070 14450 -20010
rect 14510 -20012 16732 -20010
rect 14510 -20070 14912 -20012
rect 14450 -20136 14514 -20070
rect 14906 -20072 14912 -20070
rect 14972 -20070 15366 -20012
rect 14972 -20072 14978 -20070
rect 15360 -20072 15366 -20070
rect 15426 -20070 15828 -20012
rect 15426 -20072 15432 -20070
rect 15822 -20072 15828 -20070
rect 15888 -20070 16282 -20012
rect 15888 -20072 15894 -20070
rect 16276 -20072 16282 -20070
rect 16342 -20066 16732 -20012
rect 16792 -20010 16798 -20006
rect 16792 -20066 17198 -20010
rect 16342 -20070 17198 -20066
rect 17258 -20070 17654 -20010
rect 17714 -20070 17720 -20010
rect 16342 -20072 16348 -20070
rect 14912 -20136 14976 -20072
rect 15366 -20136 15430 -20072
rect 15828 -20136 15892 -20072
rect 16282 -20136 16346 -20072
rect 16732 -20136 16796 -20070
rect 17198 -20136 17262 -20070
rect 17654 -20136 17718 -20070
rect 14378 -20142 14586 -20136
rect 14378 -20176 14390 -20142
rect 14574 -20176 14586 -20142
rect 14378 -20182 14586 -20176
rect 14836 -20142 15044 -20136
rect 14836 -20176 14848 -20142
rect 15032 -20176 15044 -20142
rect 14836 -20182 15044 -20176
rect 15294 -20142 15502 -20136
rect 15294 -20176 15306 -20142
rect 15490 -20176 15502 -20142
rect 15294 -20182 15502 -20176
rect 15752 -20142 15960 -20136
rect 15752 -20176 15764 -20142
rect 15948 -20176 15960 -20142
rect 15752 -20182 15960 -20176
rect 16210 -20142 16418 -20136
rect 16210 -20176 16222 -20142
rect 16406 -20176 16418 -20142
rect 16210 -20182 16418 -20176
rect 16668 -20142 16876 -20136
rect 16668 -20176 16680 -20142
rect 16864 -20176 16876 -20142
rect 16668 -20182 16876 -20176
rect 17126 -20142 17334 -20136
rect 17126 -20176 17138 -20142
rect 17322 -20176 17334 -20142
rect 17126 -20182 17334 -20176
rect 17584 -20142 17792 -20136
rect 17584 -20176 17596 -20142
rect 17780 -20176 17792 -20142
rect 17584 -20182 17792 -20176
rect 13812 -20366 13818 -20262
rect 14222 -20290 14236 -20226
rect 14230 -20358 14236 -20290
rect 13812 -20402 13822 -20366
rect 13762 -20556 13822 -20402
rect 14222 -20402 14236 -20358
rect 14270 -20290 14282 -20226
rect 14688 -20226 14734 -20214
rect 14270 -20358 14276 -20290
rect 14270 -20402 14282 -20358
rect 13920 -20452 14128 -20446
rect 13920 -20486 13932 -20452
rect 14116 -20486 14128 -20452
rect 13920 -20492 14128 -20486
rect 13990 -20556 14050 -20492
rect 14222 -20556 14282 -20402
rect 14688 -20402 14694 -20226
rect 14728 -20402 14734 -20226
rect 14688 -20414 14734 -20402
rect 15146 -20226 15192 -20214
rect 15146 -20402 15152 -20226
rect 15186 -20402 15192 -20226
rect 15146 -20414 15192 -20402
rect 15604 -20226 15650 -20214
rect 15604 -20402 15610 -20226
rect 15644 -20402 15650 -20226
rect 15604 -20414 15650 -20402
rect 16062 -20226 16108 -20214
rect 16062 -20402 16068 -20226
rect 16102 -20402 16108 -20226
rect 16062 -20414 16108 -20402
rect 16520 -20226 16566 -20214
rect 16520 -20402 16526 -20226
rect 16560 -20402 16566 -20226
rect 16520 -20414 16566 -20402
rect 16978 -20226 17024 -20214
rect 16978 -20402 16984 -20226
rect 17018 -20402 17024 -20226
rect 16978 -20414 17024 -20402
rect 17436 -20226 17482 -20214
rect 17436 -20402 17442 -20226
rect 17476 -20402 17482 -20226
rect 17886 -20226 17946 -19930
rect 18126 -20136 18186 -19790
rect 18042 -20142 18250 -20136
rect 18042 -20176 18054 -20142
rect 18238 -20176 18250 -20142
rect 18042 -20182 18250 -20176
rect 17886 -20268 17900 -20226
rect 17436 -20414 17482 -20402
rect 17894 -20402 17900 -20268
rect 17934 -20268 17946 -20226
rect 18344 -20226 18404 -19790
rect 18344 -20266 18358 -20226
rect 17934 -20402 17940 -20268
rect 18352 -20356 18358 -20266
rect 17894 -20414 17940 -20402
rect 18342 -20402 18358 -20356
rect 18392 -20266 18404 -20226
rect 18690 -19914 18802 -19790
rect 18392 -20356 18398 -20266
rect 18392 -20402 18402 -20356
rect 14378 -20452 14586 -20446
rect 14378 -20486 14390 -20452
rect 14574 -20486 14586 -20452
rect 14378 -20492 14586 -20486
rect 14836 -20452 15044 -20446
rect 14836 -20486 14848 -20452
rect 15032 -20486 15044 -20452
rect 14836 -20492 15044 -20486
rect 15294 -20452 15502 -20446
rect 15294 -20486 15306 -20452
rect 15490 -20486 15502 -20452
rect 15294 -20492 15502 -20486
rect 15752 -20452 15960 -20446
rect 15752 -20486 15764 -20452
rect 15948 -20486 15960 -20452
rect 15752 -20492 15960 -20486
rect 16210 -20452 16418 -20446
rect 16210 -20486 16222 -20452
rect 16406 -20486 16418 -20452
rect 16210 -20492 16418 -20486
rect 16668 -20452 16876 -20446
rect 16668 -20486 16680 -20452
rect 16864 -20486 16876 -20452
rect 16668 -20492 16876 -20486
rect 17126 -20452 17334 -20446
rect 17126 -20486 17138 -20452
rect 17322 -20486 17334 -20452
rect 17126 -20492 17334 -20486
rect 17584 -20452 17792 -20446
rect 17584 -20486 17596 -20452
rect 17780 -20486 17792 -20452
rect 17584 -20492 17792 -20486
rect 18042 -20452 18250 -20446
rect 18042 -20486 18054 -20452
rect 18238 -20486 18250 -20452
rect 18042 -20492 18250 -20486
rect 13762 -20616 14282 -20556
rect 13762 -21450 13822 -20616
rect 13990 -21450 14050 -20616
rect 14222 -21450 14282 -20616
rect 14448 -20558 14508 -20492
rect 14910 -20558 14970 -20492
rect 15364 -20558 15424 -20492
rect 15826 -20558 15886 -20492
rect 16280 -20558 16340 -20492
rect 16730 -20558 16790 -20492
rect 17196 -20558 17256 -20492
rect 17652 -20558 17712 -20492
rect 14448 -20618 17712 -20558
rect 18116 -21450 18176 -20492
rect 18342 -21450 18402 -20402
rect 8694 -21478 18464 -21450
rect 8694 -21564 8744 -21478
rect 8840 -21564 9324 -21478
rect 9420 -21564 9924 -21478
rect 10020 -21564 10524 -21478
rect 10620 -21564 11124 -21478
rect 11220 -21564 11724 -21478
rect 11820 -21564 12324 -21478
rect 12420 -21564 12924 -21478
rect 13020 -21564 13524 -21478
rect 13620 -21564 14124 -21478
rect 14220 -21564 14724 -21478
rect 14820 -21564 15324 -21478
rect 15420 -21564 15924 -21478
rect 16020 -21564 16524 -21478
rect 16620 -21564 17124 -21478
rect 17220 -21564 17724 -21478
rect 17820 -21564 18324 -21478
rect 18420 -21564 18464 -21478
rect 8694 -21594 18464 -21564
rect 8346 -22042 8458 -21918
rect 9058 -22042 9068 -21742
rect 18080 -22042 18090 -21742
rect 18690 -21918 18696 -19914
rect 18796 -21918 18802 -19914
rect 23080 -21226 23140 -5530
rect 27300 -4608 37756 -4602
rect 27300 -4708 27406 -4608
rect 37650 -4708 37756 -4608
rect 27300 -4714 37756 -4708
rect 27300 -4838 27412 -4714
rect 27300 -6842 27306 -4838
rect 27406 -6842 27412 -4838
rect 28012 -5014 28022 -4714
rect 37034 -5014 37044 -4714
rect 37644 -4838 37756 -4714
rect 27638 -5192 37408 -5162
rect 27638 -5278 27682 -5192
rect 27778 -5278 28282 -5192
rect 28378 -5278 28882 -5192
rect 28978 -5278 29482 -5192
rect 29578 -5278 30082 -5192
rect 30178 -5278 30682 -5192
rect 30778 -5278 31282 -5192
rect 31378 -5278 31882 -5192
rect 31978 -5278 32482 -5192
rect 32578 -5278 33082 -5192
rect 33178 -5278 33682 -5192
rect 33778 -5278 34282 -5192
rect 34378 -5278 34882 -5192
rect 34978 -5278 35482 -5192
rect 35578 -5278 36082 -5192
rect 36178 -5278 36682 -5192
rect 36778 -5278 37262 -5192
rect 37358 -5278 37408 -5192
rect 27638 -5306 37408 -5278
rect 27700 -6354 27760 -5306
rect 27926 -6264 27986 -5306
rect 28390 -6198 31654 -6138
rect 28390 -6264 28450 -6198
rect 28846 -6264 28906 -6198
rect 29312 -6264 29372 -6198
rect 29762 -6264 29822 -6198
rect 30216 -6264 30276 -6198
rect 30678 -6264 30738 -6198
rect 31132 -6264 31192 -6198
rect 31594 -6264 31654 -6198
rect 31820 -6140 31880 -5306
rect 32052 -6140 32112 -5306
rect 32280 -6140 32340 -5306
rect 31820 -6200 32340 -6140
rect 27852 -6270 28060 -6264
rect 27852 -6304 27864 -6270
rect 28048 -6304 28060 -6270
rect 27852 -6310 28060 -6304
rect 28310 -6270 28518 -6264
rect 28310 -6304 28322 -6270
rect 28506 -6304 28518 -6270
rect 28310 -6310 28518 -6304
rect 28768 -6270 28976 -6264
rect 28768 -6304 28780 -6270
rect 28964 -6304 28976 -6270
rect 28768 -6310 28976 -6304
rect 29226 -6270 29434 -6264
rect 29226 -6304 29238 -6270
rect 29422 -6304 29434 -6270
rect 29226 -6310 29434 -6304
rect 29684 -6270 29892 -6264
rect 29684 -6304 29696 -6270
rect 29880 -6304 29892 -6270
rect 29684 -6310 29892 -6304
rect 30142 -6270 30350 -6264
rect 30142 -6304 30154 -6270
rect 30338 -6304 30350 -6270
rect 30142 -6310 30350 -6304
rect 30600 -6270 30808 -6264
rect 30600 -6304 30612 -6270
rect 30796 -6304 30808 -6270
rect 30600 -6310 30808 -6304
rect 31058 -6270 31266 -6264
rect 31058 -6304 31070 -6270
rect 31254 -6304 31266 -6270
rect 31058 -6310 31266 -6304
rect 31516 -6270 31724 -6264
rect 31516 -6304 31528 -6270
rect 31712 -6304 31724 -6270
rect 31516 -6310 31724 -6304
rect 27700 -6400 27710 -6354
rect 27704 -6490 27710 -6400
rect 27300 -6966 27412 -6842
rect 27698 -6530 27710 -6490
rect 27744 -6400 27760 -6354
rect 28162 -6354 28208 -6342
rect 27744 -6490 27750 -6400
rect 28162 -6488 28168 -6354
rect 27744 -6530 27758 -6490
rect 27698 -6966 27758 -6530
rect 28156 -6530 28168 -6488
rect 28202 -6488 28208 -6354
rect 28620 -6354 28666 -6342
rect 28202 -6530 28216 -6488
rect 27852 -6580 28060 -6574
rect 27852 -6614 27864 -6580
rect 28048 -6614 28060 -6580
rect 27852 -6620 28060 -6614
rect 27916 -6966 27976 -6620
rect 28156 -6826 28216 -6530
rect 28620 -6530 28626 -6354
rect 28660 -6530 28666 -6354
rect 28620 -6542 28666 -6530
rect 29078 -6354 29124 -6342
rect 29078 -6530 29084 -6354
rect 29118 -6530 29124 -6354
rect 29078 -6542 29124 -6530
rect 29536 -6354 29582 -6342
rect 29536 -6530 29542 -6354
rect 29576 -6530 29582 -6354
rect 29536 -6542 29582 -6530
rect 29994 -6354 30040 -6342
rect 29994 -6530 30000 -6354
rect 30034 -6530 30040 -6354
rect 29994 -6542 30040 -6530
rect 30452 -6354 30498 -6342
rect 30452 -6530 30458 -6354
rect 30492 -6530 30498 -6354
rect 30452 -6542 30498 -6530
rect 30910 -6354 30956 -6342
rect 30910 -6530 30916 -6354
rect 30950 -6530 30956 -6354
rect 30910 -6542 30956 -6530
rect 31368 -6354 31414 -6342
rect 31368 -6530 31374 -6354
rect 31408 -6530 31414 -6354
rect 31820 -6354 31880 -6200
rect 32052 -6264 32112 -6200
rect 31974 -6270 32182 -6264
rect 31974 -6304 31986 -6270
rect 32170 -6304 32182 -6270
rect 31974 -6310 32182 -6304
rect 31820 -6398 31832 -6354
rect 31826 -6466 31832 -6398
rect 31368 -6542 31414 -6530
rect 31820 -6530 31832 -6466
rect 31866 -6398 31880 -6354
rect 32280 -6354 32340 -6200
rect 32280 -6390 32290 -6354
rect 31866 -6466 31872 -6398
rect 31866 -6530 31880 -6466
rect 32284 -6494 32290 -6390
rect 28310 -6580 28518 -6574
rect 28310 -6614 28322 -6580
rect 28506 -6614 28518 -6580
rect 28310 -6620 28518 -6614
rect 28768 -6580 28976 -6574
rect 28768 -6614 28780 -6580
rect 28964 -6614 28976 -6580
rect 28768 -6620 28976 -6614
rect 29226 -6580 29434 -6574
rect 29226 -6614 29238 -6580
rect 29422 -6614 29434 -6580
rect 29226 -6620 29434 -6614
rect 29684 -6580 29892 -6574
rect 29684 -6614 29696 -6580
rect 29880 -6614 29892 -6580
rect 29684 -6620 29892 -6614
rect 30142 -6580 30350 -6574
rect 30142 -6614 30154 -6580
rect 30338 -6614 30350 -6580
rect 30142 -6620 30350 -6614
rect 30600 -6580 30808 -6574
rect 30600 -6614 30612 -6580
rect 30796 -6614 30808 -6580
rect 30600 -6620 30808 -6614
rect 31058 -6580 31266 -6574
rect 31058 -6614 31070 -6580
rect 31254 -6614 31266 -6580
rect 31058 -6620 31266 -6614
rect 31516 -6580 31724 -6574
rect 31516 -6614 31528 -6580
rect 31712 -6614 31724 -6580
rect 31516 -6620 31724 -6614
rect 28384 -6686 28448 -6620
rect 28840 -6686 28904 -6620
rect 29306 -6686 29370 -6620
rect 29756 -6684 29820 -6620
rect 30210 -6684 30274 -6620
rect 30672 -6684 30736 -6620
rect 31126 -6684 31190 -6620
rect 29754 -6686 29760 -6684
rect 28382 -6746 28388 -6686
rect 28448 -6746 28844 -6686
rect 28904 -6690 29760 -6686
rect 28904 -6746 29310 -6690
rect 29304 -6750 29310 -6746
rect 29370 -6744 29760 -6690
rect 29820 -6686 29826 -6684
rect 30208 -6686 30214 -6684
rect 29820 -6744 30214 -6686
rect 30274 -6686 30280 -6684
rect 30670 -6686 30676 -6684
rect 30274 -6744 30676 -6686
rect 30736 -6686 30742 -6684
rect 31124 -6686 31130 -6684
rect 30736 -6744 31130 -6686
rect 31190 -6686 31196 -6684
rect 31588 -6686 31652 -6620
rect 31190 -6744 31592 -6686
rect 29370 -6746 31592 -6744
rect 31652 -6746 31658 -6686
rect 29370 -6750 29376 -6746
rect 28150 -6886 28156 -6826
rect 28216 -6886 28222 -6826
rect 31820 -6966 31880 -6530
rect 32276 -6530 32290 -6494
rect 32324 -6390 32340 -6354
rect 32696 -5686 32756 -5306
rect 32930 -5596 32990 -5306
rect 32852 -5602 33060 -5596
rect 32852 -5636 32864 -5602
rect 33048 -5636 33060 -5602
rect 32852 -5642 33060 -5636
rect 32696 -5862 32710 -5686
rect 32744 -5862 32756 -5686
rect 33156 -5686 33216 -5306
rect 33390 -5470 33450 -5464
rect 33450 -5530 36654 -5470
rect 33390 -5596 33450 -5530
rect 33846 -5596 33906 -5530
rect 34312 -5596 34372 -5530
rect 34762 -5596 34822 -5530
rect 35216 -5596 35276 -5530
rect 35678 -5596 35738 -5530
rect 36132 -5596 36192 -5530
rect 36594 -5596 36654 -5530
rect 37044 -5596 37104 -5306
rect 33310 -5602 33518 -5596
rect 33310 -5636 33322 -5602
rect 33506 -5636 33518 -5602
rect 33310 -5642 33518 -5636
rect 33768 -5602 33976 -5596
rect 33768 -5636 33780 -5602
rect 33964 -5636 33976 -5602
rect 33768 -5642 33976 -5636
rect 34226 -5602 34434 -5596
rect 34226 -5636 34238 -5602
rect 34422 -5636 34434 -5602
rect 34226 -5642 34434 -5636
rect 34684 -5602 34892 -5596
rect 34684 -5636 34696 -5602
rect 34880 -5636 34892 -5602
rect 34684 -5642 34892 -5636
rect 35142 -5602 35350 -5596
rect 35142 -5636 35154 -5602
rect 35338 -5636 35350 -5602
rect 35142 -5642 35350 -5636
rect 35600 -5602 35808 -5596
rect 35600 -5636 35612 -5602
rect 35796 -5636 35808 -5602
rect 35600 -5642 35808 -5636
rect 36058 -5602 36266 -5596
rect 36058 -5636 36070 -5602
rect 36254 -5636 36266 -5602
rect 36058 -5642 36266 -5636
rect 36516 -5602 36724 -5596
rect 36516 -5636 36528 -5602
rect 36712 -5636 36724 -5602
rect 36516 -5642 36724 -5636
rect 36974 -5602 37182 -5596
rect 36974 -5636 36986 -5602
rect 37170 -5636 37182 -5602
rect 36974 -5642 37182 -5636
rect 33156 -5714 33168 -5686
rect 32696 -6354 32756 -5862
rect 33162 -5862 33168 -5714
rect 33202 -5714 33216 -5686
rect 33620 -5686 33666 -5674
rect 33202 -5862 33208 -5714
rect 33162 -5874 33208 -5862
rect 33620 -5862 33626 -5686
rect 33660 -5862 33666 -5686
rect 33620 -5874 33666 -5862
rect 34078 -5686 34124 -5674
rect 34078 -5862 34084 -5686
rect 34118 -5862 34124 -5686
rect 34078 -5874 34124 -5862
rect 34536 -5686 34582 -5674
rect 34536 -5862 34542 -5686
rect 34576 -5862 34582 -5686
rect 34536 -5874 34582 -5862
rect 34994 -5686 35040 -5674
rect 34994 -5862 35000 -5686
rect 35034 -5862 35040 -5686
rect 34994 -5874 35040 -5862
rect 35452 -5686 35498 -5674
rect 35452 -5862 35458 -5686
rect 35492 -5862 35498 -5686
rect 35452 -5874 35498 -5862
rect 35910 -5686 35956 -5674
rect 35910 -5862 35916 -5686
rect 35950 -5862 35956 -5686
rect 35910 -5874 35956 -5862
rect 36368 -5686 36414 -5674
rect 36368 -5862 36374 -5686
rect 36408 -5862 36414 -5686
rect 36826 -5686 36872 -5674
rect 36826 -5834 36832 -5686
rect 36368 -5874 36414 -5862
rect 36820 -5862 36832 -5834
rect 36866 -5834 36872 -5686
rect 37284 -5686 37344 -5306
rect 36866 -5862 36880 -5834
rect 37284 -5842 37290 -5686
rect 32852 -5912 33060 -5906
rect 32852 -5946 32864 -5912
rect 33048 -5946 33060 -5912
rect 32852 -5952 33060 -5946
rect 33310 -5912 33518 -5906
rect 33310 -5946 33322 -5912
rect 33506 -5946 33518 -5912
rect 33310 -5952 33518 -5946
rect 33768 -5912 33976 -5906
rect 33768 -5946 33780 -5912
rect 33964 -5946 33976 -5912
rect 33768 -5952 33976 -5946
rect 34226 -5912 34434 -5906
rect 34226 -5946 34238 -5912
rect 34422 -5946 34434 -5912
rect 34226 -5952 34434 -5946
rect 34684 -5912 34892 -5906
rect 34684 -5946 34696 -5912
rect 34880 -5946 34892 -5912
rect 34684 -5952 34892 -5946
rect 35142 -5912 35350 -5906
rect 35142 -5946 35154 -5912
rect 35338 -5946 35350 -5912
rect 35142 -5952 35350 -5946
rect 35600 -5912 35808 -5906
rect 35600 -5946 35612 -5912
rect 35796 -5946 35808 -5912
rect 35600 -5952 35808 -5946
rect 36058 -5912 36266 -5906
rect 36058 -5946 36070 -5912
rect 36254 -5946 36266 -5912
rect 36058 -5952 36266 -5946
rect 36516 -5912 36724 -5906
rect 36516 -5946 36528 -5912
rect 36712 -5946 36724 -5912
rect 36516 -5952 36724 -5946
rect 32928 -6264 32988 -5952
rect 33384 -6018 33444 -5952
rect 33840 -6018 33900 -5952
rect 34306 -6018 34366 -5952
rect 34756 -6018 34816 -5952
rect 35210 -6018 35270 -5952
rect 35672 -6018 35732 -5952
rect 36126 -6018 36186 -5952
rect 36588 -6018 36648 -5952
rect 33384 -6078 36648 -6018
rect 33390 -6198 36654 -6138
rect 33390 -6264 33450 -6198
rect 33846 -6264 33906 -6198
rect 34312 -6264 34372 -6198
rect 34762 -6264 34822 -6198
rect 35216 -6264 35276 -6198
rect 35678 -6264 35738 -6198
rect 36132 -6264 36192 -6198
rect 36594 -6264 36654 -6198
rect 32852 -6270 33060 -6264
rect 32852 -6304 32864 -6270
rect 33048 -6304 33060 -6270
rect 32852 -6310 33060 -6304
rect 33310 -6270 33518 -6264
rect 33310 -6304 33322 -6270
rect 33506 -6304 33518 -6270
rect 33310 -6310 33518 -6304
rect 33768 -6270 33976 -6264
rect 33768 -6304 33780 -6270
rect 33964 -6304 33976 -6270
rect 33768 -6310 33976 -6304
rect 34226 -6270 34434 -6264
rect 34226 -6304 34238 -6270
rect 34422 -6304 34434 -6270
rect 34226 -6310 34434 -6304
rect 34684 -6270 34892 -6264
rect 34684 -6304 34696 -6270
rect 34880 -6304 34892 -6270
rect 34684 -6310 34892 -6304
rect 35142 -6270 35350 -6264
rect 35142 -6304 35154 -6270
rect 35338 -6304 35350 -6270
rect 35142 -6310 35350 -6304
rect 35600 -6270 35808 -6264
rect 35600 -6304 35612 -6270
rect 35796 -6304 35808 -6270
rect 35600 -6310 35808 -6304
rect 36058 -6270 36266 -6264
rect 36058 -6304 36070 -6270
rect 36254 -6304 36266 -6270
rect 36058 -6310 36266 -6304
rect 36516 -6270 36724 -6264
rect 36516 -6304 36528 -6270
rect 36712 -6304 36724 -6270
rect 36516 -6310 36724 -6304
rect 32324 -6494 32330 -6390
rect 32696 -6410 32710 -6354
rect 32324 -6530 32336 -6494
rect 32704 -6502 32710 -6410
rect 31974 -6580 32182 -6574
rect 31974 -6614 31986 -6580
rect 32170 -6614 32182 -6580
rect 31974 -6620 32182 -6614
rect 32042 -6966 32102 -6620
rect 32276 -6966 32336 -6530
rect 32696 -6530 32710 -6502
rect 32744 -6410 32756 -6354
rect 33162 -6354 33208 -6342
rect 32744 -6502 32750 -6410
rect 33162 -6500 33168 -6354
rect 32744 -6530 32756 -6502
rect 32696 -6966 32756 -6530
rect 33156 -6530 33168 -6500
rect 33202 -6500 33208 -6354
rect 33620 -6354 33666 -6342
rect 33202 -6530 33216 -6500
rect 32852 -6580 33060 -6574
rect 32852 -6614 32864 -6580
rect 33048 -6614 33060 -6580
rect 32852 -6620 33060 -6614
rect 32928 -6966 32988 -6620
rect 33156 -6814 33216 -6530
rect 33620 -6530 33626 -6354
rect 33660 -6530 33666 -6354
rect 33620 -6542 33666 -6530
rect 34078 -6354 34124 -6342
rect 34078 -6530 34084 -6354
rect 34118 -6530 34124 -6354
rect 34078 -6542 34124 -6530
rect 34536 -6354 34582 -6342
rect 34536 -6530 34542 -6354
rect 34576 -6530 34582 -6354
rect 34536 -6542 34582 -6530
rect 34994 -6354 35040 -6342
rect 34994 -6530 35000 -6354
rect 35034 -6530 35040 -6354
rect 34994 -6542 35040 -6530
rect 35452 -6354 35498 -6342
rect 35452 -6530 35458 -6354
rect 35492 -6530 35498 -6354
rect 35452 -6542 35498 -6530
rect 35910 -6354 35956 -6342
rect 35910 -6530 35916 -6354
rect 35950 -6530 35956 -6354
rect 35910 -6542 35956 -6530
rect 36368 -6354 36414 -6342
rect 36368 -6530 36374 -6354
rect 36408 -6530 36414 -6354
rect 36820 -6354 36880 -5862
rect 37276 -5862 37290 -5842
rect 37324 -5716 37344 -5686
rect 37324 -5842 37330 -5716
rect 37324 -5862 37336 -5842
rect 36974 -5912 37182 -5906
rect 36974 -5946 36986 -5912
rect 37170 -5946 37182 -5912
rect 36974 -5952 37182 -5946
rect 37048 -6078 37108 -5952
rect 37276 -6078 37336 -5862
rect 37048 -6138 37336 -6078
rect 37048 -6264 37108 -6138
rect 36974 -6270 37182 -6264
rect 36974 -6304 36986 -6270
rect 37170 -6304 37182 -6270
rect 36974 -6310 37182 -6304
rect 36820 -6396 36832 -6354
rect 36368 -6542 36414 -6530
rect 36826 -6530 36832 -6396
rect 36866 -6396 36880 -6354
rect 37276 -6354 37336 -6138
rect 37276 -6394 37290 -6354
rect 36866 -6530 36872 -6396
rect 37284 -6490 37290 -6394
rect 36826 -6542 36872 -6530
rect 37276 -6530 37290 -6490
rect 37324 -6394 37336 -6354
rect 37324 -6490 37330 -6394
rect 37324 -6530 37336 -6490
rect 33310 -6580 33518 -6574
rect 33310 -6614 33322 -6580
rect 33506 -6614 33518 -6580
rect 33310 -6620 33518 -6614
rect 33768 -6580 33976 -6574
rect 33768 -6614 33780 -6580
rect 33964 -6614 33976 -6580
rect 33768 -6620 33976 -6614
rect 34226 -6580 34434 -6574
rect 34226 -6614 34238 -6580
rect 34422 -6614 34434 -6580
rect 34226 -6620 34434 -6614
rect 34684 -6580 34892 -6574
rect 34684 -6614 34696 -6580
rect 34880 -6614 34892 -6580
rect 34684 -6620 34892 -6614
rect 35142 -6580 35350 -6574
rect 35142 -6614 35154 -6580
rect 35338 -6614 35350 -6580
rect 35142 -6620 35350 -6614
rect 35600 -6580 35808 -6574
rect 35600 -6614 35612 -6580
rect 35796 -6614 35808 -6580
rect 35600 -6620 35808 -6614
rect 36058 -6580 36266 -6574
rect 36058 -6614 36070 -6580
rect 36254 -6614 36266 -6580
rect 36058 -6620 36266 -6614
rect 36516 -6580 36724 -6574
rect 36516 -6614 36528 -6580
rect 36712 -6614 36724 -6580
rect 36516 -6620 36724 -6614
rect 36974 -6580 37182 -6574
rect 36974 -6614 36986 -6580
rect 37170 -6614 37182 -6580
rect 36974 -6620 37182 -6614
rect 33384 -6686 33450 -6620
rect 33840 -6680 33906 -6620
rect 33840 -6686 33846 -6680
rect 33384 -6746 33390 -6686
rect 33450 -6740 33846 -6686
rect 33906 -6686 33912 -6680
rect 34306 -6686 34372 -6620
rect 34756 -6686 34822 -6620
rect 35210 -6686 35276 -6620
rect 35672 -6680 35738 -6620
rect 35672 -6686 35678 -6680
rect 33906 -6740 34312 -6686
rect 33450 -6746 34312 -6740
rect 34372 -6746 34762 -6686
rect 34822 -6746 35216 -6686
rect 35276 -6740 35678 -6686
rect 35738 -6686 35744 -6680
rect 36126 -6686 36192 -6620
rect 36588 -6680 36654 -6620
rect 36588 -6686 36594 -6680
rect 35738 -6740 36132 -6686
rect 35276 -6746 36132 -6740
rect 36192 -6740 36594 -6686
rect 36654 -6740 36660 -6680
rect 36192 -6746 36648 -6740
rect 33156 -6880 33216 -6874
rect 37046 -6966 37106 -6620
rect 37276 -6966 37336 -6530
rect 37644 -6842 37650 -4838
rect 37750 -6842 37756 -4838
rect 37644 -6966 37756 -6842
rect 27300 -6972 37756 -6966
rect 27300 -7072 27406 -6972
rect 37650 -7072 37756 -6972
rect 27300 -7078 37756 -7072
rect 27300 -7308 37756 -7302
rect 27300 -7408 27406 -7308
rect 37650 -7408 37756 -7308
rect 27300 -7414 37756 -7408
rect 27300 -7590 27412 -7414
rect 27300 -12762 27306 -7590
rect 27406 -9384 27412 -7590
rect 27698 -7847 27758 -7414
rect 27926 -7748 27986 -7414
rect 28156 -7488 28216 -7482
rect 27851 -7754 28059 -7748
rect 27851 -7788 27863 -7754
rect 28047 -7788 28059 -7754
rect 27851 -7794 28059 -7788
rect 27698 -7880 27709 -7847
rect 27703 -8970 27709 -7880
rect 27700 -9023 27709 -8970
rect 27743 -7880 27758 -7847
rect 28156 -7847 28216 -7548
rect 28388 -7618 28448 -7612
rect 28844 -7618 28904 -7612
rect 29760 -7618 29820 -7612
rect 28448 -7678 28844 -7620
rect 29310 -7620 29370 -7618
rect 28904 -7624 29760 -7620
rect 28904 -7678 29310 -7624
rect 28388 -7680 29310 -7678
rect 28388 -7748 28448 -7680
rect 28844 -7748 28904 -7680
rect 29370 -7678 29760 -7624
rect 30214 -7618 30274 -7612
rect 29820 -7678 30214 -7620
rect 30676 -7618 30736 -7612
rect 31592 -7616 31652 -7610
rect 30274 -7678 30676 -7620
rect 31130 -7620 31190 -7618
rect 30736 -7624 31592 -7620
rect 30736 -7678 31130 -7624
rect 29370 -7680 31130 -7678
rect 29310 -7748 29370 -7684
rect 29760 -7748 29820 -7680
rect 30214 -7748 30274 -7680
rect 30676 -7748 30736 -7680
rect 31190 -7676 31592 -7624
rect 31190 -7680 31652 -7676
rect 31130 -7748 31190 -7684
rect 31592 -7748 31652 -7680
rect 28309 -7754 28517 -7748
rect 28309 -7788 28321 -7754
rect 28505 -7788 28517 -7754
rect 28309 -7794 28517 -7788
rect 28767 -7754 28975 -7748
rect 28767 -7788 28779 -7754
rect 28963 -7788 28975 -7754
rect 28767 -7794 28975 -7788
rect 29225 -7754 29433 -7748
rect 29225 -7788 29237 -7754
rect 29421 -7788 29433 -7754
rect 29225 -7794 29433 -7788
rect 29683 -7754 29891 -7748
rect 29683 -7788 29695 -7754
rect 29879 -7788 29891 -7754
rect 29683 -7794 29891 -7788
rect 30141 -7754 30349 -7748
rect 30141 -7788 30153 -7754
rect 30337 -7788 30349 -7754
rect 30141 -7794 30349 -7788
rect 30599 -7754 30807 -7748
rect 30599 -7788 30611 -7754
rect 30795 -7788 30807 -7754
rect 30599 -7794 30807 -7788
rect 31057 -7754 31265 -7748
rect 31057 -7788 31069 -7754
rect 31253 -7788 31265 -7754
rect 31057 -7794 31265 -7788
rect 31515 -7754 31723 -7748
rect 31515 -7788 31527 -7754
rect 31711 -7788 31723 -7754
rect 31515 -7794 31723 -7788
rect 28156 -7854 28167 -7847
rect 27743 -8970 27749 -7880
rect 27743 -9023 27760 -8970
rect 27700 -9384 27760 -9023
rect 28161 -9023 28167 -7854
rect 28201 -7854 28216 -7847
rect 28619 -7847 28665 -7835
rect 28201 -9023 28207 -7854
rect 28161 -9035 28207 -9023
rect 28619 -9023 28625 -7847
rect 28659 -9023 28665 -7847
rect 28619 -9035 28665 -9023
rect 29077 -7847 29123 -7835
rect 29077 -9023 29083 -7847
rect 29117 -9023 29123 -7847
rect 29077 -9035 29123 -9023
rect 29535 -7847 29581 -7835
rect 29535 -9023 29541 -7847
rect 29575 -9023 29581 -7847
rect 29535 -9035 29581 -9023
rect 29993 -7847 30039 -7835
rect 29993 -9023 29999 -7847
rect 30033 -9023 30039 -7847
rect 29993 -9035 30039 -9023
rect 30451 -7847 30497 -7835
rect 30451 -9023 30457 -7847
rect 30491 -9023 30497 -7847
rect 30451 -9035 30497 -9023
rect 30909 -7847 30955 -7835
rect 30909 -9023 30915 -7847
rect 30949 -9023 30955 -7847
rect 30909 -9035 30955 -9023
rect 31367 -7847 31413 -7835
rect 31367 -9023 31373 -7847
rect 31407 -9023 31413 -7847
rect 31820 -7847 31880 -7414
rect 32050 -7748 32110 -7414
rect 31973 -7754 32181 -7748
rect 31973 -7788 31985 -7754
rect 32169 -7788 32181 -7754
rect 31973 -7794 32181 -7788
rect 31820 -7888 31831 -7847
rect 31825 -8980 31831 -7888
rect 31367 -9035 31413 -9023
rect 31818 -9023 31831 -8980
rect 31865 -7888 31880 -7847
rect 32278 -7847 32338 -7414
rect 32278 -7882 32289 -7847
rect 31865 -8980 31871 -7888
rect 31865 -9023 31878 -8980
rect 32283 -9002 32289 -7882
rect 27851 -9082 28059 -9076
rect 27851 -9116 27863 -9082
rect 28047 -9116 28059 -9082
rect 27851 -9122 28059 -9116
rect 28309 -9082 28517 -9076
rect 28309 -9116 28321 -9082
rect 28505 -9116 28517 -9082
rect 28309 -9122 28517 -9116
rect 28767 -9082 28975 -9076
rect 28767 -9116 28779 -9082
rect 28963 -9116 28975 -9082
rect 28767 -9122 28975 -9116
rect 29225 -9082 29433 -9076
rect 29225 -9116 29237 -9082
rect 29421 -9116 29433 -9082
rect 29225 -9122 29433 -9116
rect 29683 -9082 29891 -9076
rect 29683 -9116 29695 -9082
rect 29879 -9116 29891 -9082
rect 29683 -9122 29891 -9116
rect 30141 -9082 30349 -9076
rect 30141 -9116 30153 -9082
rect 30337 -9116 30349 -9082
rect 30141 -9122 30349 -9116
rect 30599 -9082 30807 -9076
rect 30599 -9116 30611 -9082
rect 30795 -9116 30807 -9082
rect 30599 -9122 30807 -9116
rect 31057 -9082 31265 -9076
rect 31057 -9116 31069 -9082
rect 31253 -9116 31265 -9082
rect 31057 -9122 31265 -9116
rect 31515 -9082 31723 -9076
rect 31515 -9116 31527 -9082
rect 31711 -9116 31723 -9082
rect 31515 -9122 31723 -9116
rect 27926 -9384 27986 -9122
rect 28388 -9192 28448 -9122
rect 28844 -9192 28904 -9122
rect 29310 -9192 29370 -9122
rect 29760 -9192 29820 -9122
rect 30214 -9192 30274 -9122
rect 30676 -9192 30736 -9122
rect 31130 -9192 31190 -9122
rect 31592 -9192 31652 -9122
rect 28388 -9252 31652 -9192
rect 31818 -9174 31878 -9023
rect 32276 -9023 32289 -9002
rect 32323 -7882 32338 -7847
rect 32698 -7847 32758 -7414
rect 32926 -7748 32986 -7414
rect 33150 -7554 33156 -7494
rect 33216 -7554 33222 -7494
rect 32851 -7754 33059 -7748
rect 32851 -7788 32863 -7754
rect 33047 -7788 33059 -7754
rect 32851 -7794 33059 -7788
rect 32698 -7882 32709 -7847
rect 32323 -9002 32329 -7882
rect 32323 -9023 32336 -9002
rect 32703 -9008 32709 -7882
rect 31973 -9082 32181 -9076
rect 31973 -9116 31985 -9082
rect 32169 -9116 32181 -9082
rect 31973 -9122 32181 -9116
rect 32044 -9174 32104 -9122
rect 32276 -9174 32336 -9023
rect 32696 -9023 32709 -9008
rect 32743 -7882 32758 -7847
rect 33156 -7847 33216 -7554
rect 33390 -7616 33450 -7610
rect 34762 -7614 34822 -7608
rect 33846 -7620 33906 -7614
rect 34312 -7620 34372 -7614
rect 33450 -7676 33846 -7620
rect 33390 -7680 33846 -7676
rect 33906 -7680 34312 -7620
rect 34372 -7674 34762 -7620
rect 35216 -7620 35276 -7614
rect 35678 -7620 35738 -7614
rect 36132 -7616 36192 -7610
rect 34822 -7674 35216 -7620
rect 34372 -7680 35216 -7674
rect 35276 -7680 35678 -7620
rect 35738 -7676 36132 -7620
rect 36594 -7616 36654 -7610
rect 36192 -7676 36594 -7620
rect 35738 -7680 36654 -7676
rect 33390 -7748 33450 -7680
rect 33846 -7748 33906 -7680
rect 34312 -7748 34372 -7680
rect 34762 -7748 34822 -7680
rect 35216 -7748 35276 -7680
rect 35678 -7748 35738 -7680
rect 36132 -7748 36192 -7680
rect 36594 -7748 36654 -7680
rect 37048 -7748 37108 -7414
rect 33309 -7754 33517 -7748
rect 33309 -7788 33321 -7754
rect 33505 -7788 33517 -7754
rect 33309 -7794 33517 -7788
rect 33767 -7754 33975 -7748
rect 33767 -7788 33779 -7754
rect 33963 -7788 33975 -7754
rect 33767 -7794 33975 -7788
rect 34225 -7754 34433 -7748
rect 34225 -7788 34237 -7754
rect 34421 -7788 34433 -7754
rect 34225 -7794 34433 -7788
rect 34683 -7754 34891 -7748
rect 34683 -7788 34695 -7754
rect 34879 -7788 34891 -7754
rect 34683 -7794 34891 -7788
rect 35141 -7754 35349 -7748
rect 35141 -7788 35153 -7754
rect 35337 -7788 35349 -7754
rect 35141 -7794 35349 -7788
rect 35599 -7754 35807 -7748
rect 35599 -7788 35611 -7754
rect 35795 -7788 35807 -7754
rect 35599 -7794 35807 -7788
rect 36057 -7754 36265 -7748
rect 36057 -7788 36069 -7754
rect 36253 -7788 36265 -7754
rect 36057 -7794 36265 -7788
rect 36515 -7754 36723 -7748
rect 36515 -7788 36527 -7754
rect 36711 -7788 36723 -7754
rect 36515 -7794 36723 -7788
rect 36973 -7754 37181 -7748
rect 36973 -7788 36985 -7754
rect 37169 -7788 37181 -7754
rect 36973 -7794 37181 -7788
rect 32743 -9008 32749 -7882
rect 33156 -7914 33167 -7847
rect 32743 -9023 32756 -9008
rect 32696 -9174 32756 -9023
rect 33161 -9023 33167 -7914
rect 33201 -7914 33216 -7847
rect 33619 -7847 33665 -7835
rect 33201 -9023 33207 -7914
rect 33161 -9035 33207 -9023
rect 33619 -9023 33625 -7847
rect 33659 -9023 33665 -7847
rect 33619 -9035 33665 -9023
rect 34077 -7847 34123 -7835
rect 34077 -9023 34083 -7847
rect 34117 -9023 34123 -7847
rect 34077 -9035 34123 -9023
rect 34535 -7847 34581 -7835
rect 34535 -9023 34541 -7847
rect 34575 -9023 34581 -7847
rect 34535 -9035 34581 -9023
rect 34993 -7847 35039 -7835
rect 34993 -9023 34999 -7847
rect 35033 -9023 35039 -7847
rect 34993 -9035 35039 -9023
rect 35451 -7847 35497 -7835
rect 35451 -9023 35457 -7847
rect 35491 -9023 35497 -7847
rect 35451 -9035 35497 -9023
rect 35909 -7847 35955 -7835
rect 35909 -9023 35915 -7847
rect 35949 -9023 35955 -7847
rect 35909 -9035 35955 -9023
rect 36367 -7847 36413 -7835
rect 36367 -9023 36373 -7847
rect 36407 -9023 36413 -7847
rect 36825 -7847 36871 -7835
rect 36825 -8956 36831 -7847
rect 36367 -9035 36413 -9023
rect 36818 -9023 36831 -8956
rect 36865 -8956 36871 -7847
rect 37276 -7847 37336 -7414
rect 37276 -7868 37289 -7847
rect 36865 -9023 36878 -8956
rect 37283 -8976 37289 -7868
rect 32851 -9082 33059 -9076
rect 32851 -9116 32863 -9082
rect 33047 -9116 33059 -9082
rect 32851 -9122 33059 -9116
rect 33309 -9082 33517 -9076
rect 33309 -9116 33321 -9082
rect 33505 -9116 33517 -9082
rect 33309 -9122 33517 -9116
rect 33767 -9082 33975 -9076
rect 33767 -9116 33779 -9082
rect 33963 -9116 33975 -9082
rect 33767 -9122 33975 -9116
rect 34225 -9082 34433 -9076
rect 34225 -9116 34237 -9082
rect 34421 -9116 34433 -9082
rect 34225 -9122 34433 -9116
rect 34683 -9082 34891 -9076
rect 34683 -9116 34695 -9082
rect 34879 -9116 34891 -9082
rect 34683 -9122 34891 -9116
rect 35141 -9082 35349 -9076
rect 35141 -9116 35153 -9082
rect 35337 -9116 35349 -9082
rect 35141 -9122 35349 -9116
rect 35599 -9082 35807 -9076
rect 35599 -9116 35611 -9082
rect 35795 -9116 35807 -9082
rect 35599 -9122 35807 -9116
rect 36057 -9082 36265 -9076
rect 36057 -9116 36069 -9082
rect 36253 -9116 36265 -9082
rect 36057 -9122 36265 -9116
rect 36515 -9082 36723 -9076
rect 36515 -9116 36527 -9082
rect 36711 -9116 36723 -9082
rect 36515 -9122 36723 -9116
rect 32926 -9174 32986 -9122
rect 31818 -9234 32986 -9174
rect 33382 -9192 33442 -9122
rect 33838 -9192 33898 -9122
rect 34304 -9192 34364 -9122
rect 34754 -9192 34814 -9122
rect 35208 -9192 35268 -9122
rect 35670 -9192 35730 -9122
rect 36124 -9192 36184 -9122
rect 36586 -9192 36646 -9122
rect 33382 -9252 36646 -9192
rect 36818 -9294 36878 -9023
rect 37276 -9023 37289 -8976
rect 37323 -7868 37336 -7847
rect 37644 -7590 37756 -7414
rect 37323 -8976 37329 -7868
rect 37323 -9023 37336 -8976
rect 36973 -9082 37181 -9076
rect 36973 -9116 36985 -9082
rect 37169 -9116 37181 -9082
rect 36973 -9122 37181 -9116
rect 36812 -9354 36818 -9294
rect 36878 -9354 36884 -9294
rect 27406 -9444 28536 -9384
rect 27406 -9878 27412 -9444
rect 28476 -9878 28536 -9444
rect 29388 -9460 35864 -9400
rect 37048 -9448 37108 -9122
rect 37276 -9448 37336 -9023
rect 37644 -9448 37650 -7590
rect 27406 -9938 28994 -9878
rect 27406 -12762 27412 -9938
rect 28476 -10112 28536 -9938
rect 28702 -10013 28762 -9938
rect 28628 -10019 28836 -10013
rect 28628 -10053 28640 -10019
rect 28824 -10053 28836 -10019
rect 28628 -10059 28836 -10053
rect 28476 -10156 28486 -10112
rect 28480 -11618 28486 -10156
rect 28472 -11688 28486 -11618
rect 28520 -10156 28536 -10112
rect 28934 -10112 28994 -9938
rect 29158 -9940 29164 -9880
rect 29224 -9940 29230 -9880
rect 29164 -10013 29224 -9940
rect 29086 -10019 29294 -10013
rect 29086 -10053 29098 -10019
rect 29282 -10053 29294 -10019
rect 29086 -10059 29294 -10053
rect 28520 -11618 28526 -10156
rect 28934 -10174 28944 -10112
rect 28938 -11612 28944 -10174
rect 28520 -11688 28532 -11618
rect 28472 -12476 28532 -11688
rect 28930 -11688 28944 -11612
rect 28978 -10174 28994 -10112
rect 29388 -10112 29448 -9460
rect 30302 -9590 34946 -9530
rect 29618 -9940 29624 -9880
rect 29684 -9940 29690 -9880
rect 30076 -9940 30082 -9880
rect 30142 -9940 30148 -9880
rect 29624 -10013 29684 -9940
rect 30082 -10013 30142 -9940
rect 29544 -10019 29752 -10013
rect 29544 -10053 29556 -10019
rect 29740 -10053 29752 -10019
rect 29544 -10059 29752 -10053
rect 30002 -10019 30210 -10013
rect 30002 -10053 30014 -10019
rect 30198 -10053 30210 -10019
rect 30002 -10059 30210 -10053
rect 29388 -10172 29402 -10112
rect 28978 -11612 28984 -10174
rect 28978 -11688 28990 -11612
rect 28628 -11747 28836 -11741
rect 28628 -11781 28640 -11747
rect 28824 -11781 28836 -11747
rect 28628 -11787 28836 -11781
rect 28700 -12476 28760 -11787
rect 28930 -12476 28990 -11688
rect 29396 -11688 29402 -10172
rect 29436 -10172 29448 -10112
rect 29854 -10112 29900 -10100
rect 29436 -11688 29442 -10172
rect 29854 -11632 29860 -10112
rect 29396 -11700 29442 -11688
rect 29846 -11688 29860 -11632
rect 29894 -11632 29900 -10112
rect 30302 -10112 30362 -9590
rect 31222 -9716 34038 -9656
rect 30532 -9940 30538 -9880
rect 30598 -9940 30604 -9880
rect 30988 -9940 30994 -9880
rect 31054 -9940 31060 -9880
rect 30538 -10013 30598 -9940
rect 30994 -10013 31054 -9940
rect 30460 -10019 30668 -10013
rect 30460 -10053 30472 -10019
rect 30656 -10053 30668 -10019
rect 30460 -10059 30668 -10053
rect 30918 -10019 31126 -10013
rect 30918 -10053 30930 -10019
rect 31114 -10053 31126 -10019
rect 30918 -10059 31126 -10053
rect 30302 -10180 30318 -10112
rect 29894 -11688 29906 -11632
rect 29086 -11747 29294 -11741
rect 29086 -11781 29098 -11747
rect 29282 -11781 29294 -11747
rect 29086 -11787 29294 -11781
rect 29544 -11747 29752 -11741
rect 29544 -11781 29556 -11747
rect 29740 -11781 29752 -11747
rect 29544 -11787 29752 -11781
rect 29160 -11854 29220 -11787
rect 29620 -11854 29680 -11787
rect 29154 -11914 29160 -11854
rect 29220 -11914 29226 -11854
rect 29614 -11914 29620 -11854
rect 29680 -11914 29686 -11854
rect 29846 -12222 29906 -11688
rect 30312 -11688 30318 -10180
rect 30352 -10180 30362 -10112
rect 30770 -10112 30816 -10100
rect 30352 -11688 30358 -10180
rect 30770 -11630 30776 -10112
rect 30312 -11700 30358 -11688
rect 30766 -11688 30776 -11630
rect 30810 -11630 30816 -10112
rect 31222 -10112 31282 -9716
rect 32136 -9832 33114 -9772
rect 31444 -9940 31450 -9880
rect 31510 -9940 31516 -9880
rect 31904 -9940 31910 -9880
rect 31970 -9940 31976 -9880
rect 31450 -10013 31510 -9940
rect 31910 -10013 31970 -9940
rect 31376 -10019 31584 -10013
rect 31376 -10053 31388 -10019
rect 31572 -10053 31584 -10019
rect 31376 -10059 31584 -10053
rect 31834 -10019 32042 -10013
rect 31834 -10053 31846 -10019
rect 32030 -10053 32042 -10019
rect 31834 -10059 32042 -10053
rect 31222 -10144 31234 -10112
rect 30810 -11688 30826 -11630
rect 30002 -11747 30210 -11741
rect 30002 -11781 30014 -11747
rect 30198 -11781 30210 -11747
rect 30002 -11787 30210 -11781
rect 30460 -11747 30668 -11741
rect 30460 -11781 30472 -11747
rect 30656 -11781 30668 -11747
rect 30460 -11787 30668 -11781
rect 30078 -11854 30138 -11787
rect 30534 -11854 30594 -11787
rect 30072 -11914 30078 -11854
rect 30138 -11914 30144 -11854
rect 30528 -11914 30534 -11854
rect 30594 -11914 30600 -11854
rect 30766 -12088 30826 -11688
rect 31228 -11688 31234 -10144
rect 31268 -10144 31282 -10112
rect 31686 -10112 31732 -10100
rect 31268 -11688 31274 -10144
rect 31686 -11644 31692 -10112
rect 31228 -11700 31274 -11688
rect 31682 -11688 31692 -11644
rect 31726 -11644 31732 -10112
rect 32136 -10112 32196 -9832
rect 32354 -9880 32438 -9876
rect 32354 -9942 32366 -9880
rect 32426 -9942 32438 -9880
rect 32354 -9948 32438 -9942
rect 32592 -9892 32652 -9886
rect 32366 -10013 32426 -9948
rect 32820 -9940 32826 -9880
rect 32886 -9940 32892 -9880
rect 32820 -9942 32892 -9940
rect 32292 -10019 32500 -10013
rect 32292 -10053 32304 -10019
rect 32488 -10053 32500 -10019
rect 32292 -10059 32500 -10053
rect 32136 -10140 32150 -10112
rect 31726 -11688 31742 -11644
rect 30918 -11747 31126 -11741
rect 30918 -11781 30930 -11747
rect 31114 -11781 31126 -11747
rect 30918 -11787 31126 -11781
rect 31376 -11747 31584 -11741
rect 31376 -11781 31388 -11747
rect 31572 -11781 31584 -11747
rect 31376 -11787 31584 -11781
rect 30990 -11854 31050 -11787
rect 31446 -11854 31506 -11787
rect 30984 -11914 30990 -11854
rect 31050 -11914 31056 -11854
rect 31440 -11914 31446 -11854
rect 31506 -11914 31512 -11854
rect 31682 -11964 31742 -11688
rect 32144 -11688 32150 -10140
rect 32184 -10140 32196 -10112
rect 32592 -10112 32652 -9952
rect 32826 -10013 32886 -9942
rect 32750 -10019 32958 -10013
rect 32750 -10053 32762 -10019
rect 32946 -10053 32958 -10019
rect 32750 -10059 32958 -10053
rect 32592 -10134 32608 -10112
rect 32184 -11688 32190 -10140
rect 32144 -11700 32190 -11688
rect 32602 -11688 32608 -10134
rect 32642 -10134 32652 -10112
rect 33054 -10112 33114 -9832
rect 33278 -9940 33284 -9880
rect 33344 -9940 33350 -9880
rect 33732 -9940 33738 -9880
rect 33798 -9940 33804 -9880
rect 33284 -10013 33344 -9940
rect 33738 -10013 33798 -9940
rect 33208 -10019 33416 -10013
rect 33208 -10053 33220 -10019
rect 33404 -10053 33416 -10019
rect 33208 -10059 33416 -10053
rect 33666 -10019 33874 -10013
rect 33666 -10053 33678 -10019
rect 33862 -10053 33874 -10019
rect 33666 -10059 33874 -10053
rect 33978 -10100 34038 -9716
rect 34196 -9940 34202 -9880
rect 34262 -9940 34268 -9880
rect 34654 -9940 34660 -9880
rect 34720 -9940 34726 -9880
rect 34202 -10013 34262 -9940
rect 34660 -10013 34720 -9940
rect 34124 -10019 34332 -10013
rect 34124 -10053 34136 -10019
rect 34320 -10053 34332 -10019
rect 34124 -10059 34332 -10053
rect 34582 -10019 34790 -10013
rect 34582 -10053 34594 -10019
rect 34778 -10053 34790 -10019
rect 34582 -10059 34790 -10053
rect 32642 -11688 32648 -10134
rect 33054 -10192 33066 -10112
rect 32602 -11700 32648 -11688
rect 33060 -11688 33066 -10192
rect 33100 -10192 33114 -10112
rect 33518 -10112 33564 -10100
rect 33100 -11688 33106 -10192
rect 33518 -11610 33524 -10112
rect 33060 -11700 33106 -11688
rect 33512 -11688 33524 -11610
rect 33558 -11610 33564 -10112
rect 33976 -10112 34038 -10100
rect 33558 -11688 33572 -11610
rect 31834 -11747 32042 -11741
rect 31834 -11781 31846 -11747
rect 32030 -11781 32042 -11747
rect 31834 -11787 32042 -11781
rect 32292 -11747 32500 -11741
rect 32292 -11781 32304 -11747
rect 32488 -11781 32500 -11747
rect 32292 -11787 32500 -11781
rect 32750 -11747 32958 -11741
rect 32750 -11781 32762 -11747
rect 32946 -11781 32958 -11747
rect 32750 -11787 32958 -11781
rect 33208 -11747 33416 -11741
rect 33208 -11781 33220 -11747
rect 33404 -11781 33416 -11747
rect 33208 -11787 33416 -11781
rect 31902 -11854 31962 -11787
rect 32360 -11854 32420 -11787
rect 32828 -11854 32888 -11787
rect 33284 -11854 33344 -11787
rect 31896 -11914 31902 -11854
rect 31962 -11914 31968 -11854
rect 32354 -11914 32360 -11854
rect 32420 -11914 32426 -11854
rect 32822 -11914 32828 -11854
rect 32888 -11914 32894 -11854
rect 33278 -11914 33284 -11854
rect 33344 -11914 33350 -11854
rect 33512 -11964 33572 -11688
rect 33976 -11688 33982 -10112
rect 34016 -10184 34038 -10112
rect 34434 -10112 34480 -10100
rect 34016 -11688 34022 -10184
rect 34434 -11628 34440 -10112
rect 33976 -11700 34022 -11688
rect 34428 -11688 34440 -11628
rect 34474 -11628 34480 -10112
rect 34886 -10112 34946 -9590
rect 35110 -9940 35116 -9880
rect 35176 -9940 35182 -9880
rect 35570 -9940 35576 -9880
rect 35636 -9940 35642 -9880
rect 35116 -10013 35176 -9940
rect 35576 -10013 35636 -9940
rect 35040 -10019 35248 -10013
rect 35040 -10053 35052 -10019
rect 35236 -10053 35248 -10019
rect 35040 -10059 35248 -10053
rect 35498 -10019 35706 -10013
rect 35498 -10053 35510 -10019
rect 35694 -10053 35706 -10019
rect 35498 -10059 35706 -10053
rect 34886 -10190 34898 -10112
rect 34474 -11688 34488 -11628
rect 33666 -11747 33874 -11741
rect 33666 -11781 33678 -11747
rect 33862 -11781 33874 -11747
rect 33666 -11787 33874 -11781
rect 34124 -11747 34332 -11741
rect 34124 -11781 34136 -11747
rect 34320 -11781 34332 -11747
rect 34124 -11787 34332 -11781
rect 33734 -11854 33794 -11787
rect 34198 -11854 34258 -11787
rect 33728 -11914 33734 -11854
rect 33794 -11914 33800 -11854
rect 34192 -11914 34198 -11854
rect 34258 -11914 34264 -11854
rect 31682 -12024 33572 -11964
rect 34428 -12088 34488 -11688
rect 34892 -11688 34898 -10190
rect 34932 -10190 34946 -10112
rect 35350 -10112 35396 -10100
rect 34932 -11688 34938 -10190
rect 35350 -11630 35356 -10112
rect 34892 -11700 34938 -11688
rect 35344 -11688 35356 -11630
rect 35390 -11630 35396 -10112
rect 35804 -10112 35864 -9460
rect 36716 -9508 37650 -9448
rect 36716 -9880 36776 -9508
rect 37644 -9880 37650 -9508
rect 36026 -9940 36032 -9880
rect 36092 -9940 36098 -9880
rect 36262 -9940 37650 -9880
rect 36032 -10013 36092 -9940
rect 35956 -10019 36164 -10013
rect 35956 -10053 35968 -10019
rect 36152 -10053 36164 -10019
rect 35956 -10059 36164 -10053
rect 35804 -10196 35814 -10112
rect 35390 -11688 35404 -11630
rect 34582 -11747 34790 -11741
rect 34582 -11781 34594 -11747
rect 34778 -11781 34790 -11747
rect 34582 -11787 34790 -11781
rect 35040 -11747 35248 -11741
rect 35040 -11781 35052 -11747
rect 35236 -11781 35248 -11747
rect 35040 -11787 35248 -11781
rect 34656 -11854 34716 -11787
rect 35112 -11854 35172 -11787
rect 34650 -11914 34656 -11854
rect 34716 -11914 34722 -11854
rect 35106 -11914 35112 -11854
rect 35172 -11914 35178 -11854
rect 30766 -12148 34488 -12088
rect 35344 -12222 35404 -11688
rect 35808 -11688 35814 -10196
rect 35848 -10196 35864 -10112
rect 36262 -10112 36322 -9940
rect 36488 -10013 36548 -9940
rect 36414 -10019 36622 -10013
rect 36414 -10053 36426 -10019
rect 36610 -10053 36622 -10019
rect 36414 -10059 36622 -10053
rect 36262 -10156 36272 -10112
rect 35848 -11688 35854 -10196
rect 36266 -11624 36272 -10156
rect 35808 -11700 35854 -11688
rect 36260 -11688 36272 -11624
rect 36306 -10156 36322 -10112
rect 36716 -10112 36776 -9940
rect 36306 -11624 36312 -10156
rect 36716 -10172 36730 -10112
rect 36306 -11688 36320 -11624
rect 36724 -11656 36730 -10172
rect 35498 -11747 35706 -11741
rect 35498 -11781 35510 -11747
rect 35694 -11781 35706 -11747
rect 35498 -11787 35706 -11781
rect 35956 -11747 36164 -11741
rect 35956 -11781 35968 -11747
rect 36152 -11781 36164 -11747
rect 35956 -11787 36164 -11781
rect 35572 -11854 35632 -11787
rect 36028 -11854 36088 -11787
rect 35566 -11914 35572 -11854
rect 35632 -11914 35638 -11854
rect 36022 -11914 36028 -11854
rect 36088 -11914 36094 -11854
rect 29846 -12282 35404 -12222
rect 36260 -12476 36320 -11688
rect 36718 -11688 36730 -11656
rect 36764 -10172 36776 -10112
rect 36764 -11656 36770 -10172
rect 36764 -11688 36778 -11656
rect 36414 -11747 36622 -11741
rect 36414 -11781 36426 -11747
rect 36610 -11781 36622 -11747
rect 36414 -11787 36622 -11781
rect 36486 -12476 36546 -11787
rect 36718 -12476 36778 -11688
rect 28450 -12486 36806 -12476
rect 28450 -12572 28476 -12486
rect 28572 -12572 28896 -12486
rect 28992 -12572 29496 -12486
rect 29592 -12572 30096 -12486
rect 30192 -12572 30696 -12486
rect 30792 -12572 31296 -12486
rect 31392 -12572 31896 -12486
rect 31992 -12572 32496 -12486
rect 32592 -12572 33096 -12486
rect 33192 -12572 33696 -12486
rect 33792 -12572 34296 -12486
rect 34392 -12572 34896 -12486
rect 34992 -12572 35496 -12486
rect 35592 -12572 36096 -12486
rect 36192 -12572 36696 -12486
rect 36792 -12572 36806 -12486
rect 28450 -12586 36806 -12572
rect 27300 -13046 27412 -12762
rect 28012 -13046 28022 -12746
rect 37034 -13046 37044 -12746
rect 37644 -12762 37650 -9940
rect 37750 -12762 37756 -7590
rect 37644 -13046 37756 -12762
rect 27300 -13052 37756 -13046
rect 27300 -13152 27406 -13052
rect 37650 -13152 37756 -13052
rect 27300 -13158 37756 -13152
rect 23346 -13604 33802 -13598
rect 23346 -13704 23452 -13604
rect 33696 -13704 33802 -13604
rect 23346 -13710 33802 -13704
rect 23346 -13994 23458 -13710
rect 23346 -19166 23352 -13994
rect 23452 -16816 23458 -13994
rect 24058 -14010 24068 -13710
rect 33080 -14010 33090 -13710
rect 33690 -13994 33802 -13710
rect 24296 -14184 32652 -14170
rect 24296 -14270 24310 -14184
rect 24406 -14270 24910 -14184
rect 25006 -14270 25510 -14184
rect 25606 -14270 26110 -14184
rect 26206 -14270 26710 -14184
rect 26806 -14270 27310 -14184
rect 27406 -14270 27910 -14184
rect 28006 -14270 28510 -14184
rect 28606 -14270 29110 -14184
rect 29206 -14270 29710 -14184
rect 29806 -14270 30310 -14184
rect 30406 -14270 30910 -14184
rect 31006 -14270 31510 -14184
rect 31606 -14270 32110 -14184
rect 32206 -14270 32530 -14184
rect 32626 -14270 32652 -14184
rect 24296 -14280 32652 -14270
rect 24324 -15068 24384 -14280
rect 24556 -14969 24616 -14280
rect 24480 -14975 24688 -14969
rect 24480 -15009 24492 -14975
rect 24676 -15009 24688 -14975
rect 24480 -15015 24688 -15009
rect 24324 -15100 24338 -15068
rect 24332 -16584 24338 -15100
rect 24326 -16644 24338 -16584
rect 24372 -15100 24384 -15068
rect 24782 -15068 24842 -14280
rect 25698 -14534 31256 -14474
rect 25008 -14902 25014 -14842
rect 25074 -14902 25080 -14842
rect 25464 -14902 25470 -14842
rect 25530 -14902 25536 -14842
rect 25014 -14969 25074 -14902
rect 25470 -14969 25530 -14902
rect 24938 -14975 25146 -14969
rect 24938 -15009 24950 -14975
rect 25134 -15009 25146 -14975
rect 24938 -15015 25146 -15009
rect 25396 -14975 25604 -14969
rect 25396 -15009 25408 -14975
rect 25592 -15009 25604 -14975
rect 25396 -15015 25604 -15009
rect 24372 -16584 24378 -15100
rect 24782 -15132 24796 -15068
rect 24372 -16644 24386 -16584
rect 24790 -16600 24796 -15132
rect 24326 -16816 24386 -16644
rect 24780 -16644 24796 -16600
rect 24830 -15132 24842 -15068
rect 25248 -15068 25294 -15056
rect 24830 -16600 24836 -15132
rect 25248 -16560 25254 -15068
rect 24830 -16644 24840 -16600
rect 24480 -16703 24688 -16697
rect 24480 -16737 24492 -16703
rect 24676 -16737 24688 -16703
rect 24480 -16743 24688 -16737
rect 24554 -16816 24614 -16743
rect 24780 -16816 24840 -16644
rect 25238 -16644 25254 -16560
rect 25288 -16560 25294 -15068
rect 25698 -15068 25758 -14534
rect 26614 -14668 30336 -14608
rect 25924 -14902 25930 -14842
rect 25990 -14902 25996 -14842
rect 26380 -14902 26386 -14842
rect 26446 -14902 26452 -14842
rect 25930 -14969 25990 -14902
rect 26386 -14969 26446 -14902
rect 25854 -14975 26062 -14969
rect 25854 -15009 25866 -14975
rect 26050 -15009 26062 -14975
rect 25854 -15015 26062 -15009
rect 26312 -14975 26520 -14969
rect 26312 -15009 26324 -14975
rect 26508 -15009 26520 -14975
rect 26312 -15015 26520 -15009
rect 25698 -15126 25712 -15068
rect 25288 -16644 25298 -16560
rect 24938 -16703 25146 -16697
rect 24938 -16737 24950 -16703
rect 25134 -16737 25146 -16703
rect 24938 -16743 25146 -16737
rect 25010 -16816 25070 -16743
rect 23452 -16876 24840 -16816
rect 25004 -16876 25010 -16816
rect 25070 -16876 25076 -16816
rect 23452 -17248 23458 -16876
rect 24326 -17248 24386 -16876
rect 23452 -17308 24386 -17248
rect 25238 -17296 25298 -16644
rect 25706 -16644 25712 -15126
rect 25746 -15126 25758 -15068
rect 26164 -15068 26210 -15056
rect 25746 -16644 25752 -15126
rect 26164 -16566 26170 -15068
rect 25706 -16656 25752 -16644
rect 26156 -16644 26170 -16566
rect 26204 -16566 26210 -15068
rect 26614 -15068 26674 -14668
rect 27530 -14792 29420 -14732
rect 26838 -14902 26844 -14842
rect 26904 -14902 26910 -14842
rect 27302 -14902 27308 -14842
rect 27368 -14902 27374 -14842
rect 26844 -14969 26904 -14902
rect 27308 -14969 27368 -14902
rect 26770 -14975 26978 -14969
rect 26770 -15009 26782 -14975
rect 26966 -15009 26978 -14975
rect 26770 -15015 26978 -15009
rect 27228 -14975 27436 -14969
rect 27228 -15009 27240 -14975
rect 27424 -15009 27436 -14975
rect 27228 -15015 27436 -15009
rect 26614 -15128 26628 -15068
rect 26204 -16644 26216 -16566
rect 25396 -16703 25604 -16697
rect 25396 -16737 25408 -16703
rect 25592 -16737 25604 -16703
rect 25396 -16743 25604 -16737
rect 25854 -16703 26062 -16697
rect 25854 -16737 25866 -16703
rect 26050 -16737 26062 -16703
rect 25854 -16743 26062 -16737
rect 25466 -16816 25526 -16743
rect 25926 -16816 25986 -16743
rect 25460 -16876 25466 -16816
rect 25526 -16876 25532 -16816
rect 25920 -16876 25926 -16816
rect 25986 -16876 25992 -16816
rect 26156 -17166 26216 -16644
rect 26622 -16644 26628 -15128
rect 26662 -15128 26674 -15068
rect 27080 -15068 27126 -15056
rect 26662 -16644 26668 -15128
rect 27080 -16572 27086 -15068
rect 26622 -16656 26668 -16644
rect 27064 -16644 27086 -16572
rect 27120 -16644 27126 -15068
rect 27530 -15068 27590 -14792
rect 27752 -14902 27758 -14842
rect 27818 -14902 27824 -14842
rect 28208 -14902 28214 -14842
rect 28274 -14902 28280 -14842
rect 28676 -14902 28682 -14842
rect 28742 -14902 28748 -14842
rect 29134 -14902 29140 -14842
rect 29200 -14902 29206 -14842
rect 27758 -14969 27818 -14902
rect 28214 -14969 28274 -14902
rect 28682 -14969 28742 -14902
rect 29140 -14969 29200 -14902
rect 27686 -14975 27894 -14969
rect 27686 -15009 27698 -14975
rect 27882 -15009 27894 -14975
rect 27686 -15015 27894 -15009
rect 28144 -14975 28352 -14969
rect 28144 -15009 28156 -14975
rect 28340 -15009 28352 -14975
rect 28144 -15015 28352 -15009
rect 28602 -14975 28810 -14969
rect 28602 -15009 28614 -14975
rect 28798 -15009 28810 -14975
rect 28602 -15015 28810 -15009
rect 29060 -14975 29268 -14969
rect 29060 -15009 29072 -14975
rect 29256 -15009 29268 -14975
rect 29060 -15015 29268 -15009
rect 27530 -15146 27544 -15068
rect 27064 -16656 27126 -16644
rect 27538 -16644 27544 -15146
rect 27578 -15146 27590 -15068
rect 27996 -15068 28042 -15056
rect 27578 -16644 27584 -15146
rect 27996 -16564 28002 -15068
rect 27538 -16656 27584 -16644
rect 27988 -16644 28002 -16564
rect 28036 -16564 28042 -15068
rect 28454 -15068 28500 -15056
rect 28036 -16644 28048 -16564
rect 28454 -16622 28460 -15068
rect 26312 -16703 26520 -16697
rect 26312 -16737 26324 -16703
rect 26508 -16737 26520 -16703
rect 26312 -16743 26520 -16737
rect 26770 -16703 26978 -16697
rect 26770 -16737 26782 -16703
rect 26966 -16737 26978 -16703
rect 26770 -16743 26978 -16737
rect 26382 -16816 26442 -16743
rect 26840 -16816 26900 -16743
rect 26376 -16876 26382 -16816
rect 26442 -16876 26448 -16816
rect 26834 -16876 26840 -16816
rect 26900 -16876 26906 -16816
rect 27064 -17040 27124 -16656
rect 27228 -16703 27436 -16697
rect 27228 -16737 27240 -16703
rect 27424 -16737 27436 -16703
rect 27228 -16743 27436 -16737
rect 27686 -16703 27894 -16697
rect 27686 -16737 27698 -16703
rect 27882 -16737 27894 -16703
rect 27686 -16743 27894 -16737
rect 27304 -16816 27364 -16743
rect 27758 -16816 27818 -16743
rect 27298 -16876 27304 -16816
rect 27364 -16876 27370 -16816
rect 27752 -16876 27758 -16816
rect 27818 -16876 27824 -16816
rect 27988 -16924 28048 -16644
rect 28450 -16644 28460 -16622
rect 28494 -16622 28500 -15068
rect 28912 -15068 28958 -15056
rect 28912 -16616 28918 -15068
rect 28494 -16644 28510 -16622
rect 28144 -16703 28352 -16697
rect 28144 -16737 28156 -16703
rect 28340 -16737 28352 -16703
rect 28144 -16743 28352 -16737
rect 28216 -16814 28276 -16743
rect 28450 -16804 28510 -16644
rect 28906 -16644 28918 -16616
rect 28952 -16616 28958 -15068
rect 29360 -15068 29420 -14792
rect 29590 -14902 29596 -14842
rect 29656 -14902 29662 -14842
rect 30046 -14902 30052 -14842
rect 30112 -14902 30118 -14842
rect 29596 -14969 29656 -14902
rect 30052 -14969 30112 -14902
rect 29518 -14975 29726 -14969
rect 29518 -15009 29530 -14975
rect 29714 -15009 29726 -14975
rect 29518 -15015 29726 -15009
rect 29976 -14975 30184 -14969
rect 29976 -15009 29988 -14975
rect 30172 -15009 30184 -14975
rect 29976 -15015 30184 -15009
rect 29360 -15112 29376 -15068
rect 28952 -16644 28966 -16616
rect 28602 -16703 28810 -16697
rect 28602 -16737 28614 -16703
rect 28798 -16737 28810 -16703
rect 28602 -16743 28810 -16737
rect 28210 -16816 28282 -16814
rect 28210 -16876 28216 -16816
rect 28276 -16876 28282 -16816
rect 28676 -16808 28736 -16743
rect 28450 -16870 28510 -16864
rect 28664 -16814 28748 -16808
rect 28664 -16876 28676 -16814
rect 28736 -16876 28748 -16814
rect 28664 -16880 28748 -16876
rect 28906 -16924 28966 -16644
rect 29370 -16644 29376 -15112
rect 29410 -15112 29420 -15068
rect 29828 -15068 29874 -15056
rect 29410 -16644 29416 -15112
rect 29828 -16612 29834 -15068
rect 29370 -16656 29416 -16644
rect 29820 -16644 29834 -16612
rect 29868 -16612 29874 -15068
rect 30276 -15068 30336 -14668
rect 30502 -14902 30508 -14842
rect 30568 -14902 30574 -14842
rect 30958 -14902 30964 -14842
rect 31024 -14902 31030 -14842
rect 30508 -14969 30568 -14902
rect 30964 -14969 31024 -14902
rect 30434 -14975 30642 -14969
rect 30434 -15009 30446 -14975
rect 30630 -15009 30642 -14975
rect 30434 -15015 30642 -15009
rect 30892 -14975 31100 -14969
rect 30892 -15009 30904 -14975
rect 31088 -15009 31100 -14975
rect 30892 -15015 31100 -15009
rect 30276 -15126 30292 -15068
rect 29868 -16644 29880 -16612
rect 29060 -16703 29268 -16697
rect 29060 -16737 29072 -16703
rect 29256 -16737 29268 -16703
rect 29060 -16743 29268 -16737
rect 29518 -16703 29726 -16697
rect 29518 -16737 29530 -16703
rect 29714 -16737 29726 -16703
rect 29518 -16743 29726 -16737
rect 29132 -16816 29192 -16743
rect 29592 -16816 29652 -16743
rect 29126 -16876 29132 -16816
rect 29192 -16876 29198 -16816
rect 29586 -16876 29592 -16816
rect 29652 -16876 29658 -16816
rect 27988 -16984 28966 -16924
rect 29820 -17040 29880 -16644
rect 30286 -16644 30292 -15126
rect 30326 -15126 30336 -15068
rect 30744 -15068 30790 -15056
rect 30326 -16644 30332 -15126
rect 30744 -16576 30750 -15068
rect 30286 -16656 30332 -16644
rect 30740 -16644 30750 -16576
rect 30784 -16576 30790 -15068
rect 31196 -15068 31256 -14534
rect 31416 -14902 31422 -14842
rect 31482 -14902 31488 -14842
rect 31876 -14902 31882 -14842
rect 31942 -14902 31948 -14842
rect 31422 -14969 31482 -14902
rect 31882 -14969 31942 -14902
rect 31350 -14975 31558 -14969
rect 31350 -15009 31362 -14975
rect 31546 -15009 31558 -14975
rect 31350 -15015 31558 -15009
rect 31808 -14975 32016 -14969
rect 31808 -15009 31820 -14975
rect 32004 -15009 32016 -14975
rect 31808 -15015 32016 -15009
rect 31196 -15124 31208 -15068
rect 30784 -16644 30800 -16576
rect 29976 -16703 30184 -16697
rect 29976 -16737 29988 -16703
rect 30172 -16737 30184 -16703
rect 29976 -16743 30184 -16737
rect 30434 -16703 30642 -16697
rect 30434 -16737 30446 -16703
rect 30630 -16737 30642 -16703
rect 30434 -16743 30642 -16737
rect 30048 -16816 30108 -16743
rect 30504 -16816 30564 -16743
rect 30042 -16876 30048 -16816
rect 30108 -16876 30114 -16816
rect 30498 -16876 30504 -16816
rect 30564 -16876 30570 -16816
rect 27064 -17100 29880 -17040
rect 30740 -17166 30800 -16644
rect 31202 -16644 31208 -15124
rect 31242 -15124 31256 -15068
rect 31660 -15068 31706 -15056
rect 31242 -16644 31248 -15124
rect 31660 -16584 31666 -15068
rect 31202 -16656 31248 -16644
rect 31654 -16644 31666 -16584
rect 31700 -16584 31706 -15068
rect 32112 -15068 32172 -14280
rect 32342 -14969 32402 -14280
rect 32266 -14975 32474 -14969
rect 32266 -15009 32278 -14975
rect 32462 -15009 32474 -14975
rect 32266 -15015 32474 -15009
rect 32112 -15144 32124 -15068
rect 32118 -16582 32124 -15144
rect 31700 -16644 31714 -16584
rect 30892 -16703 31100 -16697
rect 30892 -16737 30904 -16703
rect 31088 -16737 31100 -16703
rect 30892 -16743 31100 -16737
rect 31350 -16703 31558 -16697
rect 31350 -16737 31362 -16703
rect 31546 -16737 31558 -16703
rect 31350 -16743 31558 -16737
rect 30960 -16816 31020 -16743
rect 31418 -16816 31478 -16743
rect 30954 -16876 30960 -16816
rect 31020 -16876 31026 -16816
rect 31412 -16876 31418 -16816
rect 31478 -16876 31484 -16816
rect 26156 -17226 30800 -17166
rect 31654 -17296 31714 -16644
rect 32108 -16644 32124 -16582
rect 32158 -15144 32172 -15068
rect 32570 -15068 32630 -14280
rect 32570 -15138 32582 -15068
rect 32158 -16582 32164 -15144
rect 32158 -16644 32168 -16582
rect 32576 -16600 32582 -15138
rect 31808 -16703 32016 -16697
rect 31808 -16737 31820 -16703
rect 32004 -16737 32016 -16703
rect 31808 -16743 32016 -16737
rect 31878 -16816 31938 -16743
rect 31872 -16876 31878 -16816
rect 31938 -16876 31944 -16816
rect 32108 -16818 32168 -16644
rect 32566 -16644 32582 -16600
rect 32616 -15138 32630 -15068
rect 32616 -16600 32622 -15138
rect 32616 -16644 32626 -16600
rect 32266 -16703 32474 -16697
rect 32266 -16737 32278 -16703
rect 32462 -16737 32474 -16703
rect 32266 -16743 32474 -16737
rect 32340 -16818 32400 -16743
rect 32566 -16818 32626 -16644
rect 33690 -16818 33696 -13994
rect 32108 -16878 33696 -16818
rect 23452 -19166 23458 -17308
rect 23766 -17733 23826 -17308
rect 23994 -17634 24054 -17308
rect 25238 -17356 31714 -17296
rect 32566 -17312 32626 -16878
rect 33690 -17312 33696 -16878
rect 32566 -17372 33696 -17312
rect 24218 -17462 24224 -17402
rect 24284 -17462 24290 -17402
rect 23921 -17640 24129 -17634
rect 23921 -17674 23933 -17640
rect 24117 -17674 24129 -17640
rect 23921 -17680 24129 -17674
rect 23766 -17780 23779 -17733
rect 23773 -18888 23779 -17780
rect 23346 -19342 23458 -19166
rect 23766 -18909 23779 -18888
rect 23813 -17780 23826 -17733
rect 24224 -17733 24284 -17462
rect 24456 -17564 27720 -17504
rect 24456 -17634 24516 -17564
rect 24918 -17634 24978 -17564
rect 25372 -17634 25432 -17564
rect 25834 -17634 25894 -17564
rect 26288 -17634 26348 -17564
rect 26738 -17634 26798 -17564
rect 27204 -17634 27264 -17564
rect 27660 -17634 27720 -17564
rect 28116 -17582 29284 -17522
rect 28116 -17634 28176 -17582
rect 24379 -17640 24587 -17634
rect 24379 -17674 24391 -17640
rect 24575 -17674 24587 -17640
rect 24379 -17680 24587 -17674
rect 24837 -17640 25045 -17634
rect 24837 -17674 24849 -17640
rect 25033 -17674 25045 -17640
rect 24837 -17680 25045 -17674
rect 25295 -17640 25503 -17634
rect 25295 -17674 25307 -17640
rect 25491 -17674 25503 -17640
rect 25295 -17680 25503 -17674
rect 25753 -17640 25961 -17634
rect 25753 -17674 25765 -17640
rect 25949 -17674 25961 -17640
rect 25753 -17680 25961 -17674
rect 26211 -17640 26419 -17634
rect 26211 -17674 26223 -17640
rect 26407 -17674 26419 -17640
rect 26211 -17680 26419 -17674
rect 26669 -17640 26877 -17634
rect 26669 -17674 26681 -17640
rect 26865 -17674 26877 -17640
rect 26669 -17680 26877 -17674
rect 27127 -17640 27335 -17634
rect 27127 -17674 27139 -17640
rect 27323 -17674 27335 -17640
rect 27127 -17680 27335 -17674
rect 27585 -17640 27793 -17634
rect 27585 -17674 27597 -17640
rect 27781 -17674 27793 -17640
rect 27585 -17680 27793 -17674
rect 28043 -17640 28251 -17634
rect 28043 -17674 28055 -17640
rect 28239 -17674 28251 -17640
rect 28043 -17680 28251 -17674
rect 23813 -18888 23819 -17780
rect 24224 -17800 24237 -17733
rect 23813 -18909 23826 -18888
rect 23766 -19342 23826 -18909
rect 24231 -18909 24237 -17800
rect 24271 -17800 24284 -17733
rect 24689 -17733 24735 -17721
rect 24271 -18909 24277 -17800
rect 24231 -18921 24277 -18909
rect 24689 -18909 24695 -17733
rect 24729 -18909 24735 -17733
rect 24689 -18921 24735 -18909
rect 25147 -17733 25193 -17721
rect 25147 -18909 25153 -17733
rect 25187 -18909 25193 -17733
rect 25147 -18921 25193 -18909
rect 25605 -17733 25651 -17721
rect 25605 -18909 25611 -17733
rect 25645 -18909 25651 -17733
rect 25605 -18921 25651 -18909
rect 26063 -17733 26109 -17721
rect 26063 -18909 26069 -17733
rect 26103 -18909 26109 -17733
rect 26063 -18921 26109 -18909
rect 26521 -17733 26567 -17721
rect 26521 -18909 26527 -17733
rect 26561 -18909 26567 -17733
rect 26521 -18921 26567 -18909
rect 26979 -17733 27025 -17721
rect 26979 -18909 26985 -17733
rect 27019 -18909 27025 -17733
rect 26979 -18921 27025 -18909
rect 27437 -17733 27483 -17721
rect 27437 -18909 27443 -17733
rect 27477 -18909 27483 -17733
rect 27895 -17733 27941 -17721
rect 27895 -18842 27901 -17733
rect 27437 -18921 27483 -18909
rect 27886 -18909 27901 -18842
rect 27935 -18842 27941 -17733
rect 28346 -17733 28406 -17582
rect 28346 -17748 28359 -17733
rect 27935 -18909 27946 -18842
rect 28353 -18874 28359 -17748
rect 23921 -18968 24129 -18962
rect 23921 -19002 23933 -18968
rect 24117 -19002 24129 -18968
rect 23921 -19008 24129 -19002
rect 24379 -18968 24587 -18962
rect 24379 -19002 24391 -18968
rect 24575 -19002 24587 -18968
rect 24379 -19008 24587 -19002
rect 24837 -18968 25045 -18962
rect 24837 -19002 24849 -18968
rect 25033 -19002 25045 -18968
rect 24837 -19008 25045 -19002
rect 25295 -18968 25503 -18962
rect 25295 -19002 25307 -18968
rect 25491 -19002 25503 -18968
rect 25295 -19008 25503 -19002
rect 25753 -18968 25961 -18962
rect 25753 -19002 25765 -18968
rect 25949 -19002 25961 -18968
rect 25753 -19008 25961 -19002
rect 26211 -18968 26419 -18962
rect 26211 -19002 26223 -18968
rect 26407 -19002 26419 -18968
rect 26211 -19008 26419 -19002
rect 26669 -18968 26877 -18962
rect 26669 -19002 26681 -18968
rect 26865 -19002 26877 -18968
rect 26669 -19008 26877 -19002
rect 27127 -18968 27335 -18962
rect 27127 -19002 27139 -18968
rect 27323 -19002 27335 -18968
rect 27127 -19008 27335 -19002
rect 27585 -18968 27793 -18962
rect 27585 -19002 27597 -18968
rect 27781 -19002 27793 -18968
rect 27585 -19008 27793 -19002
rect 23994 -19342 24054 -19008
rect 24448 -19076 24508 -19008
rect 24910 -19076 24970 -19008
rect 25364 -19076 25424 -19008
rect 25826 -19076 25886 -19008
rect 26280 -19076 26340 -19008
rect 26730 -19076 26790 -19008
rect 27196 -19076 27256 -19008
rect 27652 -19076 27712 -19008
rect 24448 -19080 25364 -19076
rect 24508 -19136 24910 -19080
rect 24448 -19146 24508 -19140
rect 24970 -19136 25364 -19080
rect 25424 -19136 25826 -19076
rect 25886 -19082 26730 -19076
rect 25886 -19136 26280 -19082
rect 24910 -19146 24970 -19140
rect 25364 -19142 25424 -19136
rect 25826 -19142 25886 -19136
rect 26340 -19136 26730 -19082
rect 26790 -19136 27196 -19076
rect 27256 -19080 27712 -19076
rect 27256 -19136 27652 -19080
rect 26730 -19142 26790 -19136
rect 27196 -19142 27256 -19136
rect 26280 -19148 26340 -19142
rect 27652 -19146 27712 -19140
rect 27886 -19202 27946 -18909
rect 28344 -18909 28359 -18874
rect 28393 -17748 28406 -17733
rect 28766 -17733 28826 -17582
rect 28998 -17634 29058 -17582
rect 28921 -17640 29129 -17634
rect 28921 -17674 28933 -17640
rect 29117 -17674 29129 -17640
rect 28921 -17680 29129 -17674
rect 28393 -18874 28399 -17748
rect 28766 -17754 28779 -17733
rect 28773 -18874 28779 -17754
rect 28393 -18909 28404 -18874
rect 28043 -18968 28251 -18962
rect 28043 -19002 28055 -18968
rect 28239 -19002 28251 -18968
rect 28043 -19008 28251 -19002
rect 27880 -19262 27886 -19202
rect 27946 -19262 27952 -19202
rect 28116 -19342 28176 -19008
rect 28344 -19342 28404 -18909
rect 28764 -18909 28779 -18874
rect 28813 -17754 28826 -17733
rect 29224 -17733 29284 -17582
rect 29450 -17564 32714 -17504
rect 29450 -17634 29510 -17564
rect 29912 -17634 29972 -17564
rect 30366 -17634 30426 -17564
rect 30828 -17634 30888 -17564
rect 31282 -17634 31342 -17564
rect 31732 -17634 31792 -17564
rect 32198 -17634 32258 -17564
rect 32654 -17634 32714 -17564
rect 33116 -17634 33176 -17372
rect 29379 -17640 29587 -17634
rect 29379 -17674 29391 -17640
rect 29575 -17674 29587 -17640
rect 29379 -17680 29587 -17674
rect 29837 -17640 30045 -17634
rect 29837 -17674 29849 -17640
rect 30033 -17674 30045 -17640
rect 29837 -17680 30045 -17674
rect 30295 -17640 30503 -17634
rect 30295 -17674 30307 -17640
rect 30491 -17674 30503 -17640
rect 30295 -17680 30503 -17674
rect 30753 -17640 30961 -17634
rect 30753 -17674 30765 -17640
rect 30949 -17674 30961 -17640
rect 30753 -17680 30961 -17674
rect 31211 -17640 31419 -17634
rect 31211 -17674 31223 -17640
rect 31407 -17674 31419 -17640
rect 31211 -17680 31419 -17674
rect 31669 -17640 31877 -17634
rect 31669 -17674 31681 -17640
rect 31865 -17674 31877 -17640
rect 31669 -17680 31877 -17674
rect 32127 -17640 32335 -17634
rect 32127 -17674 32139 -17640
rect 32323 -17674 32335 -17640
rect 32127 -17680 32335 -17674
rect 32585 -17640 32793 -17634
rect 32585 -17674 32597 -17640
rect 32781 -17674 32793 -17640
rect 32585 -17680 32793 -17674
rect 33043 -17640 33251 -17634
rect 33043 -17674 33055 -17640
rect 33239 -17674 33251 -17640
rect 33043 -17680 33251 -17674
rect 28813 -18874 28819 -17754
rect 29224 -17776 29237 -17733
rect 29231 -18868 29237 -17776
rect 28813 -18909 28824 -18874
rect 28764 -19342 28824 -18909
rect 29222 -18909 29237 -18868
rect 29271 -17776 29284 -17733
rect 29689 -17733 29735 -17721
rect 29271 -18868 29277 -17776
rect 29271 -18909 29282 -18868
rect 28921 -18968 29129 -18962
rect 28921 -19002 28933 -18968
rect 29117 -19002 29129 -18968
rect 28921 -19008 29129 -19002
rect 28992 -19342 29052 -19008
rect 29222 -19342 29282 -18909
rect 29689 -18909 29695 -17733
rect 29729 -18909 29735 -17733
rect 29689 -18921 29735 -18909
rect 30147 -17733 30193 -17721
rect 30147 -18909 30153 -17733
rect 30187 -18909 30193 -17733
rect 30147 -18921 30193 -18909
rect 30605 -17733 30651 -17721
rect 30605 -18909 30611 -17733
rect 30645 -18909 30651 -17733
rect 30605 -18921 30651 -18909
rect 31063 -17733 31109 -17721
rect 31063 -18909 31069 -17733
rect 31103 -18909 31109 -17733
rect 31063 -18921 31109 -18909
rect 31521 -17733 31567 -17721
rect 31521 -18909 31527 -17733
rect 31561 -18909 31567 -17733
rect 31521 -18921 31567 -18909
rect 31979 -17733 32025 -17721
rect 31979 -18909 31985 -17733
rect 32019 -18909 32025 -17733
rect 31979 -18921 32025 -18909
rect 32437 -17733 32483 -17721
rect 32437 -18909 32443 -17733
rect 32477 -18909 32483 -17733
rect 32895 -17733 32941 -17721
rect 32895 -18902 32901 -17733
rect 32437 -18921 32483 -18909
rect 32886 -18909 32901 -18902
rect 32935 -18902 32941 -17733
rect 33342 -17733 33402 -17372
rect 33342 -17786 33359 -17733
rect 33353 -18876 33359 -17786
rect 32935 -18909 32946 -18902
rect 29379 -18968 29587 -18962
rect 29379 -19002 29391 -18968
rect 29575 -19002 29587 -18968
rect 29379 -19008 29587 -19002
rect 29837 -18968 30045 -18962
rect 29837 -19002 29849 -18968
rect 30033 -19002 30045 -18968
rect 29837 -19008 30045 -19002
rect 30295 -18968 30503 -18962
rect 30295 -19002 30307 -18968
rect 30491 -19002 30503 -18968
rect 30295 -19008 30503 -19002
rect 30753 -18968 30961 -18962
rect 30753 -19002 30765 -18968
rect 30949 -19002 30961 -18968
rect 30753 -19008 30961 -19002
rect 31211 -18968 31419 -18962
rect 31211 -19002 31223 -18968
rect 31407 -19002 31419 -18968
rect 31211 -19008 31419 -19002
rect 31669 -18968 31877 -18962
rect 31669 -19002 31681 -18968
rect 31865 -19002 31877 -18968
rect 31669 -19008 31877 -19002
rect 32127 -18968 32335 -18962
rect 32127 -19002 32139 -18968
rect 32323 -19002 32335 -18968
rect 32127 -19008 32335 -19002
rect 32585 -18968 32793 -18962
rect 32585 -19002 32597 -18968
rect 32781 -19002 32793 -18968
rect 32585 -19008 32793 -19002
rect 29450 -19076 29510 -19008
rect 29912 -19072 29972 -19008
rect 29450 -19080 29912 -19076
rect 29510 -19132 29912 -19080
rect 30366 -19076 30426 -19008
rect 30828 -19076 30888 -19008
rect 31282 -19076 31342 -19008
rect 31732 -19072 31792 -19008
rect 29972 -19078 31732 -19076
rect 29972 -19132 30366 -19078
rect 29510 -19136 30366 -19132
rect 29912 -19138 29972 -19136
rect 30426 -19136 30828 -19078
rect 29450 -19146 29510 -19140
rect 30366 -19144 30426 -19138
rect 30888 -19136 31282 -19078
rect 30828 -19144 30888 -19138
rect 31342 -19132 31732 -19078
rect 32198 -19076 32258 -19008
rect 32654 -19076 32714 -19008
rect 31792 -19078 32714 -19076
rect 31792 -19132 32198 -19078
rect 31342 -19136 32198 -19132
rect 31732 -19138 31792 -19136
rect 32258 -19136 32654 -19078
rect 31282 -19144 31342 -19138
rect 32198 -19144 32258 -19138
rect 32654 -19144 32714 -19138
rect 32886 -19208 32946 -18909
rect 33344 -18909 33359 -18876
rect 33393 -17786 33402 -17733
rect 33393 -18876 33399 -17786
rect 33393 -18909 33404 -18876
rect 33043 -18968 33251 -18962
rect 33043 -19002 33055 -18968
rect 33239 -19002 33251 -18968
rect 33043 -19008 33251 -19002
rect 32886 -19274 32946 -19268
rect 33116 -19342 33176 -19008
rect 33344 -19342 33404 -18909
rect 33690 -19166 33696 -17372
rect 33796 -19166 33802 -13994
rect 33690 -19342 33802 -19166
rect 23346 -19348 33802 -19342
rect 23346 -19448 23452 -19348
rect 33696 -19448 33802 -19348
rect 23346 -19454 33802 -19448
rect 23346 -19684 33802 -19678
rect 23346 -19784 23452 -19684
rect 33696 -19784 33802 -19684
rect 23346 -19790 33802 -19784
rect 23346 -19914 23458 -19790
rect 23074 -21286 23080 -21226
rect 23140 -21286 23146 -21226
rect 18690 -22042 18802 -21918
rect 8346 -22048 18802 -22042
rect 8346 -22148 8452 -22048
rect 18696 -22148 18802 -22048
rect 8346 -22154 18802 -22148
rect 23346 -21918 23352 -19914
rect 23452 -21918 23458 -19914
rect 23766 -20226 23826 -19790
rect 23996 -20136 24056 -19790
rect 27886 -19882 27946 -19876
rect 24454 -20016 24910 -20010
rect 24442 -20076 24448 -20016
rect 24508 -20070 24910 -20016
rect 24970 -20016 25826 -20010
rect 24970 -20070 25364 -20016
rect 24508 -20076 24514 -20070
rect 24448 -20136 24514 -20076
rect 24910 -20136 24976 -20070
rect 25358 -20076 25364 -20070
rect 25424 -20070 25826 -20016
rect 25886 -20070 26280 -20010
rect 26340 -20070 26730 -20010
rect 26790 -20016 27652 -20010
rect 26790 -20070 27196 -20016
rect 25424 -20076 25430 -20070
rect 25364 -20136 25430 -20076
rect 25826 -20136 25892 -20070
rect 26280 -20136 26346 -20070
rect 26730 -20136 26796 -20070
rect 27190 -20076 27196 -20070
rect 27256 -20070 27652 -20016
rect 27712 -20070 27718 -20010
rect 27256 -20076 27262 -20070
rect 27196 -20136 27262 -20076
rect 27652 -20136 27718 -20070
rect 23920 -20142 24128 -20136
rect 23920 -20176 23932 -20142
rect 24116 -20176 24128 -20142
rect 23920 -20182 24128 -20176
rect 24378 -20142 24586 -20136
rect 24378 -20176 24390 -20142
rect 24574 -20176 24586 -20142
rect 24378 -20182 24586 -20176
rect 24836 -20142 25044 -20136
rect 24836 -20176 24848 -20142
rect 25032 -20176 25044 -20142
rect 24836 -20182 25044 -20176
rect 25294 -20142 25502 -20136
rect 25294 -20176 25306 -20142
rect 25490 -20176 25502 -20142
rect 25294 -20182 25502 -20176
rect 25752 -20142 25960 -20136
rect 25752 -20176 25764 -20142
rect 25948 -20176 25960 -20142
rect 25752 -20182 25960 -20176
rect 26210 -20142 26418 -20136
rect 26210 -20176 26222 -20142
rect 26406 -20176 26418 -20142
rect 26210 -20182 26418 -20176
rect 26668 -20142 26876 -20136
rect 26668 -20176 26680 -20142
rect 26864 -20176 26876 -20142
rect 26668 -20182 26876 -20176
rect 27126 -20142 27334 -20136
rect 27126 -20176 27138 -20142
rect 27322 -20176 27334 -20142
rect 27126 -20182 27334 -20176
rect 27584 -20142 27792 -20136
rect 27584 -20176 27596 -20142
rect 27780 -20176 27792 -20142
rect 27584 -20182 27792 -20176
rect 23766 -20266 23778 -20226
rect 23772 -20362 23778 -20266
rect 23766 -20402 23778 -20362
rect 23812 -20266 23826 -20226
rect 24230 -20226 24276 -20214
rect 23812 -20362 23818 -20266
rect 24230 -20360 24236 -20226
rect 23812 -20402 23826 -20362
rect 23766 -20618 23826 -20402
rect 24222 -20402 24236 -20360
rect 24270 -20360 24276 -20226
rect 24688 -20226 24734 -20214
rect 24270 -20402 24282 -20360
rect 23920 -20452 24128 -20446
rect 23920 -20486 23932 -20452
rect 24116 -20486 24128 -20452
rect 23920 -20492 24128 -20486
rect 23994 -20618 24054 -20492
rect 23766 -20678 24054 -20618
rect 23766 -20894 23826 -20678
rect 23994 -20804 24054 -20678
rect 23920 -20810 24128 -20804
rect 23920 -20844 23932 -20810
rect 24116 -20844 24128 -20810
rect 23920 -20850 24128 -20844
rect 23766 -20914 23778 -20894
rect 23772 -21040 23778 -20914
rect 23758 -21070 23778 -21040
rect 23812 -20914 23826 -20894
rect 24222 -20894 24282 -20402
rect 24688 -20402 24694 -20226
rect 24728 -20402 24734 -20226
rect 24688 -20414 24734 -20402
rect 25146 -20226 25192 -20214
rect 25146 -20402 25152 -20226
rect 25186 -20402 25192 -20226
rect 25146 -20414 25192 -20402
rect 25604 -20226 25650 -20214
rect 25604 -20402 25610 -20226
rect 25644 -20402 25650 -20226
rect 25604 -20414 25650 -20402
rect 26062 -20226 26108 -20214
rect 26062 -20402 26068 -20226
rect 26102 -20402 26108 -20226
rect 26062 -20414 26108 -20402
rect 26520 -20226 26566 -20214
rect 26520 -20402 26526 -20226
rect 26560 -20402 26566 -20226
rect 26520 -20414 26566 -20402
rect 26978 -20226 27024 -20214
rect 26978 -20402 26984 -20226
rect 27018 -20402 27024 -20226
rect 26978 -20414 27024 -20402
rect 27436 -20226 27482 -20214
rect 27436 -20402 27442 -20226
rect 27476 -20402 27482 -20226
rect 27886 -20226 27946 -19942
rect 28114 -20136 28174 -19790
rect 28042 -20142 28250 -20136
rect 28042 -20176 28054 -20142
rect 28238 -20176 28250 -20142
rect 28042 -20182 28250 -20176
rect 27886 -20256 27900 -20226
rect 27436 -20414 27482 -20402
rect 27894 -20402 27900 -20256
rect 27934 -20256 27946 -20226
rect 28346 -20226 28406 -19790
rect 28346 -20254 28358 -20226
rect 27934 -20402 27940 -20256
rect 28352 -20346 28358 -20254
rect 27894 -20414 27940 -20402
rect 28346 -20402 28358 -20346
rect 28392 -20254 28406 -20226
rect 28766 -20226 28826 -19790
rect 29000 -20136 29060 -19790
rect 28920 -20142 29128 -20136
rect 28920 -20176 28932 -20142
rect 29116 -20176 29128 -20142
rect 28920 -20182 29128 -20176
rect 28392 -20346 28398 -20254
rect 28766 -20262 28778 -20226
rect 28392 -20402 28406 -20346
rect 28772 -20366 28778 -20262
rect 24378 -20452 24586 -20446
rect 24378 -20486 24390 -20452
rect 24574 -20486 24586 -20452
rect 24378 -20492 24586 -20486
rect 24836 -20452 25044 -20446
rect 24836 -20486 24848 -20452
rect 25032 -20486 25044 -20452
rect 24836 -20492 25044 -20486
rect 25294 -20452 25502 -20446
rect 25294 -20486 25306 -20452
rect 25490 -20486 25502 -20452
rect 25294 -20492 25502 -20486
rect 25752 -20452 25960 -20446
rect 25752 -20486 25764 -20452
rect 25948 -20486 25960 -20452
rect 25752 -20492 25960 -20486
rect 26210 -20452 26418 -20446
rect 26210 -20486 26222 -20452
rect 26406 -20486 26418 -20452
rect 26210 -20492 26418 -20486
rect 26668 -20452 26876 -20446
rect 26668 -20486 26680 -20452
rect 26864 -20486 26876 -20452
rect 26668 -20492 26876 -20486
rect 27126 -20452 27334 -20446
rect 27126 -20486 27138 -20452
rect 27322 -20486 27334 -20452
rect 27126 -20492 27334 -20486
rect 27584 -20452 27792 -20446
rect 27584 -20486 27596 -20452
rect 27780 -20486 27792 -20452
rect 27584 -20492 27792 -20486
rect 28042 -20452 28250 -20446
rect 28042 -20486 28054 -20452
rect 28238 -20486 28250 -20452
rect 28042 -20492 28250 -20486
rect 24448 -20558 24508 -20492
rect 24910 -20558 24970 -20492
rect 25364 -20558 25424 -20492
rect 25826 -20558 25886 -20492
rect 26280 -20558 26340 -20492
rect 26730 -20558 26790 -20492
rect 27196 -20558 27256 -20492
rect 27652 -20558 27712 -20492
rect 24448 -20618 27712 -20558
rect 24454 -20738 27718 -20678
rect 24454 -20804 24514 -20738
rect 24916 -20804 24976 -20738
rect 25370 -20804 25430 -20738
rect 25832 -20804 25892 -20738
rect 26286 -20804 26346 -20738
rect 26736 -20804 26796 -20738
rect 27202 -20804 27262 -20738
rect 27658 -20804 27718 -20738
rect 28114 -20804 28174 -20492
rect 24378 -20810 24586 -20804
rect 24378 -20844 24390 -20810
rect 24574 -20844 24586 -20810
rect 24378 -20850 24586 -20844
rect 24836 -20810 25044 -20804
rect 24836 -20844 24848 -20810
rect 25032 -20844 25044 -20810
rect 24836 -20850 25044 -20844
rect 25294 -20810 25502 -20804
rect 25294 -20844 25306 -20810
rect 25490 -20844 25502 -20810
rect 25294 -20850 25502 -20844
rect 25752 -20810 25960 -20804
rect 25752 -20844 25764 -20810
rect 25948 -20844 25960 -20810
rect 25752 -20850 25960 -20844
rect 26210 -20810 26418 -20804
rect 26210 -20844 26222 -20810
rect 26406 -20844 26418 -20810
rect 26210 -20850 26418 -20844
rect 26668 -20810 26876 -20804
rect 26668 -20844 26680 -20810
rect 26864 -20844 26876 -20810
rect 26668 -20850 26876 -20844
rect 27126 -20810 27334 -20804
rect 27126 -20844 27138 -20810
rect 27322 -20844 27334 -20810
rect 27126 -20850 27334 -20844
rect 27584 -20810 27792 -20804
rect 27584 -20844 27596 -20810
rect 27780 -20844 27792 -20810
rect 27584 -20850 27792 -20844
rect 28042 -20810 28250 -20804
rect 28042 -20844 28054 -20810
rect 28238 -20844 28250 -20810
rect 28042 -20850 28250 -20844
rect 23812 -21070 23818 -20914
rect 24222 -20922 24236 -20894
rect 23758 -21450 23818 -21070
rect 24230 -21070 24236 -20922
rect 24270 -20922 24282 -20894
rect 24688 -20894 24734 -20882
rect 24270 -21070 24276 -20922
rect 24230 -21082 24276 -21070
rect 24688 -21070 24694 -20894
rect 24728 -21070 24734 -20894
rect 24688 -21082 24734 -21070
rect 25146 -20894 25192 -20882
rect 25146 -21070 25152 -20894
rect 25186 -21070 25192 -20894
rect 25146 -21082 25192 -21070
rect 25604 -20894 25650 -20882
rect 25604 -21070 25610 -20894
rect 25644 -21070 25650 -20894
rect 25604 -21082 25650 -21070
rect 26062 -20894 26108 -20882
rect 26062 -21070 26068 -20894
rect 26102 -21070 26108 -20894
rect 26062 -21082 26108 -21070
rect 26520 -20894 26566 -20882
rect 26520 -21070 26526 -20894
rect 26560 -21070 26566 -20894
rect 26520 -21082 26566 -21070
rect 26978 -20894 27024 -20882
rect 26978 -21070 26984 -20894
rect 27018 -21070 27024 -20894
rect 26978 -21082 27024 -21070
rect 27436 -20894 27482 -20882
rect 27436 -21070 27442 -20894
rect 27476 -21070 27482 -20894
rect 27894 -20894 27940 -20882
rect 27894 -21042 27900 -20894
rect 27436 -21082 27482 -21070
rect 27886 -21070 27900 -21042
rect 27934 -21042 27940 -20894
rect 28346 -20894 28406 -20402
rect 27934 -21070 27946 -21042
rect 23920 -21120 24128 -21114
rect 23920 -21154 23932 -21120
rect 24116 -21154 24128 -21120
rect 23920 -21160 24128 -21154
rect 24378 -21120 24586 -21114
rect 24378 -21154 24390 -21120
rect 24574 -21154 24586 -21120
rect 24378 -21160 24586 -21154
rect 24836 -21120 25044 -21114
rect 24836 -21154 24848 -21120
rect 25032 -21154 25044 -21120
rect 24836 -21160 25044 -21154
rect 25294 -21120 25502 -21114
rect 25294 -21154 25306 -21120
rect 25490 -21154 25502 -21120
rect 25294 -21160 25502 -21154
rect 25752 -21120 25960 -21114
rect 25752 -21154 25764 -21120
rect 25948 -21154 25960 -21120
rect 25752 -21160 25960 -21154
rect 26210 -21120 26418 -21114
rect 26210 -21154 26222 -21120
rect 26406 -21154 26418 -21120
rect 26210 -21160 26418 -21154
rect 26668 -21120 26876 -21114
rect 26668 -21154 26680 -21120
rect 26864 -21154 26876 -21120
rect 26668 -21160 26876 -21154
rect 27126 -21120 27334 -21114
rect 27126 -21154 27138 -21120
rect 27322 -21154 27334 -21120
rect 27126 -21160 27334 -21154
rect 27584 -21120 27792 -21114
rect 27584 -21154 27596 -21120
rect 27780 -21154 27792 -21120
rect 27584 -21160 27792 -21154
rect 23998 -21450 24058 -21160
rect 24448 -21226 24508 -21160
rect 24910 -21226 24970 -21160
rect 25364 -21226 25424 -21160
rect 25826 -21226 25886 -21160
rect 26280 -21226 26340 -21160
rect 26730 -21226 26790 -21160
rect 27196 -21226 27256 -21160
rect 27652 -21226 27712 -21160
rect 24442 -21286 24448 -21226
rect 24508 -21286 27712 -21226
rect 27886 -21450 27946 -21070
rect 28346 -21070 28358 -20894
rect 28392 -21070 28406 -20894
rect 28042 -21120 28250 -21114
rect 28042 -21154 28054 -21120
rect 28238 -21154 28250 -21120
rect 28042 -21160 28250 -21154
rect 28112 -21450 28172 -21160
rect 28346 -21450 28406 -21070
rect 28762 -20402 28778 -20366
rect 28812 -20262 28826 -20226
rect 29222 -20226 29282 -19790
rect 32880 -19930 32886 -19870
rect 32946 -19930 32952 -19870
rect 31726 -20010 31732 -20006
rect 29444 -20070 29450 -20010
rect 29510 -20012 31732 -20010
rect 29510 -20070 29912 -20012
rect 29450 -20136 29514 -20070
rect 29906 -20072 29912 -20070
rect 29972 -20070 30366 -20012
rect 29972 -20072 29978 -20070
rect 30360 -20072 30366 -20070
rect 30426 -20070 30828 -20012
rect 30426 -20072 30432 -20070
rect 30822 -20072 30828 -20070
rect 30888 -20070 31282 -20012
rect 30888 -20072 30894 -20070
rect 31276 -20072 31282 -20070
rect 31342 -20066 31732 -20012
rect 31792 -20010 31798 -20006
rect 31792 -20066 32198 -20010
rect 31342 -20070 32198 -20066
rect 32258 -20070 32654 -20010
rect 32714 -20070 32720 -20010
rect 31342 -20072 31348 -20070
rect 29912 -20136 29976 -20072
rect 30366 -20136 30430 -20072
rect 30828 -20136 30892 -20072
rect 31282 -20136 31346 -20072
rect 31732 -20136 31796 -20070
rect 32198 -20136 32262 -20070
rect 32654 -20136 32718 -20070
rect 29378 -20142 29586 -20136
rect 29378 -20176 29390 -20142
rect 29574 -20176 29586 -20142
rect 29378 -20182 29586 -20176
rect 29836 -20142 30044 -20136
rect 29836 -20176 29848 -20142
rect 30032 -20176 30044 -20142
rect 29836 -20182 30044 -20176
rect 30294 -20142 30502 -20136
rect 30294 -20176 30306 -20142
rect 30490 -20176 30502 -20142
rect 30294 -20182 30502 -20176
rect 30752 -20142 30960 -20136
rect 30752 -20176 30764 -20142
rect 30948 -20176 30960 -20142
rect 30752 -20182 30960 -20176
rect 31210 -20142 31418 -20136
rect 31210 -20176 31222 -20142
rect 31406 -20176 31418 -20142
rect 31210 -20182 31418 -20176
rect 31668 -20142 31876 -20136
rect 31668 -20176 31680 -20142
rect 31864 -20176 31876 -20142
rect 31668 -20182 31876 -20176
rect 32126 -20142 32334 -20136
rect 32126 -20176 32138 -20142
rect 32322 -20176 32334 -20142
rect 32126 -20182 32334 -20176
rect 32584 -20142 32792 -20136
rect 32584 -20176 32596 -20142
rect 32780 -20176 32792 -20142
rect 32584 -20182 32792 -20176
rect 28812 -20366 28818 -20262
rect 29222 -20290 29236 -20226
rect 29230 -20358 29236 -20290
rect 28812 -20402 28822 -20366
rect 28762 -20556 28822 -20402
rect 29222 -20402 29236 -20358
rect 29270 -20290 29282 -20226
rect 29688 -20226 29734 -20214
rect 29270 -20358 29276 -20290
rect 29270 -20402 29282 -20358
rect 28920 -20452 29128 -20446
rect 28920 -20486 28932 -20452
rect 29116 -20486 29128 -20452
rect 28920 -20492 29128 -20486
rect 28990 -20556 29050 -20492
rect 29222 -20556 29282 -20402
rect 29688 -20402 29694 -20226
rect 29728 -20402 29734 -20226
rect 29688 -20414 29734 -20402
rect 30146 -20226 30192 -20214
rect 30146 -20402 30152 -20226
rect 30186 -20402 30192 -20226
rect 30146 -20414 30192 -20402
rect 30604 -20226 30650 -20214
rect 30604 -20402 30610 -20226
rect 30644 -20402 30650 -20226
rect 30604 -20414 30650 -20402
rect 31062 -20226 31108 -20214
rect 31062 -20402 31068 -20226
rect 31102 -20402 31108 -20226
rect 31062 -20414 31108 -20402
rect 31520 -20226 31566 -20214
rect 31520 -20402 31526 -20226
rect 31560 -20402 31566 -20226
rect 31520 -20414 31566 -20402
rect 31978 -20226 32024 -20214
rect 31978 -20402 31984 -20226
rect 32018 -20402 32024 -20226
rect 31978 -20414 32024 -20402
rect 32436 -20226 32482 -20214
rect 32436 -20402 32442 -20226
rect 32476 -20402 32482 -20226
rect 32886 -20226 32946 -19930
rect 33126 -20136 33186 -19790
rect 33042 -20142 33250 -20136
rect 33042 -20176 33054 -20142
rect 33238 -20176 33250 -20142
rect 33042 -20182 33250 -20176
rect 32886 -20268 32900 -20226
rect 32436 -20414 32482 -20402
rect 32894 -20402 32900 -20268
rect 32934 -20268 32946 -20226
rect 33344 -20226 33404 -19790
rect 33344 -20266 33358 -20226
rect 32934 -20402 32940 -20268
rect 33352 -20356 33358 -20266
rect 32894 -20414 32940 -20402
rect 33342 -20402 33358 -20356
rect 33392 -20266 33404 -20226
rect 33690 -19914 33802 -19790
rect 33392 -20356 33398 -20266
rect 33392 -20402 33402 -20356
rect 29378 -20452 29586 -20446
rect 29378 -20486 29390 -20452
rect 29574 -20486 29586 -20452
rect 29378 -20492 29586 -20486
rect 29836 -20452 30044 -20446
rect 29836 -20486 29848 -20452
rect 30032 -20486 30044 -20452
rect 29836 -20492 30044 -20486
rect 30294 -20452 30502 -20446
rect 30294 -20486 30306 -20452
rect 30490 -20486 30502 -20452
rect 30294 -20492 30502 -20486
rect 30752 -20452 30960 -20446
rect 30752 -20486 30764 -20452
rect 30948 -20486 30960 -20452
rect 30752 -20492 30960 -20486
rect 31210 -20452 31418 -20446
rect 31210 -20486 31222 -20452
rect 31406 -20486 31418 -20452
rect 31210 -20492 31418 -20486
rect 31668 -20452 31876 -20446
rect 31668 -20486 31680 -20452
rect 31864 -20486 31876 -20452
rect 31668 -20492 31876 -20486
rect 32126 -20452 32334 -20446
rect 32126 -20486 32138 -20452
rect 32322 -20486 32334 -20452
rect 32126 -20492 32334 -20486
rect 32584 -20452 32792 -20446
rect 32584 -20486 32596 -20452
rect 32780 -20486 32792 -20452
rect 32584 -20492 32792 -20486
rect 33042 -20452 33250 -20446
rect 33042 -20486 33054 -20452
rect 33238 -20486 33250 -20452
rect 33042 -20492 33250 -20486
rect 28762 -20616 29282 -20556
rect 28762 -21450 28822 -20616
rect 28990 -21450 29050 -20616
rect 29222 -21450 29282 -20616
rect 29448 -20558 29508 -20492
rect 29910 -20558 29970 -20492
rect 30364 -20558 30424 -20492
rect 30826 -20558 30886 -20492
rect 31280 -20558 31340 -20492
rect 31730 -20558 31790 -20492
rect 32196 -20558 32256 -20492
rect 32652 -20558 32712 -20492
rect 29448 -20618 32712 -20558
rect 33116 -21450 33176 -20492
rect 33342 -21450 33402 -20402
rect 23694 -21478 33464 -21450
rect 23694 -21564 23744 -21478
rect 23840 -21564 24324 -21478
rect 24420 -21564 24924 -21478
rect 25020 -21564 25524 -21478
rect 25620 -21564 26124 -21478
rect 26220 -21564 26724 -21478
rect 26820 -21564 27324 -21478
rect 27420 -21564 27924 -21478
rect 28020 -21564 28524 -21478
rect 28620 -21564 29124 -21478
rect 29220 -21564 29724 -21478
rect 29820 -21564 30324 -21478
rect 30420 -21564 30924 -21478
rect 31020 -21564 31524 -21478
rect 31620 -21564 32124 -21478
rect 32220 -21564 32724 -21478
rect 32820 -21564 33324 -21478
rect 33420 -21564 33464 -21478
rect 23694 -21594 33464 -21564
rect 23346 -22042 23458 -21918
rect 24058 -22042 24068 -21742
rect 33080 -22042 33090 -21742
rect 33690 -21918 33696 -19914
rect 33796 -21918 33802 -19914
rect 33690 -22042 33802 -21918
rect 23346 -22048 33802 -22042
rect 23346 -22148 23452 -22048
rect 33696 -22148 33802 -22048
rect 23346 -22154 33802 -22148
<< via1 >>
rect 23440 17094 24040 17394
rect 32072 17094 32672 17394
rect 23562 16868 32558 16978
rect 23602 16606 23662 16666
rect 24622 16606 24682 16666
rect 24620 16006 24680 16066
rect 25060 16006 25120 16066
rect 28056 16606 28116 16666
rect 31486 16612 31546 16672
rect 25900 16006 25960 16066
rect 26336 16006 26396 16066
rect 26770 16006 26830 16066
rect 27632 16006 27692 16066
rect 28052 16006 28112 16066
rect 28484 16006 28544 16066
rect 23602 15414 23662 15474
rect 32494 16612 32554 16672
rect 29340 16006 29400 16066
rect 29770 16006 29830 16066
rect 30202 16006 30262 16066
rect 31052 16006 31112 16066
rect 31486 16006 31546 16066
rect 26340 15414 26400 15474
rect 29770 15414 29830 15474
rect 32494 15414 32554 15474
rect 24534 15078 24594 15138
rect 24664 14934 24724 14994
rect 25528 14934 25588 14994
rect 25656 14936 25716 14996
rect 23080 14100 23140 14160
rect 29994 14368 30054 14374
rect 29994 14320 30000 14368
rect 30000 14320 30048 14368
rect 30048 14320 30054 14368
rect 29994 14314 30054 14320
rect 24530 13504 24590 13564
rect 24664 13386 24724 13446
rect 27152 14096 27252 14196
rect 29356 14116 29416 14176
rect 29848 14170 29908 14176
rect 29848 14128 29856 14170
rect 29856 14128 29904 14170
rect 29904 14128 29908 14170
rect 29848 14116 29908 14128
rect 29526 14058 29586 14064
rect 29526 14010 29532 14058
rect 29532 14010 29580 14058
rect 29580 14010 29586 14058
rect 29526 14004 29586 14010
rect 26304 13382 26364 13442
rect 26442 13384 26502 13444
rect 24664 13104 24724 13164
rect 26304 13102 26364 13162
rect 25098 12990 25158 13050
rect 26808 12990 26868 13050
rect 27246 12990 27306 13050
rect 28526 12990 28586 13050
rect 30244 12990 30304 13050
rect 25096 12438 25156 12498
rect 25530 12438 25590 12498
rect 25952 12438 26012 12498
rect 26378 12438 26438 12498
rect 26812 12438 26872 12498
rect 27246 12438 27306 12498
rect 28102 12438 28162 12498
rect 28966 12438 29026 12498
rect 29386 12438 29446 12498
rect 29818 12438 29878 12498
rect 30248 12438 30308 12498
rect 30672 12438 30732 12498
rect 31104 12438 31164 12498
rect 28526 11874 28586 11934
rect 24176 11572 32038 11716
rect 23440 11162 24040 11462
rect 32072 11162 32672 11462
rect 13066 10328 13448 10628
rect 21200 10328 21878 10628
rect 15134 10064 15230 10150
rect 15714 10064 15810 10150
rect 16314 10064 16410 10150
rect 16914 10064 17010 10150
rect 17514 10064 17610 10150
rect 18114 10064 18210 10150
rect 18714 10064 18810 10150
rect 19314 10064 19410 10150
rect 19914 10064 20010 10150
rect 19048 9812 19108 9872
rect 15612 9132 15672 9192
rect 23648 10328 24248 10628
rect 28280 10328 28880 10628
rect 23896 10064 23992 10150
rect 24476 10064 24572 10150
rect 25076 10064 25172 10150
rect 25676 10064 25772 10150
rect 26276 10064 26372 10150
rect 26876 10064 26972 10150
rect 27476 10064 27572 10150
rect 28076 10064 28172 10150
rect 28676 10064 28772 10150
rect 24600 9258 24660 9318
rect 25062 9258 25122 9318
rect 25516 9260 25576 9320
rect 25978 9258 26038 9318
rect 26432 9258 26492 9318
rect 26882 9258 26942 9318
rect 27348 9258 27408 9318
rect 27804 9258 27864 9318
rect 28038 9050 28098 9110
rect 33086 8977 33182 8996
rect 33086 8943 33139 8977
rect 33139 8943 33173 8977
rect 33173 8943 33182 8977
rect 33086 8924 33182 8943
rect 28038 8708 28098 8768
rect 14008 7978 14068 8038
rect 14464 7978 14524 8038
rect 14924 7978 14984 8038
rect 15380 7978 15440 8038
rect 15838 7978 15898 8038
rect 16302 7978 16362 8038
rect 16756 7978 16816 8038
rect 14012 6004 14072 6064
rect 14468 6004 14528 6064
rect 14928 6004 14988 6064
rect 15384 6004 15444 6064
rect 17216 7978 17276 8038
rect 17446 7978 17506 8038
rect 17674 7978 17734 8038
rect 15842 6004 15902 6064
rect 16306 6004 16366 6064
rect 18130 7978 18190 8038
rect 18590 7978 18650 8038
rect 19046 7978 19106 8038
rect 19502 7978 19562 8038
rect 16756 6004 16816 6064
rect 17212 6004 17272 6064
rect 17680 6004 17740 6064
rect 18138 6004 18198 6064
rect 19958 7978 20018 8038
rect 20416 7978 20476 8038
rect 18594 6004 18654 6064
rect 19050 6004 19110 6064
rect 20876 7978 20936 8038
rect 19506 6004 19566 6064
rect 19962 6004 20022 6064
rect 20420 6004 20480 6064
rect 20880 6004 20940 6064
rect 13308 5346 13404 5432
rect 13908 5346 14004 5432
rect 14508 5346 14604 5432
rect 15108 5346 15204 5432
rect 15708 5346 15804 5432
rect 16308 5346 16404 5432
rect 16908 5346 17004 5432
rect 17508 5346 17604 5432
rect 18108 5346 18204 5432
rect 18708 5346 18804 5432
rect 19308 5346 19404 5432
rect 19908 5346 20004 5432
rect 20508 5346 20604 5432
rect 21108 5346 21204 5432
rect 21528 5346 21624 5432
rect 13066 4872 13448 5172
rect 21200 4872 21878 5172
rect 8458 3990 9058 4290
rect 18090 3990 18690 4290
rect 9310 3730 9406 3816
rect 9910 3730 10006 3816
rect 10510 3730 10606 3816
rect 11110 3730 11206 3816
rect 11710 3730 11806 3816
rect 12310 3730 12406 3816
rect 12910 3730 13006 3816
rect 13510 3730 13606 3816
rect 14110 3730 14206 3816
rect 14710 3730 14806 3816
rect 15310 3730 15406 3816
rect 15910 3730 16006 3816
rect 16510 3730 16606 3816
rect 17110 3730 17206 3816
rect 17530 3730 17626 3816
rect 10014 3098 10074 3158
rect 10470 3098 10530 3158
rect 10930 3098 10990 3158
rect 11386 3098 11446 3158
rect 10010 1124 10070 1184
rect 11844 3098 11904 3158
rect 12308 3098 12368 3158
rect 10466 1124 10526 1184
rect 10926 1124 10986 1184
rect 12758 3098 12818 3158
rect 13214 3098 13274 3158
rect 13682 3098 13742 3158
rect 14140 3098 14200 3158
rect 11382 1124 11442 1184
rect 11840 1124 11900 1184
rect 12304 1124 12364 1184
rect 12758 1124 12818 1184
rect 14596 3098 14656 3158
rect 15052 3098 15112 3158
rect 13216 1180 13276 1184
rect 13216 1132 13222 1180
rect 13222 1132 13270 1180
rect 13270 1132 13276 1180
rect 13216 1124 13276 1132
rect 13450 1136 13510 1196
rect 13676 1126 13736 1184
rect 13676 1124 13736 1126
rect 15508 3098 15568 3158
rect 15964 3098 16024 3158
rect 14132 1124 14192 1184
rect 14592 1124 14652 1184
rect 16422 3098 16482 3158
rect 16882 3098 16942 3158
rect 15048 1124 15108 1184
rect 15504 1124 15564 1184
rect 15960 1124 16020 1184
rect 16418 1124 16478 1184
rect 16878 1124 16938 1184
rect 9224 538 9284 598
rect 12658 436 12718 496
rect 9448 -1140 9508 -1080
rect 9910 -1140 9970 -1080
rect 10364 -1136 10424 -1076
rect 10826 -1136 10886 -1076
rect 11280 -1142 11340 -1082
rect 11730 -1136 11790 -1076
rect 12196 -1136 12256 -1076
rect 12652 -1140 12712 -1080
rect 12886 -1262 12946 -1202
rect 14450 -1140 14510 -1080
rect 14912 -1132 14972 -1072
rect 15366 -1138 15426 -1078
rect 15828 -1138 15888 -1078
rect 16282 -1138 16342 -1078
rect 16732 -1132 16792 -1072
rect 17198 -1138 17258 -1078
rect 17654 -1138 17714 -1078
rect 17886 -1268 17946 -1208
rect 23080 8564 23140 8624
rect 22940 6004 23000 6064
rect 22942 3098 23002 3158
rect 22768 700 22828 760
rect 12886 -1942 12946 -1882
rect 9448 -2076 9508 -2016
rect 9910 -2070 9970 -2010
rect 10364 -2076 10424 -2016
rect 10826 -2070 10886 -2010
rect 11280 -2070 11340 -2010
rect 11730 -2070 11790 -2010
rect 12196 -2076 12256 -2016
rect 12652 -2070 12712 -2010
rect 12650 -3286 12710 -3226
rect 17886 -1930 17946 -1870
rect 14450 -2070 14510 -2010
rect 14912 -2072 14972 -2012
rect 15366 -2072 15426 -2012
rect 15828 -2072 15888 -2012
rect 16282 -2072 16342 -2012
rect 16732 -2066 16792 -2006
rect 17198 -2070 17258 -2010
rect 17654 -2070 17714 -2010
rect 8744 -3564 8840 -3478
rect 9324 -3564 9420 -3478
rect 9924 -3564 10020 -3478
rect 10524 -3564 10620 -3478
rect 11124 -3564 11220 -3478
rect 11724 -3564 11820 -3478
rect 12324 -3564 12420 -3478
rect 12924 -3564 13020 -3478
rect 13524 -3564 13620 -3478
rect 14124 -3564 14220 -3478
rect 14724 -3564 14820 -3478
rect 15324 -3564 15420 -3478
rect 15924 -3564 16020 -3478
rect 16524 -3564 16620 -3478
rect 17124 -3564 17220 -3478
rect 17724 -3564 17820 -3478
rect 18324 -3564 18420 -3478
rect 8458 -4042 9058 -3742
rect 18090 -4042 18690 -3742
rect 12412 -5014 13012 -4714
rect 22044 -5014 22644 -4714
rect 12682 -5278 12778 -5192
rect 13282 -5278 13378 -5192
rect 13882 -5278 13978 -5192
rect 14482 -5278 14578 -5192
rect 15082 -5278 15178 -5192
rect 15682 -5278 15778 -5192
rect 16282 -5278 16378 -5192
rect 16882 -5278 16978 -5192
rect 17482 -5278 17578 -5192
rect 18082 -5278 18178 -5192
rect 18682 -5278 18778 -5192
rect 19282 -5278 19378 -5192
rect 19882 -5278 19978 -5192
rect 20482 -5278 20578 -5192
rect 21082 -5278 21178 -5192
rect 21682 -5278 21778 -5192
rect 22262 -5278 22358 -5192
rect 13388 -6746 13448 -6686
rect 13844 -6746 13904 -6686
rect 14310 -6750 14370 -6690
rect 14760 -6744 14820 -6684
rect 15214 -6744 15274 -6684
rect 15676 -6744 15736 -6684
rect 16130 -6744 16190 -6684
rect 16592 -6746 16652 -6686
rect 13156 -6886 13216 -6826
rect 21596 -5530 21656 -5470
rect 18390 -6746 18450 -6686
rect 18846 -6740 18906 -6680
rect 19312 -6746 19372 -6686
rect 19762 -6746 19822 -6686
rect 20216 -6746 20276 -6686
rect 20678 -6740 20738 -6680
rect 21132 -6746 21192 -6686
rect 21594 -6740 21654 -6680
rect 18156 -6874 18216 -6814
rect 13156 -7548 13216 -7488
rect 13388 -7678 13448 -7618
rect 13844 -7678 13904 -7618
rect 14310 -7684 14370 -7624
rect 14760 -7678 14820 -7618
rect 15214 -7678 15274 -7618
rect 15676 -7678 15736 -7618
rect 16130 -7684 16190 -7624
rect 16592 -7676 16652 -7616
rect 18156 -7554 18216 -7494
rect 18390 -7676 18450 -7616
rect 18846 -7680 18906 -7620
rect 19312 -7680 19372 -7620
rect 19762 -7674 19822 -7614
rect 20216 -7680 20276 -7620
rect 20678 -7680 20738 -7620
rect 21132 -7676 21192 -7616
rect 21594 -7676 21654 -7616
rect 21818 -9354 21878 -9294
rect 14164 -9940 14224 -9880
rect 14624 -9940 14684 -9880
rect 15082 -9940 15142 -9880
rect 15538 -9940 15598 -9880
rect 15994 -9940 16054 -9880
rect 14160 -11914 14220 -11854
rect 14620 -11914 14680 -11854
rect 16450 -9940 16510 -9880
rect 16910 -9940 16970 -9880
rect 15078 -11914 15138 -11854
rect 15534 -11914 15594 -11854
rect 17366 -9882 17426 -9880
rect 17366 -9940 17426 -9882
rect 17592 -9952 17652 -9892
rect 17826 -9888 17886 -9880
rect 17826 -9936 17832 -9888
rect 17832 -9936 17880 -9888
rect 17880 -9936 17886 -9888
rect 17826 -9940 17886 -9936
rect 15990 -11914 16050 -11854
rect 16446 -11914 16506 -11854
rect 18284 -9940 18344 -9880
rect 18738 -9940 18798 -9880
rect 19202 -9940 19262 -9880
rect 19660 -9940 19720 -9880
rect 16902 -11914 16962 -11854
rect 17360 -11914 17420 -11854
rect 17828 -11914 17888 -11854
rect 18284 -11914 18344 -11854
rect 20116 -9940 20176 -9880
rect 20576 -9940 20636 -9880
rect 18734 -11914 18794 -11854
rect 19198 -11914 19258 -11854
rect 21032 -9940 21092 -9880
rect 19656 -11914 19716 -11854
rect 20112 -11914 20172 -11854
rect 20572 -11914 20632 -11854
rect 21028 -11914 21088 -11854
rect 13476 -12572 13572 -12486
rect 13896 -12572 13992 -12486
rect 14496 -12572 14592 -12486
rect 15096 -12572 15192 -12486
rect 15696 -12572 15792 -12486
rect 16296 -12572 16392 -12486
rect 16896 -12572 16992 -12486
rect 17496 -12572 17592 -12486
rect 18096 -12572 18192 -12486
rect 18696 -12572 18792 -12486
rect 19296 -12572 19392 -12486
rect 19896 -12572 19992 -12486
rect 20496 -12572 20592 -12486
rect 21096 -12572 21192 -12486
rect 21696 -12572 21792 -12486
rect 12412 -13046 13012 -12746
rect 22044 -13046 22644 -12746
rect 30826 8642 30886 8648
rect 30826 8594 30832 8642
rect 30832 8594 30880 8642
rect 30880 8594 30886 8642
rect 30826 8588 30886 8594
rect 32954 8678 33014 8684
rect 32954 8630 32960 8678
rect 32960 8630 33008 8678
rect 33008 8630 33014 8678
rect 32954 8624 33014 8630
rect 24600 8390 24660 8450
rect 25062 8390 25122 8450
rect 25516 8390 25576 8450
rect 25978 8390 26038 8450
rect 26432 8390 26492 8450
rect 26882 8390 26942 8450
rect 27348 8390 27408 8450
rect 27804 8390 27864 8450
rect 28038 8396 28098 8456
rect 31930 8562 31990 8568
rect 31930 8514 31936 8562
rect 31936 8514 31984 8562
rect 31984 8514 31990 8562
rect 31930 8508 31990 8514
rect 30406 8380 30502 8452
rect 35784 8380 35880 8452
rect 27812 6818 27872 6878
rect 23824 5346 23920 5432
rect 24424 5346 24520 5432
rect 25024 5346 25120 5432
rect 25624 5346 25720 5432
rect 26224 5346 26320 5432
rect 26824 5346 26920 5432
rect 27424 5346 27520 5432
rect 28024 5346 28120 5432
rect 28624 5346 28720 5432
rect 23648 4872 24248 5172
rect 28280 4872 28880 5172
rect 34630 8314 34690 8320
rect 34630 8266 34636 8314
rect 34636 8266 34684 8314
rect 34684 8266 34690 8314
rect 34630 8260 34690 8266
rect 30570 8190 30630 8196
rect 30570 8142 30576 8190
rect 30576 8142 30624 8190
rect 30624 8142 30630 8190
rect 30570 8136 30630 8142
rect 30826 8238 30886 8244
rect 30826 8190 30832 8238
rect 30832 8190 30880 8238
rect 30880 8190 30886 8238
rect 30826 8184 30886 8190
rect 32952 8202 33012 8208
rect 32952 8154 32964 8202
rect 32964 8154 33012 8202
rect 32952 8148 33012 8154
rect 33524 8238 33584 8244
rect 33524 8190 33530 8238
rect 33530 8190 33578 8238
rect 33578 8190 33584 8238
rect 33524 8184 33584 8190
rect 33268 8148 33328 8154
rect 33268 8100 33274 8148
rect 33274 8100 33322 8148
rect 33322 8100 33328 8148
rect 33268 8094 33328 8100
rect 35652 8202 35712 8208
rect 35652 8154 35658 8202
rect 35658 8154 35706 8202
rect 35706 8154 35712 8202
rect 35652 8148 35712 8154
rect 31930 8016 31990 8022
rect 31930 7968 31936 8016
rect 31936 7968 31984 8016
rect 31984 7968 31990 8016
rect 31930 7962 31990 7968
rect 33086 7836 33182 7908
rect 34628 7776 34688 7782
rect 34628 7728 34634 7776
rect 34634 7728 34682 7776
rect 34682 7728 34688 7776
rect 34628 7722 34688 7728
rect 30570 7644 30630 7650
rect 30570 7596 30576 7644
rect 30576 7596 30624 7644
rect 30624 7596 30630 7644
rect 30570 7590 30630 7596
rect 30826 7554 30886 7560
rect 30826 7506 30832 7554
rect 30832 7506 30880 7554
rect 30880 7506 30886 7554
rect 30826 7500 30886 7506
rect 32954 7590 33014 7596
rect 32954 7542 32960 7590
rect 32960 7542 33012 7590
rect 33012 7542 33014 7590
rect 32954 7536 33014 7542
rect 33268 7604 33328 7610
rect 33268 7556 33274 7604
rect 33274 7556 33322 7604
rect 33322 7556 33328 7604
rect 33268 7550 33328 7556
rect 33524 7554 33584 7560
rect 33524 7506 33530 7554
rect 33530 7506 33578 7554
rect 33578 7506 33584 7554
rect 33524 7500 33584 7506
rect 35652 7590 35712 7596
rect 35652 7542 35658 7590
rect 35658 7542 35706 7590
rect 35706 7542 35712 7590
rect 35652 7536 35712 7542
rect 31930 7472 31990 7478
rect 31930 7424 31936 7472
rect 31936 7424 31984 7472
rect 31984 7424 31990 7472
rect 31930 7418 31990 7424
rect 30406 7292 30502 7364
rect 35784 7292 35880 7364
rect 34628 7232 34688 7238
rect 34628 7184 34634 7232
rect 34634 7184 34682 7232
rect 34682 7184 34688 7232
rect 34628 7178 34688 7184
rect 30570 7100 30630 7106
rect 30570 7052 30576 7100
rect 30576 7052 30624 7100
rect 30624 7052 30630 7100
rect 30570 7046 30630 7052
rect 30826 7150 30886 7156
rect 30826 7102 30832 7150
rect 30832 7102 30880 7150
rect 30880 7102 30886 7150
rect 30826 7096 30886 7102
rect 32954 7114 33014 7120
rect 32954 7066 32960 7114
rect 32960 7066 33008 7114
rect 33008 7066 33014 7114
rect 32954 7060 33014 7066
rect 33524 7150 33584 7156
rect 33524 7102 33530 7150
rect 33530 7102 33578 7150
rect 33578 7102 33584 7150
rect 33524 7096 33584 7102
rect 33268 7060 33328 7066
rect 33268 7012 33274 7060
rect 33274 7012 33322 7060
rect 33322 7012 33328 7060
rect 33268 7006 33328 7012
rect 35652 7114 35712 7120
rect 35652 7066 35658 7114
rect 35658 7066 35710 7114
rect 35710 7066 35712 7114
rect 35652 7060 35712 7066
rect 31930 6928 31990 6934
rect 31930 6880 31936 6928
rect 31936 6880 31984 6928
rect 31984 6880 31990 6928
rect 31930 6874 31990 6880
rect 33086 6748 33182 6820
rect 34628 6688 34688 6694
rect 34628 6640 34634 6688
rect 34634 6640 34682 6688
rect 34682 6640 34688 6688
rect 34628 6634 34688 6640
rect 30570 6556 30630 6562
rect 30570 6508 30576 6556
rect 30576 6508 30624 6556
rect 30624 6508 30630 6556
rect 30570 6502 30630 6508
rect 30826 6466 30886 6472
rect 30826 6418 30832 6466
rect 30832 6418 30880 6466
rect 30880 6418 30886 6466
rect 30826 6412 30886 6418
rect 32954 6502 33014 6508
rect 32954 6454 32960 6502
rect 32960 6454 33008 6502
rect 33008 6454 33014 6502
rect 32954 6448 33014 6454
rect 33268 6514 33328 6520
rect 33268 6466 33274 6514
rect 33274 6466 33322 6514
rect 33322 6466 33328 6514
rect 33268 6460 33328 6466
rect 33524 6466 33584 6472
rect 33524 6418 33530 6466
rect 33530 6418 33578 6466
rect 33578 6418 33584 6466
rect 33524 6412 33584 6418
rect 35650 6502 35710 6508
rect 35650 6454 35662 6502
rect 35662 6454 35710 6502
rect 35650 6448 35710 6454
rect 31930 6386 31990 6392
rect 31930 6338 31936 6386
rect 31936 6338 31984 6386
rect 31984 6338 31990 6386
rect 31930 6332 31990 6338
rect 30406 6204 30502 6276
rect 35784 6204 35880 6276
rect 34628 6142 34688 6148
rect 34628 6094 34634 6142
rect 34634 6094 34682 6142
rect 34682 6094 34688 6142
rect 34628 6088 34688 6094
rect 30570 6014 30630 6020
rect 30570 5966 30576 6014
rect 30576 5966 30624 6014
rect 30624 5966 30630 6014
rect 30570 5960 30630 5966
rect 30826 6062 30886 6068
rect 30826 6014 30832 6062
rect 30832 6014 30880 6062
rect 30880 6014 30886 6062
rect 30826 6008 30886 6014
rect 32954 6026 33014 6032
rect 32954 5978 32960 6026
rect 32960 5978 33012 6026
rect 33012 5978 33014 6026
rect 32954 5972 33014 5978
rect 33276 6032 33336 6038
rect 33276 5984 33282 6032
rect 33282 5984 33330 6032
rect 33330 5984 33336 6032
rect 33276 5978 33336 5984
rect 33524 6062 33584 6068
rect 33524 6014 33530 6062
rect 33530 6014 33578 6062
rect 33578 6014 33584 6062
rect 33524 6008 33584 6014
rect 35652 6026 35712 6032
rect 35652 5978 35658 6026
rect 35658 5978 35706 6026
rect 35706 5978 35712 6026
rect 35652 5972 35712 5978
rect 31930 5842 31990 5848
rect 31930 5794 31936 5842
rect 31936 5794 31984 5842
rect 31984 5794 31990 5842
rect 31930 5788 31990 5794
rect 33086 5660 33182 5732
rect 23458 3990 24058 4290
rect 33090 3990 33690 4290
rect 24310 3730 24406 3816
rect 24910 3730 25006 3816
rect 25510 3730 25606 3816
rect 26110 3730 26206 3816
rect 26710 3730 26806 3816
rect 27310 3730 27406 3816
rect 27910 3730 28006 3816
rect 28510 3730 28606 3816
rect 29110 3730 29206 3816
rect 29710 3730 29806 3816
rect 30310 3730 30406 3816
rect 30910 3730 31006 3816
rect 31510 3730 31606 3816
rect 32110 3730 32206 3816
rect 32530 3730 32626 3816
rect 25014 3098 25074 3158
rect 25470 3098 25530 3158
rect 25930 3098 25990 3158
rect 26386 3098 26446 3158
rect 25010 1124 25070 1184
rect 26844 3098 26904 3158
rect 27308 3098 27368 3158
rect 25466 1124 25526 1184
rect 25926 1124 25986 1184
rect 27758 3098 27818 3158
rect 28214 3098 28274 3158
rect 28682 3098 28742 3158
rect 29140 3098 29200 3158
rect 26382 1124 26442 1184
rect 26840 1124 26900 1184
rect 27304 1124 27364 1184
rect 27758 1124 27818 1184
rect 29596 3098 29656 3158
rect 30052 3098 30112 3158
rect 28216 1180 28276 1184
rect 28216 1132 28222 1180
rect 28222 1132 28270 1180
rect 28270 1132 28276 1180
rect 28216 1124 28276 1132
rect 28450 1136 28510 1196
rect 28676 1126 28736 1184
rect 28676 1124 28736 1126
rect 30508 3098 30568 3158
rect 30964 3098 31024 3158
rect 29132 1124 29192 1184
rect 29592 1124 29652 1184
rect 31422 3098 31482 3158
rect 31882 3098 31942 3158
rect 30048 1124 30108 1184
rect 30504 1124 30564 1184
rect 30960 1124 31020 1184
rect 31418 1124 31478 1184
rect 31878 1124 31938 1184
rect 24224 538 24284 598
rect 24448 -1140 24508 -1080
rect 24910 -1140 24970 -1080
rect 25364 -1136 25424 -1076
rect 25826 -1136 25886 -1076
rect 26280 -1142 26340 -1082
rect 26730 -1136 26790 -1076
rect 27196 -1136 27256 -1076
rect 27652 -1140 27712 -1080
rect 27886 -1262 27946 -1202
rect 29450 -1140 29510 -1080
rect 29912 -1132 29972 -1072
rect 30366 -1138 30426 -1078
rect 30828 -1138 30888 -1078
rect 31282 -1138 31342 -1078
rect 31732 -1132 31792 -1072
rect 32198 -1138 32258 -1078
rect 32654 -1138 32714 -1078
rect 32886 -1268 32946 -1208
rect 23080 -3286 23140 -3226
rect 22940 -9940 23000 -9880
rect 8458 -14010 9058 -13710
rect 18090 -14010 18690 -13710
rect 9310 -14270 9406 -14184
rect 9910 -14270 10006 -14184
rect 10510 -14270 10606 -14184
rect 11110 -14270 11206 -14184
rect 11710 -14270 11806 -14184
rect 12310 -14270 12406 -14184
rect 12910 -14270 13006 -14184
rect 13510 -14270 13606 -14184
rect 14110 -14270 14206 -14184
rect 14710 -14270 14806 -14184
rect 15310 -14270 15406 -14184
rect 15910 -14270 16006 -14184
rect 16510 -14270 16606 -14184
rect 17110 -14270 17206 -14184
rect 17530 -14270 17626 -14184
rect 10014 -14902 10074 -14842
rect 10470 -14902 10530 -14842
rect 10930 -14902 10990 -14842
rect 11386 -14902 11446 -14842
rect 10010 -16876 10070 -16816
rect 11844 -14902 11904 -14842
rect 12308 -14902 12368 -14842
rect 10466 -16876 10526 -16816
rect 10926 -16876 10986 -16816
rect 12758 -14902 12818 -14842
rect 13214 -14902 13274 -14842
rect 13682 -14902 13742 -14842
rect 14140 -14902 14200 -14842
rect 11382 -16876 11442 -16816
rect 11840 -16876 11900 -16816
rect 12304 -16876 12364 -16816
rect 12758 -16876 12818 -16816
rect 14596 -14902 14656 -14842
rect 15052 -14902 15112 -14842
rect 13216 -16820 13276 -16816
rect 13216 -16868 13222 -16820
rect 13222 -16868 13270 -16820
rect 13270 -16868 13276 -16820
rect 13216 -16876 13276 -16868
rect 13450 -16864 13510 -16804
rect 13676 -16874 13736 -16816
rect 13676 -16876 13736 -16874
rect 15508 -14902 15568 -14842
rect 15964 -14902 16024 -14842
rect 14132 -16876 14192 -16816
rect 14592 -16876 14652 -16816
rect 16422 -14902 16482 -14842
rect 16882 -14902 16942 -14842
rect 15048 -16876 15108 -16816
rect 15504 -16876 15564 -16816
rect 15960 -16876 16020 -16816
rect 16418 -16876 16478 -16816
rect 16878 -16876 16938 -16816
rect 9224 -17462 9284 -17402
rect 9448 -19140 9508 -19080
rect 9910 -19140 9970 -19080
rect 10364 -19136 10424 -19076
rect 10826 -19136 10886 -19076
rect 11280 -19142 11340 -19082
rect 11730 -19136 11790 -19076
rect 12196 -19136 12256 -19076
rect 12652 -19140 12712 -19080
rect 12886 -19262 12946 -19202
rect 14450 -19140 14510 -19080
rect 14912 -19132 14972 -19072
rect 15366 -19138 15426 -19078
rect 15828 -19138 15888 -19078
rect 16282 -19138 16342 -19078
rect 16732 -19132 16792 -19072
rect 17198 -19138 17258 -19078
rect 17654 -19138 17714 -19078
rect 17886 -19268 17946 -19208
rect 27886 -1942 27946 -1882
rect 24448 -2076 24508 -2016
rect 24910 -2070 24970 -2010
rect 25364 -2076 25424 -2016
rect 25826 -2070 25886 -2010
rect 26280 -2070 26340 -2010
rect 26730 -2070 26790 -2010
rect 27196 -2076 27256 -2016
rect 27652 -2070 27712 -2010
rect 24448 -3286 24508 -3226
rect 32886 -1930 32946 -1870
rect 29450 -2070 29510 -2010
rect 29912 -2072 29972 -2012
rect 30366 -2072 30426 -2012
rect 30828 -2072 30888 -2012
rect 31282 -2072 31342 -2012
rect 31732 -2066 31792 -2006
rect 32198 -2070 32258 -2010
rect 32654 -2070 32714 -2010
rect 23744 -3564 23840 -3478
rect 24324 -3564 24420 -3478
rect 24924 -3564 25020 -3478
rect 25524 -3564 25620 -3478
rect 26124 -3564 26220 -3478
rect 26724 -3564 26820 -3478
rect 27324 -3564 27420 -3478
rect 27924 -3564 28020 -3478
rect 28524 -3564 28620 -3478
rect 29124 -3564 29220 -3478
rect 29724 -3564 29820 -3478
rect 30324 -3564 30420 -3478
rect 30924 -3564 31020 -3478
rect 31524 -3564 31620 -3478
rect 32124 -3564 32220 -3478
rect 32724 -3564 32820 -3478
rect 33324 -3564 33420 -3478
rect 23458 -4042 24058 -3742
rect 33090 -4042 33690 -3742
rect 23080 -5530 23140 -5470
rect 22940 -16876 23000 -16816
rect 12886 -19942 12946 -19882
rect 9448 -20076 9508 -20016
rect 9910 -20070 9970 -20010
rect 10364 -20076 10424 -20016
rect 10826 -20070 10886 -20010
rect 11280 -20070 11340 -20010
rect 11730 -20070 11790 -20010
rect 12196 -20076 12256 -20016
rect 12652 -20070 12712 -20010
rect 12652 -21286 12712 -21226
rect 17886 -19930 17946 -19870
rect 14450 -20070 14510 -20010
rect 14912 -20072 14972 -20012
rect 15366 -20072 15426 -20012
rect 15828 -20072 15888 -20012
rect 16282 -20072 16342 -20012
rect 16732 -20066 16792 -20006
rect 17198 -20070 17258 -20010
rect 17654 -20070 17714 -20010
rect 8744 -21564 8840 -21478
rect 9324 -21564 9420 -21478
rect 9924 -21564 10020 -21478
rect 10524 -21564 10620 -21478
rect 11124 -21564 11220 -21478
rect 11724 -21564 11820 -21478
rect 12324 -21564 12420 -21478
rect 12924 -21564 13020 -21478
rect 13524 -21564 13620 -21478
rect 14124 -21564 14220 -21478
rect 14724 -21564 14820 -21478
rect 15324 -21564 15420 -21478
rect 15924 -21564 16020 -21478
rect 16524 -21564 16620 -21478
rect 17124 -21564 17220 -21478
rect 17724 -21564 17820 -21478
rect 18324 -21564 18420 -21478
rect 8458 -22042 9058 -21742
rect 18090 -22042 18690 -21742
rect 27412 -5014 28012 -4714
rect 37044 -5014 37644 -4714
rect 27682 -5278 27778 -5192
rect 28282 -5278 28378 -5192
rect 28882 -5278 28978 -5192
rect 29482 -5278 29578 -5192
rect 30082 -5278 30178 -5192
rect 30682 -5278 30778 -5192
rect 31282 -5278 31378 -5192
rect 31882 -5278 31978 -5192
rect 32482 -5278 32578 -5192
rect 33082 -5278 33178 -5192
rect 33682 -5278 33778 -5192
rect 34282 -5278 34378 -5192
rect 34882 -5278 34978 -5192
rect 35482 -5278 35578 -5192
rect 36082 -5278 36178 -5192
rect 36682 -5278 36778 -5192
rect 37262 -5278 37358 -5192
rect 28388 -6746 28448 -6686
rect 28844 -6746 28904 -6686
rect 29310 -6750 29370 -6690
rect 29760 -6744 29820 -6684
rect 30214 -6744 30274 -6684
rect 30676 -6744 30736 -6684
rect 31130 -6744 31190 -6684
rect 31592 -6746 31652 -6686
rect 28156 -6886 28216 -6826
rect 33390 -5530 33450 -5470
rect 33390 -6746 33450 -6686
rect 33846 -6740 33906 -6680
rect 34312 -6746 34372 -6686
rect 34762 -6746 34822 -6686
rect 35216 -6746 35276 -6686
rect 35678 -6740 35738 -6680
rect 36132 -6746 36192 -6686
rect 36594 -6740 36654 -6680
rect 33156 -6874 33216 -6814
rect 28156 -7548 28216 -7488
rect 28388 -7678 28448 -7618
rect 28844 -7678 28904 -7618
rect 29310 -7684 29370 -7624
rect 29760 -7678 29820 -7618
rect 30214 -7678 30274 -7618
rect 30676 -7678 30736 -7618
rect 31130 -7684 31190 -7624
rect 31592 -7676 31652 -7616
rect 33156 -7554 33216 -7494
rect 33390 -7676 33450 -7616
rect 33846 -7680 33906 -7620
rect 34312 -7680 34372 -7620
rect 34762 -7674 34822 -7614
rect 35216 -7680 35276 -7620
rect 35678 -7680 35738 -7620
rect 36132 -7676 36192 -7616
rect 36594 -7676 36654 -7616
rect 36818 -9354 36878 -9294
rect 29164 -9940 29224 -9880
rect 29624 -9940 29684 -9880
rect 30082 -9940 30142 -9880
rect 30538 -9940 30598 -9880
rect 30994 -9940 31054 -9880
rect 29160 -11914 29220 -11854
rect 29620 -11914 29680 -11854
rect 31450 -9940 31510 -9880
rect 31910 -9940 31970 -9880
rect 30078 -11914 30138 -11854
rect 30534 -11914 30594 -11854
rect 32366 -9882 32426 -9880
rect 32366 -9940 32426 -9882
rect 32592 -9952 32652 -9892
rect 32826 -9888 32886 -9880
rect 32826 -9936 32832 -9888
rect 32832 -9936 32880 -9888
rect 32880 -9936 32886 -9888
rect 32826 -9940 32886 -9936
rect 30990 -11914 31050 -11854
rect 31446 -11914 31506 -11854
rect 33284 -9940 33344 -9880
rect 33738 -9940 33798 -9880
rect 34202 -9940 34262 -9880
rect 34660 -9940 34720 -9880
rect 31902 -11914 31962 -11854
rect 32360 -11914 32420 -11854
rect 32828 -11914 32888 -11854
rect 33284 -11914 33344 -11854
rect 35116 -9940 35176 -9880
rect 35576 -9940 35636 -9880
rect 33734 -11914 33794 -11854
rect 34198 -11914 34258 -11854
rect 36032 -9940 36092 -9880
rect 34656 -11914 34716 -11854
rect 35112 -11914 35172 -11854
rect 35572 -11914 35632 -11854
rect 36028 -11914 36088 -11854
rect 28476 -12572 28572 -12486
rect 28896 -12572 28992 -12486
rect 29496 -12572 29592 -12486
rect 30096 -12572 30192 -12486
rect 30696 -12572 30792 -12486
rect 31296 -12572 31392 -12486
rect 31896 -12572 31992 -12486
rect 32496 -12572 32592 -12486
rect 33096 -12572 33192 -12486
rect 33696 -12572 33792 -12486
rect 34296 -12572 34392 -12486
rect 34896 -12572 34992 -12486
rect 35496 -12572 35592 -12486
rect 36096 -12572 36192 -12486
rect 36696 -12572 36792 -12486
rect 27412 -13046 28012 -12746
rect 37044 -13046 37644 -12746
rect 23458 -14010 24058 -13710
rect 33090 -14010 33690 -13710
rect 24310 -14270 24406 -14184
rect 24910 -14270 25006 -14184
rect 25510 -14270 25606 -14184
rect 26110 -14270 26206 -14184
rect 26710 -14270 26806 -14184
rect 27310 -14270 27406 -14184
rect 27910 -14270 28006 -14184
rect 28510 -14270 28606 -14184
rect 29110 -14270 29206 -14184
rect 29710 -14270 29806 -14184
rect 30310 -14270 30406 -14184
rect 30910 -14270 31006 -14184
rect 31510 -14270 31606 -14184
rect 32110 -14270 32206 -14184
rect 32530 -14270 32626 -14184
rect 25014 -14902 25074 -14842
rect 25470 -14902 25530 -14842
rect 25930 -14902 25990 -14842
rect 26386 -14902 26446 -14842
rect 25010 -16876 25070 -16816
rect 26844 -14902 26904 -14842
rect 27308 -14902 27368 -14842
rect 25466 -16876 25526 -16816
rect 25926 -16876 25986 -16816
rect 27758 -14902 27818 -14842
rect 28214 -14902 28274 -14842
rect 28682 -14902 28742 -14842
rect 29140 -14902 29200 -14842
rect 26382 -16876 26442 -16816
rect 26840 -16876 26900 -16816
rect 27304 -16876 27364 -16816
rect 27758 -16876 27818 -16816
rect 29596 -14902 29656 -14842
rect 30052 -14902 30112 -14842
rect 28216 -16820 28276 -16816
rect 28216 -16868 28222 -16820
rect 28222 -16868 28270 -16820
rect 28270 -16868 28276 -16820
rect 28216 -16876 28276 -16868
rect 28450 -16864 28510 -16804
rect 28676 -16874 28736 -16816
rect 28676 -16876 28736 -16874
rect 30508 -14902 30568 -14842
rect 30964 -14902 31024 -14842
rect 29132 -16876 29192 -16816
rect 29592 -16876 29652 -16816
rect 31422 -14902 31482 -14842
rect 31882 -14902 31942 -14842
rect 30048 -16876 30108 -16816
rect 30504 -16876 30564 -16816
rect 30960 -16876 31020 -16816
rect 31418 -16876 31478 -16816
rect 31878 -16876 31938 -16816
rect 24224 -17462 24284 -17402
rect 24448 -19140 24508 -19080
rect 24910 -19140 24970 -19080
rect 25364 -19136 25424 -19076
rect 25826 -19136 25886 -19076
rect 26280 -19142 26340 -19082
rect 26730 -19136 26790 -19076
rect 27196 -19136 27256 -19076
rect 27652 -19140 27712 -19080
rect 27886 -19262 27946 -19202
rect 29450 -19140 29510 -19080
rect 29912 -19132 29972 -19072
rect 30366 -19138 30426 -19078
rect 30828 -19138 30888 -19078
rect 31282 -19138 31342 -19078
rect 31732 -19132 31792 -19072
rect 32198 -19138 32258 -19078
rect 32654 -19138 32714 -19078
rect 32886 -19268 32946 -19208
rect 23080 -21286 23140 -21226
rect 27886 -19942 27946 -19882
rect 24448 -20076 24508 -20016
rect 24910 -20070 24970 -20010
rect 25364 -20076 25424 -20016
rect 25826 -20070 25886 -20010
rect 26280 -20070 26340 -20010
rect 26730 -20070 26790 -20010
rect 27196 -20076 27256 -20016
rect 27652 -20070 27712 -20010
rect 24448 -21286 24508 -21226
rect 32886 -19930 32946 -19870
rect 29450 -20070 29510 -20010
rect 29912 -20072 29972 -20012
rect 30366 -20072 30426 -20012
rect 30828 -20072 30888 -20012
rect 31282 -20072 31342 -20012
rect 31732 -20066 31792 -20006
rect 32198 -20070 32258 -20010
rect 32654 -20070 32714 -20010
rect 23744 -21564 23840 -21478
rect 24324 -21564 24420 -21478
rect 24924 -21564 25020 -21478
rect 25524 -21564 25620 -21478
rect 26124 -21564 26220 -21478
rect 26724 -21564 26820 -21478
rect 27324 -21564 27420 -21478
rect 27924 -21564 28020 -21478
rect 28524 -21564 28620 -21478
rect 29124 -21564 29220 -21478
rect 29724 -21564 29820 -21478
rect 30324 -21564 30420 -21478
rect 30924 -21564 31020 -21478
rect 31524 -21564 31620 -21478
rect 32124 -21564 32220 -21478
rect 32724 -21564 32820 -21478
rect 33324 -21564 33420 -21478
rect 23458 -22042 24058 -21742
rect 33090 -22042 33690 -21742
<< metal2 >>
rect 23440 17394 24040 17404
rect 23440 17084 24040 17094
rect 32072 17394 32672 17404
rect 32072 17084 32672 17094
rect 23526 16978 32596 17012
rect 23526 16868 23562 16978
rect 32558 16868 32596 16978
rect 23526 16830 32596 16868
rect 31486 16672 31546 16678
rect 32494 16672 32554 16678
rect 23602 16666 23662 16672
rect 24622 16666 24682 16672
rect 28056 16666 28116 16672
rect 23662 16606 24622 16666
rect 24682 16606 28056 16666
rect 31546 16612 32494 16672
rect 31486 16606 31546 16612
rect 32494 16606 32554 16612
rect 23602 16600 23662 16606
rect 24622 16600 24682 16606
rect 28056 16600 28116 16606
rect 24620 16066 24680 16072
rect 25060 16066 25120 16072
rect 25900 16066 25960 16072
rect 26336 16066 26396 16072
rect 26770 16066 26830 16072
rect 27632 16066 27692 16072
rect 28052 16066 28112 16072
rect 28484 16066 28544 16072
rect 29340 16066 29400 16072
rect 29770 16066 29830 16072
rect 30202 16066 30262 16072
rect 31052 16066 31112 16072
rect 31486 16066 31546 16072
rect 23480 16006 24620 16066
rect 24680 16006 25060 16066
rect 25120 16006 25900 16066
rect 25960 16006 26336 16066
rect 26396 16006 26770 16066
rect 26830 16006 27632 16066
rect 27692 16006 28052 16066
rect 28112 16006 28484 16066
rect 28544 16006 29340 16066
rect 29400 16006 29770 16066
rect 29830 16006 30202 16066
rect 30262 16006 31052 16066
rect 31112 16006 31486 16066
rect 23480 14870 23540 16006
rect 24620 16000 24680 16006
rect 25060 16000 25120 16006
rect 25900 16000 25960 16006
rect 26336 16000 26396 16006
rect 26770 16000 26830 16006
rect 27632 16000 27692 16006
rect 28052 16000 28112 16006
rect 28484 16000 28544 16006
rect 29340 16000 29400 16006
rect 29770 16000 29830 16006
rect 30202 16000 30262 16006
rect 31052 16000 31112 16006
rect 31486 16000 31546 16006
rect 23602 15474 23662 15480
rect 26340 15474 26400 15480
rect 29770 15474 29830 15480
rect 32494 15474 32554 15480
rect 23662 15414 26340 15474
rect 26400 15414 29770 15474
rect 29830 15414 32494 15474
rect 23602 15408 23662 15414
rect 24394 14994 24454 15414
rect 26340 15408 26400 15414
rect 29770 15408 29830 15414
rect 32494 15408 32554 15414
rect 24534 15138 24594 15144
rect 24594 15078 30054 15138
rect 24534 15072 24594 15078
rect 24664 14994 24724 15000
rect 25528 14994 25588 15000
rect 24394 14934 24664 14994
rect 24724 14934 25528 14994
rect 24664 14928 24724 14934
rect 25528 14928 25588 14934
rect 25656 14996 25716 15002
rect 25716 14936 29908 14996
rect 25656 14930 25716 14936
rect 23480 14810 23878 14870
rect 23074 14100 23080 14160
rect 23140 14100 23146 14160
rect 13066 10628 13448 10638
rect 13066 10318 13448 10328
rect 21200 10628 21878 10638
rect 21200 10318 21878 10328
rect 15084 10150 20056 10180
rect 15084 10064 15134 10150
rect 15230 10064 15714 10150
rect 15810 10064 16314 10150
rect 16410 10064 16914 10150
rect 17010 10064 17514 10150
rect 17610 10064 18114 10150
rect 18210 10064 18714 10150
rect 18810 10064 19314 10150
rect 19410 10064 19914 10150
rect 20010 10064 20056 10150
rect 15084 10036 20056 10064
rect 19048 9872 19108 9878
rect 23080 9872 23140 14100
rect 23818 11934 23878 14810
rect 27152 14196 27252 14202
rect 27148 14101 27152 14191
rect 27252 14101 27256 14191
rect 29848 14176 29908 14936
rect 29994 14374 30054 15078
rect 29988 14314 29994 14374
rect 30054 14314 30060 14374
rect 29350 14116 29356 14176
rect 29416 14116 29422 14176
rect 29842 14116 29848 14176
rect 29908 14116 29914 14176
rect 27152 14090 27252 14096
rect 29356 13788 29416 14116
rect 29520 14004 29526 14064
rect 29586 14004 29592 14064
rect 27042 13728 29416 13788
rect 24530 13564 24590 13570
rect 27042 13564 27102 13728
rect 24590 13504 27102 13564
rect 24530 13498 24590 13504
rect 24658 13386 24664 13446
rect 24724 13386 24730 13446
rect 26304 13442 26364 13448
rect 24664 13164 24724 13386
rect 24658 13104 24664 13164
rect 24724 13104 24730 13164
rect 26304 13162 26364 13382
rect 26442 13444 26502 13450
rect 29526 13444 29586 14004
rect 34621 13582 34630 13642
rect 34690 13582 34699 13642
rect 26502 13384 29586 13444
rect 26442 13378 26502 13384
rect 26298 13102 26304 13162
rect 26364 13102 26370 13162
rect 25098 13050 25158 13056
rect 26808 13050 26868 13056
rect 27246 13050 27306 13056
rect 28526 13050 28586 13056
rect 30244 13050 30304 13056
rect 25158 12990 26808 13050
rect 26868 12990 27246 13050
rect 27306 12990 28526 13050
rect 28586 12990 30244 13050
rect 25098 12984 25158 12990
rect 26808 12984 26868 12990
rect 27246 12984 27306 12990
rect 28526 12984 28586 12990
rect 30244 12984 30304 12990
rect 25096 12498 25156 12504
rect 25530 12498 25590 12504
rect 25952 12498 26012 12504
rect 26378 12498 26438 12504
rect 26812 12498 26872 12504
rect 27246 12498 27306 12504
rect 28102 12498 28162 12504
rect 28966 12498 29026 12504
rect 29386 12498 29446 12504
rect 29818 12498 29878 12504
rect 30248 12498 30308 12504
rect 30672 12498 30732 12504
rect 31104 12498 31164 12504
rect 25156 12438 25530 12498
rect 25590 12438 25952 12498
rect 26012 12438 26378 12498
rect 26438 12438 26812 12498
rect 26872 12438 27246 12498
rect 27306 12438 28102 12498
rect 28162 12438 28966 12498
rect 29026 12438 29386 12498
rect 29446 12438 29818 12498
rect 29878 12438 30248 12498
rect 30308 12438 30672 12498
rect 30732 12438 31104 12498
rect 31164 12438 32238 12498
rect 25096 12432 25156 12438
rect 25530 12432 25590 12438
rect 25952 12432 26012 12438
rect 26378 12432 26438 12438
rect 26812 12432 26872 12438
rect 27246 12432 27306 12438
rect 28102 12432 28162 12438
rect 28966 12432 29026 12438
rect 29386 12432 29446 12438
rect 29818 12432 29878 12438
rect 30248 12432 30308 12438
rect 30672 12432 30732 12438
rect 31104 12432 31164 12438
rect 28526 11934 28586 11940
rect 23818 11874 28526 11934
rect 28526 11868 28586 11874
rect 24136 11716 32076 11756
rect 24136 11572 24176 11716
rect 32038 11572 32076 11716
rect 24136 11542 32076 11572
rect 23440 11462 24040 11472
rect 23440 11152 24040 11162
rect 32072 11462 32672 11472
rect 32072 11152 32672 11162
rect 23648 10628 24248 10638
rect 23648 10318 24248 10328
rect 28280 10628 28880 10638
rect 28280 10318 28880 10328
rect 23846 10150 28818 10180
rect 23846 10064 23896 10150
rect 23992 10064 24476 10150
rect 24572 10064 25076 10150
rect 25172 10064 25676 10150
rect 25772 10064 26276 10150
rect 26372 10064 26876 10150
rect 26972 10064 27476 10150
rect 27572 10064 28076 10150
rect 28172 10064 28676 10150
rect 28772 10064 28818 10150
rect 23846 10036 28818 10064
rect 19108 9812 23140 9872
rect 19048 9806 19108 9812
rect 15606 9132 15612 9192
rect 15672 9132 15678 9192
rect 14008 8038 14068 8044
rect 14464 8038 14524 8044
rect 14924 8038 14984 8044
rect 15380 8038 15440 8044
rect 15612 8038 15672 9132
rect 23080 8624 23140 9812
rect 24600 9318 24660 9324
rect 23074 8564 23080 8624
rect 23140 8564 23146 8624
rect 24600 8450 24660 9258
rect 24600 8384 24660 8390
rect 25062 9318 25122 9324
rect 25062 8450 25122 9258
rect 25516 9320 25576 9326
rect 25516 8450 25576 9260
rect 25978 9318 26038 9324
rect 25978 8450 26038 9258
rect 26432 9318 26492 9324
rect 26432 8450 26492 9258
rect 26882 9318 26942 9324
rect 26882 8450 26942 9258
rect 27348 9318 27408 9324
rect 27348 8450 27408 9258
rect 27804 9318 27864 9324
rect 27804 8450 27864 9258
rect 28038 9110 28098 9116
rect 28038 8768 28098 9050
rect 33074 8996 33194 9008
rect 33074 8924 33086 8996
rect 33182 8924 33194 8996
rect 33074 8912 33194 8924
rect 28032 8708 28038 8768
rect 28098 8708 28104 8768
rect 28038 8456 28098 8708
rect 30826 8648 32954 8684
rect 30886 8624 32954 8648
rect 33014 8624 33020 8684
rect 30826 8582 30886 8588
rect 31930 8568 31990 8574
rect 25510 8390 25516 8450
rect 25576 8390 25582 8450
rect 25972 8390 25978 8450
rect 26038 8390 26044 8450
rect 26876 8390 26882 8450
rect 26942 8390 26948 8450
rect 27342 8390 27348 8450
rect 27408 8390 27414 8450
rect 28032 8396 28038 8456
rect 28098 8396 28104 8456
rect 30394 8452 30514 8464
rect 25062 8384 25122 8390
rect 26432 8384 26492 8390
rect 27804 8384 27864 8390
rect 30394 8380 30406 8452
rect 30502 8380 30514 8452
rect 31930 8448 31990 8508
rect 30394 8368 30514 8380
rect 30570 8388 31990 8448
rect 30570 8196 30630 8388
rect 34630 8320 34690 13582
rect 35772 8452 35892 8464
rect 35772 8380 35784 8452
rect 35880 8380 35892 8452
rect 35772 8368 35892 8380
rect 34624 8260 34630 8320
rect 34690 8260 34696 8320
rect 30826 8244 30886 8250
rect 33524 8244 33584 8250
rect 32952 8208 33018 8214
rect 30886 8184 32952 8208
rect 30826 8148 32952 8184
rect 33012 8148 33018 8208
rect 33584 8184 35652 8208
rect 32952 8142 33018 8148
rect 33268 8154 33328 8160
rect 30570 8130 30630 8136
rect 33524 8148 35652 8184
rect 35712 8148 35718 8208
rect 15838 8038 15898 8044
rect 16302 8038 16362 8044
rect 16756 8038 16816 8044
rect 17216 8038 17276 8044
rect 17446 8038 17506 8044
rect 17674 8038 17734 8044
rect 18130 8038 18190 8044
rect 18590 8038 18650 8044
rect 19046 8038 19106 8044
rect 19502 8038 19562 8044
rect 19958 8038 20018 8044
rect 20416 8038 20476 8044
rect 20876 8038 20936 8044
rect 14068 7978 14464 8038
rect 14524 7978 14924 8038
rect 14984 7978 15380 8038
rect 15440 7978 15838 8038
rect 15898 7978 16302 8038
rect 16362 7978 16756 8038
rect 16816 7978 17216 8038
rect 17276 7978 17446 8038
rect 17506 7978 17674 8038
rect 17734 7978 18130 8038
rect 18190 7978 18590 8038
rect 18650 7978 19046 8038
rect 19106 7978 19502 8038
rect 19562 7978 19958 8038
rect 20018 7978 20416 8038
rect 20476 7978 20876 8038
rect 14008 7972 14068 7978
rect 14464 7972 14524 7978
rect 14924 7972 14984 7978
rect 15380 7972 15440 7978
rect 15838 7972 15898 7978
rect 16302 7972 16362 7978
rect 16756 7972 16816 7978
rect 17216 7972 17276 7978
rect 17446 7972 17506 7978
rect 17674 7972 17734 7978
rect 18130 7972 18190 7978
rect 18590 7972 18650 7978
rect 19046 7972 19106 7978
rect 19502 7972 19562 7978
rect 19958 7972 20018 7978
rect 20416 7972 20476 7978
rect 20876 7972 20936 7978
rect 31930 8022 31990 8028
rect 31930 7902 31990 7962
rect 30570 7842 31990 7902
rect 33074 7908 33194 7920
rect 30570 7650 30630 7842
rect 33074 7836 33086 7908
rect 33182 7836 33194 7908
rect 33268 7902 33328 8094
rect 33268 7842 34688 7902
rect 33074 7824 33194 7836
rect 34628 7782 34688 7842
rect 34628 7716 34688 7722
rect 33268 7610 33328 7616
rect 30570 7584 30630 7590
rect 30826 7560 32954 7596
rect 30886 7536 32954 7560
rect 33014 7536 33020 7596
rect 30826 7494 30886 7500
rect 31930 7478 31990 7484
rect 30394 7364 30514 7376
rect 30394 7292 30406 7364
rect 30502 7292 30514 7364
rect 31930 7358 31990 7418
rect 30394 7280 30514 7292
rect 30570 7298 31990 7358
rect 33268 7358 33328 7550
rect 33524 7560 35652 7596
rect 33584 7536 35652 7560
rect 35712 7536 35718 7596
rect 33524 7494 33584 7500
rect 35772 7364 35892 7376
rect 33268 7298 34688 7358
rect 30570 7106 30630 7298
rect 34628 7238 34688 7298
rect 35772 7292 35784 7364
rect 35880 7292 35892 7364
rect 35772 7280 35892 7292
rect 34628 7172 34688 7178
rect 30826 7156 30886 7162
rect 33524 7156 33584 7162
rect 30886 7096 32954 7120
rect 30826 7060 32954 7096
rect 33014 7060 33020 7120
rect 33584 7096 35652 7120
rect 33268 7066 33328 7072
rect 30570 7040 30630 7046
rect 33524 7060 35652 7096
rect 35712 7060 35718 7120
rect 31930 6934 31990 6940
rect 27812 6878 27872 6884
rect 27872 6818 29436 6878
rect 27812 6812 27872 6818
rect 14012 6064 14072 6070
rect 14468 6064 14528 6070
rect 14928 6064 14988 6070
rect 15384 6064 15444 6070
rect 15842 6064 15902 6070
rect 16306 6064 16366 6070
rect 16756 6064 16816 6070
rect 17212 6064 17272 6070
rect 17680 6064 17740 6070
rect 18138 6064 18198 6070
rect 18594 6064 18654 6070
rect 19050 6064 19110 6070
rect 19506 6064 19566 6070
rect 19962 6064 20022 6070
rect 20420 6064 20480 6070
rect 20880 6064 20940 6070
rect 22940 6064 23000 6070
rect 14072 6004 14468 6064
rect 14528 6004 14928 6064
rect 14988 6004 15384 6064
rect 15444 6004 15842 6064
rect 15902 6004 16306 6064
rect 16366 6004 16756 6064
rect 16816 6004 17212 6064
rect 17272 6004 17680 6064
rect 17740 6004 18138 6064
rect 18198 6004 18594 6064
rect 18654 6004 19050 6064
rect 19110 6004 19506 6064
rect 19566 6004 19962 6064
rect 20022 6004 20420 6064
rect 20480 6004 20880 6064
rect 20940 6004 22940 6064
rect 14012 5998 14072 6004
rect 14468 5998 14528 6004
rect 14928 5998 14988 6004
rect 15384 5998 15444 6004
rect 15842 5998 15902 6004
rect 16306 5998 16366 6004
rect 16756 5998 16816 6004
rect 17212 5998 17272 6004
rect 17680 5998 17740 6004
rect 18138 5998 18198 6004
rect 18594 5998 18654 6004
rect 19050 5998 19110 6004
rect 19506 5998 19566 6004
rect 19962 5998 20022 6004
rect 20420 5998 20480 6004
rect 20880 5998 20940 6004
rect 22940 5998 23000 6004
rect 29336 5476 29436 6818
rect 31930 6814 31990 6874
rect 30570 6754 31990 6814
rect 33074 6820 33194 6832
rect 30570 6562 30630 6754
rect 33074 6748 33086 6820
rect 33182 6748 33194 6820
rect 33268 6814 33328 7006
rect 33268 6754 34688 6814
rect 33074 6736 33194 6748
rect 34628 6694 34688 6754
rect 34628 6628 34688 6634
rect 33268 6520 33328 6526
rect 30570 6496 30630 6502
rect 30826 6472 32954 6508
rect 30886 6448 32954 6472
rect 33014 6448 33020 6508
rect 35650 6508 35716 6514
rect 30826 6406 30886 6412
rect 31930 6392 31990 6398
rect 30394 6276 30514 6288
rect 30394 6204 30406 6276
rect 30502 6204 30514 6276
rect 31930 6272 31990 6332
rect 30394 6192 30514 6204
rect 30570 6212 31990 6272
rect 33268 6268 33328 6460
rect 33524 6472 35650 6508
rect 33584 6448 35650 6472
rect 35710 6448 35716 6508
rect 35650 6442 35716 6448
rect 33524 6406 33584 6412
rect 35772 6276 35892 6288
rect 30570 6020 30630 6212
rect 33268 6208 34688 6268
rect 34628 6148 34688 6208
rect 35772 6204 35784 6276
rect 35880 6204 35892 6276
rect 35772 6192 35892 6204
rect 34628 6082 34688 6088
rect 30826 6068 30886 6074
rect 33524 6068 33584 6074
rect 33276 6038 33336 6044
rect 30886 6008 32954 6032
rect 30826 5972 32954 6008
rect 33014 5972 33020 6032
rect 33170 5978 33276 6038
rect 30570 5954 30630 5960
rect 31930 5848 31990 5854
rect 33170 5848 33230 5978
rect 33276 5972 33336 5978
rect 33584 6008 35652 6032
rect 33524 5972 35652 6008
rect 35712 5972 35718 6032
rect 31990 5788 33230 5848
rect 31930 5782 31990 5788
rect 33074 5732 33194 5744
rect 33074 5660 33086 5732
rect 33182 5660 33194 5732
rect 33074 5648 33194 5660
rect 13294 5432 21650 5442
rect 13294 5346 13308 5432
rect 13404 5346 13908 5432
rect 14004 5346 14508 5432
rect 14604 5346 15108 5432
rect 15204 5346 15708 5432
rect 15804 5346 16308 5432
rect 16404 5346 16908 5432
rect 17004 5346 17508 5432
rect 17604 5346 18108 5432
rect 18204 5346 18708 5432
rect 18804 5346 19308 5432
rect 19404 5346 19908 5432
rect 20004 5346 20508 5432
rect 20604 5346 21108 5432
rect 21204 5346 21528 5432
rect 21624 5346 21650 5432
rect 13294 5332 21650 5346
rect 23810 5432 28808 5442
rect 23810 5346 23824 5432
rect 23920 5346 24424 5432
rect 24520 5346 25024 5432
rect 25120 5346 25624 5432
rect 25720 5346 26224 5432
rect 26320 5346 26824 5432
rect 26920 5346 27424 5432
rect 27520 5346 28024 5432
rect 28120 5346 28624 5432
rect 28720 5346 28808 5432
rect 29336 5376 33972 5476
rect 23810 5332 28808 5346
rect 13066 5172 13448 5182
rect 13066 4862 13448 4872
rect 21200 5172 21878 5182
rect 21200 4862 21878 4872
rect 23648 5172 24248 5182
rect 23648 4862 24248 4872
rect 28280 5172 28880 5182
rect 28280 4862 28880 4872
rect 8458 4290 9058 4300
rect 8458 3980 9058 3990
rect 18090 4290 18690 4300
rect 18090 3980 18690 3990
rect 23458 4290 24058 4300
rect 23458 3980 24058 3990
rect 33090 4290 33690 4300
rect 33090 3980 33690 3990
rect 9296 3816 17652 3830
rect 9296 3730 9310 3816
rect 9406 3730 9910 3816
rect 10006 3730 10510 3816
rect 10606 3730 11110 3816
rect 11206 3730 11710 3816
rect 11806 3730 12310 3816
rect 12406 3730 12910 3816
rect 13006 3730 13510 3816
rect 13606 3730 14110 3816
rect 14206 3730 14710 3816
rect 14806 3730 15310 3816
rect 15406 3730 15910 3816
rect 16006 3730 16510 3816
rect 16606 3730 17110 3816
rect 17206 3730 17530 3816
rect 17626 3730 17652 3816
rect 9296 3720 17652 3730
rect 24296 3816 32652 3830
rect 24296 3730 24310 3816
rect 24406 3730 24910 3816
rect 25006 3730 25510 3816
rect 25606 3730 26110 3816
rect 26206 3730 26710 3816
rect 26806 3730 27310 3816
rect 27406 3730 27910 3816
rect 28006 3730 28510 3816
rect 28606 3730 29110 3816
rect 29206 3730 29710 3816
rect 29806 3730 30310 3816
rect 30406 3730 30910 3816
rect 31006 3730 31510 3816
rect 31606 3730 32110 3816
rect 32206 3730 32530 3816
rect 32626 3730 32652 3816
rect 24296 3720 32652 3730
rect 10014 3158 10074 3164
rect 10470 3158 10530 3164
rect 10930 3158 10990 3164
rect 11386 3158 11446 3164
rect 11844 3158 11904 3164
rect 12308 3158 12368 3164
rect 12758 3158 12818 3164
rect 13214 3158 13274 3164
rect 13682 3158 13742 3164
rect 14140 3158 14200 3164
rect 14596 3158 14656 3164
rect 15052 3158 15112 3164
rect 15508 3158 15568 3164
rect 15964 3158 16024 3164
rect 16422 3158 16482 3164
rect 16882 3158 16942 3164
rect 25014 3158 25074 3164
rect 25470 3158 25530 3164
rect 25930 3158 25990 3164
rect 26386 3158 26446 3164
rect 26844 3158 26904 3164
rect 27308 3158 27368 3164
rect 27758 3158 27818 3164
rect 28214 3158 28274 3164
rect 28682 3158 28742 3164
rect 29140 3158 29200 3164
rect 29596 3158 29656 3164
rect 30052 3158 30112 3164
rect 30508 3158 30568 3164
rect 30964 3158 31024 3164
rect 31422 3158 31482 3164
rect 31882 3158 31942 3164
rect 10074 3098 10470 3158
rect 10530 3098 10930 3158
rect 10990 3098 11386 3158
rect 11446 3098 11844 3158
rect 11904 3098 12308 3158
rect 12368 3098 12758 3158
rect 12818 3098 13214 3158
rect 13274 3098 13682 3158
rect 13742 3098 14140 3158
rect 14200 3098 14596 3158
rect 14656 3098 15052 3158
rect 15112 3098 15508 3158
rect 15568 3098 15964 3158
rect 16024 3098 16422 3158
rect 16482 3098 16882 3158
rect 16942 3098 22942 3158
rect 23002 3098 25014 3158
rect 25074 3098 25470 3158
rect 25530 3098 25930 3158
rect 25990 3098 26386 3158
rect 26446 3098 26844 3158
rect 26904 3098 27308 3158
rect 27368 3098 27758 3158
rect 27818 3098 28214 3158
rect 28274 3098 28682 3158
rect 28742 3098 29140 3158
rect 29200 3098 29596 3158
rect 29656 3098 30052 3158
rect 30112 3098 30508 3158
rect 30568 3098 30964 3158
rect 31024 3098 31422 3158
rect 31482 3098 31882 3158
rect 10014 3092 10074 3098
rect 10470 3092 10530 3098
rect 10930 3092 10990 3098
rect 11386 3092 11446 3098
rect 11844 3092 11904 3098
rect 12308 3092 12368 3098
rect 12758 3092 12818 3098
rect 13214 3092 13274 3098
rect 13682 3092 13742 3098
rect 14140 3092 14200 3098
rect 14596 3092 14656 3098
rect 15052 3092 15112 3098
rect 15508 3092 15568 3098
rect 15964 3092 16024 3098
rect 16422 3092 16482 3098
rect 16882 3092 16942 3098
rect 25014 3092 25074 3098
rect 25470 3092 25530 3098
rect 25930 3092 25990 3098
rect 26386 3092 26446 3098
rect 26844 3092 26904 3098
rect 27308 3092 27368 3098
rect 27758 3092 27818 3098
rect 28214 3092 28274 3098
rect 28682 3092 28742 3098
rect 29140 3092 29200 3098
rect 29596 3092 29656 3098
rect 30052 3092 30112 3098
rect 30508 3092 30568 3098
rect 30964 3092 31024 3098
rect 31422 3092 31482 3098
rect 31882 3092 31942 3098
rect 10010 1184 10070 1190
rect 10466 1184 10526 1190
rect 10926 1184 10986 1190
rect 11382 1184 11442 1190
rect 11840 1184 11900 1190
rect 12304 1184 12364 1190
rect 12758 1184 12818 1190
rect 13216 1184 13276 1190
rect 10070 1124 10466 1184
rect 10526 1124 10926 1184
rect 10986 1124 11382 1184
rect 11442 1124 11840 1184
rect 11900 1124 12304 1184
rect 12364 1124 12758 1184
rect 12818 1124 13216 1184
rect 13444 1136 13450 1196
rect 13510 1136 13516 1196
rect 13676 1184 13736 1190
rect 14132 1184 14192 1190
rect 14592 1184 14652 1190
rect 15048 1184 15108 1190
rect 15504 1184 15564 1190
rect 15960 1184 16020 1190
rect 16418 1184 16478 1190
rect 16878 1184 16938 1190
rect 10010 1118 10070 1124
rect 10466 1118 10526 1124
rect 10926 1118 10986 1124
rect 11382 1118 11442 1124
rect 11840 1118 11900 1124
rect 12304 1118 12364 1124
rect 12758 1118 12818 1124
rect 13216 1118 13276 1124
rect 9224 598 9284 604
rect 13450 598 13510 1136
rect 13736 1124 14132 1184
rect 14192 1124 14592 1184
rect 14652 1124 15048 1184
rect 15108 1124 15504 1184
rect 15564 1124 15960 1184
rect 16020 1124 16418 1184
rect 16478 1124 16878 1184
rect 13676 1118 13736 1124
rect 14132 1118 14192 1124
rect 14592 1118 14652 1124
rect 15048 1118 15108 1124
rect 15504 1118 15564 1124
rect 15960 1118 16020 1124
rect 16418 1118 16478 1124
rect 16878 1118 16938 1124
rect 25010 1184 25070 1190
rect 25466 1184 25526 1190
rect 25926 1184 25986 1190
rect 26382 1184 26442 1190
rect 26840 1184 26900 1190
rect 27304 1184 27364 1190
rect 27758 1184 27818 1190
rect 28216 1184 28276 1190
rect 25070 1124 25466 1184
rect 25526 1124 25926 1184
rect 25986 1124 26382 1184
rect 26442 1124 26840 1184
rect 26900 1124 27304 1184
rect 27364 1124 27758 1184
rect 27818 1124 28216 1184
rect 28444 1136 28450 1196
rect 28510 1136 28516 1196
rect 28676 1184 28736 1190
rect 29132 1184 29192 1190
rect 29592 1184 29652 1190
rect 30048 1184 30108 1190
rect 30504 1184 30564 1190
rect 30960 1184 31020 1190
rect 31418 1184 31478 1190
rect 31878 1184 31938 1190
rect 25010 1118 25070 1124
rect 25466 1118 25526 1124
rect 25926 1118 25986 1124
rect 26382 1118 26442 1124
rect 26840 1118 26900 1124
rect 27304 1118 27364 1124
rect 27758 1118 27818 1124
rect 28216 1118 28276 1124
rect 22768 760 22828 766
rect 9284 538 13510 598
rect 13714 700 22768 760
rect 9224 532 9284 538
rect 12658 496 12718 502
rect 13714 496 13774 700
rect 22768 694 22828 700
rect 24224 598 24284 604
rect 28450 598 28510 1136
rect 28736 1124 29132 1184
rect 29192 1124 29592 1184
rect 29652 1124 30048 1184
rect 30108 1124 30504 1184
rect 30564 1124 30960 1184
rect 31020 1124 31418 1184
rect 31478 1124 31878 1184
rect 28676 1118 28736 1124
rect 29132 1118 29192 1124
rect 29592 1118 29652 1124
rect 30048 1118 30108 1124
rect 30504 1118 30564 1124
rect 30960 1118 31020 1124
rect 31418 1118 31478 1124
rect 31878 1118 31938 1124
rect 24284 538 28510 598
rect 24224 532 24284 538
rect 12718 436 13774 496
rect 12658 430 12718 436
rect 9442 -1140 9448 -1080
rect 9508 -1140 9514 -1080
rect 9904 -1140 9910 -1080
rect 9970 -1140 9976 -1080
rect 10358 -1136 10364 -1076
rect 10424 -1136 10430 -1076
rect 10820 -1136 10826 -1076
rect 10886 -1136 10892 -1076
rect 9448 -1534 9508 -1140
rect 9910 -1534 9970 -1140
rect 10364 -1534 10424 -1136
rect 10826 -1534 10886 -1136
rect 11274 -1142 11280 -1082
rect 11340 -1142 11346 -1082
rect 11724 -1136 11730 -1076
rect 11790 -1136 11796 -1076
rect 12190 -1136 12196 -1076
rect 12256 -1136 12262 -1076
rect 11280 -1534 11340 -1142
rect 11730 -1534 11790 -1136
rect 12196 -1534 12256 -1136
rect 12646 -1140 12652 -1080
rect 12712 -1140 12718 -1080
rect 14444 -1140 14450 -1080
rect 14510 -1140 14516 -1080
rect 14906 -1132 14912 -1072
rect 14972 -1132 14978 -1072
rect 12652 -1534 12712 -1140
rect 9446 -1594 12712 -1534
rect 9448 -2016 9508 -1594
rect 9910 -2010 9970 -1594
rect 9910 -2076 9970 -2070
rect 10364 -2016 10424 -1594
rect 10826 -2010 10886 -1594
rect 10826 -2076 10886 -2070
rect 11280 -2010 11340 -1594
rect 11280 -2076 11340 -2070
rect 11730 -2010 11790 -1594
rect 11730 -2076 11790 -2070
rect 12196 -2016 12256 -1594
rect 12652 -2010 12712 -1594
rect 12886 -1202 12946 -1196
rect 12886 -1540 12946 -1262
rect 14450 -1540 14510 -1140
rect 14912 -1540 14972 -1132
rect 15360 -1138 15366 -1078
rect 15426 -1138 15432 -1078
rect 15822 -1138 15828 -1078
rect 15888 -1138 15894 -1078
rect 16276 -1138 16282 -1078
rect 16342 -1138 16348 -1078
rect 16726 -1132 16732 -1072
rect 16792 -1132 16798 -1072
rect 15366 -1540 15426 -1138
rect 15828 -1540 15888 -1138
rect 16282 -1540 16342 -1138
rect 16732 -1540 16792 -1132
rect 17192 -1138 17198 -1078
rect 17258 -1138 17264 -1078
rect 17648 -1138 17654 -1078
rect 17714 -1138 17720 -1078
rect 17198 -1540 17258 -1138
rect 17654 -1540 17714 -1138
rect 24442 -1140 24448 -1080
rect 24508 -1140 24514 -1080
rect 24904 -1140 24910 -1080
rect 24970 -1140 24976 -1080
rect 25358 -1136 25364 -1076
rect 25424 -1136 25430 -1076
rect 25820 -1136 25826 -1076
rect 25886 -1136 25892 -1076
rect 17880 -1268 17886 -1208
rect 17946 -1268 17952 -1208
rect 12886 -1600 17714 -1540
rect 12886 -1882 12946 -1600
rect 12880 -1942 12886 -1882
rect 12946 -1942 12952 -1882
rect 12652 -2076 12712 -2070
rect 14450 -2010 14510 -1600
rect 14450 -2076 14510 -2070
rect 14912 -2012 14972 -1600
rect 9448 -2082 9508 -2076
rect 10364 -2082 10424 -2076
rect 12196 -2082 12256 -2076
rect 14912 -2078 14972 -2072
rect 15366 -2012 15426 -1600
rect 15366 -2078 15426 -2072
rect 15828 -2012 15888 -1600
rect 15828 -2078 15888 -2072
rect 16282 -2012 16342 -1600
rect 16732 -2006 16792 -1600
rect 16732 -2072 16792 -2066
rect 17198 -2010 17258 -1600
rect 16282 -2078 16342 -2072
rect 17198 -2076 17258 -2070
rect 17654 -2010 17714 -1600
rect 17886 -1544 17946 -1268
rect 23150 -1534 23210 -1525
rect 24448 -1534 24508 -1140
rect 24910 -1534 24970 -1140
rect 25364 -1534 25424 -1136
rect 25826 -1534 25886 -1136
rect 26274 -1142 26280 -1082
rect 26340 -1142 26346 -1082
rect 26724 -1136 26730 -1076
rect 26790 -1136 26796 -1076
rect 27190 -1136 27196 -1076
rect 27256 -1136 27262 -1076
rect 26280 -1534 26340 -1142
rect 26730 -1534 26790 -1136
rect 27196 -1534 27256 -1136
rect 27646 -1140 27652 -1080
rect 27712 -1140 27718 -1080
rect 29444 -1140 29450 -1080
rect 29510 -1140 29516 -1080
rect 29906 -1132 29912 -1072
rect 29972 -1132 29978 -1072
rect 27652 -1534 27712 -1140
rect 17886 -1604 18972 -1544
rect 23210 -1594 27712 -1534
rect 23150 -1603 23210 -1594
rect 17886 -1870 17946 -1604
rect 18872 -1733 18972 -1604
rect 18868 -1823 18877 -1733
rect 18967 -1823 18976 -1733
rect 18872 -1828 18972 -1823
rect 17886 -1936 17946 -1930
rect 17654 -2076 17714 -2070
rect 24448 -2016 24508 -1594
rect 24910 -2010 24970 -1594
rect 24910 -2076 24970 -2070
rect 25364 -2016 25424 -1594
rect 25826 -2010 25886 -1594
rect 25826 -2076 25886 -2070
rect 26280 -2010 26340 -1594
rect 26280 -2076 26340 -2070
rect 26730 -2010 26790 -1594
rect 26730 -2076 26790 -2070
rect 27196 -2016 27256 -1594
rect 27652 -2010 27712 -1594
rect 27886 -1202 27946 -1196
rect 27886 -1540 27946 -1262
rect 29450 -1540 29510 -1140
rect 29912 -1540 29972 -1132
rect 30360 -1138 30366 -1078
rect 30426 -1138 30432 -1078
rect 30822 -1138 30828 -1078
rect 30888 -1138 30894 -1078
rect 31276 -1138 31282 -1078
rect 31342 -1138 31348 -1078
rect 31726 -1132 31732 -1072
rect 31792 -1132 31798 -1072
rect 30366 -1540 30426 -1138
rect 30828 -1540 30888 -1138
rect 31282 -1540 31342 -1138
rect 31732 -1540 31792 -1132
rect 32192 -1138 32198 -1078
rect 32258 -1138 32264 -1078
rect 32648 -1138 32654 -1078
rect 32714 -1138 32720 -1078
rect 32198 -1540 32258 -1138
rect 32654 -1540 32714 -1138
rect 32880 -1268 32886 -1208
rect 32946 -1268 32952 -1208
rect 27886 -1600 32714 -1540
rect 27886 -1882 27946 -1600
rect 27880 -1942 27886 -1882
rect 27946 -1942 27952 -1882
rect 27652 -2076 27712 -2070
rect 29450 -2010 29510 -1600
rect 29450 -2076 29510 -2070
rect 29912 -2012 29972 -1600
rect 24448 -2082 24508 -2076
rect 25364 -2082 25424 -2076
rect 27196 -2082 27256 -2076
rect 29912 -2078 29972 -2072
rect 30366 -2012 30426 -1600
rect 30366 -2078 30426 -2072
rect 30828 -2012 30888 -1600
rect 30828 -2078 30888 -2072
rect 31282 -2012 31342 -1600
rect 31732 -2006 31792 -1600
rect 31732 -2072 31792 -2066
rect 32198 -2010 32258 -1600
rect 31282 -2078 31342 -2072
rect 32198 -2076 32258 -2070
rect 32654 -2010 32714 -1600
rect 32886 -1544 32946 -1268
rect 33872 -1544 33972 5376
rect 32886 -1604 33972 -1544
rect 32886 -1870 32946 -1604
rect 33872 -1733 33972 -1604
rect 33868 -1823 33877 -1733
rect 33967 -1823 33976 -1733
rect 33872 -1828 33972 -1823
rect 32886 -1936 32946 -1930
rect 32654 -2076 32714 -2070
rect 12650 -3226 12710 -3220
rect 23080 -3226 23140 -3220
rect 12710 -3286 23080 -3226
rect 23140 -3286 24448 -3226
rect 24508 -3286 24514 -3226
rect 12650 -3292 12710 -3286
rect 23080 -3292 23140 -3286
rect 8694 -3478 18464 -3450
rect 8694 -3564 8744 -3478
rect 8840 -3564 9324 -3478
rect 9420 -3564 9924 -3478
rect 10020 -3564 10524 -3478
rect 10620 -3564 11124 -3478
rect 11220 -3564 11724 -3478
rect 11820 -3564 12324 -3478
rect 12420 -3564 12924 -3478
rect 13020 -3564 13524 -3478
rect 13620 -3564 14124 -3478
rect 14220 -3564 14724 -3478
rect 14820 -3564 15324 -3478
rect 15420 -3564 15924 -3478
rect 16020 -3564 16524 -3478
rect 16620 -3564 17124 -3478
rect 17220 -3564 17724 -3478
rect 17820 -3564 18324 -3478
rect 18420 -3564 18464 -3478
rect 8694 -3594 18464 -3564
rect 23694 -3478 33464 -3450
rect 23694 -3564 23744 -3478
rect 23840 -3564 24324 -3478
rect 24420 -3564 24924 -3478
rect 25020 -3564 25524 -3478
rect 25620 -3564 26124 -3478
rect 26220 -3564 26724 -3478
rect 26820 -3564 27324 -3478
rect 27420 -3564 27924 -3478
rect 28020 -3564 28524 -3478
rect 28620 -3564 29124 -3478
rect 29220 -3564 29724 -3478
rect 29820 -3564 30324 -3478
rect 30420 -3564 30924 -3478
rect 31020 -3564 31524 -3478
rect 31620 -3564 32124 -3478
rect 32220 -3564 32724 -3478
rect 32820 -3564 33324 -3478
rect 33420 -3564 33464 -3478
rect 23694 -3594 33464 -3564
rect 8458 -3742 9058 -3732
rect 8458 -4052 9058 -4042
rect 18090 -3742 18690 -3732
rect 18090 -4052 18690 -4042
rect 23458 -3742 24058 -3732
rect 23458 -4052 24058 -4042
rect 33090 -3742 33690 -3732
rect 33090 -4052 33690 -4042
rect 12412 -4714 13012 -4704
rect 12412 -5024 13012 -5014
rect 22044 -4714 22644 -4704
rect 22044 -5024 22644 -5014
rect 27412 -4714 28012 -4704
rect 27412 -5024 28012 -5014
rect 37044 -4714 37644 -4704
rect 37044 -5024 37644 -5014
rect 12638 -5192 22408 -5162
rect 12638 -5278 12682 -5192
rect 12778 -5278 13282 -5192
rect 13378 -5278 13882 -5192
rect 13978 -5278 14482 -5192
rect 14578 -5278 15082 -5192
rect 15178 -5278 15682 -5192
rect 15778 -5278 16282 -5192
rect 16378 -5278 16882 -5192
rect 16978 -5278 17482 -5192
rect 17578 -5278 18082 -5192
rect 18178 -5278 18682 -5192
rect 18778 -5278 19282 -5192
rect 19378 -5278 19882 -5192
rect 19978 -5278 20482 -5192
rect 20578 -5278 21082 -5192
rect 21178 -5278 21682 -5192
rect 21778 -5278 22262 -5192
rect 22358 -5278 22408 -5192
rect 12638 -5306 22408 -5278
rect 27638 -5192 37408 -5162
rect 27638 -5278 27682 -5192
rect 27778 -5278 28282 -5192
rect 28378 -5278 28882 -5192
rect 28978 -5278 29482 -5192
rect 29578 -5278 30082 -5192
rect 30178 -5278 30682 -5192
rect 30778 -5278 31282 -5192
rect 31378 -5278 31882 -5192
rect 31978 -5278 32482 -5192
rect 32578 -5278 33082 -5192
rect 33178 -5278 33682 -5192
rect 33778 -5278 34282 -5192
rect 34378 -5278 34882 -5192
rect 34978 -5278 35482 -5192
rect 35578 -5278 36082 -5192
rect 36178 -5278 36682 -5192
rect 36778 -5278 37262 -5192
rect 37358 -5278 37408 -5192
rect 27638 -5306 37408 -5278
rect 21596 -5470 21656 -5464
rect 21656 -5530 23080 -5470
rect 23140 -5530 33390 -5470
rect 33450 -5530 33456 -5470
rect 21596 -5536 21656 -5530
rect 13388 -6686 13448 -6680
rect 13156 -6826 13216 -6820
rect 8164 -6933 8224 -6928
rect 12130 -6933 12230 -6928
rect 8134 -7023 8143 -6933
rect 8233 -7023 8242 -6933
rect 12126 -7023 12135 -6933
rect 12225 -7023 12234 -6933
rect 8164 -19534 8224 -7023
rect 12130 -7152 12230 -7023
rect 13156 -7152 13216 -6886
rect 12130 -7212 13216 -7152
rect 13156 -7488 13216 -7212
rect 13388 -7156 13448 -6746
rect 13844 -6686 13904 -6680
rect 14760 -6684 14820 -6678
rect 13844 -7156 13904 -6746
rect 14310 -6690 14370 -6684
rect 14310 -7156 14370 -6750
rect 14760 -7156 14820 -6744
rect 15214 -6684 15274 -6678
rect 15214 -7156 15274 -6744
rect 15676 -6684 15736 -6678
rect 15676 -7156 15736 -6744
rect 16130 -6684 16190 -6678
rect 18846 -6680 18906 -6674
rect 20678 -6680 20738 -6674
rect 21594 -6680 21654 -6674
rect 16130 -7156 16190 -6744
rect 16592 -6686 16652 -6680
rect 16592 -7156 16652 -6746
rect 18390 -6686 18450 -6680
rect 18150 -6874 18156 -6814
rect 18216 -6874 18222 -6814
rect 18156 -7156 18216 -6874
rect 13388 -7216 18216 -7156
rect 13150 -7548 13156 -7488
rect 13216 -7548 13222 -7488
rect 13388 -7618 13448 -7216
rect 13844 -7618 13904 -7216
rect 13382 -7678 13388 -7618
rect 13448 -7678 13454 -7618
rect 13838 -7678 13844 -7618
rect 13904 -7678 13910 -7618
rect 14310 -7624 14370 -7216
rect 14760 -7618 14820 -7216
rect 15214 -7618 15274 -7216
rect 15676 -7618 15736 -7216
rect 14304 -7684 14310 -7624
rect 14370 -7684 14376 -7624
rect 14754 -7678 14760 -7618
rect 14820 -7678 14826 -7618
rect 15208 -7678 15214 -7618
rect 15274 -7678 15280 -7618
rect 15670 -7678 15676 -7618
rect 15736 -7678 15742 -7618
rect 16130 -7624 16190 -7216
rect 16592 -7616 16652 -7216
rect 18156 -7494 18216 -7216
rect 18156 -7560 18216 -7554
rect 18390 -7162 18450 -6746
rect 18846 -7162 18906 -6740
rect 19312 -6686 19372 -6680
rect 19312 -7162 19372 -6746
rect 19762 -6686 19822 -6680
rect 19762 -7162 19822 -6746
rect 20216 -6686 20276 -6680
rect 20216 -7162 20276 -6746
rect 20678 -7162 20738 -6740
rect 21132 -6686 21192 -6680
rect 21132 -7162 21192 -6746
rect 21594 -7162 21654 -6740
rect 28388 -6686 28448 -6680
rect 28156 -6826 28216 -6820
rect 27130 -6933 27230 -6928
rect 27126 -7023 27135 -6933
rect 27225 -7023 27234 -6933
rect 27130 -7152 27230 -7023
rect 28156 -7152 28216 -6886
rect 22834 -7162 22894 -7153
rect 18390 -7222 22834 -7162
rect 27130 -7212 28216 -7152
rect 18390 -7616 18450 -7222
rect 16124 -7684 16130 -7624
rect 16190 -7684 16196 -7624
rect 16586 -7676 16592 -7616
rect 16652 -7676 16658 -7616
rect 18384 -7676 18390 -7616
rect 18450 -7676 18456 -7616
rect 18846 -7620 18906 -7222
rect 19312 -7620 19372 -7222
rect 19762 -7614 19822 -7222
rect 18840 -7680 18846 -7620
rect 18906 -7680 18912 -7620
rect 19306 -7680 19312 -7620
rect 19372 -7680 19378 -7620
rect 19756 -7674 19762 -7614
rect 19822 -7674 19828 -7614
rect 20216 -7620 20276 -7222
rect 20678 -7620 20738 -7222
rect 21132 -7616 21192 -7222
rect 21594 -7616 21654 -7222
rect 22834 -7231 22894 -7222
rect 28156 -7488 28216 -7212
rect 28388 -7156 28448 -6746
rect 28844 -6686 28904 -6680
rect 29760 -6684 29820 -6678
rect 28844 -7156 28904 -6746
rect 29310 -6690 29370 -6684
rect 29310 -7156 29370 -6750
rect 29760 -7156 29820 -6744
rect 30214 -6684 30274 -6678
rect 30214 -7156 30274 -6744
rect 30676 -6684 30736 -6678
rect 30676 -7156 30736 -6744
rect 31130 -6684 31190 -6678
rect 33846 -6680 33906 -6674
rect 35678 -6680 35738 -6674
rect 36594 -6680 36654 -6674
rect 31130 -7156 31190 -6744
rect 31592 -6686 31652 -6680
rect 31592 -7156 31652 -6746
rect 33390 -6686 33450 -6680
rect 33150 -6874 33156 -6814
rect 33216 -6874 33222 -6814
rect 33156 -7156 33216 -6874
rect 28388 -7216 33216 -7156
rect 28150 -7548 28156 -7488
rect 28216 -7548 28222 -7488
rect 20210 -7680 20216 -7620
rect 20276 -7680 20282 -7620
rect 20672 -7680 20678 -7620
rect 20738 -7680 20744 -7620
rect 21126 -7676 21132 -7616
rect 21192 -7676 21198 -7616
rect 21588 -7676 21594 -7616
rect 21654 -7676 21660 -7616
rect 28388 -7618 28448 -7216
rect 28844 -7618 28904 -7216
rect 28382 -7678 28388 -7618
rect 28448 -7678 28454 -7618
rect 28838 -7678 28844 -7618
rect 28904 -7678 28910 -7618
rect 29310 -7624 29370 -7216
rect 29760 -7618 29820 -7216
rect 30214 -7618 30274 -7216
rect 30676 -7618 30736 -7216
rect 29304 -7684 29310 -7624
rect 29370 -7684 29376 -7624
rect 29754 -7678 29760 -7618
rect 29820 -7678 29826 -7618
rect 30208 -7678 30214 -7618
rect 30274 -7678 30280 -7618
rect 30670 -7678 30676 -7618
rect 30736 -7678 30742 -7618
rect 31130 -7624 31190 -7216
rect 31592 -7616 31652 -7216
rect 33156 -7494 33216 -7216
rect 33156 -7560 33216 -7554
rect 33390 -7162 33450 -6746
rect 33846 -7162 33906 -6740
rect 34312 -6686 34372 -6680
rect 34312 -7162 34372 -6746
rect 34762 -6686 34822 -6680
rect 34762 -7162 34822 -6746
rect 35216 -6686 35276 -6680
rect 35216 -7162 35276 -6746
rect 35678 -7162 35738 -6740
rect 36132 -6686 36192 -6680
rect 36132 -7162 36192 -6746
rect 36594 -7162 36654 -6740
rect 33390 -7222 37914 -7162
rect 33390 -7616 33450 -7222
rect 31124 -7684 31130 -7624
rect 31190 -7684 31196 -7624
rect 31586 -7676 31592 -7616
rect 31652 -7676 31658 -7616
rect 33384 -7676 33390 -7616
rect 33450 -7676 33456 -7616
rect 33846 -7620 33906 -7222
rect 34312 -7620 34372 -7222
rect 34762 -7614 34822 -7222
rect 33840 -7680 33846 -7620
rect 33906 -7680 33912 -7620
rect 34306 -7680 34312 -7620
rect 34372 -7680 34378 -7620
rect 34756 -7674 34762 -7614
rect 34822 -7674 34828 -7614
rect 35216 -7620 35276 -7222
rect 35678 -7620 35738 -7222
rect 36132 -7616 36192 -7222
rect 36594 -7616 36654 -7222
rect 35210 -7680 35216 -7620
rect 35276 -7680 35282 -7620
rect 35672 -7680 35678 -7620
rect 35738 -7680 35744 -7620
rect 36126 -7676 36132 -7616
rect 36192 -7676 36198 -7616
rect 36588 -7676 36594 -7616
rect 36654 -7676 36660 -7616
rect 21818 -9294 21878 -9288
rect 36818 -9294 36878 -9288
rect 17592 -9354 21818 -9294
rect 14164 -9880 14224 -9874
rect 14624 -9880 14684 -9874
rect 15082 -9880 15142 -9874
rect 15538 -9880 15598 -9874
rect 15994 -9880 16054 -9874
rect 16450 -9880 16510 -9874
rect 16910 -9880 16970 -9874
rect 17366 -9880 17426 -9874
rect 14224 -9940 14624 -9880
rect 14684 -9940 15082 -9880
rect 15142 -9940 15538 -9880
rect 15598 -9940 15994 -9880
rect 16054 -9940 16450 -9880
rect 16510 -9940 16910 -9880
rect 16970 -9940 17366 -9880
rect 17592 -9892 17652 -9354
rect 21818 -9360 21878 -9354
rect 32592 -9354 36818 -9294
rect 17826 -9880 17886 -9874
rect 18284 -9880 18344 -9874
rect 18738 -9880 18798 -9874
rect 19202 -9880 19262 -9874
rect 19660 -9880 19720 -9874
rect 20116 -9880 20176 -9874
rect 20576 -9880 20636 -9874
rect 21032 -9880 21092 -9874
rect 29164 -9880 29224 -9874
rect 29624 -9880 29684 -9874
rect 30082 -9880 30142 -9874
rect 30538 -9880 30598 -9874
rect 30994 -9880 31054 -9874
rect 31450 -9880 31510 -9874
rect 31910 -9880 31970 -9874
rect 32366 -9880 32426 -9874
rect 14164 -9946 14224 -9940
rect 14624 -9946 14684 -9940
rect 15082 -9946 15142 -9940
rect 15538 -9946 15598 -9940
rect 15994 -9946 16054 -9940
rect 16450 -9946 16510 -9940
rect 16910 -9946 16970 -9940
rect 17366 -9946 17426 -9940
rect 17586 -9952 17592 -9892
rect 17652 -9952 17658 -9892
rect 17886 -9940 18284 -9880
rect 18344 -9940 18738 -9880
rect 18798 -9940 19202 -9880
rect 19262 -9940 19660 -9880
rect 19720 -9940 20116 -9880
rect 20176 -9940 20576 -9880
rect 20636 -9940 21032 -9880
rect 21092 -9940 22940 -9880
rect 23000 -9940 29164 -9880
rect 29224 -9940 29624 -9880
rect 29684 -9940 30082 -9880
rect 30142 -9940 30538 -9880
rect 30598 -9940 30994 -9880
rect 31054 -9940 31450 -9880
rect 31510 -9940 31910 -9880
rect 31970 -9940 32366 -9880
rect 32592 -9892 32652 -9354
rect 36818 -9360 36878 -9354
rect 32826 -9880 32886 -9874
rect 33284 -9880 33344 -9874
rect 33738 -9880 33798 -9874
rect 34202 -9880 34262 -9874
rect 34660 -9880 34720 -9874
rect 35116 -9880 35176 -9874
rect 35576 -9880 35636 -9874
rect 36032 -9880 36092 -9874
rect 17826 -9946 17886 -9940
rect 18284 -9946 18344 -9940
rect 18738 -9946 18798 -9940
rect 19202 -9946 19262 -9940
rect 19660 -9946 19720 -9940
rect 20116 -9946 20176 -9940
rect 20576 -9946 20636 -9940
rect 21032 -9946 21092 -9940
rect 29164 -9946 29224 -9940
rect 29624 -9946 29684 -9940
rect 30082 -9946 30142 -9940
rect 30538 -9946 30598 -9940
rect 30994 -9946 31054 -9940
rect 31450 -9946 31510 -9940
rect 31910 -9946 31970 -9940
rect 32366 -9946 32426 -9940
rect 32586 -9952 32592 -9892
rect 32652 -9952 32658 -9892
rect 32886 -9940 33284 -9880
rect 33344 -9940 33738 -9880
rect 33798 -9940 34202 -9880
rect 34262 -9940 34660 -9880
rect 34720 -9940 35116 -9880
rect 35176 -9940 35576 -9880
rect 35636 -9940 36032 -9880
rect 32826 -9946 32886 -9940
rect 33284 -9946 33344 -9940
rect 33738 -9946 33798 -9940
rect 34202 -9946 34262 -9940
rect 34660 -9946 34720 -9940
rect 35116 -9946 35176 -9940
rect 35576 -9946 35636 -9940
rect 36032 -9946 36092 -9940
rect 14160 -11854 14220 -11848
rect 14620 -11854 14680 -11848
rect 15078 -11854 15138 -11848
rect 15534 -11854 15594 -11848
rect 15990 -11854 16050 -11848
rect 16446 -11854 16506 -11848
rect 16902 -11854 16962 -11848
rect 17360 -11854 17420 -11848
rect 17828 -11854 17888 -11848
rect 18284 -11854 18344 -11848
rect 18734 -11854 18794 -11848
rect 19198 -11854 19258 -11848
rect 19656 -11854 19716 -11848
rect 20112 -11854 20172 -11848
rect 20572 -11854 20632 -11848
rect 21028 -11854 21088 -11848
rect 14220 -11914 14620 -11854
rect 14680 -11914 15078 -11854
rect 15138 -11914 15534 -11854
rect 15594 -11914 15990 -11854
rect 16050 -11914 16446 -11854
rect 16506 -11914 16902 -11854
rect 16962 -11914 17360 -11854
rect 17420 -11914 17828 -11854
rect 17888 -11914 18284 -11854
rect 18344 -11914 18734 -11854
rect 18794 -11914 19198 -11854
rect 19258 -11914 19656 -11854
rect 19716 -11914 20112 -11854
rect 20172 -11914 20572 -11854
rect 20632 -11914 21028 -11854
rect 14160 -11920 14220 -11914
rect 14620 -11920 14680 -11914
rect 15078 -11920 15138 -11914
rect 15534 -11920 15594 -11914
rect 15990 -11920 16050 -11914
rect 16446 -11920 16506 -11914
rect 16902 -11920 16962 -11914
rect 17360 -11920 17420 -11914
rect 17828 -11920 17888 -11914
rect 18284 -11920 18344 -11914
rect 18734 -11920 18794 -11914
rect 19198 -11920 19258 -11914
rect 19656 -11920 19716 -11914
rect 20112 -11920 20172 -11914
rect 20572 -11920 20632 -11914
rect 21028 -11920 21088 -11914
rect 29160 -11854 29220 -11848
rect 29620 -11854 29680 -11848
rect 30078 -11854 30138 -11848
rect 30534 -11854 30594 -11848
rect 30990 -11854 31050 -11848
rect 31446 -11854 31506 -11848
rect 31902 -11854 31962 -11848
rect 32360 -11854 32420 -11848
rect 32828 -11854 32888 -11848
rect 33284 -11854 33344 -11848
rect 33734 -11854 33794 -11848
rect 34198 -11854 34258 -11848
rect 34656 -11854 34716 -11848
rect 35112 -11854 35172 -11848
rect 35572 -11854 35632 -11848
rect 36028 -11854 36088 -11848
rect 29220 -11914 29620 -11854
rect 29680 -11914 30078 -11854
rect 30138 -11914 30534 -11854
rect 30594 -11914 30990 -11854
rect 31050 -11914 31446 -11854
rect 31506 -11914 31902 -11854
rect 31962 -11914 32360 -11854
rect 32420 -11914 32828 -11854
rect 32888 -11914 33284 -11854
rect 33344 -11914 33734 -11854
rect 33794 -11914 34198 -11854
rect 34258 -11914 34656 -11854
rect 34716 -11914 35112 -11854
rect 35172 -11914 35572 -11854
rect 35632 -11914 36028 -11854
rect 29160 -11920 29220 -11914
rect 29620 -11920 29680 -11914
rect 30078 -11920 30138 -11914
rect 30534 -11920 30594 -11914
rect 30990 -11920 31050 -11914
rect 31446 -11920 31506 -11914
rect 31902 -11920 31962 -11914
rect 32360 -11920 32420 -11914
rect 32828 -11920 32888 -11914
rect 33284 -11920 33344 -11914
rect 33734 -11920 33794 -11914
rect 34198 -11920 34258 -11914
rect 34656 -11920 34716 -11914
rect 35112 -11920 35172 -11914
rect 35572 -11920 35632 -11914
rect 36028 -11920 36088 -11914
rect 13450 -12486 21806 -12476
rect 13450 -12572 13476 -12486
rect 13572 -12572 13896 -12486
rect 13992 -12572 14496 -12486
rect 14592 -12572 15096 -12486
rect 15192 -12572 15696 -12486
rect 15792 -12572 16296 -12486
rect 16392 -12572 16896 -12486
rect 16992 -12572 17496 -12486
rect 17592 -12572 18096 -12486
rect 18192 -12572 18696 -12486
rect 18792 -12572 19296 -12486
rect 19392 -12572 19896 -12486
rect 19992 -12572 20496 -12486
rect 20592 -12572 21096 -12486
rect 21192 -12572 21696 -12486
rect 21792 -12572 21806 -12486
rect 13450 -12586 21806 -12572
rect 28450 -12486 36806 -12476
rect 28450 -12572 28476 -12486
rect 28572 -12572 28896 -12486
rect 28992 -12572 29496 -12486
rect 29592 -12572 30096 -12486
rect 30192 -12572 30696 -12486
rect 30792 -12572 31296 -12486
rect 31392 -12572 31896 -12486
rect 31992 -12572 32496 -12486
rect 32592 -12572 33096 -12486
rect 33192 -12572 33696 -12486
rect 33792 -12572 34296 -12486
rect 34392 -12572 34896 -12486
rect 34992 -12572 35496 -12486
rect 35592 -12572 36096 -12486
rect 36192 -12572 36696 -12486
rect 36792 -12572 36806 -12486
rect 28450 -12586 36806 -12572
rect 12412 -12746 13012 -12736
rect 12412 -13056 13012 -13046
rect 22044 -12746 22644 -12736
rect 22044 -13056 22644 -13046
rect 27412 -12746 28012 -12736
rect 27412 -13056 28012 -13046
rect 37044 -12746 37644 -12736
rect 37044 -13056 37644 -13046
rect 8458 -13710 9058 -13700
rect 8458 -14020 9058 -14010
rect 18090 -13710 18690 -13700
rect 18090 -14020 18690 -14010
rect 23458 -13710 24058 -13700
rect 23458 -14020 24058 -14010
rect 33090 -13710 33690 -13700
rect 33090 -14020 33690 -14010
rect 9296 -14184 17652 -14170
rect 9296 -14270 9310 -14184
rect 9406 -14270 9910 -14184
rect 10006 -14270 10510 -14184
rect 10606 -14270 11110 -14184
rect 11206 -14270 11710 -14184
rect 11806 -14270 12310 -14184
rect 12406 -14270 12910 -14184
rect 13006 -14270 13510 -14184
rect 13606 -14270 14110 -14184
rect 14206 -14270 14710 -14184
rect 14806 -14270 15310 -14184
rect 15406 -14270 15910 -14184
rect 16006 -14270 16510 -14184
rect 16606 -14270 17110 -14184
rect 17206 -14270 17530 -14184
rect 17626 -14270 17652 -14184
rect 9296 -14280 17652 -14270
rect 24296 -14184 32652 -14170
rect 24296 -14270 24310 -14184
rect 24406 -14270 24910 -14184
rect 25006 -14270 25510 -14184
rect 25606 -14270 26110 -14184
rect 26206 -14270 26710 -14184
rect 26806 -14270 27310 -14184
rect 27406 -14270 27910 -14184
rect 28006 -14270 28510 -14184
rect 28606 -14270 29110 -14184
rect 29206 -14270 29710 -14184
rect 29806 -14270 30310 -14184
rect 30406 -14270 30910 -14184
rect 31006 -14270 31510 -14184
rect 31606 -14270 32110 -14184
rect 32206 -14270 32530 -14184
rect 32626 -14270 32652 -14184
rect 24296 -14280 32652 -14270
rect 10014 -14842 10074 -14836
rect 10470 -14842 10530 -14836
rect 10930 -14842 10990 -14836
rect 11386 -14842 11446 -14836
rect 11844 -14842 11904 -14836
rect 12308 -14842 12368 -14836
rect 12758 -14842 12818 -14836
rect 13214 -14842 13274 -14836
rect 13682 -14842 13742 -14836
rect 14140 -14842 14200 -14836
rect 14596 -14842 14656 -14836
rect 15052 -14842 15112 -14836
rect 15508 -14842 15568 -14836
rect 15964 -14842 16024 -14836
rect 16422 -14842 16482 -14836
rect 16882 -14842 16942 -14836
rect 10074 -14902 10470 -14842
rect 10530 -14902 10930 -14842
rect 10990 -14902 11386 -14842
rect 11446 -14902 11844 -14842
rect 11904 -14902 12308 -14842
rect 12368 -14902 12758 -14842
rect 12818 -14902 13214 -14842
rect 13274 -14902 13682 -14842
rect 13742 -14902 14140 -14842
rect 14200 -14902 14596 -14842
rect 14656 -14902 15052 -14842
rect 15112 -14902 15508 -14842
rect 15568 -14902 15964 -14842
rect 16024 -14902 16422 -14842
rect 16482 -14902 16882 -14842
rect 10014 -14908 10074 -14902
rect 10470 -14908 10530 -14902
rect 10930 -14908 10990 -14902
rect 11386 -14908 11446 -14902
rect 11844 -14908 11904 -14902
rect 12308 -14908 12368 -14902
rect 12758 -14908 12818 -14902
rect 13214 -14908 13274 -14902
rect 13682 -14908 13742 -14902
rect 14140 -14908 14200 -14902
rect 14596 -14908 14656 -14902
rect 15052 -14908 15112 -14902
rect 15508 -14908 15568 -14902
rect 15964 -14908 16024 -14902
rect 16422 -14908 16482 -14902
rect 16882 -14908 16942 -14902
rect 25014 -14842 25074 -14836
rect 25470 -14842 25530 -14836
rect 25930 -14842 25990 -14836
rect 26386 -14842 26446 -14836
rect 26844 -14842 26904 -14836
rect 27308 -14842 27368 -14836
rect 27758 -14842 27818 -14836
rect 28214 -14842 28274 -14836
rect 28682 -14842 28742 -14836
rect 29140 -14842 29200 -14836
rect 29596 -14842 29656 -14836
rect 30052 -14842 30112 -14836
rect 30508 -14842 30568 -14836
rect 30964 -14842 31024 -14836
rect 31422 -14842 31482 -14836
rect 31882 -14842 31942 -14836
rect 25074 -14902 25470 -14842
rect 25530 -14902 25930 -14842
rect 25990 -14902 26386 -14842
rect 26446 -14902 26844 -14842
rect 26904 -14902 27308 -14842
rect 27368 -14902 27758 -14842
rect 27818 -14902 28214 -14842
rect 28274 -14902 28682 -14842
rect 28742 -14902 29140 -14842
rect 29200 -14902 29596 -14842
rect 29656 -14902 30052 -14842
rect 30112 -14902 30508 -14842
rect 30568 -14902 30964 -14842
rect 31024 -14902 31422 -14842
rect 31482 -14902 31882 -14842
rect 25014 -14908 25074 -14902
rect 25470 -14908 25530 -14902
rect 25930 -14908 25990 -14902
rect 26386 -14908 26446 -14902
rect 26844 -14908 26904 -14902
rect 27308 -14908 27368 -14902
rect 27758 -14908 27818 -14902
rect 28214 -14908 28274 -14902
rect 28682 -14908 28742 -14902
rect 29140 -14908 29200 -14902
rect 29596 -14908 29656 -14902
rect 30052 -14908 30112 -14902
rect 30508 -14908 30568 -14902
rect 30964 -14908 31024 -14902
rect 31422 -14908 31482 -14902
rect 31882 -14908 31942 -14902
rect 10010 -16816 10070 -16810
rect 10466 -16816 10526 -16810
rect 10926 -16816 10986 -16810
rect 11382 -16816 11442 -16810
rect 11840 -16816 11900 -16810
rect 12304 -16816 12364 -16810
rect 12758 -16816 12818 -16810
rect 13216 -16816 13276 -16810
rect 10070 -16876 10466 -16816
rect 10526 -16876 10926 -16816
rect 10986 -16876 11382 -16816
rect 11442 -16876 11840 -16816
rect 11900 -16876 12304 -16816
rect 12364 -16876 12758 -16816
rect 12818 -16876 13216 -16816
rect 13444 -16864 13450 -16804
rect 13510 -16864 13516 -16804
rect 13676 -16816 13736 -16810
rect 14132 -16816 14192 -16810
rect 14592 -16816 14652 -16810
rect 15048 -16816 15108 -16810
rect 15504 -16816 15564 -16810
rect 15960 -16816 16020 -16810
rect 16418 -16816 16478 -16810
rect 16878 -16816 16938 -16810
rect 22940 -16816 23000 -16810
rect 25010 -16816 25070 -16810
rect 25466 -16816 25526 -16810
rect 25926 -16816 25986 -16810
rect 26382 -16816 26442 -16810
rect 26840 -16816 26900 -16810
rect 27304 -16816 27364 -16810
rect 27758 -16816 27818 -16810
rect 28216 -16816 28276 -16810
rect 10010 -16882 10070 -16876
rect 10466 -16882 10526 -16876
rect 10926 -16882 10986 -16876
rect 11382 -16882 11442 -16876
rect 11840 -16882 11900 -16876
rect 12304 -16882 12364 -16876
rect 12758 -16882 12818 -16876
rect 13216 -16882 13276 -16876
rect 9224 -17402 9284 -17396
rect 13450 -17402 13510 -16864
rect 13736 -16876 14132 -16816
rect 14192 -16876 14592 -16816
rect 14652 -16876 15048 -16816
rect 15108 -16876 15504 -16816
rect 15564 -16876 15960 -16816
rect 16020 -16876 16418 -16816
rect 16478 -16876 16878 -16816
rect 16938 -16876 22940 -16816
rect 23000 -16876 25010 -16816
rect 25070 -16876 25466 -16816
rect 25526 -16876 25926 -16816
rect 25986 -16876 26382 -16816
rect 26442 -16876 26840 -16816
rect 26900 -16876 27304 -16816
rect 27364 -16876 27758 -16816
rect 27818 -16876 28216 -16816
rect 28444 -16864 28450 -16804
rect 28510 -16864 28516 -16804
rect 28676 -16816 28736 -16810
rect 29132 -16816 29192 -16810
rect 29592 -16816 29652 -16810
rect 30048 -16816 30108 -16810
rect 30504 -16816 30564 -16810
rect 30960 -16816 31020 -16810
rect 31418 -16816 31478 -16810
rect 31878 -16816 31938 -16810
rect 13676 -16882 13736 -16876
rect 14132 -16882 14192 -16876
rect 14592 -16882 14652 -16876
rect 15048 -16882 15108 -16876
rect 15504 -16882 15564 -16876
rect 15960 -16882 16020 -16876
rect 16418 -16882 16478 -16876
rect 16878 -16882 16938 -16876
rect 22940 -16882 23000 -16876
rect 25010 -16882 25070 -16876
rect 25466 -16882 25526 -16876
rect 25926 -16882 25986 -16876
rect 26382 -16882 26442 -16876
rect 26840 -16882 26900 -16876
rect 27304 -16882 27364 -16876
rect 27758 -16882 27818 -16876
rect 28216 -16882 28276 -16876
rect 9284 -17462 13510 -17402
rect 24224 -17402 24284 -17396
rect 28450 -17402 28510 -16864
rect 28736 -16876 29132 -16816
rect 29192 -16876 29592 -16816
rect 29652 -16876 30048 -16816
rect 30108 -16876 30504 -16816
rect 30564 -16876 30960 -16816
rect 31020 -16876 31418 -16816
rect 31478 -16876 31878 -16816
rect 28676 -16882 28736 -16876
rect 29132 -16882 29192 -16876
rect 29592 -16882 29652 -16876
rect 30048 -16882 30108 -16876
rect 30504 -16882 30564 -16876
rect 30960 -16882 31020 -16876
rect 31418 -16882 31478 -16876
rect 31878 -16882 31938 -16876
rect 24284 -17462 28510 -17402
rect 9224 -17468 9284 -17462
rect 24224 -17468 24284 -17462
rect 9442 -19140 9448 -19080
rect 9508 -19140 9514 -19080
rect 9904 -19140 9910 -19080
rect 9970 -19140 9976 -19080
rect 10358 -19136 10364 -19076
rect 10424 -19136 10430 -19076
rect 10820 -19136 10826 -19076
rect 10886 -19136 10892 -19076
rect 9448 -19534 9508 -19140
rect 9910 -19534 9970 -19140
rect 10364 -19534 10424 -19136
rect 10826 -19534 10886 -19136
rect 11274 -19142 11280 -19082
rect 11340 -19142 11346 -19082
rect 11724 -19136 11730 -19076
rect 11790 -19136 11796 -19076
rect 12190 -19136 12196 -19076
rect 12256 -19136 12262 -19076
rect 11280 -19534 11340 -19142
rect 11730 -19534 11790 -19136
rect 12196 -19534 12256 -19136
rect 12646 -19140 12652 -19080
rect 12712 -19140 12718 -19080
rect 14444 -19140 14450 -19080
rect 14510 -19140 14516 -19080
rect 14906 -19132 14912 -19072
rect 14972 -19132 14978 -19072
rect 12652 -19534 12712 -19140
rect 8164 -19594 12712 -19534
rect 9448 -20016 9508 -19594
rect 9910 -20010 9970 -19594
rect 9910 -20076 9970 -20070
rect 10364 -20016 10424 -19594
rect 10826 -20010 10886 -19594
rect 10826 -20076 10886 -20070
rect 11280 -20010 11340 -19594
rect 11280 -20076 11340 -20070
rect 11730 -20010 11790 -19594
rect 11730 -20076 11790 -20070
rect 12196 -20016 12256 -19594
rect 12652 -20010 12712 -19594
rect 12886 -19202 12946 -19196
rect 12886 -19540 12946 -19262
rect 14450 -19540 14510 -19140
rect 14912 -19540 14972 -19132
rect 15360 -19138 15366 -19078
rect 15426 -19138 15432 -19078
rect 15822 -19138 15828 -19078
rect 15888 -19138 15894 -19078
rect 16276 -19138 16282 -19078
rect 16342 -19138 16348 -19078
rect 16726 -19132 16732 -19072
rect 16792 -19132 16798 -19072
rect 15366 -19540 15426 -19138
rect 15828 -19540 15888 -19138
rect 16282 -19540 16342 -19138
rect 16732 -19540 16792 -19132
rect 17192 -19138 17198 -19078
rect 17258 -19138 17264 -19078
rect 17648 -19138 17654 -19078
rect 17714 -19138 17720 -19078
rect 17198 -19540 17258 -19138
rect 17654 -19540 17714 -19138
rect 24442 -19140 24448 -19080
rect 24508 -19140 24514 -19080
rect 24904 -19140 24910 -19080
rect 24970 -19140 24976 -19080
rect 25358 -19136 25364 -19076
rect 25424 -19136 25430 -19076
rect 25820 -19136 25826 -19076
rect 25886 -19136 25892 -19076
rect 17880 -19268 17886 -19208
rect 17946 -19268 17952 -19208
rect 12886 -19600 17714 -19540
rect 12886 -19882 12946 -19600
rect 12880 -19942 12886 -19882
rect 12946 -19942 12952 -19882
rect 12652 -20076 12712 -20070
rect 14450 -20010 14510 -19600
rect 14450 -20076 14510 -20070
rect 14912 -20012 14972 -19600
rect 9448 -20082 9508 -20076
rect 10364 -20082 10424 -20076
rect 12196 -20082 12256 -20076
rect 14912 -20078 14972 -20072
rect 15366 -20012 15426 -19600
rect 15366 -20078 15426 -20072
rect 15828 -20012 15888 -19600
rect 15828 -20078 15888 -20072
rect 16282 -20012 16342 -19600
rect 16732 -20006 16792 -19600
rect 16732 -20072 16792 -20066
rect 17198 -20010 17258 -19600
rect 16282 -20078 16342 -20072
rect 17198 -20076 17258 -20070
rect 17654 -20010 17714 -19600
rect 17886 -19544 17946 -19268
rect 24448 -19534 24508 -19140
rect 24910 -19534 24970 -19140
rect 25364 -19534 25424 -19136
rect 25826 -19534 25886 -19136
rect 26274 -19142 26280 -19082
rect 26340 -19142 26346 -19082
rect 26724 -19136 26730 -19076
rect 26790 -19136 26796 -19076
rect 27190 -19136 27196 -19076
rect 27256 -19136 27262 -19076
rect 26280 -19534 26340 -19142
rect 26730 -19534 26790 -19136
rect 27196 -19534 27256 -19136
rect 27646 -19140 27652 -19080
rect 27712 -19140 27718 -19080
rect 29444 -19140 29450 -19080
rect 29510 -19140 29516 -19080
rect 29906 -19132 29912 -19072
rect 29972 -19132 29978 -19072
rect 27652 -19534 27712 -19140
rect 17886 -19604 18972 -19544
rect 17886 -19870 17946 -19604
rect 18872 -19733 18972 -19604
rect 22954 -19594 27712 -19534
rect 22954 -19733 23014 -19594
rect 18868 -19823 18877 -19733
rect 18967 -19823 18976 -19733
rect 22932 -19823 22941 -19733
rect 23031 -19823 23040 -19733
rect 18872 -19828 18972 -19823
rect 22954 -19828 23014 -19823
rect 17886 -19936 17946 -19930
rect 17654 -20076 17714 -20070
rect 24448 -20016 24508 -19594
rect 24910 -20010 24970 -19594
rect 24910 -20076 24970 -20070
rect 25364 -20016 25424 -19594
rect 25826 -20010 25886 -19594
rect 25826 -20076 25886 -20070
rect 26280 -20010 26340 -19594
rect 26280 -20076 26340 -20070
rect 26730 -20010 26790 -19594
rect 26730 -20076 26790 -20070
rect 27196 -20016 27256 -19594
rect 27652 -20010 27712 -19594
rect 27886 -19202 27946 -19196
rect 27886 -19540 27946 -19262
rect 29450 -19540 29510 -19140
rect 29912 -19540 29972 -19132
rect 30360 -19138 30366 -19078
rect 30426 -19138 30432 -19078
rect 30822 -19138 30828 -19078
rect 30888 -19138 30894 -19078
rect 31276 -19138 31282 -19078
rect 31342 -19138 31348 -19078
rect 31726 -19132 31732 -19072
rect 31792 -19132 31798 -19072
rect 30366 -19540 30426 -19138
rect 30828 -19540 30888 -19138
rect 31282 -19540 31342 -19138
rect 31732 -19540 31792 -19132
rect 32192 -19138 32198 -19078
rect 32258 -19138 32264 -19078
rect 32648 -19138 32654 -19078
rect 32714 -19138 32720 -19078
rect 32198 -19540 32258 -19138
rect 32654 -19540 32714 -19138
rect 32880 -19268 32886 -19208
rect 32946 -19268 32952 -19208
rect 27886 -19600 32714 -19540
rect 27886 -19882 27946 -19600
rect 27880 -19942 27886 -19882
rect 27946 -19942 27952 -19882
rect 27652 -20076 27712 -20070
rect 29450 -20010 29510 -19600
rect 29450 -20076 29510 -20070
rect 29912 -20012 29972 -19600
rect 24448 -20082 24508 -20076
rect 25364 -20082 25424 -20076
rect 27196 -20082 27256 -20076
rect 29912 -20078 29972 -20072
rect 30366 -20012 30426 -19600
rect 30366 -20078 30426 -20072
rect 30828 -20012 30888 -19600
rect 30828 -20078 30888 -20072
rect 31282 -20012 31342 -19600
rect 31732 -20006 31792 -19600
rect 31732 -20072 31792 -20066
rect 32198 -20010 32258 -19600
rect 31282 -20078 31342 -20072
rect 32198 -20076 32258 -20070
rect 32654 -20010 32714 -19600
rect 32886 -19544 32946 -19268
rect 32886 -19604 33972 -19544
rect 32886 -19870 32946 -19604
rect 33872 -19733 33972 -19604
rect 37854 -19733 37914 -7222
rect 33868 -19823 33877 -19733
rect 33967 -19823 33976 -19733
rect 37830 -19823 37839 -19733
rect 37929 -19823 37938 -19733
rect 33872 -19828 33972 -19823
rect 37854 -19828 37914 -19823
rect 32886 -19936 32946 -19930
rect 32654 -20076 32714 -20070
rect 23080 -21226 23140 -21220
rect 24448 -21226 24508 -21220
rect 12646 -21286 12652 -21226
rect 12712 -21286 23080 -21226
rect 23140 -21286 24448 -21226
rect 23080 -21292 23140 -21286
rect 24448 -21292 24508 -21286
rect 8694 -21478 18464 -21450
rect 8694 -21564 8744 -21478
rect 8840 -21564 9324 -21478
rect 9420 -21564 9924 -21478
rect 10020 -21564 10524 -21478
rect 10620 -21564 11124 -21478
rect 11220 -21564 11724 -21478
rect 11820 -21564 12324 -21478
rect 12420 -21564 12924 -21478
rect 13020 -21564 13524 -21478
rect 13620 -21564 14124 -21478
rect 14220 -21564 14724 -21478
rect 14820 -21564 15324 -21478
rect 15420 -21564 15924 -21478
rect 16020 -21564 16524 -21478
rect 16620 -21564 17124 -21478
rect 17220 -21564 17724 -21478
rect 17820 -21564 18324 -21478
rect 18420 -21564 18464 -21478
rect 8694 -21594 18464 -21564
rect 23694 -21478 33464 -21450
rect 23694 -21564 23744 -21478
rect 23840 -21564 24324 -21478
rect 24420 -21564 24924 -21478
rect 25020 -21564 25524 -21478
rect 25620 -21564 26124 -21478
rect 26220 -21564 26724 -21478
rect 26820 -21564 27324 -21478
rect 27420 -21564 27924 -21478
rect 28020 -21564 28524 -21478
rect 28620 -21564 29124 -21478
rect 29220 -21564 29724 -21478
rect 29820 -21564 30324 -21478
rect 30420 -21564 30924 -21478
rect 31020 -21564 31524 -21478
rect 31620 -21564 32124 -21478
rect 32220 -21564 32724 -21478
rect 32820 -21564 33324 -21478
rect 33420 -21564 33464 -21478
rect 23694 -21594 33464 -21564
rect 8458 -21742 9058 -21732
rect 8458 -22052 9058 -22042
rect 18090 -21742 18690 -21732
rect 18090 -22052 18690 -22042
rect 23458 -21742 24058 -21732
rect 23458 -22052 24058 -22042
rect 33090 -21742 33690 -21732
rect 33090 -22052 33690 -22042
<< via2 >>
rect 23440 17094 24040 17394
rect 32072 17094 32672 17394
rect 23562 16868 32558 16978
rect 13066 10328 13448 10628
rect 21200 10328 21878 10628
rect 15134 10064 15230 10150
rect 15714 10064 15810 10150
rect 16314 10064 16410 10150
rect 16914 10064 17010 10150
rect 17514 10064 17610 10150
rect 18114 10064 18210 10150
rect 18714 10064 18810 10150
rect 19314 10064 19410 10150
rect 19914 10064 20010 10150
rect 27157 14101 27247 14191
rect 34630 13582 34690 13642
rect 24176 11572 32038 11716
rect 23440 11162 24040 11462
rect 32072 11162 32672 11462
rect 23648 10328 24248 10628
rect 28280 10328 28880 10628
rect 23896 10064 23992 10150
rect 24476 10064 24572 10150
rect 25076 10064 25172 10150
rect 25676 10064 25772 10150
rect 26276 10064 26372 10150
rect 26876 10064 26972 10150
rect 27476 10064 27572 10150
rect 28076 10064 28172 10150
rect 28676 10064 28772 10150
rect 33086 8924 33182 8996
rect 30406 8380 30502 8452
rect 35784 8380 35880 8452
rect 33086 7836 33182 7908
rect 30406 7292 30502 7364
rect 35784 7292 35880 7364
rect 33086 6748 33182 6820
rect 30406 6204 30502 6276
rect 35784 6204 35880 6276
rect 33086 5660 33182 5732
rect 13308 5346 13404 5432
rect 13908 5346 14004 5432
rect 14508 5346 14604 5432
rect 15108 5346 15204 5432
rect 15708 5346 15804 5432
rect 16308 5346 16404 5432
rect 16908 5346 17004 5432
rect 17508 5346 17604 5432
rect 18108 5346 18204 5432
rect 18708 5346 18804 5432
rect 19308 5346 19404 5432
rect 19908 5346 20004 5432
rect 20508 5346 20604 5432
rect 21108 5346 21204 5432
rect 21528 5346 21624 5432
rect 23824 5346 23920 5432
rect 24424 5346 24520 5432
rect 25024 5346 25120 5432
rect 25624 5346 25720 5432
rect 26224 5346 26320 5432
rect 26824 5346 26920 5432
rect 27424 5346 27520 5432
rect 28024 5346 28120 5432
rect 28624 5346 28720 5432
rect 13066 4872 13448 5172
rect 21200 4872 21878 5172
rect 23648 4872 24248 5172
rect 28280 4872 28880 5172
rect 8458 3990 9058 4290
rect 18090 3990 18690 4290
rect 23458 3990 24058 4290
rect 33090 3990 33690 4290
rect 9310 3730 9406 3816
rect 9910 3730 10006 3816
rect 10510 3730 10606 3816
rect 11110 3730 11206 3816
rect 11710 3730 11806 3816
rect 12310 3730 12406 3816
rect 12910 3730 13006 3816
rect 13510 3730 13606 3816
rect 14110 3730 14206 3816
rect 14710 3730 14806 3816
rect 15310 3730 15406 3816
rect 15910 3730 16006 3816
rect 16510 3730 16606 3816
rect 17110 3730 17206 3816
rect 17530 3730 17626 3816
rect 24310 3730 24406 3816
rect 24910 3730 25006 3816
rect 25510 3730 25606 3816
rect 26110 3730 26206 3816
rect 26710 3730 26806 3816
rect 27310 3730 27406 3816
rect 27910 3730 28006 3816
rect 28510 3730 28606 3816
rect 29110 3730 29206 3816
rect 29710 3730 29806 3816
rect 30310 3730 30406 3816
rect 30910 3730 31006 3816
rect 31510 3730 31606 3816
rect 32110 3730 32206 3816
rect 32530 3730 32626 3816
rect 23150 -1594 23210 -1534
rect 18877 -1823 18967 -1733
rect 33877 -1823 33967 -1733
rect 8744 -3564 8840 -3478
rect 9324 -3564 9420 -3478
rect 9924 -3564 10020 -3478
rect 10524 -3564 10620 -3478
rect 11124 -3564 11220 -3478
rect 11724 -3564 11820 -3478
rect 12324 -3564 12420 -3478
rect 12924 -3564 13020 -3478
rect 13524 -3564 13620 -3478
rect 14124 -3564 14220 -3478
rect 14724 -3564 14820 -3478
rect 15324 -3564 15420 -3478
rect 15924 -3564 16020 -3478
rect 16524 -3564 16620 -3478
rect 17124 -3564 17220 -3478
rect 17724 -3564 17820 -3478
rect 18324 -3564 18420 -3478
rect 23744 -3564 23840 -3478
rect 24324 -3564 24420 -3478
rect 24924 -3564 25020 -3478
rect 25524 -3564 25620 -3478
rect 26124 -3564 26220 -3478
rect 26724 -3564 26820 -3478
rect 27324 -3564 27420 -3478
rect 27924 -3564 28020 -3478
rect 28524 -3564 28620 -3478
rect 29124 -3564 29220 -3478
rect 29724 -3564 29820 -3478
rect 30324 -3564 30420 -3478
rect 30924 -3564 31020 -3478
rect 31524 -3564 31620 -3478
rect 32124 -3564 32220 -3478
rect 32724 -3564 32820 -3478
rect 33324 -3564 33420 -3478
rect 8458 -4042 9058 -3742
rect 18090 -4042 18690 -3742
rect 23458 -4042 24058 -3742
rect 33090 -4042 33690 -3742
rect 12412 -5014 13012 -4714
rect 22044 -5014 22644 -4714
rect 27412 -5014 28012 -4714
rect 37044 -5014 37644 -4714
rect 12682 -5278 12778 -5192
rect 13282 -5278 13378 -5192
rect 13882 -5278 13978 -5192
rect 14482 -5278 14578 -5192
rect 15082 -5278 15178 -5192
rect 15682 -5278 15778 -5192
rect 16282 -5278 16378 -5192
rect 16882 -5278 16978 -5192
rect 17482 -5278 17578 -5192
rect 18082 -5278 18178 -5192
rect 18682 -5278 18778 -5192
rect 19282 -5278 19378 -5192
rect 19882 -5278 19978 -5192
rect 20482 -5278 20578 -5192
rect 21082 -5278 21178 -5192
rect 21682 -5278 21778 -5192
rect 22262 -5278 22358 -5192
rect 27682 -5278 27778 -5192
rect 28282 -5278 28378 -5192
rect 28882 -5278 28978 -5192
rect 29482 -5278 29578 -5192
rect 30082 -5278 30178 -5192
rect 30682 -5278 30778 -5192
rect 31282 -5278 31378 -5192
rect 31882 -5278 31978 -5192
rect 32482 -5278 32578 -5192
rect 33082 -5278 33178 -5192
rect 33682 -5278 33778 -5192
rect 34282 -5278 34378 -5192
rect 34882 -5278 34978 -5192
rect 35482 -5278 35578 -5192
rect 36082 -5278 36178 -5192
rect 36682 -5278 36778 -5192
rect 37262 -5278 37358 -5192
rect 8143 -7023 8233 -6933
rect 12135 -7023 12225 -6933
rect 27135 -7023 27225 -6933
rect 22834 -7222 22894 -7162
rect 13476 -12572 13572 -12486
rect 13896 -12572 13992 -12486
rect 14496 -12572 14592 -12486
rect 15096 -12572 15192 -12486
rect 15696 -12572 15792 -12486
rect 16296 -12572 16392 -12486
rect 16896 -12572 16992 -12486
rect 17496 -12572 17592 -12486
rect 18096 -12572 18192 -12486
rect 18696 -12572 18792 -12486
rect 19296 -12572 19392 -12486
rect 19896 -12572 19992 -12486
rect 20496 -12572 20592 -12486
rect 21096 -12572 21192 -12486
rect 21696 -12572 21792 -12486
rect 28476 -12572 28572 -12486
rect 28896 -12572 28992 -12486
rect 29496 -12572 29592 -12486
rect 30096 -12572 30192 -12486
rect 30696 -12572 30792 -12486
rect 31296 -12572 31392 -12486
rect 31896 -12572 31992 -12486
rect 32496 -12572 32592 -12486
rect 33096 -12572 33192 -12486
rect 33696 -12572 33792 -12486
rect 34296 -12572 34392 -12486
rect 34896 -12572 34992 -12486
rect 35496 -12572 35592 -12486
rect 36096 -12572 36192 -12486
rect 36696 -12572 36792 -12486
rect 12412 -13046 13012 -12746
rect 22044 -13046 22644 -12746
rect 27412 -13046 28012 -12746
rect 37044 -13046 37644 -12746
rect 8458 -14010 9058 -13710
rect 18090 -14010 18690 -13710
rect 23458 -14010 24058 -13710
rect 33090 -14010 33690 -13710
rect 9310 -14270 9406 -14184
rect 9910 -14270 10006 -14184
rect 10510 -14270 10606 -14184
rect 11110 -14270 11206 -14184
rect 11710 -14270 11806 -14184
rect 12310 -14270 12406 -14184
rect 12910 -14270 13006 -14184
rect 13510 -14270 13606 -14184
rect 14110 -14270 14206 -14184
rect 14710 -14270 14806 -14184
rect 15310 -14270 15406 -14184
rect 15910 -14270 16006 -14184
rect 16510 -14270 16606 -14184
rect 17110 -14270 17206 -14184
rect 17530 -14270 17626 -14184
rect 24310 -14270 24406 -14184
rect 24910 -14270 25006 -14184
rect 25510 -14270 25606 -14184
rect 26110 -14270 26206 -14184
rect 26710 -14270 26806 -14184
rect 27310 -14270 27406 -14184
rect 27910 -14270 28006 -14184
rect 28510 -14270 28606 -14184
rect 29110 -14270 29206 -14184
rect 29710 -14270 29806 -14184
rect 30310 -14270 30406 -14184
rect 30910 -14270 31006 -14184
rect 31510 -14270 31606 -14184
rect 32110 -14270 32206 -14184
rect 32530 -14270 32626 -14184
rect 18877 -19823 18967 -19733
rect 22941 -19823 23031 -19733
rect 33877 -19823 33967 -19733
rect 37839 -19823 37929 -19733
rect 8744 -21564 8840 -21478
rect 9324 -21564 9420 -21478
rect 9924 -21564 10020 -21478
rect 10524 -21564 10620 -21478
rect 11124 -21564 11220 -21478
rect 11724 -21564 11820 -21478
rect 12324 -21564 12420 -21478
rect 12924 -21564 13020 -21478
rect 13524 -21564 13620 -21478
rect 14124 -21564 14220 -21478
rect 14724 -21564 14820 -21478
rect 15324 -21564 15420 -21478
rect 15924 -21564 16020 -21478
rect 16524 -21564 16620 -21478
rect 17124 -21564 17220 -21478
rect 17724 -21564 17820 -21478
rect 18324 -21564 18420 -21478
rect 23744 -21564 23840 -21478
rect 24324 -21564 24420 -21478
rect 24924 -21564 25020 -21478
rect 25524 -21564 25620 -21478
rect 26124 -21564 26220 -21478
rect 26724 -21564 26820 -21478
rect 27324 -21564 27420 -21478
rect 27924 -21564 28020 -21478
rect 28524 -21564 28620 -21478
rect 29124 -21564 29220 -21478
rect 29724 -21564 29820 -21478
rect 30324 -21564 30420 -21478
rect 30924 -21564 31020 -21478
rect 31524 -21564 31620 -21478
rect 32124 -21564 32220 -21478
rect 32724 -21564 32820 -21478
rect 33324 -21564 33420 -21478
rect 8458 -22042 9058 -21742
rect 18090 -22042 18690 -21742
rect 23458 -22042 24058 -21742
rect 33090 -22042 33690 -21742
<< metal3 >>
rect 23430 17394 24050 17399
rect 23430 17094 23440 17394
rect 24040 17094 24050 17394
rect 23430 17089 24050 17094
rect 32062 17394 32682 17399
rect 32062 17094 32072 17394
rect 32672 17094 32682 17394
rect 32062 17089 32682 17094
rect 23526 16978 32596 17012
rect 23526 16868 23562 16978
rect 32558 16868 32596 16978
rect 23526 16830 32596 16868
rect 27152 14191 27252 14196
rect 27152 14101 27157 14191
rect 27247 14101 27252 14191
rect 27152 13664 27252 14101
rect 27152 13642 34698 13664
rect 27152 13582 34630 13642
rect 34690 13582 34698 13642
rect 27152 13564 34698 13582
rect 24136 11716 32076 11756
rect 24136 11572 24176 11716
rect 32038 11572 32076 11716
rect 24136 11542 32076 11572
rect 23430 11462 24050 11467
rect 23430 11162 23440 11462
rect 24040 11162 24050 11462
rect 23430 11157 24050 11162
rect 32062 11462 32682 11467
rect 32062 11162 32072 11462
rect 32672 11162 32682 11462
rect 32062 11157 32682 11162
rect 13056 10628 13458 10633
rect 13056 10328 13066 10628
rect 13448 10328 13458 10628
rect 13056 10323 13458 10328
rect 21190 10628 21888 10633
rect 21190 10328 21200 10628
rect 21878 10328 21888 10628
rect 21190 10323 21888 10328
rect 23638 10628 24258 10633
rect 23638 10328 23648 10628
rect 24248 10328 24258 10628
rect 23638 10323 24258 10328
rect 28270 10628 28890 10633
rect 28270 10328 28280 10628
rect 28880 10328 28890 10628
rect 28270 10323 28890 10328
rect 15084 10150 20056 10180
rect 15084 10064 15134 10150
rect 15230 10064 15714 10150
rect 15810 10064 16314 10150
rect 16410 10064 16914 10150
rect 17010 10064 17514 10150
rect 17610 10064 18114 10150
rect 18210 10064 18714 10150
rect 18810 10064 19314 10150
rect 19410 10064 19914 10150
rect 20010 10064 20056 10150
rect 15084 10036 20056 10064
rect 23846 10150 28818 10180
rect 23846 10064 23896 10150
rect 23992 10064 24476 10150
rect 24572 10064 25076 10150
rect 25172 10064 25676 10150
rect 25772 10064 26276 10150
rect 26372 10064 26876 10150
rect 26972 10064 27476 10150
rect 27572 10064 28076 10150
rect 28172 10064 28676 10150
rect 28772 10064 28818 10150
rect 23846 10036 28818 10064
rect 33074 8996 33194 9008
rect 33074 8924 33086 8996
rect 33182 8924 33194 8996
rect 33074 8912 33194 8924
rect 30394 8452 30514 8464
rect 30394 8380 30406 8452
rect 30502 8380 30514 8452
rect 30394 8368 30514 8380
rect 35772 8452 35892 8464
rect 35772 8380 35784 8452
rect 35880 8380 35892 8452
rect 35772 8368 35892 8380
rect 33074 7908 33194 7920
rect 33074 7836 33086 7908
rect 33182 7836 33194 7908
rect 33074 7824 33194 7836
rect 30394 7364 30514 7376
rect 30394 7292 30406 7364
rect 30502 7292 30514 7364
rect 30394 7280 30514 7292
rect 35772 7364 35892 7376
rect 35772 7292 35784 7364
rect 35880 7292 35892 7364
rect 35772 7280 35892 7292
rect 33074 6820 33194 6832
rect 33074 6748 33086 6820
rect 33182 6748 33194 6820
rect 33074 6736 33194 6748
rect 30394 6276 30514 6288
rect 30394 6204 30406 6276
rect 30502 6204 30514 6276
rect 30394 6192 30514 6204
rect 35772 6276 35892 6288
rect 35772 6204 35784 6276
rect 35880 6204 35892 6276
rect 35772 6192 35892 6204
rect 33074 5732 33194 5744
rect 33074 5660 33086 5732
rect 33182 5660 33194 5732
rect 33074 5648 33194 5660
rect 13294 5432 21650 5442
rect 13294 5346 13308 5432
rect 13404 5346 13908 5432
rect 14004 5346 14508 5432
rect 14604 5346 15108 5432
rect 15204 5346 15708 5432
rect 15804 5346 16308 5432
rect 16404 5346 16908 5432
rect 17004 5346 17508 5432
rect 17604 5346 18108 5432
rect 18204 5346 18708 5432
rect 18804 5346 19308 5432
rect 19404 5346 19908 5432
rect 20004 5346 20508 5432
rect 20604 5346 21108 5432
rect 21204 5346 21528 5432
rect 21624 5346 21650 5432
rect 13294 5332 21650 5346
rect 23810 5432 28808 5442
rect 23810 5346 23824 5432
rect 23920 5346 24424 5432
rect 24520 5346 25024 5432
rect 25120 5346 25624 5432
rect 25720 5346 26224 5432
rect 26320 5346 26824 5432
rect 26920 5346 27424 5432
rect 27520 5346 28024 5432
rect 28120 5346 28624 5432
rect 28720 5346 28808 5432
rect 23810 5332 28808 5346
rect 13056 5172 13458 5177
rect 13056 4872 13066 5172
rect 13448 4872 13458 5172
rect 13056 4867 13458 4872
rect 21190 5172 21888 5177
rect 21190 4872 21200 5172
rect 21878 4872 21888 5172
rect 21190 4867 21888 4872
rect 23638 5172 24258 5177
rect 23638 4872 23648 5172
rect 24248 4872 24258 5172
rect 23638 4867 24258 4872
rect 28270 5172 28890 5177
rect 28270 4872 28280 5172
rect 28880 4872 28890 5172
rect 28270 4867 28890 4872
rect 8448 4290 9068 4295
rect 8448 3990 8458 4290
rect 9058 3990 9068 4290
rect 8448 3985 9068 3990
rect 18080 4290 18700 4295
rect 18080 3990 18090 4290
rect 18690 3990 18700 4290
rect 18080 3985 18700 3990
rect 23448 4290 24068 4295
rect 23448 3990 23458 4290
rect 24058 3990 24068 4290
rect 23448 3985 24068 3990
rect 33080 4290 33700 4295
rect 33080 3990 33090 4290
rect 33690 3990 33700 4290
rect 33080 3985 33700 3990
rect 9296 3816 17652 3830
rect 9296 3730 9310 3816
rect 9406 3730 9910 3816
rect 10006 3730 10510 3816
rect 10606 3730 11110 3816
rect 11206 3730 11710 3816
rect 11806 3730 12310 3816
rect 12406 3730 12910 3816
rect 13006 3730 13510 3816
rect 13606 3730 14110 3816
rect 14206 3730 14710 3816
rect 14806 3730 15310 3816
rect 15406 3730 15910 3816
rect 16006 3730 16510 3816
rect 16606 3730 17110 3816
rect 17206 3730 17530 3816
rect 17626 3730 17652 3816
rect 9296 3720 17652 3730
rect 24296 3816 32652 3830
rect 24296 3730 24310 3816
rect 24406 3730 24910 3816
rect 25006 3730 25510 3816
rect 25606 3730 26110 3816
rect 26206 3730 26710 3816
rect 26806 3730 27310 3816
rect 27406 3730 27910 3816
rect 28006 3730 28510 3816
rect 28606 3730 29110 3816
rect 29206 3730 29710 3816
rect 29806 3730 30310 3816
rect 30406 3730 30910 3816
rect 31006 3730 31510 3816
rect 31606 3730 32110 3816
rect 32206 3730 32530 3816
rect 32626 3730 32652 3816
rect 24296 3720 32652 3730
rect 19072 -542 22700 -408
rect 19072 -914 19709 -542
rect 19773 -544 22700 -542
rect 19773 -914 20428 -544
rect 20492 -914 21147 -544
rect 21211 -914 21866 -544
rect 21930 -914 22585 -544
rect 22649 -914 22700 -544
rect 19072 -1244 22700 -914
rect 19072 -1612 19709 -1244
rect 19773 -1612 20428 -1244
rect 20492 -1612 21147 -1244
rect 21211 -1612 21866 -1244
rect 21930 -1612 22585 -1244
rect 22649 -1612 22700 -1244
rect 34072 -542 37700 -408
rect 34072 -914 34709 -542
rect 34773 -544 37700 -542
rect 34773 -914 35428 -544
rect 35492 -914 36147 -544
rect 36211 -914 36866 -544
rect 36930 -914 37585 -544
rect 37649 -914 37700 -544
rect 34072 -1244 37700 -914
rect 23145 -1534 23215 -1529
rect 18872 -1729 18972 -1728
rect 18867 -1827 18873 -1729
rect 18971 -1827 18977 -1729
rect 18872 -1828 18972 -1827
rect 19072 -1944 22700 -1612
rect 23130 -1594 23150 -1534
rect 23210 -1594 23230 -1534
rect 22806 -1729 22906 -1728
rect 22801 -1827 22807 -1729
rect 22905 -1827 22911 -1729
rect 19072 -2312 19709 -1944
rect 19773 -2312 20428 -1944
rect 20492 -2312 21147 -1944
rect 21211 -2312 21866 -1944
rect 21930 -2312 22585 -1944
rect 22649 -2312 22700 -1944
rect 19072 -2644 22700 -2312
rect 19072 -3012 19709 -2644
rect 19773 -3012 20428 -2644
rect 20492 -3012 21147 -2644
rect 21211 -3012 21866 -2644
rect 21930 -3012 22585 -2644
rect 22649 -3012 22700 -2644
rect 19072 -3344 22700 -3012
rect 8694 -3478 18464 -3450
rect 8694 -3564 8744 -3478
rect 8840 -3564 9324 -3478
rect 9420 -3564 9924 -3478
rect 10020 -3564 10524 -3478
rect 10620 -3564 11124 -3478
rect 11220 -3564 11724 -3478
rect 11820 -3564 12324 -3478
rect 12420 -3564 12924 -3478
rect 13020 -3564 13524 -3478
rect 13620 -3564 14124 -3478
rect 14220 -3564 14724 -3478
rect 14820 -3564 15324 -3478
rect 15420 -3564 15924 -3478
rect 16020 -3564 16524 -3478
rect 16620 -3564 17124 -3478
rect 17220 -3564 17724 -3478
rect 17820 -3564 18324 -3478
rect 18420 -3564 18464 -3478
rect 8694 -3594 18464 -3564
rect 19072 -3712 19709 -3344
rect 19773 -3712 20428 -3344
rect 20492 -3712 21147 -3344
rect 21211 -3712 21866 -3344
rect 21930 -3712 22585 -3344
rect 22649 -3712 22700 -3344
rect 8448 -3742 9068 -3737
rect 8448 -4042 8458 -3742
rect 9058 -4042 9068 -3742
rect 8448 -4047 9068 -4042
rect 18080 -3742 18700 -3737
rect 18080 -4042 18090 -3742
rect 18690 -4042 18700 -3742
rect 19072 -3862 22700 -3712
rect 18080 -4047 18700 -4042
rect 12402 -4714 13022 -4709
rect 8402 -5044 12030 -4894
rect 12402 -5014 12412 -4714
rect 13012 -5014 13022 -4714
rect 12402 -5019 13022 -5014
rect 22034 -4714 22654 -4709
rect 22034 -5014 22044 -4714
rect 22644 -5014 22654 -4714
rect 22034 -5019 22654 -5014
rect 8402 -5412 8453 -5044
rect 8517 -5412 9172 -5044
rect 9236 -5412 9891 -5044
rect 9955 -5412 10610 -5044
rect 10674 -5412 11329 -5044
rect 11393 -5412 12030 -5044
rect 12638 -5192 22408 -5162
rect 12638 -5278 12682 -5192
rect 12778 -5278 13282 -5192
rect 13378 -5278 13882 -5192
rect 13978 -5278 14482 -5192
rect 14578 -5278 15082 -5192
rect 15178 -5278 15682 -5192
rect 15778 -5278 16282 -5192
rect 16378 -5278 16882 -5192
rect 16978 -5278 17482 -5192
rect 17578 -5278 18082 -5192
rect 18178 -5278 18682 -5192
rect 18778 -5278 19282 -5192
rect 19378 -5278 19882 -5192
rect 19978 -5278 20482 -5192
rect 20578 -5278 21082 -5192
rect 21178 -5278 21682 -5192
rect 21778 -5278 22262 -5192
rect 22358 -5278 22408 -5192
rect 12638 -5306 22408 -5278
rect 8402 -5744 12030 -5412
rect 8402 -6112 8453 -5744
rect 8517 -6112 9172 -5744
rect 9236 -6112 9891 -5744
rect 9955 -6112 10610 -5744
rect 10674 -6112 11329 -5744
rect 11393 -6112 12030 -5744
rect 8402 -6444 12030 -6112
rect 8402 -6812 8453 -6444
rect 8517 -6812 9172 -6444
rect 9236 -6812 9891 -6444
rect 9955 -6812 10610 -6444
rect 10674 -6812 11329 -6444
rect 11393 -6812 12030 -6444
rect 8138 -6929 8238 -6928
rect 8133 -7027 8139 -6929
rect 8237 -7027 8243 -6929
rect 8138 -7028 8238 -7027
rect 8402 -7144 12030 -6812
rect 12130 -6929 12230 -6928
rect 12125 -7027 12131 -6929
rect 12229 -7027 12235 -6929
rect 12130 -7028 12230 -7027
rect 8402 -7512 8453 -7144
rect 8517 -7512 9172 -7144
rect 9236 -7512 9891 -7144
rect 9955 -7512 10610 -7144
rect 10674 -7512 11329 -7144
rect 11393 -7512 12030 -7144
rect 22806 -7162 22906 -1827
rect 23130 -6929 23230 -1594
rect 34072 -1612 34709 -1244
rect 34773 -1612 35428 -1244
rect 35492 -1612 36147 -1244
rect 36211 -1612 36866 -1244
rect 36930 -1612 37585 -1244
rect 37649 -1612 37700 -1244
rect 33872 -1729 33972 -1728
rect 33867 -1827 33873 -1729
rect 33971 -1827 33977 -1729
rect 33872 -1828 33972 -1827
rect 34072 -1944 37700 -1612
rect 34072 -2312 34709 -1944
rect 34773 -2312 35428 -1944
rect 35492 -2312 36147 -1944
rect 36211 -2312 36866 -1944
rect 36930 -2312 37585 -1944
rect 37649 -2312 37700 -1944
rect 34072 -2644 37700 -2312
rect 34072 -3012 34709 -2644
rect 34773 -3012 35428 -2644
rect 35492 -3012 36147 -2644
rect 36211 -3012 36866 -2644
rect 36930 -3012 37585 -2644
rect 37649 -3012 37700 -2644
rect 34072 -3344 37700 -3012
rect 23694 -3478 33464 -3450
rect 23694 -3564 23744 -3478
rect 23840 -3564 24324 -3478
rect 24420 -3564 24924 -3478
rect 25020 -3564 25524 -3478
rect 25620 -3564 26124 -3478
rect 26220 -3564 26724 -3478
rect 26820 -3564 27324 -3478
rect 27420 -3564 27924 -3478
rect 28020 -3564 28524 -3478
rect 28620 -3564 29124 -3478
rect 29220 -3564 29724 -3478
rect 29820 -3564 30324 -3478
rect 30420 -3564 30924 -3478
rect 31020 -3564 31524 -3478
rect 31620 -3564 32124 -3478
rect 32220 -3564 32724 -3478
rect 32820 -3564 33324 -3478
rect 33420 -3564 33464 -3478
rect 23694 -3594 33464 -3564
rect 34072 -3712 34709 -3344
rect 34773 -3712 35428 -3344
rect 35492 -3712 36147 -3344
rect 36211 -3712 36866 -3344
rect 36930 -3712 37585 -3344
rect 37649 -3712 37700 -3344
rect 23448 -3742 24068 -3737
rect 23448 -4042 23458 -3742
rect 24058 -4042 24068 -3742
rect 23448 -4047 24068 -4042
rect 33080 -3742 33700 -3737
rect 33080 -4042 33090 -3742
rect 33690 -4042 33700 -3742
rect 34072 -3862 37700 -3712
rect 33080 -4047 33700 -4042
rect 27402 -4714 28022 -4709
rect 23402 -5044 27030 -4894
rect 27402 -5014 27412 -4714
rect 28012 -5014 28022 -4714
rect 27402 -5019 28022 -5014
rect 37034 -4714 37654 -4709
rect 37034 -5014 37044 -4714
rect 37644 -5014 37654 -4714
rect 37034 -5019 37654 -5014
rect 23402 -5412 23453 -5044
rect 23517 -5412 24172 -5044
rect 24236 -5412 24891 -5044
rect 24955 -5412 25610 -5044
rect 25674 -5412 26329 -5044
rect 26393 -5412 27030 -5044
rect 27638 -5192 37408 -5162
rect 27638 -5278 27682 -5192
rect 27778 -5278 28282 -5192
rect 28378 -5278 28882 -5192
rect 28978 -5278 29482 -5192
rect 29578 -5278 30082 -5192
rect 30178 -5278 30682 -5192
rect 30778 -5278 31282 -5192
rect 31378 -5278 31882 -5192
rect 31978 -5278 32482 -5192
rect 32578 -5278 33082 -5192
rect 33178 -5278 33682 -5192
rect 33778 -5278 34282 -5192
rect 34378 -5278 34882 -5192
rect 34978 -5278 35482 -5192
rect 35578 -5278 36082 -5192
rect 36178 -5278 36682 -5192
rect 36778 -5278 37262 -5192
rect 37358 -5278 37408 -5192
rect 27638 -5306 37408 -5278
rect 23402 -5744 27030 -5412
rect 23402 -6112 23453 -5744
rect 23517 -6112 24172 -5744
rect 24236 -6112 24891 -5744
rect 24955 -6112 25610 -5744
rect 25674 -6112 26329 -5744
rect 26393 -6112 27030 -5744
rect 23402 -6444 27030 -6112
rect 23402 -6812 23453 -6444
rect 23517 -6812 24172 -6444
rect 24236 -6812 24891 -6444
rect 24955 -6812 25610 -6444
rect 25674 -6812 26329 -6444
rect 26393 -6812 27030 -6444
rect 23125 -7027 23131 -6929
rect 23229 -7027 23235 -6929
rect 23130 -7028 23230 -7027
rect 22806 -7222 22834 -7162
rect 22894 -7222 22906 -7162
rect 22806 -7238 22906 -7222
rect 23402 -7144 27030 -6812
rect 27130 -6929 27230 -6928
rect 27125 -7027 27131 -6929
rect 27229 -7027 27235 -6929
rect 27130 -7028 27230 -7027
rect 8402 -7842 12030 -7512
rect 8402 -8212 8453 -7842
rect 8517 -8212 9172 -7842
rect 9236 -8212 9891 -7842
rect 9955 -8212 10610 -7842
rect 10674 -8212 11329 -7842
rect 8402 -8214 11329 -8212
rect 11393 -8214 12030 -7842
rect 8402 -8348 12030 -8214
rect 23402 -7512 23453 -7144
rect 23517 -7512 24172 -7144
rect 24236 -7512 24891 -7144
rect 24955 -7512 25610 -7144
rect 25674 -7512 26329 -7144
rect 26393 -7512 27030 -7144
rect 23402 -7842 27030 -7512
rect 23402 -8212 23453 -7842
rect 23517 -8212 24172 -7842
rect 24236 -8212 24891 -7842
rect 24955 -8212 25610 -7842
rect 25674 -8212 26329 -7842
rect 23402 -8214 26329 -8212
rect 26393 -8214 27030 -7842
rect 23402 -8348 27030 -8214
rect 13450 -12486 21806 -12476
rect 13450 -12572 13476 -12486
rect 13572 -12572 13896 -12486
rect 13992 -12572 14496 -12486
rect 14592 -12572 15096 -12486
rect 15192 -12572 15696 -12486
rect 15792 -12572 16296 -12486
rect 16392 -12572 16896 -12486
rect 16992 -12572 17496 -12486
rect 17592 -12572 18096 -12486
rect 18192 -12572 18696 -12486
rect 18792 -12572 19296 -12486
rect 19392 -12572 19896 -12486
rect 19992 -12572 20496 -12486
rect 20592 -12572 21096 -12486
rect 21192 -12572 21696 -12486
rect 21792 -12572 21806 -12486
rect 13450 -12586 21806 -12572
rect 28450 -12486 36806 -12476
rect 28450 -12572 28476 -12486
rect 28572 -12572 28896 -12486
rect 28992 -12572 29496 -12486
rect 29592 -12572 30096 -12486
rect 30192 -12572 30696 -12486
rect 30792 -12572 31296 -12486
rect 31392 -12572 31896 -12486
rect 31992 -12572 32496 -12486
rect 32592 -12572 33096 -12486
rect 33192 -12572 33696 -12486
rect 33792 -12572 34296 -12486
rect 34392 -12572 34896 -12486
rect 34992 -12572 35496 -12486
rect 35592 -12572 36096 -12486
rect 36192 -12572 36696 -12486
rect 36792 -12572 36806 -12486
rect 28450 -12586 36806 -12572
rect 12402 -12746 13022 -12741
rect 12402 -13046 12412 -12746
rect 13012 -13046 13022 -12746
rect 12402 -13051 13022 -13046
rect 22034 -12746 22654 -12741
rect 22034 -13046 22044 -12746
rect 22644 -13046 22654 -12746
rect 22034 -13051 22654 -13046
rect 27402 -12746 28022 -12741
rect 27402 -13046 27412 -12746
rect 28012 -13046 28022 -12746
rect 27402 -13051 28022 -13046
rect 37034 -12746 37654 -12741
rect 37034 -13046 37044 -12746
rect 37644 -13046 37654 -12746
rect 37034 -13051 37654 -13046
rect 8448 -13710 9068 -13705
rect 8448 -14010 8458 -13710
rect 9058 -14010 9068 -13710
rect 8448 -14015 9068 -14010
rect 18080 -13710 18700 -13705
rect 18080 -14010 18090 -13710
rect 18690 -14010 18700 -13710
rect 18080 -14015 18700 -14010
rect 23448 -13710 24068 -13705
rect 23448 -14010 23458 -13710
rect 24058 -14010 24068 -13710
rect 23448 -14015 24068 -14010
rect 33080 -13710 33700 -13705
rect 33080 -14010 33090 -13710
rect 33690 -14010 33700 -13710
rect 33080 -14015 33700 -14010
rect 9296 -14184 17652 -14170
rect 9296 -14270 9310 -14184
rect 9406 -14270 9910 -14184
rect 10006 -14270 10510 -14184
rect 10606 -14270 11110 -14184
rect 11206 -14270 11710 -14184
rect 11806 -14270 12310 -14184
rect 12406 -14270 12910 -14184
rect 13006 -14270 13510 -14184
rect 13606 -14270 14110 -14184
rect 14206 -14270 14710 -14184
rect 14806 -14270 15310 -14184
rect 15406 -14270 15910 -14184
rect 16006 -14270 16510 -14184
rect 16606 -14270 17110 -14184
rect 17206 -14270 17530 -14184
rect 17626 -14270 17652 -14184
rect 9296 -14280 17652 -14270
rect 24296 -14184 32652 -14170
rect 24296 -14270 24310 -14184
rect 24406 -14270 24910 -14184
rect 25006 -14270 25510 -14184
rect 25606 -14270 26110 -14184
rect 26206 -14270 26710 -14184
rect 26806 -14270 27310 -14184
rect 27406 -14270 27910 -14184
rect 28006 -14270 28510 -14184
rect 28606 -14270 29110 -14184
rect 29206 -14270 29710 -14184
rect 29806 -14270 30310 -14184
rect 30406 -14270 30910 -14184
rect 31006 -14270 31510 -14184
rect 31606 -14270 32110 -14184
rect 32206 -14270 32530 -14184
rect 32626 -14270 32652 -14184
rect 24296 -14280 32652 -14270
rect 19072 -18542 22700 -18408
rect 19072 -18914 19709 -18542
rect 19773 -18544 22700 -18542
rect 19773 -18914 20428 -18544
rect 20492 -18914 21147 -18544
rect 21211 -18914 21866 -18544
rect 21930 -18914 22585 -18544
rect 22649 -18914 22700 -18544
rect 19072 -19244 22700 -18914
rect 19072 -19612 19709 -19244
rect 19773 -19612 20428 -19244
rect 20492 -19612 21147 -19244
rect 21211 -19612 21866 -19244
rect 21930 -19612 22585 -19244
rect 22649 -19612 22700 -19244
rect 18872 -19729 18972 -19728
rect 18867 -19827 18873 -19729
rect 18971 -19827 18977 -19729
rect 18872 -19828 18972 -19827
rect 19072 -19944 22700 -19612
rect 34072 -18542 37700 -18408
rect 34072 -18914 34709 -18542
rect 34773 -18544 37700 -18542
rect 34773 -18914 35428 -18544
rect 35492 -18914 36147 -18544
rect 36211 -18914 36866 -18544
rect 36930 -18914 37585 -18544
rect 37649 -18914 37700 -18544
rect 34072 -19244 37700 -18914
rect 34072 -19612 34709 -19244
rect 34773 -19612 35428 -19244
rect 35492 -19612 36147 -19244
rect 36211 -19612 36866 -19244
rect 36930 -19612 37585 -19244
rect 37649 -19612 37700 -19244
rect 22936 -19729 23036 -19728
rect 33872 -19729 33972 -19728
rect 22931 -19827 22937 -19729
rect 23035 -19827 23041 -19729
rect 33867 -19827 33873 -19729
rect 33971 -19827 33977 -19729
rect 22936 -19828 23036 -19827
rect 33872 -19828 33972 -19827
rect 19072 -20312 19709 -19944
rect 19773 -20312 20428 -19944
rect 20492 -20312 21147 -19944
rect 21211 -20312 21866 -19944
rect 21930 -20312 22585 -19944
rect 22649 -20312 22700 -19944
rect 19072 -20644 22700 -20312
rect 19072 -21012 19709 -20644
rect 19773 -21012 20428 -20644
rect 20492 -21012 21147 -20644
rect 21211 -21012 21866 -20644
rect 21930 -21012 22585 -20644
rect 22649 -21012 22700 -20644
rect 19072 -21344 22700 -21012
rect 8694 -21478 18464 -21450
rect 8694 -21564 8744 -21478
rect 8840 -21564 9324 -21478
rect 9420 -21564 9924 -21478
rect 10020 -21564 10524 -21478
rect 10620 -21564 11124 -21478
rect 11220 -21564 11724 -21478
rect 11820 -21564 12324 -21478
rect 12420 -21564 12924 -21478
rect 13020 -21564 13524 -21478
rect 13620 -21564 14124 -21478
rect 14220 -21564 14724 -21478
rect 14820 -21564 15324 -21478
rect 15420 -21564 15924 -21478
rect 16020 -21564 16524 -21478
rect 16620 -21564 17124 -21478
rect 17220 -21564 17724 -21478
rect 17820 -21564 18324 -21478
rect 18420 -21564 18464 -21478
rect 8694 -21594 18464 -21564
rect 19072 -21712 19709 -21344
rect 19773 -21712 20428 -21344
rect 20492 -21712 21147 -21344
rect 21211 -21712 21866 -21344
rect 21930 -21712 22585 -21344
rect 22649 -21712 22700 -21344
rect 34072 -19944 37700 -19612
rect 37834 -19729 37934 -19728
rect 37829 -19827 37835 -19729
rect 37933 -19827 37939 -19729
rect 37834 -19828 37934 -19827
rect 34072 -20312 34709 -19944
rect 34773 -20312 35428 -19944
rect 35492 -20312 36147 -19944
rect 36211 -20312 36866 -19944
rect 36930 -20312 37585 -19944
rect 37649 -20312 37700 -19944
rect 34072 -20644 37700 -20312
rect 34072 -21012 34709 -20644
rect 34773 -21012 35428 -20644
rect 35492 -21012 36147 -20644
rect 36211 -21012 36866 -20644
rect 36930 -21012 37585 -20644
rect 37649 -21012 37700 -20644
rect 34072 -21344 37700 -21012
rect 23694 -21478 33464 -21450
rect 23694 -21564 23744 -21478
rect 23840 -21564 24324 -21478
rect 24420 -21564 24924 -21478
rect 25020 -21564 25524 -21478
rect 25620 -21564 26124 -21478
rect 26220 -21564 26724 -21478
rect 26820 -21564 27324 -21478
rect 27420 -21564 27924 -21478
rect 28020 -21564 28524 -21478
rect 28620 -21564 29124 -21478
rect 29220 -21564 29724 -21478
rect 29820 -21564 30324 -21478
rect 30420 -21564 30924 -21478
rect 31020 -21564 31524 -21478
rect 31620 -21564 32124 -21478
rect 32220 -21564 32724 -21478
rect 32820 -21564 33324 -21478
rect 33420 -21564 33464 -21478
rect 23694 -21594 33464 -21564
rect 8448 -21742 9068 -21737
rect 8448 -22042 8458 -21742
rect 9058 -22042 9068 -21742
rect 8448 -22047 9068 -22042
rect 18080 -21742 18700 -21737
rect 18080 -22042 18090 -21742
rect 18690 -22042 18700 -21742
rect 19072 -21862 22700 -21712
rect 34072 -21712 34709 -21344
rect 34773 -21712 35428 -21344
rect 35492 -21712 36147 -21344
rect 36211 -21712 36866 -21344
rect 36930 -21712 37585 -21344
rect 37649 -21712 37700 -21344
rect 23448 -21742 24068 -21737
rect 18080 -22047 18700 -22042
rect 23448 -22042 23458 -21742
rect 24058 -22042 24068 -21742
rect 23448 -22047 24068 -22042
rect 33080 -21742 33700 -21737
rect 33080 -22042 33090 -21742
rect 33690 -22042 33700 -21742
rect 34072 -21862 37700 -21712
rect 33080 -22047 33700 -22042
<< via3 >>
rect 23440 17094 24040 17394
rect 32072 17094 32672 17394
rect 23562 16868 32558 16978
rect 24176 11572 32038 11716
rect 23440 11162 24040 11462
rect 32072 11162 32672 11462
rect 13066 10328 13448 10628
rect 21200 10328 21878 10628
rect 23648 10328 24248 10628
rect 28280 10328 28880 10628
rect 15134 10064 15230 10150
rect 15714 10064 15810 10150
rect 16314 10064 16410 10150
rect 16914 10064 17010 10150
rect 17514 10064 17610 10150
rect 18114 10064 18210 10150
rect 18714 10064 18810 10150
rect 19314 10064 19410 10150
rect 19914 10064 20010 10150
rect 23896 10064 23992 10150
rect 24476 10064 24572 10150
rect 25076 10064 25172 10150
rect 25676 10064 25772 10150
rect 26276 10064 26372 10150
rect 26876 10064 26972 10150
rect 27476 10064 27572 10150
rect 28076 10064 28172 10150
rect 28676 10064 28772 10150
rect 33086 8924 33182 8996
rect 30406 8380 30502 8452
rect 35784 8380 35880 8452
rect 33086 7836 33182 7908
rect 30406 7292 30502 7364
rect 35784 7292 35880 7364
rect 33086 6748 33182 6820
rect 30406 6204 30502 6276
rect 35784 6204 35880 6276
rect 33086 5660 33182 5732
rect 13066 4872 13448 5172
rect 21200 4872 21878 5172
rect 23648 4872 24248 5172
rect 28280 4872 28880 5172
rect 8458 3990 9058 4290
rect 18090 3990 18690 4290
rect 23458 3990 24058 4290
rect 33090 3990 33690 4290
rect 9310 3730 9406 3816
rect 9910 3730 10006 3816
rect 10510 3730 10606 3816
rect 11110 3730 11206 3816
rect 11710 3730 11806 3816
rect 12310 3730 12406 3816
rect 12910 3730 13006 3816
rect 13510 3730 13606 3816
rect 14110 3730 14206 3816
rect 14710 3730 14806 3816
rect 15310 3730 15406 3816
rect 15910 3730 16006 3816
rect 16510 3730 16606 3816
rect 17110 3730 17206 3816
rect 17530 3730 17626 3816
rect 24310 3730 24406 3816
rect 24910 3730 25006 3816
rect 25510 3730 25606 3816
rect 26110 3730 26206 3816
rect 26710 3730 26806 3816
rect 27310 3730 27406 3816
rect 27910 3730 28006 3816
rect 28510 3730 28606 3816
rect 29110 3730 29206 3816
rect 29710 3730 29806 3816
rect 30310 3730 30406 3816
rect 30910 3730 31006 3816
rect 31510 3730 31606 3816
rect 32110 3730 32206 3816
rect 32530 3730 32626 3816
rect 19709 -914 19773 -542
rect 20428 -914 20492 -544
rect 21147 -914 21211 -544
rect 21866 -914 21930 -544
rect 22585 -914 22649 -544
rect 19709 -1612 19773 -1244
rect 20428 -1612 20492 -1244
rect 21147 -1612 21211 -1244
rect 21866 -1612 21930 -1244
rect 22585 -1612 22649 -1244
rect 34709 -914 34773 -542
rect 35428 -914 35492 -544
rect 36147 -914 36211 -544
rect 36866 -914 36930 -544
rect 37585 -914 37649 -544
rect 18873 -1733 18971 -1729
rect 18873 -1823 18877 -1733
rect 18877 -1823 18967 -1733
rect 18967 -1823 18971 -1733
rect 18873 -1827 18971 -1823
rect 22807 -1827 22905 -1729
rect 19709 -2312 19773 -1944
rect 20428 -2312 20492 -1944
rect 21147 -2312 21211 -1944
rect 21866 -2312 21930 -1944
rect 22585 -2312 22649 -1944
rect 19709 -3012 19773 -2644
rect 20428 -3012 20492 -2644
rect 21147 -3012 21211 -2644
rect 21866 -3012 21930 -2644
rect 22585 -3012 22649 -2644
rect 8744 -3564 8840 -3478
rect 9324 -3564 9420 -3478
rect 9924 -3564 10020 -3478
rect 10524 -3564 10620 -3478
rect 11124 -3564 11220 -3478
rect 11724 -3564 11820 -3478
rect 12324 -3564 12420 -3478
rect 12924 -3564 13020 -3478
rect 13524 -3564 13620 -3478
rect 14124 -3564 14220 -3478
rect 14724 -3564 14820 -3478
rect 15324 -3564 15420 -3478
rect 15924 -3564 16020 -3478
rect 16524 -3564 16620 -3478
rect 17124 -3564 17220 -3478
rect 17724 -3564 17820 -3478
rect 18324 -3564 18420 -3478
rect 19709 -3712 19773 -3344
rect 20428 -3712 20492 -3344
rect 21147 -3712 21211 -3344
rect 21866 -3712 21930 -3344
rect 22585 -3712 22649 -3344
rect 8458 -4042 9058 -3742
rect 18090 -4042 18690 -3742
rect 12412 -5014 13012 -4714
rect 22044 -5014 22644 -4714
rect 8453 -5412 8517 -5044
rect 9172 -5412 9236 -5044
rect 9891 -5412 9955 -5044
rect 10610 -5412 10674 -5044
rect 11329 -5412 11393 -5044
rect 12682 -5278 12778 -5192
rect 13282 -5278 13378 -5192
rect 13882 -5278 13978 -5192
rect 14482 -5278 14578 -5192
rect 15082 -5278 15178 -5192
rect 15682 -5278 15778 -5192
rect 16282 -5278 16378 -5192
rect 16882 -5278 16978 -5192
rect 17482 -5278 17578 -5192
rect 18082 -5278 18178 -5192
rect 18682 -5278 18778 -5192
rect 19282 -5278 19378 -5192
rect 19882 -5278 19978 -5192
rect 20482 -5278 20578 -5192
rect 21082 -5278 21178 -5192
rect 21682 -5278 21778 -5192
rect 22262 -5278 22358 -5192
rect 8453 -6112 8517 -5744
rect 9172 -6112 9236 -5744
rect 9891 -6112 9955 -5744
rect 10610 -6112 10674 -5744
rect 11329 -6112 11393 -5744
rect 8453 -6812 8517 -6444
rect 9172 -6812 9236 -6444
rect 9891 -6812 9955 -6444
rect 10610 -6812 10674 -6444
rect 11329 -6812 11393 -6444
rect 8139 -6933 8237 -6929
rect 8139 -7023 8143 -6933
rect 8143 -7023 8233 -6933
rect 8233 -7023 8237 -6933
rect 8139 -7027 8237 -7023
rect 12131 -6933 12229 -6929
rect 12131 -7023 12135 -6933
rect 12135 -7023 12225 -6933
rect 12225 -7023 12229 -6933
rect 12131 -7027 12229 -7023
rect 8453 -7512 8517 -7144
rect 9172 -7512 9236 -7144
rect 9891 -7512 9955 -7144
rect 10610 -7512 10674 -7144
rect 11329 -7512 11393 -7144
rect 34709 -1612 34773 -1244
rect 35428 -1612 35492 -1244
rect 36147 -1612 36211 -1244
rect 36866 -1612 36930 -1244
rect 37585 -1612 37649 -1244
rect 33873 -1733 33971 -1729
rect 33873 -1823 33877 -1733
rect 33877 -1823 33967 -1733
rect 33967 -1823 33971 -1733
rect 33873 -1827 33971 -1823
rect 34709 -2312 34773 -1944
rect 35428 -2312 35492 -1944
rect 36147 -2312 36211 -1944
rect 36866 -2312 36930 -1944
rect 37585 -2312 37649 -1944
rect 34709 -3012 34773 -2644
rect 35428 -3012 35492 -2644
rect 36147 -3012 36211 -2644
rect 36866 -3012 36930 -2644
rect 37585 -3012 37649 -2644
rect 23744 -3564 23840 -3478
rect 24324 -3564 24420 -3478
rect 24924 -3564 25020 -3478
rect 25524 -3564 25620 -3478
rect 26124 -3564 26220 -3478
rect 26724 -3564 26820 -3478
rect 27324 -3564 27420 -3478
rect 27924 -3564 28020 -3478
rect 28524 -3564 28620 -3478
rect 29124 -3564 29220 -3478
rect 29724 -3564 29820 -3478
rect 30324 -3564 30420 -3478
rect 30924 -3564 31020 -3478
rect 31524 -3564 31620 -3478
rect 32124 -3564 32220 -3478
rect 32724 -3564 32820 -3478
rect 33324 -3564 33420 -3478
rect 34709 -3712 34773 -3344
rect 35428 -3712 35492 -3344
rect 36147 -3712 36211 -3344
rect 36866 -3712 36930 -3344
rect 37585 -3712 37649 -3344
rect 23458 -4042 24058 -3742
rect 33090 -4042 33690 -3742
rect 27412 -5014 28012 -4714
rect 37044 -5014 37644 -4714
rect 23453 -5412 23517 -5044
rect 24172 -5412 24236 -5044
rect 24891 -5412 24955 -5044
rect 25610 -5412 25674 -5044
rect 26329 -5412 26393 -5044
rect 27682 -5278 27778 -5192
rect 28282 -5278 28378 -5192
rect 28882 -5278 28978 -5192
rect 29482 -5278 29578 -5192
rect 30082 -5278 30178 -5192
rect 30682 -5278 30778 -5192
rect 31282 -5278 31378 -5192
rect 31882 -5278 31978 -5192
rect 32482 -5278 32578 -5192
rect 33082 -5278 33178 -5192
rect 33682 -5278 33778 -5192
rect 34282 -5278 34378 -5192
rect 34882 -5278 34978 -5192
rect 35482 -5278 35578 -5192
rect 36082 -5278 36178 -5192
rect 36682 -5278 36778 -5192
rect 37262 -5278 37358 -5192
rect 23453 -6112 23517 -5744
rect 24172 -6112 24236 -5744
rect 24891 -6112 24955 -5744
rect 25610 -6112 25674 -5744
rect 26329 -6112 26393 -5744
rect 23453 -6812 23517 -6444
rect 24172 -6812 24236 -6444
rect 24891 -6812 24955 -6444
rect 25610 -6812 25674 -6444
rect 26329 -6812 26393 -6444
rect 23131 -7027 23229 -6929
rect 27131 -6933 27229 -6929
rect 27131 -7023 27135 -6933
rect 27135 -7023 27225 -6933
rect 27225 -7023 27229 -6933
rect 27131 -7027 27229 -7023
rect 8453 -8212 8517 -7842
rect 9172 -8212 9236 -7842
rect 9891 -8212 9955 -7842
rect 10610 -8212 10674 -7842
rect 11329 -8214 11393 -7842
rect 23453 -7512 23517 -7144
rect 24172 -7512 24236 -7144
rect 24891 -7512 24955 -7144
rect 25610 -7512 25674 -7144
rect 26329 -7512 26393 -7144
rect 23453 -8212 23517 -7842
rect 24172 -8212 24236 -7842
rect 24891 -8212 24955 -7842
rect 25610 -8212 25674 -7842
rect 26329 -8214 26393 -7842
rect 13476 -12572 13572 -12486
rect 13896 -12572 13992 -12486
rect 14496 -12572 14592 -12486
rect 15096 -12572 15192 -12486
rect 15696 -12572 15792 -12486
rect 16296 -12572 16392 -12486
rect 16896 -12572 16992 -12486
rect 17496 -12572 17592 -12486
rect 18096 -12572 18192 -12486
rect 18696 -12572 18792 -12486
rect 19296 -12572 19392 -12486
rect 19896 -12572 19992 -12486
rect 20496 -12572 20592 -12486
rect 21096 -12572 21192 -12486
rect 21696 -12572 21792 -12486
rect 28476 -12572 28572 -12486
rect 28896 -12572 28992 -12486
rect 29496 -12572 29592 -12486
rect 30096 -12572 30192 -12486
rect 30696 -12572 30792 -12486
rect 31296 -12572 31392 -12486
rect 31896 -12572 31992 -12486
rect 32496 -12572 32592 -12486
rect 33096 -12572 33192 -12486
rect 33696 -12572 33792 -12486
rect 34296 -12572 34392 -12486
rect 34896 -12572 34992 -12486
rect 35496 -12572 35592 -12486
rect 36096 -12572 36192 -12486
rect 36696 -12572 36792 -12486
rect 12412 -13046 13012 -12746
rect 22044 -13046 22644 -12746
rect 27412 -13046 28012 -12746
rect 37044 -13046 37644 -12746
rect 8458 -14010 9058 -13710
rect 18090 -14010 18690 -13710
rect 23458 -14010 24058 -13710
rect 33090 -14010 33690 -13710
rect 9310 -14270 9406 -14184
rect 9910 -14270 10006 -14184
rect 10510 -14270 10606 -14184
rect 11110 -14270 11206 -14184
rect 11710 -14270 11806 -14184
rect 12310 -14270 12406 -14184
rect 12910 -14270 13006 -14184
rect 13510 -14270 13606 -14184
rect 14110 -14270 14206 -14184
rect 14710 -14270 14806 -14184
rect 15310 -14270 15406 -14184
rect 15910 -14270 16006 -14184
rect 16510 -14270 16606 -14184
rect 17110 -14270 17206 -14184
rect 17530 -14270 17626 -14184
rect 24310 -14270 24406 -14184
rect 24910 -14270 25006 -14184
rect 25510 -14270 25606 -14184
rect 26110 -14270 26206 -14184
rect 26710 -14270 26806 -14184
rect 27310 -14270 27406 -14184
rect 27910 -14270 28006 -14184
rect 28510 -14270 28606 -14184
rect 29110 -14270 29206 -14184
rect 29710 -14270 29806 -14184
rect 30310 -14270 30406 -14184
rect 30910 -14270 31006 -14184
rect 31510 -14270 31606 -14184
rect 32110 -14270 32206 -14184
rect 32530 -14270 32626 -14184
rect 19709 -18914 19773 -18542
rect 20428 -18914 20492 -18544
rect 21147 -18914 21211 -18544
rect 21866 -18914 21930 -18544
rect 22585 -18914 22649 -18544
rect 19709 -19612 19773 -19244
rect 20428 -19612 20492 -19244
rect 21147 -19612 21211 -19244
rect 21866 -19612 21930 -19244
rect 22585 -19612 22649 -19244
rect 18873 -19733 18971 -19729
rect 18873 -19823 18877 -19733
rect 18877 -19823 18967 -19733
rect 18967 -19823 18971 -19733
rect 18873 -19827 18971 -19823
rect 34709 -18914 34773 -18542
rect 35428 -18914 35492 -18544
rect 36147 -18914 36211 -18544
rect 36866 -18914 36930 -18544
rect 37585 -18914 37649 -18544
rect 34709 -19612 34773 -19244
rect 35428 -19612 35492 -19244
rect 36147 -19612 36211 -19244
rect 36866 -19612 36930 -19244
rect 37585 -19612 37649 -19244
rect 22937 -19733 23035 -19729
rect 22937 -19823 22941 -19733
rect 22941 -19823 23031 -19733
rect 23031 -19823 23035 -19733
rect 22937 -19827 23035 -19823
rect 33873 -19733 33971 -19729
rect 33873 -19823 33877 -19733
rect 33877 -19823 33967 -19733
rect 33967 -19823 33971 -19733
rect 33873 -19827 33971 -19823
rect 19709 -20312 19773 -19944
rect 20428 -20312 20492 -19944
rect 21147 -20312 21211 -19944
rect 21866 -20312 21930 -19944
rect 22585 -20312 22649 -19944
rect 19709 -21012 19773 -20644
rect 20428 -21012 20492 -20644
rect 21147 -21012 21211 -20644
rect 21866 -21012 21930 -20644
rect 22585 -21012 22649 -20644
rect 8744 -21564 8840 -21478
rect 9324 -21564 9420 -21478
rect 9924 -21564 10020 -21478
rect 10524 -21564 10620 -21478
rect 11124 -21564 11220 -21478
rect 11724 -21564 11820 -21478
rect 12324 -21564 12420 -21478
rect 12924 -21564 13020 -21478
rect 13524 -21564 13620 -21478
rect 14124 -21564 14220 -21478
rect 14724 -21564 14820 -21478
rect 15324 -21564 15420 -21478
rect 15924 -21564 16020 -21478
rect 16524 -21564 16620 -21478
rect 17124 -21564 17220 -21478
rect 17724 -21564 17820 -21478
rect 18324 -21564 18420 -21478
rect 19709 -21712 19773 -21344
rect 20428 -21712 20492 -21344
rect 21147 -21712 21211 -21344
rect 21866 -21712 21930 -21344
rect 22585 -21712 22649 -21344
rect 37835 -19733 37933 -19729
rect 37835 -19823 37839 -19733
rect 37839 -19823 37929 -19733
rect 37929 -19823 37933 -19733
rect 37835 -19827 37933 -19823
rect 34709 -20312 34773 -19944
rect 35428 -20312 35492 -19944
rect 36147 -20312 36211 -19944
rect 36866 -20312 36930 -19944
rect 37585 -20312 37649 -19944
rect 34709 -21012 34773 -20644
rect 35428 -21012 35492 -20644
rect 36147 -21012 36211 -20644
rect 36866 -21012 36930 -20644
rect 37585 -21012 37649 -20644
rect 23744 -21564 23840 -21478
rect 24324 -21564 24420 -21478
rect 24924 -21564 25020 -21478
rect 25524 -21564 25620 -21478
rect 26124 -21564 26220 -21478
rect 26724 -21564 26820 -21478
rect 27324 -21564 27420 -21478
rect 27924 -21564 28020 -21478
rect 28524 -21564 28620 -21478
rect 29124 -21564 29220 -21478
rect 29724 -21564 29820 -21478
rect 30324 -21564 30420 -21478
rect 30924 -21564 31020 -21478
rect 31524 -21564 31620 -21478
rect 32124 -21564 32220 -21478
rect 32724 -21564 32820 -21478
rect 33324 -21564 33420 -21478
rect 8458 -22042 9058 -21742
rect 18090 -22042 18690 -21742
rect 34709 -21712 34773 -21344
rect 35428 -21712 35492 -21344
rect 36147 -21712 36211 -21344
rect 36866 -21712 36930 -21344
rect 37585 -21712 37649 -21344
rect 23458 -22042 24058 -21742
rect 33090 -22042 33690 -21742
<< mimcap >>
rect 19194 -566 19594 -526
rect 19194 -886 19234 -566
rect 19554 -886 19594 -566
rect 19194 -926 19594 -886
rect 19913 -566 20313 -526
rect 19913 -886 19953 -566
rect 20273 -886 20313 -566
rect 19913 -926 20313 -886
rect 20632 -566 21032 -526
rect 20632 -886 20672 -566
rect 20992 -886 21032 -566
rect 20632 -926 21032 -886
rect 21351 -566 21751 -526
rect 21351 -886 21391 -566
rect 21711 -886 21751 -566
rect 21351 -926 21751 -886
rect 22070 -566 22470 -526
rect 22070 -886 22110 -566
rect 22430 -886 22470 -566
rect 22070 -926 22470 -886
rect 34194 -566 34594 -526
rect 34194 -886 34234 -566
rect 34554 -886 34594 -566
rect 34194 -926 34594 -886
rect 34913 -566 35313 -526
rect 34913 -886 34953 -566
rect 35273 -886 35313 -566
rect 34913 -926 35313 -886
rect 35632 -566 36032 -526
rect 35632 -886 35672 -566
rect 35992 -886 36032 -566
rect 35632 -926 36032 -886
rect 36351 -566 36751 -526
rect 36351 -886 36391 -566
rect 36711 -886 36751 -566
rect 36351 -926 36751 -886
rect 37070 -566 37470 -526
rect 37070 -886 37110 -566
rect 37430 -886 37470 -566
rect 37070 -926 37470 -886
rect 19194 -1266 19594 -1226
rect 19194 -1586 19234 -1266
rect 19554 -1586 19594 -1266
rect 19194 -1626 19594 -1586
rect 19913 -1266 20313 -1226
rect 19913 -1586 19953 -1266
rect 20273 -1586 20313 -1266
rect 19913 -1626 20313 -1586
rect 20632 -1266 21032 -1226
rect 20632 -1586 20672 -1266
rect 20992 -1586 21032 -1266
rect 20632 -1626 21032 -1586
rect 21351 -1266 21751 -1226
rect 21351 -1586 21391 -1266
rect 21711 -1586 21751 -1266
rect 21351 -1626 21751 -1586
rect 22070 -1266 22470 -1226
rect 22070 -1586 22110 -1266
rect 22430 -1586 22470 -1266
rect 22070 -1626 22470 -1586
rect 34194 -1266 34594 -1226
rect 34194 -1586 34234 -1266
rect 34554 -1586 34594 -1266
rect 34194 -1626 34594 -1586
rect 34913 -1266 35313 -1226
rect 34913 -1586 34953 -1266
rect 35273 -1586 35313 -1266
rect 34913 -1626 35313 -1586
rect 35632 -1266 36032 -1226
rect 35632 -1586 35672 -1266
rect 35992 -1586 36032 -1266
rect 35632 -1626 36032 -1586
rect 36351 -1266 36751 -1226
rect 36351 -1586 36391 -1266
rect 36711 -1586 36751 -1266
rect 36351 -1626 36751 -1586
rect 37070 -1266 37470 -1226
rect 37070 -1586 37110 -1266
rect 37430 -1586 37470 -1266
rect 37070 -1626 37470 -1586
rect 19194 -1966 19594 -1926
rect 19194 -2286 19234 -1966
rect 19554 -2286 19594 -1966
rect 19194 -2326 19594 -2286
rect 19913 -1966 20313 -1926
rect 19913 -2286 19953 -1966
rect 20273 -2286 20313 -1966
rect 19913 -2326 20313 -2286
rect 20632 -1966 21032 -1926
rect 20632 -2286 20672 -1966
rect 20992 -2286 21032 -1966
rect 20632 -2326 21032 -2286
rect 21351 -1966 21751 -1926
rect 21351 -2286 21391 -1966
rect 21711 -2286 21751 -1966
rect 21351 -2326 21751 -2286
rect 22070 -1966 22470 -1926
rect 22070 -2286 22110 -1966
rect 22430 -2286 22470 -1966
rect 22070 -2326 22470 -2286
rect 34194 -1966 34594 -1926
rect 34194 -2286 34234 -1966
rect 34554 -2286 34594 -1966
rect 34194 -2326 34594 -2286
rect 34913 -1966 35313 -1926
rect 34913 -2286 34953 -1966
rect 35273 -2286 35313 -1966
rect 34913 -2326 35313 -2286
rect 35632 -1966 36032 -1926
rect 35632 -2286 35672 -1966
rect 35992 -2286 36032 -1966
rect 35632 -2326 36032 -2286
rect 36351 -1966 36751 -1926
rect 36351 -2286 36391 -1966
rect 36711 -2286 36751 -1966
rect 36351 -2326 36751 -2286
rect 37070 -1966 37470 -1926
rect 37070 -2286 37110 -1966
rect 37430 -2286 37470 -1966
rect 37070 -2326 37470 -2286
rect 19194 -2666 19594 -2626
rect 19194 -2986 19234 -2666
rect 19554 -2986 19594 -2666
rect 19194 -3026 19594 -2986
rect 19913 -2666 20313 -2626
rect 19913 -2986 19953 -2666
rect 20273 -2986 20313 -2666
rect 19913 -3026 20313 -2986
rect 20632 -2666 21032 -2626
rect 20632 -2986 20672 -2666
rect 20992 -2986 21032 -2666
rect 20632 -3026 21032 -2986
rect 21351 -2666 21751 -2626
rect 21351 -2986 21391 -2666
rect 21711 -2986 21751 -2666
rect 21351 -3026 21751 -2986
rect 22070 -2666 22470 -2626
rect 22070 -2986 22110 -2666
rect 22430 -2986 22470 -2666
rect 22070 -3026 22470 -2986
rect 34194 -2666 34594 -2626
rect 34194 -2986 34234 -2666
rect 34554 -2986 34594 -2666
rect 34194 -3026 34594 -2986
rect 34913 -2666 35313 -2626
rect 34913 -2986 34953 -2666
rect 35273 -2986 35313 -2666
rect 34913 -3026 35313 -2986
rect 35632 -2666 36032 -2626
rect 35632 -2986 35672 -2666
rect 35992 -2986 36032 -2666
rect 35632 -3026 36032 -2986
rect 36351 -2666 36751 -2626
rect 36351 -2986 36391 -2666
rect 36711 -2986 36751 -2666
rect 36351 -3026 36751 -2986
rect 37070 -2666 37470 -2626
rect 37070 -2986 37110 -2666
rect 37430 -2986 37470 -2666
rect 37070 -3026 37470 -2986
rect 19194 -3366 19594 -3326
rect 19194 -3686 19234 -3366
rect 19554 -3686 19594 -3366
rect 19194 -3726 19594 -3686
rect 19913 -3366 20313 -3326
rect 19913 -3686 19953 -3366
rect 20273 -3686 20313 -3366
rect 19913 -3726 20313 -3686
rect 20632 -3366 21032 -3326
rect 20632 -3686 20672 -3366
rect 20992 -3686 21032 -3366
rect 20632 -3726 21032 -3686
rect 21351 -3366 21751 -3326
rect 21351 -3686 21391 -3366
rect 21711 -3686 21751 -3366
rect 21351 -3726 21751 -3686
rect 22070 -3366 22470 -3326
rect 22070 -3686 22110 -3366
rect 22430 -3686 22470 -3366
rect 22070 -3726 22470 -3686
rect 34194 -3366 34594 -3326
rect 34194 -3686 34234 -3366
rect 34554 -3686 34594 -3366
rect 34194 -3726 34594 -3686
rect 34913 -3366 35313 -3326
rect 34913 -3686 34953 -3366
rect 35273 -3686 35313 -3366
rect 34913 -3726 35313 -3686
rect 35632 -3366 36032 -3326
rect 35632 -3686 35672 -3366
rect 35992 -3686 36032 -3366
rect 35632 -3726 36032 -3686
rect 36351 -3366 36751 -3326
rect 36351 -3686 36391 -3366
rect 36711 -3686 36751 -3366
rect 36351 -3726 36751 -3686
rect 37070 -3366 37470 -3326
rect 37070 -3686 37110 -3366
rect 37430 -3686 37470 -3366
rect 37070 -3726 37470 -3686
rect 8632 -5070 9032 -5030
rect 8632 -5390 8672 -5070
rect 8992 -5390 9032 -5070
rect 8632 -5430 9032 -5390
rect 9351 -5070 9751 -5030
rect 9351 -5390 9391 -5070
rect 9711 -5390 9751 -5070
rect 9351 -5430 9751 -5390
rect 10070 -5070 10470 -5030
rect 10070 -5390 10110 -5070
rect 10430 -5390 10470 -5070
rect 10070 -5430 10470 -5390
rect 10789 -5070 11189 -5030
rect 10789 -5390 10829 -5070
rect 11149 -5390 11189 -5070
rect 10789 -5430 11189 -5390
rect 11508 -5070 11908 -5030
rect 11508 -5390 11548 -5070
rect 11868 -5390 11908 -5070
rect 11508 -5430 11908 -5390
rect 23632 -5070 24032 -5030
rect 23632 -5390 23672 -5070
rect 23992 -5390 24032 -5070
rect 23632 -5430 24032 -5390
rect 24351 -5070 24751 -5030
rect 24351 -5390 24391 -5070
rect 24711 -5390 24751 -5070
rect 24351 -5430 24751 -5390
rect 25070 -5070 25470 -5030
rect 25070 -5390 25110 -5070
rect 25430 -5390 25470 -5070
rect 25070 -5430 25470 -5390
rect 25789 -5070 26189 -5030
rect 25789 -5390 25829 -5070
rect 26149 -5390 26189 -5070
rect 25789 -5430 26189 -5390
rect 26508 -5070 26908 -5030
rect 26508 -5390 26548 -5070
rect 26868 -5390 26908 -5070
rect 26508 -5430 26908 -5390
rect 8632 -5770 9032 -5730
rect 8632 -6090 8672 -5770
rect 8992 -6090 9032 -5770
rect 8632 -6130 9032 -6090
rect 9351 -5770 9751 -5730
rect 9351 -6090 9391 -5770
rect 9711 -6090 9751 -5770
rect 9351 -6130 9751 -6090
rect 10070 -5770 10470 -5730
rect 10070 -6090 10110 -5770
rect 10430 -6090 10470 -5770
rect 10070 -6130 10470 -6090
rect 10789 -5770 11189 -5730
rect 10789 -6090 10829 -5770
rect 11149 -6090 11189 -5770
rect 10789 -6130 11189 -6090
rect 11508 -5770 11908 -5730
rect 11508 -6090 11548 -5770
rect 11868 -6090 11908 -5770
rect 11508 -6130 11908 -6090
rect 23632 -5770 24032 -5730
rect 23632 -6090 23672 -5770
rect 23992 -6090 24032 -5770
rect 23632 -6130 24032 -6090
rect 24351 -5770 24751 -5730
rect 24351 -6090 24391 -5770
rect 24711 -6090 24751 -5770
rect 24351 -6130 24751 -6090
rect 25070 -5770 25470 -5730
rect 25070 -6090 25110 -5770
rect 25430 -6090 25470 -5770
rect 25070 -6130 25470 -6090
rect 25789 -5770 26189 -5730
rect 25789 -6090 25829 -5770
rect 26149 -6090 26189 -5770
rect 25789 -6130 26189 -6090
rect 26508 -5770 26908 -5730
rect 26508 -6090 26548 -5770
rect 26868 -6090 26908 -5770
rect 26508 -6130 26908 -6090
rect 8632 -6470 9032 -6430
rect 8632 -6790 8672 -6470
rect 8992 -6790 9032 -6470
rect 8632 -6830 9032 -6790
rect 9351 -6470 9751 -6430
rect 9351 -6790 9391 -6470
rect 9711 -6790 9751 -6470
rect 9351 -6830 9751 -6790
rect 10070 -6470 10470 -6430
rect 10070 -6790 10110 -6470
rect 10430 -6790 10470 -6470
rect 10070 -6830 10470 -6790
rect 10789 -6470 11189 -6430
rect 10789 -6790 10829 -6470
rect 11149 -6790 11189 -6470
rect 10789 -6830 11189 -6790
rect 11508 -6470 11908 -6430
rect 11508 -6790 11548 -6470
rect 11868 -6790 11908 -6470
rect 11508 -6830 11908 -6790
rect 23632 -6470 24032 -6430
rect 23632 -6790 23672 -6470
rect 23992 -6790 24032 -6470
rect 23632 -6830 24032 -6790
rect 24351 -6470 24751 -6430
rect 24351 -6790 24391 -6470
rect 24711 -6790 24751 -6470
rect 24351 -6830 24751 -6790
rect 25070 -6470 25470 -6430
rect 25070 -6790 25110 -6470
rect 25430 -6790 25470 -6470
rect 25070 -6830 25470 -6790
rect 25789 -6470 26189 -6430
rect 25789 -6790 25829 -6470
rect 26149 -6790 26189 -6470
rect 25789 -6830 26189 -6790
rect 26508 -6470 26908 -6430
rect 26508 -6790 26548 -6470
rect 26868 -6790 26908 -6470
rect 26508 -6830 26908 -6790
rect 8632 -7170 9032 -7130
rect 8632 -7490 8672 -7170
rect 8992 -7490 9032 -7170
rect 8632 -7530 9032 -7490
rect 9351 -7170 9751 -7130
rect 9351 -7490 9391 -7170
rect 9711 -7490 9751 -7170
rect 9351 -7530 9751 -7490
rect 10070 -7170 10470 -7130
rect 10070 -7490 10110 -7170
rect 10430 -7490 10470 -7170
rect 10070 -7530 10470 -7490
rect 10789 -7170 11189 -7130
rect 10789 -7490 10829 -7170
rect 11149 -7490 11189 -7170
rect 10789 -7530 11189 -7490
rect 11508 -7170 11908 -7130
rect 11508 -7490 11548 -7170
rect 11868 -7490 11908 -7170
rect 11508 -7530 11908 -7490
rect 23632 -7170 24032 -7130
rect 23632 -7490 23672 -7170
rect 23992 -7490 24032 -7170
rect 23632 -7530 24032 -7490
rect 24351 -7170 24751 -7130
rect 24351 -7490 24391 -7170
rect 24711 -7490 24751 -7170
rect 24351 -7530 24751 -7490
rect 25070 -7170 25470 -7130
rect 25070 -7490 25110 -7170
rect 25430 -7490 25470 -7170
rect 25070 -7530 25470 -7490
rect 25789 -7170 26189 -7130
rect 25789 -7490 25829 -7170
rect 26149 -7490 26189 -7170
rect 25789 -7530 26189 -7490
rect 26508 -7170 26908 -7130
rect 26508 -7490 26548 -7170
rect 26868 -7490 26908 -7170
rect 26508 -7530 26908 -7490
rect 8632 -7870 9032 -7830
rect 8632 -8190 8672 -7870
rect 8992 -8190 9032 -7870
rect 8632 -8230 9032 -8190
rect 9351 -7870 9751 -7830
rect 9351 -8190 9391 -7870
rect 9711 -8190 9751 -7870
rect 9351 -8230 9751 -8190
rect 10070 -7870 10470 -7830
rect 10070 -8190 10110 -7870
rect 10430 -8190 10470 -7870
rect 10070 -8230 10470 -8190
rect 10789 -7870 11189 -7830
rect 10789 -8190 10829 -7870
rect 11149 -8190 11189 -7870
rect 10789 -8230 11189 -8190
rect 11508 -7870 11908 -7830
rect 11508 -8190 11548 -7870
rect 11868 -8190 11908 -7870
rect 11508 -8230 11908 -8190
rect 23632 -7870 24032 -7830
rect 23632 -8190 23672 -7870
rect 23992 -8190 24032 -7870
rect 23632 -8230 24032 -8190
rect 24351 -7870 24751 -7830
rect 24351 -8190 24391 -7870
rect 24711 -8190 24751 -7870
rect 24351 -8230 24751 -8190
rect 25070 -7870 25470 -7830
rect 25070 -8190 25110 -7870
rect 25430 -8190 25470 -7870
rect 25070 -8230 25470 -8190
rect 25789 -7870 26189 -7830
rect 25789 -8190 25829 -7870
rect 26149 -8190 26189 -7870
rect 25789 -8230 26189 -8190
rect 26508 -7870 26908 -7830
rect 26508 -8190 26548 -7870
rect 26868 -8190 26908 -7870
rect 26508 -8230 26908 -8190
rect 19194 -18566 19594 -18526
rect 19194 -18886 19234 -18566
rect 19554 -18886 19594 -18566
rect 19194 -18926 19594 -18886
rect 19913 -18566 20313 -18526
rect 19913 -18886 19953 -18566
rect 20273 -18886 20313 -18566
rect 19913 -18926 20313 -18886
rect 20632 -18566 21032 -18526
rect 20632 -18886 20672 -18566
rect 20992 -18886 21032 -18566
rect 20632 -18926 21032 -18886
rect 21351 -18566 21751 -18526
rect 21351 -18886 21391 -18566
rect 21711 -18886 21751 -18566
rect 21351 -18926 21751 -18886
rect 22070 -18566 22470 -18526
rect 22070 -18886 22110 -18566
rect 22430 -18886 22470 -18566
rect 22070 -18926 22470 -18886
rect 34194 -18566 34594 -18526
rect 34194 -18886 34234 -18566
rect 34554 -18886 34594 -18566
rect 34194 -18926 34594 -18886
rect 34913 -18566 35313 -18526
rect 34913 -18886 34953 -18566
rect 35273 -18886 35313 -18566
rect 34913 -18926 35313 -18886
rect 35632 -18566 36032 -18526
rect 35632 -18886 35672 -18566
rect 35992 -18886 36032 -18566
rect 35632 -18926 36032 -18886
rect 36351 -18566 36751 -18526
rect 36351 -18886 36391 -18566
rect 36711 -18886 36751 -18566
rect 36351 -18926 36751 -18886
rect 37070 -18566 37470 -18526
rect 37070 -18886 37110 -18566
rect 37430 -18886 37470 -18566
rect 37070 -18926 37470 -18886
rect 19194 -19266 19594 -19226
rect 19194 -19586 19234 -19266
rect 19554 -19586 19594 -19266
rect 19194 -19626 19594 -19586
rect 19913 -19266 20313 -19226
rect 19913 -19586 19953 -19266
rect 20273 -19586 20313 -19266
rect 19913 -19626 20313 -19586
rect 20632 -19266 21032 -19226
rect 20632 -19586 20672 -19266
rect 20992 -19586 21032 -19266
rect 20632 -19626 21032 -19586
rect 21351 -19266 21751 -19226
rect 21351 -19586 21391 -19266
rect 21711 -19586 21751 -19266
rect 21351 -19626 21751 -19586
rect 22070 -19266 22470 -19226
rect 22070 -19586 22110 -19266
rect 22430 -19586 22470 -19266
rect 22070 -19626 22470 -19586
rect 34194 -19266 34594 -19226
rect 34194 -19586 34234 -19266
rect 34554 -19586 34594 -19266
rect 34194 -19626 34594 -19586
rect 34913 -19266 35313 -19226
rect 34913 -19586 34953 -19266
rect 35273 -19586 35313 -19266
rect 34913 -19626 35313 -19586
rect 35632 -19266 36032 -19226
rect 35632 -19586 35672 -19266
rect 35992 -19586 36032 -19266
rect 35632 -19626 36032 -19586
rect 36351 -19266 36751 -19226
rect 36351 -19586 36391 -19266
rect 36711 -19586 36751 -19266
rect 36351 -19626 36751 -19586
rect 37070 -19266 37470 -19226
rect 37070 -19586 37110 -19266
rect 37430 -19586 37470 -19266
rect 37070 -19626 37470 -19586
rect 19194 -19966 19594 -19926
rect 19194 -20286 19234 -19966
rect 19554 -20286 19594 -19966
rect 19194 -20326 19594 -20286
rect 19913 -19966 20313 -19926
rect 19913 -20286 19953 -19966
rect 20273 -20286 20313 -19966
rect 19913 -20326 20313 -20286
rect 20632 -19966 21032 -19926
rect 20632 -20286 20672 -19966
rect 20992 -20286 21032 -19966
rect 20632 -20326 21032 -20286
rect 21351 -19966 21751 -19926
rect 21351 -20286 21391 -19966
rect 21711 -20286 21751 -19966
rect 21351 -20326 21751 -20286
rect 22070 -19966 22470 -19926
rect 22070 -20286 22110 -19966
rect 22430 -20286 22470 -19966
rect 22070 -20326 22470 -20286
rect 34194 -19966 34594 -19926
rect 34194 -20286 34234 -19966
rect 34554 -20286 34594 -19966
rect 34194 -20326 34594 -20286
rect 34913 -19966 35313 -19926
rect 34913 -20286 34953 -19966
rect 35273 -20286 35313 -19966
rect 34913 -20326 35313 -20286
rect 35632 -19966 36032 -19926
rect 35632 -20286 35672 -19966
rect 35992 -20286 36032 -19966
rect 35632 -20326 36032 -20286
rect 36351 -19966 36751 -19926
rect 36351 -20286 36391 -19966
rect 36711 -20286 36751 -19966
rect 36351 -20326 36751 -20286
rect 37070 -19966 37470 -19926
rect 37070 -20286 37110 -19966
rect 37430 -20286 37470 -19966
rect 37070 -20326 37470 -20286
rect 19194 -20666 19594 -20626
rect 19194 -20986 19234 -20666
rect 19554 -20986 19594 -20666
rect 19194 -21026 19594 -20986
rect 19913 -20666 20313 -20626
rect 19913 -20986 19953 -20666
rect 20273 -20986 20313 -20666
rect 19913 -21026 20313 -20986
rect 20632 -20666 21032 -20626
rect 20632 -20986 20672 -20666
rect 20992 -20986 21032 -20666
rect 20632 -21026 21032 -20986
rect 21351 -20666 21751 -20626
rect 21351 -20986 21391 -20666
rect 21711 -20986 21751 -20666
rect 21351 -21026 21751 -20986
rect 22070 -20666 22470 -20626
rect 22070 -20986 22110 -20666
rect 22430 -20986 22470 -20666
rect 22070 -21026 22470 -20986
rect 34194 -20666 34594 -20626
rect 34194 -20986 34234 -20666
rect 34554 -20986 34594 -20666
rect 34194 -21026 34594 -20986
rect 34913 -20666 35313 -20626
rect 34913 -20986 34953 -20666
rect 35273 -20986 35313 -20666
rect 34913 -21026 35313 -20986
rect 35632 -20666 36032 -20626
rect 35632 -20986 35672 -20666
rect 35992 -20986 36032 -20666
rect 35632 -21026 36032 -20986
rect 36351 -20666 36751 -20626
rect 36351 -20986 36391 -20666
rect 36711 -20986 36751 -20666
rect 36351 -21026 36751 -20986
rect 37070 -20666 37470 -20626
rect 37070 -20986 37110 -20666
rect 37430 -20986 37470 -20666
rect 37070 -21026 37470 -20986
rect 19194 -21366 19594 -21326
rect 19194 -21686 19234 -21366
rect 19554 -21686 19594 -21366
rect 19194 -21726 19594 -21686
rect 19913 -21366 20313 -21326
rect 19913 -21686 19953 -21366
rect 20273 -21686 20313 -21366
rect 19913 -21726 20313 -21686
rect 20632 -21366 21032 -21326
rect 20632 -21686 20672 -21366
rect 20992 -21686 21032 -21366
rect 20632 -21726 21032 -21686
rect 21351 -21366 21751 -21326
rect 21351 -21686 21391 -21366
rect 21711 -21686 21751 -21366
rect 21351 -21726 21751 -21686
rect 22070 -21366 22470 -21326
rect 22070 -21686 22110 -21366
rect 22430 -21686 22470 -21366
rect 22070 -21726 22470 -21686
rect 34194 -21366 34594 -21326
rect 34194 -21686 34234 -21366
rect 34554 -21686 34594 -21366
rect 34194 -21726 34594 -21686
rect 34913 -21366 35313 -21326
rect 34913 -21686 34953 -21366
rect 35273 -21686 35313 -21366
rect 34913 -21726 35313 -21686
rect 35632 -21366 36032 -21326
rect 35632 -21686 35672 -21366
rect 35992 -21686 36032 -21366
rect 35632 -21726 36032 -21686
rect 36351 -21366 36751 -21326
rect 36351 -21686 36391 -21366
rect 36711 -21686 36751 -21366
rect 36351 -21726 36751 -21686
rect 37070 -21366 37470 -21326
rect 37070 -21686 37110 -21366
rect 37430 -21686 37470 -21366
rect 37070 -21726 37470 -21686
<< mimcapcontact >>
rect 19234 -886 19554 -566
rect 19953 -886 20273 -566
rect 20672 -886 20992 -566
rect 21391 -886 21711 -566
rect 22110 -886 22430 -566
rect 34234 -886 34554 -566
rect 34953 -886 35273 -566
rect 35672 -886 35992 -566
rect 36391 -886 36711 -566
rect 37110 -886 37430 -566
rect 19234 -1586 19554 -1266
rect 19953 -1586 20273 -1266
rect 20672 -1586 20992 -1266
rect 21391 -1586 21711 -1266
rect 22110 -1586 22430 -1266
rect 34234 -1586 34554 -1266
rect 34953 -1586 35273 -1266
rect 35672 -1586 35992 -1266
rect 36391 -1586 36711 -1266
rect 37110 -1586 37430 -1266
rect 19234 -2286 19554 -1966
rect 19953 -2286 20273 -1966
rect 20672 -2286 20992 -1966
rect 21391 -2286 21711 -1966
rect 22110 -2286 22430 -1966
rect 34234 -2286 34554 -1966
rect 34953 -2286 35273 -1966
rect 35672 -2286 35992 -1966
rect 36391 -2286 36711 -1966
rect 37110 -2286 37430 -1966
rect 19234 -2986 19554 -2666
rect 19953 -2986 20273 -2666
rect 20672 -2986 20992 -2666
rect 21391 -2986 21711 -2666
rect 22110 -2986 22430 -2666
rect 34234 -2986 34554 -2666
rect 34953 -2986 35273 -2666
rect 35672 -2986 35992 -2666
rect 36391 -2986 36711 -2666
rect 37110 -2986 37430 -2666
rect 19234 -3686 19554 -3366
rect 19953 -3686 20273 -3366
rect 20672 -3686 20992 -3366
rect 21391 -3686 21711 -3366
rect 22110 -3686 22430 -3366
rect 34234 -3686 34554 -3366
rect 34953 -3686 35273 -3366
rect 35672 -3686 35992 -3366
rect 36391 -3686 36711 -3366
rect 37110 -3686 37430 -3366
rect 8672 -5390 8992 -5070
rect 9391 -5390 9711 -5070
rect 10110 -5390 10430 -5070
rect 10829 -5390 11149 -5070
rect 11548 -5390 11868 -5070
rect 23672 -5390 23992 -5070
rect 24391 -5390 24711 -5070
rect 25110 -5390 25430 -5070
rect 25829 -5390 26149 -5070
rect 26548 -5390 26868 -5070
rect 8672 -6090 8992 -5770
rect 9391 -6090 9711 -5770
rect 10110 -6090 10430 -5770
rect 10829 -6090 11149 -5770
rect 11548 -6090 11868 -5770
rect 23672 -6090 23992 -5770
rect 24391 -6090 24711 -5770
rect 25110 -6090 25430 -5770
rect 25829 -6090 26149 -5770
rect 26548 -6090 26868 -5770
rect 8672 -6790 8992 -6470
rect 9391 -6790 9711 -6470
rect 10110 -6790 10430 -6470
rect 10829 -6790 11149 -6470
rect 11548 -6790 11868 -6470
rect 23672 -6790 23992 -6470
rect 24391 -6790 24711 -6470
rect 25110 -6790 25430 -6470
rect 25829 -6790 26149 -6470
rect 26548 -6790 26868 -6470
rect 8672 -7490 8992 -7170
rect 9391 -7490 9711 -7170
rect 10110 -7490 10430 -7170
rect 10829 -7490 11149 -7170
rect 11548 -7490 11868 -7170
rect 23672 -7490 23992 -7170
rect 24391 -7490 24711 -7170
rect 25110 -7490 25430 -7170
rect 25829 -7490 26149 -7170
rect 26548 -7490 26868 -7170
rect 8672 -8190 8992 -7870
rect 9391 -8190 9711 -7870
rect 10110 -8190 10430 -7870
rect 10829 -8190 11149 -7870
rect 11548 -8190 11868 -7870
rect 23672 -8190 23992 -7870
rect 24391 -8190 24711 -7870
rect 25110 -8190 25430 -7870
rect 25829 -8190 26149 -7870
rect 26548 -8190 26868 -7870
rect 19234 -18886 19554 -18566
rect 19953 -18886 20273 -18566
rect 20672 -18886 20992 -18566
rect 21391 -18886 21711 -18566
rect 22110 -18886 22430 -18566
rect 34234 -18886 34554 -18566
rect 34953 -18886 35273 -18566
rect 35672 -18886 35992 -18566
rect 36391 -18886 36711 -18566
rect 37110 -18886 37430 -18566
rect 19234 -19586 19554 -19266
rect 19953 -19586 20273 -19266
rect 20672 -19586 20992 -19266
rect 21391 -19586 21711 -19266
rect 22110 -19586 22430 -19266
rect 34234 -19586 34554 -19266
rect 34953 -19586 35273 -19266
rect 35672 -19586 35992 -19266
rect 36391 -19586 36711 -19266
rect 37110 -19586 37430 -19266
rect 19234 -20286 19554 -19966
rect 19953 -20286 20273 -19966
rect 20672 -20286 20992 -19966
rect 21391 -20286 21711 -19966
rect 22110 -20286 22430 -19966
rect 34234 -20286 34554 -19966
rect 34953 -20286 35273 -19966
rect 35672 -20286 35992 -19966
rect 36391 -20286 36711 -19966
rect 37110 -20286 37430 -19966
rect 19234 -20986 19554 -20666
rect 19953 -20986 20273 -20666
rect 20672 -20986 20992 -20666
rect 21391 -20986 21711 -20666
rect 22110 -20986 22430 -20666
rect 34234 -20986 34554 -20666
rect 34953 -20986 35273 -20666
rect 35672 -20986 35992 -20666
rect 36391 -20986 36711 -20666
rect 37110 -20986 37430 -20666
rect 19234 -21686 19554 -21366
rect 19953 -21686 20273 -21366
rect 20672 -21686 20992 -21366
rect 21391 -21686 21711 -21366
rect 22110 -21686 22430 -21366
rect 34234 -21686 34554 -21366
rect 34953 -21686 35273 -21366
rect 35672 -21686 35992 -21366
rect 36391 -21686 36711 -21366
rect 37110 -21686 37430 -21366
<< metal4 >>
rect 23256 17542 38736 17578
rect 23256 17394 37972 17542
rect 23256 17094 23440 17394
rect 24040 17094 32072 17394
rect 32672 17094 37972 17394
rect 23256 16978 37972 17094
rect 23256 16868 23562 16978
rect 32558 16868 37972 16978
rect 23256 16812 37972 16868
rect 38702 16812 38736 17542
rect 23256 16778 38736 16812
rect 23256 11716 32856 11778
rect 23256 11572 24176 11716
rect 32038 11572 32856 11716
rect 23256 11462 32856 11572
rect 23256 11162 23440 11462
rect 24040 11162 32072 11462
rect 32672 11162 32856 11462
rect 23256 10812 32856 11162
rect 8118 10628 37822 10812
rect 8118 10328 13066 10628
rect 13448 10328 21200 10628
rect 21878 10328 23648 10628
rect 24248 10328 28280 10628
rect 28880 10328 37822 10628
rect 8118 10150 37822 10328
rect 8118 10064 15134 10150
rect 15230 10064 15714 10150
rect 15810 10064 16314 10150
rect 16410 10064 16914 10150
rect 17010 10064 17514 10150
rect 17610 10064 18114 10150
rect 18210 10064 18714 10150
rect 18810 10064 19314 10150
rect 19410 10064 19914 10150
rect 20010 10064 23896 10150
rect 23992 10064 24476 10150
rect 24572 10064 25076 10150
rect 25172 10064 25676 10150
rect 25772 10064 26276 10150
rect 26372 10064 26876 10150
rect 26972 10064 27476 10150
rect 27572 10064 28076 10150
rect 28172 10064 28676 10150
rect 28772 10064 37822 10150
rect 8118 10012 37822 10064
rect 30394 8452 30514 10012
rect 30394 8380 30406 8452
rect 30502 8380 30514 8452
rect 30394 7364 30514 8380
rect 30394 7292 30406 7364
rect 30502 7292 30514 7364
rect 30394 6276 30514 7292
rect 30394 6204 30406 6276
rect 30502 6204 30514 6276
rect 30394 5648 30514 6204
rect 33074 8996 33194 9008
rect 33074 8924 33086 8996
rect 33182 8924 33194 8996
rect 33074 7908 33194 8924
rect 33074 7836 33086 7908
rect 33182 7836 33194 7908
rect 33074 6820 33194 7836
rect 33074 6748 33086 6820
rect 33182 6748 33194 6820
rect 33074 5732 33194 6748
rect 33074 5660 33086 5732
rect 33182 5660 33194 5732
rect 12882 5484 29064 5488
rect 33074 5484 33194 5660
rect 35772 8452 35892 10012
rect 35772 8380 35784 8452
rect 35880 8380 35892 8452
rect 35772 7364 35892 8380
rect 35772 7292 35784 7364
rect 35880 7292 35892 7364
rect 35772 6276 35892 7292
rect 35772 6204 35784 6276
rect 35880 6204 35892 6276
rect 35772 5648 35892 6204
rect 8278 5450 38743 5484
rect 8278 5172 37966 5450
rect 8278 4872 13066 5172
rect 13448 4872 21200 5172
rect 21878 4872 23648 5172
rect 24248 4872 28280 5172
rect 28880 4872 37966 5172
rect 8278 4474 37966 4872
rect 8274 4290 37966 4474
rect 8274 3990 8458 4290
rect 9058 3990 18090 4290
rect 18690 3990 23458 4290
rect 24058 3990 33090 4290
rect 33690 3990 37966 4290
rect 8274 3816 37966 3990
rect 8274 3730 9310 3816
rect 9406 3730 9910 3816
rect 10006 3730 10510 3816
rect 10606 3730 11110 3816
rect 11206 3730 11710 3816
rect 11806 3730 12310 3816
rect 12406 3730 12910 3816
rect 13006 3730 13510 3816
rect 13606 3730 14110 3816
rect 14206 3730 14710 3816
rect 14806 3730 15310 3816
rect 15406 3730 15910 3816
rect 16006 3730 16510 3816
rect 16606 3730 17110 3816
rect 17206 3730 17530 3816
rect 17626 3730 24310 3816
rect 24406 3730 24910 3816
rect 25006 3730 25510 3816
rect 25606 3730 26110 3816
rect 26206 3730 26710 3816
rect 26806 3730 27310 3816
rect 27406 3730 27910 3816
rect 28006 3730 28510 3816
rect 28606 3730 29110 3816
rect 29206 3730 29710 3816
rect 29806 3730 30310 3816
rect 30406 3730 30910 3816
rect 31006 3730 31510 3816
rect 31606 3730 32110 3816
rect 32206 3730 32530 3816
rect 32626 3730 37966 3816
rect 8274 3702 37966 3730
rect 38712 3702 38743 5450
rect 8274 3674 38743 3702
rect 19693 -542 19789 -526
rect 19233 -566 19555 -565
rect 19233 -886 19234 -566
rect 19554 -682 19555 -566
rect 19693 -682 19709 -542
rect 19554 -782 19709 -682
rect 19554 -886 19555 -782
rect 19233 -887 19555 -886
rect 19348 -1265 19448 -887
rect 19684 -914 19709 -782
rect 19773 -682 19789 -542
rect 20412 -544 20508 -528
rect 19952 -566 20274 -565
rect 19952 -682 19953 -566
rect 19773 -782 19953 -682
rect 19773 -914 19789 -782
rect 19952 -886 19953 -782
rect 20273 -682 20274 -566
rect 20412 -682 20428 -544
rect 20273 -782 20428 -682
rect 20273 -886 20274 -782
rect 19952 -887 20274 -886
rect 19684 -930 19789 -914
rect 20412 -914 20428 -782
rect 20492 -682 20508 -544
rect 21131 -544 21227 -528
rect 20671 -566 20993 -565
rect 20671 -682 20672 -566
rect 20492 -782 20672 -682
rect 20492 -914 20508 -782
rect 20671 -886 20672 -782
rect 20992 -682 20993 -566
rect 21131 -682 21147 -544
rect 20992 -782 21147 -682
rect 20992 -886 20993 -782
rect 20671 -887 20993 -886
rect 20412 -930 20508 -914
rect 21131 -914 21147 -782
rect 21211 -682 21227 -544
rect 21850 -544 21946 -528
rect 21390 -566 21712 -565
rect 21390 -682 21391 -566
rect 21211 -782 21391 -682
rect 21211 -914 21227 -782
rect 21390 -886 21391 -782
rect 21711 -682 21712 -566
rect 21850 -682 21866 -544
rect 21711 -782 21866 -682
rect 21711 -886 21712 -782
rect 21390 -887 21712 -886
rect 21131 -930 21227 -914
rect 21850 -914 21866 -782
rect 21930 -682 21946 -544
rect 22569 -544 22665 -528
rect 22109 -566 22431 -565
rect 22109 -682 22110 -566
rect 21930 -782 22110 -682
rect 21930 -914 21952 -782
rect 22109 -886 22110 -782
rect 22430 -682 22431 -566
rect 22569 -682 22585 -544
rect 22430 -782 22585 -682
rect 22430 -886 22431 -782
rect 22109 -887 22431 -886
rect 19684 -1228 19784 -930
rect 20062 -1136 21606 -1036
rect 19684 -1244 19789 -1228
rect 19233 -1266 19555 -1265
rect 19233 -1586 19234 -1266
rect 19554 -1372 19555 -1266
rect 19684 -1372 19709 -1244
rect 19554 -1472 19709 -1372
rect 19554 -1586 19555 -1472
rect 19684 -1586 19709 -1472
rect 19233 -1587 19555 -1586
rect 19693 -1612 19709 -1586
rect 19773 -1612 19789 -1244
rect 20062 -1265 20162 -1136
rect 20412 -1244 20508 -1228
rect 19952 -1266 20274 -1265
rect 19952 -1586 19953 -1266
rect 20273 -1586 20274 -1266
rect 19952 -1587 20274 -1586
rect 19693 -1632 19789 -1612
rect 20062 -1728 20162 -1587
rect 20412 -1612 20428 -1244
rect 20492 -1612 20508 -1244
rect 20782 -1265 20882 -1136
rect 21131 -1244 21227 -1228
rect 20671 -1266 20993 -1265
rect 20671 -1586 20672 -1266
rect 20992 -1586 20993 -1266
rect 20671 -1587 20993 -1586
rect 20412 -1632 20508 -1612
rect 20782 -1728 20882 -1587
rect 21131 -1612 21147 -1244
rect 21211 -1612 21227 -1244
rect 21504 -1265 21605 -1136
rect 21850 -1244 21952 -914
rect 21390 -1266 21712 -1265
rect 21390 -1586 21391 -1266
rect 21711 -1586 21712 -1266
rect 21390 -1587 21712 -1586
rect 21131 -1632 21227 -1612
rect 21504 -1728 21605 -1587
rect 21850 -1612 21866 -1244
rect 21930 -1376 21952 -1244
rect 22224 -1265 22324 -887
rect 22562 -914 22585 -782
rect 22649 -914 22665 -544
rect 34693 -542 34789 -526
rect 34233 -566 34555 -565
rect 34233 -886 34234 -566
rect 34554 -682 34555 -566
rect 34693 -682 34709 -542
rect 34554 -782 34709 -682
rect 34554 -886 34555 -782
rect 34233 -887 34555 -886
rect 22562 -1244 22665 -914
rect 22109 -1266 22431 -1265
rect 22109 -1376 22110 -1266
rect 21930 -1476 22110 -1376
rect 21930 -1612 21952 -1476
rect 22109 -1586 22110 -1476
rect 22430 -1376 22431 -1266
rect 22562 -1376 22585 -1244
rect 22430 -1476 22585 -1376
rect 22430 -1586 22431 -1476
rect 22109 -1587 22431 -1586
rect 22224 -1588 22324 -1587
rect 21850 -1626 21952 -1612
rect 22562 -1612 22585 -1476
rect 22649 -1612 22665 -1244
rect 34348 -1265 34448 -887
rect 34684 -914 34709 -782
rect 34773 -682 34789 -542
rect 35412 -544 35508 -528
rect 34952 -566 35274 -565
rect 34952 -682 34953 -566
rect 34773 -782 34953 -682
rect 34773 -914 34789 -782
rect 34952 -886 34953 -782
rect 35273 -682 35274 -566
rect 35412 -682 35428 -544
rect 35273 -782 35428 -682
rect 35273 -886 35274 -782
rect 34952 -887 35274 -886
rect 34684 -930 34789 -914
rect 35412 -914 35428 -782
rect 35492 -682 35508 -544
rect 36131 -544 36227 -528
rect 35671 -566 35993 -565
rect 35671 -682 35672 -566
rect 35492 -782 35672 -682
rect 35492 -914 35508 -782
rect 35671 -886 35672 -782
rect 35992 -682 35993 -566
rect 36131 -682 36147 -544
rect 35992 -782 36147 -682
rect 35992 -886 35993 -782
rect 35671 -887 35993 -886
rect 35412 -930 35508 -914
rect 36131 -914 36147 -782
rect 36211 -682 36227 -544
rect 36850 -544 36946 -528
rect 36390 -566 36712 -565
rect 36390 -682 36391 -566
rect 36211 -782 36391 -682
rect 36211 -914 36227 -782
rect 36390 -886 36391 -782
rect 36711 -682 36712 -566
rect 36850 -682 36866 -544
rect 36711 -782 36866 -682
rect 36711 -886 36712 -782
rect 36390 -887 36712 -886
rect 36131 -930 36227 -914
rect 36850 -914 36866 -782
rect 36930 -682 36946 -544
rect 37569 -544 37665 -528
rect 37109 -566 37431 -565
rect 37109 -682 37110 -566
rect 36930 -782 37110 -682
rect 36930 -914 36952 -782
rect 37109 -886 37110 -782
rect 37430 -682 37431 -566
rect 37569 -682 37585 -544
rect 37430 -782 37585 -682
rect 37430 -886 37431 -782
rect 37109 -887 37431 -886
rect 34684 -1228 34784 -930
rect 35062 -1136 36606 -1036
rect 34684 -1244 34789 -1228
rect 34233 -1266 34555 -1265
rect 34233 -1586 34234 -1266
rect 34554 -1372 34555 -1266
rect 34684 -1372 34709 -1244
rect 34554 -1472 34709 -1372
rect 34554 -1586 34555 -1472
rect 34684 -1586 34709 -1472
rect 34233 -1587 34555 -1586
rect 22562 -1626 22665 -1612
rect 21850 -1632 21946 -1626
rect 22569 -1632 22665 -1626
rect 34693 -1612 34709 -1586
rect 34773 -1612 34789 -1244
rect 35062 -1265 35162 -1136
rect 35412 -1244 35508 -1228
rect 34952 -1266 35274 -1265
rect 34952 -1586 34953 -1266
rect 35273 -1586 35274 -1266
rect 34952 -1587 35274 -1586
rect 34693 -1632 34789 -1612
rect 35062 -1728 35162 -1587
rect 35412 -1612 35428 -1244
rect 35492 -1612 35508 -1244
rect 35782 -1265 35882 -1136
rect 36131 -1244 36227 -1228
rect 35671 -1266 35993 -1265
rect 35671 -1586 35672 -1266
rect 35992 -1586 35993 -1266
rect 35671 -1587 35993 -1586
rect 35412 -1632 35508 -1612
rect 35782 -1728 35882 -1587
rect 36131 -1612 36147 -1244
rect 36211 -1612 36227 -1244
rect 36504 -1265 36605 -1136
rect 36850 -1244 36952 -914
rect 36390 -1266 36712 -1265
rect 36390 -1586 36391 -1266
rect 36711 -1586 36712 -1266
rect 36390 -1587 36712 -1586
rect 36131 -1632 36227 -1612
rect 36504 -1728 36605 -1587
rect 36850 -1612 36866 -1244
rect 36930 -1376 36952 -1244
rect 37224 -1265 37324 -887
rect 37562 -914 37585 -782
rect 37649 -914 37665 -544
rect 37562 -1244 37665 -914
rect 37109 -1266 37431 -1265
rect 37109 -1376 37110 -1266
rect 36930 -1476 37110 -1376
rect 36930 -1612 36952 -1476
rect 37109 -1586 37110 -1476
rect 37430 -1376 37431 -1266
rect 37562 -1376 37585 -1244
rect 37430 -1476 37585 -1376
rect 37430 -1586 37431 -1476
rect 37109 -1587 37431 -1586
rect 37224 -1588 37324 -1587
rect 36850 -1626 36952 -1612
rect 37562 -1612 37585 -1476
rect 37649 -1612 37665 -1244
rect 37562 -1626 37665 -1612
rect 36850 -1632 36946 -1626
rect 37569 -1632 37665 -1626
rect 18872 -1729 22906 -1728
rect 18872 -1827 18873 -1729
rect 18971 -1827 22807 -1729
rect 22905 -1827 22906 -1729
rect 18872 -1828 22906 -1827
rect 33872 -1729 37824 -1728
rect 33872 -1827 33873 -1729
rect 33971 -1827 37824 -1729
rect 33872 -1828 37824 -1827
rect 19693 -1944 19789 -1928
rect 19693 -1964 19709 -1944
rect 19348 -1965 19448 -1964
rect 19233 -1966 19555 -1965
rect 19233 -2286 19234 -1966
rect 19554 -2074 19555 -1966
rect 19684 -2074 19709 -1964
rect 19554 -2174 19709 -2074
rect 19554 -2286 19555 -2174
rect 19233 -2287 19555 -2286
rect 19348 -2665 19448 -2287
rect 19684 -2312 19709 -2174
rect 19773 -2312 19789 -1944
rect 20062 -1965 20162 -1828
rect 20412 -1944 20508 -1928
rect 19952 -1966 20274 -1965
rect 19952 -2286 19953 -1966
rect 20273 -2286 20274 -1966
rect 19952 -2287 20274 -2286
rect 19684 -2330 19789 -2312
rect 19684 -2628 19784 -2330
rect 20062 -2430 20162 -2287
rect 20412 -2312 20428 -1944
rect 20492 -2312 20508 -1944
rect 20782 -1965 20882 -1828
rect 21131 -1944 21227 -1928
rect 20671 -1966 20993 -1965
rect 20671 -2286 20672 -1966
rect 20992 -2286 20993 -1966
rect 20671 -2287 20993 -2286
rect 20412 -2330 20508 -2312
rect 20782 -2430 20882 -2287
rect 21131 -2312 21147 -1944
rect 21211 -2312 21227 -1944
rect 21504 -1965 21605 -1828
rect 21852 -1928 21952 -1926
rect 21850 -1944 21952 -1928
rect 21390 -1966 21712 -1965
rect 21390 -2286 21391 -1966
rect 21711 -2286 21712 -1966
rect 21390 -2287 21712 -2286
rect 21131 -2330 21227 -2312
rect 21504 -2430 21605 -2287
rect 21850 -2312 21866 -1944
rect 21930 -2080 21952 -1944
rect 22562 -1928 22662 -1926
rect 22562 -1944 22665 -1928
rect 22224 -1965 22324 -1964
rect 22109 -1966 22431 -1965
rect 22109 -2080 22110 -1966
rect 21930 -2180 22110 -2080
rect 21930 -2312 21952 -2180
rect 22109 -2286 22110 -2180
rect 22430 -2080 22431 -1966
rect 22562 -2080 22585 -1944
rect 22430 -2180 22585 -2080
rect 22430 -2286 22431 -2180
rect 22109 -2287 22431 -2286
rect 21850 -2330 21952 -2312
rect 20062 -2530 21605 -2430
rect 19684 -2644 19789 -2628
rect 19233 -2666 19555 -2665
rect 19233 -2986 19234 -2666
rect 19554 -2780 19555 -2666
rect 19684 -2780 19709 -2644
rect 19554 -2880 19709 -2780
rect 19554 -2986 19555 -2880
rect 19233 -2987 19555 -2986
rect 19348 -3365 19448 -2987
rect 19684 -3012 19709 -2880
rect 19773 -3012 19789 -2644
rect 20062 -2665 20162 -2530
rect 20412 -2644 20508 -2628
rect 19952 -2666 20274 -2665
rect 19952 -2986 19953 -2666
rect 20273 -2986 20274 -2666
rect 19952 -2987 20274 -2986
rect 19684 -3030 19789 -3012
rect 19684 -3328 19784 -3030
rect 20062 -3130 20162 -2987
rect 20412 -3012 20428 -2644
rect 20492 -3012 20508 -2644
rect 20782 -2665 20882 -2530
rect 21131 -2644 21227 -2628
rect 20671 -2666 20993 -2665
rect 20671 -2986 20672 -2666
rect 20992 -2986 20993 -2666
rect 20671 -2987 20993 -2986
rect 20412 -3030 20508 -3012
rect 20782 -3130 20882 -2987
rect 21131 -3012 21147 -2644
rect 21211 -3012 21227 -2644
rect 21504 -2665 21605 -2530
rect 21852 -2628 21952 -2330
rect 21850 -2644 21952 -2628
rect 21390 -2666 21712 -2665
rect 21390 -2986 21391 -2666
rect 21711 -2986 21712 -2666
rect 21390 -2987 21712 -2986
rect 21131 -3030 21227 -3012
rect 21504 -3130 21605 -2987
rect 21850 -3012 21866 -2644
rect 21930 -2772 21952 -2644
rect 22224 -2665 22324 -2287
rect 22562 -2312 22585 -2180
rect 22649 -2312 22665 -1944
rect 34693 -1944 34789 -1928
rect 34693 -1964 34709 -1944
rect 34348 -1965 34448 -1964
rect 34233 -1966 34555 -1965
rect 34233 -2286 34234 -1966
rect 34554 -2074 34555 -1966
rect 34684 -2074 34709 -1964
rect 34554 -2174 34709 -2074
rect 34554 -2286 34555 -2174
rect 34233 -2287 34555 -2286
rect 22562 -2330 22665 -2312
rect 22562 -2628 22662 -2330
rect 22562 -2644 22665 -2628
rect 22109 -2666 22431 -2665
rect 22109 -2772 22110 -2666
rect 21930 -2872 22110 -2772
rect 21930 -3012 21952 -2872
rect 22109 -2986 22110 -2872
rect 22430 -2772 22431 -2666
rect 22562 -2772 22585 -2644
rect 22430 -2872 22585 -2772
rect 22430 -2986 22431 -2872
rect 22109 -2987 22431 -2986
rect 20062 -3230 21606 -3130
rect 19684 -3344 19789 -3328
rect 19233 -3366 19555 -3365
rect 19233 -3426 19234 -3366
rect 7314 -3454 19234 -3426
rect 7314 -5298 7348 -3454
rect 8082 -3478 19234 -3454
rect 8082 -3564 8744 -3478
rect 8840 -3564 9324 -3478
rect 9420 -3564 9924 -3478
rect 10020 -3564 10524 -3478
rect 10620 -3564 11124 -3478
rect 11220 -3564 11724 -3478
rect 11820 -3564 12324 -3478
rect 12420 -3564 12924 -3478
rect 13020 -3564 13524 -3478
rect 13620 -3564 14124 -3478
rect 14220 -3564 14724 -3478
rect 14820 -3564 15324 -3478
rect 15420 -3564 15924 -3478
rect 16020 -3564 16524 -3478
rect 16620 -3564 17124 -3478
rect 17220 -3564 17724 -3478
rect 17820 -3564 18324 -3478
rect 18420 -3564 19234 -3478
rect 8082 -3686 19234 -3564
rect 19554 -3426 19555 -3366
rect 19684 -3426 19709 -3344
rect 19554 -3686 19709 -3426
rect 8082 -3712 19709 -3686
rect 19773 -3426 19789 -3344
rect 20412 -3344 20508 -3328
rect 19952 -3366 20274 -3365
rect 19952 -3426 19953 -3366
rect 19773 -3686 19953 -3426
rect 20273 -3426 20274 -3366
rect 20412 -3426 20428 -3344
rect 20273 -3686 20428 -3426
rect 19773 -3712 20428 -3686
rect 20492 -3426 20508 -3344
rect 21131 -3344 21227 -3328
rect 20671 -3366 20993 -3365
rect 20671 -3426 20672 -3366
rect 20492 -3686 20672 -3426
rect 20992 -3426 20993 -3366
rect 21131 -3426 21147 -3344
rect 20992 -3686 21147 -3426
rect 20492 -3712 21147 -3686
rect 21211 -3426 21227 -3344
rect 21850 -3344 21952 -3012
rect 21390 -3366 21712 -3365
rect 21390 -3426 21391 -3366
rect 21211 -3686 21391 -3426
rect 21711 -3426 21712 -3366
rect 21850 -3426 21866 -3344
rect 21711 -3686 21866 -3426
rect 21211 -3712 21866 -3686
rect 21930 -3426 21952 -3344
rect 22224 -3365 22324 -2987
rect 22562 -3012 22585 -2872
rect 22649 -3012 22665 -2644
rect 34348 -2665 34448 -2287
rect 34684 -2312 34709 -2174
rect 34773 -2312 34789 -1944
rect 35062 -1965 35162 -1828
rect 35412 -1944 35508 -1928
rect 34952 -1966 35274 -1965
rect 34952 -2286 34953 -1966
rect 35273 -2286 35274 -1966
rect 34952 -2287 35274 -2286
rect 34684 -2330 34789 -2312
rect 34684 -2628 34784 -2330
rect 35062 -2430 35162 -2287
rect 35412 -2312 35428 -1944
rect 35492 -2312 35508 -1944
rect 35782 -1965 35882 -1828
rect 36131 -1944 36227 -1928
rect 35671 -1966 35993 -1965
rect 35671 -2286 35672 -1966
rect 35992 -2286 35993 -1966
rect 35671 -2287 35993 -2286
rect 35412 -2330 35508 -2312
rect 35782 -2430 35882 -2287
rect 36131 -2312 36147 -1944
rect 36211 -2312 36227 -1944
rect 36504 -1965 36605 -1828
rect 36852 -1928 36952 -1926
rect 36850 -1944 36952 -1928
rect 36390 -1966 36712 -1965
rect 36390 -2286 36391 -1966
rect 36711 -2286 36712 -1966
rect 36390 -2287 36712 -2286
rect 36131 -2330 36227 -2312
rect 36504 -2430 36605 -2287
rect 36850 -2312 36866 -1944
rect 36930 -2080 36952 -1944
rect 37562 -1928 37662 -1926
rect 37562 -1944 37665 -1928
rect 37224 -1965 37324 -1964
rect 37109 -1966 37431 -1965
rect 37109 -2080 37110 -1966
rect 36930 -2180 37110 -2080
rect 36930 -2312 36952 -2180
rect 37109 -2286 37110 -2180
rect 37430 -2080 37431 -1966
rect 37562 -2080 37585 -1944
rect 37430 -2180 37585 -2080
rect 37430 -2286 37431 -2180
rect 37109 -2287 37431 -2286
rect 36850 -2330 36952 -2312
rect 35062 -2530 36605 -2430
rect 34684 -2644 34789 -2628
rect 34233 -2666 34555 -2665
rect 34233 -2986 34234 -2666
rect 34554 -2780 34555 -2666
rect 34684 -2780 34709 -2644
rect 34554 -2880 34709 -2780
rect 34554 -2986 34555 -2880
rect 34233 -2987 34555 -2986
rect 22562 -3344 22665 -3012
rect 22109 -3366 22431 -3365
rect 22109 -3426 22110 -3366
rect 21930 -3686 22110 -3426
rect 22430 -3426 22431 -3366
rect 22562 -3426 22585 -3344
rect 22430 -3686 22585 -3426
rect 21930 -3712 22585 -3686
rect 22649 -3426 22665 -3344
rect 34348 -3365 34448 -2987
rect 34684 -3012 34709 -2880
rect 34773 -3012 34789 -2644
rect 35062 -2665 35162 -2530
rect 35412 -2644 35508 -2628
rect 34952 -2666 35274 -2665
rect 34952 -2986 34953 -2666
rect 35273 -2986 35274 -2666
rect 34952 -2987 35274 -2986
rect 34684 -3030 34789 -3012
rect 34684 -3328 34784 -3030
rect 35062 -3130 35162 -2987
rect 35412 -3012 35428 -2644
rect 35492 -3012 35508 -2644
rect 35782 -2665 35882 -2530
rect 36131 -2644 36227 -2628
rect 35671 -2666 35993 -2665
rect 35671 -2986 35672 -2666
rect 35992 -2986 35993 -2666
rect 35671 -2987 35993 -2986
rect 35412 -3030 35508 -3012
rect 35782 -3130 35882 -2987
rect 36131 -3012 36147 -2644
rect 36211 -3012 36227 -2644
rect 36504 -2665 36605 -2530
rect 36852 -2628 36952 -2330
rect 36850 -2644 36952 -2628
rect 36390 -2666 36712 -2665
rect 36390 -2986 36391 -2666
rect 36711 -2986 36712 -2666
rect 36390 -2987 36712 -2986
rect 36131 -3030 36227 -3012
rect 36504 -3130 36605 -2987
rect 36850 -3012 36866 -2644
rect 36930 -2772 36952 -2644
rect 37224 -2665 37324 -2287
rect 37562 -2312 37585 -2180
rect 37649 -2312 37665 -1944
rect 37562 -2330 37665 -2312
rect 37562 -2628 37662 -2330
rect 37562 -2644 37665 -2628
rect 37109 -2666 37431 -2665
rect 37109 -2772 37110 -2666
rect 36930 -2872 37110 -2772
rect 36930 -3012 36952 -2872
rect 37109 -2986 37110 -2872
rect 37430 -2772 37431 -2666
rect 37562 -2772 37585 -2644
rect 37430 -2872 37585 -2772
rect 37430 -2986 37431 -2872
rect 37109 -2987 37431 -2986
rect 35062 -3230 36606 -3130
rect 34684 -3344 34789 -3328
rect 34233 -3366 34555 -3365
rect 34233 -3426 34234 -3366
rect 22649 -3478 34234 -3426
rect 22649 -3564 23744 -3478
rect 23840 -3564 24324 -3478
rect 24420 -3564 24924 -3478
rect 25020 -3564 25524 -3478
rect 25620 -3564 26124 -3478
rect 26220 -3564 26724 -3478
rect 26820 -3564 27324 -3478
rect 27420 -3564 27924 -3478
rect 28020 -3564 28524 -3478
rect 28620 -3564 29124 -3478
rect 29220 -3564 29724 -3478
rect 29820 -3564 30324 -3478
rect 30420 -3564 30924 -3478
rect 31020 -3564 31524 -3478
rect 31620 -3564 32124 -3478
rect 32220 -3564 32724 -3478
rect 32820 -3564 33324 -3478
rect 33420 -3564 34234 -3478
rect 22649 -3686 34234 -3564
rect 34554 -3426 34555 -3366
rect 34684 -3426 34709 -3344
rect 34554 -3686 34709 -3426
rect 22649 -3712 34709 -3686
rect 34773 -3426 34789 -3344
rect 35412 -3344 35508 -3328
rect 34952 -3366 35274 -3365
rect 34952 -3426 34953 -3366
rect 34773 -3686 34953 -3426
rect 35273 -3426 35274 -3366
rect 35412 -3426 35428 -3344
rect 35273 -3686 35428 -3426
rect 34773 -3712 35428 -3686
rect 35492 -3426 35508 -3344
rect 36131 -3344 36227 -3328
rect 35671 -3366 35993 -3365
rect 35671 -3426 35672 -3366
rect 35492 -3686 35672 -3426
rect 35992 -3426 35993 -3366
rect 36131 -3426 36147 -3344
rect 35992 -3686 36147 -3426
rect 35492 -3712 36147 -3686
rect 36211 -3426 36227 -3344
rect 36850 -3344 36952 -3012
rect 36390 -3366 36712 -3365
rect 36390 -3426 36391 -3366
rect 36211 -3686 36391 -3426
rect 36711 -3426 36712 -3366
rect 36850 -3426 36866 -3344
rect 36711 -3686 36866 -3426
rect 36211 -3712 36866 -3686
rect 36930 -3426 36952 -3344
rect 37224 -3365 37324 -2987
rect 37562 -3012 37585 -2872
rect 37649 -3012 37665 -2644
rect 37562 -3344 37665 -3012
rect 37109 -3366 37431 -3365
rect 37109 -3426 37110 -3366
rect 36930 -3686 37110 -3426
rect 37430 -3426 37431 -3366
rect 37562 -3426 37585 -3344
rect 37430 -3686 37585 -3426
rect 36930 -3712 37585 -3686
rect 37649 -3426 37665 -3344
rect 37649 -3432 37822 -3426
rect 37649 -3712 37826 -3432
rect 8082 -3742 37826 -3712
rect 8082 -4042 8458 -3742
rect 9058 -4042 18090 -3742
rect 18690 -4042 23458 -3742
rect 24058 -4042 33090 -3742
rect 33690 -4042 37826 -3742
rect 8082 -4530 37826 -4042
rect 8082 -4714 37828 -4530
rect 8082 -5014 12412 -4714
rect 13012 -5014 22044 -4714
rect 22644 -5014 27412 -4714
rect 28012 -5014 37044 -4714
rect 37644 -5014 37828 -4714
rect 8082 -5044 37828 -5014
rect 8082 -5298 8453 -5044
rect 7314 -5330 8453 -5298
rect 8437 -5412 8453 -5330
rect 8517 -5070 9172 -5044
rect 8517 -5330 8672 -5070
rect 8517 -5412 8540 -5330
rect 8671 -5390 8672 -5330
rect 8992 -5330 9172 -5070
rect 8992 -5390 8993 -5330
rect 8671 -5391 8993 -5390
rect 8437 -5744 8540 -5412
rect 8437 -6112 8453 -5744
rect 8517 -5884 8540 -5744
rect 8778 -5769 8878 -5391
rect 9150 -5412 9172 -5330
rect 9236 -5070 9891 -5044
rect 9236 -5330 9391 -5070
rect 9236 -5412 9252 -5330
rect 9390 -5390 9391 -5330
rect 9711 -5330 9891 -5070
rect 9711 -5390 9712 -5330
rect 9390 -5391 9712 -5390
rect 9150 -5744 9252 -5412
rect 9875 -5412 9891 -5330
rect 9955 -5070 10610 -5044
rect 9955 -5330 10110 -5070
rect 9955 -5412 9971 -5330
rect 10109 -5390 10110 -5330
rect 10430 -5330 10610 -5070
rect 10430 -5390 10431 -5330
rect 10109 -5391 10431 -5390
rect 9875 -5428 9971 -5412
rect 10594 -5412 10610 -5330
rect 10674 -5070 11329 -5044
rect 10674 -5330 10829 -5070
rect 10674 -5412 10690 -5330
rect 10828 -5390 10829 -5330
rect 11149 -5330 11329 -5070
rect 11149 -5390 11150 -5330
rect 10828 -5391 11150 -5390
rect 10594 -5428 10690 -5412
rect 11313 -5412 11329 -5330
rect 11393 -5070 23453 -5044
rect 11393 -5330 11548 -5070
rect 11393 -5412 11418 -5330
rect 11547 -5390 11548 -5330
rect 11868 -5192 23453 -5070
rect 11868 -5278 12682 -5192
rect 12778 -5278 13282 -5192
rect 13378 -5278 13882 -5192
rect 13978 -5278 14482 -5192
rect 14578 -5278 15082 -5192
rect 15178 -5278 15682 -5192
rect 15778 -5278 16282 -5192
rect 16378 -5278 16882 -5192
rect 16978 -5278 17482 -5192
rect 17578 -5278 18082 -5192
rect 18178 -5278 18682 -5192
rect 18778 -5278 19282 -5192
rect 19378 -5278 19882 -5192
rect 19978 -5278 20482 -5192
rect 20578 -5278 21082 -5192
rect 21178 -5278 21682 -5192
rect 21778 -5278 22262 -5192
rect 22358 -5278 23453 -5192
rect 11868 -5330 23453 -5278
rect 11868 -5390 11869 -5330
rect 11547 -5391 11869 -5390
rect 11313 -5428 11418 -5412
rect 9496 -5626 11040 -5526
rect 8671 -5770 8993 -5769
rect 8671 -5884 8672 -5770
rect 8517 -5984 8672 -5884
rect 8517 -6112 8540 -5984
rect 8671 -6090 8672 -5984
rect 8992 -5884 8993 -5770
rect 9150 -5884 9172 -5744
rect 8992 -5984 9172 -5884
rect 8992 -6090 8993 -5984
rect 8671 -6091 8993 -6090
rect 8437 -6128 8540 -6112
rect 8440 -6426 8540 -6128
rect 8437 -6444 8540 -6426
rect 8437 -6812 8453 -6444
rect 8517 -6576 8540 -6444
rect 8778 -6469 8878 -6091
rect 9150 -6112 9172 -5984
rect 9236 -6112 9252 -5744
rect 9497 -5769 9598 -5626
rect 9875 -5744 9971 -5726
rect 9390 -5770 9712 -5769
rect 9390 -6090 9391 -5770
rect 9711 -6090 9712 -5770
rect 9390 -6091 9712 -6090
rect 9150 -6128 9252 -6112
rect 9150 -6426 9250 -6128
rect 9497 -6226 9598 -6091
rect 9875 -6112 9891 -5744
rect 9955 -6112 9971 -5744
rect 10220 -5769 10320 -5626
rect 10594 -5744 10690 -5726
rect 10109 -5770 10431 -5769
rect 10109 -6090 10110 -5770
rect 10430 -6090 10431 -5770
rect 10109 -6091 10431 -6090
rect 9875 -6128 9971 -6112
rect 10220 -6226 10320 -6091
rect 10594 -6112 10610 -5744
rect 10674 -6112 10690 -5744
rect 10940 -5769 11040 -5626
rect 11318 -5726 11418 -5428
rect 11313 -5744 11418 -5726
rect 10828 -5770 11150 -5769
rect 10828 -6090 10829 -5770
rect 11149 -6090 11150 -5770
rect 10828 -6091 11150 -6090
rect 10594 -6128 10690 -6112
rect 10940 -6226 11040 -6091
rect 11313 -6112 11329 -5744
rect 11393 -5876 11418 -5744
rect 11654 -5769 11754 -5391
rect 23437 -5412 23453 -5330
rect 23517 -5070 24172 -5044
rect 23517 -5330 23672 -5070
rect 23517 -5412 23540 -5330
rect 23671 -5390 23672 -5330
rect 23992 -5330 24172 -5070
rect 23992 -5390 23993 -5330
rect 23671 -5391 23993 -5390
rect 23437 -5744 23540 -5412
rect 11547 -5770 11869 -5769
rect 11547 -5876 11548 -5770
rect 11393 -5976 11548 -5876
rect 11393 -6112 11418 -5976
rect 11547 -6090 11548 -5976
rect 11868 -6090 11869 -5770
rect 11547 -6091 11869 -6090
rect 11313 -6128 11418 -6112
rect 9497 -6326 11040 -6226
rect 9150 -6444 9252 -6426
rect 8671 -6470 8993 -6469
rect 8671 -6576 8672 -6470
rect 8517 -6676 8672 -6576
rect 8517 -6812 8540 -6676
rect 8671 -6790 8672 -6676
rect 8992 -6576 8993 -6470
rect 9150 -6576 9172 -6444
rect 8992 -6676 9172 -6576
rect 8992 -6790 8993 -6676
rect 8671 -6791 8993 -6790
rect 8778 -6792 8878 -6791
rect 8437 -6828 8540 -6812
rect 8440 -6830 8540 -6828
rect 9150 -6812 9172 -6676
rect 9236 -6812 9252 -6444
rect 9497 -6469 9598 -6326
rect 9875 -6444 9971 -6426
rect 9390 -6470 9712 -6469
rect 9390 -6790 9391 -6470
rect 9711 -6790 9712 -6470
rect 9390 -6791 9712 -6790
rect 9150 -6828 9252 -6812
rect 9150 -6830 9250 -6828
rect 9497 -6928 9598 -6791
rect 9875 -6812 9891 -6444
rect 9955 -6812 9971 -6444
rect 10220 -6469 10320 -6326
rect 10594 -6444 10690 -6426
rect 10109 -6470 10431 -6469
rect 10109 -6790 10110 -6470
rect 10430 -6790 10431 -6470
rect 10109 -6791 10431 -6790
rect 9875 -6828 9971 -6812
rect 10220 -6928 10320 -6791
rect 10594 -6812 10610 -6444
rect 10674 -6812 10690 -6444
rect 10940 -6469 11040 -6326
rect 11318 -6426 11418 -6128
rect 11313 -6444 11418 -6426
rect 10828 -6470 11150 -6469
rect 10828 -6790 10829 -6470
rect 11149 -6790 11150 -6470
rect 10828 -6791 11150 -6790
rect 10594 -6828 10690 -6812
rect 10940 -6928 11040 -6791
rect 11313 -6812 11329 -6444
rect 11393 -6582 11418 -6444
rect 11654 -6469 11754 -6091
rect 23437 -6112 23453 -5744
rect 23517 -5884 23540 -5744
rect 23778 -5769 23878 -5391
rect 24150 -5412 24172 -5330
rect 24236 -5070 24891 -5044
rect 24236 -5330 24391 -5070
rect 24236 -5412 24252 -5330
rect 24390 -5390 24391 -5330
rect 24711 -5330 24891 -5070
rect 24711 -5390 24712 -5330
rect 24390 -5391 24712 -5390
rect 24150 -5744 24252 -5412
rect 24875 -5412 24891 -5330
rect 24955 -5070 25610 -5044
rect 24955 -5330 25110 -5070
rect 24955 -5412 24971 -5330
rect 25109 -5390 25110 -5330
rect 25430 -5330 25610 -5070
rect 25430 -5390 25431 -5330
rect 25109 -5391 25431 -5390
rect 24875 -5428 24971 -5412
rect 25594 -5412 25610 -5330
rect 25674 -5070 26329 -5044
rect 25674 -5330 25829 -5070
rect 25674 -5412 25690 -5330
rect 25828 -5390 25829 -5330
rect 26149 -5330 26329 -5070
rect 26149 -5390 26150 -5330
rect 25828 -5391 26150 -5390
rect 25594 -5428 25690 -5412
rect 26313 -5412 26329 -5330
rect 26393 -5070 37828 -5044
rect 26393 -5330 26548 -5070
rect 26393 -5412 26418 -5330
rect 26547 -5390 26548 -5330
rect 26868 -5192 37828 -5070
rect 26868 -5278 27682 -5192
rect 27778 -5278 28282 -5192
rect 28378 -5278 28882 -5192
rect 28978 -5278 29482 -5192
rect 29578 -5278 30082 -5192
rect 30178 -5278 30682 -5192
rect 30778 -5278 31282 -5192
rect 31378 -5278 31882 -5192
rect 31978 -5278 32482 -5192
rect 32578 -5278 33082 -5192
rect 33178 -5278 33682 -5192
rect 33778 -5278 34282 -5192
rect 34378 -5278 34882 -5192
rect 34978 -5278 35482 -5192
rect 35578 -5278 36082 -5192
rect 36178 -5278 36682 -5192
rect 36778 -5278 37262 -5192
rect 37358 -5278 37828 -5192
rect 26868 -5330 37828 -5278
rect 26868 -5390 26869 -5330
rect 26547 -5391 26869 -5390
rect 26313 -5428 26418 -5412
rect 24496 -5626 26040 -5526
rect 23671 -5770 23993 -5769
rect 23671 -5884 23672 -5770
rect 23517 -5984 23672 -5884
rect 23517 -6112 23540 -5984
rect 23671 -6090 23672 -5984
rect 23992 -5884 23993 -5770
rect 24150 -5884 24172 -5744
rect 23992 -5984 24172 -5884
rect 23992 -6090 23993 -5984
rect 23671 -6091 23993 -6090
rect 23437 -6128 23540 -6112
rect 23440 -6426 23540 -6128
rect 23437 -6444 23540 -6426
rect 11547 -6470 11869 -6469
rect 11547 -6582 11548 -6470
rect 11393 -6682 11548 -6582
rect 11393 -6792 11418 -6682
rect 11547 -6790 11548 -6682
rect 11868 -6790 11869 -6470
rect 11547 -6791 11869 -6790
rect 11654 -6792 11754 -6791
rect 11393 -6812 11409 -6792
rect 11313 -6828 11409 -6812
rect 23437 -6812 23453 -6444
rect 23517 -6576 23540 -6444
rect 23778 -6469 23878 -6091
rect 24150 -6112 24172 -5984
rect 24236 -6112 24252 -5744
rect 24497 -5769 24598 -5626
rect 24875 -5744 24971 -5726
rect 24390 -5770 24712 -5769
rect 24390 -6090 24391 -5770
rect 24711 -6090 24712 -5770
rect 24390 -6091 24712 -6090
rect 24150 -6128 24252 -6112
rect 24150 -6426 24250 -6128
rect 24497 -6226 24598 -6091
rect 24875 -6112 24891 -5744
rect 24955 -6112 24971 -5744
rect 25220 -5769 25320 -5626
rect 25594 -5744 25690 -5726
rect 25109 -5770 25431 -5769
rect 25109 -6090 25110 -5770
rect 25430 -6090 25431 -5770
rect 25109 -6091 25431 -6090
rect 24875 -6128 24971 -6112
rect 25220 -6226 25320 -6091
rect 25594 -6112 25610 -5744
rect 25674 -6112 25690 -5744
rect 25940 -5769 26040 -5626
rect 26318 -5726 26418 -5428
rect 26313 -5744 26418 -5726
rect 25828 -5770 26150 -5769
rect 25828 -6090 25829 -5770
rect 26149 -6090 26150 -5770
rect 25828 -6091 26150 -6090
rect 25594 -6128 25690 -6112
rect 25940 -6226 26040 -6091
rect 26313 -6112 26329 -5744
rect 26393 -5876 26418 -5744
rect 26654 -5769 26754 -5391
rect 26547 -5770 26869 -5769
rect 26547 -5876 26548 -5770
rect 26393 -5976 26548 -5876
rect 26393 -6112 26418 -5976
rect 26547 -6090 26548 -5976
rect 26868 -6090 26869 -5770
rect 26547 -6091 26869 -6090
rect 26313 -6128 26418 -6112
rect 24497 -6326 26040 -6226
rect 24150 -6444 24252 -6426
rect 23671 -6470 23993 -6469
rect 23671 -6576 23672 -6470
rect 23517 -6676 23672 -6576
rect 23517 -6812 23540 -6676
rect 23671 -6790 23672 -6676
rect 23992 -6576 23993 -6470
rect 24150 -6576 24172 -6444
rect 23992 -6676 24172 -6576
rect 23992 -6790 23993 -6676
rect 23671 -6791 23993 -6790
rect 23778 -6792 23878 -6791
rect 23437 -6828 23540 -6812
rect 23440 -6830 23540 -6828
rect 24150 -6812 24172 -6676
rect 24236 -6812 24252 -6444
rect 24497 -6469 24598 -6326
rect 24875 -6444 24971 -6426
rect 24390 -6470 24712 -6469
rect 24390 -6790 24391 -6470
rect 24711 -6790 24712 -6470
rect 24390 -6791 24712 -6790
rect 24150 -6828 24252 -6812
rect 24150 -6830 24250 -6828
rect 24497 -6928 24598 -6791
rect 24875 -6812 24891 -6444
rect 24955 -6812 24971 -6444
rect 25220 -6469 25320 -6326
rect 25594 -6444 25690 -6426
rect 25109 -6470 25431 -6469
rect 25109 -6790 25110 -6470
rect 25430 -6790 25431 -6470
rect 25109 -6791 25431 -6790
rect 24875 -6828 24971 -6812
rect 25220 -6928 25320 -6791
rect 25594 -6812 25610 -6444
rect 25674 -6812 25690 -6444
rect 25940 -6469 26040 -6326
rect 26318 -6426 26418 -6128
rect 26313 -6444 26418 -6426
rect 25828 -6470 26150 -6469
rect 25828 -6790 25829 -6470
rect 26149 -6790 26150 -6470
rect 25828 -6791 26150 -6790
rect 25594 -6828 25690 -6812
rect 25940 -6928 26040 -6791
rect 26313 -6812 26329 -6444
rect 26393 -6582 26418 -6444
rect 26654 -6469 26754 -6091
rect 26547 -6470 26869 -6469
rect 26547 -6582 26548 -6470
rect 26393 -6682 26548 -6582
rect 26393 -6792 26418 -6682
rect 26547 -6790 26548 -6682
rect 26868 -6790 26869 -6470
rect 26547 -6791 26869 -6790
rect 26654 -6792 26754 -6791
rect 26393 -6812 26409 -6792
rect 26313 -6828 26409 -6812
rect 8138 -6929 12230 -6928
rect 8138 -7027 8139 -6929
rect 8237 -7027 12131 -6929
rect 12229 -7027 12230 -6929
rect 8138 -7028 12230 -7027
rect 23130 -6929 27230 -6928
rect 23130 -7027 23131 -6929
rect 23229 -7027 27131 -6929
rect 27229 -7027 27230 -6929
rect 23130 -7028 27230 -7027
rect 8437 -7130 8533 -7124
rect 9156 -7130 9252 -7124
rect 8437 -7144 8540 -7130
rect 8437 -7512 8453 -7144
rect 8517 -7280 8540 -7144
rect 9150 -7144 9252 -7130
rect 8778 -7169 8878 -7168
rect 8671 -7170 8993 -7169
rect 8671 -7280 8672 -7170
rect 8517 -7380 8672 -7280
rect 8517 -7512 8540 -7380
rect 8671 -7490 8672 -7380
rect 8992 -7280 8993 -7170
rect 9150 -7280 9172 -7144
rect 8992 -7380 9172 -7280
rect 8992 -7490 8993 -7380
rect 8671 -7491 8993 -7490
rect 8437 -7842 8540 -7512
rect 8437 -8212 8453 -7842
rect 8517 -7974 8540 -7842
rect 8778 -7869 8878 -7491
rect 9150 -7512 9172 -7380
rect 9236 -7512 9252 -7144
rect 9497 -7169 9598 -7028
rect 9875 -7144 9971 -7124
rect 9390 -7170 9712 -7169
rect 9390 -7490 9391 -7170
rect 9711 -7490 9712 -7170
rect 9390 -7491 9712 -7490
rect 9150 -7842 9252 -7512
rect 9497 -7620 9598 -7491
rect 9875 -7512 9891 -7144
rect 9955 -7512 9971 -7144
rect 10220 -7169 10320 -7028
rect 10594 -7144 10690 -7124
rect 10109 -7170 10431 -7169
rect 10109 -7490 10110 -7170
rect 10430 -7490 10431 -7170
rect 10109 -7491 10431 -7490
rect 9875 -7528 9971 -7512
rect 10220 -7620 10320 -7491
rect 10594 -7512 10610 -7144
rect 10674 -7512 10690 -7144
rect 10940 -7169 11040 -7028
rect 11313 -7144 11409 -7124
rect 10828 -7170 11150 -7169
rect 10828 -7490 10829 -7170
rect 11149 -7490 11150 -7170
rect 10828 -7491 11150 -7490
rect 10594 -7528 10690 -7512
rect 10940 -7620 11040 -7491
rect 11313 -7512 11329 -7144
rect 11393 -7170 11409 -7144
rect 23437 -7130 23533 -7124
rect 24156 -7130 24252 -7124
rect 23437 -7144 23540 -7130
rect 11547 -7170 11869 -7169
rect 11393 -7284 11418 -7170
rect 11547 -7284 11548 -7170
rect 11393 -7384 11548 -7284
rect 11393 -7512 11418 -7384
rect 11547 -7490 11548 -7384
rect 11868 -7490 11869 -7170
rect 11547 -7491 11869 -7490
rect 11313 -7528 11418 -7512
rect 9496 -7720 11040 -7620
rect 11318 -7826 11418 -7528
rect 8671 -7870 8993 -7869
rect 8671 -7974 8672 -7870
rect 8517 -8074 8672 -7974
rect 8517 -8212 8533 -8074
rect 8671 -8190 8672 -8074
rect 8992 -7974 8993 -7870
rect 9150 -7974 9172 -7842
rect 8992 -8074 9172 -7974
rect 8992 -8190 8993 -8074
rect 8671 -8191 8993 -8190
rect 8437 -8228 8533 -8212
rect 9156 -8212 9172 -8074
rect 9236 -7974 9252 -7842
rect 9875 -7842 9971 -7826
rect 9390 -7870 9712 -7869
rect 9390 -7974 9391 -7870
rect 9236 -8074 9391 -7974
rect 9236 -8212 9252 -8074
rect 9390 -8190 9391 -8074
rect 9711 -7974 9712 -7870
rect 9875 -7974 9891 -7842
rect 9711 -8074 9891 -7974
rect 9711 -8190 9712 -8074
rect 9390 -8191 9712 -8190
rect 9156 -8228 9252 -8212
rect 9875 -8212 9891 -8074
rect 9955 -7974 9971 -7842
rect 10594 -7842 10690 -7826
rect 10109 -7870 10431 -7869
rect 10109 -7974 10110 -7870
rect 9955 -8074 10110 -7974
rect 9955 -8212 9971 -8074
rect 10109 -8190 10110 -8074
rect 10430 -7974 10431 -7870
rect 10594 -7974 10610 -7842
rect 10430 -8074 10610 -7974
rect 10430 -8190 10431 -8074
rect 10109 -8191 10431 -8190
rect 9875 -8228 9971 -8212
rect 10594 -8212 10610 -8074
rect 10674 -7974 10690 -7842
rect 11313 -7842 11418 -7826
rect 10828 -7870 11150 -7869
rect 10828 -7974 10829 -7870
rect 10674 -8074 10829 -7974
rect 10674 -8212 10690 -8074
rect 10828 -8190 10829 -8074
rect 11149 -7974 11150 -7870
rect 11313 -7974 11329 -7842
rect 11149 -8074 11329 -7974
rect 11149 -8190 11150 -8074
rect 10828 -8191 11150 -8190
rect 10594 -8228 10690 -8212
rect 11313 -8214 11329 -8074
rect 11393 -7974 11418 -7842
rect 11654 -7869 11754 -7491
rect 23437 -7512 23453 -7144
rect 23517 -7280 23540 -7144
rect 24150 -7144 24252 -7130
rect 23778 -7169 23878 -7168
rect 23671 -7170 23993 -7169
rect 23671 -7280 23672 -7170
rect 23517 -7380 23672 -7280
rect 23517 -7512 23540 -7380
rect 23671 -7490 23672 -7380
rect 23992 -7280 23993 -7170
rect 24150 -7280 24172 -7144
rect 23992 -7380 24172 -7280
rect 23992 -7490 23993 -7380
rect 23671 -7491 23993 -7490
rect 23437 -7842 23540 -7512
rect 11547 -7870 11869 -7869
rect 11547 -7974 11548 -7870
rect 11393 -8074 11548 -7974
rect 11393 -8214 11409 -8074
rect 11547 -8190 11548 -8074
rect 11868 -8190 11869 -7870
rect 11547 -8191 11869 -8190
rect 11313 -8230 11409 -8214
rect 23437 -8212 23453 -7842
rect 23517 -7974 23540 -7842
rect 23778 -7869 23878 -7491
rect 24150 -7512 24172 -7380
rect 24236 -7512 24252 -7144
rect 24497 -7169 24598 -7028
rect 24875 -7144 24971 -7124
rect 24390 -7170 24712 -7169
rect 24390 -7490 24391 -7170
rect 24711 -7490 24712 -7170
rect 24390 -7491 24712 -7490
rect 24150 -7842 24252 -7512
rect 24497 -7620 24598 -7491
rect 24875 -7512 24891 -7144
rect 24955 -7512 24971 -7144
rect 25220 -7169 25320 -7028
rect 25594 -7144 25690 -7124
rect 25109 -7170 25431 -7169
rect 25109 -7490 25110 -7170
rect 25430 -7490 25431 -7170
rect 25109 -7491 25431 -7490
rect 24875 -7528 24971 -7512
rect 25220 -7620 25320 -7491
rect 25594 -7512 25610 -7144
rect 25674 -7512 25690 -7144
rect 25940 -7169 26040 -7028
rect 26313 -7144 26409 -7124
rect 25828 -7170 26150 -7169
rect 25828 -7490 25829 -7170
rect 26149 -7490 26150 -7170
rect 25828 -7491 26150 -7490
rect 25594 -7528 25690 -7512
rect 25940 -7620 26040 -7491
rect 26313 -7512 26329 -7144
rect 26393 -7170 26409 -7144
rect 26547 -7170 26869 -7169
rect 26393 -7284 26418 -7170
rect 26547 -7284 26548 -7170
rect 26393 -7384 26548 -7284
rect 26393 -7512 26418 -7384
rect 26547 -7490 26548 -7384
rect 26868 -7490 26869 -7170
rect 26547 -7491 26869 -7490
rect 26313 -7528 26418 -7512
rect 24496 -7720 26040 -7620
rect 26318 -7826 26418 -7528
rect 23671 -7870 23993 -7869
rect 23671 -7974 23672 -7870
rect 23517 -8074 23672 -7974
rect 23517 -8212 23533 -8074
rect 23671 -8190 23672 -8074
rect 23992 -7974 23993 -7870
rect 24150 -7974 24172 -7842
rect 23992 -8074 24172 -7974
rect 23992 -8190 23993 -8074
rect 23671 -8191 23993 -8190
rect 23437 -8228 23533 -8212
rect 24156 -8212 24172 -8074
rect 24236 -7974 24252 -7842
rect 24875 -7842 24971 -7826
rect 24390 -7870 24712 -7869
rect 24390 -7974 24391 -7870
rect 24236 -8074 24391 -7974
rect 24236 -8212 24252 -8074
rect 24390 -8190 24391 -8074
rect 24711 -7974 24712 -7870
rect 24875 -7974 24891 -7842
rect 24711 -8074 24891 -7974
rect 24711 -8190 24712 -8074
rect 24390 -8191 24712 -8190
rect 24156 -8228 24252 -8212
rect 24875 -8212 24891 -8074
rect 24955 -7974 24971 -7842
rect 25594 -7842 25690 -7826
rect 25109 -7870 25431 -7869
rect 25109 -7974 25110 -7870
rect 24955 -8074 25110 -7974
rect 24955 -8212 24971 -8074
rect 25109 -8190 25110 -8074
rect 25430 -7974 25431 -7870
rect 25594 -7974 25610 -7842
rect 25430 -8074 25610 -7974
rect 25430 -8190 25431 -8074
rect 25109 -8191 25431 -8190
rect 24875 -8228 24971 -8212
rect 25594 -8212 25610 -8074
rect 25674 -7974 25690 -7842
rect 26313 -7842 26418 -7826
rect 25828 -7870 26150 -7869
rect 25828 -7974 25829 -7870
rect 25674 -8074 25829 -7974
rect 25674 -8212 25690 -8074
rect 25828 -8190 25829 -8074
rect 26149 -7974 26150 -7870
rect 26313 -7974 26329 -7842
rect 26149 -8074 26329 -7974
rect 26149 -8190 26150 -8074
rect 25828 -8191 26150 -8190
rect 25594 -8228 25690 -8212
rect 26313 -8214 26329 -8074
rect 26393 -7974 26418 -7842
rect 26654 -7869 26754 -7491
rect 26547 -7870 26869 -7869
rect 26547 -7974 26548 -7870
rect 26393 -8074 26548 -7974
rect 26393 -8214 26409 -8074
rect 26547 -8190 26548 -8074
rect 26868 -8190 26869 -7870
rect 26547 -8191 26869 -8190
rect 26313 -8230 26409 -8214
rect 8274 -12456 38738 -12426
rect 8274 -12486 37966 -12456
rect 8274 -12572 13476 -12486
rect 13572 -12572 13896 -12486
rect 13992 -12572 14496 -12486
rect 14592 -12572 15096 -12486
rect 15192 -12572 15696 -12486
rect 15792 -12572 16296 -12486
rect 16392 -12572 16896 -12486
rect 16992 -12572 17496 -12486
rect 17592 -12572 18096 -12486
rect 18192 -12572 18696 -12486
rect 18792 -12572 19296 -12486
rect 19392 -12572 19896 -12486
rect 19992 -12572 20496 -12486
rect 20592 -12572 21096 -12486
rect 21192 -12572 21696 -12486
rect 21792 -12572 28476 -12486
rect 28572 -12572 28896 -12486
rect 28992 -12572 29496 -12486
rect 29592 -12572 30096 -12486
rect 30192 -12572 30696 -12486
rect 30792 -12572 31296 -12486
rect 31392 -12572 31896 -12486
rect 31992 -12572 32496 -12486
rect 32592 -12572 33096 -12486
rect 33192 -12572 33696 -12486
rect 33792 -12572 34296 -12486
rect 34392 -12572 34896 -12486
rect 34992 -12572 35496 -12486
rect 35592 -12572 36096 -12486
rect 36192 -12572 36696 -12486
rect 36792 -12572 37966 -12486
rect 8274 -12746 37966 -12572
rect 8274 -13046 12412 -12746
rect 13012 -13046 22044 -12746
rect 22644 -13046 27412 -12746
rect 28012 -13046 37044 -12746
rect 37644 -13046 37966 -12746
rect 8274 -13710 37966 -13046
rect 8274 -14010 8458 -13710
rect 9058 -14010 18090 -13710
rect 18690 -14010 23458 -13710
rect 24058 -14010 33090 -13710
rect 33690 -14010 37966 -13710
rect 8274 -14184 37966 -14010
rect 8274 -14270 9310 -14184
rect 9406 -14270 9910 -14184
rect 10006 -14270 10510 -14184
rect 10606 -14270 11110 -14184
rect 11206 -14270 11710 -14184
rect 11806 -14270 12310 -14184
rect 12406 -14270 12910 -14184
rect 13006 -14270 13510 -14184
rect 13606 -14270 14110 -14184
rect 14206 -14270 14710 -14184
rect 14806 -14270 15310 -14184
rect 15406 -14270 15910 -14184
rect 16006 -14270 16510 -14184
rect 16606 -14270 17110 -14184
rect 17206 -14270 17530 -14184
rect 17626 -14270 24310 -14184
rect 24406 -14270 24910 -14184
rect 25006 -14270 25510 -14184
rect 25606 -14270 26110 -14184
rect 26206 -14270 26710 -14184
rect 26806 -14270 27310 -14184
rect 27406 -14270 27910 -14184
rect 28006 -14270 28510 -14184
rect 28606 -14270 29110 -14184
rect 29206 -14270 29710 -14184
rect 29806 -14270 30310 -14184
rect 30406 -14270 30910 -14184
rect 31006 -14270 31510 -14184
rect 31606 -14270 32110 -14184
rect 32206 -14270 32530 -14184
rect 32626 -14270 37966 -14184
rect 8274 -14302 37966 -14270
rect 38700 -14302 38738 -12456
rect 8274 -14328 38738 -14302
rect 19693 -18542 19789 -18526
rect 19233 -18566 19555 -18565
rect 19233 -18886 19234 -18566
rect 19554 -18682 19555 -18566
rect 19693 -18682 19709 -18542
rect 19554 -18782 19709 -18682
rect 19554 -18886 19555 -18782
rect 19233 -18887 19555 -18886
rect 19348 -19265 19448 -18887
rect 19684 -18914 19709 -18782
rect 19773 -18682 19789 -18542
rect 20412 -18544 20508 -18528
rect 19952 -18566 20274 -18565
rect 19952 -18682 19953 -18566
rect 19773 -18782 19953 -18682
rect 19773 -18914 19789 -18782
rect 19952 -18886 19953 -18782
rect 20273 -18682 20274 -18566
rect 20412 -18682 20428 -18544
rect 20273 -18782 20428 -18682
rect 20273 -18886 20274 -18782
rect 19952 -18887 20274 -18886
rect 19684 -18930 19789 -18914
rect 20412 -18914 20428 -18782
rect 20492 -18682 20508 -18544
rect 21131 -18544 21227 -18528
rect 20671 -18566 20993 -18565
rect 20671 -18682 20672 -18566
rect 20492 -18782 20672 -18682
rect 20492 -18914 20508 -18782
rect 20671 -18886 20672 -18782
rect 20992 -18682 20993 -18566
rect 21131 -18682 21147 -18544
rect 20992 -18782 21147 -18682
rect 20992 -18886 20993 -18782
rect 20671 -18887 20993 -18886
rect 20412 -18930 20508 -18914
rect 21131 -18914 21147 -18782
rect 21211 -18682 21227 -18544
rect 21850 -18544 21946 -18528
rect 21390 -18566 21712 -18565
rect 21390 -18682 21391 -18566
rect 21211 -18782 21391 -18682
rect 21211 -18914 21227 -18782
rect 21390 -18886 21391 -18782
rect 21711 -18682 21712 -18566
rect 21850 -18682 21866 -18544
rect 21711 -18782 21866 -18682
rect 21711 -18886 21712 -18782
rect 21390 -18887 21712 -18886
rect 21131 -18930 21227 -18914
rect 21850 -18914 21866 -18782
rect 21930 -18682 21946 -18544
rect 22569 -18544 22665 -18528
rect 22109 -18566 22431 -18565
rect 22109 -18682 22110 -18566
rect 21930 -18782 22110 -18682
rect 21930 -18914 21952 -18782
rect 22109 -18886 22110 -18782
rect 22430 -18682 22431 -18566
rect 22569 -18682 22585 -18544
rect 22430 -18782 22585 -18682
rect 22430 -18886 22431 -18782
rect 22109 -18887 22431 -18886
rect 19684 -19228 19784 -18930
rect 20062 -19136 21606 -19036
rect 19684 -19244 19789 -19228
rect 19233 -19266 19555 -19265
rect 19233 -19586 19234 -19266
rect 19554 -19372 19555 -19266
rect 19684 -19372 19709 -19244
rect 19554 -19472 19709 -19372
rect 19554 -19586 19555 -19472
rect 19684 -19586 19709 -19472
rect 19233 -19587 19555 -19586
rect 19693 -19612 19709 -19586
rect 19773 -19612 19789 -19244
rect 20062 -19265 20162 -19136
rect 20412 -19244 20508 -19228
rect 19952 -19266 20274 -19265
rect 19952 -19586 19953 -19266
rect 20273 -19586 20274 -19266
rect 19952 -19587 20274 -19586
rect 19693 -19632 19789 -19612
rect 20062 -19728 20162 -19587
rect 20412 -19612 20428 -19244
rect 20492 -19612 20508 -19244
rect 20782 -19265 20882 -19136
rect 21131 -19244 21227 -19228
rect 20671 -19266 20993 -19265
rect 20671 -19586 20672 -19266
rect 20992 -19586 20993 -19266
rect 20671 -19587 20993 -19586
rect 20412 -19632 20508 -19612
rect 20782 -19728 20882 -19587
rect 21131 -19612 21147 -19244
rect 21211 -19612 21227 -19244
rect 21504 -19265 21605 -19136
rect 21850 -19244 21952 -18914
rect 21390 -19266 21712 -19265
rect 21390 -19586 21391 -19266
rect 21711 -19586 21712 -19266
rect 21390 -19587 21712 -19586
rect 21131 -19632 21227 -19612
rect 21504 -19728 21605 -19587
rect 21850 -19612 21866 -19244
rect 21930 -19376 21952 -19244
rect 22224 -19265 22324 -18887
rect 22562 -18914 22585 -18782
rect 22649 -18914 22665 -18544
rect 34693 -18542 34789 -18526
rect 34233 -18566 34555 -18565
rect 34233 -18886 34234 -18566
rect 34554 -18682 34555 -18566
rect 34693 -18682 34709 -18542
rect 34554 -18782 34709 -18682
rect 34554 -18886 34555 -18782
rect 34233 -18887 34555 -18886
rect 22562 -19244 22665 -18914
rect 22109 -19266 22431 -19265
rect 22109 -19376 22110 -19266
rect 21930 -19476 22110 -19376
rect 21930 -19612 21952 -19476
rect 22109 -19586 22110 -19476
rect 22430 -19376 22431 -19266
rect 22562 -19376 22585 -19244
rect 22430 -19476 22585 -19376
rect 22430 -19586 22431 -19476
rect 22109 -19587 22431 -19586
rect 22224 -19588 22324 -19587
rect 21850 -19626 21952 -19612
rect 22562 -19612 22585 -19476
rect 22649 -19612 22665 -19244
rect 34348 -19265 34448 -18887
rect 34684 -18914 34709 -18782
rect 34773 -18682 34789 -18542
rect 35412 -18544 35508 -18528
rect 34952 -18566 35274 -18565
rect 34952 -18682 34953 -18566
rect 34773 -18782 34953 -18682
rect 34773 -18914 34789 -18782
rect 34952 -18886 34953 -18782
rect 35273 -18682 35274 -18566
rect 35412 -18682 35428 -18544
rect 35273 -18782 35428 -18682
rect 35273 -18886 35274 -18782
rect 34952 -18887 35274 -18886
rect 34684 -18930 34789 -18914
rect 35412 -18914 35428 -18782
rect 35492 -18682 35508 -18544
rect 36131 -18544 36227 -18528
rect 35671 -18566 35993 -18565
rect 35671 -18682 35672 -18566
rect 35492 -18782 35672 -18682
rect 35492 -18914 35508 -18782
rect 35671 -18886 35672 -18782
rect 35992 -18682 35993 -18566
rect 36131 -18682 36147 -18544
rect 35992 -18782 36147 -18682
rect 35992 -18886 35993 -18782
rect 35671 -18887 35993 -18886
rect 35412 -18930 35508 -18914
rect 36131 -18914 36147 -18782
rect 36211 -18682 36227 -18544
rect 36850 -18544 36946 -18528
rect 36390 -18566 36712 -18565
rect 36390 -18682 36391 -18566
rect 36211 -18782 36391 -18682
rect 36211 -18914 36227 -18782
rect 36390 -18886 36391 -18782
rect 36711 -18682 36712 -18566
rect 36850 -18682 36866 -18544
rect 36711 -18782 36866 -18682
rect 36711 -18886 36712 -18782
rect 36390 -18887 36712 -18886
rect 36131 -18930 36227 -18914
rect 36850 -18914 36866 -18782
rect 36930 -18682 36946 -18544
rect 37569 -18544 37665 -18528
rect 37109 -18566 37431 -18565
rect 37109 -18682 37110 -18566
rect 36930 -18782 37110 -18682
rect 36930 -18914 36952 -18782
rect 37109 -18886 37110 -18782
rect 37430 -18682 37431 -18566
rect 37569 -18682 37585 -18544
rect 37430 -18782 37585 -18682
rect 37430 -18886 37431 -18782
rect 37109 -18887 37431 -18886
rect 34684 -19228 34784 -18930
rect 35062 -19136 36606 -19036
rect 34684 -19244 34789 -19228
rect 34233 -19266 34555 -19265
rect 34233 -19586 34234 -19266
rect 34554 -19372 34555 -19266
rect 34684 -19372 34709 -19244
rect 34554 -19472 34709 -19372
rect 34554 -19586 34555 -19472
rect 34684 -19586 34709 -19472
rect 34233 -19587 34555 -19586
rect 22562 -19626 22665 -19612
rect 21850 -19632 21946 -19626
rect 22569 -19632 22665 -19626
rect 34693 -19612 34709 -19586
rect 34773 -19612 34789 -19244
rect 35062 -19265 35162 -19136
rect 35412 -19244 35508 -19228
rect 34952 -19266 35274 -19265
rect 34952 -19586 34953 -19266
rect 35273 -19586 35274 -19266
rect 34952 -19587 35274 -19586
rect 34693 -19632 34789 -19612
rect 35062 -19728 35162 -19587
rect 35412 -19612 35428 -19244
rect 35492 -19612 35508 -19244
rect 35782 -19265 35882 -19136
rect 36131 -19244 36227 -19228
rect 35671 -19266 35993 -19265
rect 35671 -19586 35672 -19266
rect 35992 -19586 35993 -19266
rect 35671 -19587 35993 -19586
rect 35412 -19632 35508 -19612
rect 35782 -19728 35882 -19587
rect 36131 -19612 36147 -19244
rect 36211 -19612 36227 -19244
rect 36504 -19265 36605 -19136
rect 36850 -19244 36952 -18914
rect 36390 -19266 36712 -19265
rect 36390 -19586 36391 -19266
rect 36711 -19586 36712 -19266
rect 36390 -19587 36712 -19586
rect 36131 -19632 36227 -19612
rect 36504 -19728 36605 -19587
rect 36850 -19612 36866 -19244
rect 36930 -19376 36952 -19244
rect 37224 -19265 37324 -18887
rect 37562 -18914 37585 -18782
rect 37649 -18914 37665 -18544
rect 37562 -19244 37665 -18914
rect 37109 -19266 37431 -19265
rect 37109 -19376 37110 -19266
rect 36930 -19476 37110 -19376
rect 36930 -19612 36952 -19476
rect 37109 -19586 37110 -19476
rect 37430 -19376 37431 -19266
rect 37562 -19376 37585 -19244
rect 37430 -19476 37585 -19376
rect 37430 -19586 37431 -19476
rect 37109 -19587 37431 -19586
rect 37224 -19588 37324 -19587
rect 36850 -19626 36952 -19612
rect 37562 -19612 37585 -19476
rect 37649 -19612 37665 -19244
rect 37562 -19626 37665 -19612
rect 36850 -19632 36946 -19626
rect 37569 -19632 37665 -19626
rect 18872 -19729 23036 -19728
rect 18872 -19827 18873 -19729
rect 18971 -19827 22937 -19729
rect 23035 -19827 23036 -19729
rect 18872 -19828 23036 -19827
rect 33872 -19729 37934 -19728
rect 33872 -19827 33873 -19729
rect 33971 -19827 37835 -19729
rect 37933 -19827 37934 -19729
rect 33872 -19828 37934 -19827
rect 19693 -19944 19789 -19928
rect 19693 -19964 19709 -19944
rect 19348 -19965 19448 -19964
rect 19233 -19966 19555 -19965
rect 19233 -20286 19234 -19966
rect 19554 -20074 19555 -19966
rect 19684 -20074 19709 -19964
rect 19554 -20174 19709 -20074
rect 19554 -20286 19555 -20174
rect 19233 -20287 19555 -20286
rect 19348 -20665 19448 -20287
rect 19684 -20312 19709 -20174
rect 19773 -20312 19789 -19944
rect 20062 -19965 20162 -19828
rect 20412 -19944 20508 -19928
rect 19952 -19966 20274 -19965
rect 19952 -20286 19953 -19966
rect 20273 -20286 20274 -19966
rect 19952 -20287 20274 -20286
rect 19684 -20330 19789 -20312
rect 19684 -20628 19784 -20330
rect 20062 -20430 20162 -20287
rect 20412 -20312 20428 -19944
rect 20492 -20312 20508 -19944
rect 20782 -19965 20882 -19828
rect 21131 -19944 21227 -19928
rect 20671 -19966 20993 -19965
rect 20671 -20286 20672 -19966
rect 20992 -20286 20993 -19966
rect 20671 -20287 20993 -20286
rect 20412 -20330 20508 -20312
rect 20782 -20430 20882 -20287
rect 21131 -20312 21147 -19944
rect 21211 -20312 21227 -19944
rect 21504 -19965 21605 -19828
rect 21852 -19928 21952 -19926
rect 21850 -19944 21952 -19928
rect 21390 -19966 21712 -19965
rect 21390 -20286 21391 -19966
rect 21711 -20286 21712 -19966
rect 21390 -20287 21712 -20286
rect 21131 -20330 21227 -20312
rect 21504 -20430 21605 -20287
rect 21850 -20312 21866 -19944
rect 21930 -20080 21952 -19944
rect 22562 -19928 22662 -19926
rect 22562 -19944 22665 -19928
rect 22224 -19965 22324 -19964
rect 22109 -19966 22431 -19965
rect 22109 -20080 22110 -19966
rect 21930 -20180 22110 -20080
rect 21930 -20312 21952 -20180
rect 22109 -20286 22110 -20180
rect 22430 -20080 22431 -19966
rect 22562 -20080 22585 -19944
rect 22430 -20180 22585 -20080
rect 22430 -20286 22431 -20180
rect 22109 -20287 22431 -20286
rect 21850 -20330 21952 -20312
rect 20062 -20530 21605 -20430
rect 19684 -20644 19789 -20628
rect 19233 -20666 19555 -20665
rect 19233 -20986 19234 -20666
rect 19554 -20780 19555 -20666
rect 19684 -20780 19709 -20644
rect 19554 -20880 19709 -20780
rect 19554 -20986 19555 -20880
rect 19233 -20987 19555 -20986
rect 19348 -21365 19448 -20987
rect 19684 -21012 19709 -20880
rect 19773 -21012 19789 -20644
rect 20062 -20665 20162 -20530
rect 20412 -20644 20508 -20628
rect 19952 -20666 20274 -20665
rect 19952 -20986 19953 -20666
rect 20273 -20986 20274 -20666
rect 19952 -20987 20274 -20986
rect 19684 -21030 19789 -21012
rect 19684 -21328 19784 -21030
rect 20062 -21130 20162 -20987
rect 20412 -21012 20428 -20644
rect 20492 -21012 20508 -20644
rect 20782 -20665 20882 -20530
rect 21131 -20644 21227 -20628
rect 20671 -20666 20993 -20665
rect 20671 -20986 20672 -20666
rect 20992 -20986 20993 -20666
rect 20671 -20987 20993 -20986
rect 20412 -21030 20508 -21012
rect 20782 -21130 20882 -20987
rect 21131 -21012 21147 -20644
rect 21211 -21012 21227 -20644
rect 21504 -20665 21605 -20530
rect 21852 -20628 21952 -20330
rect 21850 -20644 21952 -20628
rect 21390 -20666 21712 -20665
rect 21390 -20986 21391 -20666
rect 21711 -20986 21712 -20666
rect 21390 -20987 21712 -20986
rect 21131 -21030 21227 -21012
rect 21504 -21130 21605 -20987
rect 21850 -21012 21866 -20644
rect 21930 -20772 21952 -20644
rect 22224 -20665 22324 -20287
rect 22562 -20312 22585 -20180
rect 22649 -20312 22665 -19944
rect 34693 -19944 34789 -19928
rect 34693 -19964 34709 -19944
rect 34348 -19965 34448 -19964
rect 34233 -19966 34555 -19965
rect 34233 -20286 34234 -19966
rect 34554 -20074 34555 -19966
rect 34684 -20074 34709 -19964
rect 34554 -20174 34709 -20074
rect 34554 -20286 34555 -20174
rect 34233 -20287 34555 -20286
rect 22562 -20330 22665 -20312
rect 22562 -20628 22662 -20330
rect 22562 -20644 22665 -20628
rect 22109 -20666 22431 -20665
rect 22109 -20772 22110 -20666
rect 21930 -20872 22110 -20772
rect 21930 -21012 21952 -20872
rect 22109 -20986 22110 -20872
rect 22430 -20772 22431 -20666
rect 22562 -20772 22585 -20644
rect 22430 -20872 22585 -20772
rect 22430 -20986 22431 -20872
rect 22109 -20987 22431 -20986
rect 20062 -21230 21606 -21130
rect 19684 -21344 19789 -21328
rect 19233 -21366 19555 -21365
rect 19233 -21426 19234 -21366
rect 8120 -21478 19234 -21426
rect 8120 -21564 8744 -21478
rect 8840 -21564 9324 -21478
rect 9420 -21564 9924 -21478
rect 10020 -21564 10524 -21478
rect 10620 -21564 11124 -21478
rect 11220 -21564 11724 -21478
rect 11820 -21564 12324 -21478
rect 12420 -21564 12924 -21478
rect 13020 -21564 13524 -21478
rect 13620 -21564 14124 -21478
rect 14220 -21564 14724 -21478
rect 14820 -21564 15324 -21478
rect 15420 -21564 15924 -21478
rect 16020 -21564 16524 -21478
rect 16620 -21564 17124 -21478
rect 17220 -21564 17724 -21478
rect 17820 -21564 18324 -21478
rect 18420 -21564 19234 -21478
rect 8120 -21686 19234 -21564
rect 19554 -21426 19555 -21366
rect 19684 -21426 19709 -21344
rect 19554 -21686 19709 -21426
rect 8120 -21712 19709 -21686
rect 19773 -21426 19789 -21344
rect 20412 -21344 20508 -21328
rect 19952 -21366 20274 -21365
rect 19952 -21426 19953 -21366
rect 19773 -21686 19953 -21426
rect 20273 -21426 20274 -21366
rect 20412 -21426 20428 -21344
rect 20273 -21686 20428 -21426
rect 19773 -21712 20428 -21686
rect 20492 -21426 20508 -21344
rect 21131 -21344 21227 -21328
rect 20671 -21366 20993 -21365
rect 20671 -21426 20672 -21366
rect 20492 -21686 20672 -21426
rect 20992 -21426 20993 -21366
rect 21131 -21426 21147 -21344
rect 20992 -21686 21147 -21426
rect 20492 -21712 21147 -21686
rect 21211 -21426 21227 -21344
rect 21850 -21344 21952 -21012
rect 21390 -21366 21712 -21365
rect 21390 -21426 21391 -21366
rect 21211 -21686 21391 -21426
rect 21711 -21426 21712 -21366
rect 21850 -21426 21866 -21344
rect 21711 -21686 21866 -21426
rect 21211 -21712 21866 -21686
rect 21930 -21426 21952 -21344
rect 22224 -21365 22324 -20987
rect 22562 -21012 22585 -20872
rect 22649 -21012 22665 -20644
rect 34348 -20665 34448 -20287
rect 34684 -20312 34709 -20174
rect 34773 -20312 34789 -19944
rect 35062 -19965 35162 -19828
rect 35412 -19944 35508 -19928
rect 34952 -19966 35274 -19965
rect 34952 -20286 34953 -19966
rect 35273 -20286 35274 -19966
rect 34952 -20287 35274 -20286
rect 34684 -20330 34789 -20312
rect 34684 -20628 34784 -20330
rect 35062 -20430 35162 -20287
rect 35412 -20312 35428 -19944
rect 35492 -20312 35508 -19944
rect 35782 -19965 35882 -19828
rect 36131 -19944 36227 -19928
rect 35671 -19966 35993 -19965
rect 35671 -20286 35672 -19966
rect 35992 -20286 35993 -19966
rect 35671 -20287 35993 -20286
rect 35412 -20330 35508 -20312
rect 35782 -20430 35882 -20287
rect 36131 -20312 36147 -19944
rect 36211 -20312 36227 -19944
rect 36504 -19965 36605 -19828
rect 36852 -19928 36952 -19926
rect 36850 -19944 36952 -19928
rect 36390 -19966 36712 -19965
rect 36390 -20286 36391 -19966
rect 36711 -20286 36712 -19966
rect 36390 -20287 36712 -20286
rect 36131 -20330 36227 -20312
rect 36504 -20430 36605 -20287
rect 36850 -20312 36866 -19944
rect 36930 -20080 36952 -19944
rect 37562 -19928 37662 -19926
rect 37562 -19944 37665 -19928
rect 37224 -19965 37324 -19964
rect 37109 -19966 37431 -19965
rect 37109 -20080 37110 -19966
rect 36930 -20180 37110 -20080
rect 36930 -20312 36952 -20180
rect 37109 -20286 37110 -20180
rect 37430 -20080 37431 -19966
rect 37562 -20080 37585 -19944
rect 37430 -20180 37585 -20080
rect 37430 -20286 37431 -20180
rect 37109 -20287 37431 -20286
rect 36850 -20330 36952 -20312
rect 35062 -20530 36605 -20430
rect 34684 -20644 34789 -20628
rect 34233 -20666 34555 -20665
rect 34233 -20986 34234 -20666
rect 34554 -20780 34555 -20666
rect 34684 -20780 34709 -20644
rect 34554 -20880 34709 -20780
rect 34554 -20986 34555 -20880
rect 34233 -20987 34555 -20986
rect 22562 -21344 22665 -21012
rect 22109 -21366 22431 -21365
rect 22109 -21426 22110 -21366
rect 21930 -21686 22110 -21426
rect 22430 -21426 22431 -21366
rect 22562 -21426 22585 -21344
rect 22430 -21686 22585 -21426
rect 21930 -21712 22585 -21686
rect 22649 -21426 22665 -21344
rect 34348 -21365 34448 -20987
rect 34684 -21012 34709 -20880
rect 34773 -21012 34789 -20644
rect 35062 -20665 35162 -20530
rect 35412 -20644 35508 -20628
rect 34952 -20666 35274 -20665
rect 34952 -20986 34953 -20666
rect 35273 -20986 35274 -20666
rect 34952 -20987 35274 -20986
rect 34684 -21030 34789 -21012
rect 34684 -21328 34784 -21030
rect 35062 -21130 35162 -20987
rect 35412 -21012 35428 -20644
rect 35492 -21012 35508 -20644
rect 35782 -20665 35882 -20530
rect 36131 -20644 36227 -20628
rect 35671 -20666 35993 -20665
rect 35671 -20986 35672 -20666
rect 35992 -20986 35993 -20666
rect 35671 -20987 35993 -20986
rect 35412 -21030 35508 -21012
rect 35782 -21130 35882 -20987
rect 36131 -21012 36147 -20644
rect 36211 -21012 36227 -20644
rect 36504 -20665 36605 -20530
rect 36852 -20628 36952 -20330
rect 36850 -20644 36952 -20628
rect 36390 -20666 36712 -20665
rect 36390 -20986 36391 -20666
rect 36711 -20986 36712 -20666
rect 36390 -20987 36712 -20986
rect 36131 -21030 36227 -21012
rect 36504 -21130 36605 -20987
rect 36850 -21012 36866 -20644
rect 36930 -20772 36952 -20644
rect 37224 -20665 37324 -20287
rect 37562 -20312 37585 -20180
rect 37649 -20312 37665 -19944
rect 37562 -20330 37665 -20312
rect 37562 -20628 37662 -20330
rect 37562 -20644 37665 -20628
rect 37109 -20666 37431 -20665
rect 37109 -20772 37110 -20666
rect 36930 -20872 37110 -20772
rect 36930 -21012 36952 -20872
rect 37109 -20986 37110 -20872
rect 37430 -20772 37431 -20666
rect 37562 -20772 37585 -20644
rect 37430 -20872 37585 -20772
rect 37430 -20986 37431 -20872
rect 37109 -20987 37431 -20986
rect 35062 -21230 36606 -21130
rect 34684 -21344 34789 -21328
rect 34233 -21366 34555 -21365
rect 34233 -21426 34234 -21366
rect 22649 -21478 34234 -21426
rect 22649 -21564 23744 -21478
rect 23840 -21564 24324 -21478
rect 24420 -21564 24924 -21478
rect 25020 -21564 25524 -21478
rect 25620 -21564 26124 -21478
rect 26220 -21564 26724 -21478
rect 26820 -21564 27324 -21478
rect 27420 -21564 27924 -21478
rect 28020 -21564 28524 -21478
rect 28620 -21564 29124 -21478
rect 29220 -21564 29724 -21478
rect 29820 -21564 30324 -21478
rect 30420 -21564 30924 -21478
rect 31020 -21564 31524 -21478
rect 31620 -21564 32124 -21478
rect 32220 -21564 32724 -21478
rect 32820 -21564 33324 -21478
rect 33420 -21564 34234 -21478
rect 22649 -21686 34234 -21564
rect 34554 -21426 34555 -21366
rect 34684 -21426 34709 -21344
rect 34554 -21686 34709 -21426
rect 22649 -21712 34709 -21686
rect 34773 -21426 34789 -21344
rect 35412 -21344 35508 -21328
rect 34952 -21366 35274 -21365
rect 34952 -21426 34953 -21366
rect 34773 -21686 34953 -21426
rect 35273 -21426 35274 -21366
rect 35412 -21426 35428 -21344
rect 35273 -21686 35428 -21426
rect 34773 -21712 35428 -21686
rect 35492 -21426 35508 -21344
rect 36131 -21344 36227 -21328
rect 35671 -21366 35993 -21365
rect 35671 -21426 35672 -21366
rect 35492 -21686 35672 -21426
rect 35992 -21426 35993 -21366
rect 36131 -21426 36147 -21344
rect 35992 -21686 36147 -21426
rect 35492 -21712 36147 -21686
rect 36211 -21426 36227 -21344
rect 36850 -21344 36952 -21012
rect 36390 -21366 36712 -21365
rect 36390 -21426 36391 -21366
rect 36211 -21686 36391 -21426
rect 36711 -21426 36712 -21366
rect 36850 -21426 36866 -21344
rect 36711 -21686 36866 -21426
rect 36211 -21712 36866 -21686
rect 36930 -21426 36952 -21344
rect 37224 -21365 37324 -20987
rect 37562 -21012 37585 -20872
rect 37649 -21012 37665 -20644
rect 37562 -21344 37665 -21012
rect 37109 -21366 37431 -21365
rect 37109 -21426 37110 -21366
rect 36930 -21686 37110 -21426
rect 37430 -21426 37431 -21366
rect 37562 -21426 37585 -21344
rect 37430 -21686 37585 -21426
rect 36930 -21712 37585 -21686
rect 37649 -21426 37665 -21344
rect 37649 -21712 37822 -21426
rect 8120 -21742 37822 -21712
rect 8120 -22042 8458 -21742
rect 9058 -22042 18090 -21742
rect 18690 -22042 23458 -21742
rect 24058 -22042 33090 -21742
rect 33690 -22042 37822 -21742
rect 8120 -22226 37822 -22042
rect 21852 -22230 21952 -22226
rect 36852 -22230 36952 -22226
<< via4 >>
rect 37972 16812 38702 17542
rect 7318 10012 8118 10812
rect 37966 3702 38712 5450
rect 7348 -5298 8082 -3454
rect 37966 -14302 38700 -12456
rect 7320 -22226 8120 -21426
<< metal5 >>
rect 37936 17542 38736 17578
rect 37936 16812 37972 17542
rect 38702 16812 38736 17542
rect 7320 10836 8120 10896
rect 7294 10812 8142 10836
rect 7294 10012 7318 10812
rect 8118 10012 8142 10812
rect 7294 9988 8142 10012
rect 7320 -3454 8120 9988
rect 7320 -5298 7348 -3454
rect 8082 -5298 8120 -3454
rect 7320 -21402 8120 -5298
rect 37936 5450 38736 16812
rect 37936 3702 37966 5450
rect 38712 3702 38736 5450
rect 37936 -12456 38736 3702
rect 37936 -14302 37966 -12456
rect 38700 -14302 38736 -12456
rect 7296 -21426 8144 -21402
rect 7296 -22226 7320 -21426
rect 8120 -22226 8144 -21426
rect 7296 -22250 8144 -22226
rect 7320 -22262 8120 -22250
rect 37936 -22262 38736 -14302
<< labels >>
flabel metal1 32888 14140 32900 14154 1 FreeSans 480 0 0 0 vsigin
port 3 n
flabel metal2 32196 12456 32208 12470 1 FreeSans 480 0 0 0 ibiasn
port 4 n
flabel metal4 30452 9650 30462 9664 1 FreeSans 480 0 0 0 VSS
port 2 n ground bidirectional
flabel metal4 33486 17114 33506 17132 1 FreeSans 480 0 0 0 VDD
port 1 n power bidirectional
flabel metal1 23198 14118 23210 14134 1 FreeSans 480 0 0 0 vcp
port 5 n
rlabel comment 30552 7328 30552 7328 4 freq_div_0/dfxbp_1
rlabel comment 30552 6240 30552 6240 4 freq_div_0/dfxbp_1
flabel metal1 30232 7863 30285 7892 0 FreeSans 200 0 0 0 freq_div_0/VPWR
rlabel comment 30210 8416 30210 8416 2 freq_div_0/tapvpwrvgnd_1
flabel metal1 30232 7852 30285 7881 0 FreeSans 200 0 0 0 freq_div_0/VPWR
flabel metal1 30232 6775 30285 6804 0 FreeSans 200 0 0 0 freq_div_0/VPWR
rlabel comment 30210 7328 30210 7328 2 freq_div_0/tapvpwrvgnd_1
flabel metal1 30232 6764 30285 6793 0 FreeSans 200 0 0 0 freq_div_0/VPWR
flabel metal1 30232 5687 30285 5716 0 FreeSans 200 0 0 0 freq_div_0/VPWR
rlabel comment 30210 6240 30210 6240 2 freq_div_0/tapvpwrvgnd_1
rlabel comment 36076 6240 36076 6240 8 freq_div_0/tapvpwrvgnd_1
flabel metal1 36001 5687 36054 5716 0 FreeSans 200 180 0 0 freq_div_0/VPWR
flabel metal1 36001 6764 36054 6793 0 FreeSans 200 180 0 0 freq_div_0/VPWR
rlabel comment 36076 7328 36076 7328 8 freq_div_0/tapvpwrvgnd_1
flabel metal1 36001 6775 36054 6804 0 FreeSans 200 180 0 0 freq_div_0/VPWR
flabel metal1 36001 7852 36054 7881 0 FreeSans 200 180 0 0 freq_div_0/VPWR
rlabel comment 36076 8416 36076 8416 8 freq_div_0/tapvpwrvgnd_1
flabel metal1 36001 7863 36054 7892 0 FreeSans 200 180 0 0 freq_div_0/VPWR
flabel metal1 30134 8670 30140 8676 1 FreeSans 480 0 0 0 freq_div_0/vin
flabel metal1 36004 7310 36055 7348 0 FreeSans 200 180 0 0 freq_div_0/VGND
flabel metal1 36004 7308 36055 7346 0 FreeSans 200 180 0 0 freq_div_0/VGND
flabel metal1 36004 6222 36055 6260 0 FreeSans 200 180 0 0 freq_div_0/VGND
flabel metal1 36004 6220 36055 6258 0 FreeSans 200 180 0 0 freq_div_0/VGND
flabel metal1 30231 6220 30282 6258 0 FreeSans 200 0 0 0 freq_div_0/VGND
flabel metal1 30231 6222 30282 6260 0 FreeSans 200 0 0 0 freq_div_0/VGND
flabel metal1 30231 7308 30282 7346 0 FreeSans 200 0 0 0 freq_div_0/VGND
flabel metal1 30231 7310 30282 7348 0 FreeSans 200 0 0 0 freq_div_0/VGND
flabel metal1 30231 8396 30282 8434 0 FreeSans 200 0 0 0 freq_div_0/VGND
flabel metal1 36004 8396 36055 8434 0 FreeSans 200 180 0 0 freq_div_0/VGND
flabel metal4 30446 8180 30450 8184 1 FreeSans 480 0 0 0 freq_div_0/VSS
flabel metal4 33126 8176 33136 8184 1 FreeSans 480 0 0 0 freq_div_0/VDD
flabel metal2 34650 8634 34660 8642 1 FreeSans 480 0 0 0 freq_div_0/vout
flabel metal1 36001 8940 36054 8969 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__tapvpwrvgnd_1_12/VPWR
flabel metal1 36004 8398 36055 8436 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__tapvpwrvgnd_1_12/VGND
rlabel comment 36076 8416 36076 8416 6 freq_div_0/sky130_fd_sc_hd__tapvpwrvgnd_1_12/tapvpwrvgnd_1
flabel metal1 33132 8940 33185 8969 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__tapvpwrvgnd_1_0/VPWR
flabel metal1 33131 8398 33182 8436 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__tapvpwrvgnd_1_0/VGND
rlabel comment 33110 8416 33110 8416 4 freq_div_0/sky130_fd_sc_hd__tapvpwrvgnd_1_0/tapvpwrvgnd_1
flabel locali 32464 8705 32498 8739 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_0/Y
flabel locali 32464 8637 32498 8671 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_0/Y
flabel locali 32372 8637 32406 8671 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_0/A
flabel nwell 32329 8943 32363 8977 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_0/VPB
flabel pwell 32329 8399 32363 8433 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_0/VNB
flabel metal1 32329 8399 32363 8433 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_0/VGND
flabel metal1 32329 8943 32363 8977 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_0/VPWR
rlabel comment 32300 8416 32300 8416 4 freq_div_0/sky130_fd_sc_hd__inv_1_0/inv_1
flabel locali 32973 8569 33007 8603 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_0/Y
flabel locali 32973 8637 33007 8671 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_0/Y
flabel locali 32973 8705 33007 8739 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_0/Y
flabel locali 32605 8637 32639 8671 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_0/A
flabel locali 32697 8637 32731 8671 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_0/A
flabel locali 32789 8637 32823 8671 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_0/A
flabel locali 32881 8637 32915 8671 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_0/A
flabel nwell 32605 8943 32639 8977 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_0/VPB
flabel pwell 32605 8399 32639 8433 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_0/VNB
flabel metal1 32605 8943 32639 8977 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_0/VPWR
flabel metal1 32605 8399 32639 8433 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_0/VGND
rlabel comment 32576 8416 32576 8416 4 freq_div_0/sky130_fd_sc_hd__inv_4_0/inv_4
flabel metal1 30232 8940 30285 8969 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__tapvpwrvgnd_1_1/VPWR
flabel metal1 30231 8398 30282 8436 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__tapvpwrvgnd_1_1/VGND
rlabel comment 30210 8416 30210 8416 4 freq_div_0/sky130_fd_sc_hd__tapvpwrvgnd_1_1/tapvpwrvgnd_1
flabel metal1 30581 8399 30615 8433 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_0/VGND
flabel metal1 30581 8943 30615 8977 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_0/VPWR
flabel locali 32237 8720 32271 8754 0 FreeSans 400 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_0/Q_N
flabel locali 30841 8637 30875 8671 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_0/D
flabel locali 30581 8637 30615 8671 0 FreeSans 400 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_0/CLK
flabel locali 31942 8501 31976 8535 0 FreeSans 400 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_0/Q
flabel pwell 30581 8399 30615 8433 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_0/VNB
flabel pwell 30598 8416 30598 8416 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_0/VNB
flabel nwell 30581 8943 30615 8977 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_0/VPB
flabel nwell 30598 8960 30598 8960 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_0/VPB
rlabel comment 30552 8416 30552 8416 4 freq_div_0/sky130_fd_sc_hd__dfxbp_1_0/dfxbp_1
flabel metal1 36001 7863 36054 7892 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__tapvpwrvgnd_1_11/VPWR
flabel metal1 36004 8396 36055 8434 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__tapvpwrvgnd_1_11/VGND
rlabel comment 36076 8416 36076 8416 8 freq_div_0/sky130_fd_sc_hd__tapvpwrvgnd_1_11/tapvpwrvgnd_1
flabel locali 35162 8093 35196 8127 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_6/Y
flabel locali 35162 8161 35196 8195 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_6/Y
flabel locali 35070 8161 35104 8195 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_6/A
flabel nwell 35027 7855 35061 7889 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_6/VPB
flabel pwell 35027 8399 35061 8433 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_6/VNB
flabel metal1 35027 8399 35061 8433 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_6/VGND
flabel metal1 35027 7855 35061 7889 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_6/VPWR
rlabel comment 34998 8416 34998 8416 2 freq_div_0/sky130_fd_sc_hd__inv_1_6/inv_1
flabel locali 35671 8229 35705 8263 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_6/Y
flabel locali 35671 8161 35705 8195 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_6/Y
flabel locali 35671 8093 35705 8127 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_6/Y
flabel locali 35303 8161 35337 8195 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_6/A
flabel locali 35395 8161 35429 8195 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_6/A
flabel locali 35487 8161 35521 8195 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_6/A
flabel locali 35579 8161 35613 8195 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_6/A
flabel nwell 35303 7855 35337 7889 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_6/VPB
flabel pwell 35303 8399 35337 8433 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_6/VNB
flabel metal1 35303 7855 35337 7889 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_6/VPWR
flabel metal1 35303 8399 35337 8433 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_6/VGND
rlabel comment 35274 8416 35274 8416 2 freq_div_0/sky130_fd_sc_hd__inv_4_6/inv_4
flabel metal1 33279 8399 33313 8433 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_6/VGND
flabel metal1 33279 7855 33313 7889 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_6/VPWR
flabel locali 34935 8078 34969 8112 0 FreeSans 400 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_6/Q_N
flabel locali 33539 8161 33573 8195 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_6/D
flabel locali 33279 8161 33313 8195 0 FreeSans 400 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_6/CLK
flabel locali 34640 8297 34674 8331 0 FreeSans 400 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_6/Q
flabel pwell 33279 8399 33313 8433 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_6/VNB
flabel pwell 33296 8416 33296 8416 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_6/VNB
flabel nwell 33279 7855 33313 7889 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_6/VPB
flabel nwell 33296 7872 33296 7872 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_6/VPB
rlabel comment 33250 8416 33250 8416 2 freq_div_0/sky130_fd_sc_hd__dfxbp_1_6/dfxbp_1
flabel locali 32464 8093 32498 8127 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_1/Y
flabel locali 32464 8161 32498 8195 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_1/Y
flabel locali 32372 8161 32406 8195 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_1/A
flabel nwell 32329 7855 32363 7889 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_1/VPB
flabel pwell 32329 8399 32363 8433 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_1/VNB
flabel metal1 32329 8399 32363 8433 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_1/VGND
flabel metal1 32329 7855 32363 7889 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_1/VPWR
rlabel comment 32300 8416 32300 8416 2 freq_div_0/sky130_fd_sc_hd__inv_1_1/inv_1
flabel locali 32973 8229 33007 8263 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_1/Y
flabel locali 32973 8161 33007 8195 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_1/Y
flabel locali 32973 8093 33007 8127 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_1/Y
flabel locali 32605 8161 32639 8195 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_1/A
flabel locali 32697 8161 32731 8195 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_1/A
flabel locali 32789 8161 32823 8195 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_1/A
flabel locali 32881 8161 32915 8195 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_1/A
flabel nwell 32605 7855 32639 7889 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_1/VPB
flabel pwell 32605 8399 32639 8433 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_1/VNB
flabel metal1 32605 7855 32639 7889 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_1/VPWR
flabel metal1 32605 8399 32639 8433 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_1/VGND
rlabel comment 32576 8416 32576 8416 2 freq_div_0/sky130_fd_sc_hd__inv_4_1/inv_4
flabel metal1 30232 7863 30285 7892 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__tapvpwrvgnd_1_2/VPWR
flabel metal1 30231 8396 30282 8434 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__tapvpwrvgnd_1_2/VGND
rlabel comment 30210 8416 30210 8416 2 freq_div_0/sky130_fd_sc_hd__tapvpwrvgnd_1_2/tapvpwrvgnd_1
flabel metal1 30581 8399 30615 8433 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_1/VGND
flabel metal1 30581 7855 30615 7889 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_1/VPWR
flabel locali 32237 8078 32271 8112 0 FreeSans 400 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_1/Q_N
flabel locali 30841 8161 30875 8195 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_1/D
flabel locali 30581 8161 30615 8195 0 FreeSans 400 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_1/CLK
flabel locali 31942 8297 31976 8331 0 FreeSans 400 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_1/Q
flabel pwell 30581 8399 30615 8433 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_1/VNB
flabel pwell 30598 8416 30598 8416 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_1/VNB
flabel nwell 30581 7855 30615 7889 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_1/VPB
flabel nwell 30598 7872 30598 7872 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_1/VPB
rlabel comment 30552 8416 30552 8416 2 freq_div_0/sky130_fd_sc_hd__dfxbp_1_1/dfxbp_1
flabel metal1 36001 7852 36054 7881 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__tapvpwrvgnd_1_10/VPWR
flabel metal1 36004 7310 36055 7348 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__tapvpwrvgnd_1_10/VGND
rlabel comment 36076 7328 36076 7328 6 freq_div_0/sky130_fd_sc_hd__tapvpwrvgnd_1_10/tapvpwrvgnd_1
flabel locali 35162 7617 35196 7651 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_7/Y
flabel locali 35162 7549 35196 7583 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_7/Y
flabel locali 35070 7549 35104 7583 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_7/A
flabel nwell 35027 7855 35061 7889 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_7/VPB
flabel pwell 35027 7311 35061 7345 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_7/VNB
flabel metal1 35027 7311 35061 7345 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_7/VGND
flabel metal1 35027 7855 35061 7889 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_7/VPWR
rlabel comment 34998 7328 34998 7328 4 freq_div_0/sky130_fd_sc_hd__inv_1_7/inv_1
flabel locali 35671 7481 35705 7515 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_7/Y
flabel locali 35671 7549 35705 7583 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_7/Y
flabel locali 35671 7617 35705 7651 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_7/Y
flabel locali 35303 7549 35337 7583 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_7/A
flabel locali 35395 7549 35429 7583 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_7/A
flabel locali 35487 7549 35521 7583 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_7/A
flabel locali 35579 7549 35613 7583 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_7/A
flabel nwell 35303 7855 35337 7889 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_7/VPB
flabel pwell 35303 7311 35337 7345 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_7/VNB
flabel metal1 35303 7855 35337 7889 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_7/VPWR
flabel metal1 35303 7311 35337 7345 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_7/VGND
rlabel comment 35274 7328 35274 7328 4 freq_div_0/sky130_fd_sc_hd__inv_4_7/inv_4
flabel metal1 33279 7311 33313 7345 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_7/VGND
flabel metal1 33279 7855 33313 7889 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_7/VPWR
flabel locali 34935 7632 34969 7666 0 FreeSans 400 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_7/Q_N
flabel locali 33539 7549 33573 7583 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_7/D
flabel locali 33279 7549 33313 7583 0 FreeSans 400 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_7/CLK
flabel locali 34640 7413 34674 7447 0 FreeSans 400 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_7/Q
flabel pwell 33279 7311 33313 7345 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_7/VNB
flabel pwell 33296 7328 33296 7328 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_7/VNB
flabel nwell 33279 7855 33313 7889 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_7/VPB
flabel nwell 33296 7872 33296 7872 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_7/VPB
rlabel comment 33250 7328 33250 7328 4 freq_div_0/sky130_fd_sc_hd__dfxbp_1_7/dfxbp_1
flabel locali 32464 7617 32498 7651 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_3/Y
flabel locali 32464 7549 32498 7583 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_3/Y
flabel locali 32372 7549 32406 7583 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_3/A
flabel nwell 32329 7855 32363 7889 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_3/VPB
flabel pwell 32329 7311 32363 7345 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_3/VNB
flabel metal1 32329 7311 32363 7345 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_3/VGND
flabel metal1 32329 7855 32363 7889 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_3/VPWR
rlabel comment 32300 7328 32300 7328 4 freq_div_0/sky130_fd_sc_hd__inv_1_3/inv_1
flabel locali 32973 7481 33007 7515 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_3/Y
flabel locali 32973 7549 33007 7583 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_3/Y
flabel locali 32973 7617 33007 7651 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_3/Y
flabel locali 32605 7549 32639 7583 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_3/A
flabel locali 32697 7549 32731 7583 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_3/A
flabel locali 32789 7549 32823 7583 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_3/A
flabel locali 32881 7549 32915 7583 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_3/A
flabel nwell 32605 7855 32639 7889 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_3/VPB
flabel pwell 32605 7311 32639 7345 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_3/VNB
flabel metal1 32605 7855 32639 7889 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_3/VPWR
flabel metal1 32605 7311 32639 7345 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_3/VGND
rlabel comment 32576 7328 32576 7328 4 freq_div_0/sky130_fd_sc_hd__inv_4_3/inv_4
flabel metal1 30232 7852 30285 7881 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__tapvpwrvgnd_1_3/VPWR
flabel metal1 30231 7310 30282 7348 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__tapvpwrvgnd_1_3/VGND
rlabel comment 30210 7328 30210 7328 4 freq_div_0/sky130_fd_sc_hd__tapvpwrvgnd_1_3/tapvpwrvgnd_1
flabel metal1 30581 7311 30615 7345 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_3/VGND
flabel metal1 30581 7855 30615 7889 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_3/VPWR
flabel locali 32237 7632 32271 7666 0 FreeSans 400 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_3/Q_N
flabel locali 30841 7549 30875 7583 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_3/D
flabel locali 30581 7549 30615 7583 0 FreeSans 400 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_3/CLK
flabel locali 31942 7413 31976 7447 0 FreeSans 400 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_3/Q
flabel pwell 30581 7311 30615 7345 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_3/VNB
flabel pwell 30598 7328 30598 7328 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_3/VNB
flabel nwell 30581 7855 30615 7889 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_3/VPB
flabel nwell 30598 7872 30598 7872 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_3/VPB
rlabel comment 30552 7328 30552 7328 4 freq_div_0/sky130_fd_sc_hd__dfxbp_1_3/dfxbp_1
flabel metal1 36001 6775 36054 6804 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__tapvpwrvgnd_1_9/VPWR
flabel metal1 36004 7308 36055 7346 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__tapvpwrvgnd_1_9/VGND
rlabel comment 36076 7328 36076 7328 8 freq_div_0/sky130_fd_sc_hd__tapvpwrvgnd_1_9/tapvpwrvgnd_1
flabel locali 35162 7005 35196 7039 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_8/Y
flabel locali 35162 7073 35196 7107 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_8/Y
flabel locali 35070 7073 35104 7107 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_8/A
flabel nwell 35027 6767 35061 6801 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_8/VPB
flabel pwell 35027 7311 35061 7345 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_8/VNB
flabel metal1 35027 7311 35061 7345 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_8/VGND
flabel metal1 35027 6767 35061 6801 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_8/VPWR
rlabel comment 34998 7328 34998 7328 2 freq_div_0/sky130_fd_sc_hd__inv_1_8/inv_1
flabel locali 35671 7141 35705 7175 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_8/Y
flabel locali 35671 7073 35705 7107 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_8/Y
flabel locali 35671 7005 35705 7039 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_8/Y
flabel locali 35303 7073 35337 7107 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_8/A
flabel locali 35395 7073 35429 7107 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_8/A
flabel locali 35487 7073 35521 7107 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_8/A
flabel locali 35579 7073 35613 7107 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_8/A
flabel nwell 35303 6767 35337 6801 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_8/VPB
flabel pwell 35303 7311 35337 7345 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_8/VNB
flabel metal1 35303 6767 35337 6801 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_8/VPWR
flabel metal1 35303 7311 35337 7345 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_8/VGND
rlabel comment 35274 7328 35274 7328 2 freq_div_0/sky130_fd_sc_hd__inv_4_8/inv_4
flabel metal1 33279 7311 33313 7345 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_8/VGND
flabel metal1 33279 6767 33313 6801 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_8/VPWR
flabel locali 34935 6990 34969 7024 0 FreeSans 400 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_8/Q_N
flabel locali 33539 7073 33573 7107 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_8/D
flabel locali 33279 7073 33313 7107 0 FreeSans 400 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_8/CLK
flabel locali 34640 7209 34674 7243 0 FreeSans 400 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_8/Q
flabel pwell 33279 7311 33313 7345 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_8/VNB
flabel pwell 33296 7328 33296 7328 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_8/VNB
flabel nwell 33279 6767 33313 6801 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_8/VPB
flabel nwell 33296 6784 33296 6784 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_8/VPB
rlabel comment 33250 7328 33250 7328 2 freq_div_0/sky130_fd_sc_hd__dfxbp_1_8/dfxbp_1
flabel locali 32464 7005 32498 7039 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_2/Y
flabel locali 32464 7073 32498 7107 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_2/Y
flabel locali 32372 7073 32406 7107 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_2/A
flabel nwell 32329 6767 32363 6801 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_2/VPB
flabel pwell 32329 7311 32363 7345 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_2/VNB
flabel metal1 32329 7311 32363 7345 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_2/VGND
flabel metal1 32329 6767 32363 6801 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_2/VPWR
rlabel comment 32300 7328 32300 7328 2 freq_div_0/sky130_fd_sc_hd__inv_1_2/inv_1
flabel locali 32973 7141 33007 7175 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_2/Y
flabel locali 32973 7073 33007 7107 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_2/Y
flabel locali 32973 7005 33007 7039 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_2/Y
flabel locali 32605 7073 32639 7107 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_2/A
flabel locali 32697 7073 32731 7107 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_2/A
flabel locali 32789 7073 32823 7107 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_2/A
flabel locali 32881 7073 32915 7107 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_2/A
flabel nwell 32605 6767 32639 6801 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_2/VPB
flabel pwell 32605 7311 32639 7345 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_2/VNB
flabel metal1 32605 6767 32639 6801 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_2/VPWR
flabel metal1 32605 7311 32639 7345 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_2/VGND
rlabel comment 32576 7328 32576 7328 2 freq_div_0/sky130_fd_sc_hd__inv_4_2/inv_4
flabel metal1 30232 6775 30285 6804 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__tapvpwrvgnd_1_4/VPWR
flabel metal1 30231 7308 30282 7346 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__tapvpwrvgnd_1_4/VGND
rlabel comment 30210 7328 30210 7328 2 freq_div_0/sky130_fd_sc_hd__tapvpwrvgnd_1_4/tapvpwrvgnd_1
flabel metal1 30581 7311 30615 7345 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_2/VGND
flabel metal1 30581 6767 30615 6801 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_2/VPWR
flabel locali 32237 6990 32271 7024 0 FreeSans 400 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_2/Q_N
flabel locali 30841 7073 30875 7107 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_2/D
flabel locali 30581 7073 30615 7107 0 FreeSans 400 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_2/CLK
flabel locali 31942 7209 31976 7243 0 FreeSans 400 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_2/Q
flabel pwell 30581 7311 30615 7345 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_2/VNB
flabel pwell 30598 7328 30598 7328 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_2/VNB
flabel nwell 30581 6767 30615 6801 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_2/VPB
flabel nwell 30598 6784 30598 6784 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_2/VPB
rlabel comment 30552 7328 30552 7328 2 freq_div_0/sky130_fd_sc_hd__dfxbp_1_2/dfxbp_1
flabel metal1 36001 6764 36054 6793 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__tapvpwrvgnd_1_8/VPWR
flabel metal1 36004 6222 36055 6260 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__tapvpwrvgnd_1_8/VGND
rlabel comment 36076 6240 36076 6240 6 freq_div_0/sky130_fd_sc_hd__tapvpwrvgnd_1_8/tapvpwrvgnd_1
flabel metal1 36001 5687 36054 5716 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__tapvpwrvgnd_1_7/VPWR
flabel metal1 36004 6220 36055 6258 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__tapvpwrvgnd_1_7/VGND
rlabel comment 36076 6240 36076 6240 8 freq_div_0/sky130_fd_sc_hd__tapvpwrvgnd_1_7/tapvpwrvgnd_1
flabel locali 35162 6529 35196 6563 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_9/Y
flabel locali 35162 6461 35196 6495 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_9/Y
flabel locali 35070 6461 35104 6495 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_9/A
flabel nwell 35027 6767 35061 6801 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_9/VPB
flabel pwell 35027 6223 35061 6257 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_9/VNB
flabel metal1 35027 6223 35061 6257 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_9/VGND
flabel metal1 35027 6767 35061 6801 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_9/VPWR
rlabel comment 34998 6240 34998 6240 4 freq_div_0/sky130_fd_sc_hd__inv_1_9/inv_1
flabel locali 35162 5917 35196 5951 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_10/Y
flabel locali 35162 5985 35196 6019 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_10/Y
flabel locali 35070 5985 35104 6019 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_10/A
flabel nwell 35027 5679 35061 5713 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_10/VPB
flabel pwell 35027 6223 35061 6257 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_10/VNB
flabel metal1 35027 6223 35061 6257 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_10/VGND
flabel metal1 35027 5679 35061 5713 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_10/VPWR
rlabel comment 34998 6240 34998 6240 2 freq_div_0/sky130_fd_sc_hd__inv_1_10/inv_1
flabel locali 35671 6393 35705 6427 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_9/Y
flabel locali 35671 6461 35705 6495 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_9/Y
flabel locali 35671 6529 35705 6563 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_9/Y
flabel locali 35303 6461 35337 6495 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_9/A
flabel locali 35395 6461 35429 6495 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_9/A
flabel locali 35487 6461 35521 6495 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_9/A
flabel locali 35579 6461 35613 6495 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_9/A
flabel nwell 35303 6767 35337 6801 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_9/VPB
flabel pwell 35303 6223 35337 6257 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_9/VNB
flabel metal1 35303 6767 35337 6801 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_9/VPWR
flabel metal1 35303 6223 35337 6257 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_9/VGND
rlabel comment 35274 6240 35274 6240 4 freq_div_0/sky130_fd_sc_hd__inv_4_9/inv_4
flabel locali 35671 6053 35705 6087 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_10/Y
flabel locali 35671 5985 35705 6019 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_10/Y
flabel locali 35671 5917 35705 5951 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_10/Y
flabel locali 35303 5985 35337 6019 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_10/A
flabel locali 35395 5985 35429 6019 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_10/A
flabel locali 35487 5985 35521 6019 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_10/A
flabel locali 35579 5985 35613 6019 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_10/A
flabel nwell 35303 5679 35337 5713 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_10/VPB
flabel pwell 35303 6223 35337 6257 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_10/VNB
flabel metal1 35303 5679 35337 5713 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_10/VPWR
flabel metal1 35303 6223 35337 6257 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_10/VGND
rlabel comment 35274 6240 35274 6240 2 freq_div_0/sky130_fd_sc_hd__inv_4_10/inv_4
flabel metal1 33279 6223 33313 6257 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_9/VGND
flabel metal1 33279 6767 33313 6801 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_9/VPWR
flabel locali 34935 6544 34969 6578 0 FreeSans 400 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_9/Q_N
flabel locali 33539 6461 33573 6495 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_9/D
flabel locali 33279 6461 33313 6495 0 FreeSans 400 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_9/CLK
flabel locali 34640 6325 34674 6359 0 FreeSans 400 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_9/Q
flabel pwell 33279 6223 33313 6257 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_9/VNB
flabel pwell 33296 6240 33296 6240 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_9/VNB
flabel nwell 33279 6767 33313 6801 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_9/VPB
flabel nwell 33296 6784 33296 6784 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_9/VPB
rlabel comment 33250 6240 33250 6240 4 freq_div_0/sky130_fd_sc_hd__dfxbp_1_9/dfxbp_1
flabel metal1 33279 6223 33313 6257 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_10/VGND
flabel metal1 33279 5679 33313 5713 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_10/VPWR
flabel locali 34935 5902 34969 5936 0 FreeSans 400 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_10/Q_N
flabel locali 33539 5985 33573 6019 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_10/D
flabel locali 33279 5985 33313 6019 0 FreeSans 400 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_10/CLK
flabel locali 34640 6121 34674 6155 0 FreeSans 400 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_10/Q
flabel pwell 33279 6223 33313 6257 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_10/VNB
flabel pwell 33296 6240 33296 6240 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_10/VNB
flabel nwell 33279 5679 33313 5713 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_10/VPB
flabel nwell 33296 5696 33296 5696 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_10/VPB
rlabel comment 33250 6240 33250 6240 2 freq_div_0/sky130_fd_sc_hd__dfxbp_1_10/dfxbp_1
flabel locali 32464 6529 32498 6563 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_4/Y
flabel locali 32464 6461 32498 6495 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_4/Y
flabel locali 32372 6461 32406 6495 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_4/A
flabel nwell 32329 6767 32363 6801 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_4/VPB
flabel pwell 32329 6223 32363 6257 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_4/VNB
flabel metal1 32329 6223 32363 6257 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_4/VGND
flabel metal1 32329 6767 32363 6801 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_4/VPWR
rlabel comment 32300 6240 32300 6240 4 freq_div_0/sky130_fd_sc_hd__inv_1_4/inv_1
flabel locali 32464 5917 32498 5951 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_5/Y
flabel locali 32464 5985 32498 6019 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_5/Y
flabel locali 32372 5985 32406 6019 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_5/A
flabel nwell 32329 5679 32363 5713 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_5/VPB
flabel pwell 32329 6223 32363 6257 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_5/VNB
flabel metal1 32329 6223 32363 6257 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_5/VGND
flabel metal1 32329 5679 32363 5713 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_1_5/VPWR
rlabel comment 32300 6240 32300 6240 2 freq_div_0/sky130_fd_sc_hd__inv_1_5/inv_1
flabel locali 32973 6393 33007 6427 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_4/Y
flabel locali 32973 6461 33007 6495 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_4/Y
flabel locali 32973 6529 33007 6563 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_4/Y
flabel locali 32605 6461 32639 6495 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_4/A
flabel locali 32697 6461 32731 6495 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_4/A
flabel locali 32789 6461 32823 6495 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_4/A
flabel locali 32881 6461 32915 6495 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_4/A
flabel nwell 32605 6767 32639 6801 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_4/VPB
flabel pwell 32605 6223 32639 6257 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_4/VNB
flabel metal1 32605 6767 32639 6801 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_4/VPWR
flabel metal1 32605 6223 32639 6257 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_4/VGND
rlabel comment 32576 6240 32576 6240 4 freq_div_0/sky130_fd_sc_hd__inv_4_4/inv_4
flabel locali 32973 6053 33007 6087 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_5/Y
flabel locali 32973 5985 33007 6019 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_5/Y
flabel locali 32973 5917 33007 5951 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_5/Y
flabel locali 32605 5985 32639 6019 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_5/A
flabel locali 32697 5985 32731 6019 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_5/A
flabel locali 32789 5985 32823 6019 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_5/A
flabel locali 32881 5985 32915 6019 0 FreeSans 340 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_5/A
flabel nwell 32605 5679 32639 5713 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_5/VPB
flabel pwell 32605 6223 32639 6257 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_5/VNB
flabel metal1 32605 5679 32639 5713 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_5/VPWR
flabel metal1 32605 6223 32639 6257 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__inv_4_5/VGND
rlabel comment 32576 6240 32576 6240 2 freq_div_0/sky130_fd_sc_hd__inv_4_5/inv_4
flabel metal1 30232 6764 30285 6793 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__tapvpwrvgnd_1_5/VPWR
flabel metal1 30231 6222 30282 6260 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__tapvpwrvgnd_1_5/VGND
rlabel comment 30210 6240 30210 6240 4 freq_div_0/sky130_fd_sc_hd__tapvpwrvgnd_1_5/tapvpwrvgnd_1
flabel metal1 30232 5687 30285 5716 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__tapvpwrvgnd_1_6/VPWR
flabel metal1 30231 6220 30282 6258 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__tapvpwrvgnd_1_6/VGND
rlabel comment 30210 6240 30210 6240 2 freq_div_0/sky130_fd_sc_hd__tapvpwrvgnd_1_6/tapvpwrvgnd_1
flabel metal1 30581 6223 30615 6257 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_4/VGND
flabel metal1 30581 6767 30615 6801 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_4/VPWR
flabel locali 32237 6544 32271 6578 0 FreeSans 400 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_4/Q_N
flabel locali 30841 6461 30875 6495 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_4/D
flabel locali 30581 6461 30615 6495 0 FreeSans 400 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_4/CLK
flabel locali 31942 6325 31976 6359 0 FreeSans 400 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_4/Q
flabel pwell 30581 6223 30615 6257 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_4/VNB
flabel pwell 30598 6240 30598 6240 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_4/VNB
flabel nwell 30581 6767 30615 6801 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_4/VPB
flabel nwell 30598 6784 30598 6784 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_4/VPB
rlabel comment 30552 6240 30552 6240 4 freq_div_0/sky130_fd_sc_hd__dfxbp_1_4/dfxbp_1
flabel metal1 30581 6223 30615 6257 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_5/VGND
flabel metal1 30581 5679 30615 5713 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_5/VPWR
flabel locali 32237 5902 32271 5936 0 FreeSans 400 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_5/Q_N
flabel locali 30841 5985 30875 6019 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_5/D
flabel locali 30581 5985 30615 6019 0 FreeSans 400 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_5/CLK
flabel locali 31942 6121 31976 6155 0 FreeSans 400 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_5/Q
flabel pwell 30581 6223 30615 6257 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_5/VNB
flabel pwell 30598 6240 30598 6240 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_5/VNB
flabel nwell 30581 5679 30615 5713 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_5/VPB
flabel nwell 30598 5696 30598 5696 0 FreeSans 200 0 0 0 freq_div_0/sky130_fd_sc_hd__dfxbp_1_5/VPB
rlabel comment 30552 6240 30552 6240 2 freq_div_0/sky130_fd_sc_hd__dfxbp_1_5/dfxbp_1
flabel metal1 27696 12958 27708 12964 1 FreeSans 480 0 0 0 pfd_cp_lpf_0/vswitchl
flabel metal2 28552 12460 28562 12472 1 FreeSans 480 0 0 0 pfd_cp_lpf_0/ibiasn
flabel metal1 26590 13976 26600 13984 1 FreeSans 480 0 0 0 pfd_cp_lpf_0/vpdiode
flabel metal1 24692 13612 24704 13630 1 FreeSans 480 0 0 0 pfd_cp_lpf_0/vswitchl
flabel metal2 25280 14952 25294 14970 1 FreeSans 480 0 0 0 pfd_cp_lpf_0/vswitchh
flabel metal2 29136 15434 29152 15448 1 FreeSans 480 0 0 0 pfd_cp_lpf_0/vswitchh
flabel metal1 24434 13998 24444 14008 1 FreeSans 480 0 0 0 pfd_cp_lpf_0/vcp
flabel metal1 29632 14146 29636 14150 1 FreeSans 480 0 0 0 pfd_cp_lpf_0/vQB
flabel metal1 29956 14138 29962 14146 1 FreeSans 480 0 0 0 pfd_cp_lpf_0/vQA
flabel metal1 32450 14146 32456 14150 1 FreeSans 480 0 0 0 pfd_cp_lpf_0/vsig_in
flabel metal1 27178 14158 27186 14162 1 FreeSans 480 0 0 0 pfd_cp_lpf_0/vin_div
flabel metal1 29952 14246 29956 14250 1 FreeSans 480 0 0 0 pfd_cp_lpf_0/vRSTN
flabel metal2 29304 13418 29312 13426 1 FreeSans 480 0 0 0 pfd_cp_lpf_0/VQBb
flabel metal2 30028 14692 30036 14700 1 FreeSans 480 0 0 0 pfd_cp_lpf_0/vQAb
flabel metal2 28658 16032 28674 16042 1 FreeSans 480 0 0 0 pfd_cp_lpf_0/vpbias
flabel metal2 28042 11894 28052 11902 1 FreeSans 480 0 0 0 pfd_cp_lpf_0/vpbias
flabel metal4 29358 17044 29370 17060 1 FreeSans 480 0 0 0 pfd_cp_lpf_0/VDD
flabel metal4 28978 11416 29004 11442 1 FreeSans 480 0 0 0 pfd_cp_lpf_0/VSS
flabel metal1 25814 14258 25820 14268 1 FreeSans 480 0 0 0 pfd_cp_lpf_0/vndiode
flabel locali 30006 14203 30040 14237 0 FreeSans 340 0 0 0 pfd_cp_lpf_0/sky130_fd_sc_hd__inv_1_1/Y
flabel locali 30006 14135 30040 14169 0 FreeSans 340 0 0 0 pfd_cp_lpf_0/sky130_fd_sc_hd__inv_1_1/Y
flabel locali 30098 14135 30132 14169 0 FreeSans 340 0 0 0 pfd_cp_lpf_0/sky130_fd_sc_hd__inv_1_1/A
flabel nwell 30141 14441 30175 14475 0 FreeSans 200 0 0 0 pfd_cp_lpf_0/sky130_fd_sc_hd__inv_1_1/VPB
flabel pwell 30141 13897 30175 13931 0 FreeSans 200 0 0 0 pfd_cp_lpf_0/sky130_fd_sc_hd__inv_1_1/VNB
flabel metal1 30141 13897 30175 13931 0 FreeSans 200 0 0 0 pfd_cp_lpf_0/sky130_fd_sc_hd__inv_1_1/VGND
flabel metal1 30141 14441 30175 14475 0 FreeSans 200 0 0 0 pfd_cp_lpf_0/sky130_fd_sc_hd__inv_1_1/VPWR
rlabel comment 30204 13914 30204 13914 6 pfd_cp_lpf_0/sky130_fd_sc_hd__inv_1_1/inv_1
flabel locali 29540 14203 29574 14237 0 FreeSans 340 0 0 0 pfd_cp_lpf_0/sky130_fd_sc_hd__inv_1_0/Y
flabel locali 29540 14135 29574 14169 0 FreeSans 340 0 0 0 pfd_cp_lpf_0/sky130_fd_sc_hd__inv_1_0/Y
flabel locali 29448 14135 29482 14169 0 FreeSans 340 0 0 0 pfd_cp_lpf_0/sky130_fd_sc_hd__inv_1_0/A
flabel nwell 29405 14441 29439 14475 0 FreeSans 200 0 0 0 pfd_cp_lpf_0/sky130_fd_sc_hd__inv_1_0/VPB
flabel pwell 29405 13897 29439 13931 0 FreeSans 200 0 0 0 pfd_cp_lpf_0/sky130_fd_sc_hd__inv_1_0/VNB
flabel metal1 29405 13897 29439 13931 0 FreeSans 200 0 0 0 pfd_cp_lpf_0/sky130_fd_sc_hd__inv_1_0/VGND
flabel metal1 29405 14441 29439 14475 0 FreeSans 200 0 0 0 pfd_cp_lpf_0/sky130_fd_sc_hd__inv_1_0/VPWR
rlabel comment 29376 13914 29376 13914 4 pfd_cp_lpf_0/sky130_fd_sc_hd__inv_1_0/inv_1
flabel locali 30537 14132 30566 14167 0 FreeSans 200 0 0 0 pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_1/Q
flabel locali 30242 14135 30264 14168 0 FreeSans 200 0 0 0 pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_1/Q_N
flabel locali 30805 14067 30839 14101 0 FreeSans 400 0 0 0 pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_1/RESET_B
flabel locali 31981 14203 32015 14237 0 FreeSans 400 0 0 0 pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_1/D
flabel locali 32256 14203 32290 14237 0 FreeSans 400 0 0 0 pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_1/CLK
flabel locali 32256 14135 32290 14169 0 FreeSans 400 0 0 0 pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_1/CLK
flabel locali 30805 14135 30839 14169 0 FreeSans 400 0 0 0 pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_1/RESET_B
flabel metal1 32257 13897 32291 13931 0 FreeSans 200 0 0 0 pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_1/VGND
flabel metal1 32257 14441 32291 14475 0 FreeSans 200 0 0 0 pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_1/VPWR
flabel nwell 32257 14441 32291 14475 0 FreeSans 200 0 0 0 pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_1/VPB
flabel pwell 32257 13897 32291 13931 0 FreeSans 200 0 0 0 pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_1/VNB
rlabel comment 32320 13914 32320 13914 6 pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_1/dfrbp_1
rlabel viali 30805 14067 30839 14101 1 pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_1/RESET_B
rlabel viali 30865 14130 30899 14164 1 pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_1/RESET_B
rlabel locali 30791 14041 30839 14121 1 pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_1/RESET_B
rlabel locali 30791 14121 30899 14195 1 pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_1/RESET_B
rlabel metal1 30793 14061 30851 14070 1 pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_1/RESET_B
rlabel metal1 30853 14107 30911 14170 1 pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_1/RESET_B
rlabel metal1 30793 14098 30911 14107 1 pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_1/RESET_B
rlabel metal1 31441 14098 31571 14107 1 pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_1/RESET_B
rlabel metal1 30793 14070 31571 14098 1 pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_1/RESET_B
rlabel metal1 31441 14061 31571 14070 1 pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_1/RESET_B
flabel locali 29014 14132 29043 14167 0 FreeSans 200 0 0 0 pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_0/Q
flabel locali 29316 14135 29338 14168 0 FreeSans 200 0 0 0 pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_0/Q_N
flabel locali 28741 14067 28775 14101 0 FreeSans 400 0 0 0 pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_0/RESET_B
flabel locali 27565 14203 27599 14237 0 FreeSans 400 0 0 0 pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_0/D
flabel locali 27290 14203 27324 14237 0 FreeSans 400 0 0 0 pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_0/CLK
flabel locali 27290 14135 27324 14169 0 FreeSans 400 0 0 0 pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_0/CLK
flabel locali 28741 14135 28775 14169 0 FreeSans 400 0 0 0 pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_0/RESET_B
flabel metal1 27289 13897 27323 13931 0 FreeSans 200 0 0 0 pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_0/VGND
flabel metal1 27289 14441 27323 14475 0 FreeSans 200 0 0 0 pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_0/VPWR
flabel nwell 27289 14441 27323 14475 0 FreeSans 200 0 0 0 pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_0/VPB
flabel pwell 27289 13897 27323 13931 0 FreeSans 200 0 0 0 pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_0/VNB
rlabel comment 27260 13914 27260 13914 4 pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_0/dfrbp_1
rlabel viali 28741 14067 28775 14101 1 pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_0/RESET_B
rlabel viali 28681 14130 28715 14164 1 pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_0/RESET_B
rlabel locali 28741 14041 28789 14121 1 pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_0/RESET_B
rlabel locali 28681 14121 28789 14195 1 pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_0/RESET_B
rlabel metal1 28729 14061 28787 14070 1 pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_0/RESET_B
rlabel metal1 28669 14107 28727 14170 1 pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_0/RESET_B
rlabel metal1 28669 14098 28787 14107 1 pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_0/RESET_B
rlabel metal1 28009 14098 28139 14107 1 pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_0/RESET_B
rlabel metal1 28009 14070 28787 14098 1 pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_0/RESET_B
rlabel metal1 28009 14061 28139 14070 1 pfd_cp_lpf_0/sky130_fd_sc_hd__dfrbp_1_0/RESET_B
flabel locali 29772 13999 29806 14033 0 FreeSans 250 0 0 0 pfd_cp_lpf_0/sky130_fd_sc_hd__nand2_1_0/Y
flabel locali 29772 14067 29806 14101 0 FreeSans 250 0 0 0 pfd_cp_lpf_0/sky130_fd_sc_hd__nand2_1_0/Y
flabel locali 29772 14135 29806 14169 0 FreeSans 250 0 0 0 pfd_cp_lpf_0/sky130_fd_sc_hd__nand2_1_0/Y
flabel locali 29680 14135 29714 14169 0 FreeSans 250 0 0 0 pfd_cp_lpf_0/sky130_fd_sc_hd__nand2_1_0/B
flabel locali 29864 14135 29898 14169 0 FreeSans 250 0 0 0 pfd_cp_lpf_0/sky130_fd_sc_hd__nand2_1_0/A
flabel nwell 29680 14441 29714 14475 0 FreeSans 200 0 0 0 pfd_cp_lpf_0/sky130_fd_sc_hd__nand2_1_0/VPB
flabel pwell 29680 13897 29714 13931 0 FreeSans 200 0 0 0 pfd_cp_lpf_0/sky130_fd_sc_hd__nand2_1_0/VNB
flabel metal1 29680 13897 29714 13931 0 FreeSans 200 0 0 0 pfd_cp_lpf_0/sky130_fd_sc_hd__nand2_1_0/VGND
flabel metal1 29680 14441 29714 14475 0 FreeSans 200 0 0 0 pfd_cp_lpf_0/sky130_fd_sc_hd__nand2_1_0/VPWR
rlabel comment 29652 13914 29652 13914 4 pfd_cp_lpf_0/sky130_fd_sc_hd__nand2_1_0/nand2_1
flabel metal2 14130 8006 14138 8012 5 FreeSans 480 0 0 0 cs_ring_osc_0/vpbias
flabel metal1 16032 9838 16038 9846 5 FreeSans 480 0 0 0 cs_ring_osc_0/vctrl
flabel metal1 29932 8670 29948 8684 1 FreeSans 480 0 0 0 cs_ring_osc_0/voscbuf
flabel metal1 28632 8728 28648 8740 1 FreeSans 480 0 0 0 cs_ring_osc_0/vosc
flabel metal1 29330 8680 29338 8684 1 FreeSans 480 0 0 0 cs_ring_osc_0/vosc2
flabel metal4 11146 10354 11166 10372 1 FreeSans 480 0 0 0 cs_ring_osc_0/VSS
flabel metal4 10806 4882 10818 4900 1 FreeSans 480 0 0 0 cs_ring_osc_0/VDD
flabel locali 29240 8591 29274 8625 0 FreeSans 340 0 0 0 cs_ring_osc_0/sky130_fd_sc_hd__inv_1_0/Y
flabel locali 29240 8659 29274 8693 0 FreeSans 340 0 0 0 cs_ring_osc_0/sky130_fd_sc_hd__inv_1_0/Y
flabel locali 29148 8659 29182 8693 0 FreeSans 340 0 0 0 cs_ring_osc_0/sky130_fd_sc_hd__inv_1_0/A
flabel nwell 29105 8353 29139 8387 0 FreeSans 200 0 0 0 cs_ring_osc_0/sky130_fd_sc_hd__inv_1_0/VPB
flabel pwell 29105 8897 29139 8931 0 FreeSans 200 0 0 0 cs_ring_osc_0/sky130_fd_sc_hd__inv_1_0/VNB
flabel metal1 29105 8897 29139 8931 0 FreeSans 200 0 0 0 cs_ring_osc_0/sky130_fd_sc_hd__inv_1_0/VGND
flabel metal1 29105 8353 29139 8387 0 FreeSans 200 0 0 0 cs_ring_osc_0/sky130_fd_sc_hd__inv_1_0/VPWR
rlabel comment 29076 8914 29076 8914 2 cs_ring_osc_0/sky130_fd_sc_hd__inv_1_0/inv_1
flabel locali 29749 8727 29783 8761 0 FreeSans 340 0 0 0 cs_ring_osc_0/sky130_fd_sc_hd__inv_4_0/Y
flabel locali 29749 8659 29783 8693 0 FreeSans 340 0 0 0 cs_ring_osc_0/sky130_fd_sc_hd__inv_4_0/Y
flabel locali 29749 8591 29783 8625 0 FreeSans 340 0 0 0 cs_ring_osc_0/sky130_fd_sc_hd__inv_4_0/Y
flabel locali 29381 8659 29415 8693 0 FreeSans 340 0 0 0 cs_ring_osc_0/sky130_fd_sc_hd__inv_4_0/A
flabel locali 29473 8659 29507 8693 0 FreeSans 340 0 0 0 cs_ring_osc_0/sky130_fd_sc_hd__inv_4_0/A
flabel locali 29565 8659 29599 8693 0 FreeSans 340 0 0 0 cs_ring_osc_0/sky130_fd_sc_hd__inv_4_0/A
flabel locali 29657 8659 29691 8693 0 FreeSans 340 0 0 0 cs_ring_osc_0/sky130_fd_sc_hd__inv_4_0/A
flabel nwell 29381 8353 29415 8387 0 FreeSans 200 0 0 0 cs_ring_osc_0/sky130_fd_sc_hd__inv_4_0/VPB
flabel pwell 29381 8897 29415 8931 0 FreeSans 200 0 0 0 cs_ring_osc_0/sky130_fd_sc_hd__inv_4_0/VNB
flabel metal1 29381 8353 29415 8387 0 FreeSans 200 0 0 0 cs_ring_osc_0/sky130_fd_sc_hd__inv_4_0/VPWR
flabel metal1 29381 8897 29415 8931 0 FreeSans 200 0 0 0 cs_ring_osc_0/sky130_fd_sc_hd__inv_4_0/VGND
rlabel comment 29352 8914 29352 8914 2 cs_ring_osc_0/sky130_fd_sc_hd__inv_4_0/inv_4
flabel metal4 26074 -3824 26094 -3804 1 FreeSans 480 0 0 0 cs_ring_osc_0/cs_ring_osc_stage_5/VSS
flabel metal4 25840 4080 25874 4104 1 FreeSans 480 0 0 0 cs_ring_osc_0/cs_ring_osc_stage_5/VDD
flabel metal2 24674 -1570 24688 -1556 1 FreeSans 480 0 0 0 cs_ring_osc_0/cs_ring_osc_stage_5/vin
flabel metal1 24676 -3264 24684 -3254 1 FreeSans 480 0 0 0 cs_ring_osc_0/cs_ring_osc_stage_5/vbiasn
flabel metal2 25146 1152 25156 1158 1 FreeSans 480 0 0 0 cs_ring_osc_0/cs_ring_osc_stage_5/vbiasp
flabel metal2 32500 -1576 32512 -1562 1 FreeSans 480 0 0 0 cs_ring_osc_0/cs_ring_osc_stage_5/voutcs
flabel metal2 32906 -1546 32918 -1536 1 FreeSans 480 0 0 0 cs_ring_osc_0/cs_ring_osc_stage_5/vout
flabel metal1 24240 -2674 24252 -2656 1 FreeSans 480 0 0 0 cs_ring_osc_0/cs_ring_osc_stage_5/csinvn
flabel metal2 24790 554 24800 568 1 FreeSans 480 0 0 0 cs_ring_osc_0/cs_ring_osc_stage_5/csinvp
flabel metal4 11074 -3824 11094 -3804 1 FreeSans 480 0 0 0 cs_ring_osc_0/cs_ring_osc_stage_0/VSS
flabel metal4 10840 4080 10874 4104 1 FreeSans 480 0 0 0 cs_ring_osc_0/cs_ring_osc_stage_0/VDD
flabel metal2 9674 -1570 9688 -1556 1 FreeSans 480 0 0 0 cs_ring_osc_0/cs_ring_osc_stage_0/vin
flabel metal1 9676 -3264 9684 -3254 1 FreeSans 480 0 0 0 cs_ring_osc_0/cs_ring_osc_stage_0/vbiasn
flabel metal2 10146 1152 10156 1158 1 FreeSans 480 0 0 0 cs_ring_osc_0/cs_ring_osc_stage_0/vbiasp
flabel metal2 17500 -1576 17512 -1562 1 FreeSans 480 0 0 0 cs_ring_osc_0/cs_ring_osc_stage_0/voutcs
flabel metal2 17906 -1546 17918 -1536 1 FreeSans 480 0 0 0 cs_ring_osc_0/cs_ring_osc_stage_0/vout
flabel metal1 9240 -2674 9252 -2656 1 FreeSans 480 0 0 0 cs_ring_osc_0/cs_ring_osc_stage_0/csinvn
flabel metal2 9790 554 9800 568 1 FreeSans 480 0 0 0 cs_ring_osc_0/cs_ring_osc_stage_0/csinvp
flabel metal4 35008 -4952 35028 -4932 5 FreeSans 480 0 0 0 cs_ring_osc_0/cs_ring_osc_stage_4/VSS
flabel metal4 35228 -12860 35262 -12836 5 FreeSans 480 0 0 0 cs_ring_osc_0/cs_ring_osc_stage_4/VDD
flabel metal2 36414 -7200 36428 -7186 5 FreeSans 480 0 0 0 cs_ring_osc_0/cs_ring_osc_stage_4/vin
flabel metal1 36418 -5502 36426 -5492 5 FreeSans 480 0 0 0 cs_ring_osc_0/cs_ring_osc_stage_4/vbiasn
flabel metal2 35946 -9914 35956 -9908 5 FreeSans 480 0 0 0 cs_ring_osc_0/cs_ring_osc_stage_4/vbiasp
flabel metal2 28590 -7194 28602 -7180 5 FreeSans 480 0 0 0 cs_ring_osc_0/cs_ring_osc_stage_4/voutcs
flabel metal2 28184 -7220 28196 -7210 5 FreeSans 480 0 0 0 cs_ring_osc_0/cs_ring_osc_stage_4/vout
flabel metal1 36850 -6100 36862 -6082 5 FreeSans 480 0 0 0 cs_ring_osc_0/cs_ring_osc_stage_4/csinvn
flabel metal2 36302 -9324 36312 -9310 5 FreeSans 480 0 0 0 cs_ring_osc_0/cs_ring_osc_stage_4/csinvp
flabel metal4 20008 -4952 20028 -4932 5 FreeSans 480 0 0 0 cs_ring_osc_0/cs_ring_osc_stage_1/VSS
flabel metal4 20228 -12860 20262 -12836 5 FreeSans 480 0 0 0 cs_ring_osc_0/cs_ring_osc_stage_1/VDD
flabel metal2 21414 -7200 21428 -7186 5 FreeSans 480 0 0 0 cs_ring_osc_0/cs_ring_osc_stage_1/vin
flabel metal1 21418 -5502 21426 -5492 5 FreeSans 480 0 0 0 cs_ring_osc_0/cs_ring_osc_stage_1/vbiasn
flabel metal2 20946 -9914 20956 -9908 5 FreeSans 480 0 0 0 cs_ring_osc_0/cs_ring_osc_stage_1/vbiasp
flabel metal2 13590 -7194 13602 -7180 5 FreeSans 480 0 0 0 cs_ring_osc_0/cs_ring_osc_stage_1/voutcs
flabel metal2 13184 -7220 13196 -7210 5 FreeSans 480 0 0 0 cs_ring_osc_0/cs_ring_osc_stage_1/vout
flabel metal1 21850 -6100 21862 -6082 5 FreeSans 480 0 0 0 cs_ring_osc_0/cs_ring_osc_stage_1/csinvn
flabel metal2 21302 -9324 21312 -9310 5 FreeSans 480 0 0 0 cs_ring_osc_0/cs_ring_osc_stage_1/csinvp
flabel metal4 26074 -21824 26094 -21804 1 FreeSans 480 0 0 0 cs_ring_osc_0/cs_ring_osc_stage_3/VSS
flabel metal4 25840 -13920 25874 -13896 1 FreeSans 480 0 0 0 cs_ring_osc_0/cs_ring_osc_stage_3/VDD
flabel metal2 24674 -19570 24688 -19556 1 FreeSans 480 0 0 0 cs_ring_osc_0/cs_ring_osc_stage_3/vin
flabel metal1 24676 -21264 24684 -21254 1 FreeSans 480 0 0 0 cs_ring_osc_0/cs_ring_osc_stage_3/vbiasn
flabel metal2 25146 -16848 25156 -16842 1 FreeSans 480 0 0 0 cs_ring_osc_0/cs_ring_osc_stage_3/vbiasp
flabel metal2 32500 -19576 32512 -19562 1 FreeSans 480 0 0 0 cs_ring_osc_0/cs_ring_osc_stage_3/voutcs
flabel metal2 32906 -19546 32918 -19536 1 FreeSans 480 0 0 0 cs_ring_osc_0/cs_ring_osc_stage_3/vout
flabel metal1 24240 -20674 24252 -20656 1 FreeSans 480 0 0 0 cs_ring_osc_0/cs_ring_osc_stage_3/csinvn
flabel metal2 24790 -17446 24800 -17432 1 FreeSans 480 0 0 0 cs_ring_osc_0/cs_ring_osc_stage_3/csinvp
flabel metal4 11074 -21824 11094 -21804 1 FreeSans 480 0 0 0 cs_ring_osc_0/cs_ring_osc_stage_2/VSS
flabel metal4 10840 -13920 10874 -13896 1 FreeSans 480 0 0 0 cs_ring_osc_0/cs_ring_osc_stage_2/VDD
flabel metal2 9674 -19570 9688 -19556 1 FreeSans 480 0 0 0 cs_ring_osc_0/cs_ring_osc_stage_2/vin
flabel metal1 9676 -21264 9684 -21254 1 FreeSans 480 0 0 0 cs_ring_osc_0/cs_ring_osc_stage_2/vbiasn
flabel metal2 10146 -16848 10156 -16842 1 FreeSans 480 0 0 0 cs_ring_osc_0/cs_ring_osc_stage_2/vbiasp
flabel metal2 17500 -19576 17512 -19562 1 FreeSans 480 0 0 0 cs_ring_osc_0/cs_ring_osc_stage_2/voutcs
flabel metal2 17906 -19546 17918 -19536 1 FreeSans 480 0 0 0 cs_ring_osc_0/cs_ring_osc_stage_2/vout
flabel metal1 9240 -20674 9252 -20656 1 FreeSans 480 0 0 0 cs_ring_osc_0/cs_ring_osc_stage_2/csinvn
flabel metal2 9790 -17446 9800 -17432 1 FreeSans 480 0 0 0 cs_ring_osc_0/cs_ring_osc_stage_2/csinvp
<< end >>
