magic
tech sky130A
magscale 1 2
timestamp 1624477805
<< pwell >>
rect -941 -310 941 310
<< nmos >>
rect -745 -100 -545 100
rect -487 -100 -287 100
rect -229 -100 -29 100
rect 29 -100 229 100
rect 287 -100 487 100
rect 545 -100 745 100
<< ndiff >>
rect -803 88 -745 100
rect -803 -88 -791 88
rect -757 -88 -745 88
rect -803 -100 -745 -88
rect -545 88 -487 100
rect -545 -88 -533 88
rect -499 -88 -487 88
rect -545 -100 -487 -88
rect -287 88 -229 100
rect -287 -88 -275 88
rect -241 -88 -229 88
rect -287 -100 -229 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 229 88 287 100
rect 229 -88 241 88
rect 275 -88 287 88
rect 229 -100 287 -88
rect 487 88 545 100
rect 487 -88 499 88
rect 533 -88 545 88
rect 487 -100 545 -88
rect 745 88 803 100
rect 745 -88 757 88
rect 791 -88 803 88
rect 745 -100 803 -88
<< ndiffc >>
rect -791 -88 -757 88
rect -533 -88 -499 88
rect -275 -88 -241 88
rect -17 -88 17 88
rect 241 -88 275 88
rect 499 -88 533 88
rect 757 -88 791 88
<< psubdiff >>
rect -905 240 -809 274
rect 809 240 905 274
rect -905 178 -871 240
rect 871 178 905 240
rect -905 -240 -871 -178
rect 871 -240 905 -178
rect -905 -274 -809 -240
rect 809 -274 905 -240
<< psubdiffcont >>
rect -809 240 809 274
rect -905 -178 -871 178
rect 871 -178 905 178
rect -809 -274 809 -240
<< poly >>
rect -711 172 -579 188
rect -711 155 -695 172
rect -745 138 -695 155
rect -595 155 -579 172
rect -453 172 -321 188
rect -453 155 -437 172
rect -595 138 -545 155
rect -745 100 -545 138
rect -487 138 -437 155
rect -337 155 -321 172
rect -195 172 -63 188
rect -195 155 -179 172
rect -337 138 -287 155
rect -487 100 -287 138
rect -229 138 -179 155
rect -79 155 -63 172
rect 63 172 195 188
rect 63 155 79 172
rect -79 138 -29 155
rect -229 100 -29 138
rect 29 138 79 155
rect 179 155 195 172
rect 321 172 453 188
rect 321 155 337 172
rect 179 138 229 155
rect 29 100 229 138
rect 287 138 337 155
rect 437 155 453 172
rect 579 172 711 188
rect 579 155 595 172
rect 437 138 487 155
rect 287 100 487 138
rect 545 138 595 155
rect 695 155 711 172
rect 695 138 745 155
rect 545 100 745 138
rect -745 -138 -545 -100
rect -745 -155 -695 -138
rect -711 -172 -695 -155
rect -595 -155 -545 -138
rect -487 -138 -287 -100
rect -487 -155 -437 -138
rect -595 -172 -579 -155
rect -711 -188 -579 -172
rect -453 -172 -437 -155
rect -337 -155 -287 -138
rect -229 -138 -29 -100
rect -229 -155 -179 -138
rect -337 -172 -321 -155
rect -453 -188 -321 -172
rect -195 -172 -179 -155
rect -79 -155 -29 -138
rect 29 -138 229 -100
rect 29 -155 79 -138
rect -79 -172 -63 -155
rect -195 -188 -63 -172
rect 63 -172 79 -155
rect 179 -155 229 -138
rect 287 -138 487 -100
rect 287 -155 337 -138
rect 179 -172 195 -155
rect 63 -188 195 -172
rect 321 -172 337 -155
rect 437 -155 487 -138
rect 545 -138 745 -100
rect 545 -155 595 -138
rect 437 -172 453 -155
rect 321 -188 453 -172
rect 579 -172 595 -155
rect 695 -155 745 -138
rect 695 -172 711 -155
rect 579 -188 711 -172
<< polycont >>
rect -695 138 -595 172
rect -437 138 -337 172
rect -179 138 -79 172
rect 79 138 179 172
rect 337 138 437 172
rect 595 138 695 172
rect -695 -172 -595 -138
rect -437 -172 -337 -138
rect -179 -172 -79 -138
rect 79 -172 179 -138
rect 337 -172 437 -138
rect 595 -172 695 -138
<< locali >>
rect -905 240 -809 274
rect 809 240 905 274
rect -905 178 -871 240
rect 871 178 905 240
rect -711 138 -695 172
rect -595 138 -579 172
rect -453 138 -437 172
rect -337 138 -321 172
rect -195 138 -179 172
rect -79 138 -63 172
rect 63 138 79 172
rect 179 138 195 172
rect 321 138 337 172
rect 437 138 453 172
rect 579 138 595 172
rect 695 138 711 172
rect -791 88 -757 104
rect -791 -104 -757 -88
rect -533 88 -499 104
rect -533 -104 -499 -88
rect -275 88 -241 104
rect -275 -104 -241 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 241 88 275 104
rect 241 -104 275 -88
rect 499 88 533 104
rect 499 -104 533 -88
rect 757 88 791 104
rect 757 -104 791 -88
rect -711 -172 -695 -138
rect -595 -172 -579 -138
rect -453 -172 -437 -138
rect -337 -172 -321 -138
rect -195 -172 -179 -138
rect -79 -172 -63 -138
rect 63 -172 79 -138
rect 179 -172 195 -138
rect 321 -172 337 -138
rect 437 -172 453 -138
rect 579 -172 595 -138
rect 695 -172 711 -138
rect -905 -240 -871 -178
rect 871 -240 905 -178
rect -905 -274 -809 -240
rect 809 -274 905 -240
<< viali >>
rect -687 138 -603 172
rect -429 138 -345 172
rect -171 138 -87 172
rect 87 138 171 172
rect 345 138 429 172
rect 603 138 687 172
rect -791 -88 -757 88
rect -533 -88 -499 88
rect -275 -88 -241 88
rect -17 -88 17 88
rect 241 -88 275 88
rect 499 -88 533 88
rect 757 -88 791 88
rect -687 -172 -603 -138
rect -429 -172 -345 -138
rect -171 -172 -87 -138
rect 87 -172 171 -138
rect 345 -172 429 -138
rect 603 -172 687 -138
<< metal1 >>
rect -699 172 -591 178
rect -699 138 -687 172
rect -603 138 -591 172
rect -699 132 -591 138
rect -441 172 -333 178
rect -441 138 -429 172
rect -345 138 -333 172
rect -441 132 -333 138
rect -183 172 -75 178
rect -183 138 -171 172
rect -87 138 -75 172
rect -183 132 -75 138
rect 75 172 183 178
rect 75 138 87 172
rect 171 138 183 172
rect 75 132 183 138
rect 333 172 441 178
rect 333 138 345 172
rect 429 138 441 172
rect 333 132 441 138
rect 591 172 699 178
rect 591 138 603 172
rect 687 138 699 172
rect 591 132 699 138
rect -797 88 -751 100
rect -797 -88 -791 88
rect -757 -88 -751 88
rect -797 -100 -751 -88
rect -539 88 -493 100
rect -539 -88 -533 88
rect -499 -88 -493 88
rect -539 -100 -493 -88
rect -281 88 -235 100
rect -281 -88 -275 88
rect -241 -88 -235 88
rect -281 -100 -235 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 235 88 281 100
rect 235 -88 241 88
rect 275 -88 281 88
rect 235 -100 281 -88
rect 493 88 539 100
rect 493 -88 499 88
rect 533 -88 539 88
rect 493 -100 539 -88
rect 751 88 797 100
rect 751 -88 757 88
rect 791 -88 797 88
rect 751 -100 797 -88
rect -699 -138 -591 -132
rect -699 -172 -687 -138
rect -603 -172 -591 -138
rect -699 -178 -591 -172
rect -441 -138 -333 -132
rect -441 -172 -429 -138
rect -345 -172 -333 -138
rect -441 -178 -333 -172
rect -183 -138 -75 -132
rect -183 -172 -171 -138
rect -87 -172 -75 -138
rect -183 -178 -75 -172
rect 75 -138 183 -132
rect 75 -172 87 -138
rect 171 -172 183 -138
rect 75 -178 183 -172
rect 333 -138 441 -132
rect 333 -172 345 -138
rect 429 -172 441 -138
rect 333 -178 441 -172
rect 591 -138 699 -132
rect 591 -172 603 -138
rect 687 -172 699 -138
rect 591 -178 699 -172
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -888 -257 888 257
string parameters w 1 l 1 m 1 nf 6 diffcov 100 polycov 60 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
