magic
tech sky130A
magscale 1 2
timestamp 1624252453
<< nwell >>
rect -2000 400 2000 2400
rect -2400 -400 2400 -40
rect -2400 -2400 -2000 -400
rect 2000 -2400 2400 -400
rect -2400 -2800 2400 -2400
<< pwell >>
rect -2400 2400 2400 2800
rect -2400 400 -2000 2400
rect 2000 400 2400 2400
rect -2400 40 2400 400
rect -2000 -2400 2000 -400
<< mvnmos >>
rect -1551 -1900 -1451 -900
rect -1393 -1900 -1293 -900
rect -1235 -1900 -1135 -900
rect -1077 -1900 -977 -900
rect -919 -1900 -819 -900
rect -761 -1900 -661 -900
rect -603 -1900 -503 -900
rect -445 -1900 -345 -900
rect -287 -1900 -187 -900
rect -129 -1900 -29 -900
rect 29 -1900 129 -900
rect 187 -1900 287 -900
rect 345 -1900 445 -900
rect 503 -1900 603 -900
rect 661 -1900 761 -900
rect 819 -1900 919 -900
rect 977 -1900 1077 -900
rect 1135 -1900 1235 -900
rect 1293 -1900 1393 -900
rect 1451 -1900 1551 -900
<< mvpmos >>
rect -1551 900 -1451 1900
rect -1393 900 -1293 1900
rect -1235 900 -1135 1900
rect -1077 900 -977 1900
rect -919 900 -819 1900
rect -761 900 -661 1900
rect -603 900 -503 1900
rect -445 900 -345 1900
rect -287 900 -187 1900
rect -129 900 -29 1900
rect 29 900 129 1900
rect 187 900 287 1900
rect 345 900 445 1900
rect 503 900 603 1900
rect 661 900 761 1900
rect 819 900 919 1900
rect 977 900 1077 1900
rect 1135 900 1235 1900
rect 1293 900 1393 1900
rect 1451 900 1551 1900
<< mvndiff >>
rect -1609 -912 -1551 -900
rect -1609 -1888 -1597 -912
rect -1563 -1888 -1551 -912
rect -1609 -1900 -1551 -1888
rect -1451 -912 -1393 -900
rect -1451 -1888 -1439 -912
rect -1405 -1888 -1393 -912
rect -1451 -1900 -1393 -1888
rect -1293 -912 -1235 -900
rect -1293 -1888 -1281 -912
rect -1247 -1888 -1235 -912
rect -1293 -1900 -1235 -1888
rect -1135 -912 -1077 -900
rect -1135 -1888 -1123 -912
rect -1089 -1888 -1077 -912
rect -1135 -1900 -1077 -1888
rect -977 -912 -919 -900
rect -977 -1888 -965 -912
rect -931 -1888 -919 -912
rect -977 -1900 -919 -1888
rect -819 -912 -761 -900
rect -819 -1888 -807 -912
rect -773 -1888 -761 -912
rect -819 -1900 -761 -1888
rect -661 -912 -603 -900
rect -661 -1888 -649 -912
rect -615 -1888 -603 -912
rect -661 -1900 -603 -1888
rect -503 -912 -445 -900
rect -503 -1888 -491 -912
rect -457 -1888 -445 -912
rect -503 -1900 -445 -1888
rect -345 -912 -287 -900
rect -345 -1888 -333 -912
rect -299 -1888 -287 -912
rect -345 -1900 -287 -1888
rect -187 -912 -129 -900
rect -187 -1888 -175 -912
rect -141 -1888 -129 -912
rect -187 -1900 -129 -1888
rect -29 -912 29 -900
rect -29 -1888 -17 -912
rect 17 -1888 29 -912
rect -29 -1900 29 -1888
rect 129 -912 187 -900
rect 129 -1888 141 -912
rect 175 -1888 187 -912
rect 129 -1900 187 -1888
rect 287 -912 345 -900
rect 287 -1888 299 -912
rect 333 -1888 345 -912
rect 287 -1900 345 -1888
rect 445 -912 503 -900
rect 445 -1888 457 -912
rect 491 -1888 503 -912
rect 445 -1900 503 -1888
rect 603 -912 661 -900
rect 603 -1888 615 -912
rect 649 -1888 661 -912
rect 603 -1900 661 -1888
rect 761 -912 819 -900
rect 761 -1888 773 -912
rect 807 -1888 819 -912
rect 761 -1900 819 -1888
rect 919 -912 977 -900
rect 919 -1888 931 -912
rect 965 -1888 977 -912
rect 919 -1900 977 -1888
rect 1077 -912 1135 -900
rect 1077 -1888 1089 -912
rect 1123 -1888 1135 -912
rect 1077 -1900 1135 -1888
rect 1235 -912 1293 -900
rect 1235 -1888 1247 -912
rect 1281 -1888 1293 -912
rect 1235 -1900 1293 -1888
rect 1393 -912 1451 -900
rect 1393 -1888 1405 -912
rect 1439 -1888 1451 -912
rect 1393 -1900 1451 -1888
rect 1551 -912 1609 -900
rect 1551 -1888 1563 -912
rect 1597 -1888 1609 -912
rect 1551 -1900 1609 -1888
<< mvpdiff >>
rect -1609 1888 -1551 1900
rect -1609 912 -1597 1888
rect -1563 912 -1551 1888
rect -1609 900 -1551 912
rect -1451 1888 -1393 1900
rect -1451 912 -1439 1888
rect -1405 912 -1393 1888
rect -1451 900 -1393 912
rect -1293 1888 -1235 1900
rect -1293 912 -1281 1888
rect -1247 912 -1235 1888
rect -1293 900 -1235 912
rect -1135 1888 -1077 1900
rect -1135 912 -1123 1888
rect -1089 912 -1077 1888
rect -1135 900 -1077 912
rect -977 1888 -919 1900
rect -977 912 -965 1888
rect -931 912 -919 1888
rect -977 900 -919 912
rect -819 1888 -761 1900
rect -819 912 -807 1888
rect -773 912 -761 1888
rect -819 900 -761 912
rect -661 1888 -603 1900
rect -661 912 -649 1888
rect -615 912 -603 1888
rect -661 900 -603 912
rect -503 1888 -445 1900
rect -503 912 -491 1888
rect -457 912 -445 1888
rect -503 900 -445 912
rect -345 1888 -287 1900
rect -345 912 -333 1888
rect -299 912 -287 1888
rect -345 900 -287 912
rect -187 1888 -129 1900
rect -187 912 -175 1888
rect -141 912 -129 1888
rect -187 900 -129 912
rect -29 1888 29 1900
rect -29 912 -17 1888
rect 17 912 29 1888
rect -29 900 29 912
rect 129 1888 187 1900
rect 129 912 141 1888
rect 175 912 187 1888
rect 129 900 187 912
rect 287 1888 345 1900
rect 287 912 299 1888
rect 333 912 345 1888
rect 287 900 345 912
rect 445 1888 503 1900
rect 445 912 457 1888
rect 491 912 503 1888
rect 445 900 503 912
rect 603 1888 661 1900
rect 603 912 615 1888
rect 649 912 661 1888
rect 603 900 661 912
rect 761 1888 819 1900
rect 761 912 773 1888
rect 807 912 819 1888
rect 761 900 819 912
rect 919 1888 977 1900
rect 919 912 931 1888
rect 965 912 977 1888
rect 919 900 977 912
rect 1077 1888 1135 1900
rect 1077 912 1089 1888
rect 1123 912 1135 1888
rect 1077 900 1135 912
rect 1235 1888 1293 1900
rect 1235 912 1247 1888
rect 1281 912 1293 1888
rect 1235 900 1293 912
rect 1393 1888 1451 1900
rect 1393 912 1405 1888
rect 1439 912 1451 1888
rect 1393 900 1451 912
rect 1551 1888 1609 1900
rect 1551 912 1563 1888
rect 1597 912 1609 1888
rect 1551 900 1609 912
<< mvndiffc >>
rect -1597 -1888 -1563 -912
rect -1439 -1888 -1405 -912
rect -1281 -1888 -1247 -912
rect -1123 -1888 -1089 -912
rect -965 -1888 -931 -912
rect -807 -1888 -773 -912
rect -649 -1888 -615 -912
rect -491 -1888 -457 -912
rect -333 -1888 -299 -912
rect -175 -1888 -141 -912
rect -17 -1888 17 -912
rect 141 -1888 175 -912
rect 299 -1888 333 -912
rect 457 -1888 491 -912
rect 615 -1888 649 -912
rect 773 -1888 807 -912
rect 931 -1888 965 -912
rect 1089 -1888 1123 -912
rect 1247 -1888 1281 -912
rect 1405 -1888 1439 -912
rect 1563 -1888 1597 -912
<< mvpdiffc >>
rect -1597 912 -1563 1888
rect -1439 912 -1405 1888
rect -1281 912 -1247 1888
rect -1123 912 -1089 1888
rect -965 912 -931 1888
rect -807 912 -773 1888
rect -649 912 -615 1888
rect -491 912 -457 1888
rect -333 912 -299 1888
rect -175 912 -141 1888
rect -17 912 17 1888
rect 141 912 175 1888
rect 299 912 333 1888
rect 457 912 491 1888
rect 615 912 649 1888
rect 773 912 807 1888
rect 931 912 965 1888
rect 1089 912 1123 1888
rect 1247 912 1281 1888
rect 1405 912 1439 1888
rect 1563 912 1597 1888
<< mvpsubdiff >>
rect -2334 2722 2334 2734
rect -2334 2562 -2100 2722
rect 2100 2562 2334 2722
rect -2334 2550 2334 2562
rect -2334 2500 -2150 2550
rect -2334 340 -2322 2500
rect -2162 340 -2150 2500
rect 2150 2500 2334 2550
rect -2334 290 -2150 340
rect 2150 340 2162 2500
rect 2322 340 2334 2500
rect 2150 290 2334 340
rect -2334 278 2334 290
rect -2334 118 -2100 278
rect 2100 118 2334 278
rect -2334 106 2334 118
rect -1934 -478 1934 -466
rect -1934 -638 -1700 -478
rect 1700 -638 1934 -478
rect -1934 -650 1934 -638
rect -1934 -700 -1750 -650
rect -1934 -2100 -1922 -700
rect -1762 -2100 -1750 -700
rect 1750 -700 1934 -650
rect -1934 -2150 -1750 -2100
rect 1750 -2100 1762 -700
rect 1922 -2100 1934 -700
rect 1750 -2150 1934 -2100
rect -1934 -2162 1934 -2150
rect -1934 -2322 -1700 -2162
rect 1700 -2322 1934 -2162
rect -1934 -2334 1934 -2322
<< mvnsubdiff >>
rect -1934 2322 1934 2334
rect -1934 2162 -1700 2322
rect 1700 2162 1934 2322
rect -1934 2150 1934 2162
rect -1934 2100 -1750 2150
rect -1934 700 -1922 2100
rect -1762 700 -1750 2100
rect 1750 2100 1934 2150
rect -1934 650 -1750 700
rect 1750 700 1762 2100
rect 1922 700 1934 2100
rect 1750 650 1934 700
rect -1934 638 1934 650
rect -1934 478 -1700 638
rect 1700 478 1934 638
rect -1934 466 1934 478
rect -2334 -118 2334 -106
rect -2334 -278 -2100 -118
rect 2100 -278 2334 -118
rect -2334 -290 2334 -278
rect -2334 -340 -2150 -290
rect -2334 -2500 -2322 -340
rect -2162 -2500 -2150 -340
rect 2150 -340 2334 -290
rect -2334 -2550 -2150 -2500
rect 2150 -2500 2162 -340
rect 2322 -2500 2334 -340
rect 2150 -2550 2334 -2500
rect -2334 -2562 2334 -2550
rect -2334 -2722 -2100 -2562
rect 2100 -2722 2334 -2562
rect -2334 -2734 2334 -2722
<< mvpsubdiffcont >>
rect -2100 2562 2100 2722
rect -2322 340 -2162 2500
rect 2162 340 2322 2500
rect -2100 118 2100 278
rect -1700 -638 1700 -478
rect -1922 -2100 -1762 -700
rect 1762 -2100 1922 -700
rect -1700 -2322 1700 -2162
<< mvnsubdiffcont >>
rect -1700 2162 1700 2322
rect -1922 700 -1762 2100
rect 1762 700 1922 2100
rect -1700 478 1700 638
rect -2100 -278 2100 -118
rect -2322 -2500 -2162 -340
rect 2162 -2500 2322 -340
rect -2100 -2722 2100 -2562
<< poly >>
rect -1537 1981 -1465 1997
rect -1537 1964 -1521 1981
rect -1551 1947 -1521 1964
rect -1481 1964 -1465 1981
rect -1379 1981 -1307 1997
rect -1379 1964 -1363 1981
rect -1481 1947 -1451 1964
rect -1551 1900 -1451 1947
rect -1393 1947 -1363 1964
rect -1323 1964 -1307 1981
rect -1221 1981 -1149 1997
rect -1221 1964 -1205 1981
rect -1323 1947 -1293 1964
rect -1393 1900 -1293 1947
rect -1235 1947 -1205 1964
rect -1165 1964 -1149 1981
rect -1063 1981 -991 1997
rect -1063 1964 -1047 1981
rect -1165 1947 -1135 1964
rect -1235 1900 -1135 1947
rect -1077 1947 -1047 1964
rect -1007 1964 -991 1981
rect -905 1981 -833 1997
rect -905 1964 -889 1981
rect -1007 1947 -977 1964
rect -1077 1900 -977 1947
rect -919 1947 -889 1964
rect -849 1964 -833 1981
rect -747 1981 -675 1997
rect -747 1964 -731 1981
rect -849 1947 -819 1964
rect -919 1900 -819 1947
rect -761 1947 -731 1964
rect -691 1964 -675 1981
rect -589 1981 -517 1997
rect -589 1964 -573 1981
rect -691 1947 -661 1964
rect -761 1900 -661 1947
rect -603 1947 -573 1964
rect -533 1964 -517 1981
rect -431 1981 -359 1997
rect -431 1964 -415 1981
rect -533 1947 -503 1964
rect -603 1900 -503 1947
rect -445 1947 -415 1964
rect -375 1964 -359 1981
rect -273 1981 -201 1997
rect -273 1964 -257 1981
rect -375 1947 -345 1964
rect -445 1900 -345 1947
rect -287 1947 -257 1964
rect -217 1964 -201 1981
rect -115 1981 -43 1997
rect -115 1964 -99 1981
rect -217 1947 -187 1964
rect -287 1900 -187 1947
rect -129 1947 -99 1964
rect -59 1964 -43 1981
rect 43 1981 115 1997
rect 43 1964 59 1981
rect -59 1947 -29 1964
rect -129 1900 -29 1947
rect 29 1947 59 1964
rect 99 1964 115 1981
rect 201 1981 273 1997
rect 201 1964 217 1981
rect 99 1947 129 1964
rect 29 1900 129 1947
rect 187 1947 217 1964
rect 257 1964 273 1981
rect 359 1981 431 1997
rect 359 1964 375 1981
rect 257 1947 287 1964
rect 187 1900 287 1947
rect 345 1947 375 1964
rect 415 1964 431 1981
rect 517 1981 589 1997
rect 517 1964 533 1981
rect 415 1947 445 1964
rect 345 1900 445 1947
rect 503 1947 533 1964
rect 573 1964 589 1981
rect 675 1981 747 1997
rect 675 1964 691 1981
rect 573 1947 603 1964
rect 503 1900 603 1947
rect 661 1947 691 1964
rect 731 1964 747 1981
rect 833 1981 905 1997
rect 833 1964 849 1981
rect 731 1947 761 1964
rect 661 1900 761 1947
rect 819 1947 849 1964
rect 889 1964 905 1981
rect 991 1981 1063 1997
rect 991 1964 1007 1981
rect 889 1947 919 1964
rect 819 1900 919 1947
rect 977 1947 1007 1964
rect 1047 1964 1063 1981
rect 1149 1981 1221 1997
rect 1149 1964 1165 1981
rect 1047 1947 1077 1964
rect 977 1900 1077 1947
rect 1135 1947 1165 1964
rect 1205 1964 1221 1981
rect 1307 1981 1379 1997
rect 1307 1964 1323 1981
rect 1205 1947 1235 1964
rect 1135 1900 1235 1947
rect 1293 1947 1323 1964
rect 1363 1964 1379 1981
rect 1465 1981 1537 1997
rect 1465 1964 1481 1981
rect 1363 1947 1393 1964
rect 1293 1900 1393 1947
rect 1451 1947 1481 1964
rect 1521 1964 1537 1981
rect 1521 1947 1551 1964
rect 1451 1900 1551 1947
rect -1551 853 -1451 900
rect -1551 836 -1521 853
rect -1537 819 -1521 836
rect -1481 836 -1451 853
rect -1393 853 -1293 900
rect -1393 836 -1363 853
rect -1481 819 -1465 836
rect -1537 803 -1465 819
rect -1379 819 -1363 836
rect -1323 836 -1293 853
rect -1235 853 -1135 900
rect -1235 836 -1205 853
rect -1323 819 -1307 836
rect -1379 803 -1307 819
rect -1221 819 -1205 836
rect -1165 836 -1135 853
rect -1077 853 -977 900
rect -1077 836 -1047 853
rect -1165 819 -1149 836
rect -1221 803 -1149 819
rect -1063 819 -1047 836
rect -1007 836 -977 853
rect -919 853 -819 900
rect -919 836 -889 853
rect -1007 819 -991 836
rect -1063 803 -991 819
rect -905 819 -889 836
rect -849 836 -819 853
rect -761 853 -661 900
rect -761 836 -731 853
rect -849 819 -833 836
rect -905 803 -833 819
rect -747 819 -731 836
rect -691 836 -661 853
rect -603 853 -503 900
rect -603 836 -573 853
rect -691 819 -675 836
rect -747 803 -675 819
rect -589 819 -573 836
rect -533 836 -503 853
rect -445 853 -345 900
rect -445 836 -415 853
rect -533 819 -517 836
rect -589 803 -517 819
rect -431 819 -415 836
rect -375 836 -345 853
rect -287 853 -187 900
rect -287 836 -257 853
rect -375 819 -359 836
rect -431 803 -359 819
rect -273 819 -257 836
rect -217 836 -187 853
rect -129 853 -29 900
rect -129 836 -99 853
rect -217 819 -201 836
rect -273 803 -201 819
rect -115 819 -99 836
rect -59 836 -29 853
rect 29 853 129 900
rect 29 836 59 853
rect -59 819 -43 836
rect -115 803 -43 819
rect 43 819 59 836
rect 99 836 129 853
rect 187 853 287 900
rect 187 836 217 853
rect 99 819 115 836
rect 43 803 115 819
rect 201 819 217 836
rect 257 836 287 853
rect 345 853 445 900
rect 345 836 375 853
rect 257 819 273 836
rect 201 803 273 819
rect 359 819 375 836
rect 415 836 445 853
rect 503 853 603 900
rect 503 836 533 853
rect 415 819 431 836
rect 359 803 431 819
rect 517 819 533 836
rect 573 836 603 853
rect 661 853 761 900
rect 661 836 691 853
rect 573 819 589 836
rect 517 803 589 819
rect 675 819 691 836
rect 731 836 761 853
rect 819 853 919 900
rect 819 836 849 853
rect 731 819 747 836
rect 675 803 747 819
rect 833 819 849 836
rect 889 836 919 853
rect 977 853 1077 900
rect 977 836 1007 853
rect 889 819 905 836
rect 833 803 905 819
rect 991 819 1007 836
rect 1047 836 1077 853
rect 1135 853 1235 900
rect 1135 836 1165 853
rect 1047 819 1063 836
rect 991 803 1063 819
rect 1149 819 1165 836
rect 1205 836 1235 853
rect 1293 853 1393 900
rect 1293 836 1323 853
rect 1205 819 1221 836
rect 1149 803 1221 819
rect 1307 819 1323 836
rect 1363 836 1393 853
rect 1451 853 1551 900
rect 1451 836 1481 853
rect 1363 819 1379 836
rect 1307 803 1379 819
rect 1465 819 1481 836
rect 1521 836 1551 853
rect 1521 819 1537 836
rect 1465 803 1537 819
rect -1537 -828 -1465 -812
rect -1537 -845 -1521 -828
rect -1551 -862 -1521 -845
rect -1481 -845 -1465 -828
rect -1379 -828 -1307 -812
rect -1379 -845 -1363 -828
rect -1481 -862 -1451 -845
rect -1551 -900 -1451 -862
rect -1393 -862 -1363 -845
rect -1323 -845 -1307 -828
rect -1221 -828 -1149 -812
rect -1221 -845 -1205 -828
rect -1323 -862 -1293 -845
rect -1393 -900 -1293 -862
rect -1235 -862 -1205 -845
rect -1165 -845 -1149 -828
rect -1063 -828 -991 -812
rect -1063 -845 -1047 -828
rect -1165 -862 -1135 -845
rect -1235 -900 -1135 -862
rect -1077 -862 -1047 -845
rect -1007 -845 -991 -828
rect -905 -828 -833 -812
rect -905 -845 -889 -828
rect -1007 -862 -977 -845
rect -1077 -900 -977 -862
rect -919 -862 -889 -845
rect -849 -845 -833 -828
rect -747 -828 -675 -812
rect -747 -845 -731 -828
rect -849 -862 -819 -845
rect -919 -900 -819 -862
rect -761 -862 -731 -845
rect -691 -845 -675 -828
rect -589 -828 -517 -812
rect -589 -845 -573 -828
rect -691 -862 -661 -845
rect -761 -900 -661 -862
rect -603 -862 -573 -845
rect -533 -845 -517 -828
rect -431 -828 -359 -812
rect -431 -845 -415 -828
rect -533 -862 -503 -845
rect -603 -900 -503 -862
rect -445 -862 -415 -845
rect -375 -845 -359 -828
rect -273 -828 -201 -812
rect -273 -845 -257 -828
rect -375 -862 -345 -845
rect -445 -900 -345 -862
rect -287 -862 -257 -845
rect -217 -845 -201 -828
rect -115 -828 -43 -812
rect -115 -845 -99 -828
rect -217 -862 -187 -845
rect -287 -900 -187 -862
rect -129 -862 -99 -845
rect -59 -845 -43 -828
rect 43 -828 115 -812
rect 43 -845 59 -828
rect -59 -862 -29 -845
rect -129 -900 -29 -862
rect 29 -862 59 -845
rect 99 -845 115 -828
rect 201 -828 273 -812
rect 201 -845 217 -828
rect 99 -862 129 -845
rect 29 -900 129 -862
rect 187 -862 217 -845
rect 257 -845 273 -828
rect 359 -828 431 -812
rect 359 -845 375 -828
rect 257 -862 287 -845
rect 187 -900 287 -862
rect 345 -862 375 -845
rect 415 -845 431 -828
rect 517 -828 589 -812
rect 517 -845 533 -828
rect 415 -862 445 -845
rect 345 -900 445 -862
rect 503 -862 533 -845
rect 573 -845 589 -828
rect 675 -828 747 -812
rect 675 -845 691 -828
rect 573 -862 603 -845
rect 503 -900 603 -862
rect 661 -862 691 -845
rect 731 -845 747 -828
rect 833 -828 905 -812
rect 833 -845 849 -828
rect 731 -862 761 -845
rect 661 -900 761 -862
rect 819 -862 849 -845
rect 889 -845 905 -828
rect 991 -828 1063 -812
rect 991 -845 1007 -828
rect 889 -862 919 -845
rect 819 -900 919 -862
rect 977 -862 1007 -845
rect 1047 -845 1063 -828
rect 1149 -828 1221 -812
rect 1149 -845 1165 -828
rect 1047 -862 1077 -845
rect 977 -900 1077 -862
rect 1135 -862 1165 -845
rect 1205 -845 1221 -828
rect 1307 -828 1379 -812
rect 1307 -845 1323 -828
rect 1205 -862 1235 -845
rect 1135 -900 1235 -862
rect 1293 -862 1323 -845
rect 1363 -845 1379 -828
rect 1465 -828 1537 -812
rect 1465 -845 1481 -828
rect 1363 -862 1393 -845
rect 1293 -900 1393 -862
rect 1451 -862 1481 -845
rect 1521 -845 1537 -828
rect 1521 -862 1551 -845
rect 1451 -900 1551 -862
rect -1551 -1938 -1451 -1900
rect -1551 -1955 -1521 -1938
rect -1537 -1972 -1521 -1955
rect -1481 -1955 -1451 -1938
rect -1393 -1938 -1293 -1900
rect -1393 -1955 -1363 -1938
rect -1481 -1972 -1465 -1955
rect -1537 -1988 -1465 -1972
rect -1379 -1972 -1363 -1955
rect -1323 -1955 -1293 -1938
rect -1235 -1938 -1135 -1900
rect -1235 -1955 -1205 -1938
rect -1323 -1972 -1307 -1955
rect -1379 -1988 -1307 -1972
rect -1221 -1972 -1205 -1955
rect -1165 -1955 -1135 -1938
rect -1077 -1938 -977 -1900
rect -1077 -1955 -1047 -1938
rect -1165 -1972 -1149 -1955
rect -1221 -1988 -1149 -1972
rect -1063 -1972 -1047 -1955
rect -1007 -1955 -977 -1938
rect -919 -1938 -819 -1900
rect -919 -1955 -889 -1938
rect -1007 -1972 -991 -1955
rect -1063 -1988 -991 -1972
rect -905 -1972 -889 -1955
rect -849 -1955 -819 -1938
rect -761 -1938 -661 -1900
rect -761 -1955 -731 -1938
rect -849 -1972 -833 -1955
rect -905 -1988 -833 -1972
rect -747 -1972 -731 -1955
rect -691 -1955 -661 -1938
rect -603 -1938 -503 -1900
rect -603 -1955 -573 -1938
rect -691 -1972 -675 -1955
rect -747 -1988 -675 -1972
rect -589 -1972 -573 -1955
rect -533 -1955 -503 -1938
rect -445 -1938 -345 -1900
rect -445 -1955 -415 -1938
rect -533 -1972 -517 -1955
rect -589 -1988 -517 -1972
rect -431 -1972 -415 -1955
rect -375 -1955 -345 -1938
rect -287 -1938 -187 -1900
rect -287 -1955 -257 -1938
rect -375 -1972 -359 -1955
rect -431 -1988 -359 -1972
rect -273 -1972 -257 -1955
rect -217 -1955 -187 -1938
rect -129 -1938 -29 -1900
rect -129 -1955 -99 -1938
rect -217 -1972 -201 -1955
rect -273 -1988 -201 -1972
rect -115 -1972 -99 -1955
rect -59 -1955 -29 -1938
rect 29 -1938 129 -1900
rect 29 -1955 59 -1938
rect -59 -1972 -43 -1955
rect -115 -1988 -43 -1972
rect 43 -1972 59 -1955
rect 99 -1955 129 -1938
rect 187 -1938 287 -1900
rect 187 -1955 217 -1938
rect 99 -1972 115 -1955
rect 43 -1988 115 -1972
rect 201 -1972 217 -1955
rect 257 -1955 287 -1938
rect 345 -1938 445 -1900
rect 345 -1955 375 -1938
rect 257 -1972 273 -1955
rect 201 -1988 273 -1972
rect 359 -1972 375 -1955
rect 415 -1955 445 -1938
rect 503 -1938 603 -1900
rect 503 -1955 533 -1938
rect 415 -1972 431 -1955
rect 359 -1988 431 -1972
rect 517 -1972 533 -1955
rect 573 -1955 603 -1938
rect 661 -1938 761 -1900
rect 661 -1955 691 -1938
rect 573 -1972 589 -1955
rect 517 -1988 589 -1972
rect 675 -1972 691 -1955
rect 731 -1955 761 -1938
rect 819 -1938 919 -1900
rect 819 -1955 849 -1938
rect 731 -1972 747 -1955
rect 675 -1988 747 -1972
rect 833 -1972 849 -1955
rect 889 -1955 919 -1938
rect 977 -1938 1077 -1900
rect 977 -1955 1007 -1938
rect 889 -1972 905 -1955
rect 833 -1988 905 -1972
rect 991 -1972 1007 -1955
rect 1047 -1955 1077 -1938
rect 1135 -1938 1235 -1900
rect 1135 -1955 1165 -1938
rect 1047 -1972 1063 -1955
rect 991 -1988 1063 -1972
rect 1149 -1972 1165 -1955
rect 1205 -1955 1235 -1938
rect 1293 -1938 1393 -1900
rect 1293 -1955 1323 -1938
rect 1205 -1972 1221 -1955
rect 1149 -1988 1221 -1972
rect 1307 -1972 1323 -1955
rect 1363 -1955 1393 -1938
rect 1451 -1938 1551 -1900
rect 1451 -1955 1481 -1938
rect 1363 -1972 1379 -1955
rect 1307 -1988 1379 -1972
rect 1465 -1972 1481 -1955
rect 1521 -1955 1551 -1938
rect 1521 -1972 1537 -1955
rect 1465 -1988 1537 -1972
<< polycont >>
rect -1521 1947 -1481 1981
rect -1363 1947 -1323 1981
rect -1205 1947 -1165 1981
rect -1047 1947 -1007 1981
rect -889 1947 -849 1981
rect -731 1947 -691 1981
rect -573 1947 -533 1981
rect -415 1947 -375 1981
rect -257 1947 -217 1981
rect -99 1947 -59 1981
rect 59 1947 99 1981
rect 217 1947 257 1981
rect 375 1947 415 1981
rect 533 1947 573 1981
rect 691 1947 731 1981
rect 849 1947 889 1981
rect 1007 1947 1047 1981
rect 1165 1947 1205 1981
rect 1323 1947 1363 1981
rect 1481 1947 1521 1981
rect -1521 819 -1481 853
rect -1363 819 -1323 853
rect -1205 819 -1165 853
rect -1047 819 -1007 853
rect -889 819 -849 853
rect -731 819 -691 853
rect -573 819 -533 853
rect -415 819 -375 853
rect -257 819 -217 853
rect -99 819 -59 853
rect 59 819 99 853
rect 217 819 257 853
rect 375 819 415 853
rect 533 819 573 853
rect 691 819 731 853
rect 849 819 889 853
rect 1007 819 1047 853
rect 1165 819 1205 853
rect 1323 819 1363 853
rect 1481 819 1521 853
rect -1521 -862 -1481 -828
rect -1363 -862 -1323 -828
rect -1205 -862 -1165 -828
rect -1047 -862 -1007 -828
rect -889 -862 -849 -828
rect -731 -862 -691 -828
rect -573 -862 -533 -828
rect -415 -862 -375 -828
rect -257 -862 -217 -828
rect -99 -862 -59 -828
rect 59 -862 99 -828
rect 217 -862 257 -828
rect 375 -862 415 -828
rect 533 -862 573 -828
rect 691 -862 731 -828
rect 849 -862 889 -828
rect 1007 -862 1047 -828
rect 1165 -862 1205 -828
rect 1323 -862 1363 -828
rect 1481 -862 1521 -828
rect -1521 -1972 -1481 -1938
rect -1363 -1972 -1323 -1938
rect -1205 -1972 -1165 -1938
rect -1047 -1972 -1007 -1938
rect -889 -1972 -849 -1938
rect -731 -1972 -691 -1938
rect -573 -1972 -533 -1938
rect -415 -1972 -375 -1938
rect -257 -1972 -217 -1938
rect -99 -1972 -59 -1938
rect 59 -1972 99 -1938
rect 217 -1972 257 -1938
rect 375 -1972 415 -1938
rect 533 -1972 573 -1938
rect 691 -1972 731 -1938
rect 849 -1972 889 -1938
rect 1007 -1972 1047 -1938
rect 1165 -1972 1205 -1938
rect 1323 -1972 1363 -1938
rect 1481 -1972 1521 -1938
<< locali >>
rect -2322 2500 -2162 2722
rect 2162 2500 2322 2722
rect -1922 2100 -1762 2322
rect 1762 2100 1922 2322
rect -1597 1888 -1563 1904
rect -1597 896 -1563 912
rect -1439 1888 -1405 1904
rect -1439 896 -1405 912
rect -1281 1888 -1247 1904
rect -1281 896 -1247 912
rect -1123 1888 -1089 1904
rect -1123 896 -1089 912
rect -965 1888 -931 1904
rect -965 896 -931 912
rect -807 1888 -773 1904
rect -807 896 -773 912
rect -649 1888 -615 1904
rect -649 896 -615 912
rect -491 1888 -457 1904
rect -491 896 -457 912
rect -333 1888 -299 1904
rect -333 896 -299 912
rect -175 1888 -141 1904
rect -175 896 -141 912
rect -17 1888 17 1904
rect -17 896 17 912
rect 141 1888 175 1904
rect 141 896 175 912
rect 299 1888 333 1904
rect 299 896 333 912
rect 457 1888 491 1904
rect 457 896 491 912
rect 615 1888 649 1904
rect 615 896 649 912
rect 773 1888 807 1904
rect 773 896 807 912
rect 931 1888 965 1904
rect 931 896 965 912
rect 1089 1888 1123 1904
rect 1089 896 1123 912
rect 1247 1888 1281 1904
rect 1247 896 1281 912
rect 1405 1888 1439 1904
rect 1405 896 1439 912
rect 1563 1888 1597 1904
rect 1563 896 1597 912
rect -1537 819 -1521 853
rect -1481 819 -1465 853
rect -1379 819 -1363 853
rect -1323 819 -1307 853
rect -1221 819 -1205 853
rect -1165 819 -1149 853
rect -1063 819 -1047 853
rect -1007 819 -991 853
rect -905 819 -889 853
rect -849 819 -833 853
rect -747 819 -731 853
rect -691 819 -675 853
rect -589 819 -573 853
rect -533 819 -517 853
rect -431 819 -415 853
rect -375 819 -359 853
rect -273 819 -257 853
rect -217 819 -201 853
rect -115 819 -99 853
rect -59 819 -43 853
rect 43 819 59 853
rect 99 819 115 853
rect 201 819 217 853
rect 257 819 273 853
rect 359 819 375 853
rect 415 819 431 853
rect 517 819 533 853
rect 573 819 589 853
rect 675 819 691 853
rect 731 819 747 853
rect 833 819 849 853
rect 889 819 905 853
rect 991 819 1007 853
rect 1047 819 1063 853
rect 1149 819 1165 853
rect 1205 819 1221 853
rect 1307 819 1323 853
rect 1363 819 1379 853
rect 1465 819 1481 853
rect 1521 819 1537 853
rect -1922 478 -1762 700
rect 1762 478 1922 700
rect -2322 118 -2162 340
rect 2162 118 2322 340
rect -2322 -340 -2162 -118
rect 2162 -340 2322 -118
rect -1922 -700 -1762 -478
rect 1762 -700 1922 -478
rect -1537 -862 -1521 -828
rect -1481 -862 -1465 -828
rect -1379 -862 -1363 -828
rect -1323 -862 -1307 -828
rect -1221 -862 -1205 -828
rect -1165 -862 -1149 -828
rect -1063 -862 -1047 -828
rect -1007 -862 -991 -828
rect -905 -862 -889 -828
rect -849 -862 -833 -828
rect -747 -862 -731 -828
rect -691 -862 -675 -828
rect -589 -862 -573 -828
rect -533 -862 -517 -828
rect -431 -862 -415 -828
rect -375 -862 -359 -828
rect -273 -862 -257 -828
rect -217 -862 -201 -828
rect -115 -862 -99 -828
rect -59 -862 -43 -828
rect 43 -862 59 -828
rect 99 -862 115 -828
rect 201 -862 217 -828
rect 257 -862 273 -828
rect 359 -862 375 -828
rect 415 -862 431 -828
rect 517 -862 533 -828
rect 573 -862 589 -828
rect 675 -862 691 -828
rect 731 -862 747 -828
rect 833 -862 849 -828
rect 889 -862 905 -828
rect 991 -862 1007 -828
rect 1047 -862 1063 -828
rect 1149 -862 1165 -828
rect 1205 -862 1221 -828
rect 1307 -862 1323 -828
rect 1363 -862 1379 -828
rect 1465 -862 1481 -828
rect 1521 -862 1537 -828
rect -1597 -912 -1563 -896
rect -1597 -1904 -1563 -1888
rect -1439 -912 -1405 -896
rect -1439 -1904 -1405 -1888
rect -1281 -912 -1247 -896
rect -1281 -1904 -1247 -1888
rect -1123 -912 -1089 -896
rect -1123 -1904 -1089 -1888
rect -965 -912 -931 -896
rect -965 -1904 -931 -1888
rect -807 -912 -773 -896
rect -807 -1904 -773 -1888
rect -649 -912 -615 -896
rect -649 -1904 -615 -1888
rect -491 -912 -457 -896
rect -491 -1904 -457 -1888
rect -333 -912 -299 -896
rect -333 -1904 -299 -1888
rect -175 -912 -141 -896
rect -175 -1904 -141 -1888
rect -17 -912 17 -896
rect -17 -1904 17 -1888
rect 141 -912 175 -896
rect 141 -1904 175 -1888
rect 299 -912 333 -896
rect 299 -1904 333 -1888
rect 457 -912 491 -896
rect 457 -1904 491 -1888
rect 615 -912 649 -896
rect 615 -1904 649 -1888
rect 773 -912 807 -896
rect 773 -1904 807 -1888
rect 931 -912 965 -896
rect 931 -1904 965 -1888
rect 1089 -912 1123 -896
rect 1089 -1904 1123 -1888
rect 1247 -912 1281 -896
rect 1247 -1904 1281 -1888
rect 1405 -912 1439 -896
rect 1405 -1904 1439 -1888
rect 1563 -912 1597 -896
rect 1563 -1904 1597 -1888
rect -1922 -2322 -1762 -2100
rect 1762 -2322 1922 -2100
rect -2322 -2722 -2162 -2500
rect 2162 -2722 2322 -2500
<< viali >>
rect -2162 2562 -2100 2722
rect -2100 2562 2100 2722
rect 2100 2562 2162 2722
rect -2322 392 -2162 2448
rect -1762 2162 -1700 2322
rect -1700 2162 1700 2322
rect 1700 2162 1762 2322
rect -1922 714 -1762 2086
rect -1603 1947 -1521 1981
rect -1521 1947 -1481 1981
rect -1481 1947 -1363 1981
rect -1363 1947 -1323 1981
rect -1323 1947 -1205 1981
rect -1205 1947 -1165 1981
rect -1165 1947 -1047 1981
rect -1047 1947 -1007 1981
rect -1007 1947 -889 1981
rect -889 1947 -849 1981
rect -849 1947 -731 1981
rect -731 1947 -691 1981
rect -691 1947 -573 1981
rect -573 1947 -533 1981
rect -533 1947 -415 1981
rect -415 1947 -375 1981
rect -375 1947 -257 1981
rect -257 1947 -217 1981
rect -217 1947 -99 1981
rect -99 1947 -59 1981
rect -59 1947 59 1981
rect 59 1947 99 1981
rect 99 1947 217 1981
rect 217 1947 257 1981
rect 257 1947 375 1981
rect 375 1947 415 1981
rect 415 1947 533 1981
rect 533 1947 573 1981
rect 573 1947 691 1981
rect 691 1947 731 1981
rect 731 1947 849 1981
rect 849 1947 889 1981
rect 889 1947 1007 1981
rect 1007 1947 1047 1981
rect 1047 1947 1165 1981
rect 1165 1947 1205 1981
rect 1205 1947 1323 1981
rect 1323 1947 1363 1981
rect 1363 1947 1481 1981
rect 1481 1947 1521 1981
rect 1521 1947 1603 1981
rect -1597 912 -1563 1888
rect -1439 912 -1405 1888
rect -1281 912 -1247 1888
rect -1123 912 -1089 1888
rect -965 912 -931 1888
rect -807 912 -773 1888
rect -649 912 -615 1888
rect -491 912 -457 1888
rect -333 912 -299 1888
rect -175 912 -141 1888
rect -17 912 17 1888
rect 141 912 175 1888
rect 299 912 333 1888
rect 457 912 491 1888
rect 615 912 649 1888
rect 773 912 807 1888
rect 931 912 965 1888
rect 1089 912 1123 1888
rect 1247 912 1281 1888
rect 1405 912 1439 1888
rect 1563 912 1597 1888
rect 1762 714 1922 2086
rect -1762 478 -1700 638
rect -1700 478 1700 638
rect 1700 478 1762 638
rect 2162 392 2322 2448
rect -2162 118 -2100 278
rect -2100 118 2100 278
rect 2100 118 2162 278
rect -2162 -278 -2100 -118
rect -2100 -278 2100 -118
rect 2100 -278 2162 -118
rect -2322 -2448 -2162 -392
rect -1762 -638 -1700 -478
rect -1700 -638 1700 -478
rect 1700 -638 1762 -478
rect -1922 -2086 -1762 -714
rect -1597 -1888 -1563 -912
rect -1439 -1888 -1405 -912
rect -1281 -1888 -1247 -912
rect -1123 -1888 -1089 -912
rect -965 -1888 -931 -912
rect -807 -1888 -773 -912
rect -649 -1888 -615 -912
rect -491 -1888 -457 -912
rect -333 -1888 -299 -912
rect -175 -1888 -141 -912
rect -17 -1888 17 -912
rect 141 -1888 175 -912
rect 299 -1888 333 -912
rect 457 -1888 491 -912
rect 615 -1888 649 -912
rect 773 -1888 807 -912
rect 931 -1888 965 -912
rect 1089 -1888 1123 -912
rect 1247 -1888 1281 -912
rect 1405 -1888 1439 -912
rect 1563 -1888 1597 -912
rect -1603 -1972 -1521 -1938
rect -1521 -1972 -1481 -1938
rect -1481 -1972 -1363 -1938
rect -1363 -1972 -1323 -1938
rect -1323 -1972 -1205 -1938
rect -1205 -1972 -1165 -1938
rect -1165 -1972 -1047 -1938
rect -1047 -1972 -1007 -1938
rect -1007 -1972 -889 -1938
rect -889 -1972 -849 -1938
rect -849 -1972 -731 -1938
rect -731 -1972 -691 -1938
rect -691 -1972 -573 -1938
rect -573 -1972 -533 -1938
rect -533 -1972 -415 -1938
rect -415 -1972 -375 -1938
rect -375 -1972 -257 -1938
rect -257 -1972 -217 -1938
rect -217 -1972 -99 -1938
rect -99 -1972 -59 -1938
rect -59 -1972 59 -1938
rect 59 -1972 99 -1938
rect 99 -1972 217 -1938
rect 217 -1972 257 -1938
rect 257 -1972 375 -1938
rect 375 -1972 415 -1938
rect 415 -1972 533 -1938
rect 533 -1972 573 -1938
rect 573 -1972 691 -1938
rect 691 -1972 731 -1938
rect 731 -1972 849 -1938
rect 849 -1972 889 -1938
rect 889 -1972 1007 -1938
rect 1007 -1972 1047 -1938
rect 1047 -1972 1165 -1938
rect 1165 -1972 1205 -1938
rect 1205 -1972 1323 -1938
rect 1323 -1972 1363 -1938
rect 1363 -1972 1481 -1938
rect 1481 -1972 1521 -1938
rect 1521 -1972 1603 -1938
rect 1762 -2086 1922 -714
rect -1762 -2322 -1700 -2162
rect -1700 -2322 1700 -2162
rect 1700 -2322 1762 -2162
rect 2162 -2448 2322 -392
rect -2162 -2722 -2100 -2562
rect -2100 -2722 2100 -2562
rect 2100 -2722 2162 -2562
<< metal1 >>
rect -2400 3118 2400 3178
rect -2400 2838 -2340 3118
rect 2340 2838 2400 3118
rect -2400 2824 2400 2838
rect -2328 2722 2328 2728
rect -2328 2562 -2162 2722
rect 2162 2562 2328 2722
rect -2328 2460 2328 2562
rect -2328 2448 -2060 2460
rect -2328 392 -2322 2448
rect -2162 392 -2060 2448
rect 2061 2448 2328 2460
rect -2000 2328 2000 2400
rect -2000 2156 -1928 2328
rect 1928 2156 2000 2328
rect -2000 2086 -1756 2156
rect -2000 714 -1922 2086
rect -1762 714 -1756 2086
rect -1603 1987 -1557 2156
rect -1287 1987 -1241 2156
rect -971 1987 -925 2156
rect -655 1987 -609 2156
rect -339 1987 -293 2156
rect -23 1987 23 2156
rect 293 1987 339 2156
rect 609 1987 655 2156
rect 925 1987 971 2156
rect 1241 1987 1287 2156
rect 1557 1987 1603 2156
rect 1756 2086 2000 2156
rect -1615 1981 1615 1987
rect -1615 1947 -1603 1981
rect 1603 1947 1615 1981
rect -1615 1941 1615 1947
rect -1603 1888 -1557 1941
rect -1603 912 -1597 1888
rect -1563 912 -1557 1888
rect -1603 900 -1557 912
rect -1445 1888 -1399 1900
rect -1445 912 -1439 1888
rect -1405 912 -1399 1888
rect -1445 860 -1399 912
rect -1287 1888 -1241 1941
rect -1287 912 -1281 1888
rect -1247 912 -1241 1888
rect -1287 900 -1241 912
rect -1129 1888 -1083 1900
rect -1129 912 -1123 1888
rect -1089 912 -1083 1888
rect -1129 860 -1083 912
rect -971 1888 -925 1941
rect -971 912 -965 1888
rect -931 912 -925 1888
rect -971 900 -925 912
rect -813 1888 -767 1900
rect -813 912 -807 1888
rect -773 912 -767 1888
rect -813 860 -767 912
rect -655 1888 -609 1941
rect -655 912 -649 1888
rect -615 912 -609 1888
rect -655 900 -609 912
rect -497 1888 -451 1900
rect -497 912 -491 1888
rect -457 912 -451 1888
rect -497 860 -451 912
rect -339 1888 -293 1941
rect -339 912 -333 1888
rect -299 912 -293 1888
rect -339 900 -293 912
rect -181 1888 -135 1900
rect -181 912 -175 1888
rect -141 912 -135 1888
rect -181 860 -135 912
rect -23 1888 23 1941
rect -23 912 -17 1888
rect 17 912 23 1888
rect -23 900 23 912
rect 135 1888 181 1900
rect 135 912 141 1888
rect 175 912 181 1888
rect 135 860 181 912
rect 293 1888 339 1941
rect 293 912 299 1888
rect 333 912 339 1888
rect 293 900 339 912
rect 451 1888 497 1900
rect 451 912 457 1888
rect 491 912 497 1888
rect 451 860 497 912
rect 609 1888 655 1941
rect 609 912 615 1888
rect 649 912 655 1888
rect 609 900 655 912
rect 767 1888 813 1900
rect 767 912 773 1888
rect 807 912 813 1888
rect 767 860 813 912
rect 925 1888 971 1941
rect 925 912 931 1888
rect 965 912 971 1888
rect 925 900 971 912
rect 1083 1888 1129 1900
rect 1083 912 1089 1888
rect 1123 912 1129 1888
rect 1083 860 1129 912
rect 1241 1888 1287 1941
rect 1241 912 1247 1888
rect 1281 912 1287 1888
rect 1241 900 1287 912
rect 1399 1888 1445 1900
rect 1399 912 1405 1888
rect 1439 912 1445 1888
rect 1399 860 1445 912
rect 1557 1888 1603 1941
rect 1557 912 1563 1888
rect 1597 912 1603 1888
rect 1557 900 1603 912
rect -2000 644 -1756 714
rect -1455 700 -1445 860
rect -1045 700 1045 860
rect 1445 700 1455 860
rect 1756 714 1762 2086
rect 1922 714 2000 2086
rect 1756 644 2000 714
rect -2000 638 35 644
rect 955 638 2000 644
rect -2000 478 -1762 638
rect 1762 478 2000 638
rect -2000 472 35 478
rect 955 472 2000 478
rect -2000 400 2000 472
rect -2328 340 -2060 392
rect 2061 392 2162 2448
rect 2322 392 2328 2448
rect 2061 340 2328 392
rect -2328 284 2328 340
rect -2328 278 -965 284
rect -45 278 2328 284
rect -2328 118 -2162 278
rect 2162 118 2328 278
rect -2328 112 -965 118
rect -45 112 2328 118
rect -2328 40 2328 112
rect -2360 -112 2360 -40
rect -2360 -118 35 -112
rect 955 -118 2360 -112
rect -2360 -278 -2162 -118
rect 2162 -278 2360 -118
rect -2360 -284 35 -278
rect 955 -284 2360 -278
rect -2360 -340 2360 -284
rect -2360 -392 -2060 -340
rect -2360 -2448 -2322 -392
rect -2162 -2448 -2060 -392
rect 2060 -392 2360 -340
rect -2000 -472 2000 -400
rect -2000 -478 -965 -472
rect -45 -478 2000 -472
rect -2000 -638 -1762 -478
rect 1762 -638 2000 -478
rect -2000 -644 -965 -638
rect -45 -644 2000 -638
rect -2000 -714 -1750 -644
rect -2000 -2086 -1922 -714
rect -1762 -2086 -1750 -714
rect -1455 -860 -1445 -700
rect -1045 -860 1045 -700
rect 1445 -860 1455 -700
rect 1756 -714 2000 -644
rect -1603 -912 -1557 -900
rect -1603 -1888 -1597 -912
rect -1563 -1888 -1557 -912
rect -1603 -1932 -1557 -1888
rect -1445 -912 -1399 -860
rect -1445 -1888 -1439 -912
rect -1405 -1888 -1399 -912
rect -1445 -1900 -1399 -1888
rect -1287 -912 -1241 -900
rect -1287 -1888 -1281 -912
rect -1247 -1888 -1241 -912
rect -1287 -1932 -1241 -1888
rect -1129 -912 -1083 -860
rect -1129 -1888 -1123 -912
rect -1089 -1888 -1083 -912
rect -1129 -1900 -1083 -1888
rect -971 -912 -925 -900
rect -971 -1888 -965 -912
rect -931 -1888 -925 -912
rect -971 -1932 -925 -1888
rect -813 -912 -767 -860
rect -813 -1888 -807 -912
rect -773 -1888 -767 -912
rect -813 -1900 -767 -1888
rect -655 -912 -609 -900
rect -655 -1888 -649 -912
rect -615 -1888 -609 -912
rect -655 -1932 -609 -1888
rect -497 -912 -451 -860
rect -497 -1888 -491 -912
rect -457 -1888 -451 -912
rect -497 -1900 -451 -1888
rect -339 -912 -293 -900
rect -339 -1888 -333 -912
rect -299 -1888 -293 -912
rect -339 -1932 -293 -1888
rect -181 -912 -135 -860
rect -181 -1888 -175 -912
rect -141 -1888 -135 -912
rect -181 -1900 -135 -1888
rect -23 -912 23 -900
rect -23 -1888 -17 -912
rect 17 -1888 23 -912
rect -23 -1932 23 -1888
rect 135 -912 181 -860
rect 135 -1888 141 -912
rect 175 -1888 181 -912
rect 135 -1900 181 -1888
rect 293 -912 339 -900
rect 293 -1888 299 -912
rect 333 -1888 339 -912
rect 293 -1932 339 -1888
rect 451 -912 497 -860
rect 451 -1888 457 -912
rect 491 -1888 497 -912
rect 451 -1900 497 -1888
rect 609 -912 655 -900
rect 609 -1888 615 -912
rect 649 -1888 655 -912
rect 609 -1932 655 -1888
rect 767 -912 813 -860
rect 767 -1888 773 -912
rect 807 -1888 813 -912
rect 767 -1900 813 -1888
rect 925 -912 971 -900
rect 925 -1888 931 -912
rect 965 -1888 971 -912
rect 925 -1932 971 -1888
rect 1083 -912 1129 -860
rect 1083 -1888 1089 -912
rect 1123 -1888 1129 -912
rect 1083 -1900 1129 -1888
rect 1241 -912 1287 -900
rect 1241 -1888 1247 -912
rect 1281 -1888 1287 -912
rect 1241 -1932 1287 -1888
rect 1399 -912 1445 -860
rect 1399 -1888 1405 -912
rect 1439 -1888 1445 -912
rect 1399 -1900 1445 -1888
rect 1557 -912 1603 -900
rect 1557 -1888 1563 -912
rect 1597 -1888 1603 -912
rect 1557 -1932 1603 -1888
rect -1615 -1938 1615 -1932
rect -1615 -1972 -1603 -1938
rect 1603 -1972 1615 -1938
rect -1615 -1978 1615 -1972
rect -2000 -2156 -1750 -2086
rect -1603 -2156 -1557 -1978
rect -1287 -2156 -1241 -1978
rect -971 -2156 -925 -1978
rect -655 -2156 -609 -1978
rect -339 -2156 -293 -1978
rect -23 -2156 23 -1978
rect 293 -2156 339 -1978
rect 609 -2156 655 -1978
rect 925 -2156 971 -1978
rect 1241 -2156 1287 -1978
rect 1557 -2156 1603 -1978
rect 1756 -2086 1762 -714
rect 1922 -2086 2000 -714
rect 1756 -2156 2000 -2086
rect -2000 -2328 -1928 -2156
rect 1928 -2328 2000 -2156
rect -2000 -2400 2000 -2328
rect -2360 -2460 -2060 -2448
rect 2060 -2448 2162 -392
rect 2322 -2448 2360 -392
rect 2060 -2460 2360 -2448
rect -2360 -2562 2360 -2460
rect -2360 -2722 -2162 -2562
rect 2162 -2722 2360 -2562
rect -2360 -2728 2360 -2722
rect -2400 -2838 2400 -2825
rect -2400 -3118 -2340 -2838
rect 2340 -3118 2400 -2838
rect -2400 -3178 2400 -3118
<< via1 >>
rect -2340 2838 2340 3118
rect -1928 2322 1928 2328
rect -1928 2162 -1762 2322
rect -1762 2162 1762 2322
rect 1762 2162 1928 2322
rect -1928 2156 1928 2162
rect -1445 700 -1045 860
rect 1045 700 1445 860
rect 35 638 955 644
rect 35 478 955 638
rect 35 472 955 478
rect -965 278 -45 284
rect -965 118 -45 278
rect -965 112 -45 118
rect 35 -118 955 -112
rect 35 -278 955 -118
rect 35 -284 955 -278
rect -965 -478 -45 -472
rect -965 -638 -45 -478
rect -965 -644 -45 -638
rect -1445 -860 -1045 -700
rect 1045 -860 1445 -700
rect -1928 -2162 1928 -2156
rect -1928 -2322 -1762 -2162
rect -1762 -2322 1762 -2162
rect 1762 -2322 1928 -2162
rect -1928 -2328 1928 -2322
rect -2340 -3118 2340 -2838
<< metal2 >>
rect -2400 3118 2400 3178
rect -2400 2838 -2340 3118
rect 2340 2838 2400 3118
rect -2400 2328 2400 2838
rect -2400 2156 -1928 2328
rect 1928 2156 2400 2328
rect -2400 2150 2400 2156
rect -1928 2146 1928 2150
rect -1445 860 -1045 870
rect -1445 284 -1045 700
rect 1045 860 1445 870
rect 35 644 955 654
rect -2400 -284 -1045 284
rect -1445 -700 -1045 -284
rect -965 284 -45 294
rect -965 -472 -45 112
rect 35 -112 955 472
rect 35 -294 955 -284
rect 1045 284 1445 700
rect 1045 -284 2400 284
rect -965 -654 -45 -644
rect -1445 -870 -1045 -860
rect 1045 -700 1445 -284
rect 1045 -870 1445 -860
rect -1928 -2150 1928 -2146
rect -2400 -2156 2400 -2150
rect -2400 -2328 -1928 -2156
rect 1928 -2328 2400 -2156
rect -2400 -2838 2400 -2328
rect -2400 -3118 -2340 -2838
rect 2340 -3118 2400 -2838
rect -2400 -3178 2400 -3118
<< labels >>
flabel metal2 -2400 -284 -2397 284 3 FreeSans 400 0 0 0 clamp
port 1 e
flabel metal2 -2392 -2814 -2386 -2808 1 FreeSans 480 0 0 0 VSS
port 3 n ground bidirectional
flabel metal2 -2376 2812 -2370 2816 1 FreeSans 480 0 0 0 VDD
port 2 n power bidirectional
<< end >>
