magic
tech sky130A
magscale 1 2
timestamp 1622534145
<< pwell >>
rect -63642 -40598 63642 40598
<< psubdiff >>
rect -63606 40528 -63510 40562
rect 63510 40528 63606 40562
rect -63606 40466 -63572 40528
rect 63572 40466 63606 40528
rect -63606 -40528 -63572 -40466
rect 63572 -40528 63606 -40466
rect -63606 -40562 -63510 -40528
rect 63510 -40562 63606 -40528
<< psubdiffcont >>
rect -63510 40528 63510 40562
rect -63606 -40466 -63572 40466
rect 63572 -40466 63606 40466
rect -63510 -40562 63510 -40528
<< xpolycontact >>
rect -63476 40000 -63406 40432
rect -63476 -40432 -63406 -40000
rect -63158 40000 -63088 40432
rect -63158 -40432 -63088 -40000
rect -62840 40000 -62770 40432
rect -62840 -40432 -62770 -40000
rect -62522 40000 -62452 40432
rect -62522 -40432 -62452 -40000
rect -62204 40000 -62134 40432
rect -62204 -40432 -62134 -40000
rect -61886 40000 -61816 40432
rect -61886 -40432 -61816 -40000
rect -61568 40000 -61498 40432
rect -61568 -40432 -61498 -40000
rect -61250 40000 -61180 40432
rect -61250 -40432 -61180 -40000
rect -60932 40000 -60862 40432
rect -60932 -40432 -60862 -40000
rect -60614 40000 -60544 40432
rect -60614 -40432 -60544 -40000
rect -60296 40000 -60226 40432
rect -60296 -40432 -60226 -40000
rect -59978 40000 -59908 40432
rect -59978 -40432 -59908 -40000
rect -59660 40000 -59590 40432
rect -59660 -40432 -59590 -40000
rect -59342 40000 -59272 40432
rect -59342 -40432 -59272 -40000
rect -59024 40000 -58954 40432
rect -59024 -40432 -58954 -40000
rect -58706 40000 -58636 40432
rect -58706 -40432 -58636 -40000
rect -58388 40000 -58318 40432
rect -58388 -40432 -58318 -40000
rect -58070 40000 -58000 40432
rect -58070 -40432 -58000 -40000
rect -57752 40000 -57682 40432
rect -57752 -40432 -57682 -40000
rect -57434 40000 -57364 40432
rect -57434 -40432 -57364 -40000
rect -57116 40000 -57046 40432
rect -57116 -40432 -57046 -40000
rect -56798 40000 -56728 40432
rect -56798 -40432 -56728 -40000
rect -56480 40000 -56410 40432
rect -56480 -40432 -56410 -40000
rect -56162 40000 -56092 40432
rect -56162 -40432 -56092 -40000
rect -55844 40000 -55774 40432
rect -55844 -40432 -55774 -40000
rect -55526 40000 -55456 40432
rect -55526 -40432 -55456 -40000
rect -55208 40000 -55138 40432
rect -55208 -40432 -55138 -40000
rect -54890 40000 -54820 40432
rect -54890 -40432 -54820 -40000
rect -54572 40000 -54502 40432
rect -54572 -40432 -54502 -40000
rect -54254 40000 -54184 40432
rect -54254 -40432 -54184 -40000
rect -53936 40000 -53866 40432
rect -53936 -40432 -53866 -40000
rect -53618 40000 -53548 40432
rect -53618 -40432 -53548 -40000
rect -53300 40000 -53230 40432
rect -53300 -40432 -53230 -40000
rect -52982 40000 -52912 40432
rect -52982 -40432 -52912 -40000
rect -52664 40000 -52594 40432
rect -52664 -40432 -52594 -40000
rect -52346 40000 -52276 40432
rect -52346 -40432 -52276 -40000
rect -52028 40000 -51958 40432
rect -52028 -40432 -51958 -40000
rect -51710 40000 -51640 40432
rect -51710 -40432 -51640 -40000
rect -51392 40000 -51322 40432
rect -51392 -40432 -51322 -40000
rect -51074 40000 -51004 40432
rect -51074 -40432 -51004 -40000
rect -50756 40000 -50686 40432
rect -50756 -40432 -50686 -40000
rect -50438 40000 -50368 40432
rect -50438 -40432 -50368 -40000
rect -50120 40000 -50050 40432
rect -50120 -40432 -50050 -40000
rect -49802 40000 -49732 40432
rect -49802 -40432 -49732 -40000
rect -49484 40000 -49414 40432
rect -49484 -40432 -49414 -40000
rect -49166 40000 -49096 40432
rect -49166 -40432 -49096 -40000
rect -48848 40000 -48778 40432
rect -48848 -40432 -48778 -40000
rect -48530 40000 -48460 40432
rect -48530 -40432 -48460 -40000
rect -48212 40000 -48142 40432
rect -48212 -40432 -48142 -40000
rect -47894 40000 -47824 40432
rect -47894 -40432 -47824 -40000
rect -47576 40000 -47506 40432
rect -47576 -40432 -47506 -40000
rect -47258 40000 -47188 40432
rect -47258 -40432 -47188 -40000
rect -46940 40000 -46870 40432
rect -46940 -40432 -46870 -40000
rect -46622 40000 -46552 40432
rect -46622 -40432 -46552 -40000
rect -46304 40000 -46234 40432
rect -46304 -40432 -46234 -40000
rect -45986 40000 -45916 40432
rect -45986 -40432 -45916 -40000
rect -45668 40000 -45598 40432
rect -45668 -40432 -45598 -40000
rect -45350 40000 -45280 40432
rect -45350 -40432 -45280 -40000
rect -45032 40000 -44962 40432
rect -45032 -40432 -44962 -40000
rect -44714 40000 -44644 40432
rect -44714 -40432 -44644 -40000
rect -44396 40000 -44326 40432
rect -44396 -40432 -44326 -40000
rect -44078 40000 -44008 40432
rect -44078 -40432 -44008 -40000
rect -43760 40000 -43690 40432
rect -43760 -40432 -43690 -40000
rect -43442 40000 -43372 40432
rect -43442 -40432 -43372 -40000
rect -43124 40000 -43054 40432
rect -43124 -40432 -43054 -40000
rect -42806 40000 -42736 40432
rect -42806 -40432 -42736 -40000
rect -42488 40000 -42418 40432
rect -42488 -40432 -42418 -40000
rect -42170 40000 -42100 40432
rect -42170 -40432 -42100 -40000
rect -41852 40000 -41782 40432
rect -41852 -40432 -41782 -40000
rect -41534 40000 -41464 40432
rect -41534 -40432 -41464 -40000
rect -41216 40000 -41146 40432
rect -41216 -40432 -41146 -40000
rect -40898 40000 -40828 40432
rect -40898 -40432 -40828 -40000
rect -40580 40000 -40510 40432
rect -40580 -40432 -40510 -40000
rect -40262 40000 -40192 40432
rect -40262 -40432 -40192 -40000
rect -39944 40000 -39874 40432
rect -39944 -40432 -39874 -40000
rect -39626 40000 -39556 40432
rect -39626 -40432 -39556 -40000
rect -39308 40000 -39238 40432
rect -39308 -40432 -39238 -40000
rect -38990 40000 -38920 40432
rect -38990 -40432 -38920 -40000
rect -38672 40000 -38602 40432
rect -38672 -40432 -38602 -40000
rect -38354 40000 -38284 40432
rect -38354 -40432 -38284 -40000
rect -38036 40000 -37966 40432
rect -38036 -40432 -37966 -40000
rect -37718 40000 -37648 40432
rect -37718 -40432 -37648 -40000
rect -37400 40000 -37330 40432
rect -37400 -40432 -37330 -40000
rect -37082 40000 -37012 40432
rect -37082 -40432 -37012 -40000
rect -36764 40000 -36694 40432
rect -36764 -40432 -36694 -40000
rect -36446 40000 -36376 40432
rect -36446 -40432 -36376 -40000
rect -36128 40000 -36058 40432
rect -36128 -40432 -36058 -40000
rect -35810 40000 -35740 40432
rect -35810 -40432 -35740 -40000
rect -35492 40000 -35422 40432
rect -35492 -40432 -35422 -40000
rect -35174 40000 -35104 40432
rect -35174 -40432 -35104 -40000
rect -34856 40000 -34786 40432
rect -34856 -40432 -34786 -40000
rect -34538 40000 -34468 40432
rect -34538 -40432 -34468 -40000
rect -34220 40000 -34150 40432
rect -34220 -40432 -34150 -40000
rect -33902 40000 -33832 40432
rect -33902 -40432 -33832 -40000
rect -33584 40000 -33514 40432
rect -33584 -40432 -33514 -40000
rect -33266 40000 -33196 40432
rect -33266 -40432 -33196 -40000
rect -32948 40000 -32878 40432
rect -32948 -40432 -32878 -40000
rect -32630 40000 -32560 40432
rect -32630 -40432 -32560 -40000
rect -32312 40000 -32242 40432
rect -32312 -40432 -32242 -40000
rect -31994 40000 -31924 40432
rect -31994 -40432 -31924 -40000
rect -31676 40000 -31606 40432
rect -31676 -40432 -31606 -40000
rect -31358 40000 -31288 40432
rect -31358 -40432 -31288 -40000
rect -31040 40000 -30970 40432
rect -31040 -40432 -30970 -40000
rect -30722 40000 -30652 40432
rect -30722 -40432 -30652 -40000
rect -30404 40000 -30334 40432
rect -30404 -40432 -30334 -40000
rect -30086 40000 -30016 40432
rect -30086 -40432 -30016 -40000
rect -29768 40000 -29698 40432
rect -29768 -40432 -29698 -40000
rect -29450 40000 -29380 40432
rect -29450 -40432 -29380 -40000
rect -29132 40000 -29062 40432
rect -29132 -40432 -29062 -40000
rect -28814 40000 -28744 40432
rect -28814 -40432 -28744 -40000
rect -28496 40000 -28426 40432
rect -28496 -40432 -28426 -40000
rect -28178 40000 -28108 40432
rect -28178 -40432 -28108 -40000
rect -27860 40000 -27790 40432
rect -27860 -40432 -27790 -40000
rect -27542 40000 -27472 40432
rect -27542 -40432 -27472 -40000
rect -27224 40000 -27154 40432
rect -27224 -40432 -27154 -40000
rect -26906 40000 -26836 40432
rect -26906 -40432 -26836 -40000
rect -26588 40000 -26518 40432
rect -26588 -40432 -26518 -40000
rect -26270 40000 -26200 40432
rect -26270 -40432 -26200 -40000
rect -25952 40000 -25882 40432
rect -25952 -40432 -25882 -40000
rect -25634 40000 -25564 40432
rect -25634 -40432 -25564 -40000
rect -25316 40000 -25246 40432
rect -25316 -40432 -25246 -40000
rect -24998 40000 -24928 40432
rect -24998 -40432 -24928 -40000
rect -24680 40000 -24610 40432
rect -24680 -40432 -24610 -40000
rect -24362 40000 -24292 40432
rect -24362 -40432 -24292 -40000
rect -24044 40000 -23974 40432
rect -24044 -40432 -23974 -40000
rect -23726 40000 -23656 40432
rect -23726 -40432 -23656 -40000
rect -23408 40000 -23338 40432
rect -23408 -40432 -23338 -40000
rect -23090 40000 -23020 40432
rect -23090 -40432 -23020 -40000
rect -22772 40000 -22702 40432
rect -22772 -40432 -22702 -40000
rect -22454 40000 -22384 40432
rect -22454 -40432 -22384 -40000
rect -22136 40000 -22066 40432
rect -22136 -40432 -22066 -40000
rect -21818 40000 -21748 40432
rect -21818 -40432 -21748 -40000
rect -21500 40000 -21430 40432
rect -21500 -40432 -21430 -40000
rect -21182 40000 -21112 40432
rect -21182 -40432 -21112 -40000
rect -20864 40000 -20794 40432
rect -20864 -40432 -20794 -40000
rect -20546 40000 -20476 40432
rect -20546 -40432 -20476 -40000
rect -20228 40000 -20158 40432
rect -20228 -40432 -20158 -40000
rect -19910 40000 -19840 40432
rect -19910 -40432 -19840 -40000
rect -19592 40000 -19522 40432
rect -19592 -40432 -19522 -40000
rect -19274 40000 -19204 40432
rect -19274 -40432 -19204 -40000
rect -18956 40000 -18886 40432
rect -18956 -40432 -18886 -40000
rect -18638 40000 -18568 40432
rect -18638 -40432 -18568 -40000
rect -18320 40000 -18250 40432
rect -18320 -40432 -18250 -40000
rect -18002 40000 -17932 40432
rect -18002 -40432 -17932 -40000
rect -17684 40000 -17614 40432
rect -17684 -40432 -17614 -40000
rect -17366 40000 -17296 40432
rect -17366 -40432 -17296 -40000
rect -17048 40000 -16978 40432
rect -17048 -40432 -16978 -40000
rect -16730 40000 -16660 40432
rect -16730 -40432 -16660 -40000
rect -16412 40000 -16342 40432
rect -16412 -40432 -16342 -40000
rect -16094 40000 -16024 40432
rect -16094 -40432 -16024 -40000
rect -15776 40000 -15706 40432
rect -15776 -40432 -15706 -40000
rect -15458 40000 -15388 40432
rect -15458 -40432 -15388 -40000
rect -15140 40000 -15070 40432
rect -15140 -40432 -15070 -40000
rect -14822 40000 -14752 40432
rect -14822 -40432 -14752 -40000
rect -14504 40000 -14434 40432
rect -14504 -40432 -14434 -40000
rect -14186 40000 -14116 40432
rect -14186 -40432 -14116 -40000
rect -13868 40000 -13798 40432
rect -13868 -40432 -13798 -40000
rect -13550 40000 -13480 40432
rect -13550 -40432 -13480 -40000
rect -13232 40000 -13162 40432
rect -13232 -40432 -13162 -40000
rect -12914 40000 -12844 40432
rect -12914 -40432 -12844 -40000
rect -12596 40000 -12526 40432
rect -12596 -40432 -12526 -40000
rect -12278 40000 -12208 40432
rect -12278 -40432 -12208 -40000
rect -11960 40000 -11890 40432
rect -11960 -40432 -11890 -40000
rect -11642 40000 -11572 40432
rect -11642 -40432 -11572 -40000
rect -11324 40000 -11254 40432
rect -11324 -40432 -11254 -40000
rect -11006 40000 -10936 40432
rect -11006 -40432 -10936 -40000
rect -10688 40000 -10618 40432
rect -10688 -40432 -10618 -40000
rect -10370 40000 -10300 40432
rect -10370 -40432 -10300 -40000
rect -10052 40000 -9982 40432
rect -10052 -40432 -9982 -40000
rect -9734 40000 -9664 40432
rect -9734 -40432 -9664 -40000
rect -9416 40000 -9346 40432
rect -9416 -40432 -9346 -40000
rect -9098 40000 -9028 40432
rect -9098 -40432 -9028 -40000
rect -8780 40000 -8710 40432
rect -8780 -40432 -8710 -40000
rect -8462 40000 -8392 40432
rect -8462 -40432 -8392 -40000
rect -8144 40000 -8074 40432
rect -8144 -40432 -8074 -40000
rect -7826 40000 -7756 40432
rect -7826 -40432 -7756 -40000
rect -7508 40000 -7438 40432
rect -7508 -40432 -7438 -40000
rect -7190 40000 -7120 40432
rect -7190 -40432 -7120 -40000
rect -6872 40000 -6802 40432
rect -6872 -40432 -6802 -40000
rect -6554 40000 -6484 40432
rect -6554 -40432 -6484 -40000
rect -6236 40000 -6166 40432
rect -6236 -40432 -6166 -40000
rect -5918 40000 -5848 40432
rect -5918 -40432 -5848 -40000
rect -5600 40000 -5530 40432
rect -5600 -40432 -5530 -40000
rect -5282 40000 -5212 40432
rect -5282 -40432 -5212 -40000
rect -4964 40000 -4894 40432
rect -4964 -40432 -4894 -40000
rect -4646 40000 -4576 40432
rect -4646 -40432 -4576 -40000
rect -4328 40000 -4258 40432
rect -4328 -40432 -4258 -40000
rect -4010 40000 -3940 40432
rect -4010 -40432 -3940 -40000
rect -3692 40000 -3622 40432
rect -3692 -40432 -3622 -40000
rect -3374 40000 -3304 40432
rect -3374 -40432 -3304 -40000
rect -3056 40000 -2986 40432
rect -3056 -40432 -2986 -40000
rect -2738 40000 -2668 40432
rect -2738 -40432 -2668 -40000
rect -2420 40000 -2350 40432
rect -2420 -40432 -2350 -40000
rect -2102 40000 -2032 40432
rect -2102 -40432 -2032 -40000
rect -1784 40000 -1714 40432
rect -1784 -40432 -1714 -40000
rect -1466 40000 -1396 40432
rect -1466 -40432 -1396 -40000
rect -1148 40000 -1078 40432
rect -1148 -40432 -1078 -40000
rect -830 40000 -760 40432
rect -830 -40432 -760 -40000
rect -512 40000 -442 40432
rect -512 -40432 -442 -40000
rect -194 40000 -124 40432
rect -194 -40432 -124 -40000
rect 124 40000 194 40432
rect 124 -40432 194 -40000
rect 442 40000 512 40432
rect 442 -40432 512 -40000
rect 760 40000 830 40432
rect 760 -40432 830 -40000
rect 1078 40000 1148 40432
rect 1078 -40432 1148 -40000
rect 1396 40000 1466 40432
rect 1396 -40432 1466 -40000
rect 1714 40000 1784 40432
rect 1714 -40432 1784 -40000
rect 2032 40000 2102 40432
rect 2032 -40432 2102 -40000
rect 2350 40000 2420 40432
rect 2350 -40432 2420 -40000
rect 2668 40000 2738 40432
rect 2668 -40432 2738 -40000
rect 2986 40000 3056 40432
rect 2986 -40432 3056 -40000
rect 3304 40000 3374 40432
rect 3304 -40432 3374 -40000
rect 3622 40000 3692 40432
rect 3622 -40432 3692 -40000
rect 3940 40000 4010 40432
rect 3940 -40432 4010 -40000
rect 4258 40000 4328 40432
rect 4258 -40432 4328 -40000
rect 4576 40000 4646 40432
rect 4576 -40432 4646 -40000
rect 4894 40000 4964 40432
rect 4894 -40432 4964 -40000
rect 5212 40000 5282 40432
rect 5212 -40432 5282 -40000
rect 5530 40000 5600 40432
rect 5530 -40432 5600 -40000
rect 5848 40000 5918 40432
rect 5848 -40432 5918 -40000
rect 6166 40000 6236 40432
rect 6166 -40432 6236 -40000
rect 6484 40000 6554 40432
rect 6484 -40432 6554 -40000
rect 6802 40000 6872 40432
rect 6802 -40432 6872 -40000
rect 7120 40000 7190 40432
rect 7120 -40432 7190 -40000
rect 7438 40000 7508 40432
rect 7438 -40432 7508 -40000
rect 7756 40000 7826 40432
rect 7756 -40432 7826 -40000
rect 8074 40000 8144 40432
rect 8074 -40432 8144 -40000
rect 8392 40000 8462 40432
rect 8392 -40432 8462 -40000
rect 8710 40000 8780 40432
rect 8710 -40432 8780 -40000
rect 9028 40000 9098 40432
rect 9028 -40432 9098 -40000
rect 9346 40000 9416 40432
rect 9346 -40432 9416 -40000
rect 9664 40000 9734 40432
rect 9664 -40432 9734 -40000
rect 9982 40000 10052 40432
rect 9982 -40432 10052 -40000
rect 10300 40000 10370 40432
rect 10300 -40432 10370 -40000
rect 10618 40000 10688 40432
rect 10618 -40432 10688 -40000
rect 10936 40000 11006 40432
rect 10936 -40432 11006 -40000
rect 11254 40000 11324 40432
rect 11254 -40432 11324 -40000
rect 11572 40000 11642 40432
rect 11572 -40432 11642 -40000
rect 11890 40000 11960 40432
rect 11890 -40432 11960 -40000
rect 12208 40000 12278 40432
rect 12208 -40432 12278 -40000
rect 12526 40000 12596 40432
rect 12526 -40432 12596 -40000
rect 12844 40000 12914 40432
rect 12844 -40432 12914 -40000
rect 13162 40000 13232 40432
rect 13162 -40432 13232 -40000
rect 13480 40000 13550 40432
rect 13480 -40432 13550 -40000
rect 13798 40000 13868 40432
rect 13798 -40432 13868 -40000
rect 14116 40000 14186 40432
rect 14116 -40432 14186 -40000
rect 14434 40000 14504 40432
rect 14434 -40432 14504 -40000
rect 14752 40000 14822 40432
rect 14752 -40432 14822 -40000
rect 15070 40000 15140 40432
rect 15070 -40432 15140 -40000
rect 15388 40000 15458 40432
rect 15388 -40432 15458 -40000
rect 15706 40000 15776 40432
rect 15706 -40432 15776 -40000
rect 16024 40000 16094 40432
rect 16024 -40432 16094 -40000
rect 16342 40000 16412 40432
rect 16342 -40432 16412 -40000
rect 16660 40000 16730 40432
rect 16660 -40432 16730 -40000
rect 16978 40000 17048 40432
rect 16978 -40432 17048 -40000
rect 17296 40000 17366 40432
rect 17296 -40432 17366 -40000
rect 17614 40000 17684 40432
rect 17614 -40432 17684 -40000
rect 17932 40000 18002 40432
rect 17932 -40432 18002 -40000
rect 18250 40000 18320 40432
rect 18250 -40432 18320 -40000
rect 18568 40000 18638 40432
rect 18568 -40432 18638 -40000
rect 18886 40000 18956 40432
rect 18886 -40432 18956 -40000
rect 19204 40000 19274 40432
rect 19204 -40432 19274 -40000
rect 19522 40000 19592 40432
rect 19522 -40432 19592 -40000
rect 19840 40000 19910 40432
rect 19840 -40432 19910 -40000
rect 20158 40000 20228 40432
rect 20158 -40432 20228 -40000
rect 20476 40000 20546 40432
rect 20476 -40432 20546 -40000
rect 20794 40000 20864 40432
rect 20794 -40432 20864 -40000
rect 21112 40000 21182 40432
rect 21112 -40432 21182 -40000
rect 21430 40000 21500 40432
rect 21430 -40432 21500 -40000
rect 21748 40000 21818 40432
rect 21748 -40432 21818 -40000
rect 22066 40000 22136 40432
rect 22066 -40432 22136 -40000
rect 22384 40000 22454 40432
rect 22384 -40432 22454 -40000
rect 22702 40000 22772 40432
rect 22702 -40432 22772 -40000
rect 23020 40000 23090 40432
rect 23020 -40432 23090 -40000
rect 23338 40000 23408 40432
rect 23338 -40432 23408 -40000
rect 23656 40000 23726 40432
rect 23656 -40432 23726 -40000
rect 23974 40000 24044 40432
rect 23974 -40432 24044 -40000
rect 24292 40000 24362 40432
rect 24292 -40432 24362 -40000
rect 24610 40000 24680 40432
rect 24610 -40432 24680 -40000
rect 24928 40000 24998 40432
rect 24928 -40432 24998 -40000
rect 25246 40000 25316 40432
rect 25246 -40432 25316 -40000
rect 25564 40000 25634 40432
rect 25564 -40432 25634 -40000
rect 25882 40000 25952 40432
rect 25882 -40432 25952 -40000
rect 26200 40000 26270 40432
rect 26200 -40432 26270 -40000
rect 26518 40000 26588 40432
rect 26518 -40432 26588 -40000
rect 26836 40000 26906 40432
rect 26836 -40432 26906 -40000
rect 27154 40000 27224 40432
rect 27154 -40432 27224 -40000
rect 27472 40000 27542 40432
rect 27472 -40432 27542 -40000
rect 27790 40000 27860 40432
rect 27790 -40432 27860 -40000
rect 28108 40000 28178 40432
rect 28108 -40432 28178 -40000
rect 28426 40000 28496 40432
rect 28426 -40432 28496 -40000
rect 28744 40000 28814 40432
rect 28744 -40432 28814 -40000
rect 29062 40000 29132 40432
rect 29062 -40432 29132 -40000
rect 29380 40000 29450 40432
rect 29380 -40432 29450 -40000
rect 29698 40000 29768 40432
rect 29698 -40432 29768 -40000
rect 30016 40000 30086 40432
rect 30016 -40432 30086 -40000
rect 30334 40000 30404 40432
rect 30334 -40432 30404 -40000
rect 30652 40000 30722 40432
rect 30652 -40432 30722 -40000
rect 30970 40000 31040 40432
rect 30970 -40432 31040 -40000
rect 31288 40000 31358 40432
rect 31288 -40432 31358 -40000
rect 31606 40000 31676 40432
rect 31606 -40432 31676 -40000
rect 31924 40000 31994 40432
rect 31924 -40432 31994 -40000
rect 32242 40000 32312 40432
rect 32242 -40432 32312 -40000
rect 32560 40000 32630 40432
rect 32560 -40432 32630 -40000
rect 32878 40000 32948 40432
rect 32878 -40432 32948 -40000
rect 33196 40000 33266 40432
rect 33196 -40432 33266 -40000
rect 33514 40000 33584 40432
rect 33514 -40432 33584 -40000
rect 33832 40000 33902 40432
rect 33832 -40432 33902 -40000
rect 34150 40000 34220 40432
rect 34150 -40432 34220 -40000
rect 34468 40000 34538 40432
rect 34468 -40432 34538 -40000
rect 34786 40000 34856 40432
rect 34786 -40432 34856 -40000
rect 35104 40000 35174 40432
rect 35104 -40432 35174 -40000
rect 35422 40000 35492 40432
rect 35422 -40432 35492 -40000
rect 35740 40000 35810 40432
rect 35740 -40432 35810 -40000
rect 36058 40000 36128 40432
rect 36058 -40432 36128 -40000
rect 36376 40000 36446 40432
rect 36376 -40432 36446 -40000
rect 36694 40000 36764 40432
rect 36694 -40432 36764 -40000
rect 37012 40000 37082 40432
rect 37012 -40432 37082 -40000
rect 37330 40000 37400 40432
rect 37330 -40432 37400 -40000
rect 37648 40000 37718 40432
rect 37648 -40432 37718 -40000
rect 37966 40000 38036 40432
rect 37966 -40432 38036 -40000
rect 38284 40000 38354 40432
rect 38284 -40432 38354 -40000
rect 38602 40000 38672 40432
rect 38602 -40432 38672 -40000
rect 38920 40000 38990 40432
rect 38920 -40432 38990 -40000
rect 39238 40000 39308 40432
rect 39238 -40432 39308 -40000
rect 39556 40000 39626 40432
rect 39556 -40432 39626 -40000
rect 39874 40000 39944 40432
rect 39874 -40432 39944 -40000
rect 40192 40000 40262 40432
rect 40192 -40432 40262 -40000
rect 40510 40000 40580 40432
rect 40510 -40432 40580 -40000
rect 40828 40000 40898 40432
rect 40828 -40432 40898 -40000
rect 41146 40000 41216 40432
rect 41146 -40432 41216 -40000
rect 41464 40000 41534 40432
rect 41464 -40432 41534 -40000
rect 41782 40000 41852 40432
rect 41782 -40432 41852 -40000
rect 42100 40000 42170 40432
rect 42100 -40432 42170 -40000
rect 42418 40000 42488 40432
rect 42418 -40432 42488 -40000
rect 42736 40000 42806 40432
rect 42736 -40432 42806 -40000
rect 43054 40000 43124 40432
rect 43054 -40432 43124 -40000
rect 43372 40000 43442 40432
rect 43372 -40432 43442 -40000
rect 43690 40000 43760 40432
rect 43690 -40432 43760 -40000
rect 44008 40000 44078 40432
rect 44008 -40432 44078 -40000
rect 44326 40000 44396 40432
rect 44326 -40432 44396 -40000
rect 44644 40000 44714 40432
rect 44644 -40432 44714 -40000
rect 44962 40000 45032 40432
rect 44962 -40432 45032 -40000
rect 45280 40000 45350 40432
rect 45280 -40432 45350 -40000
rect 45598 40000 45668 40432
rect 45598 -40432 45668 -40000
rect 45916 40000 45986 40432
rect 45916 -40432 45986 -40000
rect 46234 40000 46304 40432
rect 46234 -40432 46304 -40000
rect 46552 40000 46622 40432
rect 46552 -40432 46622 -40000
rect 46870 40000 46940 40432
rect 46870 -40432 46940 -40000
rect 47188 40000 47258 40432
rect 47188 -40432 47258 -40000
rect 47506 40000 47576 40432
rect 47506 -40432 47576 -40000
rect 47824 40000 47894 40432
rect 47824 -40432 47894 -40000
rect 48142 40000 48212 40432
rect 48142 -40432 48212 -40000
rect 48460 40000 48530 40432
rect 48460 -40432 48530 -40000
rect 48778 40000 48848 40432
rect 48778 -40432 48848 -40000
rect 49096 40000 49166 40432
rect 49096 -40432 49166 -40000
rect 49414 40000 49484 40432
rect 49414 -40432 49484 -40000
rect 49732 40000 49802 40432
rect 49732 -40432 49802 -40000
rect 50050 40000 50120 40432
rect 50050 -40432 50120 -40000
rect 50368 40000 50438 40432
rect 50368 -40432 50438 -40000
rect 50686 40000 50756 40432
rect 50686 -40432 50756 -40000
rect 51004 40000 51074 40432
rect 51004 -40432 51074 -40000
rect 51322 40000 51392 40432
rect 51322 -40432 51392 -40000
rect 51640 40000 51710 40432
rect 51640 -40432 51710 -40000
rect 51958 40000 52028 40432
rect 51958 -40432 52028 -40000
rect 52276 40000 52346 40432
rect 52276 -40432 52346 -40000
rect 52594 40000 52664 40432
rect 52594 -40432 52664 -40000
rect 52912 40000 52982 40432
rect 52912 -40432 52982 -40000
rect 53230 40000 53300 40432
rect 53230 -40432 53300 -40000
rect 53548 40000 53618 40432
rect 53548 -40432 53618 -40000
rect 53866 40000 53936 40432
rect 53866 -40432 53936 -40000
rect 54184 40000 54254 40432
rect 54184 -40432 54254 -40000
rect 54502 40000 54572 40432
rect 54502 -40432 54572 -40000
rect 54820 40000 54890 40432
rect 54820 -40432 54890 -40000
rect 55138 40000 55208 40432
rect 55138 -40432 55208 -40000
rect 55456 40000 55526 40432
rect 55456 -40432 55526 -40000
rect 55774 40000 55844 40432
rect 55774 -40432 55844 -40000
rect 56092 40000 56162 40432
rect 56092 -40432 56162 -40000
rect 56410 40000 56480 40432
rect 56410 -40432 56480 -40000
rect 56728 40000 56798 40432
rect 56728 -40432 56798 -40000
rect 57046 40000 57116 40432
rect 57046 -40432 57116 -40000
rect 57364 40000 57434 40432
rect 57364 -40432 57434 -40000
rect 57682 40000 57752 40432
rect 57682 -40432 57752 -40000
rect 58000 40000 58070 40432
rect 58000 -40432 58070 -40000
rect 58318 40000 58388 40432
rect 58318 -40432 58388 -40000
rect 58636 40000 58706 40432
rect 58636 -40432 58706 -40000
rect 58954 40000 59024 40432
rect 58954 -40432 59024 -40000
rect 59272 40000 59342 40432
rect 59272 -40432 59342 -40000
rect 59590 40000 59660 40432
rect 59590 -40432 59660 -40000
rect 59908 40000 59978 40432
rect 59908 -40432 59978 -40000
rect 60226 40000 60296 40432
rect 60226 -40432 60296 -40000
rect 60544 40000 60614 40432
rect 60544 -40432 60614 -40000
rect 60862 40000 60932 40432
rect 60862 -40432 60932 -40000
rect 61180 40000 61250 40432
rect 61180 -40432 61250 -40000
rect 61498 40000 61568 40432
rect 61498 -40432 61568 -40000
rect 61816 40000 61886 40432
rect 61816 -40432 61886 -40000
rect 62134 40000 62204 40432
rect 62134 -40432 62204 -40000
rect 62452 40000 62522 40432
rect 62452 -40432 62522 -40000
rect 62770 40000 62840 40432
rect 62770 -40432 62840 -40000
rect 63088 40000 63158 40432
rect 63088 -40432 63158 -40000
rect 63406 40000 63476 40432
rect 63406 -40432 63476 -40000
<< xpolyres >>
rect -63476 -40000 -63406 40000
rect -63158 -40000 -63088 40000
rect -62840 -40000 -62770 40000
rect -62522 -40000 -62452 40000
rect -62204 -40000 -62134 40000
rect -61886 -40000 -61816 40000
rect -61568 -40000 -61498 40000
rect -61250 -40000 -61180 40000
rect -60932 -40000 -60862 40000
rect -60614 -40000 -60544 40000
rect -60296 -40000 -60226 40000
rect -59978 -40000 -59908 40000
rect -59660 -40000 -59590 40000
rect -59342 -40000 -59272 40000
rect -59024 -40000 -58954 40000
rect -58706 -40000 -58636 40000
rect -58388 -40000 -58318 40000
rect -58070 -40000 -58000 40000
rect -57752 -40000 -57682 40000
rect -57434 -40000 -57364 40000
rect -57116 -40000 -57046 40000
rect -56798 -40000 -56728 40000
rect -56480 -40000 -56410 40000
rect -56162 -40000 -56092 40000
rect -55844 -40000 -55774 40000
rect -55526 -40000 -55456 40000
rect -55208 -40000 -55138 40000
rect -54890 -40000 -54820 40000
rect -54572 -40000 -54502 40000
rect -54254 -40000 -54184 40000
rect -53936 -40000 -53866 40000
rect -53618 -40000 -53548 40000
rect -53300 -40000 -53230 40000
rect -52982 -40000 -52912 40000
rect -52664 -40000 -52594 40000
rect -52346 -40000 -52276 40000
rect -52028 -40000 -51958 40000
rect -51710 -40000 -51640 40000
rect -51392 -40000 -51322 40000
rect -51074 -40000 -51004 40000
rect -50756 -40000 -50686 40000
rect -50438 -40000 -50368 40000
rect -50120 -40000 -50050 40000
rect -49802 -40000 -49732 40000
rect -49484 -40000 -49414 40000
rect -49166 -40000 -49096 40000
rect -48848 -40000 -48778 40000
rect -48530 -40000 -48460 40000
rect -48212 -40000 -48142 40000
rect -47894 -40000 -47824 40000
rect -47576 -40000 -47506 40000
rect -47258 -40000 -47188 40000
rect -46940 -40000 -46870 40000
rect -46622 -40000 -46552 40000
rect -46304 -40000 -46234 40000
rect -45986 -40000 -45916 40000
rect -45668 -40000 -45598 40000
rect -45350 -40000 -45280 40000
rect -45032 -40000 -44962 40000
rect -44714 -40000 -44644 40000
rect -44396 -40000 -44326 40000
rect -44078 -40000 -44008 40000
rect -43760 -40000 -43690 40000
rect -43442 -40000 -43372 40000
rect -43124 -40000 -43054 40000
rect -42806 -40000 -42736 40000
rect -42488 -40000 -42418 40000
rect -42170 -40000 -42100 40000
rect -41852 -40000 -41782 40000
rect -41534 -40000 -41464 40000
rect -41216 -40000 -41146 40000
rect -40898 -40000 -40828 40000
rect -40580 -40000 -40510 40000
rect -40262 -40000 -40192 40000
rect -39944 -40000 -39874 40000
rect -39626 -40000 -39556 40000
rect -39308 -40000 -39238 40000
rect -38990 -40000 -38920 40000
rect -38672 -40000 -38602 40000
rect -38354 -40000 -38284 40000
rect -38036 -40000 -37966 40000
rect -37718 -40000 -37648 40000
rect -37400 -40000 -37330 40000
rect -37082 -40000 -37012 40000
rect -36764 -40000 -36694 40000
rect -36446 -40000 -36376 40000
rect -36128 -40000 -36058 40000
rect -35810 -40000 -35740 40000
rect -35492 -40000 -35422 40000
rect -35174 -40000 -35104 40000
rect -34856 -40000 -34786 40000
rect -34538 -40000 -34468 40000
rect -34220 -40000 -34150 40000
rect -33902 -40000 -33832 40000
rect -33584 -40000 -33514 40000
rect -33266 -40000 -33196 40000
rect -32948 -40000 -32878 40000
rect -32630 -40000 -32560 40000
rect -32312 -40000 -32242 40000
rect -31994 -40000 -31924 40000
rect -31676 -40000 -31606 40000
rect -31358 -40000 -31288 40000
rect -31040 -40000 -30970 40000
rect -30722 -40000 -30652 40000
rect -30404 -40000 -30334 40000
rect -30086 -40000 -30016 40000
rect -29768 -40000 -29698 40000
rect -29450 -40000 -29380 40000
rect -29132 -40000 -29062 40000
rect -28814 -40000 -28744 40000
rect -28496 -40000 -28426 40000
rect -28178 -40000 -28108 40000
rect -27860 -40000 -27790 40000
rect -27542 -40000 -27472 40000
rect -27224 -40000 -27154 40000
rect -26906 -40000 -26836 40000
rect -26588 -40000 -26518 40000
rect -26270 -40000 -26200 40000
rect -25952 -40000 -25882 40000
rect -25634 -40000 -25564 40000
rect -25316 -40000 -25246 40000
rect -24998 -40000 -24928 40000
rect -24680 -40000 -24610 40000
rect -24362 -40000 -24292 40000
rect -24044 -40000 -23974 40000
rect -23726 -40000 -23656 40000
rect -23408 -40000 -23338 40000
rect -23090 -40000 -23020 40000
rect -22772 -40000 -22702 40000
rect -22454 -40000 -22384 40000
rect -22136 -40000 -22066 40000
rect -21818 -40000 -21748 40000
rect -21500 -40000 -21430 40000
rect -21182 -40000 -21112 40000
rect -20864 -40000 -20794 40000
rect -20546 -40000 -20476 40000
rect -20228 -40000 -20158 40000
rect -19910 -40000 -19840 40000
rect -19592 -40000 -19522 40000
rect -19274 -40000 -19204 40000
rect -18956 -40000 -18886 40000
rect -18638 -40000 -18568 40000
rect -18320 -40000 -18250 40000
rect -18002 -40000 -17932 40000
rect -17684 -40000 -17614 40000
rect -17366 -40000 -17296 40000
rect -17048 -40000 -16978 40000
rect -16730 -40000 -16660 40000
rect -16412 -40000 -16342 40000
rect -16094 -40000 -16024 40000
rect -15776 -40000 -15706 40000
rect -15458 -40000 -15388 40000
rect -15140 -40000 -15070 40000
rect -14822 -40000 -14752 40000
rect -14504 -40000 -14434 40000
rect -14186 -40000 -14116 40000
rect -13868 -40000 -13798 40000
rect -13550 -40000 -13480 40000
rect -13232 -40000 -13162 40000
rect -12914 -40000 -12844 40000
rect -12596 -40000 -12526 40000
rect -12278 -40000 -12208 40000
rect -11960 -40000 -11890 40000
rect -11642 -40000 -11572 40000
rect -11324 -40000 -11254 40000
rect -11006 -40000 -10936 40000
rect -10688 -40000 -10618 40000
rect -10370 -40000 -10300 40000
rect -10052 -40000 -9982 40000
rect -9734 -40000 -9664 40000
rect -9416 -40000 -9346 40000
rect -9098 -40000 -9028 40000
rect -8780 -40000 -8710 40000
rect -8462 -40000 -8392 40000
rect -8144 -40000 -8074 40000
rect -7826 -40000 -7756 40000
rect -7508 -40000 -7438 40000
rect -7190 -40000 -7120 40000
rect -6872 -40000 -6802 40000
rect -6554 -40000 -6484 40000
rect -6236 -40000 -6166 40000
rect -5918 -40000 -5848 40000
rect -5600 -40000 -5530 40000
rect -5282 -40000 -5212 40000
rect -4964 -40000 -4894 40000
rect -4646 -40000 -4576 40000
rect -4328 -40000 -4258 40000
rect -4010 -40000 -3940 40000
rect -3692 -40000 -3622 40000
rect -3374 -40000 -3304 40000
rect -3056 -40000 -2986 40000
rect -2738 -40000 -2668 40000
rect -2420 -40000 -2350 40000
rect -2102 -40000 -2032 40000
rect -1784 -40000 -1714 40000
rect -1466 -40000 -1396 40000
rect -1148 -40000 -1078 40000
rect -830 -40000 -760 40000
rect -512 -40000 -442 40000
rect -194 -40000 -124 40000
rect 124 -40000 194 40000
rect 442 -40000 512 40000
rect 760 -40000 830 40000
rect 1078 -40000 1148 40000
rect 1396 -40000 1466 40000
rect 1714 -40000 1784 40000
rect 2032 -40000 2102 40000
rect 2350 -40000 2420 40000
rect 2668 -40000 2738 40000
rect 2986 -40000 3056 40000
rect 3304 -40000 3374 40000
rect 3622 -40000 3692 40000
rect 3940 -40000 4010 40000
rect 4258 -40000 4328 40000
rect 4576 -40000 4646 40000
rect 4894 -40000 4964 40000
rect 5212 -40000 5282 40000
rect 5530 -40000 5600 40000
rect 5848 -40000 5918 40000
rect 6166 -40000 6236 40000
rect 6484 -40000 6554 40000
rect 6802 -40000 6872 40000
rect 7120 -40000 7190 40000
rect 7438 -40000 7508 40000
rect 7756 -40000 7826 40000
rect 8074 -40000 8144 40000
rect 8392 -40000 8462 40000
rect 8710 -40000 8780 40000
rect 9028 -40000 9098 40000
rect 9346 -40000 9416 40000
rect 9664 -40000 9734 40000
rect 9982 -40000 10052 40000
rect 10300 -40000 10370 40000
rect 10618 -40000 10688 40000
rect 10936 -40000 11006 40000
rect 11254 -40000 11324 40000
rect 11572 -40000 11642 40000
rect 11890 -40000 11960 40000
rect 12208 -40000 12278 40000
rect 12526 -40000 12596 40000
rect 12844 -40000 12914 40000
rect 13162 -40000 13232 40000
rect 13480 -40000 13550 40000
rect 13798 -40000 13868 40000
rect 14116 -40000 14186 40000
rect 14434 -40000 14504 40000
rect 14752 -40000 14822 40000
rect 15070 -40000 15140 40000
rect 15388 -40000 15458 40000
rect 15706 -40000 15776 40000
rect 16024 -40000 16094 40000
rect 16342 -40000 16412 40000
rect 16660 -40000 16730 40000
rect 16978 -40000 17048 40000
rect 17296 -40000 17366 40000
rect 17614 -40000 17684 40000
rect 17932 -40000 18002 40000
rect 18250 -40000 18320 40000
rect 18568 -40000 18638 40000
rect 18886 -40000 18956 40000
rect 19204 -40000 19274 40000
rect 19522 -40000 19592 40000
rect 19840 -40000 19910 40000
rect 20158 -40000 20228 40000
rect 20476 -40000 20546 40000
rect 20794 -40000 20864 40000
rect 21112 -40000 21182 40000
rect 21430 -40000 21500 40000
rect 21748 -40000 21818 40000
rect 22066 -40000 22136 40000
rect 22384 -40000 22454 40000
rect 22702 -40000 22772 40000
rect 23020 -40000 23090 40000
rect 23338 -40000 23408 40000
rect 23656 -40000 23726 40000
rect 23974 -40000 24044 40000
rect 24292 -40000 24362 40000
rect 24610 -40000 24680 40000
rect 24928 -40000 24998 40000
rect 25246 -40000 25316 40000
rect 25564 -40000 25634 40000
rect 25882 -40000 25952 40000
rect 26200 -40000 26270 40000
rect 26518 -40000 26588 40000
rect 26836 -40000 26906 40000
rect 27154 -40000 27224 40000
rect 27472 -40000 27542 40000
rect 27790 -40000 27860 40000
rect 28108 -40000 28178 40000
rect 28426 -40000 28496 40000
rect 28744 -40000 28814 40000
rect 29062 -40000 29132 40000
rect 29380 -40000 29450 40000
rect 29698 -40000 29768 40000
rect 30016 -40000 30086 40000
rect 30334 -40000 30404 40000
rect 30652 -40000 30722 40000
rect 30970 -40000 31040 40000
rect 31288 -40000 31358 40000
rect 31606 -40000 31676 40000
rect 31924 -40000 31994 40000
rect 32242 -40000 32312 40000
rect 32560 -40000 32630 40000
rect 32878 -40000 32948 40000
rect 33196 -40000 33266 40000
rect 33514 -40000 33584 40000
rect 33832 -40000 33902 40000
rect 34150 -40000 34220 40000
rect 34468 -40000 34538 40000
rect 34786 -40000 34856 40000
rect 35104 -40000 35174 40000
rect 35422 -40000 35492 40000
rect 35740 -40000 35810 40000
rect 36058 -40000 36128 40000
rect 36376 -40000 36446 40000
rect 36694 -40000 36764 40000
rect 37012 -40000 37082 40000
rect 37330 -40000 37400 40000
rect 37648 -40000 37718 40000
rect 37966 -40000 38036 40000
rect 38284 -40000 38354 40000
rect 38602 -40000 38672 40000
rect 38920 -40000 38990 40000
rect 39238 -40000 39308 40000
rect 39556 -40000 39626 40000
rect 39874 -40000 39944 40000
rect 40192 -40000 40262 40000
rect 40510 -40000 40580 40000
rect 40828 -40000 40898 40000
rect 41146 -40000 41216 40000
rect 41464 -40000 41534 40000
rect 41782 -40000 41852 40000
rect 42100 -40000 42170 40000
rect 42418 -40000 42488 40000
rect 42736 -40000 42806 40000
rect 43054 -40000 43124 40000
rect 43372 -40000 43442 40000
rect 43690 -40000 43760 40000
rect 44008 -40000 44078 40000
rect 44326 -40000 44396 40000
rect 44644 -40000 44714 40000
rect 44962 -40000 45032 40000
rect 45280 -40000 45350 40000
rect 45598 -40000 45668 40000
rect 45916 -40000 45986 40000
rect 46234 -40000 46304 40000
rect 46552 -40000 46622 40000
rect 46870 -40000 46940 40000
rect 47188 -40000 47258 40000
rect 47506 -40000 47576 40000
rect 47824 -40000 47894 40000
rect 48142 -40000 48212 40000
rect 48460 -40000 48530 40000
rect 48778 -40000 48848 40000
rect 49096 -40000 49166 40000
rect 49414 -40000 49484 40000
rect 49732 -40000 49802 40000
rect 50050 -40000 50120 40000
rect 50368 -40000 50438 40000
rect 50686 -40000 50756 40000
rect 51004 -40000 51074 40000
rect 51322 -40000 51392 40000
rect 51640 -40000 51710 40000
rect 51958 -40000 52028 40000
rect 52276 -40000 52346 40000
rect 52594 -40000 52664 40000
rect 52912 -40000 52982 40000
rect 53230 -40000 53300 40000
rect 53548 -40000 53618 40000
rect 53866 -40000 53936 40000
rect 54184 -40000 54254 40000
rect 54502 -40000 54572 40000
rect 54820 -40000 54890 40000
rect 55138 -40000 55208 40000
rect 55456 -40000 55526 40000
rect 55774 -40000 55844 40000
rect 56092 -40000 56162 40000
rect 56410 -40000 56480 40000
rect 56728 -40000 56798 40000
rect 57046 -40000 57116 40000
rect 57364 -40000 57434 40000
rect 57682 -40000 57752 40000
rect 58000 -40000 58070 40000
rect 58318 -40000 58388 40000
rect 58636 -40000 58706 40000
rect 58954 -40000 59024 40000
rect 59272 -40000 59342 40000
rect 59590 -40000 59660 40000
rect 59908 -40000 59978 40000
rect 60226 -40000 60296 40000
rect 60544 -40000 60614 40000
rect 60862 -40000 60932 40000
rect 61180 -40000 61250 40000
rect 61498 -40000 61568 40000
rect 61816 -40000 61886 40000
rect 62134 -40000 62204 40000
rect 62452 -40000 62522 40000
rect 62770 -40000 62840 40000
rect 63088 -40000 63158 40000
rect 63406 -40000 63476 40000
<< locali >>
rect -63606 40528 -63510 40562
rect 63510 40528 63606 40562
rect -63606 40466 -63572 40528
rect 63572 40466 63606 40528
rect -63606 -40528 -63572 -40466
rect 63572 -40528 63606 -40466
rect -63606 -40562 -63510 -40528
rect 63510 -40562 63606 -40528
<< viali >>
rect -63460 40017 -63422 40414
rect -63142 40017 -63104 40414
rect -62824 40017 -62786 40414
rect -62506 40017 -62468 40414
rect -62188 40017 -62150 40414
rect -61870 40017 -61832 40414
rect -61552 40017 -61514 40414
rect -61234 40017 -61196 40414
rect -60916 40017 -60878 40414
rect -60598 40017 -60560 40414
rect -60280 40017 -60242 40414
rect -59962 40017 -59924 40414
rect -59644 40017 -59606 40414
rect -59326 40017 -59288 40414
rect -59008 40017 -58970 40414
rect -58690 40017 -58652 40414
rect -58372 40017 -58334 40414
rect -58054 40017 -58016 40414
rect -57736 40017 -57698 40414
rect -57418 40017 -57380 40414
rect -57100 40017 -57062 40414
rect -56782 40017 -56744 40414
rect -56464 40017 -56426 40414
rect -56146 40017 -56108 40414
rect -55828 40017 -55790 40414
rect -55510 40017 -55472 40414
rect -55192 40017 -55154 40414
rect -54874 40017 -54836 40414
rect -54556 40017 -54518 40414
rect -54238 40017 -54200 40414
rect -53920 40017 -53882 40414
rect -53602 40017 -53564 40414
rect -53284 40017 -53246 40414
rect -52966 40017 -52928 40414
rect -52648 40017 -52610 40414
rect -52330 40017 -52292 40414
rect -52012 40017 -51974 40414
rect -51694 40017 -51656 40414
rect -51376 40017 -51338 40414
rect -51058 40017 -51020 40414
rect -50740 40017 -50702 40414
rect -50422 40017 -50384 40414
rect -50104 40017 -50066 40414
rect -49786 40017 -49748 40414
rect -49468 40017 -49430 40414
rect -49150 40017 -49112 40414
rect -48832 40017 -48794 40414
rect -48514 40017 -48476 40414
rect -48196 40017 -48158 40414
rect -47878 40017 -47840 40414
rect -47560 40017 -47522 40414
rect -47242 40017 -47204 40414
rect -46924 40017 -46886 40414
rect -46606 40017 -46568 40414
rect -46288 40017 -46250 40414
rect -45970 40017 -45932 40414
rect -45652 40017 -45614 40414
rect -45334 40017 -45296 40414
rect -45016 40017 -44978 40414
rect -44698 40017 -44660 40414
rect -44380 40017 -44342 40414
rect -44062 40017 -44024 40414
rect -43744 40017 -43706 40414
rect -43426 40017 -43388 40414
rect -43108 40017 -43070 40414
rect -42790 40017 -42752 40414
rect -42472 40017 -42434 40414
rect -42154 40017 -42116 40414
rect -41836 40017 -41798 40414
rect -41518 40017 -41480 40414
rect -41200 40017 -41162 40414
rect -40882 40017 -40844 40414
rect -40564 40017 -40526 40414
rect -40246 40017 -40208 40414
rect -39928 40017 -39890 40414
rect -39610 40017 -39572 40414
rect -39292 40017 -39254 40414
rect -38974 40017 -38936 40414
rect -38656 40017 -38618 40414
rect -38338 40017 -38300 40414
rect -38020 40017 -37982 40414
rect -37702 40017 -37664 40414
rect -37384 40017 -37346 40414
rect -37066 40017 -37028 40414
rect -36748 40017 -36710 40414
rect -36430 40017 -36392 40414
rect -36112 40017 -36074 40414
rect -35794 40017 -35756 40414
rect -35476 40017 -35438 40414
rect -35158 40017 -35120 40414
rect -34840 40017 -34802 40414
rect -34522 40017 -34484 40414
rect -34204 40017 -34166 40414
rect -33886 40017 -33848 40414
rect -33568 40017 -33530 40414
rect -33250 40017 -33212 40414
rect -32932 40017 -32894 40414
rect -32614 40017 -32576 40414
rect -32296 40017 -32258 40414
rect -31978 40017 -31940 40414
rect -31660 40017 -31622 40414
rect -31342 40017 -31304 40414
rect -31024 40017 -30986 40414
rect -30706 40017 -30668 40414
rect -30388 40017 -30350 40414
rect -30070 40017 -30032 40414
rect -29752 40017 -29714 40414
rect -29434 40017 -29396 40414
rect -29116 40017 -29078 40414
rect -28798 40017 -28760 40414
rect -28480 40017 -28442 40414
rect -28162 40017 -28124 40414
rect -27844 40017 -27806 40414
rect -27526 40017 -27488 40414
rect -27208 40017 -27170 40414
rect -26890 40017 -26852 40414
rect -26572 40017 -26534 40414
rect -26254 40017 -26216 40414
rect -25936 40017 -25898 40414
rect -25618 40017 -25580 40414
rect -25300 40017 -25262 40414
rect -24982 40017 -24944 40414
rect -24664 40017 -24626 40414
rect -24346 40017 -24308 40414
rect -24028 40017 -23990 40414
rect -23710 40017 -23672 40414
rect -23392 40017 -23354 40414
rect -23074 40017 -23036 40414
rect -22756 40017 -22718 40414
rect -22438 40017 -22400 40414
rect -22120 40017 -22082 40414
rect -21802 40017 -21764 40414
rect -21484 40017 -21446 40414
rect -21166 40017 -21128 40414
rect -20848 40017 -20810 40414
rect -20530 40017 -20492 40414
rect -20212 40017 -20174 40414
rect -19894 40017 -19856 40414
rect -19576 40017 -19538 40414
rect -19258 40017 -19220 40414
rect -18940 40017 -18902 40414
rect -18622 40017 -18584 40414
rect -18304 40017 -18266 40414
rect -17986 40017 -17948 40414
rect -17668 40017 -17630 40414
rect -17350 40017 -17312 40414
rect -17032 40017 -16994 40414
rect -16714 40017 -16676 40414
rect -16396 40017 -16358 40414
rect -16078 40017 -16040 40414
rect -15760 40017 -15722 40414
rect -15442 40017 -15404 40414
rect -15124 40017 -15086 40414
rect -14806 40017 -14768 40414
rect -14488 40017 -14450 40414
rect -14170 40017 -14132 40414
rect -13852 40017 -13814 40414
rect -13534 40017 -13496 40414
rect -13216 40017 -13178 40414
rect -12898 40017 -12860 40414
rect -12580 40017 -12542 40414
rect -12262 40017 -12224 40414
rect -11944 40017 -11906 40414
rect -11626 40017 -11588 40414
rect -11308 40017 -11270 40414
rect -10990 40017 -10952 40414
rect -10672 40017 -10634 40414
rect -10354 40017 -10316 40414
rect -10036 40017 -9998 40414
rect -9718 40017 -9680 40414
rect -9400 40017 -9362 40414
rect -9082 40017 -9044 40414
rect -8764 40017 -8726 40414
rect -8446 40017 -8408 40414
rect -8128 40017 -8090 40414
rect -7810 40017 -7772 40414
rect -7492 40017 -7454 40414
rect -7174 40017 -7136 40414
rect -6856 40017 -6818 40414
rect -6538 40017 -6500 40414
rect -6220 40017 -6182 40414
rect -5902 40017 -5864 40414
rect -5584 40017 -5546 40414
rect -5266 40017 -5228 40414
rect -4948 40017 -4910 40414
rect -4630 40017 -4592 40414
rect -4312 40017 -4274 40414
rect -3994 40017 -3956 40414
rect -3676 40017 -3638 40414
rect -3358 40017 -3320 40414
rect -3040 40017 -3002 40414
rect -2722 40017 -2684 40414
rect -2404 40017 -2366 40414
rect -2086 40017 -2048 40414
rect -1768 40017 -1730 40414
rect -1450 40017 -1412 40414
rect -1132 40017 -1094 40414
rect -814 40017 -776 40414
rect -496 40017 -458 40414
rect -178 40017 -140 40414
rect 140 40017 178 40414
rect 458 40017 496 40414
rect 776 40017 814 40414
rect 1094 40017 1132 40414
rect 1412 40017 1450 40414
rect 1730 40017 1768 40414
rect 2048 40017 2086 40414
rect 2366 40017 2404 40414
rect 2684 40017 2722 40414
rect 3002 40017 3040 40414
rect 3320 40017 3358 40414
rect 3638 40017 3676 40414
rect 3956 40017 3994 40414
rect 4274 40017 4312 40414
rect 4592 40017 4630 40414
rect 4910 40017 4948 40414
rect 5228 40017 5266 40414
rect 5546 40017 5584 40414
rect 5864 40017 5902 40414
rect 6182 40017 6220 40414
rect 6500 40017 6538 40414
rect 6818 40017 6856 40414
rect 7136 40017 7174 40414
rect 7454 40017 7492 40414
rect 7772 40017 7810 40414
rect 8090 40017 8128 40414
rect 8408 40017 8446 40414
rect 8726 40017 8764 40414
rect 9044 40017 9082 40414
rect 9362 40017 9400 40414
rect 9680 40017 9718 40414
rect 9998 40017 10036 40414
rect 10316 40017 10354 40414
rect 10634 40017 10672 40414
rect 10952 40017 10990 40414
rect 11270 40017 11308 40414
rect 11588 40017 11626 40414
rect 11906 40017 11944 40414
rect 12224 40017 12262 40414
rect 12542 40017 12580 40414
rect 12860 40017 12898 40414
rect 13178 40017 13216 40414
rect 13496 40017 13534 40414
rect 13814 40017 13852 40414
rect 14132 40017 14170 40414
rect 14450 40017 14488 40414
rect 14768 40017 14806 40414
rect 15086 40017 15124 40414
rect 15404 40017 15442 40414
rect 15722 40017 15760 40414
rect 16040 40017 16078 40414
rect 16358 40017 16396 40414
rect 16676 40017 16714 40414
rect 16994 40017 17032 40414
rect 17312 40017 17350 40414
rect 17630 40017 17668 40414
rect 17948 40017 17986 40414
rect 18266 40017 18304 40414
rect 18584 40017 18622 40414
rect 18902 40017 18940 40414
rect 19220 40017 19258 40414
rect 19538 40017 19576 40414
rect 19856 40017 19894 40414
rect 20174 40017 20212 40414
rect 20492 40017 20530 40414
rect 20810 40017 20848 40414
rect 21128 40017 21166 40414
rect 21446 40017 21484 40414
rect 21764 40017 21802 40414
rect 22082 40017 22120 40414
rect 22400 40017 22438 40414
rect 22718 40017 22756 40414
rect 23036 40017 23074 40414
rect 23354 40017 23392 40414
rect 23672 40017 23710 40414
rect 23990 40017 24028 40414
rect 24308 40017 24346 40414
rect 24626 40017 24664 40414
rect 24944 40017 24982 40414
rect 25262 40017 25300 40414
rect 25580 40017 25618 40414
rect 25898 40017 25936 40414
rect 26216 40017 26254 40414
rect 26534 40017 26572 40414
rect 26852 40017 26890 40414
rect 27170 40017 27208 40414
rect 27488 40017 27526 40414
rect 27806 40017 27844 40414
rect 28124 40017 28162 40414
rect 28442 40017 28480 40414
rect 28760 40017 28798 40414
rect 29078 40017 29116 40414
rect 29396 40017 29434 40414
rect 29714 40017 29752 40414
rect 30032 40017 30070 40414
rect 30350 40017 30388 40414
rect 30668 40017 30706 40414
rect 30986 40017 31024 40414
rect 31304 40017 31342 40414
rect 31622 40017 31660 40414
rect 31940 40017 31978 40414
rect 32258 40017 32296 40414
rect 32576 40017 32614 40414
rect 32894 40017 32932 40414
rect 33212 40017 33250 40414
rect 33530 40017 33568 40414
rect 33848 40017 33886 40414
rect 34166 40017 34204 40414
rect 34484 40017 34522 40414
rect 34802 40017 34840 40414
rect 35120 40017 35158 40414
rect 35438 40017 35476 40414
rect 35756 40017 35794 40414
rect 36074 40017 36112 40414
rect 36392 40017 36430 40414
rect 36710 40017 36748 40414
rect 37028 40017 37066 40414
rect 37346 40017 37384 40414
rect 37664 40017 37702 40414
rect 37982 40017 38020 40414
rect 38300 40017 38338 40414
rect 38618 40017 38656 40414
rect 38936 40017 38974 40414
rect 39254 40017 39292 40414
rect 39572 40017 39610 40414
rect 39890 40017 39928 40414
rect 40208 40017 40246 40414
rect 40526 40017 40564 40414
rect 40844 40017 40882 40414
rect 41162 40017 41200 40414
rect 41480 40017 41518 40414
rect 41798 40017 41836 40414
rect 42116 40017 42154 40414
rect 42434 40017 42472 40414
rect 42752 40017 42790 40414
rect 43070 40017 43108 40414
rect 43388 40017 43426 40414
rect 43706 40017 43744 40414
rect 44024 40017 44062 40414
rect 44342 40017 44380 40414
rect 44660 40017 44698 40414
rect 44978 40017 45016 40414
rect 45296 40017 45334 40414
rect 45614 40017 45652 40414
rect 45932 40017 45970 40414
rect 46250 40017 46288 40414
rect 46568 40017 46606 40414
rect 46886 40017 46924 40414
rect 47204 40017 47242 40414
rect 47522 40017 47560 40414
rect 47840 40017 47878 40414
rect 48158 40017 48196 40414
rect 48476 40017 48514 40414
rect 48794 40017 48832 40414
rect 49112 40017 49150 40414
rect 49430 40017 49468 40414
rect 49748 40017 49786 40414
rect 50066 40017 50104 40414
rect 50384 40017 50422 40414
rect 50702 40017 50740 40414
rect 51020 40017 51058 40414
rect 51338 40017 51376 40414
rect 51656 40017 51694 40414
rect 51974 40017 52012 40414
rect 52292 40017 52330 40414
rect 52610 40017 52648 40414
rect 52928 40017 52966 40414
rect 53246 40017 53284 40414
rect 53564 40017 53602 40414
rect 53882 40017 53920 40414
rect 54200 40017 54238 40414
rect 54518 40017 54556 40414
rect 54836 40017 54874 40414
rect 55154 40017 55192 40414
rect 55472 40017 55510 40414
rect 55790 40017 55828 40414
rect 56108 40017 56146 40414
rect 56426 40017 56464 40414
rect 56744 40017 56782 40414
rect 57062 40017 57100 40414
rect 57380 40017 57418 40414
rect 57698 40017 57736 40414
rect 58016 40017 58054 40414
rect 58334 40017 58372 40414
rect 58652 40017 58690 40414
rect 58970 40017 59008 40414
rect 59288 40017 59326 40414
rect 59606 40017 59644 40414
rect 59924 40017 59962 40414
rect 60242 40017 60280 40414
rect 60560 40017 60598 40414
rect 60878 40017 60916 40414
rect 61196 40017 61234 40414
rect 61514 40017 61552 40414
rect 61832 40017 61870 40414
rect 62150 40017 62188 40414
rect 62468 40017 62506 40414
rect 62786 40017 62824 40414
rect 63104 40017 63142 40414
rect 63422 40017 63460 40414
rect -63460 -40414 -63422 -40017
rect -63142 -40414 -63104 -40017
rect -62824 -40414 -62786 -40017
rect -62506 -40414 -62468 -40017
rect -62188 -40414 -62150 -40017
rect -61870 -40414 -61832 -40017
rect -61552 -40414 -61514 -40017
rect -61234 -40414 -61196 -40017
rect -60916 -40414 -60878 -40017
rect -60598 -40414 -60560 -40017
rect -60280 -40414 -60242 -40017
rect -59962 -40414 -59924 -40017
rect -59644 -40414 -59606 -40017
rect -59326 -40414 -59288 -40017
rect -59008 -40414 -58970 -40017
rect -58690 -40414 -58652 -40017
rect -58372 -40414 -58334 -40017
rect -58054 -40414 -58016 -40017
rect -57736 -40414 -57698 -40017
rect -57418 -40414 -57380 -40017
rect -57100 -40414 -57062 -40017
rect -56782 -40414 -56744 -40017
rect -56464 -40414 -56426 -40017
rect -56146 -40414 -56108 -40017
rect -55828 -40414 -55790 -40017
rect -55510 -40414 -55472 -40017
rect -55192 -40414 -55154 -40017
rect -54874 -40414 -54836 -40017
rect -54556 -40414 -54518 -40017
rect -54238 -40414 -54200 -40017
rect -53920 -40414 -53882 -40017
rect -53602 -40414 -53564 -40017
rect -53284 -40414 -53246 -40017
rect -52966 -40414 -52928 -40017
rect -52648 -40414 -52610 -40017
rect -52330 -40414 -52292 -40017
rect -52012 -40414 -51974 -40017
rect -51694 -40414 -51656 -40017
rect -51376 -40414 -51338 -40017
rect -51058 -40414 -51020 -40017
rect -50740 -40414 -50702 -40017
rect -50422 -40414 -50384 -40017
rect -50104 -40414 -50066 -40017
rect -49786 -40414 -49748 -40017
rect -49468 -40414 -49430 -40017
rect -49150 -40414 -49112 -40017
rect -48832 -40414 -48794 -40017
rect -48514 -40414 -48476 -40017
rect -48196 -40414 -48158 -40017
rect -47878 -40414 -47840 -40017
rect -47560 -40414 -47522 -40017
rect -47242 -40414 -47204 -40017
rect -46924 -40414 -46886 -40017
rect -46606 -40414 -46568 -40017
rect -46288 -40414 -46250 -40017
rect -45970 -40414 -45932 -40017
rect -45652 -40414 -45614 -40017
rect -45334 -40414 -45296 -40017
rect -45016 -40414 -44978 -40017
rect -44698 -40414 -44660 -40017
rect -44380 -40414 -44342 -40017
rect -44062 -40414 -44024 -40017
rect -43744 -40414 -43706 -40017
rect -43426 -40414 -43388 -40017
rect -43108 -40414 -43070 -40017
rect -42790 -40414 -42752 -40017
rect -42472 -40414 -42434 -40017
rect -42154 -40414 -42116 -40017
rect -41836 -40414 -41798 -40017
rect -41518 -40414 -41480 -40017
rect -41200 -40414 -41162 -40017
rect -40882 -40414 -40844 -40017
rect -40564 -40414 -40526 -40017
rect -40246 -40414 -40208 -40017
rect -39928 -40414 -39890 -40017
rect -39610 -40414 -39572 -40017
rect -39292 -40414 -39254 -40017
rect -38974 -40414 -38936 -40017
rect -38656 -40414 -38618 -40017
rect -38338 -40414 -38300 -40017
rect -38020 -40414 -37982 -40017
rect -37702 -40414 -37664 -40017
rect -37384 -40414 -37346 -40017
rect -37066 -40414 -37028 -40017
rect -36748 -40414 -36710 -40017
rect -36430 -40414 -36392 -40017
rect -36112 -40414 -36074 -40017
rect -35794 -40414 -35756 -40017
rect -35476 -40414 -35438 -40017
rect -35158 -40414 -35120 -40017
rect -34840 -40414 -34802 -40017
rect -34522 -40414 -34484 -40017
rect -34204 -40414 -34166 -40017
rect -33886 -40414 -33848 -40017
rect -33568 -40414 -33530 -40017
rect -33250 -40414 -33212 -40017
rect -32932 -40414 -32894 -40017
rect -32614 -40414 -32576 -40017
rect -32296 -40414 -32258 -40017
rect -31978 -40414 -31940 -40017
rect -31660 -40414 -31622 -40017
rect -31342 -40414 -31304 -40017
rect -31024 -40414 -30986 -40017
rect -30706 -40414 -30668 -40017
rect -30388 -40414 -30350 -40017
rect -30070 -40414 -30032 -40017
rect -29752 -40414 -29714 -40017
rect -29434 -40414 -29396 -40017
rect -29116 -40414 -29078 -40017
rect -28798 -40414 -28760 -40017
rect -28480 -40414 -28442 -40017
rect -28162 -40414 -28124 -40017
rect -27844 -40414 -27806 -40017
rect -27526 -40414 -27488 -40017
rect -27208 -40414 -27170 -40017
rect -26890 -40414 -26852 -40017
rect -26572 -40414 -26534 -40017
rect -26254 -40414 -26216 -40017
rect -25936 -40414 -25898 -40017
rect -25618 -40414 -25580 -40017
rect -25300 -40414 -25262 -40017
rect -24982 -40414 -24944 -40017
rect -24664 -40414 -24626 -40017
rect -24346 -40414 -24308 -40017
rect -24028 -40414 -23990 -40017
rect -23710 -40414 -23672 -40017
rect -23392 -40414 -23354 -40017
rect -23074 -40414 -23036 -40017
rect -22756 -40414 -22718 -40017
rect -22438 -40414 -22400 -40017
rect -22120 -40414 -22082 -40017
rect -21802 -40414 -21764 -40017
rect -21484 -40414 -21446 -40017
rect -21166 -40414 -21128 -40017
rect -20848 -40414 -20810 -40017
rect -20530 -40414 -20492 -40017
rect -20212 -40414 -20174 -40017
rect -19894 -40414 -19856 -40017
rect -19576 -40414 -19538 -40017
rect -19258 -40414 -19220 -40017
rect -18940 -40414 -18902 -40017
rect -18622 -40414 -18584 -40017
rect -18304 -40414 -18266 -40017
rect -17986 -40414 -17948 -40017
rect -17668 -40414 -17630 -40017
rect -17350 -40414 -17312 -40017
rect -17032 -40414 -16994 -40017
rect -16714 -40414 -16676 -40017
rect -16396 -40414 -16358 -40017
rect -16078 -40414 -16040 -40017
rect -15760 -40414 -15722 -40017
rect -15442 -40414 -15404 -40017
rect -15124 -40414 -15086 -40017
rect -14806 -40414 -14768 -40017
rect -14488 -40414 -14450 -40017
rect -14170 -40414 -14132 -40017
rect -13852 -40414 -13814 -40017
rect -13534 -40414 -13496 -40017
rect -13216 -40414 -13178 -40017
rect -12898 -40414 -12860 -40017
rect -12580 -40414 -12542 -40017
rect -12262 -40414 -12224 -40017
rect -11944 -40414 -11906 -40017
rect -11626 -40414 -11588 -40017
rect -11308 -40414 -11270 -40017
rect -10990 -40414 -10952 -40017
rect -10672 -40414 -10634 -40017
rect -10354 -40414 -10316 -40017
rect -10036 -40414 -9998 -40017
rect -9718 -40414 -9680 -40017
rect -9400 -40414 -9362 -40017
rect -9082 -40414 -9044 -40017
rect -8764 -40414 -8726 -40017
rect -8446 -40414 -8408 -40017
rect -8128 -40414 -8090 -40017
rect -7810 -40414 -7772 -40017
rect -7492 -40414 -7454 -40017
rect -7174 -40414 -7136 -40017
rect -6856 -40414 -6818 -40017
rect -6538 -40414 -6500 -40017
rect -6220 -40414 -6182 -40017
rect -5902 -40414 -5864 -40017
rect -5584 -40414 -5546 -40017
rect -5266 -40414 -5228 -40017
rect -4948 -40414 -4910 -40017
rect -4630 -40414 -4592 -40017
rect -4312 -40414 -4274 -40017
rect -3994 -40414 -3956 -40017
rect -3676 -40414 -3638 -40017
rect -3358 -40414 -3320 -40017
rect -3040 -40414 -3002 -40017
rect -2722 -40414 -2684 -40017
rect -2404 -40414 -2366 -40017
rect -2086 -40414 -2048 -40017
rect -1768 -40414 -1730 -40017
rect -1450 -40414 -1412 -40017
rect -1132 -40414 -1094 -40017
rect -814 -40414 -776 -40017
rect -496 -40414 -458 -40017
rect -178 -40414 -140 -40017
rect 140 -40414 178 -40017
rect 458 -40414 496 -40017
rect 776 -40414 814 -40017
rect 1094 -40414 1132 -40017
rect 1412 -40414 1450 -40017
rect 1730 -40414 1768 -40017
rect 2048 -40414 2086 -40017
rect 2366 -40414 2404 -40017
rect 2684 -40414 2722 -40017
rect 3002 -40414 3040 -40017
rect 3320 -40414 3358 -40017
rect 3638 -40414 3676 -40017
rect 3956 -40414 3994 -40017
rect 4274 -40414 4312 -40017
rect 4592 -40414 4630 -40017
rect 4910 -40414 4948 -40017
rect 5228 -40414 5266 -40017
rect 5546 -40414 5584 -40017
rect 5864 -40414 5902 -40017
rect 6182 -40414 6220 -40017
rect 6500 -40414 6538 -40017
rect 6818 -40414 6856 -40017
rect 7136 -40414 7174 -40017
rect 7454 -40414 7492 -40017
rect 7772 -40414 7810 -40017
rect 8090 -40414 8128 -40017
rect 8408 -40414 8446 -40017
rect 8726 -40414 8764 -40017
rect 9044 -40414 9082 -40017
rect 9362 -40414 9400 -40017
rect 9680 -40414 9718 -40017
rect 9998 -40414 10036 -40017
rect 10316 -40414 10354 -40017
rect 10634 -40414 10672 -40017
rect 10952 -40414 10990 -40017
rect 11270 -40414 11308 -40017
rect 11588 -40414 11626 -40017
rect 11906 -40414 11944 -40017
rect 12224 -40414 12262 -40017
rect 12542 -40414 12580 -40017
rect 12860 -40414 12898 -40017
rect 13178 -40414 13216 -40017
rect 13496 -40414 13534 -40017
rect 13814 -40414 13852 -40017
rect 14132 -40414 14170 -40017
rect 14450 -40414 14488 -40017
rect 14768 -40414 14806 -40017
rect 15086 -40414 15124 -40017
rect 15404 -40414 15442 -40017
rect 15722 -40414 15760 -40017
rect 16040 -40414 16078 -40017
rect 16358 -40414 16396 -40017
rect 16676 -40414 16714 -40017
rect 16994 -40414 17032 -40017
rect 17312 -40414 17350 -40017
rect 17630 -40414 17668 -40017
rect 17948 -40414 17986 -40017
rect 18266 -40414 18304 -40017
rect 18584 -40414 18622 -40017
rect 18902 -40414 18940 -40017
rect 19220 -40414 19258 -40017
rect 19538 -40414 19576 -40017
rect 19856 -40414 19894 -40017
rect 20174 -40414 20212 -40017
rect 20492 -40414 20530 -40017
rect 20810 -40414 20848 -40017
rect 21128 -40414 21166 -40017
rect 21446 -40414 21484 -40017
rect 21764 -40414 21802 -40017
rect 22082 -40414 22120 -40017
rect 22400 -40414 22438 -40017
rect 22718 -40414 22756 -40017
rect 23036 -40414 23074 -40017
rect 23354 -40414 23392 -40017
rect 23672 -40414 23710 -40017
rect 23990 -40414 24028 -40017
rect 24308 -40414 24346 -40017
rect 24626 -40414 24664 -40017
rect 24944 -40414 24982 -40017
rect 25262 -40414 25300 -40017
rect 25580 -40414 25618 -40017
rect 25898 -40414 25936 -40017
rect 26216 -40414 26254 -40017
rect 26534 -40414 26572 -40017
rect 26852 -40414 26890 -40017
rect 27170 -40414 27208 -40017
rect 27488 -40414 27526 -40017
rect 27806 -40414 27844 -40017
rect 28124 -40414 28162 -40017
rect 28442 -40414 28480 -40017
rect 28760 -40414 28798 -40017
rect 29078 -40414 29116 -40017
rect 29396 -40414 29434 -40017
rect 29714 -40414 29752 -40017
rect 30032 -40414 30070 -40017
rect 30350 -40414 30388 -40017
rect 30668 -40414 30706 -40017
rect 30986 -40414 31024 -40017
rect 31304 -40414 31342 -40017
rect 31622 -40414 31660 -40017
rect 31940 -40414 31978 -40017
rect 32258 -40414 32296 -40017
rect 32576 -40414 32614 -40017
rect 32894 -40414 32932 -40017
rect 33212 -40414 33250 -40017
rect 33530 -40414 33568 -40017
rect 33848 -40414 33886 -40017
rect 34166 -40414 34204 -40017
rect 34484 -40414 34522 -40017
rect 34802 -40414 34840 -40017
rect 35120 -40414 35158 -40017
rect 35438 -40414 35476 -40017
rect 35756 -40414 35794 -40017
rect 36074 -40414 36112 -40017
rect 36392 -40414 36430 -40017
rect 36710 -40414 36748 -40017
rect 37028 -40414 37066 -40017
rect 37346 -40414 37384 -40017
rect 37664 -40414 37702 -40017
rect 37982 -40414 38020 -40017
rect 38300 -40414 38338 -40017
rect 38618 -40414 38656 -40017
rect 38936 -40414 38974 -40017
rect 39254 -40414 39292 -40017
rect 39572 -40414 39610 -40017
rect 39890 -40414 39928 -40017
rect 40208 -40414 40246 -40017
rect 40526 -40414 40564 -40017
rect 40844 -40414 40882 -40017
rect 41162 -40414 41200 -40017
rect 41480 -40414 41518 -40017
rect 41798 -40414 41836 -40017
rect 42116 -40414 42154 -40017
rect 42434 -40414 42472 -40017
rect 42752 -40414 42790 -40017
rect 43070 -40414 43108 -40017
rect 43388 -40414 43426 -40017
rect 43706 -40414 43744 -40017
rect 44024 -40414 44062 -40017
rect 44342 -40414 44380 -40017
rect 44660 -40414 44698 -40017
rect 44978 -40414 45016 -40017
rect 45296 -40414 45334 -40017
rect 45614 -40414 45652 -40017
rect 45932 -40414 45970 -40017
rect 46250 -40414 46288 -40017
rect 46568 -40414 46606 -40017
rect 46886 -40414 46924 -40017
rect 47204 -40414 47242 -40017
rect 47522 -40414 47560 -40017
rect 47840 -40414 47878 -40017
rect 48158 -40414 48196 -40017
rect 48476 -40414 48514 -40017
rect 48794 -40414 48832 -40017
rect 49112 -40414 49150 -40017
rect 49430 -40414 49468 -40017
rect 49748 -40414 49786 -40017
rect 50066 -40414 50104 -40017
rect 50384 -40414 50422 -40017
rect 50702 -40414 50740 -40017
rect 51020 -40414 51058 -40017
rect 51338 -40414 51376 -40017
rect 51656 -40414 51694 -40017
rect 51974 -40414 52012 -40017
rect 52292 -40414 52330 -40017
rect 52610 -40414 52648 -40017
rect 52928 -40414 52966 -40017
rect 53246 -40414 53284 -40017
rect 53564 -40414 53602 -40017
rect 53882 -40414 53920 -40017
rect 54200 -40414 54238 -40017
rect 54518 -40414 54556 -40017
rect 54836 -40414 54874 -40017
rect 55154 -40414 55192 -40017
rect 55472 -40414 55510 -40017
rect 55790 -40414 55828 -40017
rect 56108 -40414 56146 -40017
rect 56426 -40414 56464 -40017
rect 56744 -40414 56782 -40017
rect 57062 -40414 57100 -40017
rect 57380 -40414 57418 -40017
rect 57698 -40414 57736 -40017
rect 58016 -40414 58054 -40017
rect 58334 -40414 58372 -40017
rect 58652 -40414 58690 -40017
rect 58970 -40414 59008 -40017
rect 59288 -40414 59326 -40017
rect 59606 -40414 59644 -40017
rect 59924 -40414 59962 -40017
rect 60242 -40414 60280 -40017
rect 60560 -40414 60598 -40017
rect 60878 -40414 60916 -40017
rect 61196 -40414 61234 -40017
rect 61514 -40414 61552 -40017
rect 61832 -40414 61870 -40017
rect 62150 -40414 62188 -40017
rect 62468 -40414 62506 -40017
rect 62786 -40414 62824 -40017
rect 63104 -40414 63142 -40017
rect 63422 -40414 63460 -40017
<< metal1 >>
rect -63466 40414 -63416 40426
rect -63466 40017 -63460 40414
rect -63422 40017 -63416 40414
rect -63466 40005 -63416 40017
rect -63148 40414 -63098 40426
rect -63148 40017 -63142 40414
rect -63104 40017 -63098 40414
rect -63148 40005 -63098 40017
rect -62830 40414 -62780 40426
rect -62830 40017 -62824 40414
rect -62786 40017 -62780 40414
rect -62830 40005 -62780 40017
rect -62512 40414 -62462 40426
rect -62512 40017 -62506 40414
rect -62468 40017 -62462 40414
rect -62512 40005 -62462 40017
rect -62194 40414 -62144 40426
rect -62194 40017 -62188 40414
rect -62150 40017 -62144 40414
rect -62194 40005 -62144 40017
rect -61876 40414 -61826 40426
rect -61876 40017 -61870 40414
rect -61832 40017 -61826 40414
rect -61876 40005 -61826 40017
rect -61558 40414 -61508 40426
rect -61558 40017 -61552 40414
rect -61514 40017 -61508 40414
rect -61558 40005 -61508 40017
rect -61240 40414 -61190 40426
rect -61240 40017 -61234 40414
rect -61196 40017 -61190 40414
rect -61240 40005 -61190 40017
rect -60922 40414 -60872 40426
rect -60922 40017 -60916 40414
rect -60878 40017 -60872 40414
rect -60922 40005 -60872 40017
rect -60604 40414 -60554 40426
rect -60604 40017 -60598 40414
rect -60560 40017 -60554 40414
rect -60604 40005 -60554 40017
rect -60286 40414 -60236 40426
rect -60286 40017 -60280 40414
rect -60242 40017 -60236 40414
rect -60286 40005 -60236 40017
rect -59968 40414 -59918 40426
rect -59968 40017 -59962 40414
rect -59924 40017 -59918 40414
rect -59968 40005 -59918 40017
rect -59650 40414 -59600 40426
rect -59650 40017 -59644 40414
rect -59606 40017 -59600 40414
rect -59650 40005 -59600 40017
rect -59332 40414 -59282 40426
rect -59332 40017 -59326 40414
rect -59288 40017 -59282 40414
rect -59332 40005 -59282 40017
rect -59014 40414 -58964 40426
rect -59014 40017 -59008 40414
rect -58970 40017 -58964 40414
rect -59014 40005 -58964 40017
rect -58696 40414 -58646 40426
rect -58696 40017 -58690 40414
rect -58652 40017 -58646 40414
rect -58696 40005 -58646 40017
rect -58378 40414 -58328 40426
rect -58378 40017 -58372 40414
rect -58334 40017 -58328 40414
rect -58378 40005 -58328 40017
rect -58060 40414 -58010 40426
rect -58060 40017 -58054 40414
rect -58016 40017 -58010 40414
rect -58060 40005 -58010 40017
rect -57742 40414 -57692 40426
rect -57742 40017 -57736 40414
rect -57698 40017 -57692 40414
rect -57742 40005 -57692 40017
rect -57424 40414 -57374 40426
rect -57424 40017 -57418 40414
rect -57380 40017 -57374 40414
rect -57424 40005 -57374 40017
rect -57106 40414 -57056 40426
rect -57106 40017 -57100 40414
rect -57062 40017 -57056 40414
rect -57106 40005 -57056 40017
rect -56788 40414 -56738 40426
rect -56788 40017 -56782 40414
rect -56744 40017 -56738 40414
rect -56788 40005 -56738 40017
rect -56470 40414 -56420 40426
rect -56470 40017 -56464 40414
rect -56426 40017 -56420 40414
rect -56470 40005 -56420 40017
rect -56152 40414 -56102 40426
rect -56152 40017 -56146 40414
rect -56108 40017 -56102 40414
rect -56152 40005 -56102 40017
rect -55834 40414 -55784 40426
rect -55834 40017 -55828 40414
rect -55790 40017 -55784 40414
rect -55834 40005 -55784 40017
rect -55516 40414 -55466 40426
rect -55516 40017 -55510 40414
rect -55472 40017 -55466 40414
rect -55516 40005 -55466 40017
rect -55198 40414 -55148 40426
rect -55198 40017 -55192 40414
rect -55154 40017 -55148 40414
rect -55198 40005 -55148 40017
rect -54880 40414 -54830 40426
rect -54880 40017 -54874 40414
rect -54836 40017 -54830 40414
rect -54880 40005 -54830 40017
rect -54562 40414 -54512 40426
rect -54562 40017 -54556 40414
rect -54518 40017 -54512 40414
rect -54562 40005 -54512 40017
rect -54244 40414 -54194 40426
rect -54244 40017 -54238 40414
rect -54200 40017 -54194 40414
rect -54244 40005 -54194 40017
rect -53926 40414 -53876 40426
rect -53926 40017 -53920 40414
rect -53882 40017 -53876 40414
rect -53926 40005 -53876 40017
rect -53608 40414 -53558 40426
rect -53608 40017 -53602 40414
rect -53564 40017 -53558 40414
rect -53608 40005 -53558 40017
rect -53290 40414 -53240 40426
rect -53290 40017 -53284 40414
rect -53246 40017 -53240 40414
rect -53290 40005 -53240 40017
rect -52972 40414 -52922 40426
rect -52972 40017 -52966 40414
rect -52928 40017 -52922 40414
rect -52972 40005 -52922 40017
rect -52654 40414 -52604 40426
rect -52654 40017 -52648 40414
rect -52610 40017 -52604 40414
rect -52654 40005 -52604 40017
rect -52336 40414 -52286 40426
rect -52336 40017 -52330 40414
rect -52292 40017 -52286 40414
rect -52336 40005 -52286 40017
rect -52018 40414 -51968 40426
rect -52018 40017 -52012 40414
rect -51974 40017 -51968 40414
rect -52018 40005 -51968 40017
rect -51700 40414 -51650 40426
rect -51700 40017 -51694 40414
rect -51656 40017 -51650 40414
rect -51700 40005 -51650 40017
rect -51382 40414 -51332 40426
rect -51382 40017 -51376 40414
rect -51338 40017 -51332 40414
rect -51382 40005 -51332 40017
rect -51064 40414 -51014 40426
rect -51064 40017 -51058 40414
rect -51020 40017 -51014 40414
rect -51064 40005 -51014 40017
rect -50746 40414 -50696 40426
rect -50746 40017 -50740 40414
rect -50702 40017 -50696 40414
rect -50746 40005 -50696 40017
rect -50428 40414 -50378 40426
rect -50428 40017 -50422 40414
rect -50384 40017 -50378 40414
rect -50428 40005 -50378 40017
rect -50110 40414 -50060 40426
rect -50110 40017 -50104 40414
rect -50066 40017 -50060 40414
rect -50110 40005 -50060 40017
rect -49792 40414 -49742 40426
rect -49792 40017 -49786 40414
rect -49748 40017 -49742 40414
rect -49792 40005 -49742 40017
rect -49474 40414 -49424 40426
rect -49474 40017 -49468 40414
rect -49430 40017 -49424 40414
rect -49474 40005 -49424 40017
rect -49156 40414 -49106 40426
rect -49156 40017 -49150 40414
rect -49112 40017 -49106 40414
rect -49156 40005 -49106 40017
rect -48838 40414 -48788 40426
rect -48838 40017 -48832 40414
rect -48794 40017 -48788 40414
rect -48838 40005 -48788 40017
rect -48520 40414 -48470 40426
rect -48520 40017 -48514 40414
rect -48476 40017 -48470 40414
rect -48520 40005 -48470 40017
rect -48202 40414 -48152 40426
rect -48202 40017 -48196 40414
rect -48158 40017 -48152 40414
rect -48202 40005 -48152 40017
rect -47884 40414 -47834 40426
rect -47884 40017 -47878 40414
rect -47840 40017 -47834 40414
rect -47884 40005 -47834 40017
rect -47566 40414 -47516 40426
rect -47566 40017 -47560 40414
rect -47522 40017 -47516 40414
rect -47566 40005 -47516 40017
rect -47248 40414 -47198 40426
rect -47248 40017 -47242 40414
rect -47204 40017 -47198 40414
rect -47248 40005 -47198 40017
rect -46930 40414 -46880 40426
rect -46930 40017 -46924 40414
rect -46886 40017 -46880 40414
rect -46930 40005 -46880 40017
rect -46612 40414 -46562 40426
rect -46612 40017 -46606 40414
rect -46568 40017 -46562 40414
rect -46612 40005 -46562 40017
rect -46294 40414 -46244 40426
rect -46294 40017 -46288 40414
rect -46250 40017 -46244 40414
rect -46294 40005 -46244 40017
rect -45976 40414 -45926 40426
rect -45976 40017 -45970 40414
rect -45932 40017 -45926 40414
rect -45976 40005 -45926 40017
rect -45658 40414 -45608 40426
rect -45658 40017 -45652 40414
rect -45614 40017 -45608 40414
rect -45658 40005 -45608 40017
rect -45340 40414 -45290 40426
rect -45340 40017 -45334 40414
rect -45296 40017 -45290 40414
rect -45340 40005 -45290 40017
rect -45022 40414 -44972 40426
rect -45022 40017 -45016 40414
rect -44978 40017 -44972 40414
rect -45022 40005 -44972 40017
rect -44704 40414 -44654 40426
rect -44704 40017 -44698 40414
rect -44660 40017 -44654 40414
rect -44704 40005 -44654 40017
rect -44386 40414 -44336 40426
rect -44386 40017 -44380 40414
rect -44342 40017 -44336 40414
rect -44386 40005 -44336 40017
rect -44068 40414 -44018 40426
rect -44068 40017 -44062 40414
rect -44024 40017 -44018 40414
rect -44068 40005 -44018 40017
rect -43750 40414 -43700 40426
rect -43750 40017 -43744 40414
rect -43706 40017 -43700 40414
rect -43750 40005 -43700 40017
rect -43432 40414 -43382 40426
rect -43432 40017 -43426 40414
rect -43388 40017 -43382 40414
rect -43432 40005 -43382 40017
rect -43114 40414 -43064 40426
rect -43114 40017 -43108 40414
rect -43070 40017 -43064 40414
rect -43114 40005 -43064 40017
rect -42796 40414 -42746 40426
rect -42796 40017 -42790 40414
rect -42752 40017 -42746 40414
rect -42796 40005 -42746 40017
rect -42478 40414 -42428 40426
rect -42478 40017 -42472 40414
rect -42434 40017 -42428 40414
rect -42478 40005 -42428 40017
rect -42160 40414 -42110 40426
rect -42160 40017 -42154 40414
rect -42116 40017 -42110 40414
rect -42160 40005 -42110 40017
rect -41842 40414 -41792 40426
rect -41842 40017 -41836 40414
rect -41798 40017 -41792 40414
rect -41842 40005 -41792 40017
rect -41524 40414 -41474 40426
rect -41524 40017 -41518 40414
rect -41480 40017 -41474 40414
rect -41524 40005 -41474 40017
rect -41206 40414 -41156 40426
rect -41206 40017 -41200 40414
rect -41162 40017 -41156 40414
rect -41206 40005 -41156 40017
rect -40888 40414 -40838 40426
rect -40888 40017 -40882 40414
rect -40844 40017 -40838 40414
rect -40888 40005 -40838 40017
rect -40570 40414 -40520 40426
rect -40570 40017 -40564 40414
rect -40526 40017 -40520 40414
rect -40570 40005 -40520 40017
rect -40252 40414 -40202 40426
rect -40252 40017 -40246 40414
rect -40208 40017 -40202 40414
rect -40252 40005 -40202 40017
rect -39934 40414 -39884 40426
rect -39934 40017 -39928 40414
rect -39890 40017 -39884 40414
rect -39934 40005 -39884 40017
rect -39616 40414 -39566 40426
rect -39616 40017 -39610 40414
rect -39572 40017 -39566 40414
rect -39616 40005 -39566 40017
rect -39298 40414 -39248 40426
rect -39298 40017 -39292 40414
rect -39254 40017 -39248 40414
rect -39298 40005 -39248 40017
rect -38980 40414 -38930 40426
rect -38980 40017 -38974 40414
rect -38936 40017 -38930 40414
rect -38980 40005 -38930 40017
rect -38662 40414 -38612 40426
rect -38662 40017 -38656 40414
rect -38618 40017 -38612 40414
rect -38662 40005 -38612 40017
rect -38344 40414 -38294 40426
rect -38344 40017 -38338 40414
rect -38300 40017 -38294 40414
rect -38344 40005 -38294 40017
rect -38026 40414 -37976 40426
rect -38026 40017 -38020 40414
rect -37982 40017 -37976 40414
rect -38026 40005 -37976 40017
rect -37708 40414 -37658 40426
rect -37708 40017 -37702 40414
rect -37664 40017 -37658 40414
rect -37708 40005 -37658 40017
rect -37390 40414 -37340 40426
rect -37390 40017 -37384 40414
rect -37346 40017 -37340 40414
rect -37390 40005 -37340 40017
rect -37072 40414 -37022 40426
rect -37072 40017 -37066 40414
rect -37028 40017 -37022 40414
rect -37072 40005 -37022 40017
rect -36754 40414 -36704 40426
rect -36754 40017 -36748 40414
rect -36710 40017 -36704 40414
rect -36754 40005 -36704 40017
rect -36436 40414 -36386 40426
rect -36436 40017 -36430 40414
rect -36392 40017 -36386 40414
rect -36436 40005 -36386 40017
rect -36118 40414 -36068 40426
rect -36118 40017 -36112 40414
rect -36074 40017 -36068 40414
rect -36118 40005 -36068 40017
rect -35800 40414 -35750 40426
rect -35800 40017 -35794 40414
rect -35756 40017 -35750 40414
rect -35800 40005 -35750 40017
rect -35482 40414 -35432 40426
rect -35482 40017 -35476 40414
rect -35438 40017 -35432 40414
rect -35482 40005 -35432 40017
rect -35164 40414 -35114 40426
rect -35164 40017 -35158 40414
rect -35120 40017 -35114 40414
rect -35164 40005 -35114 40017
rect -34846 40414 -34796 40426
rect -34846 40017 -34840 40414
rect -34802 40017 -34796 40414
rect -34846 40005 -34796 40017
rect -34528 40414 -34478 40426
rect -34528 40017 -34522 40414
rect -34484 40017 -34478 40414
rect -34528 40005 -34478 40017
rect -34210 40414 -34160 40426
rect -34210 40017 -34204 40414
rect -34166 40017 -34160 40414
rect -34210 40005 -34160 40017
rect -33892 40414 -33842 40426
rect -33892 40017 -33886 40414
rect -33848 40017 -33842 40414
rect -33892 40005 -33842 40017
rect -33574 40414 -33524 40426
rect -33574 40017 -33568 40414
rect -33530 40017 -33524 40414
rect -33574 40005 -33524 40017
rect -33256 40414 -33206 40426
rect -33256 40017 -33250 40414
rect -33212 40017 -33206 40414
rect -33256 40005 -33206 40017
rect -32938 40414 -32888 40426
rect -32938 40017 -32932 40414
rect -32894 40017 -32888 40414
rect -32938 40005 -32888 40017
rect -32620 40414 -32570 40426
rect -32620 40017 -32614 40414
rect -32576 40017 -32570 40414
rect -32620 40005 -32570 40017
rect -32302 40414 -32252 40426
rect -32302 40017 -32296 40414
rect -32258 40017 -32252 40414
rect -32302 40005 -32252 40017
rect -31984 40414 -31934 40426
rect -31984 40017 -31978 40414
rect -31940 40017 -31934 40414
rect -31984 40005 -31934 40017
rect -31666 40414 -31616 40426
rect -31666 40017 -31660 40414
rect -31622 40017 -31616 40414
rect -31666 40005 -31616 40017
rect -31348 40414 -31298 40426
rect -31348 40017 -31342 40414
rect -31304 40017 -31298 40414
rect -31348 40005 -31298 40017
rect -31030 40414 -30980 40426
rect -31030 40017 -31024 40414
rect -30986 40017 -30980 40414
rect -31030 40005 -30980 40017
rect -30712 40414 -30662 40426
rect -30712 40017 -30706 40414
rect -30668 40017 -30662 40414
rect -30712 40005 -30662 40017
rect -30394 40414 -30344 40426
rect -30394 40017 -30388 40414
rect -30350 40017 -30344 40414
rect -30394 40005 -30344 40017
rect -30076 40414 -30026 40426
rect -30076 40017 -30070 40414
rect -30032 40017 -30026 40414
rect -30076 40005 -30026 40017
rect -29758 40414 -29708 40426
rect -29758 40017 -29752 40414
rect -29714 40017 -29708 40414
rect -29758 40005 -29708 40017
rect -29440 40414 -29390 40426
rect -29440 40017 -29434 40414
rect -29396 40017 -29390 40414
rect -29440 40005 -29390 40017
rect -29122 40414 -29072 40426
rect -29122 40017 -29116 40414
rect -29078 40017 -29072 40414
rect -29122 40005 -29072 40017
rect -28804 40414 -28754 40426
rect -28804 40017 -28798 40414
rect -28760 40017 -28754 40414
rect -28804 40005 -28754 40017
rect -28486 40414 -28436 40426
rect -28486 40017 -28480 40414
rect -28442 40017 -28436 40414
rect -28486 40005 -28436 40017
rect -28168 40414 -28118 40426
rect -28168 40017 -28162 40414
rect -28124 40017 -28118 40414
rect -28168 40005 -28118 40017
rect -27850 40414 -27800 40426
rect -27850 40017 -27844 40414
rect -27806 40017 -27800 40414
rect -27850 40005 -27800 40017
rect -27532 40414 -27482 40426
rect -27532 40017 -27526 40414
rect -27488 40017 -27482 40414
rect -27532 40005 -27482 40017
rect -27214 40414 -27164 40426
rect -27214 40017 -27208 40414
rect -27170 40017 -27164 40414
rect -27214 40005 -27164 40017
rect -26896 40414 -26846 40426
rect -26896 40017 -26890 40414
rect -26852 40017 -26846 40414
rect -26896 40005 -26846 40017
rect -26578 40414 -26528 40426
rect -26578 40017 -26572 40414
rect -26534 40017 -26528 40414
rect -26578 40005 -26528 40017
rect -26260 40414 -26210 40426
rect -26260 40017 -26254 40414
rect -26216 40017 -26210 40414
rect -26260 40005 -26210 40017
rect -25942 40414 -25892 40426
rect -25942 40017 -25936 40414
rect -25898 40017 -25892 40414
rect -25942 40005 -25892 40017
rect -25624 40414 -25574 40426
rect -25624 40017 -25618 40414
rect -25580 40017 -25574 40414
rect -25624 40005 -25574 40017
rect -25306 40414 -25256 40426
rect -25306 40017 -25300 40414
rect -25262 40017 -25256 40414
rect -25306 40005 -25256 40017
rect -24988 40414 -24938 40426
rect -24988 40017 -24982 40414
rect -24944 40017 -24938 40414
rect -24988 40005 -24938 40017
rect -24670 40414 -24620 40426
rect -24670 40017 -24664 40414
rect -24626 40017 -24620 40414
rect -24670 40005 -24620 40017
rect -24352 40414 -24302 40426
rect -24352 40017 -24346 40414
rect -24308 40017 -24302 40414
rect -24352 40005 -24302 40017
rect -24034 40414 -23984 40426
rect -24034 40017 -24028 40414
rect -23990 40017 -23984 40414
rect -24034 40005 -23984 40017
rect -23716 40414 -23666 40426
rect -23716 40017 -23710 40414
rect -23672 40017 -23666 40414
rect -23716 40005 -23666 40017
rect -23398 40414 -23348 40426
rect -23398 40017 -23392 40414
rect -23354 40017 -23348 40414
rect -23398 40005 -23348 40017
rect -23080 40414 -23030 40426
rect -23080 40017 -23074 40414
rect -23036 40017 -23030 40414
rect -23080 40005 -23030 40017
rect -22762 40414 -22712 40426
rect -22762 40017 -22756 40414
rect -22718 40017 -22712 40414
rect -22762 40005 -22712 40017
rect -22444 40414 -22394 40426
rect -22444 40017 -22438 40414
rect -22400 40017 -22394 40414
rect -22444 40005 -22394 40017
rect -22126 40414 -22076 40426
rect -22126 40017 -22120 40414
rect -22082 40017 -22076 40414
rect -22126 40005 -22076 40017
rect -21808 40414 -21758 40426
rect -21808 40017 -21802 40414
rect -21764 40017 -21758 40414
rect -21808 40005 -21758 40017
rect -21490 40414 -21440 40426
rect -21490 40017 -21484 40414
rect -21446 40017 -21440 40414
rect -21490 40005 -21440 40017
rect -21172 40414 -21122 40426
rect -21172 40017 -21166 40414
rect -21128 40017 -21122 40414
rect -21172 40005 -21122 40017
rect -20854 40414 -20804 40426
rect -20854 40017 -20848 40414
rect -20810 40017 -20804 40414
rect -20854 40005 -20804 40017
rect -20536 40414 -20486 40426
rect -20536 40017 -20530 40414
rect -20492 40017 -20486 40414
rect -20536 40005 -20486 40017
rect -20218 40414 -20168 40426
rect -20218 40017 -20212 40414
rect -20174 40017 -20168 40414
rect -20218 40005 -20168 40017
rect -19900 40414 -19850 40426
rect -19900 40017 -19894 40414
rect -19856 40017 -19850 40414
rect -19900 40005 -19850 40017
rect -19582 40414 -19532 40426
rect -19582 40017 -19576 40414
rect -19538 40017 -19532 40414
rect -19582 40005 -19532 40017
rect -19264 40414 -19214 40426
rect -19264 40017 -19258 40414
rect -19220 40017 -19214 40414
rect -19264 40005 -19214 40017
rect -18946 40414 -18896 40426
rect -18946 40017 -18940 40414
rect -18902 40017 -18896 40414
rect -18946 40005 -18896 40017
rect -18628 40414 -18578 40426
rect -18628 40017 -18622 40414
rect -18584 40017 -18578 40414
rect -18628 40005 -18578 40017
rect -18310 40414 -18260 40426
rect -18310 40017 -18304 40414
rect -18266 40017 -18260 40414
rect -18310 40005 -18260 40017
rect -17992 40414 -17942 40426
rect -17992 40017 -17986 40414
rect -17948 40017 -17942 40414
rect -17992 40005 -17942 40017
rect -17674 40414 -17624 40426
rect -17674 40017 -17668 40414
rect -17630 40017 -17624 40414
rect -17674 40005 -17624 40017
rect -17356 40414 -17306 40426
rect -17356 40017 -17350 40414
rect -17312 40017 -17306 40414
rect -17356 40005 -17306 40017
rect -17038 40414 -16988 40426
rect -17038 40017 -17032 40414
rect -16994 40017 -16988 40414
rect -17038 40005 -16988 40017
rect -16720 40414 -16670 40426
rect -16720 40017 -16714 40414
rect -16676 40017 -16670 40414
rect -16720 40005 -16670 40017
rect -16402 40414 -16352 40426
rect -16402 40017 -16396 40414
rect -16358 40017 -16352 40414
rect -16402 40005 -16352 40017
rect -16084 40414 -16034 40426
rect -16084 40017 -16078 40414
rect -16040 40017 -16034 40414
rect -16084 40005 -16034 40017
rect -15766 40414 -15716 40426
rect -15766 40017 -15760 40414
rect -15722 40017 -15716 40414
rect -15766 40005 -15716 40017
rect -15448 40414 -15398 40426
rect -15448 40017 -15442 40414
rect -15404 40017 -15398 40414
rect -15448 40005 -15398 40017
rect -15130 40414 -15080 40426
rect -15130 40017 -15124 40414
rect -15086 40017 -15080 40414
rect -15130 40005 -15080 40017
rect -14812 40414 -14762 40426
rect -14812 40017 -14806 40414
rect -14768 40017 -14762 40414
rect -14812 40005 -14762 40017
rect -14494 40414 -14444 40426
rect -14494 40017 -14488 40414
rect -14450 40017 -14444 40414
rect -14494 40005 -14444 40017
rect -14176 40414 -14126 40426
rect -14176 40017 -14170 40414
rect -14132 40017 -14126 40414
rect -14176 40005 -14126 40017
rect -13858 40414 -13808 40426
rect -13858 40017 -13852 40414
rect -13814 40017 -13808 40414
rect -13858 40005 -13808 40017
rect -13540 40414 -13490 40426
rect -13540 40017 -13534 40414
rect -13496 40017 -13490 40414
rect -13540 40005 -13490 40017
rect -13222 40414 -13172 40426
rect -13222 40017 -13216 40414
rect -13178 40017 -13172 40414
rect -13222 40005 -13172 40017
rect -12904 40414 -12854 40426
rect -12904 40017 -12898 40414
rect -12860 40017 -12854 40414
rect -12904 40005 -12854 40017
rect -12586 40414 -12536 40426
rect -12586 40017 -12580 40414
rect -12542 40017 -12536 40414
rect -12586 40005 -12536 40017
rect -12268 40414 -12218 40426
rect -12268 40017 -12262 40414
rect -12224 40017 -12218 40414
rect -12268 40005 -12218 40017
rect -11950 40414 -11900 40426
rect -11950 40017 -11944 40414
rect -11906 40017 -11900 40414
rect -11950 40005 -11900 40017
rect -11632 40414 -11582 40426
rect -11632 40017 -11626 40414
rect -11588 40017 -11582 40414
rect -11632 40005 -11582 40017
rect -11314 40414 -11264 40426
rect -11314 40017 -11308 40414
rect -11270 40017 -11264 40414
rect -11314 40005 -11264 40017
rect -10996 40414 -10946 40426
rect -10996 40017 -10990 40414
rect -10952 40017 -10946 40414
rect -10996 40005 -10946 40017
rect -10678 40414 -10628 40426
rect -10678 40017 -10672 40414
rect -10634 40017 -10628 40414
rect -10678 40005 -10628 40017
rect -10360 40414 -10310 40426
rect -10360 40017 -10354 40414
rect -10316 40017 -10310 40414
rect -10360 40005 -10310 40017
rect -10042 40414 -9992 40426
rect -10042 40017 -10036 40414
rect -9998 40017 -9992 40414
rect -10042 40005 -9992 40017
rect -9724 40414 -9674 40426
rect -9724 40017 -9718 40414
rect -9680 40017 -9674 40414
rect -9724 40005 -9674 40017
rect -9406 40414 -9356 40426
rect -9406 40017 -9400 40414
rect -9362 40017 -9356 40414
rect -9406 40005 -9356 40017
rect -9088 40414 -9038 40426
rect -9088 40017 -9082 40414
rect -9044 40017 -9038 40414
rect -9088 40005 -9038 40017
rect -8770 40414 -8720 40426
rect -8770 40017 -8764 40414
rect -8726 40017 -8720 40414
rect -8770 40005 -8720 40017
rect -8452 40414 -8402 40426
rect -8452 40017 -8446 40414
rect -8408 40017 -8402 40414
rect -8452 40005 -8402 40017
rect -8134 40414 -8084 40426
rect -8134 40017 -8128 40414
rect -8090 40017 -8084 40414
rect -8134 40005 -8084 40017
rect -7816 40414 -7766 40426
rect -7816 40017 -7810 40414
rect -7772 40017 -7766 40414
rect -7816 40005 -7766 40017
rect -7498 40414 -7448 40426
rect -7498 40017 -7492 40414
rect -7454 40017 -7448 40414
rect -7498 40005 -7448 40017
rect -7180 40414 -7130 40426
rect -7180 40017 -7174 40414
rect -7136 40017 -7130 40414
rect -7180 40005 -7130 40017
rect -6862 40414 -6812 40426
rect -6862 40017 -6856 40414
rect -6818 40017 -6812 40414
rect -6862 40005 -6812 40017
rect -6544 40414 -6494 40426
rect -6544 40017 -6538 40414
rect -6500 40017 -6494 40414
rect -6544 40005 -6494 40017
rect -6226 40414 -6176 40426
rect -6226 40017 -6220 40414
rect -6182 40017 -6176 40414
rect -6226 40005 -6176 40017
rect -5908 40414 -5858 40426
rect -5908 40017 -5902 40414
rect -5864 40017 -5858 40414
rect -5908 40005 -5858 40017
rect -5590 40414 -5540 40426
rect -5590 40017 -5584 40414
rect -5546 40017 -5540 40414
rect -5590 40005 -5540 40017
rect -5272 40414 -5222 40426
rect -5272 40017 -5266 40414
rect -5228 40017 -5222 40414
rect -5272 40005 -5222 40017
rect -4954 40414 -4904 40426
rect -4954 40017 -4948 40414
rect -4910 40017 -4904 40414
rect -4954 40005 -4904 40017
rect -4636 40414 -4586 40426
rect -4636 40017 -4630 40414
rect -4592 40017 -4586 40414
rect -4636 40005 -4586 40017
rect -4318 40414 -4268 40426
rect -4318 40017 -4312 40414
rect -4274 40017 -4268 40414
rect -4318 40005 -4268 40017
rect -4000 40414 -3950 40426
rect -4000 40017 -3994 40414
rect -3956 40017 -3950 40414
rect -4000 40005 -3950 40017
rect -3682 40414 -3632 40426
rect -3682 40017 -3676 40414
rect -3638 40017 -3632 40414
rect -3682 40005 -3632 40017
rect -3364 40414 -3314 40426
rect -3364 40017 -3358 40414
rect -3320 40017 -3314 40414
rect -3364 40005 -3314 40017
rect -3046 40414 -2996 40426
rect -3046 40017 -3040 40414
rect -3002 40017 -2996 40414
rect -3046 40005 -2996 40017
rect -2728 40414 -2678 40426
rect -2728 40017 -2722 40414
rect -2684 40017 -2678 40414
rect -2728 40005 -2678 40017
rect -2410 40414 -2360 40426
rect -2410 40017 -2404 40414
rect -2366 40017 -2360 40414
rect -2410 40005 -2360 40017
rect -2092 40414 -2042 40426
rect -2092 40017 -2086 40414
rect -2048 40017 -2042 40414
rect -2092 40005 -2042 40017
rect -1774 40414 -1724 40426
rect -1774 40017 -1768 40414
rect -1730 40017 -1724 40414
rect -1774 40005 -1724 40017
rect -1456 40414 -1406 40426
rect -1456 40017 -1450 40414
rect -1412 40017 -1406 40414
rect -1456 40005 -1406 40017
rect -1138 40414 -1088 40426
rect -1138 40017 -1132 40414
rect -1094 40017 -1088 40414
rect -1138 40005 -1088 40017
rect -820 40414 -770 40426
rect -820 40017 -814 40414
rect -776 40017 -770 40414
rect -820 40005 -770 40017
rect -502 40414 -452 40426
rect -502 40017 -496 40414
rect -458 40017 -452 40414
rect -502 40005 -452 40017
rect -184 40414 -134 40426
rect -184 40017 -178 40414
rect -140 40017 -134 40414
rect -184 40005 -134 40017
rect 134 40414 184 40426
rect 134 40017 140 40414
rect 178 40017 184 40414
rect 134 40005 184 40017
rect 452 40414 502 40426
rect 452 40017 458 40414
rect 496 40017 502 40414
rect 452 40005 502 40017
rect 770 40414 820 40426
rect 770 40017 776 40414
rect 814 40017 820 40414
rect 770 40005 820 40017
rect 1088 40414 1138 40426
rect 1088 40017 1094 40414
rect 1132 40017 1138 40414
rect 1088 40005 1138 40017
rect 1406 40414 1456 40426
rect 1406 40017 1412 40414
rect 1450 40017 1456 40414
rect 1406 40005 1456 40017
rect 1724 40414 1774 40426
rect 1724 40017 1730 40414
rect 1768 40017 1774 40414
rect 1724 40005 1774 40017
rect 2042 40414 2092 40426
rect 2042 40017 2048 40414
rect 2086 40017 2092 40414
rect 2042 40005 2092 40017
rect 2360 40414 2410 40426
rect 2360 40017 2366 40414
rect 2404 40017 2410 40414
rect 2360 40005 2410 40017
rect 2678 40414 2728 40426
rect 2678 40017 2684 40414
rect 2722 40017 2728 40414
rect 2678 40005 2728 40017
rect 2996 40414 3046 40426
rect 2996 40017 3002 40414
rect 3040 40017 3046 40414
rect 2996 40005 3046 40017
rect 3314 40414 3364 40426
rect 3314 40017 3320 40414
rect 3358 40017 3364 40414
rect 3314 40005 3364 40017
rect 3632 40414 3682 40426
rect 3632 40017 3638 40414
rect 3676 40017 3682 40414
rect 3632 40005 3682 40017
rect 3950 40414 4000 40426
rect 3950 40017 3956 40414
rect 3994 40017 4000 40414
rect 3950 40005 4000 40017
rect 4268 40414 4318 40426
rect 4268 40017 4274 40414
rect 4312 40017 4318 40414
rect 4268 40005 4318 40017
rect 4586 40414 4636 40426
rect 4586 40017 4592 40414
rect 4630 40017 4636 40414
rect 4586 40005 4636 40017
rect 4904 40414 4954 40426
rect 4904 40017 4910 40414
rect 4948 40017 4954 40414
rect 4904 40005 4954 40017
rect 5222 40414 5272 40426
rect 5222 40017 5228 40414
rect 5266 40017 5272 40414
rect 5222 40005 5272 40017
rect 5540 40414 5590 40426
rect 5540 40017 5546 40414
rect 5584 40017 5590 40414
rect 5540 40005 5590 40017
rect 5858 40414 5908 40426
rect 5858 40017 5864 40414
rect 5902 40017 5908 40414
rect 5858 40005 5908 40017
rect 6176 40414 6226 40426
rect 6176 40017 6182 40414
rect 6220 40017 6226 40414
rect 6176 40005 6226 40017
rect 6494 40414 6544 40426
rect 6494 40017 6500 40414
rect 6538 40017 6544 40414
rect 6494 40005 6544 40017
rect 6812 40414 6862 40426
rect 6812 40017 6818 40414
rect 6856 40017 6862 40414
rect 6812 40005 6862 40017
rect 7130 40414 7180 40426
rect 7130 40017 7136 40414
rect 7174 40017 7180 40414
rect 7130 40005 7180 40017
rect 7448 40414 7498 40426
rect 7448 40017 7454 40414
rect 7492 40017 7498 40414
rect 7448 40005 7498 40017
rect 7766 40414 7816 40426
rect 7766 40017 7772 40414
rect 7810 40017 7816 40414
rect 7766 40005 7816 40017
rect 8084 40414 8134 40426
rect 8084 40017 8090 40414
rect 8128 40017 8134 40414
rect 8084 40005 8134 40017
rect 8402 40414 8452 40426
rect 8402 40017 8408 40414
rect 8446 40017 8452 40414
rect 8402 40005 8452 40017
rect 8720 40414 8770 40426
rect 8720 40017 8726 40414
rect 8764 40017 8770 40414
rect 8720 40005 8770 40017
rect 9038 40414 9088 40426
rect 9038 40017 9044 40414
rect 9082 40017 9088 40414
rect 9038 40005 9088 40017
rect 9356 40414 9406 40426
rect 9356 40017 9362 40414
rect 9400 40017 9406 40414
rect 9356 40005 9406 40017
rect 9674 40414 9724 40426
rect 9674 40017 9680 40414
rect 9718 40017 9724 40414
rect 9674 40005 9724 40017
rect 9992 40414 10042 40426
rect 9992 40017 9998 40414
rect 10036 40017 10042 40414
rect 9992 40005 10042 40017
rect 10310 40414 10360 40426
rect 10310 40017 10316 40414
rect 10354 40017 10360 40414
rect 10310 40005 10360 40017
rect 10628 40414 10678 40426
rect 10628 40017 10634 40414
rect 10672 40017 10678 40414
rect 10628 40005 10678 40017
rect 10946 40414 10996 40426
rect 10946 40017 10952 40414
rect 10990 40017 10996 40414
rect 10946 40005 10996 40017
rect 11264 40414 11314 40426
rect 11264 40017 11270 40414
rect 11308 40017 11314 40414
rect 11264 40005 11314 40017
rect 11582 40414 11632 40426
rect 11582 40017 11588 40414
rect 11626 40017 11632 40414
rect 11582 40005 11632 40017
rect 11900 40414 11950 40426
rect 11900 40017 11906 40414
rect 11944 40017 11950 40414
rect 11900 40005 11950 40017
rect 12218 40414 12268 40426
rect 12218 40017 12224 40414
rect 12262 40017 12268 40414
rect 12218 40005 12268 40017
rect 12536 40414 12586 40426
rect 12536 40017 12542 40414
rect 12580 40017 12586 40414
rect 12536 40005 12586 40017
rect 12854 40414 12904 40426
rect 12854 40017 12860 40414
rect 12898 40017 12904 40414
rect 12854 40005 12904 40017
rect 13172 40414 13222 40426
rect 13172 40017 13178 40414
rect 13216 40017 13222 40414
rect 13172 40005 13222 40017
rect 13490 40414 13540 40426
rect 13490 40017 13496 40414
rect 13534 40017 13540 40414
rect 13490 40005 13540 40017
rect 13808 40414 13858 40426
rect 13808 40017 13814 40414
rect 13852 40017 13858 40414
rect 13808 40005 13858 40017
rect 14126 40414 14176 40426
rect 14126 40017 14132 40414
rect 14170 40017 14176 40414
rect 14126 40005 14176 40017
rect 14444 40414 14494 40426
rect 14444 40017 14450 40414
rect 14488 40017 14494 40414
rect 14444 40005 14494 40017
rect 14762 40414 14812 40426
rect 14762 40017 14768 40414
rect 14806 40017 14812 40414
rect 14762 40005 14812 40017
rect 15080 40414 15130 40426
rect 15080 40017 15086 40414
rect 15124 40017 15130 40414
rect 15080 40005 15130 40017
rect 15398 40414 15448 40426
rect 15398 40017 15404 40414
rect 15442 40017 15448 40414
rect 15398 40005 15448 40017
rect 15716 40414 15766 40426
rect 15716 40017 15722 40414
rect 15760 40017 15766 40414
rect 15716 40005 15766 40017
rect 16034 40414 16084 40426
rect 16034 40017 16040 40414
rect 16078 40017 16084 40414
rect 16034 40005 16084 40017
rect 16352 40414 16402 40426
rect 16352 40017 16358 40414
rect 16396 40017 16402 40414
rect 16352 40005 16402 40017
rect 16670 40414 16720 40426
rect 16670 40017 16676 40414
rect 16714 40017 16720 40414
rect 16670 40005 16720 40017
rect 16988 40414 17038 40426
rect 16988 40017 16994 40414
rect 17032 40017 17038 40414
rect 16988 40005 17038 40017
rect 17306 40414 17356 40426
rect 17306 40017 17312 40414
rect 17350 40017 17356 40414
rect 17306 40005 17356 40017
rect 17624 40414 17674 40426
rect 17624 40017 17630 40414
rect 17668 40017 17674 40414
rect 17624 40005 17674 40017
rect 17942 40414 17992 40426
rect 17942 40017 17948 40414
rect 17986 40017 17992 40414
rect 17942 40005 17992 40017
rect 18260 40414 18310 40426
rect 18260 40017 18266 40414
rect 18304 40017 18310 40414
rect 18260 40005 18310 40017
rect 18578 40414 18628 40426
rect 18578 40017 18584 40414
rect 18622 40017 18628 40414
rect 18578 40005 18628 40017
rect 18896 40414 18946 40426
rect 18896 40017 18902 40414
rect 18940 40017 18946 40414
rect 18896 40005 18946 40017
rect 19214 40414 19264 40426
rect 19214 40017 19220 40414
rect 19258 40017 19264 40414
rect 19214 40005 19264 40017
rect 19532 40414 19582 40426
rect 19532 40017 19538 40414
rect 19576 40017 19582 40414
rect 19532 40005 19582 40017
rect 19850 40414 19900 40426
rect 19850 40017 19856 40414
rect 19894 40017 19900 40414
rect 19850 40005 19900 40017
rect 20168 40414 20218 40426
rect 20168 40017 20174 40414
rect 20212 40017 20218 40414
rect 20168 40005 20218 40017
rect 20486 40414 20536 40426
rect 20486 40017 20492 40414
rect 20530 40017 20536 40414
rect 20486 40005 20536 40017
rect 20804 40414 20854 40426
rect 20804 40017 20810 40414
rect 20848 40017 20854 40414
rect 20804 40005 20854 40017
rect 21122 40414 21172 40426
rect 21122 40017 21128 40414
rect 21166 40017 21172 40414
rect 21122 40005 21172 40017
rect 21440 40414 21490 40426
rect 21440 40017 21446 40414
rect 21484 40017 21490 40414
rect 21440 40005 21490 40017
rect 21758 40414 21808 40426
rect 21758 40017 21764 40414
rect 21802 40017 21808 40414
rect 21758 40005 21808 40017
rect 22076 40414 22126 40426
rect 22076 40017 22082 40414
rect 22120 40017 22126 40414
rect 22076 40005 22126 40017
rect 22394 40414 22444 40426
rect 22394 40017 22400 40414
rect 22438 40017 22444 40414
rect 22394 40005 22444 40017
rect 22712 40414 22762 40426
rect 22712 40017 22718 40414
rect 22756 40017 22762 40414
rect 22712 40005 22762 40017
rect 23030 40414 23080 40426
rect 23030 40017 23036 40414
rect 23074 40017 23080 40414
rect 23030 40005 23080 40017
rect 23348 40414 23398 40426
rect 23348 40017 23354 40414
rect 23392 40017 23398 40414
rect 23348 40005 23398 40017
rect 23666 40414 23716 40426
rect 23666 40017 23672 40414
rect 23710 40017 23716 40414
rect 23666 40005 23716 40017
rect 23984 40414 24034 40426
rect 23984 40017 23990 40414
rect 24028 40017 24034 40414
rect 23984 40005 24034 40017
rect 24302 40414 24352 40426
rect 24302 40017 24308 40414
rect 24346 40017 24352 40414
rect 24302 40005 24352 40017
rect 24620 40414 24670 40426
rect 24620 40017 24626 40414
rect 24664 40017 24670 40414
rect 24620 40005 24670 40017
rect 24938 40414 24988 40426
rect 24938 40017 24944 40414
rect 24982 40017 24988 40414
rect 24938 40005 24988 40017
rect 25256 40414 25306 40426
rect 25256 40017 25262 40414
rect 25300 40017 25306 40414
rect 25256 40005 25306 40017
rect 25574 40414 25624 40426
rect 25574 40017 25580 40414
rect 25618 40017 25624 40414
rect 25574 40005 25624 40017
rect 25892 40414 25942 40426
rect 25892 40017 25898 40414
rect 25936 40017 25942 40414
rect 25892 40005 25942 40017
rect 26210 40414 26260 40426
rect 26210 40017 26216 40414
rect 26254 40017 26260 40414
rect 26210 40005 26260 40017
rect 26528 40414 26578 40426
rect 26528 40017 26534 40414
rect 26572 40017 26578 40414
rect 26528 40005 26578 40017
rect 26846 40414 26896 40426
rect 26846 40017 26852 40414
rect 26890 40017 26896 40414
rect 26846 40005 26896 40017
rect 27164 40414 27214 40426
rect 27164 40017 27170 40414
rect 27208 40017 27214 40414
rect 27164 40005 27214 40017
rect 27482 40414 27532 40426
rect 27482 40017 27488 40414
rect 27526 40017 27532 40414
rect 27482 40005 27532 40017
rect 27800 40414 27850 40426
rect 27800 40017 27806 40414
rect 27844 40017 27850 40414
rect 27800 40005 27850 40017
rect 28118 40414 28168 40426
rect 28118 40017 28124 40414
rect 28162 40017 28168 40414
rect 28118 40005 28168 40017
rect 28436 40414 28486 40426
rect 28436 40017 28442 40414
rect 28480 40017 28486 40414
rect 28436 40005 28486 40017
rect 28754 40414 28804 40426
rect 28754 40017 28760 40414
rect 28798 40017 28804 40414
rect 28754 40005 28804 40017
rect 29072 40414 29122 40426
rect 29072 40017 29078 40414
rect 29116 40017 29122 40414
rect 29072 40005 29122 40017
rect 29390 40414 29440 40426
rect 29390 40017 29396 40414
rect 29434 40017 29440 40414
rect 29390 40005 29440 40017
rect 29708 40414 29758 40426
rect 29708 40017 29714 40414
rect 29752 40017 29758 40414
rect 29708 40005 29758 40017
rect 30026 40414 30076 40426
rect 30026 40017 30032 40414
rect 30070 40017 30076 40414
rect 30026 40005 30076 40017
rect 30344 40414 30394 40426
rect 30344 40017 30350 40414
rect 30388 40017 30394 40414
rect 30344 40005 30394 40017
rect 30662 40414 30712 40426
rect 30662 40017 30668 40414
rect 30706 40017 30712 40414
rect 30662 40005 30712 40017
rect 30980 40414 31030 40426
rect 30980 40017 30986 40414
rect 31024 40017 31030 40414
rect 30980 40005 31030 40017
rect 31298 40414 31348 40426
rect 31298 40017 31304 40414
rect 31342 40017 31348 40414
rect 31298 40005 31348 40017
rect 31616 40414 31666 40426
rect 31616 40017 31622 40414
rect 31660 40017 31666 40414
rect 31616 40005 31666 40017
rect 31934 40414 31984 40426
rect 31934 40017 31940 40414
rect 31978 40017 31984 40414
rect 31934 40005 31984 40017
rect 32252 40414 32302 40426
rect 32252 40017 32258 40414
rect 32296 40017 32302 40414
rect 32252 40005 32302 40017
rect 32570 40414 32620 40426
rect 32570 40017 32576 40414
rect 32614 40017 32620 40414
rect 32570 40005 32620 40017
rect 32888 40414 32938 40426
rect 32888 40017 32894 40414
rect 32932 40017 32938 40414
rect 32888 40005 32938 40017
rect 33206 40414 33256 40426
rect 33206 40017 33212 40414
rect 33250 40017 33256 40414
rect 33206 40005 33256 40017
rect 33524 40414 33574 40426
rect 33524 40017 33530 40414
rect 33568 40017 33574 40414
rect 33524 40005 33574 40017
rect 33842 40414 33892 40426
rect 33842 40017 33848 40414
rect 33886 40017 33892 40414
rect 33842 40005 33892 40017
rect 34160 40414 34210 40426
rect 34160 40017 34166 40414
rect 34204 40017 34210 40414
rect 34160 40005 34210 40017
rect 34478 40414 34528 40426
rect 34478 40017 34484 40414
rect 34522 40017 34528 40414
rect 34478 40005 34528 40017
rect 34796 40414 34846 40426
rect 34796 40017 34802 40414
rect 34840 40017 34846 40414
rect 34796 40005 34846 40017
rect 35114 40414 35164 40426
rect 35114 40017 35120 40414
rect 35158 40017 35164 40414
rect 35114 40005 35164 40017
rect 35432 40414 35482 40426
rect 35432 40017 35438 40414
rect 35476 40017 35482 40414
rect 35432 40005 35482 40017
rect 35750 40414 35800 40426
rect 35750 40017 35756 40414
rect 35794 40017 35800 40414
rect 35750 40005 35800 40017
rect 36068 40414 36118 40426
rect 36068 40017 36074 40414
rect 36112 40017 36118 40414
rect 36068 40005 36118 40017
rect 36386 40414 36436 40426
rect 36386 40017 36392 40414
rect 36430 40017 36436 40414
rect 36386 40005 36436 40017
rect 36704 40414 36754 40426
rect 36704 40017 36710 40414
rect 36748 40017 36754 40414
rect 36704 40005 36754 40017
rect 37022 40414 37072 40426
rect 37022 40017 37028 40414
rect 37066 40017 37072 40414
rect 37022 40005 37072 40017
rect 37340 40414 37390 40426
rect 37340 40017 37346 40414
rect 37384 40017 37390 40414
rect 37340 40005 37390 40017
rect 37658 40414 37708 40426
rect 37658 40017 37664 40414
rect 37702 40017 37708 40414
rect 37658 40005 37708 40017
rect 37976 40414 38026 40426
rect 37976 40017 37982 40414
rect 38020 40017 38026 40414
rect 37976 40005 38026 40017
rect 38294 40414 38344 40426
rect 38294 40017 38300 40414
rect 38338 40017 38344 40414
rect 38294 40005 38344 40017
rect 38612 40414 38662 40426
rect 38612 40017 38618 40414
rect 38656 40017 38662 40414
rect 38612 40005 38662 40017
rect 38930 40414 38980 40426
rect 38930 40017 38936 40414
rect 38974 40017 38980 40414
rect 38930 40005 38980 40017
rect 39248 40414 39298 40426
rect 39248 40017 39254 40414
rect 39292 40017 39298 40414
rect 39248 40005 39298 40017
rect 39566 40414 39616 40426
rect 39566 40017 39572 40414
rect 39610 40017 39616 40414
rect 39566 40005 39616 40017
rect 39884 40414 39934 40426
rect 39884 40017 39890 40414
rect 39928 40017 39934 40414
rect 39884 40005 39934 40017
rect 40202 40414 40252 40426
rect 40202 40017 40208 40414
rect 40246 40017 40252 40414
rect 40202 40005 40252 40017
rect 40520 40414 40570 40426
rect 40520 40017 40526 40414
rect 40564 40017 40570 40414
rect 40520 40005 40570 40017
rect 40838 40414 40888 40426
rect 40838 40017 40844 40414
rect 40882 40017 40888 40414
rect 40838 40005 40888 40017
rect 41156 40414 41206 40426
rect 41156 40017 41162 40414
rect 41200 40017 41206 40414
rect 41156 40005 41206 40017
rect 41474 40414 41524 40426
rect 41474 40017 41480 40414
rect 41518 40017 41524 40414
rect 41474 40005 41524 40017
rect 41792 40414 41842 40426
rect 41792 40017 41798 40414
rect 41836 40017 41842 40414
rect 41792 40005 41842 40017
rect 42110 40414 42160 40426
rect 42110 40017 42116 40414
rect 42154 40017 42160 40414
rect 42110 40005 42160 40017
rect 42428 40414 42478 40426
rect 42428 40017 42434 40414
rect 42472 40017 42478 40414
rect 42428 40005 42478 40017
rect 42746 40414 42796 40426
rect 42746 40017 42752 40414
rect 42790 40017 42796 40414
rect 42746 40005 42796 40017
rect 43064 40414 43114 40426
rect 43064 40017 43070 40414
rect 43108 40017 43114 40414
rect 43064 40005 43114 40017
rect 43382 40414 43432 40426
rect 43382 40017 43388 40414
rect 43426 40017 43432 40414
rect 43382 40005 43432 40017
rect 43700 40414 43750 40426
rect 43700 40017 43706 40414
rect 43744 40017 43750 40414
rect 43700 40005 43750 40017
rect 44018 40414 44068 40426
rect 44018 40017 44024 40414
rect 44062 40017 44068 40414
rect 44018 40005 44068 40017
rect 44336 40414 44386 40426
rect 44336 40017 44342 40414
rect 44380 40017 44386 40414
rect 44336 40005 44386 40017
rect 44654 40414 44704 40426
rect 44654 40017 44660 40414
rect 44698 40017 44704 40414
rect 44654 40005 44704 40017
rect 44972 40414 45022 40426
rect 44972 40017 44978 40414
rect 45016 40017 45022 40414
rect 44972 40005 45022 40017
rect 45290 40414 45340 40426
rect 45290 40017 45296 40414
rect 45334 40017 45340 40414
rect 45290 40005 45340 40017
rect 45608 40414 45658 40426
rect 45608 40017 45614 40414
rect 45652 40017 45658 40414
rect 45608 40005 45658 40017
rect 45926 40414 45976 40426
rect 45926 40017 45932 40414
rect 45970 40017 45976 40414
rect 45926 40005 45976 40017
rect 46244 40414 46294 40426
rect 46244 40017 46250 40414
rect 46288 40017 46294 40414
rect 46244 40005 46294 40017
rect 46562 40414 46612 40426
rect 46562 40017 46568 40414
rect 46606 40017 46612 40414
rect 46562 40005 46612 40017
rect 46880 40414 46930 40426
rect 46880 40017 46886 40414
rect 46924 40017 46930 40414
rect 46880 40005 46930 40017
rect 47198 40414 47248 40426
rect 47198 40017 47204 40414
rect 47242 40017 47248 40414
rect 47198 40005 47248 40017
rect 47516 40414 47566 40426
rect 47516 40017 47522 40414
rect 47560 40017 47566 40414
rect 47516 40005 47566 40017
rect 47834 40414 47884 40426
rect 47834 40017 47840 40414
rect 47878 40017 47884 40414
rect 47834 40005 47884 40017
rect 48152 40414 48202 40426
rect 48152 40017 48158 40414
rect 48196 40017 48202 40414
rect 48152 40005 48202 40017
rect 48470 40414 48520 40426
rect 48470 40017 48476 40414
rect 48514 40017 48520 40414
rect 48470 40005 48520 40017
rect 48788 40414 48838 40426
rect 48788 40017 48794 40414
rect 48832 40017 48838 40414
rect 48788 40005 48838 40017
rect 49106 40414 49156 40426
rect 49106 40017 49112 40414
rect 49150 40017 49156 40414
rect 49106 40005 49156 40017
rect 49424 40414 49474 40426
rect 49424 40017 49430 40414
rect 49468 40017 49474 40414
rect 49424 40005 49474 40017
rect 49742 40414 49792 40426
rect 49742 40017 49748 40414
rect 49786 40017 49792 40414
rect 49742 40005 49792 40017
rect 50060 40414 50110 40426
rect 50060 40017 50066 40414
rect 50104 40017 50110 40414
rect 50060 40005 50110 40017
rect 50378 40414 50428 40426
rect 50378 40017 50384 40414
rect 50422 40017 50428 40414
rect 50378 40005 50428 40017
rect 50696 40414 50746 40426
rect 50696 40017 50702 40414
rect 50740 40017 50746 40414
rect 50696 40005 50746 40017
rect 51014 40414 51064 40426
rect 51014 40017 51020 40414
rect 51058 40017 51064 40414
rect 51014 40005 51064 40017
rect 51332 40414 51382 40426
rect 51332 40017 51338 40414
rect 51376 40017 51382 40414
rect 51332 40005 51382 40017
rect 51650 40414 51700 40426
rect 51650 40017 51656 40414
rect 51694 40017 51700 40414
rect 51650 40005 51700 40017
rect 51968 40414 52018 40426
rect 51968 40017 51974 40414
rect 52012 40017 52018 40414
rect 51968 40005 52018 40017
rect 52286 40414 52336 40426
rect 52286 40017 52292 40414
rect 52330 40017 52336 40414
rect 52286 40005 52336 40017
rect 52604 40414 52654 40426
rect 52604 40017 52610 40414
rect 52648 40017 52654 40414
rect 52604 40005 52654 40017
rect 52922 40414 52972 40426
rect 52922 40017 52928 40414
rect 52966 40017 52972 40414
rect 52922 40005 52972 40017
rect 53240 40414 53290 40426
rect 53240 40017 53246 40414
rect 53284 40017 53290 40414
rect 53240 40005 53290 40017
rect 53558 40414 53608 40426
rect 53558 40017 53564 40414
rect 53602 40017 53608 40414
rect 53558 40005 53608 40017
rect 53876 40414 53926 40426
rect 53876 40017 53882 40414
rect 53920 40017 53926 40414
rect 53876 40005 53926 40017
rect 54194 40414 54244 40426
rect 54194 40017 54200 40414
rect 54238 40017 54244 40414
rect 54194 40005 54244 40017
rect 54512 40414 54562 40426
rect 54512 40017 54518 40414
rect 54556 40017 54562 40414
rect 54512 40005 54562 40017
rect 54830 40414 54880 40426
rect 54830 40017 54836 40414
rect 54874 40017 54880 40414
rect 54830 40005 54880 40017
rect 55148 40414 55198 40426
rect 55148 40017 55154 40414
rect 55192 40017 55198 40414
rect 55148 40005 55198 40017
rect 55466 40414 55516 40426
rect 55466 40017 55472 40414
rect 55510 40017 55516 40414
rect 55466 40005 55516 40017
rect 55784 40414 55834 40426
rect 55784 40017 55790 40414
rect 55828 40017 55834 40414
rect 55784 40005 55834 40017
rect 56102 40414 56152 40426
rect 56102 40017 56108 40414
rect 56146 40017 56152 40414
rect 56102 40005 56152 40017
rect 56420 40414 56470 40426
rect 56420 40017 56426 40414
rect 56464 40017 56470 40414
rect 56420 40005 56470 40017
rect 56738 40414 56788 40426
rect 56738 40017 56744 40414
rect 56782 40017 56788 40414
rect 56738 40005 56788 40017
rect 57056 40414 57106 40426
rect 57056 40017 57062 40414
rect 57100 40017 57106 40414
rect 57056 40005 57106 40017
rect 57374 40414 57424 40426
rect 57374 40017 57380 40414
rect 57418 40017 57424 40414
rect 57374 40005 57424 40017
rect 57692 40414 57742 40426
rect 57692 40017 57698 40414
rect 57736 40017 57742 40414
rect 57692 40005 57742 40017
rect 58010 40414 58060 40426
rect 58010 40017 58016 40414
rect 58054 40017 58060 40414
rect 58010 40005 58060 40017
rect 58328 40414 58378 40426
rect 58328 40017 58334 40414
rect 58372 40017 58378 40414
rect 58328 40005 58378 40017
rect 58646 40414 58696 40426
rect 58646 40017 58652 40414
rect 58690 40017 58696 40414
rect 58646 40005 58696 40017
rect 58964 40414 59014 40426
rect 58964 40017 58970 40414
rect 59008 40017 59014 40414
rect 58964 40005 59014 40017
rect 59282 40414 59332 40426
rect 59282 40017 59288 40414
rect 59326 40017 59332 40414
rect 59282 40005 59332 40017
rect 59600 40414 59650 40426
rect 59600 40017 59606 40414
rect 59644 40017 59650 40414
rect 59600 40005 59650 40017
rect 59918 40414 59968 40426
rect 59918 40017 59924 40414
rect 59962 40017 59968 40414
rect 59918 40005 59968 40017
rect 60236 40414 60286 40426
rect 60236 40017 60242 40414
rect 60280 40017 60286 40414
rect 60236 40005 60286 40017
rect 60554 40414 60604 40426
rect 60554 40017 60560 40414
rect 60598 40017 60604 40414
rect 60554 40005 60604 40017
rect 60872 40414 60922 40426
rect 60872 40017 60878 40414
rect 60916 40017 60922 40414
rect 60872 40005 60922 40017
rect 61190 40414 61240 40426
rect 61190 40017 61196 40414
rect 61234 40017 61240 40414
rect 61190 40005 61240 40017
rect 61508 40414 61558 40426
rect 61508 40017 61514 40414
rect 61552 40017 61558 40414
rect 61508 40005 61558 40017
rect 61826 40414 61876 40426
rect 61826 40017 61832 40414
rect 61870 40017 61876 40414
rect 61826 40005 61876 40017
rect 62144 40414 62194 40426
rect 62144 40017 62150 40414
rect 62188 40017 62194 40414
rect 62144 40005 62194 40017
rect 62462 40414 62512 40426
rect 62462 40017 62468 40414
rect 62506 40017 62512 40414
rect 62462 40005 62512 40017
rect 62780 40414 62830 40426
rect 62780 40017 62786 40414
rect 62824 40017 62830 40414
rect 62780 40005 62830 40017
rect 63098 40414 63148 40426
rect 63098 40017 63104 40414
rect 63142 40017 63148 40414
rect 63098 40005 63148 40017
rect 63416 40414 63466 40426
rect 63416 40017 63422 40414
rect 63460 40017 63466 40414
rect 63416 40005 63466 40017
rect -63466 -40017 -63416 -40005
rect -63466 -40414 -63460 -40017
rect -63422 -40414 -63416 -40017
rect -63466 -40426 -63416 -40414
rect -63148 -40017 -63098 -40005
rect -63148 -40414 -63142 -40017
rect -63104 -40414 -63098 -40017
rect -63148 -40426 -63098 -40414
rect -62830 -40017 -62780 -40005
rect -62830 -40414 -62824 -40017
rect -62786 -40414 -62780 -40017
rect -62830 -40426 -62780 -40414
rect -62512 -40017 -62462 -40005
rect -62512 -40414 -62506 -40017
rect -62468 -40414 -62462 -40017
rect -62512 -40426 -62462 -40414
rect -62194 -40017 -62144 -40005
rect -62194 -40414 -62188 -40017
rect -62150 -40414 -62144 -40017
rect -62194 -40426 -62144 -40414
rect -61876 -40017 -61826 -40005
rect -61876 -40414 -61870 -40017
rect -61832 -40414 -61826 -40017
rect -61876 -40426 -61826 -40414
rect -61558 -40017 -61508 -40005
rect -61558 -40414 -61552 -40017
rect -61514 -40414 -61508 -40017
rect -61558 -40426 -61508 -40414
rect -61240 -40017 -61190 -40005
rect -61240 -40414 -61234 -40017
rect -61196 -40414 -61190 -40017
rect -61240 -40426 -61190 -40414
rect -60922 -40017 -60872 -40005
rect -60922 -40414 -60916 -40017
rect -60878 -40414 -60872 -40017
rect -60922 -40426 -60872 -40414
rect -60604 -40017 -60554 -40005
rect -60604 -40414 -60598 -40017
rect -60560 -40414 -60554 -40017
rect -60604 -40426 -60554 -40414
rect -60286 -40017 -60236 -40005
rect -60286 -40414 -60280 -40017
rect -60242 -40414 -60236 -40017
rect -60286 -40426 -60236 -40414
rect -59968 -40017 -59918 -40005
rect -59968 -40414 -59962 -40017
rect -59924 -40414 -59918 -40017
rect -59968 -40426 -59918 -40414
rect -59650 -40017 -59600 -40005
rect -59650 -40414 -59644 -40017
rect -59606 -40414 -59600 -40017
rect -59650 -40426 -59600 -40414
rect -59332 -40017 -59282 -40005
rect -59332 -40414 -59326 -40017
rect -59288 -40414 -59282 -40017
rect -59332 -40426 -59282 -40414
rect -59014 -40017 -58964 -40005
rect -59014 -40414 -59008 -40017
rect -58970 -40414 -58964 -40017
rect -59014 -40426 -58964 -40414
rect -58696 -40017 -58646 -40005
rect -58696 -40414 -58690 -40017
rect -58652 -40414 -58646 -40017
rect -58696 -40426 -58646 -40414
rect -58378 -40017 -58328 -40005
rect -58378 -40414 -58372 -40017
rect -58334 -40414 -58328 -40017
rect -58378 -40426 -58328 -40414
rect -58060 -40017 -58010 -40005
rect -58060 -40414 -58054 -40017
rect -58016 -40414 -58010 -40017
rect -58060 -40426 -58010 -40414
rect -57742 -40017 -57692 -40005
rect -57742 -40414 -57736 -40017
rect -57698 -40414 -57692 -40017
rect -57742 -40426 -57692 -40414
rect -57424 -40017 -57374 -40005
rect -57424 -40414 -57418 -40017
rect -57380 -40414 -57374 -40017
rect -57424 -40426 -57374 -40414
rect -57106 -40017 -57056 -40005
rect -57106 -40414 -57100 -40017
rect -57062 -40414 -57056 -40017
rect -57106 -40426 -57056 -40414
rect -56788 -40017 -56738 -40005
rect -56788 -40414 -56782 -40017
rect -56744 -40414 -56738 -40017
rect -56788 -40426 -56738 -40414
rect -56470 -40017 -56420 -40005
rect -56470 -40414 -56464 -40017
rect -56426 -40414 -56420 -40017
rect -56470 -40426 -56420 -40414
rect -56152 -40017 -56102 -40005
rect -56152 -40414 -56146 -40017
rect -56108 -40414 -56102 -40017
rect -56152 -40426 -56102 -40414
rect -55834 -40017 -55784 -40005
rect -55834 -40414 -55828 -40017
rect -55790 -40414 -55784 -40017
rect -55834 -40426 -55784 -40414
rect -55516 -40017 -55466 -40005
rect -55516 -40414 -55510 -40017
rect -55472 -40414 -55466 -40017
rect -55516 -40426 -55466 -40414
rect -55198 -40017 -55148 -40005
rect -55198 -40414 -55192 -40017
rect -55154 -40414 -55148 -40017
rect -55198 -40426 -55148 -40414
rect -54880 -40017 -54830 -40005
rect -54880 -40414 -54874 -40017
rect -54836 -40414 -54830 -40017
rect -54880 -40426 -54830 -40414
rect -54562 -40017 -54512 -40005
rect -54562 -40414 -54556 -40017
rect -54518 -40414 -54512 -40017
rect -54562 -40426 -54512 -40414
rect -54244 -40017 -54194 -40005
rect -54244 -40414 -54238 -40017
rect -54200 -40414 -54194 -40017
rect -54244 -40426 -54194 -40414
rect -53926 -40017 -53876 -40005
rect -53926 -40414 -53920 -40017
rect -53882 -40414 -53876 -40017
rect -53926 -40426 -53876 -40414
rect -53608 -40017 -53558 -40005
rect -53608 -40414 -53602 -40017
rect -53564 -40414 -53558 -40017
rect -53608 -40426 -53558 -40414
rect -53290 -40017 -53240 -40005
rect -53290 -40414 -53284 -40017
rect -53246 -40414 -53240 -40017
rect -53290 -40426 -53240 -40414
rect -52972 -40017 -52922 -40005
rect -52972 -40414 -52966 -40017
rect -52928 -40414 -52922 -40017
rect -52972 -40426 -52922 -40414
rect -52654 -40017 -52604 -40005
rect -52654 -40414 -52648 -40017
rect -52610 -40414 -52604 -40017
rect -52654 -40426 -52604 -40414
rect -52336 -40017 -52286 -40005
rect -52336 -40414 -52330 -40017
rect -52292 -40414 -52286 -40017
rect -52336 -40426 -52286 -40414
rect -52018 -40017 -51968 -40005
rect -52018 -40414 -52012 -40017
rect -51974 -40414 -51968 -40017
rect -52018 -40426 -51968 -40414
rect -51700 -40017 -51650 -40005
rect -51700 -40414 -51694 -40017
rect -51656 -40414 -51650 -40017
rect -51700 -40426 -51650 -40414
rect -51382 -40017 -51332 -40005
rect -51382 -40414 -51376 -40017
rect -51338 -40414 -51332 -40017
rect -51382 -40426 -51332 -40414
rect -51064 -40017 -51014 -40005
rect -51064 -40414 -51058 -40017
rect -51020 -40414 -51014 -40017
rect -51064 -40426 -51014 -40414
rect -50746 -40017 -50696 -40005
rect -50746 -40414 -50740 -40017
rect -50702 -40414 -50696 -40017
rect -50746 -40426 -50696 -40414
rect -50428 -40017 -50378 -40005
rect -50428 -40414 -50422 -40017
rect -50384 -40414 -50378 -40017
rect -50428 -40426 -50378 -40414
rect -50110 -40017 -50060 -40005
rect -50110 -40414 -50104 -40017
rect -50066 -40414 -50060 -40017
rect -50110 -40426 -50060 -40414
rect -49792 -40017 -49742 -40005
rect -49792 -40414 -49786 -40017
rect -49748 -40414 -49742 -40017
rect -49792 -40426 -49742 -40414
rect -49474 -40017 -49424 -40005
rect -49474 -40414 -49468 -40017
rect -49430 -40414 -49424 -40017
rect -49474 -40426 -49424 -40414
rect -49156 -40017 -49106 -40005
rect -49156 -40414 -49150 -40017
rect -49112 -40414 -49106 -40017
rect -49156 -40426 -49106 -40414
rect -48838 -40017 -48788 -40005
rect -48838 -40414 -48832 -40017
rect -48794 -40414 -48788 -40017
rect -48838 -40426 -48788 -40414
rect -48520 -40017 -48470 -40005
rect -48520 -40414 -48514 -40017
rect -48476 -40414 -48470 -40017
rect -48520 -40426 -48470 -40414
rect -48202 -40017 -48152 -40005
rect -48202 -40414 -48196 -40017
rect -48158 -40414 -48152 -40017
rect -48202 -40426 -48152 -40414
rect -47884 -40017 -47834 -40005
rect -47884 -40414 -47878 -40017
rect -47840 -40414 -47834 -40017
rect -47884 -40426 -47834 -40414
rect -47566 -40017 -47516 -40005
rect -47566 -40414 -47560 -40017
rect -47522 -40414 -47516 -40017
rect -47566 -40426 -47516 -40414
rect -47248 -40017 -47198 -40005
rect -47248 -40414 -47242 -40017
rect -47204 -40414 -47198 -40017
rect -47248 -40426 -47198 -40414
rect -46930 -40017 -46880 -40005
rect -46930 -40414 -46924 -40017
rect -46886 -40414 -46880 -40017
rect -46930 -40426 -46880 -40414
rect -46612 -40017 -46562 -40005
rect -46612 -40414 -46606 -40017
rect -46568 -40414 -46562 -40017
rect -46612 -40426 -46562 -40414
rect -46294 -40017 -46244 -40005
rect -46294 -40414 -46288 -40017
rect -46250 -40414 -46244 -40017
rect -46294 -40426 -46244 -40414
rect -45976 -40017 -45926 -40005
rect -45976 -40414 -45970 -40017
rect -45932 -40414 -45926 -40017
rect -45976 -40426 -45926 -40414
rect -45658 -40017 -45608 -40005
rect -45658 -40414 -45652 -40017
rect -45614 -40414 -45608 -40017
rect -45658 -40426 -45608 -40414
rect -45340 -40017 -45290 -40005
rect -45340 -40414 -45334 -40017
rect -45296 -40414 -45290 -40017
rect -45340 -40426 -45290 -40414
rect -45022 -40017 -44972 -40005
rect -45022 -40414 -45016 -40017
rect -44978 -40414 -44972 -40017
rect -45022 -40426 -44972 -40414
rect -44704 -40017 -44654 -40005
rect -44704 -40414 -44698 -40017
rect -44660 -40414 -44654 -40017
rect -44704 -40426 -44654 -40414
rect -44386 -40017 -44336 -40005
rect -44386 -40414 -44380 -40017
rect -44342 -40414 -44336 -40017
rect -44386 -40426 -44336 -40414
rect -44068 -40017 -44018 -40005
rect -44068 -40414 -44062 -40017
rect -44024 -40414 -44018 -40017
rect -44068 -40426 -44018 -40414
rect -43750 -40017 -43700 -40005
rect -43750 -40414 -43744 -40017
rect -43706 -40414 -43700 -40017
rect -43750 -40426 -43700 -40414
rect -43432 -40017 -43382 -40005
rect -43432 -40414 -43426 -40017
rect -43388 -40414 -43382 -40017
rect -43432 -40426 -43382 -40414
rect -43114 -40017 -43064 -40005
rect -43114 -40414 -43108 -40017
rect -43070 -40414 -43064 -40017
rect -43114 -40426 -43064 -40414
rect -42796 -40017 -42746 -40005
rect -42796 -40414 -42790 -40017
rect -42752 -40414 -42746 -40017
rect -42796 -40426 -42746 -40414
rect -42478 -40017 -42428 -40005
rect -42478 -40414 -42472 -40017
rect -42434 -40414 -42428 -40017
rect -42478 -40426 -42428 -40414
rect -42160 -40017 -42110 -40005
rect -42160 -40414 -42154 -40017
rect -42116 -40414 -42110 -40017
rect -42160 -40426 -42110 -40414
rect -41842 -40017 -41792 -40005
rect -41842 -40414 -41836 -40017
rect -41798 -40414 -41792 -40017
rect -41842 -40426 -41792 -40414
rect -41524 -40017 -41474 -40005
rect -41524 -40414 -41518 -40017
rect -41480 -40414 -41474 -40017
rect -41524 -40426 -41474 -40414
rect -41206 -40017 -41156 -40005
rect -41206 -40414 -41200 -40017
rect -41162 -40414 -41156 -40017
rect -41206 -40426 -41156 -40414
rect -40888 -40017 -40838 -40005
rect -40888 -40414 -40882 -40017
rect -40844 -40414 -40838 -40017
rect -40888 -40426 -40838 -40414
rect -40570 -40017 -40520 -40005
rect -40570 -40414 -40564 -40017
rect -40526 -40414 -40520 -40017
rect -40570 -40426 -40520 -40414
rect -40252 -40017 -40202 -40005
rect -40252 -40414 -40246 -40017
rect -40208 -40414 -40202 -40017
rect -40252 -40426 -40202 -40414
rect -39934 -40017 -39884 -40005
rect -39934 -40414 -39928 -40017
rect -39890 -40414 -39884 -40017
rect -39934 -40426 -39884 -40414
rect -39616 -40017 -39566 -40005
rect -39616 -40414 -39610 -40017
rect -39572 -40414 -39566 -40017
rect -39616 -40426 -39566 -40414
rect -39298 -40017 -39248 -40005
rect -39298 -40414 -39292 -40017
rect -39254 -40414 -39248 -40017
rect -39298 -40426 -39248 -40414
rect -38980 -40017 -38930 -40005
rect -38980 -40414 -38974 -40017
rect -38936 -40414 -38930 -40017
rect -38980 -40426 -38930 -40414
rect -38662 -40017 -38612 -40005
rect -38662 -40414 -38656 -40017
rect -38618 -40414 -38612 -40017
rect -38662 -40426 -38612 -40414
rect -38344 -40017 -38294 -40005
rect -38344 -40414 -38338 -40017
rect -38300 -40414 -38294 -40017
rect -38344 -40426 -38294 -40414
rect -38026 -40017 -37976 -40005
rect -38026 -40414 -38020 -40017
rect -37982 -40414 -37976 -40017
rect -38026 -40426 -37976 -40414
rect -37708 -40017 -37658 -40005
rect -37708 -40414 -37702 -40017
rect -37664 -40414 -37658 -40017
rect -37708 -40426 -37658 -40414
rect -37390 -40017 -37340 -40005
rect -37390 -40414 -37384 -40017
rect -37346 -40414 -37340 -40017
rect -37390 -40426 -37340 -40414
rect -37072 -40017 -37022 -40005
rect -37072 -40414 -37066 -40017
rect -37028 -40414 -37022 -40017
rect -37072 -40426 -37022 -40414
rect -36754 -40017 -36704 -40005
rect -36754 -40414 -36748 -40017
rect -36710 -40414 -36704 -40017
rect -36754 -40426 -36704 -40414
rect -36436 -40017 -36386 -40005
rect -36436 -40414 -36430 -40017
rect -36392 -40414 -36386 -40017
rect -36436 -40426 -36386 -40414
rect -36118 -40017 -36068 -40005
rect -36118 -40414 -36112 -40017
rect -36074 -40414 -36068 -40017
rect -36118 -40426 -36068 -40414
rect -35800 -40017 -35750 -40005
rect -35800 -40414 -35794 -40017
rect -35756 -40414 -35750 -40017
rect -35800 -40426 -35750 -40414
rect -35482 -40017 -35432 -40005
rect -35482 -40414 -35476 -40017
rect -35438 -40414 -35432 -40017
rect -35482 -40426 -35432 -40414
rect -35164 -40017 -35114 -40005
rect -35164 -40414 -35158 -40017
rect -35120 -40414 -35114 -40017
rect -35164 -40426 -35114 -40414
rect -34846 -40017 -34796 -40005
rect -34846 -40414 -34840 -40017
rect -34802 -40414 -34796 -40017
rect -34846 -40426 -34796 -40414
rect -34528 -40017 -34478 -40005
rect -34528 -40414 -34522 -40017
rect -34484 -40414 -34478 -40017
rect -34528 -40426 -34478 -40414
rect -34210 -40017 -34160 -40005
rect -34210 -40414 -34204 -40017
rect -34166 -40414 -34160 -40017
rect -34210 -40426 -34160 -40414
rect -33892 -40017 -33842 -40005
rect -33892 -40414 -33886 -40017
rect -33848 -40414 -33842 -40017
rect -33892 -40426 -33842 -40414
rect -33574 -40017 -33524 -40005
rect -33574 -40414 -33568 -40017
rect -33530 -40414 -33524 -40017
rect -33574 -40426 -33524 -40414
rect -33256 -40017 -33206 -40005
rect -33256 -40414 -33250 -40017
rect -33212 -40414 -33206 -40017
rect -33256 -40426 -33206 -40414
rect -32938 -40017 -32888 -40005
rect -32938 -40414 -32932 -40017
rect -32894 -40414 -32888 -40017
rect -32938 -40426 -32888 -40414
rect -32620 -40017 -32570 -40005
rect -32620 -40414 -32614 -40017
rect -32576 -40414 -32570 -40017
rect -32620 -40426 -32570 -40414
rect -32302 -40017 -32252 -40005
rect -32302 -40414 -32296 -40017
rect -32258 -40414 -32252 -40017
rect -32302 -40426 -32252 -40414
rect -31984 -40017 -31934 -40005
rect -31984 -40414 -31978 -40017
rect -31940 -40414 -31934 -40017
rect -31984 -40426 -31934 -40414
rect -31666 -40017 -31616 -40005
rect -31666 -40414 -31660 -40017
rect -31622 -40414 -31616 -40017
rect -31666 -40426 -31616 -40414
rect -31348 -40017 -31298 -40005
rect -31348 -40414 -31342 -40017
rect -31304 -40414 -31298 -40017
rect -31348 -40426 -31298 -40414
rect -31030 -40017 -30980 -40005
rect -31030 -40414 -31024 -40017
rect -30986 -40414 -30980 -40017
rect -31030 -40426 -30980 -40414
rect -30712 -40017 -30662 -40005
rect -30712 -40414 -30706 -40017
rect -30668 -40414 -30662 -40017
rect -30712 -40426 -30662 -40414
rect -30394 -40017 -30344 -40005
rect -30394 -40414 -30388 -40017
rect -30350 -40414 -30344 -40017
rect -30394 -40426 -30344 -40414
rect -30076 -40017 -30026 -40005
rect -30076 -40414 -30070 -40017
rect -30032 -40414 -30026 -40017
rect -30076 -40426 -30026 -40414
rect -29758 -40017 -29708 -40005
rect -29758 -40414 -29752 -40017
rect -29714 -40414 -29708 -40017
rect -29758 -40426 -29708 -40414
rect -29440 -40017 -29390 -40005
rect -29440 -40414 -29434 -40017
rect -29396 -40414 -29390 -40017
rect -29440 -40426 -29390 -40414
rect -29122 -40017 -29072 -40005
rect -29122 -40414 -29116 -40017
rect -29078 -40414 -29072 -40017
rect -29122 -40426 -29072 -40414
rect -28804 -40017 -28754 -40005
rect -28804 -40414 -28798 -40017
rect -28760 -40414 -28754 -40017
rect -28804 -40426 -28754 -40414
rect -28486 -40017 -28436 -40005
rect -28486 -40414 -28480 -40017
rect -28442 -40414 -28436 -40017
rect -28486 -40426 -28436 -40414
rect -28168 -40017 -28118 -40005
rect -28168 -40414 -28162 -40017
rect -28124 -40414 -28118 -40017
rect -28168 -40426 -28118 -40414
rect -27850 -40017 -27800 -40005
rect -27850 -40414 -27844 -40017
rect -27806 -40414 -27800 -40017
rect -27850 -40426 -27800 -40414
rect -27532 -40017 -27482 -40005
rect -27532 -40414 -27526 -40017
rect -27488 -40414 -27482 -40017
rect -27532 -40426 -27482 -40414
rect -27214 -40017 -27164 -40005
rect -27214 -40414 -27208 -40017
rect -27170 -40414 -27164 -40017
rect -27214 -40426 -27164 -40414
rect -26896 -40017 -26846 -40005
rect -26896 -40414 -26890 -40017
rect -26852 -40414 -26846 -40017
rect -26896 -40426 -26846 -40414
rect -26578 -40017 -26528 -40005
rect -26578 -40414 -26572 -40017
rect -26534 -40414 -26528 -40017
rect -26578 -40426 -26528 -40414
rect -26260 -40017 -26210 -40005
rect -26260 -40414 -26254 -40017
rect -26216 -40414 -26210 -40017
rect -26260 -40426 -26210 -40414
rect -25942 -40017 -25892 -40005
rect -25942 -40414 -25936 -40017
rect -25898 -40414 -25892 -40017
rect -25942 -40426 -25892 -40414
rect -25624 -40017 -25574 -40005
rect -25624 -40414 -25618 -40017
rect -25580 -40414 -25574 -40017
rect -25624 -40426 -25574 -40414
rect -25306 -40017 -25256 -40005
rect -25306 -40414 -25300 -40017
rect -25262 -40414 -25256 -40017
rect -25306 -40426 -25256 -40414
rect -24988 -40017 -24938 -40005
rect -24988 -40414 -24982 -40017
rect -24944 -40414 -24938 -40017
rect -24988 -40426 -24938 -40414
rect -24670 -40017 -24620 -40005
rect -24670 -40414 -24664 -40017
rect -24626 -40414 -24620 -40017
rect -24670 -40426 -24620 -40414
rect -24352 -40017 -24302 -40005
rect -24352 -40414 -24346 -40017
rect -24308 -40414 -24302 -40017
rect -24352 -40426 -24302 -40414
rect -24034 -40017 -23984 -40005
rect -24034 -40414 -24028 -40017
rect -23990 -40414 -23984 -40017
rect -24034 -40426 -23984 -40414
rect -23716 -40017 -23666 -40005
rect -23716 -40414 -23710 -40017
rect -23672 -40414 -23666 -40017
rect -23716 -40426 -23666 -40414
rect -23398 -40017 -23348 -40005
rect -23398 -40414 -23392 -40017
rect -23354 -40414 -23348 -40017
rect -23398 -40426 -23348 -40414
rect -23080 -40017 -23030 -40005
rect -23080 -40414 -23074 -40017
rect -23036 -40414 -23030 -40017
rect -23080 -40426 -23030 -40414
rect -22762 -40017 -22712 -40005
rect -22762 -40414 -22756 -40017
rect -22718 -40414 -22712 -40017
rect -22762 -40426 -22712 -40414
rect -22444 -40017 -22394 -40005
rect -22444 -40414 -22438 -40017
rect -22400 -40414 -22394 -40017
rect -22444 -40426 -22394 -40414
rect -22126 -40017 -22076 -40005
rect -22126 -40414 -22120 -40017
rect -22082 -40414 -22076 -40017
rect -22126 -40426 -22076 -40414
rect -21808 -40017 -21758 -40005
rect -21808 -40414 -21802 -40017
rect -21764 -40414 -21758 -40017
rect -21808 -40426 -21758 -40414
rect -21490 -40017 -21440 -40005
rect -21490 -40414 -21484 -40017
rect -21446 -40414 -21440 -40017
rect -21490 -40426 -21440 -40414
rect -21172 -40017 -21122 -40005
rect -21172 -40414 -21166 -40017
rect -21128 -40414 -21122 -40017
rect -21172 -40426 -21122 -40414
rect -20854 -40017 -20804 -40005
rect -20854 -40414 -20848 -40017
rect -20810 -40414 -20804 -40017
rect -20854 -40426 -20804 -40414
rect -20536 -40017 -20486 -40005
rect -20536 -40414 -20530 -40017
rect -20492 -40414 -20486 -40017
rect -20536 -40426 -20486 -40414
rect -20218 -40017 -20168 -40005
rect -20218 -40414 -20212 -40017
rect -20174 -40414 -20168 -40017
rect -20218 -40426 -20168 -40414
rect -19900 -40017 -19850 -40005
rect -19900 -40414 -19894 -40017
rect -19856 -40414 -19850 -40017
rect -19900 -40426 -19850 -40414
rect -19582 -40017 -19532 -40005
rect -19582 -40414 -19576 -40017
rect -19538 -40414 -19532 -40017
rect -19582 -40426 -19532 -40414
rect -19264 -40017 -19214 -40005
rect -19264 -40414 -19258 -40017
rect -19220 -40414 -19214 -40017
rect -19264 -40426 -19214 -40414
rect -18946 -40017 -18896 -40005
rect -18946 -40414 -18940 -40017
rect -18902 -40414 -18896 -40017
rect -18946 -40426 -18896 -40414
rect -18628 -40017 -18578 -40005
rect -18628 -40414 -18622 -40017
rect -18584 -40414 -18578 -40017
rect -18628 -40426 -18578 -40414
rect -18310 -40017 -18260 -40005
rect -18310 -40414 -18304 -40017
rect -18266 -40414 -18260 -40017
rect -18310 -40426 -18260 -40414
rect -17992 -40017 -17942 -40005
rect -17992 -40414 -17986 -40017
rect -17948 -40414 -17942 -40017
rect -17992 -40426 -17942 -40414
rect -17674 -40017 -17624 -40005
rect -17674 -40414 -17668 -40017
rect -17630 -40414 -17624 -40017
rect -17674 -40426 -17624 -40414
rect -17356 -40017 -17306 -40005
rect -17356 -40414 -17350 -40017
rect -17312 -40414 -17306 -40017
rect -17356 -40426 -17306 -40414
rect -17038 -40017 -16988 -40005
rect -17038 -40414 -17032 -40017
rect -16994 -40414 -16988 -40017
rect -17038 -40426 -16988 -40414
rect -16720 -40017 -16670 -40005
rect -16720 -40414 -16714 -40017
rect -16676 -40414 -16670 -40017
rect -16720 -40426 -16670 -40414
rect -16402 -40017 -16352 -40005
rect -16402 -40414 -16396 -40017
rect -16358 -40414 -16352 -40017
rect -16402 -40426 -16352 -40414
rect -16084 -40017 -16034 -40005
rect -16084 -40414 -16078 -40017
rect -16040 -40414 -16034 -40017
rect -16084 -40426 -16034 -40414
rect -15766 -40017 -15716 -40005
rect -15766 -40414 -15760 -40017
rect -15722 -40414 -15716 -40017
rect -15766 -40426 -15716 -40414
rect -15448 -40017 -15398 -40005
rect -15448 -40414 -15442 -40017
rect -15404 -40414 -15398 -40017
rect -15448 -40426 -15398 -40414
rect -15130 -40017 -15080 -40005
rect -15130 -40414 -15124 -40017
rect -15086 -40414 -15080 -40017
rect -15130 -40426 -15080 -40414
rect -14812 -40017 -14762 -40005
rect -14812 -40414 -14806 -40017
rect -14768 -40414 -14762 -40017
rect -14812 -40426 -14762 -40414
rect -14494 -40017 -14444 -40005
rect -14494 -40414 -14488 -40017
rect -14450 -40414 -14444 -40017
rect -14494 -40426 -14444 -40414
rect -14176 -40017 -14126 -40005
rect -14176 -40414 -14170 -40017
rect -14132 -40414 -14126 -40017
rect -14176 -40426 -14126 -40414
rect -13858 -40017 -13808 -40005
rect -13858 -40414 -13852 -40017
rect -13814 -40414 -13808 -40017
rect -13858 -40426 -13808 -40414
rect -13540 -40017 -13490 -40005
rect -13540 -40414 -13534 -40017
rect -13496 -40414 -13490 -40017
rect -13540 -40426 -13490 -40414
rect -13222 -40017 -13172 -40005
rect -13222 -40414 -13216 -40017
rect -13178 -40414 -13172 -40017
rect -13222 -40426 -13172 -40414
rect -12904 -40017 -12854 -40005
rect -12904 -40414 -12898 -40017
rect -12860 -40414 -12854 -40017
rect -12904 -40426 -12854 -40414
rect -12586 -40017 -12536 -40005
rect -12586 -40414 -12580 -40017
rect -12542 -40414 -12536 -40017
rect -12586 -40426 -12536 -40414
rect -12268 -40017 -12218 -40005
rect -12268 -40414 -12262 -40017
rect -12224 -40414 -12218 -40017
rect -12268 -40426 -12218 -40414
rect -11950 -40017 -11900 -40005
rect -11950 -40414 -11944 -40017
rect -11906 -40414 -11900 -40017
rect -11950 -40426 -11900 -40414
rect -11632 -40017 -11582 -40005
rect -11632 -40414 -11626 -40017
rect -11588 -40414 -11582 -40017
rect -11632 -40426 -11582 -40414
rect -11314 -40017 -11264 -40005
rect -11314 -40414 -11308 -40017
rect -11270 -40414 -11264 -40017
rect -11314 -40426 -11264 -40414
rect -10996 -40017 -10946 -40005
rect -10996 -40414 -10990 -40017
rect -10952 -40414 -10946 -40017
rect -10996 -40426 -10946 -40414
rect -10678 -40017 -10628 -40005
rect -10678 -40414 -10672 -40017
rect -10634 -40414 -10628 -40017
rect -10678 -40426 -10628 -40414
rect -10360 -40017 -10310 -40005
rect -10360 -40414 -10354 -40017
rect -10316 -40414 -10310 -40017
rect -10360 -40426 -10310 -40414
rect -10042 -40017 -9992 -40005
rect -10042 -40414 -10036 -40017
rect -9998 -40414 -9992 -40017
rect -10042 -40426 -9992 -40414
rect -9724 -40017 -9674 -40005
rect -9724 -40414 -9718 -40017
rect -9680 -40414 -9674 -40017
rect -9724 -40426 -9674 -40414
rect -9406 -40017 -9356 -40005
rect -9406 -40414 -9400 -40017
rect -9362 -40414 -9356 -40017
rect -9406 -40426 -9356 -40414
rect -9088 -40017 -9038 -40005
rect -9088 -40414 -9082 -40017
rect -9044 -40414 -9038 -40017
rect -9088 -40426 -9038 -40414
rect -8770 -40017 -8720 -40005
rect -8770 -40414 -8764 -40017
rect -8726 -40414 -8720 -40017
rect -8770 -40426 -8720 -40414
rect -8452 -40017 -8402 -40005
rect -8452 -40414 -8446 -40017
rect -8408 -40414 -8402 -40017
rect -8452 -40426 -8402 -40414
rect -8134 -40017 -8084 -40005
rect -8134 -40414 -8128 -40017
rect -8090 -40414 -8084 -40017
rect -8134 -40426 -8084 -40414
rect -7816 -40017 -7766 -40005
rect -7816 -40414 -7810 -40017
rect -7772 -40414 -7766 -40017
rect -7816 -40426 -7766 -40414
rect -7498 -40017 -7448 -40005
rect -7498 -40414 -7492 -40017
rect -7454 -40414 -7448 -40017
rect -7498 -40426 -7448 -40414
rect -7180 -40017 -7130 -40005
rect -7180 -40414 -7174 -40017
rect -7136 -40414 -7130 -40017
rect -7180 -40426 -7130 -40414
rect -6862 -40017 -6812 -40005
rect -6862 -40414 -6856 -40017
rect -6818 -40414 -6812 -40017
rect -6862 -40426 -6812 -40414
rect -6544 -40017 -6494 -40005
rect -6544 -40414 -6538 -40017
rect -6500 -40414 -6494 -40017
rect -6544 -40426 -6494 -40414
rect -6226 -40017 -6176 -40005
rect -6226 -40414 -6220 -40017
rect -6182 -40414 -6176 -40017
rect -6226 -40426 -6176 -40414
rect -5908 -40017 -5858 -40005
rect -5908 -40414 -5902 -40017
rect -5864 -40414 -5858 -40017
rect -5908 -40426 -5858 -40414
rect -5590 -40017 -5540 -40005
rect -5590 -40414 -5584 -40017
rect -5546 -40414 -5540 -40017
rect -5590 -40426 -5540 -40414
rect -5272 -40017 -5222 -40005
rect -5272 -40414 -5266 -40017
rect -5228 -40414 -5222 -40017
rect -5272 -40426 -5222 -40414
rect -4954 -40017 -4904 -40005
rect -4954 -40414 -4948 -40017
rect -4910 -40414 -4904 -40017
rect -4954 -40426 -4904 -40414
rect -4636 -40017 -4586 -40005
rect -4636 -40414 -4630 -40017
rect -4592 -40414 -4586 -40017
rect -4636 -40426 -4586 -40414
rect -4318 -40017 -4268 -40005
rect -4318 -40414 -4312 -40017
rect -4274 -40414 -4268 -40017
rect -4318 -40426 -4268 -40414
rect -4000 -40017 -3950 -40005
rect -4000 -40414 -3994 -40017
rect -3956 -40414 -3950 -40017
rect -4000 -40426 -3950 -40414
rect -3682 -40017 -3632 -40005
rect -3682 -40414 -3676 -40017
rect -3638 -40414 -3632 -40017
rect -3682 -40426 -3632 -40414
rect -3364 -40017 -3314 -40005
rect -3364 -40414 -3358 -40017
rect -3320 -40414 -3314 -40017
rect -3364 -40426 -3314 -40414
rect -3046 -40017 -2996 -40005
rect -3046 -40414 -3040 -40017
rect -3002 -40414 -2996 -40017
rect -3046 -40426 -2996 -40414
rect -2728 -40017 -2678 -40005
rect -2728 -40414 -2722 -40017
rect -2684 -40414 -2678 -40017
rect -2728 -40426 -2678 -40414
rect -2410 -40017 -2360 -40005
rect -2410 -40414 -2404 -40017
rect -2366 -40414 -2360 -40017
rect -2410 -40426 -2360 -40414
rect -2092 -40017 -2042 -40005
rect -2092 -40414 -2086 -40017
rect -2048 -40414 -2042 -40017
rect -2092 -40426 -2042 -40414
rect -1774 -40017 -1724 -40005
rect -1774 -40414 -1768 -40017
rect -1730 -40414 -1724 -40017
rect -1774 -40426 -1724 -40414
rect -1456 -40017 -1406 -40005
rect -1456 -40414 -1450 -40017
rect -1412 -40414 -1406 -40017
rect -1456 -40426 -1406 -40414
rect -1138 -40017 -1088 -40005
rect -1138 -40414 -1132 -40017
rect -1094 -40414 -1088 -40017
rect -1138 -40426 -1088 -40414
rect -820 -40017 -770 -40005
rect -820 -40414 -814 -40017
rect -776 -40414 -770 -40017
rect -820 -40426 -770 -40414
rect -502 -40017 -452 -40005
rect -502 -40414 -496 -40017
rect -458 -40414 -452 -40017
rect -502 -40426 -452 -40414
rect -184 -40017 -134 -40005
rect -184 -40414 -178 -40017
rect -140 -40414 -134 -40017
rect -184 -40426 -134 -40414
rect 134 -40017 184 -40005
rect 134 -40414 140 -40017
rect 178 -40414 184 -40017
rect 134 -40426 184 -40414
rect 452 -40017 502 -40005
rect 452 -40414 458 -40017
rect 496 -40414 502 -40017
rect 452 -40426 502 -40414
rect 770 -40017 820 -40005
rect 770 -40414 776 -40017
rect 814 -40414 820 -40017
rect 770 -40426 820 -40414
rect 1088 -40017 1138 -40005
rect 1088 -40414 1094 -40017
rect 1132 -40414 1138 -40017
rect 1088 -40426 1138 -40414
rect 1406 -40017 1456 -40005
rect 1406 -40414 1412 -40017
rect 1450 -40414 1456 -40017
rect 1406 -40426 1456 -40414
rect 1724 -40017 1774 -40005
rect 1724 -40414 1730 -40017
rect 1768 -40414 1774 -40017
rect 1724 -40426 1774 -40414
rect 2042 -40017 2092 -40005
rect 2042 -40414 2048 -40017
rect 2086 -40414 2092 -40017
rect 2042 -40426 2092 -40414
rect 2360 -40017 2410 -40005
rect 2360 -40414 2366 -40017
rect 2404 -40414 2410 -40017
rect 2360 -40426 2410 -40414
rect 2678 -40017 2728 -40005
rect 2678 -40414 2684 -40017
rect 2722 -40414 2728 -40017
rect 2678 -40426 2728 -40414
rect 2996 -40017 3046 -40005
rect 2996 -40414 3002 -40017
rect 3040 -40414 3046 -40017
rect 2996 -40426 3046 -40414
rect 3314 -40017 3364 -40005
rect 3314 -40414 3320 -40017
rect 3358 -40414 3364 -40017
rect 3314 -40426 3364 -40414
rect 3632 -40017 3682 -40005
rect 3632 -40414 3638 -40017
rect 3676 -40414 3682 -40017
rect 3632 -40426 3682 -40414
rect 3950 -40017 4000 -40005
rect 3950 -40414 3956 -40017
rect 3994 -40414 4000 -40017
rect 3950 -40426 4000 -40414
rect 4268 -40017 4318 -40005
rect 4268 -40414 4274 -40017
rect 4312 -40414 4318 -40017
rect 4268 -40426 4318 -40414
rect 4586 -40017 4636 -40005
rect 4586 -40414 4592 -40017
rect 4630 -40414 4636 -40017
rect 4586 -40426 4636 -40414
rect 4904 -40017 4954 -40005
rect 4904 -40414 4910 -40017
rect 4948 -40414 4954 -40017
rect 4904 -40426 4954 -40414
rect 5222 -40017 5272 -40005
rect 5222 -40414 5228 -40017
rect 5266 -40414 5272 -40017
rect 5222 -40426 5272 -40414
rect 5540 -40017 5590 -40005
rect 5540 -40414 5546 -40017
rect 5584 -40414 5590 -40017
rect 5540 -40426 5590 -40414
rect 5858 -40017 5908 -40005
rect 5858 -40414 5864 -40017
rect 5902 -40414 5908 -40017
rect 5858 -40426 5908 -40414
rect 6176 -40017 6226 -40005
rect 6176 -40414 6182 -40017
rect 6220 -40414 6226 -40017
rect 6176 -40426 6226 -40414
rect 6494 -40017 6544 -40005
rect 6494 -40414 6500 -40017
rect 6538 -40414 6544 -40017
rect 6494 -40426 6544 -40414
rect 6812 -40017 6862 -40005
rect 6812 -40414 6818 -40017
rect 6856 -40414 6862 -40017
rect 6812 -40426 6862 -40414
rect 7130 -40017 7180 -40005
rect 7130 -40414 7136 -40017
rect 7174 -40414 7180 -40017
rect 7130 -40426 7180 -40414
rect 7448 -40017 7498 -40005
rect 7448 -40414 7454 -40017
rect 7492 -40414 7498 -40017
rect 7448 -40426 7498 -40414
rect 7766 -40017 7816 -40005
rect 7766 -40414 7772 -40017
rect 7810 -40414 7816 -40017
rect 7766 -40426 7816 -40414
rect 8084 -40017 8134 -40005
rect 8084 -40414 8090 -40017
rect 8128 -40414 8134 -40017
rect 8084 -40426 8134 -40414
rect 8402 -40017 8452 -40005
rect 8402 -40414 8408 -40017
rect 8446 -40414 8452 -40017
rect 8402 -40426 8452 -40414
rect 8720 -40017 8770 -40005
rect 8720 -40414 8726 -40017
rect 8764 -40414 8770 -40017
rect 8720 -40426 8770 -40414
rect 9038 -40017 9088 -40005
rect 9038 -40414 9044 -40017
rect 9082 -40414 9088 -40017
rect 9038 -40426 9088 -40414
rect 9356 -40017 9406 -40005
rect 9356 -40414 9362 -40017
rect 9400 -40414 9406 -40017
rect 9356 -40426 9406 -40414
rect 9674 -40017 9724 -40005
rect 9674 -40414 9680 -40017
rect 9718 -40414 9724 -40017
rect 9674 -40426 9724 -40414
rect 9992 -40017 10042 -40005
rect 9992 -40414 9998 -40017
rect 10036 -40414 10042 -40017
rect 9992 -40426 10042 -40414
rect 10310 -40017 10360 -40005
rect 10310 -40414 10316 -40017
rect 10354 -40414 10360 -40017
rect 10310 -40426 10360 -40414
rect 10628 -40017 10678 -40005
rect 10628 -40414 10634 -40017
rect 10672 -40414 10678 -40017
rect 10628 -40426 10678 -40414
rect 10946 -40017 10996 -40005
rect 10946 -40414 10952 -40017
rect 10990 -40414 10996 -40017
rect 10946 -40426 10996 -40414
rect 11264 -40017 11314 -40005
rect 11264 -40414 11270 -40017
rect 11308 -40414 11314 -40017
rect 11264 -40426 11314 -40414
rect 11582 -40017 11632 -40005
rect 11582 -40414 11588 -40017
rect 11626 -40414 11632 -40017
rect 11582 -40426 11632 -40414
rect 11900 -40017 11950 -40005
rect 11900 -40414 11906 -40017
rect 11944 -40414 11950 -40017
rect 11900 -40426 11950 -40414
rect 12218 -40017 12268 -40005
rect 12218 -40414 12224 -40017
rect 12262 -40414 12268 -40017
rect 12218 -40426 12268 -40414
rect 12536 -40017 12586 -40005
rect 12536 -40414 12542 -40017
rect 12580 -40414 12586 -40017
rect 12536 -40426 12586 -40414
rect 12854 -40017 12904 -40005
rect 12854 -40414 12860 -40017
rect 12898 -40414 12904 -40017
rect 12854 -40426 12904 -40414
rect 13172 -40017 13222 -40005
rect 13172 -40414 13178 -40017
rect 13216 -40414 13222 -40017
rect 13172 -40426 13222 -40414
rect 13490 -40017 13540 -40005
rect 13490 -40414 13496 -40017
rect 13534 -40414 13540 -40017
rect 13490 -40426 13540 -40414
rect 13808 -40017 13858 -40005
rect 13808 -40414 13814 -40017
rect 13852 -40414 13858 -40017
rect 13808 -40426 13858 -40414
rect 14126 -40017 14176 -40005
rect 14126 -40414 14132 -40017
rect 14170 -40414 14176 -40017
rect 14126 -40426 14176 -40414
rect 14444 -40017 14494 -40005
rect 14444 -40414 14450 -40017
rect 14488 -40414 14494 -40017
rect 14444 -40426 14494 -40414
rect 14762 -40017 14812 -40005
rect 14762 -40414 14768 -40017
rect 14806 -40414 14812 -40017
rect 14762 -40426 14812 -40414
rect 15080 -40017 15130 -40005
rect 15080 -40414 15086 -40017
rect 15124 -40414 15130 -40017
rect 15080 -40426 15130 -40414
rect 15398 -40017 15448 -40005
rect 15398 -40414 15404 -40017
rect 15442 -40414 15448 -40017
rect 15398 -40426 15448 -40414
rect 15716 -40017 15766 -40005
rect 15716 -40414 15722 -40017
rect 15760 -40414 15766 -40017
rect 15716 -40426 15766 -40414
rect 16034 -40017 16084 -40005
rect 16034 -40414 16040 -40017
rect 16078 -40414 16084 -40017
rect 16034 -40426 16084 -40414
rect 16352 -40017 16402 -40005
rect 16352 -40414 16358 -40017
rect 16396 -40414 16402 -40017
rect 16352 -40426 16402 -40414
rect 16670 -40017 16720 -40005
rect 16670 -40414 16676 -40017
rect 16714 -40414 16720 -40017
rect 16670 -40426 16720 -40414
rect 16988 -40017 17038 -40005
rect 16988 -40414 16994 -40017
rect 17032 -40414 17038 -40017
rect 16988 -40426 17038 -40414
rect 17306 -40017 17356 -40005
rect 17306 -40414 17312 -40017
rect 17350 -40414 17356 -40017
rect 17306 -40426 17356 -40414
rect 17624 -40017 17674 -40005
rect 17624 -40414 17630 -40017
rect 17668 -40414 17674 -40017
rect 17624 -40426 17674 -40414
rect 17942 -40017 17992 -40005
rect 17942 -40414 17948 -40017
rect 17986 -40414 17992 -40017
rect 17942 -40426 17992 -40414
rect 18260 -40017 18310 -40005
rect 18260 -40414 18266 -40017
rect 18304 -40414 18310 -40017
rect 18260 -40426 18310 -40414
rect 18578 -40017 18628 -40005
rect 18578 -40414 18584 -40017
rect 18622 -40414 18628 -40017
rect 18578 -40426 18628 -40414
rect 18896 -40017 18946 -40005
rect 18896 -40414 18902 -40017
rect 18940 -40414 18946 -40017
rect 18896 -40426 18946 -40414
rect 19214 -40017 19264 -40005
rect 19214 -40414 19220 -40017
rect 19258 -40414 19264 -40017
rect 19214 -40426 19264 -40414
rect 19532 -40017 19582 -40005
rect 19532 -40414 19538 -40017
rect 19576 -40414 19582 -40017
rect 19532 -40426 19582 -40414
rect 19850 -40017 19900 -40005
rect 19850 -40414 19856 -40017
rect 19894 -40414 19900 -40017
rect 19850 -40426 19900 -40414
rect 20168 -40017 20218 -40005
rect 20168 -40414 20174 -40017
rect 20212 -40414 20218 -40017
rect 20168 -40426 20218 -40414
rect 20486 -40017 20536 -40005
rect 20486 -40414 20492 -40017
rect 20530 -40414 20536 -40017
rect 20486 -40426 20536 -40414
rect 20804 -40017 20854 -40005
rect 20804 -40414 20810 -40017
rect 20848 -40414 20854 -40017
rect 20804 -40426 20854 -40414
rect 21122 -40017 21172 -40005
rect 21122 -40414 21128 -40017
rect 21166 -40414 21172 -40017
rect 21122 -40426 21172 -40414
rect 21440 -40017 21490 -40005
rect 21440 -40414 21446 -40017
rect 21484 -40414 21490 -40017
rect 21440 -40426 21490 -40414
rect 21758 -40017 21808 -40005
rect 21758 -40414 21764 -40017
rect 21802 -40414 21808 -40017
rect 21758 -40426 21808 -40414
rect 22076 -40017 22126 -40005
rect 22076 -40414 22082 -40017
rect 22120 -40414 22126 -40017
rect 22076 -40426 22126 -40414
rect 22394 -40017 22444 -40005
rect 22394 -40414 22400 -40017
rect 22438 -40414 22444 -40017
rect 22394 -40426 22444 -40414
rect 22712 -40017 22762 -40005
rect 22712 -40414 22718 -40017
rect 22756 -40414 22762 -40017
rect 22712 -40426 22762 -40414
rect 23030 -40017 23080 -40005
rect 23030 -40414 23036 -40017
rect 23074 -40414 23080 -40017
rect 23030 -40426 23080 -40414
rect 23348 -40017 23398 -40005
rect 23348 -40414 23354 -40017
rect 23392 -40414 23398 -40017
rect 23348 -40426 23398 -40414
rect 23666 -40017 23716 -40005
rect 23666 -40414 23672 -40017
rect 23710 -40414 23716 -40017
rect 23666 -40426 23716 -40414
rect 23984 -40017 24034 -40005
rect 23984 -40414 23990 -40017
rect 24028 -40414 24034 -40017
rect 23984 -40426 24034 -40414
rect 24302 -40017 24352 -40005
rect 24302 -40414 24308 -40017
rect 24346 -40414 24352 -40017
rect 24302 -40426 24352 -40414
rect 24620 -40017 24670 -40005
rect 24620 -40414 24626 -40017
rect 24664 -40414 24670 -40017
rect 24620 -40426 24670 -40414
rect 24938 -40017 24988 -40005
rect 24938 -40414 24944 -40017
rect 24982 -40414 24988 -40017
rect 24938 -40426 24988 -40414
rect 25256 -40017 25306 -40005
rect 25256 -40414 25262 -40017
rect 25300 -40414 25306 -40017
rect 25256 -40426 25306 -40414
rect 25574 -40017 25624 -40005
rect 25574 -40414 25580 -40017
rect 25618 -40414 25624 -40017
rect 25574 -40426 25624 -40414
rect 25892 -40017 25942 -40005
rect 25892 -40414 25898 -40017
rect 25936 -40414 25942 -40017
rect 25892 -40426 25942 -40414
rect 26210 -40017 26260 -40005
rect 26210 -40414 26216 -40017
rect 26254 -40414 26260 -40017
rect 26210 -40426 26260 -40414
rect 26528 -40017 26578 -40005
rect 26528 -40414 26534 -40017
rect 26572 -40414 26578 -40017
rect 26528 -40426 26578 -40414
rect 26846 -40017 26896 -40005
rect 26846 -40414 26852 -40017
rect 26890 -40414 26896 -40017
rect 26846 -40426 26896 -40414
rect 27164 -40017 27214 -40005
rect 27164 -40414 27170 -40017
rect 27208 -40414 27214 -40017
rect 27164 -40426 27214 -40414
rect 27482 -40017 27532 -40005
rect 27482 -40414 27488 -40017
rect 27526 -40414 27532 -40017
rect 27482 -40426 27532 -40414
rect 27800 -40017 27850 -40005
rect 27800 -40414 27806 -40017
rect 27844 -40414 27850 -40017
rect 27800 -40426 27850 -40414
rect 28118 -40017 28168 -40005
rect 28118 -40414 28124 -40017
rect 28162 -40414 28168 -40017
rect 28118 -40426 28168 -40414
rect 28436 -40017 28486 -40005
rect 28436 -40414 28442 -40017
rect 28480 -40414 28486 -40017
rect 28436 -40426 28486 -40414
rect 28754 -40017 28804 -40005
rect 28754 -40414 28760 -40017
rect 28798 -40414 28804 -40017
rect 28754 -40426 28804 -40414
rect 29072 -40017 29122 -40005
rect 29072 -40414 29078 -40017
rect 29116 -40414 29122 -40017
rect 29072 -40426 29122 -40414
rect 29390 -40017 29440 -40005
rect 29390 -40414 29396 -40017
rect 29434 -40414 29440 -40017
rect 29390 -40426 29440 -40414
rect 29708 -40017 29758 -40005
rect 29708 -40414 29714 -40017
rect 29752 -40414 29758 -40017
rect 29708 -40426 29758 -40414
rect 30026 -40017 30076 -40005
rect 30026 -40414 30032 -40017
rect 30070 -40414 30076 -40017
rect 30026 -40426 30076 -40414
rect 30344 -40017 30394 -40005
rect 30344 -40414 30350 -40017
rect 30388 -40414 30394 -40017
rect 30344 -40426 30394 -40414
rect 30662 -40017 30712 -40005
rect 30662 -40414 30668 -40017
rect 30706 -40414 30712 -40017
rect 30662 -40426 30712 -40414
rect 30980 -40017 31030 -40005
rect 30980 -40414 30986 -40017
rect 31024 -40414 31030 -40017
rect 30980 -40426 31030 -40414
rect 31298 -40017 31348 -40005
rect 31298 -40414 31304 -40017
rect 31342 -40414 31348 -40017
rect 31298 -40426 31348 -40414
rect 31616 -40017 31666 -40005
rect 31616 -40414 31622 -40017
rect 31660 -40414 31666 -40017
rect 31616 -40426 31666 -40414
rect 31934 -40017 31984 -40005
rect 31934 -40414 31940 -40017
rect 31978 -40414 31984 -40017
rect 31934 -40426 31984 -40414
rect 32252 -40017 32302 -40005
rect 32252 -40414 32258 -40017
rect 32296 -40414 32302 -40017
rect 32252 -40426 32302 -40414
rect 32570 -40017 32620 -40005
rect 32570 -40414 32576 -40017
rect 32614 -40414 32620 -40017
rect 32570 -40426 32620 -40414
rect 32888 -40017 32938 -40005
rect 32888 -40414 32894 -40017
rect 32932 -40414 32938 -40017
rect 32888 -40426 32938 -40414
rect 33206 -40017 33256 -40005
rect 33206 -40414 33212 -40017
rect 33250 -40414 33256 -40017
rect 33206 -40426 33256 -40414
rect 33524 -40017 33574 -40005
rect 33524 -40414 33530 -40017
rect 33568 -40414 33574 -40017
rect 33524 -40426 33574 -40414
rect 33842 -40017 33892 -40005
rect 33842 -40414 33848 -40017
rect 33886 -40414 33892 -40017
rect 33842 -40426 33892 -40414
rect 34160 -40017 34210 -40005
rect 34160 -40414 34166 -40017
rect 34204 -40414 34210 -40017
rect 34160 -40426 34210 -40414
rect 34478 -40017 34528 -40005
rect 34478 -40414 34484 -40017
rect 34522 -40414 34528 -40017
rect 34478 -40426 34528 -40414
rect 34796 -40017 34846 -40005
rect 34796 -40414 34802 -40017
rect 34840 -40414 34846 -40017
rect 34796 -40426 34846 -40414
rect 35114 -40017 35164 -40005
rect 35114 -40414 35120 -40017
rect 35158 -40414 35164 -40017
rect 35114 -40426 35164 -40414
rect 35432 -40017 35482 -40005
rect 35432 -40414 35438 -40017
rect 35476 -40414 35482 -40017
rect 35432 -40426 35482 -40414
rect 35750 -40017 35800 -40005
rect 35750 -40414 35756 -40017
rect 35794 -40414 35800 -40017
rect 35750 -40426 35800 -40414
rect 36068 -40017 36118 -40005
rect 36068 -40414 36074 -40017
rect 36112 -40414 36118 -40017
rect 36068 -40426 36118 -40414
rect 36386 -40017 36436 -40005
rect 36386 -40414 36392 -40017
rect 36430 -40414 36436 -40017
rect 36386 -40426 36436 -40414
rect 36704 -40017 36754 -40005
rect 36704 -40414 36710 -40017
rect 36748 -40414 36754 -40017
rect 36704 -40426 36754 -40414
rect 37022 -40017 37072 -40005
rect 37022 -40414 37028 -40017
rect 37066 -40414 37072 -40017
rect 37022 -40426 37072 -40414
rect 37340 -40017 37390 -40005
rect 37340 -40414 37346 -40017
rect 37384 -40414 37390 -40017
rect 37340 -40426 37390 -40414
rect 37658 -40017 37708 -40005
rect 37658 -40414 37664 -40017
rect 37702 -40414 37708 -40017
rect 37658 -40426 37708 -40414
rect 37976 -40017 38026 -40005
rect 37976 -40414 37982 -40017
rect 38020 -40414 38026 -40017
rect 37976 -40426 38026 -40414
rect 38294 -40017 38344 -40005
rect 38294 -40414 38300 -40017
rect 38338 -40414 38344 -40017
rect 38294 -40426 38344 -40414
rect 38612 -40017 38662 -40005
rect 38612 -40414 38618 -40017
rect 38656 -40414 38662 -40017
rect 38612 -40426 38662 -40414
rect 38930 -40017 38980 -40005
rect 38930 -40414 38936 -40017
rect 38974 -40414 38980 -40017
rect 38930 -40426 38980 -40414
rect 39248 -40017 39298 -40005
rect 39248 -40414 39254 -40017
rect 39292 -40414 39298 -40017
rect 39248 -40426 39298 -40414
rect 39566 -40017 39616 -40005
rect 39566 -40414 39572 -40017
rect 39610 -40414 39616 -40017
rect 39566 -40426 39616 -40414
rect 39884 -40017 39934 -40005
rect 39884 -40414 39890 -40017
rect 39928 -40414 39934 -40017
rect 39884 -40426 39934 -40414
rect 40202 -40017 40252 -40005
rect 40202 -40414 40208 -40017
rect 40246 -40414 40252 -40017
rect 40202 -40426 40252 -40414
rect 40520 -40017 40570 -40005
rect 40520 -40414 40526 -40017
rect 40564 -40414 40570 -40017
rect 40520 -40426 40570 -40414
rect 40838 -40017 40888 -40005
rect 40838 -40414 40844 -40017
rect 40882 -40414 40888 -40017
rect 40838 -40426 40888 -40414
rect 41156 -40017 41206 -40005
rect 41156 -40414 41162 -40017
rect 41200 -40414 41206 -40017
rect 41156 -40426 41206 -40414
rect 41474 -40017 41524 -40005
rect 41474 -40414 41480 -40017
rect 41518 -40414 41524 -40017
rect 41474 -40426 41524 -40414
rect 41792 -40017 41842 -40005
rect 41792 -40414 41798 -40017
rect 41836 -40414 41842 -40017
rect 41792 -40426 41842 -40414
rect 42110 -40017 42160 -40005
rect 42110 -40414 42116 -40017
rect 42154 -40414 42160 -40017
rect 42110 -40426 42160 -40414
rect 42428 -40017 42478 -40005
rect 42428 -40414 42434 -40017
rect 42472 -40414 42478 -40017
rect 42428 -40426 42478 -40414
rect 42746 -40017 42796 -40005
rect 42746 -40414 42752 -40017
rect 42790 -40414 42796 -40017
rect 42746 -40426 42796 -40414
rect 43064 -40017 43114 -40005
rect 43064 -40414 43070 -40017
rect 43108 -40414 43114 -40017
rect 43064 -40426 43114 -40414
rect 43382 -40017 43432 -40005
rect 43382 -40414 43388 -40017
rect 43426 -40414 43432 -40017
rect 43382 -40426 43432 -40414
rect 43700 -40017 43750 -40005
rect 43700 -40414 43706 -40017
rect 43744 -40414 43750 -40017
rect 43700 -40426 43750 -40414
rect 44018 -40017 44068 -40005
rect 44018 -40414 44024 -40017
rect 44062 -40414 44068 -40017
rect 44018 -40426 44068 -40414
rect 44336 -40017 44386 -40005
rect 44336 -40414 44342 -40017
rect 44380 -40414 44386 -40017
rect 44336 -40426 44386 -40414
rect 44654 -40017 44704 -40005
rect 44654 -40414 44660 -40017
rect 44698 -40414 44704 -40017
rect 44654 -40426 44704 -40414
rect 44972 -40017 45022 -40005
rect 44972 -40414 44978 -40017
rect 45016 -40414 45022 -40017
rect 44972 -40426 45022 -40414
rect 45290 -40017 45340 -40005
rect 45290 -40414 45296 -40017
rect 45334 -40414 45340 -40017
rect 45290 -40426 45340 -40414
rect 45608 -40017 45658 -40005
rect 45608 -40414 45614 -40017
rect 45652 -40414 45658 -40017
rect 45608 -40426 45658 -40414
rect 45926 -40017 45976 -40005
rect 45926 -40414 45932 -40017
rect 45970 -40414 45976 -40017
rect 45926 -40426 45976 -40414
rect 46244 -40017 46294 -40005
rect 46244 -40414 46250 -40017
rect 46288 -40414 46294 -40017
rect 46244 -40426 46294 -40414
rect 46562 -40017 46612 -40005
rect 46562 -40414 46568 -40017
rect 46606 -40414 46612 -40017
rect 46562 -40426 46612 -40414
rect 46880 -40017 46930 -40005
rect 46880 -40414 46886 -40017
rect 46924 -40414 46930 -40017
rect 46880 -40426 46930 -40414
rect 47198 -40017 47248 -40005
rect 47198 -40414 47204 -40017
rect 47242 -40414 47248 -40017
rect 47198 -40426 47248 -40414
rect 47516 -40017 47566 -40005
rect 47516 -40414 47522 -40017
rect 47560 -40414 47566 -40017
rect 47516 -40426 47566 -40414
rect 47834 -40017 47884 -40005
rect 47834 -40414 47840 -40017
rect 47878 -40414 47884 -40017
rect 47834 -40426 47884 -40414
rect 48152 -40017 48202 -40005
rect 48152 -40414 48158 -40017
rect 48196 -40414 48202 -40017
rect 48152 -40426 48202 -40414
rect 48470 -40017 48520 -40005
rect 48470 -40414 48476 -40017
rect 48514 -40414 48520 -40017
rect 48470 -40426 48520 -40414
rect 48788 -40017 48838 -40005
rect 48788 -40414 48794 -40017
rect 48832 -40414 48838 -40017
rect 48788 -40426 48838 -40414
rect 49106 -40017 49156 -40005
rect 49106 -40414 49112 -40017
rect 49150 -40414 49156 -40017
rect 49106 -40426 49156 -40414
rect 49424 -40017 49474 -40005
rect 49424 -40414 49430 -40017
rect 49468 -40414 49474 -40017
rect 49424 -40426 49474 -40414
rect 49742 -40017 49792 -40005
rect 49742 -40414 49748 -40017
rect 49786 -40414 49792 -40017
rect 49742 -40426 49792 -40414
rect 50060 -40017 50110 -40005
rect 50060 -40414 50066 -40017
rect 50104 -40414 50110 -40017
rect 50060 -40426 50110 -40414
rect 50378 -40017 50428 -40005
rect 50378 -40414 50384 -40017
rect 50422 -40414 50428 -40017
rect 50378 -40426 50428 -40414
rect 50696 -40017 50746 -40005
rect 50696 -40414 50702 -40017
rect 50740 -40414 50746 -40017
rect 50696 -40426 50746 -40414
rect 51014 -40017 51064 -40005
rect 51014 -40414 51020 -40017
rect 51058 -40414 51064 -40017
rect 51014 -40426 51064 -40414
rect 51332 -40017 51382 -40005
rect 51332 -40414 51338 -40017
rect 51376 -40414 51382 -40017
rect 51332 -40426 51382 -40414
rect 51650 -40017 51700 -40005
rect 51650 -40414 51656 -40017
rect 51694 -40414 51700 -40017
rect 51650 -40426 51700 -40414
rect 51968 -40017 52018 -40005
rect 51968 -40414 51974 -40017
rect 52012 -40414 52018 -40017
rect 51968 -40426 52018 -40414
rect 52286 -40017 52336 -40005
rect 52286 -40414 52292 -40017
rect 52330 -40414 52336 -40017
rect 52286 -40426 52336 -40414
rect 52604 -40017 52654 -40005
rect 52604 -40414 52610 -40017
rect 52648 -40414 52654 -40017
rect 52604 -40426 52654 -40414
rect 52922 -40017 52972 -40005
rect 52922 -40414 52928 -40017
rect 52966 -40414 52972 -40017
rect 52922 -40426 52972 -40414
rect 53240 -40017 53290 -40005
rect 53240 -40414 53246 -40017
rect 53284 -40414 53290 -40017
rect 53240 -40426 53290 -40414
rect 53558 -40017 53608 -40005
rect 53558 -40414 53564 -40017
rect 53602 -40414 53608 -40017
rect 53558 -40426 53608 -40414
rect 53876 -40017 53926 -40005
rect 53876 -40414 53882 -40017
rect 53920 -40414 53926 -40017
rect 53876 -40426 53926 -40414
rect 54194 -40017 54244 -40005
rect 54194 -40414 54200 -40017
rect 54238 -40414 54244 -40017
rect 54194 -40426 54244 -40414
rect 54512 -40017 54562 -40005
rect 54512 -40414 54518 -40017
rect 54556 -40414 54562 -40017
rect 54512 -40426 54562 -40414
rect 54830 -40017 54880 -40005
rect 54830 -40414 54836 -40017
rect 54874 -40414 54880 -40017
rect 54830 -40426 54880 -40414
rect 55148 -40017 55198 -40005
rect 55148 -40414 55154 -40017
rect 55192 -40414 55198 -40017
rect 55148 -40426 55198 -40414
rect 55466 -40017 55516 -40005
rect 55466 -40414 55472 -40017
rect 55510 -40414 55516 -40017
rect 55466 -40426 55516 -40414
rect 55784 -40017 55834 -40005
rect 55784 -40414 55790 -40017
rect 55828 -40414 55834 -40017
rect 55784 -40426 55834 -40414
rect 56102 -40017 56152 -40005
rect 56102 -40414 56108 -40017
rect 56146 -40414 56152 -40017
rect 56102 -40426 56152 -40414
rect 56420 -40017 56470 -40005
rect 56420 -40414 56426 -40017
rect 56464 -40414 56470 -40017
rect 56420 -40426 56470 -40414
rect 56738 -40017 56788 -40005
rect 56738 -40414 56744 -40017
rect 56782 -40414 56788 -40017
rect 56738 -40426 56788 -40414
rect 57056 -40017 57106 -40005
rect 57056 -40414 57062 -40017
rect 57100 -40414 57106 -40017
rect 57056 -40426 57106 -40414
rect 57374 -40017 57424 -40005
rect 57374 -40414 57380 -40017
rect 57418 -40414 57424 -40017
rect 57374 -40426 57424 -40414
rect 57692 -40017 57742 -40005
rect 57692 -40414 57698 -40017
rect 57736 -40414 57742 -40017
rect 57692 -40426 57742 -40414
rect 58010 -40017 58060 -40005
rect 58010 -40414 58016 -40017
rect 58054 -40414 58060 -40017
rect 58010 -40426 58060 -40414
rect 58328 -40017 58378 -40005
rect 58328 -40414 58334 -40017
rect 58372 -40414 58378 -40017
rect 58328 -40426 58378 -40414
rect 58646 -40017 58696 -40005
rect 58646 -40414 58652 -40017
rect 58690 -40414 58696 -40017
rect 58646 -40426 58696 -40414
rect 58964 -40017 59014 -40005
rect 58964 -40414 58970 -40017
rect 59008 -40414 59014 -40017
rect 58964 -40426 59014 -40414
rect 59282 -40017 59332 -40005
rect 59282 -40414 59288 -40017
rect 59326 -40414 59332 -40017
rect 59282 -40426 59332 -40414
rect 59600 -40017 59650 -40005
rect 59600 -40414 59606 -40017
rect 59644 -40414 59650 -40017
rect 59600 -40426 59650 -40414
rect 59918 -40017 59968 -40005
rect 59918 -40414 59924 -40017
rect 59962 -40414 59968 -40017
rect 59918 -40426 59968 -40414
rect 60236 -40017 60286 -40005
rect 60236 -40414 60242 -40017
rect 60280 -40414 60286 -40017
rect 60236 -40426 60286 -40414
rect 60554 -40017 60604 -40005
rect 60554 -40414 60560 -40017
rect 60598 -40414 60604 -40017
rect 60554 -40426 60604 -40414
rect 60872 -40017 60922 -40005
rect 60872 -40414 60878 -40017
rect 60916 -40414 60922 -40017
rect 60872 -40426 60922 -40414
rect 61190 -40017 61240 -40005
rect 61190 -40414 61196 -40017
rect 61234 -40414 61240 -40017
rect 61190 -40426 61240 -40414
rect 61508 -40017 61558 -40005
rect 61508 -40414 61514 -40017
rect 61552 -40414 61558 -40017
rect 61508 -40426 61558 -40414
rect 61826 -40017 61876 -40005
rect 61826 -40414 61832 -40017
rect 61870 -40414 61876 -40017
rect 61826 -40426 61876 -40414
rect 62144 -40017 62194 -40005
rect 62144 -40414 62150 -40017
rect 62188 -40414 62194 -40017
rect 62144 -40426 62194 -40414
rect 62462 -40017 62512 -40005
rect 62462 -40414 62468 -40017
rect 62506 -40414 62512 -40017
rect 62462 -40426 62512 -40414
rect 62780 -40017 62830 -40005
rect 62780 -40414 62786 -40017
rect 62824 -40414 62830 -40017
rect 62780 -40426 62830 -40414
rect 63098 -40017 63148 -40005
rect 63098 -40414 63104 -40017
rect 63142 -40414 63148 -40017
rect 63098 -40426 63148 -40414
rect 63416 -40017 63466 -40005
rect 63416 -40414 63422 -40017
rect 63460 -40414 63466 -40017
rect 63416 -40426 63466 -40414
<< res0p35 >>
rect -63478 -40002 -63404 40002
rect -63160 -40002 -63086 40002
rect -62842 -40002 -62768 40002
rect -62524 -40002 -62450 40002
rect -62206 -40002 -62132 40002
rect -61888 -40002 -61814 40002
rect -61570 -40002 -61496 40002
rect -61252 -40002 -61178 40002
rect -60934 -40002 -60860 40002
rect -60616 -40002 -60542 40002
rect -60298 -40002 -60224 40002
rect -59980 -40002 -59906 40002
rect -59662 -40002 -59588 40002
rect -59344 -40002 -59270 40002
rect -59026 -40002 -58952 40002
rect -58708 -40002 -58634 40002
rect -58390 -40002 -58316 40002
rect -58072 -40002 -57998 40002
rect -57754 -40002 -57680 40002
rect -57436 -40002 -57362 40002
rect -57118 -40002 -57044 40002
rect -56800 -40002 -56726 40002
rect -56482 -40002 -56408 40002
rect -56164 -40002 -56090 40002
rect -55846 -40002 -55772 40002
rect -55528 -40002 -55454 40002
rect -55210 -40002 -55136 40002
rect -54892 -40002 -54818 40002
rect -54574 -40002 -54500 40002
rect -54256 -40002 -54182 40002
rect -53938 -40002 -53864 40002
rect -53620 -40002 -53546 40002
rect -53302 -40002 -53228 40002
rect -52984 -40002 -52910 40002
rect -52666 -40002 -52592 40002
rect -52348 -40002 -52274 40002
rect -52030 -40002 -51956 40002
rect -51712 -40002 -51638 40002
rect -51394 -40002 -51320 40002
rect -51076 -40002 -51002 40002
rect -50758 -40002 -50684 40002
rect -50440 -40002 -50366 40002
rect -50122 -40002 -50048 40002
rect -49804 -40002 -49730 40002
rect -49486 -40002 -49412 40002
rect -49168 -40002 -49094 40002
rect -48850 -40002 -48776 40002
rect -48532 -40002 -48458 40002
rect -48214 -40002 -48140 40002
rect -47896 -40002 -47822 40002
rect -47578 -40002 -47504 40002
rect -47260 -40002 -47186 40002
rect -46942 -40002 -46868 40002
rect -46624 -40002 -46550 40002
rect -46306 -40002 -46232 40002
rect -45988 -40002 -45914 40002
rect -45670 -40002 -45596 40002
rect -45352 -40002 -45278 40002
rect -45034 -40002 -44960 40002
rect -44716 -40002 -44642 40002
rect -44398 -40002 -44324 40002
rect -44080 -40002 -44006 40002
rect -43762 -40002 -43688 40002
rect -43444 -40002 -43370 40002
rect -43126 -40002 -43052 40002
rect -42808 -40002 -42734 40002
rect -42490 -40002 -42416 40002
rect -42172 -40002 -42098 40002
rect -41854 -40002 -41780 40002
rect -41536 -40002 -41462 40002
rect -41218 -40002 -41144 40002
rect -40900 -40002 -40826 40002
rect -40582 -40002 -40508 40002
rect -40264 -40002 -40190 40002
rect -39946 -40002 -39872 40002
rect -39628 -40002 -39554 40002
rect -39310 -40002 -39236 40002
rect -38992 -40002 -38918 40002
rect -38674 -40002 -38600 40002
rect -38356 -40002 -38282 40002
rect -38038 -40002 -37964 40002
rect -37720 -40002 -37646 40002
rect -37402 -40002 -37328 40002
rect -37084 -40002 -37010 40002
rect -36766 -40002 -36692 40002
rect -36448 -40002 -36374 40002
rect -36130 -40002 -36056 40002
rect -35812 -40002 -35738 40002
rect -35494 -40002 -35420 40002
rect -35176 -40002 -35102 40002
rect -34858 -40002 -34784 40002
rect -34540 -40002 -34466 40002
rect -34222 -40002 -34148 40002
rect -33904 -40002 -33830 40002
rect -33586 -40002 -33512 40002
rect -33268 -40002 -33194 40002
rect -32950 -40002 -32876 40002
rect -32632 -40002 -32558 40002
rect -32314 -40002 -32240 40002
rect -31996 -40002 -31922 40002
rect -31678 -40002 -31604 40002
rect -31360 -40002 -31286 40002
rect -31042 -40002 -30968 40002
rect -30724 -40002 -30650 40002
rect -30406 -40002 -30332 40002
rect -30088 -40002 -30014 40002
rect -29770 -40002 -29696 40002
rect -29452 -40002 -29378 40002
rect -29134 -40002 -29060 40002
rect -28816 -40002 -28742 40002
rect -28498 -40002 -28424 40002
rect -28180 -40002 -28106 40002
rect -27862 -40002 -27788 40002
rect -27544 -40002 -27470 40002
rect -27226 -40002 -27152 40002
rect -26908 -40002 -26834 40002
rect -26590 -40002 -26516 40002
rect -26272 -40002 -26198 40002
rect -25954 -40002 -25880 40002
rect -25636 -40002 -25562 40002
rect -25318 -40002 -25244 40002
rect -25000 -40002 -24926 40002
rect -24682 -40002 -24608 40002
rect -24364 -40002 -24290 40002
rect -24046 -40002 -23972 40002
rect -23728 -40002 -23654 40002
rect -23410 -40002 -23336 40002
rect -23092 -40002 -23018 40002
rect -22774 -40002 -22700 40002
rect -22456 -40002 -22382 40002
rect -22138 -40002 -22064 40002
rect -21820 -40002 -21746 40002
rect -21502 -40002 -21428 40002
rect -21184 -40002 -21110 40002
rect -20866 -40002 -20792 40002
rect -20548 -40002 -20474 40002
rect -20230 -40002 -20156 40002
rect -19912 -40002 -19838 40002
rect -19594 -40002 -19520 40002
rect -19276 -40002 -19202 40002
rect -18958 -40002 -18884 40002
rect -18640 -40002 -18566 40002
rect -18322 -40002 -18248 40002
rect -18004 -40002 -17930 40002
rect -17686 -40002 -17612 40002
rect -17368 -40002 -17294 40002
rect -17050 -40002 -16976 40002
rect -16732 -40002 -16658 40002
rect -16414 -40002 -16340 40002
rect -16096 -40002 -16022 40002
rect -15778 -40002 -15704 40002
rect -15460 -40002 -15386 40002
rect -15142 -40002 -15068 40002
rect -14824 -40002 -14750 40002
rect -14506 -40002 -14432 40002
rect -14188 -40002 -14114 40002
rect -13870 -40002 -13796 40002
rect -13552 -40002 -13478 40002
rect -13234 -40002 -13160 40002
rect -12916 -40002 -12842 40002
rect -12598 -40002 -12524 40002
rect -12280 -40002 -12206 40002
rect -11962 -40002 -11888 40002
rect -11644 -40002 -11570 40002
rect -11326 -40002 -11252 40002
rect -11008 -40002 -10934 40002
rect -10690 -40002 -10616 40002
rect -10372 -40002 -10298 40002
rect -10054 -40002 -9980 40002
rect -9736 -40002 -9662 40002
rect -9418 -40002 -9344 40002
rect -9100 -40002 -9026 40002
rect -8782 -40002 -8708 40002
rect -8464 -40002 -8390 40002
rect -8146 -40002 -8072 40002
rect -7828 -40002 -7754 40002
rect -7510 -40002 -7436 40002
rect -7192 -40002 -7118 40002
rect -6874 -40002 -6800 40002
rect -6556 -40002 -6482 40002
rect -6238 -40002 -6164 40002
rect -5920 -40002 -5846 40002
rect -5602 -40002 -5528 40002
rect -5284 -40002 -5210 40002
rect -4966 -40002 -4892 40002
rect -4648 -40002 -4574 40002
rect -4330 -40002 -4256 40002
rect -4012 -40002 -3938 40002
rect -3694 -40002 -3620 40002
rect -3376 -40002 -3302 40002
rect -3058 -40002 -2984 40002
rect -2740 -40002 -2666 40002
rect -2422 -40002 -2348 40002
rect -2104 -40002 -2030 40002
rect -1786 -40002 -1712 40002
rect -1468 -40002 -1394 40002
rect -1150 -40002 -1076 40002
rect -832 -40002 -758 40002
rect -514 -40002 -440 40002
rect -196 -40002 -122 40002
rect 122 -40002 196 40002
rect 440 -40002 514 40002
rect 758 -40002 832 40002
rect 1076 -40002 1150 40002
rect 1394 -40002 1468 40002
rect 1712 -40002 1786 40002
rect 2030 -40002 2104 40002
rect 2348 -40002 2422 40002
rect 2666 -40002 2740 40002
rect 2984 -40002 3058 40002
rect 3302 -40002 3376 40002
rect 3620 -40002 3694 40002
rect 3938 -40002 4012 40002
rect 4256 -40002 4330 40002
rect 4574 -40002 4648 40002
rect 4892 -40002 4966 40002
rect 5210 -40002 5284 40002
rect 5528 -40002 5602 40002
rect 5846 -40002 5920 40002
rect 6164 -40002 6238 40002
rect 6482 -40002 6556 40002
rect 6800 -40002 6874 40002
rect 7118 -40002 7192 40002
rect 7436 -40002 7510 40002
rect 7754 -40002 7828 40002
rect 8072 -40002 8146 40002
rect 8390 -40002 8464 40002
rect 8708 -40002 8782 40002
rect 9026 -40002 9100 40002
rect 9344 -40002 9418 40002
rect 9662 -40002 9736 40002
rect 9980 -40002 10054 40002
rect 10298 -40002 10372 40002
rect 10616 -40002 10690 40002
rect 10934 -40002 11008 40002
rect 11252 -40002 11326 40002
rect 11570 -40002 11644 40002
rect 11888 -40002 11962 40002
rect 12206 -40002 12280 40002
rect 12524 -40002 12598 40002
rect 12842 -40002 12916 40002
rect 13160 -40002 13234 40002
rect 13478 -40002 13552 40002
rect 13796 -40002 13870 40002
rect 14114 -40002 14188 40002
rect 14432 -40002 14506 40002
rect 14750 -40002 14824 40002
rect 15068 -40002 15142 40002
rect 15386 -40002 15460 40002
rect 15704 -40002 15778 40002
rect 16022 -40002 16096 40002
rect 16340 -40002 16414 40002
rect 16658 -40002 16732 40002
rect 16976 -40002 17050 40002
rect 17294 -40002 17368 40002
rect 17612 -40002 17686 40002
rect 17930 -40002 18004 40002
rect 18248 -40002 18322 40002
rect 18566 -40002 18640 40002
rect 18884 -40002 18958 40002
rect 19202 -40002 19276 40002
rect 19520 -40002 19594 40002
rect 19838 -40002 19912 40002
rect 20156 -40002 20230 40002
rect 20474 -40002 20548 40002
rect 20792 -40002 20866 40002
rect 21110 -40002 21184 40002
rect 21428 -40002 21502 40002
rect 21746 -40002 21820 40002
rect 22064 -40002 22138 40002
rect 22382 -40002 22456 40002
rect 22700 -40002 22774 40002
rect 23018 -40002 23092 40002
rect 23336 -40002 23410 40002
rect 23654 -40002 23728 40002
rect 23972 -40002 24046 40002
rect 24290 -40002 24364 40002
rect 24608 -40002 24682 40002
rect 24926 -40002 25000 40002
rect 25244 -40002 25318 40002
rect 25562 -40002 25636 40002
rect 25880 -40002 25954 40002
rect 26198 -40002 26272 40002
rect 26516 -40002 26590 40002
rect 26834 -40002 26908 40002
rect 27152 -40002 27226 40002
rect 27470 -40002 27544 40002
rect 27788 -40002 27862 40002
rect 28106 -40002 28180 40002
rect 28424 -40002 28498 40002
rect 28742 -40002 28816 40002
rect 29060 -40002 29134 40002
rect 29378 -40002 29452 40002
rect 29696 -40002 29770 40002
rect 30014 -40002 30088 40002
rect 30332 -40002 30406 40002
rect 30650 -40002 30724 40002
rect 30968 -40002 31042 40002
rect 31286 -40002 31360 40002
rect 31604 -40002 31678 40002
rect 31922 -40002 31996 40002
rect 32240 -40002 32314 40002
rect 32558 -40002 32632 40002
rect 32876 -40002 32950 40002
rect 33194 -40002 33268 40002
rect 33512 -40002 33586 40002
rect 33830 -40002 33904 40002
rect 34148 -40002 34222 40002
rect 34466 -40002 34540 40002
rect 34784 -40002 34858 40002
rect 35102 -40002 35176 40002
rect 35420 -40002 35494 40002
rect 35738 -40002 35812 40002
rect 36056 -40002 36130 40002
rect 36374 -40002 36448 40002
rect 36692 -40002 36766 40002
rect 37010 -40002 37084 40002
rect 37328 -40002 37402 40002
rect 37646 -40002 37720 40002
rect 37964 -40002 38038 40002
rect 38282 -40002 38356 40002
rect 38600 -40002 38674 40002
rect 38918 -40002 38992 40002
rect 39236 -40002 39310 40002
rect 39554 -40002 39628 40002
rect 39872 -40002 39946 40002
rect 40190 -40002 40264 40002
rect 40508 -40002 40582 40002
rect 40826 -40002 40900 40002
rect 41144 -40002 41218 40002
rect 41462 -40002 41536 40002
rect 41780 -40002 41854 40002
rect 42098 -40002 42172 40002
rect 42416 -40002 42490 40002
rect 42734 -40002 42808 40002
rect 43052 -40002 43126 40002
rect 43370 -40002 43444 40002
rect 43688 -40002 43762 40002
rect 44006 -40002 44080 40002
rect 44324 -40002 44398 40002
rect 44642 -40002 44716 40002
rect 44960 -40002 45034 40002
rect 45278 -40002 45352 40002
rect 45596 -40002 45670 40002
rect 45914 -40002 45988 40002
rect 46232 -40002 46306 40002
rect 46550 -40002 46624 40002
rect 46868 -40002 46942 40002
rect 47186 -40002 47260 40002
rect 47504 -40002 47578 40002
rect 47822 -40002 47896 40002
rect 48140 -40002 48214 40002
rect 48458 -40002 48532 40002
rect 48776 -40002 48850 40002
rect 49094 -40002 49168 40002
rect 49412 -40002 49486 40002
rect 49730 -40002 49804 40002
rect 50048 -40002 50122 40002
rect 50366 -40002 50440 40002
rect 50684 -40002 50758 40002
rect 51002 -40002 51076 40002
rect 51320 -40002 51394 40002
rect 51638 -40002 51712 40002
rect 51956 -40002 52030 40002
rect 52274 -40002 52348 40002
rect 52592 -40002 52666 40002
rect 52910 -40002 52984 40002
rect 53228 -40002 53302 40002
rect 53546 -40002 53620 40002
rect 53864 -40002 53938 40002
rect 54182 -40002 54256 40002
rect 54500 -40002 54574 40002
rect 54818 -40002 54892 40002
rect 55136 -40002 55210 40002
rect 55454 -40002 55528 40002
rect 55772 -40002 55846 40002
rect 56090 -40002 56164 40002
rect 56408 -40002 56482 40002
rect 56726 -40002 56800 40002
rect 57044 -40002 57118 40002
rect 57362 -40002 57436 40002
rect 57680 -40002 57754 40002
rect 57998 -40002 58072 40002
rect 58316 -40002 58390 40002
rect 58634 -40002 58708 40002
rect 58952 -40002 59026 40002
rect 59270 -40002 59344 40002
rect 59588 -40002 59662 40002
rect 59906 -40002 59980 40002
rect 60224 -40002 60298 40002
rect 60542 -40002 60616 40002
rect 60860 -40002 60934 40002
rect 61178 -40002 61252 40002
rect 61496 -40002 61570 40002
rect 61814 -40002 61888 40002
rect 62132 -40002 62206 40002
rect 62450 -40002 62524 40002
rect 62768 -40002 62842 40002
rect 63086 -40002 63160 40002
rect 63404 -40002 63478 40002
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string FIXED_BBOX -63589 -40545 63589 40545
string parameters w 0.350 l 400 m 1 nx 400 wmin 0.350 lmin 0.50 rho 2000 val 2.285meg dummy 0 dw 0.0 term 19.188 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string library sky130
<< end >>
