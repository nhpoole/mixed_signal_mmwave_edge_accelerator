magic
tech sky130A
magscale 1 2
timestamp 1624494425
<< nwell >>
rect 0 0 624 754
<< poly >>
rect 128 360 258 390
rect 128 274 158 360
rect 128 10 158 112
<< metal1 >>
rect 66 0 94 754
rect 530 504 558 754
rect 167 439 219 503
rect 293 438 558 504
rect 530 226 558 438
rect 193 160 558 226
rect 126 -1 190 51
rect 530 0 558 160
<< metal2 >>
rect 0 740 624 768
rect 179 668 207 740
rect 165 620 221 668
rect 179 471 207 620
rect 0 11 624 39
<< metal3 >>
rect 144 595 242 693
use contact_15  contact_15_0
timestamp 1624494425
transform 1 0 125 0 1 -8
box 0 0 66 66
use contact_7  contact_7_1
timestamp 1624494425
transform 1 0 129 0 1 -8
box 0 0 58 66
use contact_8  contact_8_0
timestamp 1624494425
transform 1 0 126 0 1 -7
box 0 0 64 64
use pmos_m1_w0_550_sli_dli  pmos_m1_w0_550_sli_dli_2
timestamp 1624494425
transform 1 0 68 0 1 138
box -59 -54 209 164
use contact_22  contact_22_2
timestamp 1624494425
transform 1 0 170 0 1 160
box 0 0 46 66
use contact_22  contact_22_3
timestamp 1624494425
transform 1 0 70 0 1 160
box 0 0 46 66
use pmos_m1_w0_550_sli_dli  pmos_m1_w0_550_sli_dli_0
timestamp 1624494425
transform 1 0 168 0 1 416
box -59 -54 209 164
use pmos_m1_w0_550_sli_dli  pmos_m1_w0_550_sli_dli_1
timestamp 1624494425
transform 1 0 68 0 1 416
box -59 -54 209 164
use contact_13  contact_13_0
timestamp 1624494425
transform 1 0 168 0 1 603
box -59 -43 109 125
use contact_7  contact_7_0
timestamp 1624494425
transform 1 0 164 0 1 611
box 0 0 58 66
use contact_20  contact_20_1
timestamp 1624494425
transform 1 0 167 0 1 612
box 0 0 52 64
use contact_21  contact_21_0
timestamp 1624494425
transform 1 0 160 0 1 607
box 0 0 66 74
use contact_20  contact_20_0
timestamp 1624494425
transform 1 0 167 0 1 439
box 0 0 52 64
use contact_22  contact_22_0
timestamp 1624494425
transform 1 0 270 0 1 438
box 0 0 46 66
use contact_22  contact_22_1
timestamp 1624494425
transform 1 0 70 0 1 438
box 0 0 46 66
use contact_22  contact_22_4
timestamp 1624494425
transform 1 0 170 0 1 438
box 0 0 46 66
<< labels >>
rlabel metal2 s 0 11 624 39 4 en_bar
rlabel metal3 s 144 595 242 693 4 vdd
rlabel metal1 s 66 0 94 754 4 bl
rlabel metal1 s 530 0 558 754 4 br
<< properties >>
string FIXED_BBOX 0 0 624 754
<< end >>
