magic
tech sky130A
timestamp 1626486988
<< checkpaint >>
rect -717 -717 717 717
<< metal3 >>
rect -87 76 87 87
rect -87 -76 -76 76
rect 76 -76 87 76
rect -87 -87 87 -76
<< via3 >>
rect -76 -76 76 76
<< metal4 >>
rect -87 76 87 87
rect -87 -76 -76 76
rect 76 -76 87 76
rect -87 -87 87 -76
<< end >>
