magic
tech sky130A
magscale 1 2
timestamp 1624477805
<< error_p >>
rect -1871 -200 1871 200
<< nwell >>
rect -1871 -200 1871 200
<< pmos >>
rect -1777 -100 -1577 100
rect -1519 -100 -1319 100
rect -1261 -100 -1061 100
rect -1003 -100 -803 100
rect -745 -100 -545 100
rect -487 -100 -287 100
rect -229 -100 -29 100
rect 29 -100 229 100
rect 287 -100 487 100
rect 545 -100 745 100
rect 803 -100 1003 100
rect 1061 -100 1261 100
rect 1319 -100 1519 100
rect 1577 -100 1777 100
<< pdiff >>
rect -1835 88 -1777 100
rect -1835 -88 -1823 88
rect -1789 -88 -1777 88
rect -1835 -100 -1777 -88
rect -1577 88 -1519 100
rect -1577 -88 -1565 88
rect -1531 -88 -1519 88
rect -1577 -100 -1519 -88
rect -1319 88 -1261 100
rect -1319 -88 -1307 88
rect -1273 -88 -1261 88
rect -1319 -100 -1261 -88
rect -1061 88 -1003 100
rect -1061 -88 -1049 88
rect -1015 -88 -1003 88
rect -1061 -100 -1003 -88
rect -803 88 -745 100
rect -803 -88 -791 88
rect -757 -88 -745 88
rect -803 -100 -745 -88
rect -545 88 -487 100
rect -545 -88 -533 88
rect -499 -88 -487 88
rect -545 -100 -487 -88
rect -287 88 -229 100
rect -287 -88 -275 88
rect -241 -88 -229 88
rect -287 -100 -229 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 229 88 287 100
rect 229 -88 241 88
rect 275 -88 287 88
rect 229 -100 287 -88
rect 487 88 545 100
rect 487 -88 499 88
rect 533 -88 545 88
rect 487 -100 545 -88
rect 745 88 803 100
rect 745 -88 757 88
rect 791 -88 803 88
rect 745 -100 803 -88
rect 1003 88 1061 100
rect 1003 -88 1015 88
rect 1049 -88 1061 88
rect 1003 -100 1061 -88
rect 1261 88 1319 100
rect 1261 -88 1273 88
rect 1307 -88 1319 88
rect 1261 -100 1319 -88
rect 1519 88 1577 100
rect 1519 -88 1531 88
rect 1565 -88 1577 88
rect 1519 -100 1577 -88
rect 1777 88 1835 100
rect 1777 -88 1789 88
rect 1823 -88 1835 88
rect 1777 -100 1835 -88
<< pdiffc >>
rect -1823 -88 -1789 88
rect -1565 -88 -1531 88
rect -1307 -88 -1273 88
rect -1049 -88 -1015 88
rect -791 -88 -757 88
rect -533 -88 -499 88
rect -275 -88 -241 88
rect -17 -88 17 88
rect 241 -88 275 88
rect 499 -88 533 88
rect 757 -88 791 88
rect 1015 -88 1049 88
rect 1273 -88 1307 88
rect 1531 -88 1565 88
rect 1789 -88 1823 88
<< poly >>
rect -1743 181 -1611 197
rect -1743 164 -1727 181
rect -1777 147 -1727 164
rect -1627 164 -1611 181
rect -1485 181 -1353 197
rect -1485 164 -1469 181
rect -1627 147 -1577 164
rect -1777 100 -1577 147
rect -1519 147 -1469 164
rect -1369 164 -1353 181
rect -1227 181 -1095 197
rect -1227 164 -1211 181
rect -1369 147 -1319 164
rect -1519 100 -1319 147
rect -1261 147 -1211 164
rect -1111 164 -1095 181
rect -969 181 -837 197
rect -969 164 -953 181
rect -1111 147 -1061 164
rect -1261 100 -1061 147
rect -1003 147 -953 164
rect -853 164 -837 181
rect -711 181 -579 197
rect -711 164 -695 181
rect -853 147 -803 164
rect -1003 100 -803 147
rect -745 147 -695 164
rect -595 164 -579 181
rect -453 181 -321 197
rect -453 164 -437 181
rect -595 147 -545 164
rect -745 100 -545 147
rect -487 147 -437 164
rect -337 164 -321 181
rect -195 181 -63 197
rect -195 164 -179 181
rect -337 147 -287 164
rect -487 100 -287 147
rect -229 147 -179 164
rect -79 164 -63 181
rect 63 181 195 197
rect 63 164 79 181
rect -79 147 -29 164
rect -229 100 -29 147
rect 29 147 79 164
rect 179 164 195 181
rect 321 181 453 197
rect 321 164 337 181
rect 179 147 229 164
rect 29 100 229 147
rect 287 147 337 164
rect 437 164 453 181
rect 579 181 711 197
rect 579 164 595 181
rect 437 147 487 164
rect 287 100 487 147
rect 545 147 595 164
rect 695 164 711 181
rect 837 181 969 197
rect 837 164 853 181
rect 695 147 745 164
rect 545 100 745 147
rect 803 147 853 164
rect 953 164 969 181
rect 1095 181 1227 197
rect 1095 164 1111 181
rect 953 147 1003 164
rect 803 100 1003 147
rect 1061 147 1111 164
rect 1211 164 1227 181
rect 1353 181 1485 197
rect 1353 164 1369 181
rect 1211 147 1261 164
rect 1061 100 1261 147
rect 1319 147 1369 164
rect 1469 164 1485 181
rect 1611 181 1743 197
rect 1611 164 1627 181
rect 1469 147 1519 164
rect 1319 100 1519 147
rect 1577 147 1627 164
rect 1727 164 1743 181
rect 1727 147 1777 164
rect 1577 100 1777 147
rect -1777 -147 -1577 -100
rect -1777 -164 -1727 -147
rect -1743 -181 -1727 -164
rect -1627 -164 -1577 -147
rect -1519 -147 -1319 -100
rect -1519 -164 -1469 -147
rect -1627 -181 -1611 -164
rect -1743 -197 -1611 -181
rect -1485 -181 -1469 -164
rect -1369 -164 -1319 -147
rect -1261 -147 -1061 -100
rect -1261 -164 -1211 -147
rect -1369 -181 -1353 -164
rect -1485 -197 -1353 -181
rect -1227 -181 -1211 -164
rect -1111 -164 -1061 -147
rect -1003 -147 -803 -100
rect -1003 -164 -953 -147
rect -1111 -181 -1095 -164
rect -1227 -197 -1095 -181
rect -969 -181 -953 -164
rect -853 -164 -803 -147
rect -745 -147 -545 -100
rect -745 -164 -695 -147
rect -853 -181 -837 -164
rect -969 -197 -837 -181
rect -711 -181 -695 -164
rect -595 -164 -545 -147
rect -487 -147 -287 -100
rect -487 -164 -437 -147
rect -595 -181 -579 -164
rect -711 -197 -579 -181
rect -453 -181 -437 -164
rect -337 -164 -287 -147
rect -229 -147 -29 -100
rect -229 -164 -179 -147
rect -337 -181 -321 -164
rect -453 -197 -321 -181
rect -195 -181 -179 -164
rect -79 -164 -29 -147
rect 29 -147 229 -100
rect 29 -164 79 -147
rect -79 -181 -63 -164
rect -195 -197 -63 -181
rect 63 -181 79 -164
rect 179 -164 229 -147
rect 287 -147 487 -100
rect 287 -164 337 -147
rect 179 -181 195 -164
rect 63 -197 195 -181
rect 321 -181 337 -164
rect 437 -164 487 -147
rect 545 -147 745 -100
rect 545 -164 595 -147
rect 437 -181 453 -164
rect 321 -197 453 -181
rect 579 -181 595 -164
rect 695 -164 745 -147
rect 803 -147 1003 -100
rect 803 -164 853 -147
rect 695 -181 711 -164
rect 579 -197 711 -181
rect 837 -181 853 -164
rect 953 -164 1003 -147
rect 1061 -147 1261 -100
rect 1061 -164 1111 -147
rect 953 -181 969 -164
rect 837 -197 969 -181
rect 1095 -181 1111 -164
rect 1211 -164 1261 -147
rect 1319 -147 1519 -100
rect 1319 -164 1369 -147
rect 1211 -181 1227 -164
rect 1095 -197 1227 -181
rect 1353 -181 1369 -164
rect 1469 -164 1519 -147
rect 1577 -147 1777 -100
rect 1577 -164 1627 -147
rect 1469 -181 1485 -164
rect 1353 -197 1485 -181
rect 1611 -181 1627 -164
rect 1727 -164 1777 -147
rect 1727 -181 1743 -164
rect 1611 -197 1743 -181
<< polycont >>
rect -1727 147 -1627 181
rect -1469 147 -1369 181
rect -1211 147 -1111 181
rect -953 147 -853 181
rect -695 147 -595 181
rect -437 147 -337 181
rect -179 147 -79 181
rect 79 147 179 181
rect 337 147 437 181
rect 595 147 695 181
rect 853 147 953 181
rect 1111 147 1211 181
rect 1369 147 1469 181
rect 1627 147 1727 181
rect -1727 -181 -1627 -147
rect -1469 -181 -1369 -147
rect -1211 -181 -1111 -147
rect -953 -181 -853 -147
rect -695 -181 -595 -147
rect -437 -181 -337 -147
rect -179 -181 -79 -147
rect 79 -181 179 -147
rect 337 -181 437 -147
rect 595 -181 695 -147
rect 853 -181 953 -147
rect 1111 -181 1211 -147
rect 1369 -181 1469 -147
rect 1627 -181 1727 -147
<< locali >>
rect -1743 147 -1727 181
rect -1627 147 -1611 181
rect -1485 147 -1469 181
rect -1369 147 -1353 181
rect -1227 147 -1211 181
rect -1111 147 -1095 181
rect -969 147 -953 181
rect -853 147 -837 181
rect -711 147 -695 181
rect -595 147 -579 181
rect -453 147 -437 181
rect -337 147 -321 181
rect -195 147 -179 181
rect -79 147 -63 181
rect 63 147 79 181
rect 179 147 195 181
rect 321 147 337 181
rect 437 147 453 181
rect 579 147 595 181
rect 695 147 711 181
rect 837 147 853 181
rect 953 147 969 181
rect 1095 147 1111 181
rect 1211 147 1227 181
rect 1353 147 1369 181
rect 1469 147 1485 181
rect 1611 147 1627 181
rect 1727 147 1743 181
rect -1823 88 -1789 104
rect -1823 -104 -1789 -88
rect -1565 88 -1531 104
rect -1565 -104 -1531 -88
rect -1307 88 -1273 104
rect -1307 -104 -1273 -88
rect -1049 88 -1015 104
rect -1049 -104 -1015 -88
rect -791 88 -757 104
rect -791 -104 -757 -88
rect -533 88 -499 104
rect -533 -104 -499 -88
rect -275 88 -241 104
rect -275 -104 -241 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 241 88 275 104
rect 241 -104 275 -88
rect 499 88 533 104
rect 499 -104 533 -88
rect 757 88 791 104
rect 757 -104 791 -88
rect 1015 88 1049 104
rect 1015 -104 1049 -88
rect 1273 88 1307 104
rect 1273 -104 1307 -88
rect 1531 88 1565 104
rect 1531 -104 1565 -88
rect 1789 88 1823 104
rect 1789 -104 1823 -88
rect -1743 -181 -1727 -147
rect -1627 -181 -1611 -147
rect -1485 -181 -1469 -147
rect -1369 -181 -1353 -147
rect -1227 -181 -1211 -147
rect -1111 -181 -1095 -147
rect -969 -181 -953 -147
rect -853 -181 -837 -147
rect -711 -181 -695 -147
rect -595 -181 -579 -147
rect -453 -181 -437 -147
rect -337 -181 -321 -147
rect -195 -181 -179 -147
rect -79 -181 -63 -147
rect 63 -181 79 -147
rect 179 -181 195 -147
rect 321 -181 337 -147
rect 437 -181 453 -147
rect 579 -181 595 -147
rect 695 -181 711 -147
rect 837 -181 853 -147
rect 953 -181 969 -147
rect 1095 -181 1111 -147
rect 1211 -181 1227 -147
rect 1353 -181 1369 -147
rect 1469 -181 1485 -147
rect 1611 -181 1627 -147
rect 1727 -181 1743 -147
<< viali >>
rect -1719 147 -1635 181
rect -1461 147 -1377 181
rect -1203 147 -1119 181
rect -945 147 -861 181
rect -687 147 -603 181
rect -429 147 -345 181
rect -171 147 -87 181
rect 87 147 171 181
rect 345 147 429 181
rect 603 147 687 181
rect 861 147 945 181
rect 1119 147 1203 181
rect 1377 147 1461 181
rect 1635 147 1719 181
rect -1823 -88 -1789 88
rect -1565 -88 -1531 88
rect -1307 -88 -1273 88
rect -1049 -88 -1015 88
rect -791 -88 -757 88
rect -533 -88 -499 88
rect -275 -88 -241 88
rect -17 -88 17 88
rect 241 -88 275 88
rect 499 -88 533 88
rect 757 -88 791 88
rect 1015 -88 1049 88
rect 1273 -88 1307 88
rect 1531 -88 1565 88
rect 1789 -88 1823 88
rect -1719 -181 -1635 -147
rect -1461 -181 -1377 -147
rect -1203 -181 -1119 -147
rect -945 -181 -861 -147
rect -687 -181 -603 -147
rect -429 -181 -345 -147
rect -171 -181 -87 -147
rect 87 -181 171 -147
rect 345 -181 429 -147
rect 603 -181 687 -147
rect 861 -181 945 -147
rect 1119 -181 1203 -147
rect 1377 -181 1461 -147
rect 1635 -181 1719 -147
<< metal1 >>
rect -1731 181 -1623 187
rect -1731 147 -1719 181
rect -1635 147 -1623 181
rect -1731 141 -1623 147
rect -1473 181 -1365 187
rect -1473 147 -1461 181
rect -1377 147 -1365 181
rect -1473 141 -1365 147
rect -1215 181 -1107 187
rect -1215 147 -1203 181
rect -1119 147 -1107 181
rect -1215 141 -1107 147
rect -957 181 -849 187
rect -957 147 -945 181
rect -861 147 -849 181
rect -957 141 -849 147
rect -699 181 -591 187
rect -699 147 -687 181
rect -603 147 -591 181
rect -699 141 -591 147
rect -441 181 -333 187
rect -441 147 -429 181
rect -345 147 -333 181
rect -441 141 -333 147
rect -183 181 -75 187
rect -183 147 -171 181
rect -87 147 -75 181
rect -183 141 -75 147
rect 75 181 183 187
rect 75 147 87 181
rect 171 147 183 181
rect 75 141 183 147
rect 333 181 441 187
rect 333 147 345 181
rect 429 147 441 181
rect 333 141 441 147
rect 591 181 699 187
rect 591 147 603 181
rect 687 147 699 181
rect 591 141 699 147
rect 849 181 957 187
rect 849 147 861 181
rect 945 147 957 181
rect 849 141 957 147
rect 1107 181 1215 187
rect 1107 147 1119 181
rect 1203 147 1215 181
rect 1107 141 1215 147
rect 1365 181 1473 187
rect 1365 147 1377 181
rect 1461 147 1473 181
rect 1365 141 1473 147
rect 1623 181 1731 187
rect 1623 147 1635 181
rect 1719 147 1731 181
rect 1623 141 1731 147
rect -1829 88 -1783 100
rect -1829 -88 -1823 88
rect -1789 -88 -1783 88
rect -1829 -100 -1783 -88
rect -1571 88 -1525 100
rect -1571 -88 -1565 88
rect -1531 -88 -1525 88
rect -1571 -100 -1525 -88
rect -1313 88 -1267 100
rect -1313 -88 -1307 88
rect -1273 -88 -1267 88
rect -1313 -100 -1267 -88
rect -1055 88 -1009 100
rect -1055 -88 -1049 88
rect -1015 -88 -1009 88
rect -1055 -100 -1009 -88
rect -797 88 -751 100
rect -797 -88 -791 88
rect -757 -88 -751 88
rect -797 -100 -751 -88
rect -539 88 -493 100
rect -539 -88 -533 88
rect -499 -88 -493 88
rect -539 -100 -493 -88
rect -281 88 -235 100
rect -281 -88 -275 88
rect -241 -88 -235 88
rect -281 -100 -235 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 235 88 281 100
rect 235 -88 241 88
rect 275 -88 281 88
rect 235 -100 281 -88
rect 493 88 539 100
rect 493 -88 499 88
rect 533 -88 539 88
rect 493 -100 539 -88
rect 751 88 797 100
rect 751 -88 757 88
rect 791 -88 797 88
rect 751 -100 797 -88
rect 1009 88 1055 100
rect 1009 -88 1015 88
rect 1049 -88 1055 88
rect 1009 -100 1055 -88
rect 1267 88 1313 100
rect 1267 -88 1273 88
rect 1307 -88 1313 88
rect 1267 -100 1313 -88
rect 1525 88 1571 100
rect 1525 -88 1531 88
rect 1565 -88 1571 88
rect 1525 -100 1571 -88
rect 1783 88 1829 100
rect 1783 -88 1789 88
rect 1823 -88 1829 88
rect 1783 -100 1829 -88
rect -1731 -147 -1623 -141
rect -1731 -181 -1719 -147
rect -1635 -181 -1623 -147
rect -1731 -187 -1623 -181
rect -1473 -147 -1365 -141
rect -1473 -181 -1461 -147
rect -1377 -181 -1365 -147
rect -1473 -187 -1365 -181
rect -1215 -147 -1107 -141
rect -1215 -181 -1203 -147
rect -1119 -181 -1107 -147
rect -1215 -187 -1107 -181
rect -957 -147 -849 -141
rect -957 -181 -945 -147
rect -861 -181 -849 -147
rect -957 -187 -849 -181
rect -699 -147 -591 -141
rect -699 -181 -687 -147
rect -603 -181 -591 -147
rect -699 -187 -591 -181
rect -441 -147 -333 -141
rect -441 -181 -429 -147
rect -345 -181 -333 -147
rect -441 -187 -333 -181
rect -183 -147 -75 -141
rect -183 -181 -171 -147
rect -87 -181 -75 -147
rect -183 -187 -75 -181
rect 75 -147 183 -141
rect 75 -181 87 -147
rect 171 -181 183 -147
rect 75 -187 183 -181
rect 333 -147 441 -141
rect 333 -181 345 -147
rect 429 -181 441 -147
rect 333 -187 441 -181
rect 591 -147 699 -141
rect 591 -181 603 -147
rect 687 -181 699 -147
rect 591 -187 699 -181
rect 849 -147 957 -141
rect 849 -181 861 -147
rect 945 -181 957 -147
rect 849 -187 957 -181
rect 1107 -147 1215 -141
rect 1107 -181 1119 -147
rect 1203 -181 1215 -147
rect 1107 -187 1215 -181
rect 1365 -147 1473 -141
rect 1365 -181 1377 -147
rect 1461 -181 1473 -147
rect 1365 -187 1473 -181
rect 1623 -147 1731 -141
rect 1623 -181 1635 -147
rect 1719 -181 1731 -147
rect 1623 -187 1731 -181
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string parameters w 1 l 1 m 1 nf 14 diffcov 100 polycov 60 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
