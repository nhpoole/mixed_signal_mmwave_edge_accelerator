magic
tech sky130A
magscale 1 2
timestamp 1622597354
<< metal3 >>
rect -1250 1172 1249 1200
rect -1250 -1172 1165 1172
rect 1229 -1172 1249 1172
rect -1250 -1200 1249 -1172
<< via3 >>
rect 1165 -1172 1229 1172
<< mimcap >>
rect -1150 1060 1050 1100
rect -1150 -1060 -1110 1060
rect 1010 -1060 1050 1060
rect -1150 -1100 1050 -1060
<< mimcapcontact >>
rect -1110 -1060 1010 1060
<< metal4 >>
rect 1149 1172 1245 1188
rect -1111 1060 1011 1061
rect -1111 -1060 -1110 1060
rect 1010 -1060 1011 1060
rect -1111 -1061 1011 -1060
rect 1149 -1172 1165 1172
rect 1229 -1172 1245 1172
rect 1149 -1188 1245 -1172
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_1
string FIXED_BBOX -1250 -1200 1150 1200
string parameters w 11.00 l 11.00 val 250.36 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 0 tconnect 0 ccov 100
string library sky130
<< end >>
