magic
tech sky130A
magscale 1 2
timestamp 1624494425
<< metal1 >>
rect 1570 1130 1604 2256
rect 1646 1142 1674 2256
rect 4066 1130 4100 2256
rect 4142 1142 4170 2256
rect 6562 1130 6596 2256
rect 6638 1142 6666 2256
rect 9058 1130 9092 2256
rect 9134 1142 9162 2256
rect 11554 1130 11588 2256
rect 11630 1142 11658 2256
rect 14050 1130 14084 2256
rect 14126 1142 14154 2256
rect 16546 1130 16580 2256
rect 16622 1142 16650 2256
rect 19042 1130 19076 2256
rect 19118 1142 19146 2256
rect 21538 1130 21572 2256
rect 21614 1142 21642 2256
rect 24034 1130 24068 2256
rect 24110 1142 24138 2256
rect 26530 1130 26564 2256
rect 26606 1142 26634 2256
rect 29026 1130 29060 2256
rect 29102 1142 29130 2256
rect 31522 1130 31556 2256
rect 31598 1142 31626 2256
rect 34018 1130 34052 2256
rect 34094 1142 34122 2256
rect 36514 1130 36548 2256
rect 36590 1142 36618 2256
rect 39010 1130 39044 2256
rect 39086 1142 39114 2256
rect 41506 1130 41540 2256
rect 41582 1142 41610 2256
rect 44002 1130 44036 2256
rect 44078 1142 44106 2256
rect 46498 1130 46532 2256
rect 46574 1142 46602 2256
rect 48994 1130 49028 2256
rect 49070 1142 49098 2256
rect 51490 1130 51524 2256
rect 51566 1142 51594 2256
rect 53986 1130 54020 2256
rect 54062 1142 54090 2256
rect 56482 1130 56516 2256
rect 56558 1142 56586 2256
rect 58978 1130 59012 2256
rect 59054 1142 59082 2256
rect 61474 1130 61508 2256
rect 61550 1142 61578 2256
rect 63970 1130 64004 2256
rect 64046 1142 64074 2256
rect 66466 1130 66500 2256
rect 66542 1142 66570 2256
rect 68962 1130 68996 2256
rect 69038 1142 69066 2256
rect 71458 1130 71492 2256
rect 71534 1142 71562 2256
rect 73954 1130 73988 2256
rect 74030 1142 74058 2256
rect 76450 1130 76484 2256
rect 76526 1142 76554 2256
rect 78946 1130 78980 2256
rect 79022 1142 79050 2256
rect 1478 0 1524 254
rect 3974 0 4020 254
rect 6470 0 6516 254
rect 8966 0 9012 254
rect 11462 0 11508 254
rect 13958 0 14004 254
rect 16454 0 16500 254
rect 18950 0 18996 254
rect 21446 0 21492 254
rect 23942 0 23988 254
rect 26438 0 26484 254
rect 28934 0 28980 254
rect 31430 0 31476 254
rect 33926 0 33972 254
rect 36422 0 36468 254
rect 38918 0 38964 254
rect 41414 0 41460 254
rect 43910 0 43956 254
rect 46406 0 46452 254
rect 48902 0 48948 254
rect 51398 0 51444 254
rect 53894 0 53940 254
rect 56390 0 56436 254
rect 58886 0 58932 254
rect 61382 0 61428 254
rect 63878 0 63924 254
rect 66374 0 66420 254
rect 68870 0 68916 254
rect 71366 0 71412 254
rect 73862 0 73908 254
rect 76358 0 76404 254
rect 78854 0 78900 254
<< metal2 >>
rect 1469 2170 1525 2218
rect 3965 2170 4021 2218
rect 6461 2170 6517 2218
rect 8957 2170 9013 2218
rect 11453 2170 11509 2218
rect 13949 2170 14005 2218
rect 16445 2170 16501 2218
rect 18941 2170 18997 2218
rect 21437 2170 21493 2218
rect 23933 2170 23989 2218
rect 26429 2170 26485 2218
rect 28925 2170 28981 2218
rect 31421 2170 31477 2218
rect 33917 2170 33973 2218
rect 36413 2170 36469 2218
rect 38909 2170 38965 2218
rect 41405 2170 41461 2218
rect 43901 2170 43957 2218
rect 46397 2170 46453 2218
rect 48893 2170 48949 2218
rect 51389 2170 51445 2218
rect 53885 2170 53941 2218
rect 56381 2170 56437 2218
rect 58877 2170 58933 2218
rect 61373 2170 61429 2218
rect 63869 2170 63925 2218
rect 66365 2170 66421 2218
rect 68861 2170 68917 2218
rect 71357 2170 71413 2218
rect 73853 2170 73909 2218
rect 76349 2170 76405 2218
rect 78845 2170 78901 2218
rect 1797 2018 1853 2066
rect 4293 2018 4349 2066
rect 6789 2018 6845 2066
rect 9285 2018 9341 2066
rect 11781 2018 11837 2066
rect 14277 2018 14333 2066
rect 16773 2018 16829 2066
rect 19269 2018 19325 2066
rect 21765 2018 21821 2066
rect 24261 2018 24317 2066
rect 26757 2018 26813 2066
rect 29253 2018 29309 2066
rect 31749 2018 31805 2066
rect 34245 2018 34301 2066
rect 36741 2018 36797 2066
rect 39237 2018 39293 2066
rect 41733 2018 41789 2066
rect 44229 2018 44285 2066
rect 46725 2018 46781 2066
rect 49221 2018 49277 2066
rect 51717 2018 51773 2066
rect 54213 2018 54269 2066
rect 56709 2018 56765 2066
rect 59205 2018 59261 2066
rect 61701 2018 61757 2066
rect 64197 2018 64253 2066
rect 66693 2018 66749 2066
rect 69189 2018 69245 2066
rect 71685 2018 71741 2066
rect 74181 2018 74237 2066
rect 76677 2018 76733 2066
rect 79173 2018 79229 2066
rect 1715 1244 1771 1292
rect 4211 1244 4267 1292
rect 6707 1244 6763 1292
rect 9203 1244 9259 1292
rect 11699 1244 11755 1292
rect 14195 1244 14251 1292
rect 16691 1244 16747 1292
rect 19187 1244 19243 1292
rect 21683 1244 21739 1292
rect 24179 1244 24235 1292
rect 26675 1244 26731 1292
rect 29171 1244 29227 1292
rect 31667 1244 31723 1292
rect 34163 1244 34219 1292
rect 36659 1244 36715 1292
rect 39155 1244 39211 1292
rect 41651 1244 41707 1292
rect 44147 1244 44203 1292
rect 46643 1244 46699 1292
rect 49139 1244 49195 1292
rect 51635 1244 51691 1292
rect 54131 1244 54187 1292
rect 56627 1244 56683 1292
rect 59123 1244 59179 1292
rect 61619 1244 61675 1292
rect 64115 1244 64171 1292
rect 66611 1244 66667 1292
rect 69107 1244 69163 1292
rect 71603 1244 71659 1292
rect 74099 1244 74155 1292
rect 76595 1244 76651 1292
rect 79091 1244 79147 1292
rect 1727 406 1783 454
rect 4223 406 4279 454
rect 6719 406 6775 454
rect 9215 406 9271 454
rect 11711 406 11767 454
rect 14207 406 14263 454
rect 16703 406 16759 454
rect 19199 406 19255 454
rect 21695 406 21751 454
rect 24191 406 24247 454
rect 26687 406 26743 454
rect 29183 406 29239 454
rect 31679 406 31735 454
rect 34175 406 34231 454
rect 36671 406 36727 454
rect 39167 406 39223 454
rect 41663 406 41719 454
rect 44159 406 44215 454
rect 46655 406 46711 454
rect 49151 406 49207 454
rect 51647 406 51703 454
rect 54143 406 54199 454
rect 56639 406 56695 454
rect 59135 406 59191 454
rect 61631 406 61687 454
rect 64127 406 64183 454
rect 66623 406 66679 454
rect 69119 406 69175 454
rect 71615 406 71671 454
rect 74111 406 74167 454
rect 76607 406 76663 454
rect 79103 406 79159 454
rect 1727 84 1783 132
rect 4223 84 4279 132
rect 6719 84 6775 132
rect 9215 84 9271 132
rect 11711 84 11767 132
rect 14207 84 14263 132
rect 16703 84 16759 132
rect 19199 84 19255 132
rect 21695 84 21751 132
rect 24191 84 24247 132
rect 26687 84 26743 132
rect 29183 84 29239 132
rect 31679 84 31735 132
rect 34175 84 34231 132
rect 36671 84 36727 132
rect 39167 84 39223 132
rect 41663 84 41719 132
rect 44159 84 44215 132
rect 46655 84 46711 132
rect 49151 84 49207 132
rect 51647 84 51703 132
rect 54143 84 54199 132
rect 56639 84 56695 132
rect 59135 84 59191 132
rect 61631 84 61687 132
rect 64127 84 64183 132
rect 66623 84 66679 132
rect 69119 84 69175 132
rect 71615 84 71671 132
rect 74111 84 74167 132
rect 76607 84 76663 132
rect 79103 84 79159 132
<< metal3 >>
rect 0 2164 79250 2224
rect 1776 1993 1874 2091
rect 4272 1993 4370 2091
rect 6768 1993 6866 2091
rect 9264 1993 9362 2091
rect 11760 1993 11858 2091
rect 14256 1993 14354 2091
rect 16752 1993 16850 2091
rect 19248 1993 19346 2091
rect 21744 1993 21842 2091
rect 24240 1993 24338 2091
rect 26736 1993 26834 2091
rect 29232 1993 29330 2091
rect 31728 1993 31826 2091
rect 34224 1993 34322 2091
rect 36720 1993 36818 2091
rect 39216 1993 39314 2091
rect 41712 1993 41810 2091
rect 44208 1993 44306 2091
rect 46704 1993 46802 2091
rect 49200 1993 49298 2091
rect 51696 1993 51794 2091
rect 54192 1993 54290 2091
rect 56688 1993 56786 2091
rect 59184 1993 59282 2091
rect 61680 1993 61778 2091
rect 64176 1993 64274 2091
rect 66672 1993 66770 2091
rect 69168 1993 69266 2091
rect 71664 1993 71762 2091
rect 74160 1993 74258 2091
rect 76656 1993 76754 2091
rect 79152 1993 79250 2091
rect 1694 1219 1792 1317
rect 4190 1219 4288 1317
rect 6686 1219 6784 1317
rect 9182 1219 9280 1317
rect 11678 1219 11776 1317
rect 14174 1219 14272 1317
rect 16670 1219 16768 1317
rect 19166 1219 19264 1317
rect 21662 1219 21760 1317
rect 24158 1219 24256 1317
rect 26654 1219 26752 1317
rect 29150 1219 29248 1317
rect 31646 1219 31744 1317
rect 34142 1219 34240 1317
rect 36638 1219 36736 1317
rect 39134 1219 39232 1317
rect 41630 1219 41728 1317
rect 44126 1219 44224 1317
rect 46622 1219 46720 1317
rect 49118 1219 49216 1317
rect 51614 1219 51712 1317
rect 54110 1219 54208 1317
rect 56606 1219 56704 1317
rect 59102 1219 59200 1317
rect 61598 1219 61696 1317
rect 64094 1219 64192 1317
rect 66590 1219 66688 1317
rect 69086 1219 69184 1317
rect 71582 1219 71680 1317
rect 74078 1219 74176 1317
rect 76574 1219 76672 1317
rect 79070 1219 79168 1317
rect 1706 381 1804 479
rect 4202 381 4300 479
rect 6698 381 6796 479
rect 9194 381 9292 479
rect 11690 381 11788 479
rect 14186 381 14284 479
rect 16682 381 16780 479
rect 19178 381 19276 479
rect 21674 381 21772 479
rect 24170 381 24268 479
rect 26666 381 26764 479
rect 29162 381 29260 479
rect 31658 381 31756 479
rect 34154 381 34252 479
rect 36650 381 36748 479
rect 39146 381 39244 479
rect 41642 381 41740 479
rect 44138 381 44236 479
rect 46634 381 46732 479
rect 49130 381 49228 479
rect 51626 381 51724 479
rect 54122 381 54220 479
rect 56618 381 56716 479
rect 59114 381 59212 479
rect 61610 381 61708 479
rect 64106 381 64204 479
rect 66602 381 66700 479
rect 69098 381 69196 479
rect 71594 381 71692 479
rect 74090 381 74188 479
rect 76586 381 76684 479
rect 79082 381 79180 479
rect 1706 59 1804 157
rect 4202 59 4300 157
rect 6698 59 6796 157
rect 9194 59 9292 157
rect 11690 59 11788 157
rect 14186 59 14284 157
rect 16682 59 16780 157
rect 19178 59 19276 157
rect 21674 59 21772 157
rect 24170 59 24268 157
rect 26666 59 26764 157
rect 29162 59 29260 157
rect 31658 59 31756 157
rect 34154 59 34252 157
rect 36650 59 36748 157
rect 39146 59 39244 157
rect 41642 59 41740 157
rect 44138 59 44236 157
rect 46634 59 46732 157
rect 49130 59 49228 157
rect 51626 59 51724 157
rect 54122 59 54220 157
rect 56618 59 56716 157
rect 59114 59 59212 157
rect 61610 59 61708 157
rect 64106 59 64204 157
rect 66602 59 66700 157
rect 69098 59 69196 157
rect 71594 59 71692 157
rect 74090 59 74188 157
rect 76586 59 76684 157
rect 79082 59 79180 157
use contact_9  contact_9_156
timestamp 1624494425
transform 1 0 1722 0 1 393
box 0 0 66 74
use contact_8  contact_8_156
timestamp 1624494425
transform 1 0 1723 0 1 398
box 0 0 64 64
use contact_9  contact_9_158
timestamp 1624494425
transform 1 0 1722 0 1 71
box 0 0 66 74
use contact_8  contact_8_158
timestamp 1624494425
transform 1 0 1723 0 1 76
box 0 0 64 64
use contact_9  contact_9_31
timestamp 1624494425
transform 1 0 1464 0 1 2157
box 0 0 66 74
use contact_8  contact_8_31
timestamp 1624494425
transform 1 0 1465 0 1 2162
box 0 0 64 64
use contact_9  contact_9_157
timestamp 1624494425
transform 1 0 1710 0 1 1231
box 0 0 66 74
use contact_8  contact_8_157
timestamp 1624494425
transform 1 0 1711 0 1 1236
box 0 0 64 64
use contact_9  contact_9_159
timestamp 1624494425
transform 1 0 1792 0 1 2005
box 0 0 66 74
use contact_8  contact_8_159
timestamp 1624494425
transform 1 0 1793 0 1 2010
box 0 0 64 64
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_31
timestamp 1624494425
transform 1 0 1374 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_30
timestamp 1624494425
transform 1 0 3870 0 1 0
box -541 0 937 2256
use contact_9  contact_9_152
timestamp 1624494425
transform 1 0 4218 0 1 393
box 0 0 66 74
use contact_8  contact_8_152
timestamp 1624494425
transform 1 0 4219 0 1 398
box 0 0 64 64
use contact_9  contact_9_154
timestamp 1624494425
transform 1 0 4218 0 1 71
box 0 0 66 74
use contact_8  contact_8_154
timestamp 1624494425
transform 1 0 4219 0 1 76
box 0 0 64 64
use contact_9  contact_9_153
timestamp 1624494425
transform 1 0 4206 0 1 1231
box 0 0 66 74
use contact_8  contact_8_153
timestamp 1624494425
transform 1 0 4207 0 1 1236
box 0 0 64 64
use contact_9  contact_9_30
timestamp 1624494425
transform 1 0 3960 0 1 2157
box 0 0 66 74
use contact_8  contact_8_30
timestamp 1624494425
transform 1 0 3961 0 1 2162
box 0 0 64 64
use contact_9  contact_9_155
timestamp 1624494425
transform 1 0 4288 0 1 2005
box 0 0 66 74
use contact_8  contact_8_155
timestamp 1624494425
transform 1 0 4289 0 1 2010
box 0 0 64 64
use contact_8  contact_8_150
timestamp 1624494425
transform 1 0 6715 0 1 76
box 0 0 64 64
use contact_9  contact_9_150
timestamp 1624494425
transform 1 0 6714 0 1 71
box 0 0 66 74
use contact_8  contact_8_149
timestamp 1624494425
transform 1 0 6703 0 1 1236
box 0 0 64 64
use contact_9  contact_9_149
timestamp 1624494425
transform 1 0 6702 0 1 1231
box 0 0 66 74
use contact_8  contact_8_148
timestamp 1624494425
transform 1 0 6715 0 1 398
box 0 0 64 64
use contact_9  contact_9_148
timestamp 1624494425
transform 1 0 6714 0 1 393
box 0 0 66 74
use contact_8  contact_8_29
timestamp 1624494425
transform 1 0 6457 0 1 2162
box 0 0 64 64
use contact_9  contact_9_29
timestamp 1624494425
transform 1 0 6456 0 1 2157
box 0 0 66 74
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_29
timestamp 1624494425
transform 1 0 6366 0 1 0
box -541 0 937 2256
use contact_8  contact_8_151
timestamp 1624494425
transform 1 0 6785 0 1 2010
box 0 0 64 64
use contact_9  contact_9_151
timestamp 1624494425
transform 1 0 6784 0 1 2005
box 0 0 66 74
use contact_9  contact_9_144
timestamp 1624494425
transform 1 0 9210 0 1 393
box 0 0 66 74
use contact_8  contact_8_144
timestamp 1624494425
transform 1 0 9211 0 1 398
box 0 0 64 64
use contact_9  contact_9_146
timestamp 1624494425
transform 1 0 9210 0 1 71
box 0 0 66 74
use contact_8  contact_8_146
timestamp 1624494425
transform 1 0 9211 0 1 76
box 0 0 64 64
use contact_9  contact_9_28
timestamp 1624494425
transform 1 0 8952 0 1 2157
box 0 0 66 74
use contact_8  contact_8_28
timestamp 1624494425
transform 1 0 8953 0 1 2162
box 0 0 64 64
use contact_9  contact_9_145
timestamp 1624494425
transform 1 0 9198 0 1 1231
box 0 0 66 74
use contact_8  contact_8_145
timestamp 1624494425
transform 1 0 9199 0 1 1236
box 0 0 64 64
use contact_9  contact_9_147
timestamp 1624494425
transform 1 0 9280 0 1 2005
box 0 0 66 74
use contact_8  contact_8_147
timestamp 1624494425
transform 1 0 9281 0 1 2010
box 0 0 64 64
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_28
timestamp 1624494425
transform 1 0 8862 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_27
timestamp 1624494425
transform 1 0 11358 0 1 0
box -541 0 937 2256
use contact_9  contact_9_140
timestamp 1624494425
transform 1 0 11706 0 1 393
box 0 0 66 74
use contact_8  contact_8_140
timestamp 1624494425
transform 1 0 11707 0 1 398
box 0 0 64 64
use contact_9  contact_9_142
timestamp 1624494425
transform 1 0 11706 0 1 71
box 0 0 66 74
use contact_8  contact_8_142
timestamp 1624494425
transform 1 0 11707 0 1 76
box 0 0 64 64
use contact_9  contact_9_141
timestamp 1624494425
transform 1 0 11694 0 1 1231
box 0 0 66 74
use contact_8  contact_8_141
timestamp 1624494425
transform 1 0 11695 0 1 1236
box 0 0 64 64
use contact_9  contact_9_27
timestamp 1624494425
transform 1 0 11448 0 1 2157
box 0 0 66 74
use contact_8  contact_8_27
timestamp 1624494425
transform 1 0 11449 0 1 2162
box 0 0 64 64
use contact_9  contact_9_143
timestamp 1624494425
transform 1 0 11776 0 1 2005
box 0 0 66 74
use contact_8  contact_8_143
timestamp 1624494425
transform 1 0 11777 0 1 2010
box 0 0 64 64
use contact_8  contact_8_26
timestamp 1624494425
transform 1 0 13945 0 1 2162
box 0 0 64 64
use contact_9  contact_9_26
timestamp 1624494425
transform 1 0 13944 0 1 2157
box 0 0 66 74
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_26
timestamp 1624494425
transform 1 0 13854 0 1 0
box -541 0 937 2256
use contact_8  contact_8_139
timestamp 1624494425
transform 1 0 14273 0 1 2010
box 0 0 64 64
use contact_9  contact_9_139
timestamp 1624494425
transform 1 0 14272 0 1 2005
box 0 0 66 74
use contact_8  contact_8_138
timestamp 1624494425
transform 1 0 14203 0 1 76
box 0 0 64 64
use contact_9  contact_9_138
timestamp 1624494425
transform 1 0 14202 0 1 71
box 0 0 66 74
use contact_8  contact_8_137
timestamp 1624494425
transform 1 0 14191 0 1 1236
box 0 0 64 64
use contact_9  contact_9_137
timestamp 1624494425
transform 1 0 14190 0 1 1231
box 0 0 66 74
use contact_8  contact_8_136
timestamp 1624494425
transform 1 0 14203 0 1 398
box 0 0 64 64
use contact_9  contact_9_136
timestamp 1624494425
transform 1 0 14202 0 1 393
box 0 0 66 74
use contact_9  contact_9_132
timestamp 1624494425
transform 1 0 16698 0 1 393
box 0 0 66 74
use contact_8  contact_8_132
timestamp 1624494425
transform 1 0 16699 0 1 398
box 0 0 64 64
use contact_9  contact_9_134
timestamp 1624494425
transform 1 0 16698 0 1 71
box 0 0 66 74
use contact_8  contact_8_134
timestamp 1624494425
transform 1 0 16699 0 1 76
box 0 0 64 64
use contact_9  contact_9_25
timestamp 1624494425
transform 1 0 16440 0 1 2157
box 0 0 66 74
use contact_8  contact_8_25
timestamp 1624494425
transform 1 0 16441 0 1 2162
box 0 0 64 64
use contact_9  contact_9_133
timestamp 1624494425
transform 1 0 16686 0 1 1231
box 0 0 66 74
use contact_8  contact_8_133
timestamp 1624494425
transform 1 0 16687 0 1 1236
box 0 0 64 64
use contact_9  contact_9_135
timestamp 1624494425
transform 1 0 16768 0 1 2005
box 0 0 66 74
use contact_8  contact_8_135
timestamp 1624494425
transform 1 0 16769 0 1 2010
box 0 0 64 64
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_25
timestamp 1624494425
transform 1 0 16350 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_24
timestamp 1624494425
transform 1 0 18846 0 1 0
box -541 0 937 2256
use contact_9  contact_9_128
timestamp 1624494425
transform 1 0 19194 0 1 393
box 0 0 66 74
use contact_8  contact_8_128
timestamp 1624494425
transform 1 0 19195 0 1 398
box 0 0 64 64
use contact_9  contact_9_130
timestamp 1624494425
transform 1 0 19194 0 1 71
box 0 0 66 74
use contact_8  contact_8_130
timestamp 1624494425
transform 1 0 19195 0 1 76
box 0 0 64 64
use contact_9  contact_9_129
timestamp 1624494425
transform 1 0 19182 0 1 1231
box 0 0 66 74
use contact_8  contact_8_129
timestamp 1624494425
transform 1 0 19183 0 1 1236
box 0 0 64 64
use contact_9  contact_9_24
timestamp 1624494425
transform 1 0 18936 0 1 2157
box 0 0 66 74
use contact_8  contact_8_24
timestamp 1624494425
transform 1 0 18937 0 1 2162
box 0 0 64 64
use contact_9  contact_9_131
timestamp 1624494425
transform 1 0 19264 0 1 2005
box 0 0 66 74
use contact_8  contact_8_131
timestamp 1624494425
transform 1 0 19265 0 1 2010
box 0 0 64 64
use contact_8  contact_8_23
timestamp 1624494425
transform 1 0 21433 0 1 2162
box 0 0 64 64
use contact_9  contact_9_23
timestamp 1624494425
transform 1 0 21432 0 1 2157
box 0 0 66 74
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_23
timestamp 1624494425
transform 1 0 21342 0 1 0
box -541 0 937 2256
use contact_8  contact_8_127
timestamp 1624494425
transform 1 0 21761 0 1 2010
box 0 0 64 64
use contact_9  contact_9_127
timestamp 1624494425
transform 1 0 21760 0 1 2005
box 0 0 66 74
use contact_8  contact_8_126
timestamp 1624494425
transform 1 0 21691 0 1 76
box 0 0 64 64
use contact_9  contact_9_126
timestamp 1624494425
transform 1 0 21690 0 1 71
box 0 0 66 74
use contact_8  contact_8_125
timestamp 1624494425
transform 1 0 21679 0 1 1236
box 0 0 64 64
use contact_9  contact_9_125
timestamp 1624494425
transform 1 0 21678 0 1 1231
box 0 0 66 74
use contact_8  contact_8_124
timestamp 1624494425
transform 1 0 21691 0 1 398
box 0 0 64 64
use contact_9  contact_9_124
timestamp 1624494425
transform 1 0 21690 0 1 393
box 0 0 66 74
use contact_9  contact_9_120
timestamp 1624494425
transform 1 0 24186 0 1 393
box 0 0 66 74
use contact_8  contact_8_120
timestamp 1624494425
transform 1 0 24187 0 1 398
box 0 0 64 64
use contact_9  contact_9_122
timestamp 1624494425
transform 1 0 24186 0 1 71
box 0 0 66 74
use contact_8  contact_8_122
timestamp 1624494425
transform 1 0 24187 0 1 76
box 0 0 64 64
use contact_9  contact_9_22
timestamp 1624494425
transform 1 0 23928 0 1 2157
box 0 0 66 74
use contact_8  contact_8_22
timestamp 1624494425
transform 1 0 23929 0 1 2162
box 0 0 64 64
use contact_9  contact_9_121
timestamp 1624494425
transform 1 0 24174 0 1 1231
box 0 0 66 74
use contact_8  contact_8_121
timestamp 1624494425
transform 1 0 24175 0 1 1236
box 0 0 64 64
use contact_9  contact_9_123
timestamp 1624494425
transform 1 0 24256 0 1 2005
box 0 0 66 74
use contact_8  contact_8_123
timestamp 1624494425
transform 1 0 24257 0 1 2010
box 0 0 64 64
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_22
timestamp 1624494425
transform 1 0 23838 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_21
timestamp 1624494425
transform 1 0 26334 0 1 0
box -541 0 937 2256
use contact_9  contact_9_116
timestamp 1624494425
transform 1 0 26682 0 1 393
box 0 0 66 74
use contact_8  contact_8_116
timestamp 1624494425
transform 1 0 26683 0 1 398
box 0 0 64 64
use contact_9  contact_9_118
timestamp 1624494425
transform 1 0 26682 0 1 71
box 0 0 66 74
use contact_8  contact_8_118
timestamp 1624494425
transform 1 0 26683 0 1 76
box 0 0 64 64
use contact_9  contact_9_117
timestamp 1624494425
transform 1 0 26670 0 1 1231
box 0 0 66 74
use contact_8  contact_8_117
timestamp 1624494425
transform 1 0 26671 0 1 1236
box 0 0 64 64
use contact_9  contact_9_21
timestamp 1624494425
transform 1 0 26424 0 1 2157
box 0 0 66 74
use contact_8  contact_8_21
timestamp 1624494425
transform 1 0 26425 0 1 2162
box 0 0 64 64
use contact_9  contact_9_119
timestamp 1624494425
transform 1 0 26752 0 1 2005
box 0 0 66 74
use contact_8  contact_8_119
timestamp 1624494425
transform 1 0 26753 0 1 2010
box 0 0 64 64
use contact_8  contact_8_20
timestamp 1624494425
transform 1 0 28921 0 1 2162
box 0 0 64 64
use contact_9  contact_9_20
timestamp 1624494425
transform 1 0 28920 0 1 2157
box 0 0 66 74
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_20
timestamp 1624494425
transform 1 0 28830 0 1 0
box -541 0 937 2256
use contact_8  contact_8_115
timestamp 1624494425
transform 1 0 29249 0 1 2010
box 0 0 64 64
use contact_9  contact_9_115
timestamp 1624494425
transform 1 0 29248 0 1 2005
box 0 0 66 74
use contact_8  contact_8_114
timestamp 1624494425
transform 1 0 29179 0 1 76
box 0 0 64 64
use contact_9  contact_9_114
timestamp 1624494425
transform 1 0 29178 0 1 71
box 0 0 66 74
use contact_8  contact_8_113
timestamp 1624494425
transform 1 0 29167 0 1 1236
box 0 0 64 64
use contact_9  contact_9_113
timestamp 1624494425
transform 1 0 29166 0 1 1231
box 0 0 66 74
use contact_8  contact_8_112
timestamp 1624494425
transform 1 0 29179 0 1 398
box 0 0 64 64
use contact_9  contact_9_112
timestamp 1624494425
transform 1 0 29178 0 1 393
box 0 0 66 74
use contact_9  contact_9_108
timestamp 1624494425
transform 1 0 31674 0 1 393
box 0 0 66 74
use contact_8  contact_8_108
timestamp 1624494425
transform 1 0 31675 0 1 398
box 0 0 64 64
use contact_9  contact_9_110
timestamp 1624494425
transform 1 0 31674 0 1 71
box 0 0 66 74
use contact_8  contact_8_110
timestamp 1624494425
transform 1 0 31675 0 1 76
box 0 0 64 64
use contact_9  contact_9_19
timestamp 1624494425
transform 1 0 31416 0 1 2157
box 0 0 66 74
use contact_8  contact_8_19
timestamp 1624494425
transform 1 0 31417 0 1 2162
box 0 0 64 64
use contact_9  contact_9_109
timestamp 1624494425
transform 1 0 31662 0 1 1231
box 0 0 66 74
use contact_8  contact_8_109
timestamp 1624494425
transform 1 0 31663 0 1 1236
box 0 0 64 64
use contact_9  contact_9_111
timestamp 1624494425
transform 1 0 31744 0 1 2005
box 0 0 66 74
use contact_8  contact_8_111
timestamp 1624494425
transform 1 0 31745 0 1 2010
box 0 0 64 64
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_19
timestamp 1624494425
transform 1 0 31326 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_18
timestamp 1624494425
transform 1 0 33822 0 1 0
box -541 0 937 2256
use contact_9  contact_9_104
timestamp 1624494425
transform 1 0 34170 0 1 393
box 0 0 66 74
use contact_8  contact_8_104
timestamp 1624494425
transform 1 0 34171 0 1 398
box 0 0 64 64
use contact_9  contact_9_106
timestamp 1624494425
transform 1 0 34170 0 1 71
box 0 0 66 74
use contact_8  contact_8_106
timestamp 1624494425
transform 1 0 34171 0 1 76
box 0 0 64 64
use contact_9  contact_9_105
timestamp 1624494425
transform 1 0 34158 0 1 1231
box 0 0 66 74
use contact_8  contact_8_105
timestamp 1624494425
transform 1 0 34159 0 1 1236
box 0 0 64 64
use contact_9  contact_9_18
timestamp 1624494425
transform 1 0 33912 0 1 2157
box 0 0 66 74
use contact_8  contact_8_18
timestamp 1624494425
transform 1 0 33913 0 1 2162
box 0 0 64 64
use contact_9  contact_9_107
timestamp 1624494425
transform 1 0 34240 0 1 2005
box 0 0 66 74
use contact_8  contact_8_107
timestamp 1624494425
transform 1 0 34241 0 1 2010
box 0 0 64 64
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_17
timestamp 1624494425
transform 1 0 36318 0 1 0
box -541 0 937 2256
use contact_9  contact_9_100
timestamp 1624494425
transform 1 0 36666 0 1 393
box 0 0 66 74
use contact_8  contact_8_100
timestamp 1624494425
transform 1 0 36667 0 1 398
box 0 0 64 64
use contact_9  contact_9_102
timestamp 1624494425
transform 1 0 36666 0 1 71
box 0 0 66 74
use contact_8  contact_8_102
timestamp 1624494425
transform 1 0 36667 0 1 76
box 0 0 64 64
use contact_9  contact_9_101
timestamp 1624494425
transform 1 0 36654 0 1 1231
box 0 0 66 74
use contact_8  contact_8_101
timestamp 1624494425
transform 1 0 36655 0 1 1236
box 0 0 64 64
use contact_9  contact_9_17
timestamp 1624494425
transform 1 0 36408 0 1 2157
box 0 0 66 74
use contact_8  contact_8_17
timestamp 1624494425
transform 1 0 36409 0 1 2162
box 0 0 64 64
use contact_9  contact_9_103
timestamp 1624494425
transform 1 0 36736 0 1 2005
box 0 0 66 74
use contact_8  contact_8_103
timestamp 1624494425
transform 1 0 36737 0 1 2010
box 0 0 64 64
use contact_9  contact_9_96
timestamp 1624494425
transform 1 0 39162 0 1 393
box 0 0 66 74
use contact_8  contact_8_96
timestamp 1624494425
transform 1 0 39163 0 1 398
box 0 0 64 64
use contact_9  contact_9_98
timestamp 1624494425
transform 1 0 39162 0 1 71
box 0 0 66 74
use contact_8  contact_8_98
timestamp 1624494425
transform 1 0 39163 0 1 76
box 0 0 64 64
use contact_9  contact_9_16
timestamp 1624494425
transform 1 0 38904 0 1 2157
box 0 0 66 74
use contact_8  contact_8_16
timestamp 1624494425
transform 1 0 38905 0 1 2162
box 0 0 64 64
use contact_9  contact_9_97
timestamp 1624494425
transform 1 0 39150 0 1 1231
box 0 0 66 74
use contact_8  contact_8_97
timestamp 1624494425
transform 1 0 39151 0 1 1236
box 0 0 64 64
use contact_9  contact_9_99
timestamp 1624494425
transform 1 0 39232 0 1 2005
box 0 0 66 74
use contact_8  contact_8_99
timestamp 1624494425
transform 1 0 39233 0 1 2010
box 0 0 64 64
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_16
timestamp 1624494425
transform 1 0 38814 0 1 0
box -541 0 937 2256
use contact_9  contact_9_92
timestamp 1624494425
transform 1 0 41658 0 1 393
box 0 0 66 74
use contact_8  contact_8_92
timestamp 1624494425
transform 1 0 41659 0 1 398
box 0 0 64 64
use contact_9  contact_9_94
timestamp 1624494425
transform 1 0 41658 0 1 71
box 0 0 66 74
use contact_8  contact_8_94
timestamp 1624494425
transform 1 0 41659 0 1 76
box 0 0 64 64
use contact_9  contact_9_15
timestamp 1624494425
transform 1 0 41400 0 1 2157
box 0 0 66 74
use contact_8  contact_8_15
timestamp 1624494425
transform 1 0 41401 0 1 2162
box 0 0 64 64
use contact_9  contact_9_93
timestamp 1624494425
transform 1 0 41646 0 1 1231
box 0 0 66 74
use contact_8  contact_8_93
timestamp 1624494425
transform 1 0 41647 0 1 1236
box 0 0 64 64
use contact_9  contact_9_95
timestamp 1624494425
transform 1 0 41728 0 1 2005
box 0 0 66 74
use contact_8  contact_8_95
timestamp 1624494425
transform 1 0 41729 0 1 2010
box 0 0 64 64
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_15
timestamp 1624494425
transform 1 0 41310 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_14
timestamp 1624494425
transform 1 0 43806 0 1 0
box -541 0 937 2256
use contact_9  contact_9_88
timestamp 1624494425
transform 1 0 44154 0 1 393
box 0 0 66 74
use contact_8  contact_8_88
timestamp 1624494425
transform 1 0 44155 0 1 398
box 0 0 64 64
use contact_9  contact_9_90
timestamp 1624494425
transform 1 0 44154 0 1 71
box 0 0 66 74
use contact_8  contact_8_90
timestamp 1624494425
transform 1 0 44155 0 1 76
box 0 0 64 64
use contact_9  contact_9_89
timestamp 1624494425
transform 1 0 44142 0 1 1231
box 0 0 66 74
use contact_8  contact_8_89
timestamp 1624494425
transform 1 0 44143 0 1 1236
box 0 0 64 64
use contact_9  contact_9_14
timestamp 1624494425
transform 1 0 43896 0 1 2157
box 0 0 66 74
use contact_8  contact_8_14
timestamp 1624494425
transform 1 0 43897 0 1 2162
box 0 0 64 64
use contact_9  contact_9_91
timestamp 1624494425
transform 1 0 44224 0 1 2005
box 0 0 66 74
use contact_8  contact_8_91
timestamp 1624494425
transform 1 0 44225 0 1 2010
box 0 0 64 64
use contact_8  contact_8_86
timestamp 1624494425
transform 1 0 46651 0 1 76
box 0 0 64 64
use contact_9  contact_9_86
timestamp 1624494425
transform 1 0 46650 0 1 71
box 0 0 66 74
use contact_8  contact_8_85
timestamp 1624494425
transform 1 0 46639 0 1 1236
box 0 0 64 64
use contact_9  contact_9_85
timestamp 1624494425
transform 1 0 46638 0 1 1231
box 0 0 66 74
use contact_8  contact_8_84
timestamp 1624494425
transform 1 0 46651 0 1 398
box 0 0 64 64
use contact_9  contact_9_84
timestamp 1624494425
transform 1 0 46650 0 1 393
box 0 0 66 74
use contact_8  contact_8_13
timestamp 1624494425
transform 1 0 46393 0 1 2162
box 0 0 64 64
use contact_9  contact_9_13
timestamp 1624494425
transform 1 0 46392 0 1 2157
box 0 0 66 74
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_13
timestamp 1624494425
transform 1 0 46302 0 1 0
box -541 0 937 2256
use contact_8  contact_8_87
timestamp 1624494425
transform 1 0 46721 0 1 2010
box 0 0 64 64
use contact_9  contact_9_87
timestamp 1624494425
transform 1 0 46720 0 1 2005
box 0 0 66 74
use contact_9  contact_9_80
timestamp 1624494425
transform 1 0 49146 0 1 393
box 0 0 66 74
use contact_8  contact_8_80
timestamp 1624494425
transform 1 0 49147 0 1 398
box 0 0 64 64
use contact_9  contact_9_82
timestamp 1624494425
transform 1 0 49146 0 1 71
box 0 0 66 74
use contact_8  contact_8_82
timestamp 1624494425
transform 1 0 49147 0 1 76
box 0 0 64 64
use contact_9  contact_9_12
timestamp 1624494425
transform 1 0 48888 0 1 2157
box 0 0 66 74
use contact_8  contact_8_12
timestamp 1624494425
transform 1 0 48889 0 1 2162
box 0 0 64 64
use contact_9  contact_9_81
timestamp 1624494425
transform 1 0 49134 0 1 1231
box 0 0 66 74
use contact_8  contact_8_81
timestamp 1624494425
transform 1 0 49135 0 1 1236
box 0 0 64 64
use contact_9  contact_9_83
timestamp 1624494425
transform 1 0 49216 0 1 2005
box 0 0 66 74
use contact_8  contact_8_83
timestamp 1624494425
transform 1 0 49217 0 1 2010
box 0 0 64 64
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_12
timestamp 1624494425
transform 1 0 48798 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_11
timestamp 1624494425
transform 1 0 51294 0 1 0
box -541 0 937 2256
use contact_9  contact_9_76
timestamp 1624494425
transform 1 0 51642 0 1 393
box 0 0 66 74
use contact_8  contact_8_76
timestamp 1624494425
transform 1 0 51643 0 1 398
box 0 0 64 64
use contact_9  contact_9_78
timestamp 1624494425
transform 1 0 51642 0 1 71
box 0 0 66 74
use contact_8  contact_8_78
timestamp 1624494425
transform 1 0 51643 0 1 76
box 0 0 64 64
use contact_9  contact_9_77
timestamp 1624494425
transform 1 0 51630 0 1 1231
box 0 0 66 74
use contact_8  contact_8_77
timestamp 1624494425
transform 1 0 51631 0 1 1236
box 0 0 64 64
use contact_9  contact_9_11
timestamp 1624494425
transform 1 0 51384 0 1 2157
box 0 0 66 74
use contact_8  contact_8_11
timestamp 1624494425
transform 1 0 51385 0 1 2162
box 0 0 64 64
use contact_9  contact_9_79
timestamp 1624494425
transform 1 0 51712 0 1 2005
box 0 0 66 74
use contact_8  contact_8_79
timestamp 1624494425
transform 1 0 51713 0 1 2010
box 0 0 64 64
use contact_8  contact_8_10
timestamp 1624494425
transform 1 0 53881 0 1 2162
box 0 0 64 64
use contact_9  contact_9_10
timestamp 1624494425
transform 1 0 53880 0 1 2157
box 0 0 66 74
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_10
timestamp 1624494425
transform 1 0 53790 0 1 0
box -541 0 937 2256
use contact_8  contact_8_75
timestamp 1624494425
transform 1 0 54209 0 1 2010
box 0 0 64 64
use contact_9  contact_9_75
timestamp 1624494425
transform 1 0 54208 0 1 2005
box 0 0 66 74
use contact_8  contact_8_74
timestamp 1624494425
transform 1 0 54139 0 1 76
box 0 0 64 64
use contact_9  contact_9_74
timestamp 1624494425
transform 1 0 54138 0 1 71
box 0 0 66 74
use contact_8  contact_8_73
timestamp 1624494425
transform 1 0 54127 0 1 1236
box 0 0 64 64
use contact_9  contact_9_73
timestamp 1624494425
transform 1 0 54126 0 1 1231
box 0 0 66 74
use contact_8  contact_8_72
timestamp 1624494425
transform 1 0 54139 0 1 398
box 0 0 64 64
use contact_9  contact_9_72
timestamp 1624494425
transform 1 0 54138 0 1 393
box 0 0 66 74
use contact_9  contact_9_68
timestamp 1624494425
transform 1 0 56634 0 1 393
box 0 0 66 74
use contact_8  contact_8_68
timestamp 1624494425
transform 1 0 56635 0 1 398
box 0 0 64 64
use contact_9  contact_9_70
timestamp 1624494425
transform 1 0 56634 0 1 71
box 0 0 66 74
use contact_8  contact_8_70
timestamp 1624494425
transform 1 0 56635 0 1 76
box 0 0 64 64
use contact_9  contact_9_9
timestamp 1624494425
transform 1 0 56376 0 1 2157
box 0 0 66 74
use contact_8  contact_8_9
timestamp 1624494425
transform 1 0 56377 0 1 2162
box 0 0 64 64
use contact_9  contact_9_69
timestamp 1624494425
transform 1 0 56622 0 1 1231
box 0 0 66 74
use contact_8  contact_8_69
timestamp 1624494425
transform 1 0 56623 0 1 1236
box 0 0 64 64
use contact_9  contact_9_71
timestamp 1624494425
transform 1 0 56704 0 1 2005
box 0 0 66 74
use contact_8  contact_8_71
timestamp 1624494425
transform 1 0 56705 0 1 2010
box 0 0 64 64
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_9
timestamp 1624494425
transform 1 0 56286 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_8
timestamp 1624494425
transform 1 0 58782 0 1 0
box -541 0 937 2256
use contact_9  contact_9_64
timestamp 1624494425
transform 1 0 59130 0 1 393
box 0 0 66 74
use contact_8  contact_8_64
timestamp 1624494425
transform 1 0 59131 0 1 398
box 0 0 64 64
use contact_9  contact_9_66
timestamp 1624494425
transform 1 0 59130 0 1 71
box 0 0 66 74
use contact_8  contact_8_66
timestamp 1624494425
transform 1 0 59131 0 1 76
box 0 0 64 64
use contact_9  contact_9_65
timestamp 1624494425
transform 1 0 59118 0 1 1231
box 0 0 66 74
use contact_8  contact_8_65
timestamp 1624494425
transform 1 0 59119 0 1 1236
box 0 0 64 64
use contact_9  contact_9_8
timestamp 1624494425
transform 1 0 58872 0 1 2157
box 0 0 66 74
use contact_8  contact_8_8
timestamp 1624494425
transform 1 0 58873 0 1 2162
box 0 0 64 64
use contact_9  contact_9_67
timestamp 1624494425
transform 1 0 59200 0 1 2005
box 0 0 66 74
use contact_8  contact_8_67
timestamp 1624494425
transform 1 0 59201 0 1 2010
box 0 0 64 64
use contact_8  contact_8_7
timestamp 1624494425
transform 1 0 61369 0 1 2162
box 0 0 64 64
use contact_9  contact_9_7
timestamp 1624494425
transform 1 0 61368 0 1 2157
box 0 0 66 74
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_7
timestamp 1624494425
transform 1 0 61278 0 1 0
box -541 0 937 2256
use contact_8  contact_8_63
timestamp 1624494425
transform 1 0 61697 0 1 2010
box 0 0 64 64
use contact_9  contact_9_63
timestamp 1624494425
transform 1 0 61696 0 1 2005
box 0 0 66 74
use contact_8  contact_8_62
timestamp 1624494425
transform 1 0 61627 0 1 76
box 0 0 64 64
use contact_9  contact_9_62
timestamp 1624494425
transform 1 0 61626 0 1 71
box 0 0 66 74
use contact_8  contact_8_61
timestamp 1624494425
transform 1 0 61615 0 1 1236
box 0 0 64 64
use contact_9  contact_9_61
timestamp 1624494425
transform 1 0 61614 0 1 1231
box 0 0 66 74
use contact_8  contact_8_60
timestamp 1624494425
transform 1 0 61627 0 1 398
box 0 0 64 64
use contact_9  contact_9_60
timestamp 1624494425
transform 1 0 61626 0 1 393
box 0 0 66 74
use contact_9  contact_9_56
timestamp 1624494425
transform 1 0 64122 0 1 393
box 0 0 66 74
use contact_8  contact_8_56
timestamp 1624494425
transform 1 0 64123 0 1 398
box 0 0 64 64
use contact_9  contact_9_58
timestamp 1624494425
transform 1 0 64122 0 1 71
box 0 0 66 74
use contact_8  contact_8_58
timestamp 1624494425
transform 1 0 64123 0 1 76
box 0 0 64 64
use contact_9  contact_9_6
timestamp 1624494425
transform 1 0 63864 0 1 2157
box 0 0 66 74
use contact_8  contact_8_6
timestamp 1624494425
transform 1 0 63865 0 1 2162
box 0 0 64 64
use contact_9  contact_9_57
timestamp 1624494425
transform 1 0 64110 0 1 1231
box 0 0 66 74
use contact_8  contact_8_57
timestamp 1624494425
transform 1 0 64111 0 1 1236
box 0 0 64 64
use contact_9  contact_9_59
timestamp 1624494425
transform 1 0 64192 0 1 2005
box 0 0 66 74
use contact_8  contact_8_59
timestamp 1624494425
transform 1 0 64193 0 1 2010
box 0 0 64 64
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_6
timestamp 1624494425
transform 1 0 63774 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_5
timestamp 1624494425
transform 1 0 66270 0 1 0
box -541 0 937 2256
use contact_9  contact_9_52
timestamp 1624494425
transform 1 0 66618 0 1 393
box 0 0 66 74
use contact_8  contact_8_52
timestamp 1624494425
transform 1 0 66619 0 1 398
box 0 0 64 64
use contact_9  contact_9_54
timestamp 1624494425
transform 1 0 66618 0 1 71
box 0 0 66 74
use contact_8  contact_8_54
timestamp 1624494425
transform 1 0 66619 0 1 76
box 0 0 64 64
use contact_9  contact_9_53
timestamp 1624494425
transform 1 0 66606 0 1 1231
box 0 0 66 74
use contact_8  contact_8_53
timestamp 1624494425
transform 1 0 66607 0 1 1236
box 0 0 64 64
use contact_9  contact_9_5
timestamp 1624494425
transform 1 0 66360 0 1 2157
box 0 0 66 74
use contact_8  contact_8_5
timestamp 1624494425
transform 1 0 66361 0 1 2162
box 0 0 64 64
use contact_9  contact_9_55
timestamp 1624494425
transform 1 0 66688 0 1 2005
box 0 0 66 74
use contact_8  contact_8_55
timestamp 1624494425
transform 1 0 66689 0 1 2010
box 0 0 64 64
use contact_8  contact_8_4
timestamp 1624494425
transform 1 0 68857 0 1 2162
box 0 0 64 64
use contact_9  contact_9_4
timestamp 1624494425
transform 1 0 68856 0 1 2157
box 0 0 66 74
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_4
timestamp 1624494425
transform 1 0 68766 0 1 0
box -541 0 937 2256
use contact_8  contact_8_51
timestamp 1624494425
transform 1 0 69185 0 1 2010
box 0 0 64 64
use contact_9  contact_9_51
timestamp 1624494425
transform 1 0 69184 0 1 2005
box 0 0 66 74
use contact_8  contact_8_50
timestamp 1624494425
transform 1 0 69115 0 1 76
box 0 0 64 64
use contact_9  contact_9_50
timestamp 1624494425
transform 1 0 69114 0 1 71
box 0 0 66 74
use contact_8  contact_8_49
timestamp 1624494425
transform 1 0 69103 0 1 1236
box 0 0 64 64
use contact_9  contact_9_49
timestamp 1624494425
transform 1 0 69102 0 1 1231
box 0 0 66 74
use contact_8  contact_8_48
timestamp 1624494425
transform 1 0 69115 0 1 398
box 0 0 64 64
use contact_9  contact_9_48
timestamp 1624494425
transform 1 0 69114 0 1 393
box 0 0 66 74
use contact_9  contact_9_44
timestamp 1624494425
transform 1 0 71610 0 1 393
box 0 0 66 74
use contact_8  contact_8_44
timestamp 1624494425
transform 1 0 71611 0 1 398
box 0 0 64 64
use contact_9  contact_9_46
timestamp 1624494425
transform 1 0 71610 0 1 71
box 0 0 66 74
use contact_8  contact_8_46
timestamp 1624494425
transform 1 0 71611 0 1 76
box 0 0 64 64
use contact_9  contact_9_3
timestamp 1624494425
transform 1 0 71352 0 1 2157
box 0 0 66 74
use contact_8  contact_8_3
timestamp 1624494425
transform 1 0 71353 0 1 2162
box 0 0 64 64
use contact_9  contact_9_45
timestamp 1624494425
transform 1 0 71598 0 1 1231
box 0 0 66 74
use contact_8  contact_8_45
timestamp 1624494425
transform 1 0 71599 0 1 1236
box 0 0 64 64
use contact_9  contact_9_47
timestamp 1624494425
transform 1 0 71680 0 1 2005
box 0 0 66 74
use contact_8  contact_8_47
timestamp 1624494425
transform 1 0 71681 0 1 2010
box 0 0 64 64
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_3
timestamp 1624494425
transform 1 0 71262 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_2
timestamp 1624494425
transform 1 0 73758 0 1 0
box -541 0 937 2256
use contact_9  contact_9_40
timestamp 1624494425
transform 1 0 74106 0 1 393
box 0 0 66 74
use contact_8  contact_8_40
timestamp 1624494425
transform 1 0 74107 0 1 398
box 0 0 64 64
use contact_9  contact_9_42
timestamp 1624494425
transform 1 0 74106 0 1 71
box 0 0 66 74
use contact_8  contact_8_42
timestamp 1624494425
transform 1 0 74107 0 1 76
box 0 0 64 64
use contact_9  contact_9_41
timestamp 1624494425
transform 1 0 74094 0 1 1231
box 0 0 66 74
use contact_8  contact_8_41
timestamp 1624494425
transform 1 0 74095 0 1 1236
box 0 0 64 64
use contact_9  contact_9_2
timestamp 1624494425
transform 1 0 73848 0 1 2157
box 0 0 66 74
use contact_8  contact_8_2
timestamp 1624494425
transform 1 0 73849 0 1 2162
box 0 0 64 64
use contact_9  contact_9_43
timestamp 1624494425
transform 1 0 74176 0 1 2005
box 0 0 66 74
use contact_8  contact_8_43
timestamp 1624494425
transform 1 0 74177 0 1 2010
box 0 0 64 64
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_1
timestamp 1624494425
transform 1 0 76254 0 1 0
box -541 0 937 2256
use contact_9  contact_9_36
timestamp 1624494425
transform 1 0 76602 0 1 393
box 0 0 66 74
use contact_8  contact_8_36
timestamp 1624494425
transform 1 0 76603 0 1 398
box 0 0 64 64
use contact_9  contact_9_38
timestamp 1624494425
transform 1 0 76602 0 1 71
box 0 0 66 74
use contact_8  contact_8_38
timestamp 1624494425
transform 1 0 76603 0 1 76
box 0 0 64 64
use contact_9  contact_9_37
timestamp 1624494425
transform 1 0 76590 0 1 1231
box 0 0 66 74
use contact_8  contact_8_37
timestamp 1624494425
transform 1 0 76591 0 1 1236
box 0 0 64 64
use contact_9  contact_9_1
timestamp 1624494425
transform 1 0 76344 0 1 2157
box 0 0 66 74
use contact_8  contact_8_1
timestamp 1624494425
transform 1 0 76345 0 1 2162
box 0 0 64 64
use contact_9  contact_9_39
timestamp 1624494425
transform 1 0 76672 0 1 2005
box 0 0 66 74
use contact_8  contact_8_39
timestamp 1624494425
transform 1 0 76673 0 1 2010
box 0 0 64 64
use contact_9  contact_9_32
timestamp 1624494425
transform 1 0 79098 0 1 393
box 0 0 66 74
use contact_8  contact_8_32
timestamp 1624494425
transform 1 0 79099 0 1 398
box 0 0 64 64
use contact_9  contact_9_34
timestamp 1624494425
transform 1 0 79098 0 1 71
box 0 0 66 74
use contact_8  contact_8_34
timestamp 1624494425
transform 1 0 79099 0 1 76
box 0 0 64 64
use contact_9  contact_9_0
timestamp 1624494425
transform 1 0 78840 0 1 2157
box 0 0 66 74
use contact_8  contact_8_0
timestamp 1624494425
transform 1 0 78841 0 1 2162
box 0 0 64 64
use contact_9  contact_9_33
timestamp 1624494425
transform 1 0 79086 0 1 1231
box 0 0 66 74
use contact_8  contact_8_33
timestamp 1624494425
transform 1 0 79087 0 1 1236
box 0 0 64 64
use contact_9  contact_9_35
timestamp 1624494425
transform 1 0 79168 0 1 2005
box 0 0 66 74
use contact_8  contact_8_35
timestamp 1624494425
transform 1 0 79169 0 1 2010
box 0 0 64 64
use sky130_fd_bd_sram__openram_sense_amp  sky130_fd_bd_sram__openram_sense_amp_0
timestamp 1624494425
transform 1 0 78750 0 1 0
box -541 0 937 2256
<< labels >>
rlabel metal3 s 79152 1993 79250 2091 4 gnd
rlabel metal3 s 21744 1993 21842 2091 4 gnd
rlabel metal3 s 49200 1993 49298 2091 4 gnd
rlabel metal3 s 74090 59 74188 157 4 gnd
rlabel metal3 s 4272 1993 4370 2091 4 gnd
rlabel metal3 s 31658 59 31756 157 4 gnd
rlabel metal3 s 6768 1993 6866 2091 4 gnd
rlabel metal3 s 51626 59 51724 157 4 gnd
rlabel metal3 s 9264 1993 9362 2091 4 gnd
rlabel metal3 s 14186 59 14284 157 4 gnd
rlabel metal3 s 24240 1993 24338 2091 4 gnd
rlabel metal3 s 14256 1993 14354 2091 4 gnd
rlabel metal3 s 34154 59 34252 157 4 gnd
rlabel metal3 s 39146 59 39244 157 4 gnd
rlabel metal3 s 1776 1993 1874 2091 4 gnd
rlabel metal3 s 61680 1993 61778 2091 4 gnd
rlabel metal3 s 66602 59 66700 157 4 gnd
rlabel metal3 s 71664 1993 71762 2091 4 gnd
rlabel metal3 s 26666 59 26764 157 4 gnd
rlabel metal3 s 41712 1993 41810 2091 4 gnd
rlabel metal3 s 44208 1993 44306 2091 4 gnd
rlabel metal3 s 36720 1993 36818 2091 4 gnd
rlabel metal3 s 71594 59 71692 157 4 gnd
rlabel metal3 s 19178 59 19276 157 4 gnd
rlabel metal3 s 66672 1993 66770 2091 4 gnd
rlabel metal3 s 79082 59 79180 157 4 gnd
rlabel metal3 s 51696 1993 51794 2091 4 gnd
rlabel metal3 s 21674 59 21772 157 4 gnd
rlabel metal3 s 64106 59 64204 157 4 gnd
rlabel metal3 s 19248 1993 19346 2091 4 gnd
rlabel metal3 s 76586 59 76684 157 4 gnd
rlabel metal3 s 64176 1993 64274 2091 4 gnd
rlabel metal3 s 76656 1993 76754 2091 4 gnd
rlabel metal3 s 11760 1993 11858 2091 4 gnd
rlabel metal3 s 39216 1993 39314 2091 4 gnd
rlabel metal3 s 41642 59 41740 157 4 gnd
rlabel metal3 s 1706 59 1804 157 4 gnd
rlabel metal3 s 46704 1993 46802 2091 4 gnd
rlabel metal3 s 16752 1993 16850 2091 4 gnd
rlabel metal3 s 54122 59 54220 157 4 gnd
rlabel metal3 s 31728 1993 31826 2091 4 gnd
rlabel metal3 s 34224 1993 34322 2091 4 gnd
rlabel metal3 s 69098 59 69196 157 4 gnd
rlabel metal3 s 11690 59 11788 157 4 gnd
rlabel metal3 s 29162 59 29260 157 4 gnd
rlabel metal3 s 46634 59 46732 157 4 gnd
rlabel metal3 s 24170 59 24268 157 4 gnd
rlabel metal3 s 56618 59 56716 157 4 gnd
rlabel metal3 s 69168 1993 69266 2091 4 gnd
rlabel metal3 s 59114 59 59212 157 4 gnd
rlabel metal3 s 4202 59 4300 157 4 gnd
rlabel metal3 s 9194 59 9292 157 4 gnd
rlabel metal3 s 36650 59 36748 157 4 gnd
rlabel metal3 s 44138 59 44236 157 4 gnd
rlabel metal3 s 54192 1993 54290 2091 4 gnd
rlabel metal3 s 6698 59 6796 157 4 gnd
rlabel metal3 s 61610 59 61708 157 4 gnd
rlabel metal3 s 16682 59 16780 157 4 gnd
rlabel metal3 s 26736 1993 26834 2091 4 gnd
rlabel metal3 s 29232 1993 29330 2091 4 gnd
rlabel metal3 s 49130 59 49228 157 4 gnd
rlabel metal3 s 59184 1993 59282 2091 4 gnd
rlabel metal3 s 74160 1993 74258 2091 4 gnd
rlabel metal3 s 56688 1993 56786 2091 4 gnd
rlabel metal3 s 41630 1219 41728 1317 4 vdd
rlabel metal3 s 79070 1219 79168 1317 4 vdd
rlabel metal3 s 71582 1219 71680 1317 4 vdd
rlabel metal3 s 54122 381 54220 479 4 vdd
rlabel metal3 s 11678 1219 11776 1317 4 vdd
rlabel metal3 s 11690 381 11788 479 4 vdd
rlabel metal3 s 74090 381 74188 479 4 vdd
rlabel metal3 s 19178 381 19276 479 4 vdd
rlabel metal3 s 21674 381 21772 479 4 vdd
rlabel metal3 s 21662 1219 21760 1317 4 vdd
rlabel metal3 s 61598 1219 61696 1317 4 vdd
rlabel metal3 s 44138 381 44236 479 4 vdd
rlabel metal3 s 46634 381 46732 479 4 vdd
rlabel metal3 s 29150 1219 29248 1317 4 vdd
rlabel metal3 s 51626 381 51724 479 4 vdd
rlabel metal3 s 4190 1219 4288 1317 4 vdd
rlabel metal3 s 1706 381 1804 479 4 vdd
rlabel metal3 s 6698 381 6796 479 4 vdd
rlabel metal3 s 9194 381 9292 479 4 vdd
rlabel metal3 s 26654 1219 26752 1317 4 vdd
rlabel metal3 s 16682 381 16780 479 4 vdd
rlabel metal3 s 6686 1219 6784 1317 4 vdd
rlabel metal3 s 34142 1219 34240 1317 4 vdd
rlabel metal3 s 51614 1219 51712 1317 4 vdd
rlabel metal3 s 64106 381 64204 479 4 vdd
rlabel metal3 s 74078 1219 74176 1317 4 vdd
rlabel metal3 s 4202 381 4300 479 4 vdd
rlabel metal3 s 1694 1219 1792 1317 4 vdd
rlabel metal3 s 36638 1219 36736 1317 4 vdd
rlabel metal3 s 39146 381 39244 479 4 vdd
rlabel metal3 s 31658 381 31756 479 4 vdd
rlabel metal3 s 56618 381 56716 479 4 vdd
rlabel metal3 s 46622 1219 46720 1317 4 vdd
rlabel metal3 s 64094 1219 64192 1317 4 vdd
rlabel metal3 s 49118 1219 49216 1317 4 vdd
rlabel metal3 s 61610 381 61708 479 4 vdd
rlabel metal3 s 59102 1219 59200 1317 4 vdd
rlabel metal3 s 59114 381 59212 479 4 vdd
rlabel metal3 s 54110 1219 54208 1317 4 vdd
rlabel metal3 s 9182 1219 9280 1317 4 vdd
rlabel metal3 s 76586 381 76684 479 4 vdd
rlabel metal3 s 24158 1219 24256 1317 4 vdd
rlabel metal3 s 56606 1219 56704 1317 4 vdd
rlabel metal3 s 79082 381 79180 479 4 vdd
rlabel metal3 s 71594 381 71692 479 4 vdd
rlabel metal3 s 41642 381 41740 479 4 vdd
rlabel metal3 s 66590 1219 66688 1317 4 vdd
rlabel metal3 s 49130 381 49228 479 4 vdd
rlabel metal3 s 26666 381 26764 479 4 vdd
rlabel metal3 s 76574 1219 76672 1317 4 vdd
rlabel metal3 s 31646 1219 31744 1317 4 vdd
rlabel metal3 s 34154 381 34252 479 4 vdd
rlabel metal3 s 24170 381 24268 479 4 vdd
rlabel metal3 s 39134 1219 39232 1317 4 vdd
rlabel metal3 s 14186 381 14284 479 4 vdd
rlabel metal3 s 44126 1219 44224 1317 4 vdd
rlabel metal3 s 69086 1219 69184 1317 4 vdd
rlabel metal3 s 14174 1219 14272 1317 4 vdd
rlabel metal3 s 66602 381 66700 479 4 vdd
rlabel metal3 s 36650 381 36748 479 4 vdd
rlabel metal3 s 69098 381 69196 479 4 vdd
rlabel metal3 s 16670 1219 16768 1317 4 vdd
rlabel metal3 s 29162 381 29260 479 4 vdd
rlabel metal3 s 19166 1219 19264 1317 4 vdd
rlabel metal1 s 1570 1130 1604 2256 4 bl_0
rlabel metal1 s 1646 1142 1674 2256 4 br_0
rlabel metal1 s 1478 0 1524 254 4 data_0
rlabel metal1 s 4066 1130 4100 2256 4 bl_1
rlabel metal1 s 4142 1142 4170 2256 4 br_1
rlabel metal1 s 3974 0 4020 254 4 data_1
rlabel metal1 s 6562 1130 6596 2256 4 bl_2
rlabel metal1 s 6638 1142 6666 2256 4 br_2
rlabel metal1 s 6470 0 6516 254 4 data_2
rlabel metal1 s 9058 1130 9092 2256 4 bl_3
rlabel metal1 s 9134 1142 9162 2256 4 br_3
rlabel metal1 s 8966 0 9012 254 4 data_3
rlabel metal1 s 11554 1130 11588 2256 4 bl_4
rlabel metal1 s 11630 1142 11658 2256 4 br_4
rlabel metal1 s 11462 0 11508 254 4 data_4
rlabel metal1 s 14050 1130 14084 2256 4 bl_5
rlabel metal1 s 14126 1142 14154 2256 4 br_5
rlabel metal1 s 13958 0 14004 254 4 data_5
rlabel metal1 s 16546 1130 16580 2256 4 bl_6
rlabel metal1 s 16622 1142 16650 2256 4 br_6
rlabel metal1 s 16454 0 16500 254 4 data_6
rlabel metal1 s 19042 1130 19076 2256 4 bl_7
rlabel metal1 s 19118 1142 19146 2256 4 br_7
rlabel metal1 s 18950 0 18996 254 4 data_7
rlabel metal1 s 21538 1130 21572 2256 4 bl_8
rlabel metal1 s 21614 1142 21642 2256 4 br_8
rlabel metal1 s 21446 0 21492 254 4 data_8
rlabel metal1 s 24034 1130 24068 2256 4 bl_9
rlabel metal1 s 24110 1142 24138 2256 4 br_9
rlabel metal1 s 23942 0 23988 254 4 data_9
rlabel metal1 s 26530 1130 26564 2256 4 bl_10
rlabel metal1 s 26606 1142 26634 2256 4 br_10
rlabel metal1 s 26438 0 26484 254 4 data_10
rlabel metal1 s 29026 1130 29060 2256 4 bl_11
rlabel metal1 s 29102 1142 29130 2256 4 br_11
rlabel metal1 s 28934 0 28980 254 4 data_11
rlabel metal1 s 31522 1130 31556 2256 4 bl_12
rlabel metal1 s 31598 1142 31626 2256 4 br_12
rlabel metal1 s 31430 0 31476 254 4 data_12
rlabel metal1 s 34018 1130 34052 2256 4 bl_13
rlabel metal1 s 34094 1142 34122 2256 4 br_13
rlabel metal1 s 33926 0 33972 254 4 data_13
rlabel metal1 s 36514 1130 36548 2256 4 bl_14
rlabel metal1 s 36590 1142 36618 2256 4 br_14
rlabel metal1 s 36422 0 36468 254 4 data_14
rlabel metal1 s 39010 1130 39044 2256 4 bl_15
rlabel metal1 s 39086 1142 39114 2256 4 br_15
rlabel metal1 s 38918 0 38964 254 4 data_15
rlabel metal1 s 41506 1130 41540 2256 4 bl_16
rlabel metal1 s 41582 1142 41610 2256 4 br_16
rlabel metal1 s 41414 0 41460 254 4 data_16
rlabel metal1 s 44002 1130 44036 2256 4 bl_17
rlabel metal1 s 44078 1142 44106 2256 4 br_17
rlabel metal1 s 43910 0 43956 254 4 data_17
rlabel metal1 s 46498 1130 46532 2256 4 bl_18
rlabel metal1 s 46574 1142 46602 2256 4 br_18
rlabel metal1 s 46406 0 46452 254 4 data_18
rlabel metal1 s 48994 1130 49028 2256 4 bl_19
rlabel metal1 s 49070 1142 49098 2256 4 br_19
rlabel metal1 s 48902 0 48948 254 4 data_19
rlabel metal1 s 51490 1130 51524 2256 4 bl_20
rlabel metal1 s 51566 1142 51594 2256 4 br_20
rlabel metal1 s 51398 0 51444 254 4 data_20
rlabel metal1 s 53986 1130 54020 2256 4 bl_21
rlabel metal1 s 54062 1142 54090 2256 4 br_21
rlabel metal1 s 53894 0 53940 254 4 data_21
rlabel metal1 s 56482 1130 56516 2256 4 bl_22
rlabel metal1 s 56558 1142 56586 2256 4 br_22
rlabel metal1 s 56390 0 56436 254 4 data_22
rlabel metal1 s 58978 1130 59012 2256 4 bl_23
rlabel metal1 s 59054 1142 59082 2256 4 br_23
rlabel metal1 s 58886 0 58932 254 4 data_23
rlabel metal1 s 61474 1130 61508 2256 4 bl_24
rlabel metal1 s 61550 1142 61578 2256 4 br_24
rlabel metal1 s 61382 0 61428 254 4 data_24
rlabel metal1 s 63970 1130 64004 2256 4 bl_25
rlabel metal1 s 64046 1142 64074 2256 4 br_25
rlabel metal1 s 63878 0 63924 254 4 data_25
rlabel metal1 s 66466 1130 66500 2256 4 bl_26
rlabel metal1 s 66542 1142 66570 2256 4 br_26
rlabel metal1 s 66374 0 66420 254 4 data_26
rlabel metal1 s 68962 1130 68996 2256 4 bl_27
rlabel metal1 s 69038 1142 69066 2256 4 br_27
rlabel metal1 s 68870 0 68916 254 4 data_27
rlabel metal1 s 71458 1130 71492 2256 4 bl_28
rlabel metal1 s 71534 1142 71562 2256 4 br_28
rlabel metal1 s 71366 0 71412 254 4 data_28
rlabel metal1 s 73954 1130 73988 2256 4 bl_29
rlabel metal1 s 74030 1142 74058 2256 4 br_29
rlabel metal1 s 73862 0 73908 254 4 data_29
rlabel metal1 s 76450 1130 76484 2256 4 bl_30
rlabel metal1 s 76526 1142 76554 2256 4 br_30
rlabel metal1 s 76358 0 76404 254 4 data_30
rlabel metal1 s 78946 1130 78980 2256 4 bl_31
rlabel metal1 s 79022 1142 79050 2256 4 br_31
rlabel metal1 s 78854 0 78900 254 4 data_31
rlabel metal3 s 0 2164 79250 2224 4 en
<< properties >>
string FIXED_BBOX 0 0 79250 2256
<< end >>
