magic
tech sky130A
timestamp 1626065694
<< checkpaint >>
rect -720 -720 720 720
<< metal4 >>
rect -90 59 90 90
rect -90 -59 -59 59
rect 59 -59 90 59
rect -90 -90 90 -59
<< via4 >>
rect -59 -59 59 59
<< metal5 >>
rect -90 59 90 90
rect -90 -59 -59 59
rect 59 -59 90 59
rect -90 -90 90 -59
<< end >>
