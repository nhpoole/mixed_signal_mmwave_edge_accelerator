magic
tech sky130A
magscale 1 2
timestamp 1624477805
<< error_p >>
rect -1355 -200 1355 200
<< nwell >>
rect -1355 -200 1355 200
<< pmos >>
rect -1261 -100 -1061 100
rect -1003 -100 -803 100
rect -745 -100 -545 100
rect -487 -100 -287 100
rect -229 -100 -29 100
rect 29 -100 229 100
rect 287 -100 487 100
rect 545 -100 745 100
rect 803 -100 1003 100
rect 1061 -100 1261 100
<< pdiff >>
rect -1319 88 -1261 100
rect -1319 -88 -1307 88
rect -1273 -88 -1261 88
rect -1319 -100 -1261 -88
rect -1061 88 -1003 100
rect -1061 -88 -1049 88
rect -1015 -88 -1003 88
rect -1061 -100 -1003 -88
rect -803 88 -745 100
rect -803 -88 -791 88
rect -757 -88 -745 88
rect -803 -100 -745 -88
rect -545 88 -487 100
rect -545 -88 -533 88
rect -499 -88 -487 88
rect -545 -100 -487 -88
rect -287 88 -229 100
rect -287 -88 -275 88
rect -241 -88 -229 88
rect -287 -100 -229 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 229 88 287 100
rect 229 -88 241 88
rect 275 -88 287 88
rect 229 -100 287 -88
rect 487 88 545 100
rect 487 -88 499 88
rect 533 -88 545 88
rect 487 -100 545 -88
rect 745 88 803 100
rect 745 -88 757 88
rect 791 -88 803 88
rect 745 -100 803 -88
rect 1003 88 1061 100
rect 1003 -88 1015 88
rect 1049 -88 1061 88
rect 1003 -100 1061 -88
rect 1261 88 1319 100
rect 1261 -88 1273 88
rect 1307 -88 1319 88
rect 1261 -100 1319 -88
<< pdiffc >>
rect -1307 -88 -1273 88
rect -1049 -88 -1015 88
rect -791 -88 -757 88
rect -533 -88 -499 88
rect -275 -88 -241 88
rect -17 -88 17 88
rect 241 -88 275 88
rect 499 -88 533 88
rect 757 -88 791 88
rect 1015 -88 1049 88
rect 1273 -88 1307 88
<< poly >>
rect -1261 181 -1061 197
rect -1261 147 -1245 181
rect -1077 147 -1061 181
rect -1261 100 -1061 147
rect -1003 181 -803 197
rect -1003 147 -987 181
rect -819 147 -803 181
rect -1003 100 -803 147
rect -745 181 -545 197
rect -745 147 -729 181
rect -561 147 -545 181
rect -745 100 -545 147
rect -487 181 -287 197
rect -487 147 -471 181
rect -303 147 -287 181
rect -487 100 -287 147
rect -229 181 -29 197
rect -229 147 -213 181
rect -45 147 -29 181
rect -229 100 -29 147
rect 29 181 229 197
rect 29 147 45 181
rect 213 147 229 181
rect 29 100 229 147
rect 287 181 487 197
rect 287 147 303 181
rect 471 147 487 181
rect 287 100 487 147
rect 545 181 745 197
rect 545 147 561 181
rect 729 147 745 181
rect 545 100 745 147
rect 803 181 1003 197
rect 803 147 819 181
rect 987 147 1003 181
rect 803 100 1003 147
rect 1061 181 1261 197
rect 1061 147 1077 181
rect 1245 147 1261 181
rect 1061 100 1261 147
rect -1261 -147 -1061 -100
rect -1261 -181 -1245 -147
rect -1077 -181 -1061 -147
rect -1261 -197 -1061 -181
rect -1003 -147 -803 -100
rect -1003 -181 -987 -147
rect -819 -181 -803 -147
rect -1003 -197 -803 -181
rect -745 -147 -545 -100
rect -745 -181 -729 -147
rect -561 -181 -545 -147
rect -745 -197 -545 -181
rect -487 -147 -287 -100
rect -487 -181 -471 -147
rect -303 -181 -287 -147
rect -487 -197 -287 -181
rect -229 -147 -29 -100
rect -229 -181 -213 -147
rect -45 -181 -29 -147
rect -229 -197 -29 -181
rect 29 -147 229 -100
rect 29 -181 45 -147
rect 213 -181 229 -147
rect 29 -197 229 -181
rect 287 -147 487 -100
rect 287 -181 303 -147
rect 471 -181 487 -147
rect 287 -197 487 -181
rect 545 -147 745 -100
rect 545 -181 561 -147
rect 729 -181 745 -147
rect 545 -197 745 -181
rect 803 -147 1003 -100
rect 803 -181 819 -147
rect 987 -181 1003 -147
rect 803 -197 1003 -181
rect 1061 -147 1261 -100
rect 1061 -181 1077 -147
rect 1245 -181 1261 -147
rect 1061 -197 1261 -181
<< polycont >>
rect -1245 147 -1077 181
rect -987 147 -819 181
rect -729 147 -561 181
rect -471 147 -303 181
rect -213 147 -45 181
rect 45 147 213 181
rect 303 147 471 181
rect 561 147 729 181
rect 819 147 987 181
rect 1077 147 1245 181
rect -1245 -181 -1077 -147
rect -987 -181 -819 -147
rect -729 -181 -561 -147
rect -471 -181 -303 -147
rect -213 -181 -45 -147
rect 45 -181 213 -147
rect 303 -181 471 -147
rect 561 -181 729 -147
rect 819 -181 987 -147
rect 1077 -181 1245 -147
<< locali >>
rect -1261 147 -1245 181
rect -1077 147 -1061 181
rect -1003 147 -987 181
rect -819 147 -803 181
rect -745 147 -729 181
rect -561 147 -545 181
rect -487 147 -471 181
rect -303 147 -287 181
rect -229 147 -213 181
rect -45 147 -29 181
rect 29 147 45 181
rect 213 147 229 181
rect 287 147 303 181
rect 471 147 487 181
rect 545 147 561 181
rect 729 147 745 181
rect 803 147 819 181
rect 987 147 1003 181
rect 1061 147 1077 181
rect 1245 147 1261 181
rect -1307 88 -1273 104
rect -1307 -104 -1273 -88
rect -1049 88 -1015 104
rect -1049 -104 -1015 -88
rect -791 88 -757 104
rect -791 -104 -757 -88
rect -533 88 -499 104
rect -533 -104 -499 -88
rect -275 88 -241 104
rect -275 -104 -241 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 241 88 275 104
rect 241 -104 275 -88
rect 499 88 533 104
rect 499 -104 533 -88
rect 757 88 791 104
rect 757 -104 791 -88
rect 1015 88 1049 104
rect 1015 -104 1049 -88
rect 1273 88 1307 104
rect 1273 -104 1307 -88
rect -1261 -181 -1245 -147
rect -1077 -181 -1061 -147
rect -1003 -181 -987 -147
rect -819 -181 -803 -147
rect -745 -181 -729 -147
rect -561 -181 -545 -147
rect -487 -181 -471 -147
rect -303 -181 -287 -147
rect -229 -181 -213 -147
rect -45 -181 -29 -147
rect 29 -181 45 -147
rect 213 -181 229 -147
rect 287 -181 303 -147
rect 471 -181 487 -147
rect 545 -181 561 -147
rect 729 -181 745 -147
rect 803 -181 819 -147
rect 987 -181 1003 -147
rect 1061 -181 1077 -147
rect 1245 -181 1261 -147
<< viali >>
rect -1203 147 -1119 181
rect -945 147 -861 181
rect -687 147 -603 181
rect -429 147 -345 181
rect -171 147 -87 181
rect 87 147 171 181
rect 345 147 429 181
rect 603 147 687 181
rect 861 147 945 181
rect 1119 147 1203 181
rect -1307 -88 -1273 88
rect -1049 -88 -1015 88
rect -791 -88 -757 88
rect -533 -88 -499 88
rect -275 -88 -241 88
rect -17 -88 17 88
rect 241 -88 275 88
rect 499 -88 533 88
rect 757 -88 791 88
rect 1015 -88 1049 88
rect 1273 -88 1307 88
rect -1203 -181 -1119 -147
rect -945 -181 -861 -147
rect -687 -181 -603 -147
rect -429 -181 -345 -147
rect -171 -181 -87 -147
rect 87 -181 171 -147
rect 345 -181 429 -147
rect 603 -181 687 -147
rect 861 -181 945 -147
rect 1119 -181 1203 -147
<< metal1 >>
rect -1215 181 -1107 187
rect -1215 147 -1203 181
rect -1119 147 -1107 181
rect -1215 141 -1107 147
rect -957 181 -849 187
rect -957 147 -945 181
rect -861 147 -849 181
rect -957 141 -849 147
rect -699 181 -591 187
rect -699 147 -687 181
rect -603 147 -591 181
rect -699 141 -591 147
rect -441 181 -333 187
rect -441 147 -429 181
rect -345 147 -333 181
rect -441 141 -333 147
rect -183 181 -75 187
rect -183 147 -171 181
rect -87 147 -75 181
rect -183 141 -75 147
rect 75 181 183 187
rect 75 147 87 181
rect 171 147 183 181
rect 75 141 183 147
rect 333 181 441 187
rect 333 147 345 181
rect 429 147 441 181
rect 333 141 441 147
rect 591 181 699 187
rect 591 147 603 181
rect 687 147 699 181
rect 591 141 699 147
rect 849 181 957 187
rect 849 147 861 181
rect 945 147 957 181
rect 849 141 957 147
rect 1107 181 1215 187
rect 1107 147 1119 181
rect 1203 147 1215 181
rect 1107 141 1215 147
rect -1313 88 -1267 100
rect -1313 -88 -1307 88
rect -1273 -88 -1267 88
rect -1313 -100 -1267 -88
rect -1055 88 -1009 100
rect -1055 -88 -1049 88
rect -1015 -88 -1009 88
rect -1055 -100 -1009 -88
rect -797 88 -751 100
rect -797 -88 -791 88
rect -757 -88 -751 88
rect -797 -100 -751 -88
rect -539 88 -493 100
rect -539 -88 -533 88
rect -499 -88 -493 88
rect -539 -100 -493 -88
rect -281 88 -235 100
rect -281 -88 -275 88
rect -241 -88 -235 88
rect -281 -100 -235 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 235 88 281 100
rect 235 -88 241 88
rect 275 -88 281 88
rect 235 -100 281 -88
rect 493 88 539 100
rect 493 -88 499 88
rect 533 -88 539 88
rect 493 -100 539 -88
rect 751 88 797 100
rect 751 -88 757 88
rect 791 -88 797 88
rect 751 -100 797 -88
rect 1009 88 1055 100
rect 1009 -88 1015 88
rect 1049 -88 1055 88
rect 1009 -100 1055 -88
rect 1267 88 1313 100
rect 1267 -88 1273 88
rect 1307 -88 1313 88
rect 1267 -100 1313 -88
rect -1215 -147 -1107 -141
rect -1215 -181 -1203 -147
rect -1119 -181 -1107 -147
rect -1215 -187 -1107 -181
rect -957 -147 -849 -141
rect -957 -181 -945 -147
rect -861 -181 -849 -147
rect -957 -187 -849 -181
rect -699 -147 -591 -141
rect -699 -181 -687 -147
rect -603 -181 -591 -147
rect -699 -187 -591 -181
rect -441 -147 -333 -141
rect -441 -181 -429 -147
rect -345 -181 -333 -147
rect -441 -187 -333 -181
rect -183 -147 -75 -141
rect -183 -181 -171 -147
rect -87 -181 -75 -147
rect -183 -187 -75 -181
rect 75 -147 183 -141
rect 75 -181 87 -147
rect 171 -181 183 -147
rect 75 -187 183 -181
rect 333 -147 441 -141
rect 333 -181 345 -147
rect 429 -181 441 -147
rect 333 -187 441 -181
rect 591 -147 699 -141
rect 591 -181 603 -147
rect 687 -181 699 -147
rect 591 -187 699 -181
rect 849 -147 957 -141
rect 849 -181 861 -147
rect 945 -181 957 -147
rect 849 -187 957 -181
rect 1107 -147 1215 -141
rect 1107 -181 1119 -147
rect 1203 -181 1215 -147
rect 1107 -187 1215 -181
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string parameters w 1 l 1 m 1 nf 10 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 60 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
