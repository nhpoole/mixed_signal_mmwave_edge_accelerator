magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect -2610 -1560 2492 1560
<< metal3 >>
rect -1350 -300 1232 300
<< mimcap >>
rect -1250 152 1150 200
rect -1250 -152 -1202 152
rect 1102 -152 1150 152
rect -1250 -200 1150 -152
<< mimcapcontact >>
rect -1202 -152 1102 152
<< metal4 >>
rect -1211 152 1111 161
rect -1211 -152 -1202 152
rect 1102 -152 1111 152
rect -1211 -161 1111 -152
<< properties >>
string FIXED_BBOX -1350 -300 1250 300
<< end >>
