* NGSPICE file created from biquad_gm_c_filter_flat.ext - technology: sky130A

.subckt biquad_gm_c_filter_flat VDD VSS vip vim ibiasn1 vocm vfiltp vfiltm vintp vintm
+ ibiasn2 ibiasn3 ibiasn4
X0 gm_c_stage_2/vcmcn2 vocm gm_c_stage_2/vcmn_tail2 VSS sky130_fd_pr__nfet_01v8 ad=1.74e+12p pd=1.374e+07u as=2.61e+12p ps=2.09e+07u w=2e+06u l=1e+06u
X1 gm_c_stage_1/vtail_diff vintm vintm VSS sky130_fd_pr__nfet_01v8_lvt ad=2.9e+12p pd=2.348e+07u as=4.64e+12p ps=3.664e+07u w=2e+06u l=1e+06u
X2 vintm vfiltp gm_c_stage_2/vtail_diff VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.9e+12p ps=2.348e+07u w=2e+06u l=1e+06u
X3 VDD gm_c_stage_3/vbiasp gm_c_stage_3/vbiasp VDD sky130_fd_pr__pfet_01v8 ad=9.28e+12p pd=8.256e+07u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X4 gm_c_stage_0/vcmcn gm_c_stage_0/vcmcn VDD VDD sky130_fd_pr__pfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
X5 gm_c_stage_1/vcmcn vintp gm_c_stage_1/vcmn_tail1 VSS sky130_fd_pr__nfet_01v8 ad=2.9e+12p pd=2.29e+07u as=2.61e+12p ps=2.09e+07u w=2e+06u l=1e+06u
X6 ibiasn1 ibiasn1 VSS VSS sky130_fd_pr__nfet_01v8 ad=1.74e+12p pd=1.548e+07u as=3.016e+13p ps=2.544e+08u w=1e+06u l=4e+06u
X7 ibiasn4 VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=1.74e+12p pd=1.548e+07u as=0p ps=0u w=1e+06u l=4e+06u
X8 VSS VSS gm_c_stage_2/vcmn_tail2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X9 gm_c_stage_1/vcmcn VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10 ibiasn3 ibiasn3 VSS VSS sky130_fd_pr__nfet_01v8 ad=1.74e+12p pd=1.548e+07u as=0p ps=0u w=1e+06u l=4e+06u
X11 gm_c_stage_2/vcmcn1 vocm gm_c_stage_2/vcmn_tail1 VSS sky130_fd_pr__nfet_01v8 ad=1.16e+12p pd=9.16e+06u as=2.61e+12p ps=2.09e+07u w=2e+06u l=1e+06u
X12 VSS ibiasn2 ibiasn2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.74e+12p ps=1.548e+07u w=1e+06u l=4e+06u
X13 gm_c_stage_2/vtail_diff vfiltm vintp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.06e+12p ps=3.206e+07u w=2e+06u l=1e+06u
X14 gm_c_stage_2/vtail_diff ibiasn4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X15 gm_c_stage_0/vcmn_tail1 vocm gm_c_stage_0/vcmcn1 VSS sky130_fd_pr__nfet_01v8 ad=2.61e+12p pd=2.09e+07u as=1.16e+12p ps=9.16e+06u w=2e+06u l=1e+06u
X16 vintm VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X17 VSS ibiasn4 gm_c_stage_2/vcmn_tail1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X18 gm_c_stage_2/vcmcn vintp gm_c_stage_2/vcmn_tail1 VSS sky130_fd_pr__nfet_01v8 ad=2.9e+12p pd=2.29e+07u as=0p ps=0u w=2e+06u l=1e+06u
X19 gm_c_stage_3/vcmn_tail1 vfiltp gm_c_stage_3/vcmcn VSS sky130_fd_pr__nfet_01v8 ad=2.61e+12p pd=2.09e+07u as=2.9e+12p ps=2.29e+07u w=2e+06u l=1e+06u
X20 VSS ibiasn3 ibiasn3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X21 gm_c_stage_0/vcmn_tail1 vintm gm_c_stage_0/vcmcn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+12p ps=2.29e+07u w=2e+06u l=1e+06u
X22 vintm vim gm_c_stage_0/vtail_diff VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.9e+12p ps=2.348e+07u w=2e+06u l=1e+06u
X23 gm_c_stage_3/vcmcn2 VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=1.74e+12p pd=1.374e+07u as=0p ps=0u w=2e+06u l=1e+06u
X24 ibiasn4 ibiasn4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X25 gm_c_stage_3/vtail_diff vintm vfiltm VSS sky130_fd_pr__nfet_01v8_lvt ad=2.9e+12p pd=2.348e+07u as=1.74e+12p ps=1.374e+07u w=2e+06u l=1e+06u
X26 VSS VSS gm_c_stage_2/vbiasp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=4e+06u
X27 VSS VSS gm_c_stage_3/vcmcn2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X28 gm_c_stage_3/vcmcn vfiltp gm_c_stage_3/vcmn_tail1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X29 gm_c_stage_1/vcmcn vintm gm_c_stage_1/vcmn_tail2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.61e+12p ps=2.09e+07u w=2e+06u l=1e+06u
X30 gm_c_stage_2/vbiasp VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
X31 VSS VSS ibiasn2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X32 VSS VSS gm_c_stage_3/vbiasp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=4e+06u
X33 gm_c_stage_1/vtail_diff vintp vintp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X34 gm_c_stage_0/vcmcn2 vocm gm_c_stage_0/vcmn_tail2 VSS sky130_fd_pr__nfet_01v8 ad=1.74e+12p pd=1.374e+07u as=2.61e+12p ps=2.09e+07u w=2e+06u l=1e+06u
X35 vfiltm VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X36 VDD gm_c_stage_2/vcmcn gm_c_stage_2/vcmc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X37 gm_c_stage_3/vcmcn2 vocm gm_c_stage_3/vcmn_tail2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.61e+12p ps=2.09e+07u w=2e+06u l=1e+06u
X38 VSS VSS gm_c_stage_0/vbiasp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=4e+06u
X39 gm_c_stage_1/vcmn_tail2 vocm gm_c_stage_1/vcmcn2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.74e+12p ps=1.374e+07u w=2e+06u l=1e+06u
X40 gm_c_stage_0/vcmn_tail2 vintp gm_c_stage_0/vcmcn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X41 gm_c_stage_0/vtail_diff ibiasn1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X42 VSS VSS ibiasn1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X43 gm_c_stage_3/vcmcn2 vocm gm_c_stage_3/vcmn_tail2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X44 VSS ibiasn4 ibiasn4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X45 gm_c_stage_1/vbiasp ibiasn2 VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=4e+06u
X46 VDD VDD gm_c_stage_1/vcmcn2 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X47 vintp vintp gm_c_stage_1/vtail_diff VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X48 VDD VDD vintp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=1e+06u
X49 ibiasn1 ibiasn1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X50 VDD VDD gm_c_stage_1/vcmcn VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X51 gm_c_stage_0/vcmcn vintp gm_c_stage_0/vcmn_tail2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X52 ibiasn1 ibiasn1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X53 gm_c_stage_3/vcmn_tail2 vfiltm gm_c_stage_3/vcmcn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X54 gm_c_stage_0/vcmcn1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
X55 gm_c_stage_0/vcmn_tail2 vocm gm_c_stage_0/vcmcn2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X56 VDD gm_c_stage_0/vbiasp gm_c_stage_0/vbiasp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X57 VDD VDD gm_c_stage_0/vcmcn VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X58 gm_c_stage_1/vcmcn gm_c_stage_1/vcmcn VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X59 gm_c_stage_0/vbiasp ibiasn1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X60 gm_c_stage_2/vcmcn2 vocm gm_c_stage_2/vcmn_tail2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X61 gm_c_stage_3/vtail_diff vintp vfiltp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.16e+12p ps=9.16e+06u w=2e+06u l=1e+06u
X62 gm_c_stage_3/vcmcn VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X63 VSS ibiasn3 ibiasn3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X64 VSS VSS ibiasn3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X65 VSS gm_c_stage_0/vcmc gm_c_stage_0/vcmc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=4e+06u
X66 gm_c_stage_2/vcmn_tail1 vocm gm_c_stage_2/vcmcn1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X67 gm_c_stage_2/vcmn_tail2 vintm gm_c_stage_2/vcmcn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X68 VSS ibiasn2 ibiasn2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X69 gm_c_stage_0/vtail_diff vip vintp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X70 VSS VSS vintp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X71 gm_c_stage_2/vcmcn vintm gm_c_stage_2/vcmn_tail2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X72 gm_c_stage_2/vcmn_tail1 VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X73 VDD VDD gm_c_stage_3/vcmcn2 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X74 vintp VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X75 vintp vintp gm_c_stage_1/vtail_diff VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X76 VDD VDD gm_c_stage_3/vcmcn VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X77 vintp vip gm_c_stage_0/vtail_diff VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X78 gm_c_stage_0/vcmn_tail2 ibiasn1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X79 gm_c_stage_2/vcmn_tail1 vintp gm_c_stage_2/vcmcn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X80 gm_c_stage_2/vcmn_tail2 ibiasn4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X81 VSS ibiasn1 ibiasn1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X82 VSS ibiasn2 gm_c_stage_1/vcmn_tail1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X83 gm_c_stage_0/vtail_diff vim vintm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X84 gm_c_stage_1/vcmc VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=4e+06u
X85 gm_c_stage_1/vcmn_tail2 vintm gm_c_stage_1/vcmcn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X86 gm_c_stage_0/vcmn_tail1 vintm gm_c_stage_0/vcmcn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X87 gm_c_stage_2/vbiasp ibiasn4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X88 gm_c_stage_1/vtail_diff vintm vintm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X89 vintp gm_c_stage_1/vbiasp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X90 gm_c_stage_3/vcmc VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=4e+06u
X91 gm_c_stage_0/vcmcn vintm gm_c_stage_0/vcmn_tail1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X92 gm_c_stage_1/vcmcn vintm gm_c_stage_1/vcmn_tail2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X93 VSS ibiasn1 ibiasn1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X94 VSS ibiasn4 ibiasn4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X95 ibiasn2 ibiasn2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X96 VDD VDD vintm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+11p ps=7.74e+06u w=1e+06u l=1e+06u
X97 gm_c_stage_3/vcmn_tail2 vocm gm_c_stage_3/vcmcn2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X98 gm_c_stage_0/vcmcn2 VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X99 VSS ibiasn1 gm_c_stage_0/vcmn_tail1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X100 VSS VSS gm_c_stage_1/vcmn_tail2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X101 VDD VDD vintm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X102 vfiltp vintp gm_c_stage_3/vtail_diff VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X103 VSS ibiasn1 ibiasn1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X104 ibiasn4 ibiasn4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X105 vfiltp vintp gm_c_stage_3/vtail_diff VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X106 VSS VSS gm_c_stage_1/vtail_diff VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X107 vintm gm_c_stage_0/vbiasp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X108 gm_c_stage_2/vcmcn1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
X109 VSS ibiasn3 gm_c_stage_3/vcmn_tail1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X110 vintm vintm gm_c_stage_1/vtail_diff VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X111 gm_c_stage_1/vcmn_tail1 VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X112 gm_c_stage_3/vcmn_tail2 ibiasn3 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X113 VDD gm_c_stage_0/vcmcn1 gm_c_stage_0/vcmcn1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X114 VDD gm_c_stage_2/vbiasp gm_c_stage_2/vbiasp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X115 VDD VDD gm_c_stage_2/vcmcn VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X116 gm_c_stage_2/vcmc VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=4e+06u
X117 ibiasn2 ibiasn2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X118 VDD gm_c_stage_1/vcmcn1 gm_c_stage_1/vcmcn1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X119 gm_c_stage_0/vcmc VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X120 gm_c_stage_3/vcmcn gm_c_stage_3/vcmcn VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X121 gm_c_stage_3/vtail_diff vintm vfiltm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X122 vintp gm_c_stage_0/vbiasp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X123 vfiltp gm_c_stage_3/vbiasp VDD VDD sky130_fd_pr__pfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
X124 gm_c_stage_3/vcmn_tail2 vocm gm_c_stage_3/vcmcn2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X125 VSS ibiasn1 ibiasn1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X126 VSS VSS gm_c_stage_2/vcmcn2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X127 VSS ibiasn4 ibiasn4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X128 gm_c_stage_1/vcmn_tail1 vocm gm_c_stage_1/vcmcn1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.16e+12p ps=9.16e+06u w=2e+06u l=1e+06u
X129 VDD VDD gm_c_stage_0/vcmcn2 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X130 gm_c_stage_2/vcmcn VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X131 gm_c_stage_2/vtail_diff vfiltp vintm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X132 VSS VSS vintm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X133 gm_c_stage_1/vtail_diff vintp vintp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X134 gm_c_stage_1/vcmcn1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X135 vintm VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X136 vintm vim gm_c_stage_0/vtail_diff VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X137 vintm vfiltp gm_c_stage_2/vtail_diff VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X138 VDD VDD vfiltm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X139 ibiasn4 ibiasn4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X140 gm_c_stage_1/vcmcn1 vocm gm_c_stage_1/vcmn_tail1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X141 ibiasn1 ibiasn1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X142 gm_c_stage_1/vcmcn1 vocm gm_c_stage_1/vcmn_tail1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X143 VSS VSS gm_c_stage_3/vtail_diff VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X144 VSS VSS gm_c_stage_0/vcmcn2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X145 gm_c_stage_2/vtail_diff vfiltm vintp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X146 VSS ibiasn2 ibiasn2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X147 VDD VDD vintp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X148 vfiltm vintm gm_c_stage_3/vtail_diff VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X149 gm_c_stage_3/vcmn_tail1 VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X150 gm_c_stage_0/vcmn_tail1 vocm gm_c_stage_0/vcmcn1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X151 gm_c_stage_2/vcmn_tail1 vintp gm_c_stage_2/vcmcn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X152 VSS gm_c_stage_1/vcmc gm_c_stage_1/vcmc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X153 VDD gm_c_stage_3/vcmcn1 gm_c_stage_3/vcmcn1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X154 ibiasn3 ibiasn3 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X155 gm_c_stage_0/vcmcn1 vocm gm_c_stage_0/vcmn_tail1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X156 gm_c_stage_2/vcmcn vintp gm_c_stage_2/vcmn_tail1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X157 gm_c_stage_1/vcmn_tail1 vintp gm_c_stage_1/vcmcn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X158 VSS ibiasn4 ibiasn4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X159 VSS ibiasn1 ibiasn1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X160 gm_c_stage_2/vcmn_tail2 vocm gm_c_stage_2/vcmcn2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X161 gm_c_stage_3/vcmn_tail1 vocm gm_c_stage_3/vcmcn1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.16e+12p ps=9.16e+06u w=2e+06u l=1e+06u
X162 VSS VSS gm_c_stage_0/vcmcn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X163 gm_c_stage_3/vtail_diff vintp vfiltp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X164 VSS gm_c_stage_0/vcmc gm_c_stage_0/vtail_diff VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X165 VSS ibiasn2 ibiasn2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X166 gm_c_stage_3/vcmcn1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X167 ibiasn3 ibiasn3 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X168 gm_c_stage_2/vcmcn2 VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X169 gm_c_stage_1/vtail_diff VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X170 gm_c_stage_0/vcmcn VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X171 VSS ibiasn4 ibiasn4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X172 VSS VSS gm_c_stage_1/vcmcn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X173 vintp gm_c_stage_2/vbiasp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X174 ibiasn2 ibiasn2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X175 gm_c_stage_3/vcmcn1 vocm gm_c_stage_3/vcmn_tail1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X176 gm_c_stage_1/vcmcn2 vocm gm_c_stage_1/vcmn_tail2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X177 gm_c_stage_2/vcmcn2 gm_c_stage_2/vcmcn2 VDD VDD sky130_fd_pr__pfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
X178 gm_c_stage_0/vcmn_tail1 VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X179 gm_c_stage_1/vcmcn2 gm_c_stage_1/vcmcn2 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X180 gm_c_stage_3/vcmcn1 vocm gm_c_stage_3/vcmn_tail1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X181 gm_c_stage_1/vcmcn2 vocm gm_c_stage_1/vcmn_tail2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X182 gm_c_stage_3/vtail_diff VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X183 VSS VSS vintm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X184 VDD VDD vfiltp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X185 gm_c_stage_3/vcmcn vfiltm gm_c_stage_3/vcmn_tail2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X186 VDD gm_c_stage_2/vcmcn1 gm_c_stage_2/vcmcn1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X187 gm_c_stage_1/vcmcn vintp gm_c_stage_1/vcmn_tail1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X188 ibiasn4 ibiasn4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X189 gm_c_stage_1/vtail_diff ibiasn2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X190 VSS gm_c_stage_3/vcmc gm_c_stage_3/vcmc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X191 VSS VSS gm_c_stage_1/vcmcn2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X192 vintm gm_c_stage_2/vbiasp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X193 gm_c_stage_0/vcmn_tail2 vintp gm_c_stage_0/vcmcn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X194 gm_c_stage_1/vcmn_tail2 vintm gm_c_stage_1/vcmcn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X195 VSS VSS gm_c_stage_1/vbiasp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X196 gm_c_stage_3/vcmn_tail1 vfiltp gm_c_stage_3/vcmcn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X197 VDD VDD gm_c_stage_2/vcmcn2 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X198 gm_c_stage_0/vcmcn vintp gm_c_stage_0/vcmn_tail2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X199 VSS VSS gm_c_stage_0/vtail_diff VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X200 gm_c_stage_2/vtail_diff VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X201 vintm vintm gm_c_stage_1/vtail_diff VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X202 gm_c_stage_1/vbiasp VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
X203 vintp vfiltm gm_c_stage_2/vtail_diff VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X204 ibiasn2 VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X205 VSS ibiasn3 ibiasn3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X206 gm_c_stage_0/vcmc VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
X207 gm_c_stage_0/vcmn_tail2 vocm gm_c_stage_0/vcmcn2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X208 gm_c_stage_3/vbiasp ibiasn3 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X209 ibiasn4 ibiasn4 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X210 ibiasn2 ibiasn2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X211 VSS VSS gm_c_stage_3/vcmcn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X212 VDD VDD vintm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X213 ibiasn3 ibiasn3 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X214 VSS VSS gm_c_stage_0/vcmn_tail2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X215 VSS ibiasn2 ibiasn2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X216 VSS VSS vfiltm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X217 gm_c_stage_2/vcmn_tail1 vocm gm_c_stage_2/vcmcn1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X218 gm_c_stage_0/vcmcn2 gm_c_stage_0/vcmcn2 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X219 gm_c_stage_2/vcmn_tail2 vintm gm_c_stage_2/vcmcn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X220 gm_c_stage_3/vcmcn vfiltp gm_c_stage_3/vcmn_tail1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X221 gm_c_stage_0/vtail_diff vip vintp VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X222 gm_c_stage_2/vcmcn1 vocm gm_c_stage_2/vcmn_tail1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X223 gm_c_stage_2/vcmcn vintm gm_c_stage_2/vcmn_tail2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X224 vintp vip gm_c_stage_0/vtail_diff VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X225 VDD gm_c_stage_1/vcmcn gm_c_stage_1/vcmc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X226 VSS ibiasn3 ibiasn3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X227 ibiasn1 VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X228 VSS VSS gm_c_stage_2/vcmcn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X229 VSS gm_c_stage_2/vcmc gm_c_stage_2/vtail_diff VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X230 vfiltm vintm gm_c_stage_3/vtail_diff VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X231 gm_c_stage_3/vbiasp VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X232 gm_c_stage_0/vcmcn1 vocm gm_c_stage_0/vcmn_tail1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X233 gm_c_stage_1/vcmn_tail1 vocm gm_c_stage_1/vcmcn1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X234 ibiasn3 VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X235 gm_c_stage_1/vcmn_tail2 vocm gm_c_stage_1/vcmcn2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X236 gm_c_stage_0/vtail_diff vim vintm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X237 VSS VSS ibiasn4 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X238 ibiasn3 ibiasn3 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X239 VSS gm_c_stage_1/vcmc gm_c_stage_1/vtail_diff VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X240 gm_c_stage_1/vcmc VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X241 gm_c_stage_3/vcmcn2 gm_c_stage_3/vcmcn2 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X242 vintm gm_c_stage_1/vbiasp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X243 VSS VSS gm_c_stage_3/vcmn_tail2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X244 gm_c_stage_0/vtail_diff VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X245 ibiasn1 ibiasn1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X246 gm_c_stage_3/vcmn_tail2 vfiltm gm_c_stage_3/vcmcn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X247 gm_c_stage_0/vcmcn vintm gm_c_stage_0/vcmn_tail1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X248 gm_c_stage_2/vcmcn gm_c_stage_2/vcmcn VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X249 gm_c_stage_3/vtail_diff ibiasn3 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X250 VDD gm_c_stage_1/vbiasp gm_c_stage_1/vbiasp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X251 gm_c_stage_0/vcmcn2 vocm gm_c_stage_0/vcmn_tail2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X252 VSS VSS gm_c_stage_2/vtail_diff VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X253 gm_c_stage_1/vcmn_tail2 ibiasn2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X254 VSS gm_c_stage_2/vcmc gm_c_stage_2/vcmc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X255 ibiasn2 ibiasn2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X256 VDD gm_c_stage_3/vcmcn gm_c_stage_3/vcmc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X257 gm_c_stage_3/vcmcn vfiltm gm_c_stage_3/vcmn_tail2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X258 gm_c_stage_0/vbiasp VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X259 gm_c_stage_2/vcmc VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X260 gm_c_stage_3/vcmn_tail1 vocm gm_c_stage_3/vcmcn1 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X261 VDD gm_c_stage_0/vcmcn gm_c_stage_0/vcmc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X262 VDD VDD vintp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X263 gm_c_stage_3/vcmc VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X264 VSS gm_c_stage_3/vcmc gm_c_stage_3/vtail_diff VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X265 vintp vfiltm gm_c_stage_2/vtail_diff VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X266 vfiltm gm_c_stage_3/vbiasp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X267 VSS ibiasn3 ibiasn3 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X268 gm_c_stage_1/vcmn_tail1 vintp gm_c_stage_1/vcmcn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X269 gm_c_stage_2/vcmn_tail2 vocm gm_c_stage_2/vcmcn2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X270 gm_c_stage_2/vtail_diff vfiltp vintm VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X271 gm_c_stage_1/vcmcn2 VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
C0 gm_c_stage_1/vcmn_tail2 vintm 0.32fF
C1 gm_c_stage_0/vcmcn2 gm_c_stage_0/vbiasp 0.88fF
C2 gm_c_stage_0/vcmn_tail1 gm_c_stage_0/vtail_diff 0.49fF
C3 gm_c_stage_2/vtail_diff gm_c_stage_2/vcmc 0.03fF
C4 vintp gm_c_stage_2/vbiasp 0.32fF
C5 vocm gm_c_stage_2/vcmc 0.24fF
C6 gm_c_stage_1/vcmcn gm_c_stage_1/vcmn_tail2 0.58fF
C7 VDD gm_c_stage_0/vbiasp 3.04fF
C8 gm_c_stage_3/vcmcn gm_c_stage_3/vcmc 0.05fF
C9 gm_c_stage_3/vcmn_tail1 gm_c_stage_3/vcmc 0.15fF
C10 gm_c_stage_1/vcmcn1 gm_c_stage_1/vcmcn2 0.17fF
C11 gm_c_stage_1/vcmc vintm 0.10fF
C12 vintm vim 1.21fF
C13 gm_c_stage_0/vcmcn2 vintp 2.15fF
C14 vfiltp vintm 0.71fF
C15 vfiltm vintp 3.06fF
C16 vocm gm_c_stage_1/vtail_diff 1.19fF
C17 gm_c_stage_1/vcmcn gm_c_stage_1/vcmc 0.05fF
C18 vintm gm_c_stage_0/vtail_diff 2.75fF
C19 vfiltp gm_c_stage_3/vcmn_tail2 0.07fF
C20 gm_c_stage_2/vcmcn2 gm_c_stage_2/vcmcn1 0.17fF
C21 vintp VDD 2.28fF
C22 gm_c_stage_3/vcmcn1 VDD 3.44fF
C23 vintp gm_c_stage_2/vcmc 0.10fF
C24 vintm gm_c_stage_1/vcmn_tail1 0.07fF
C25 gm_c_stage_1/vcmcn1 gm_c_stage_1/vcmcn 1.18fF
C26 gm_c_stage_3/vtail_diff vocm 1.19fF
C27 gm_c_stage_0/vcmn_tail1 gm_c_stage_0/vcmc 0.15fF
C28 gm_c_stage_1/vcmcn gm_c_stage_1/vcmn_tail1 0.58fF
C29 vintp gm_c_stage_1/vtail_diff 3.07fF
C30 gm_c_stage_0/vcmcn2 gm_c_stage_0/vcmcn 1.28fF
C31 gm_c_stage_2/vcmcn1 vocm 1.07fF
C32 gm_c_stage_0/vcmc vintm 0.10fF
C33 gm_c_stage_0/vcmcn VDD 4.05fF
C34 gm_c_stage_2/vbiasp gm_c_stage_2/vcmn_tail2 0.90fF
C35 gm_c_stage_3/vtail_diff vintp 0.33fF
C36 gm_c_stage_3/vcmcn gm_c_stage_3/vbiasp 0.53fF
C37 ibiasn2 gm_c_stage_1/vbiasp 0.04fF
C38 vintp gm_c_stage_2/vcmcn1 0.13fF
C39 gm_c_stage_1/vcmn_tail2 ibiasn2 0.06fF
C40 vfiltm gm_c_stage_2/vbiasp 0.10fF
C41 ibiasn1 gm_c_stage_0/vbiasp 0.04fF
C42 gm_c_stage_0/vcmn_tail1 vintm 2.84fF
C43 gm_c_stage_0/vcmcn1 vocm 1.07fF
C44 vfiltp gm_c_stage_3/vbiasp 0.38fF
C45 gm_c_stage_1/vcmcn2 vintm 2.12fF
C46 gm_c_stage_2/vbiasp VDD 3.04fF
C47 gm_c_stage_1/vcmc ibiasn2 0.11fF
C48 gm_c_stage_0/vcmcn1 gm_c_stage_0/vbiasp 0.19fF
C49 gm_c_stage_1/vcmcn2 gm_c_stage_1/vcmcn 1.28fF
C50 vip vim 0.51fF
C51 gm_c_stage_0/vcmcn2 VDD 1.51fF
C52 gm_c_stage_3/vcmn_tail2 gm_c_stage_3/vcmcn2 0.58fF
C53 vfiltm VDD 0.59fF
C54 gm_c_stage_3/vcmcn vocm 2.07fF
C55 vip gm_c_stage_0/vtail_diff 2.65fF
C56 vocm gm_c_stage_1/vbiasp 0.10fF
C57 gm_c_stage_3/vcmn_tail1 vocm 2.22fF
C58 gm_c_stage_1/vcmcn vintm 1.20fF
C59 gm_c_stage_0/vcmcn1 vintp 0.91fF
C60 gm_c_stage_1/vcmn_tail1 ibiasn2 0.07fF
C61 gm_c_stage_1/vcmn_tail2 vocm 4.74fF
C62 gm_c_stage_2/vcmc VDD 2.70fF
C63 gm_c_stage_2/vcmcn vintm 2.62fF
C64 gm_c_stage_3/vcmc vintm 0.10fF
C65 gm_c_stage_3/vcmcn vintp 0.11fF
C66 vintp gm_c_stage_1/vbiasp 0.42fF
C67 vfiltp gm_c_stage_2/vtail_diff 2.64fF
C68 gm_c_stage_0/vcmn_tail2 vocm 4.74fF
C69 vfiltp vocm 2.82fF
C70 gm_c_stage_3/vcmcn1 gm_c_stage_3/vcmcn 1.18fF
C71 gm_c_stage_3/vcmn_tail1 gm_c_stage_3/vcmcn1 0.58fF
C72 vocm gm_c_stage_0/vtail_diff 1.19fF
C73 gm_c_stage_0/vcmn_tail2 gm_c_stage_0/vbiasp 0.90fF
C74 vfiltm gm_c_stage_3/vtail_diff 0.58fF
C75 gm_c_stage_1/vcmcn1 vocm 1.07fF
C76 gm_c_stage_2/vcmcn1 gm_c_stage_2/vbiasp 0.19fF
C77 gm_c_stage_0/vcmcn1 gm_c_stage_0/vcmcn 1.18fF
C78 gm_c_stage_1/vcmn_tail1 vocm 0.32fF
C79 gm_c_stage_1/vcmc vintp 0.10fF
C80 vintp vim 1.61fF
C81 gm_c_stage_0/vcmn_tail2 vintp 0.32fF
C82 gm_c_stage_2/vcmn_tail1 gm_c_stage_2/vcmcn 0.58fF
C83 vfiltp vintp 1.72fF
C84 vfiltp gm_c_stage_3/vcmcn1 0.03fF
C85 vintp gm_c_stage_0/vtail_diff 0.58fF
C86 gm_c_stage_2/vcmcn1 VDD 3.44fF
C87 gm_c_stage_1/vcmcn1 vintp 0.15fF
C88 ibiasn3 gm_c_stage_3/vtail_diff 0.06fF
C89 gm_c_stage_2/vcmcn1 gm_c_stage_2/vcmc 2.37fF
C90 vintp gm_c_stage_1/vcmn_tail1 2.83fF
C91 gm_c_stage_3/vbiasp gm_c_stage_3/vcmcn2 0.88fF
C92 gm_c_stage_2/vcmn_tail1 ibiasn4 0.07fF
C93 gm_c_stage_3/vbiasp gm_c_stage_3/vcmn_tail2 0.90fF
C94 gm_c_stage_0/vcmcn gm_c_stage_0/vcmn_tail2 0.58fF
C95 vip vintm 0.30fF
C96 gm_c_stage_0/vcmcn1 gm_c_stage_0/vcmcn2 0.17fF
C97 gm_c_stage_2/vcmcn2 vintm 2.05fF
C98 vintp gm_c_stage_0/vcmc 0.10fF
C99 gm_c_stage_0/vcmcn1 VDD 3.44fF
C100 gm_c_stage_0/vcmn_tail1 vocm 0.32fF
C101 gm_c_stage_1/vcmcn2 vocm 0.28fF
C102 vfiltp gm_c_stage_2/vcmn_tail2 0.07fF
C103 vfiltm gm_c_stage_3/vcmcn 1.20fF
C104 gm_c_stage_2/vcmcn2 gm_c_stage_2/vcmcn 1.28fF
C105 vocm gm_c_stage_3/vcmcn2 0.28fF
C106 gm_c_stage_3/vcmcn VDD 4.05fF
C107 gm_c_stage_1/vbiasp VDD 3.04fF
C108 vintm gm_c_stage_2/vtail_diff 0.58fF
C109 vintm vocm 6.20fF
C110 vfiltp gm_c_stage_2/vbiasp 0.10fF
C111 gm_c_stage_3/vcmn_tail2 vocm 2.82fF
C112 gm_c_stage_0/vcmcn gm_c_stage_0/vcmc 0.05fF
C113 gm_c_stage_1/vcmcn vocm 2.07fF
C114 vintm gm_c_stage_0/vbiasp 0.51fF
C115 gm_c_stage_1/vcmcn2 vintp 0.10fF
C116 gm_c_stage_0/vcmcn2 gm_c_stage_0/vcmn_tail2 0.58fF
C117 ibiasn3 gm_c_stage_3/vcmn_tail1 0.07fF
C118 vfiltp vfiltm 3.22fF
C119 gm_c_stage_2/vcmcn vocm 2.07fF
C120 gm_c_stage_3/vcmc vocm 0.24fF
C121 gm_c_stage_1/vcmc VDD 2.70fF
C122 gm_c_stage_3/vcmcn1 gm_c_stage_3/vcmcn2 0.17fF
C123 vfiltp VDD 0.82fF
C124 vintp vintm 13.75fF
C125 gm_c_stage_3/vcmcn1 vintm 0.12fF
C126 gm_c_stage_2/vcmn_tail1 gm_c_stage_2/vtail_diff 0.49fF
C127 gm_c_stage_1/vcmcn vintp 1.45fF
C128 gm_c_stage_2/vcmn_tail1 vocm 2.22fF
C129 gm_c_stage_1/vcmcn1 VDD 3.44fF
C130 gm_c_stage_3/vcmn_tail1 gm_c_stage_3/vtail_diff 0.49fF
C131 ibiasn4 gm_c_stage_2/vtail_diff 0.06fF
C132 gm_c_stage_1/vcmc gm_c_stage_1/vtail_diff 0.03fF
C133 gm_c_stage_0/vcmn_tail1 gm_c_stage_0/vcmcn 0.58fF
C134 vintp gm_c_stage_2/vcmcn 1.12fF
C135 gm_c_stage_3/vcmc vintp 0.51fF
C136 gm_c_stage_3/vcmcn1 gm_c_stage_3/vcmc 2.37fF
C137 gm_c_stage_0/vcmcn vintm 0.42fF
C138 gm_c_stage_2/vcmn_tail1 vintp 2.83fF
C139 gm_c_stage_1/vcmn_tail1 gm_c_stage_1/vtail_diff 0.49fF
C140 vfiltp gm_c_stage_3/vtail_diff 2.76fF
C141 gm_c_stage_0/vcmc VDD 2.70fF
C142 vintm gm_c_stage_2/vcmn_tail2 0.32fF
C143 gm_c_stage_2/vcmcn2 vocm 0.28fF
C144 gm_c_stage_2/vbiasp vintm 0.34fF
C145 gm_c_stage_2/vcmcn gm_c_stage_2/vcmn_tail2 0.58fF
C146 gm_c_stage_0/vcmn_tail2 ibiasn1 0.06fF
C147 vfiltm gm_c_stage_3/vcmcn2 2.12fF
C148 gm_c_stage_1/vcmcn2 VDD 1.51fF
C149 gm_c_stage_3/vcmcn1 gm_c_stage_3/vbiasp 0.19fF
C150 gm_c_stage_3/vcmn_tail1 gm_c_stage_3/vcmcn 0.58fF
C151 vfiltm vintm 3.38fF
C152 ibiasn1 gm_c_stage_0/vtail_diff 0.06fF
C153 gm_c_stage_3/vcmcn2 VDD 1.51fF
C154 vfiltm gm_c_stage_3/vcmn_tail2 0.32fF
C155 vip vintp 0.28fF
C156 gm_c_stage_2/vcmcn gm_c_stage_2/vbiasp 0.53fF
C157 vintm VDD 2.01fF
C158 gm_c_stage_1/vcmn_tail2 gm_c_stage_1/vbiasp 0.90fF
C159 vocm gm_c_stage_2/vtail_diff 1.19fF
C160 ibiasn4 gm_c_stage_2/vcmn_tail2 0.06fF
C161 vintm gm_c_stage_2/vcmc 0.54fF
C162 gm_c_stage_1/vcmcn VDD 4.05fF
C163 vfiltm gm_c_stage_2/vcmcn 0.12fF
C164 vocm gm_c_stage_0/vbiasp 0.10fF
C165 vfiltp gm_c_stage_3/vcmcn 0.42fF
C166 vintm gm_c_stage_1/vtail_diff 4.99fF
C167 vfiltp gm_c_stage_3/vcmn_tail1 2.83fF
C168 ibiasn4 gm_c_stage_2/vbiasp 0.04fF
C169 gm_c_stage_2/vcmcn VDD 4.05fF
C170 gm_c_stage_3/vcmc VDD 2.70fF
C171 ibiasn3 gm_c_stage_3/vcmn_tail2 0.06fF
C172 gm_c_stage_2/vcmcn gm_c_stage_2/vcmc 0.05fF
C173 gm_c_stage_1/vcmcn1 gm_c_stage_1/vbiasp 0.19fF
C174 ibiasn1 gm_c_stage_0/vcmc 0.11fF
C175 vintp gm_c_stage_2/vtail_diff 2.75fF
C176 vintp vocm 3.46fF
C177 gm_c_stage_3/vcmcn1 vocm 1.07fF
C178 gm_c_stage_3/vtail_diff vintm 2.72fF
C179 gm_c_stage_0/vcmcn1 gm_c_stage_0/vcmc 2.37fF
C180 vintp gm_c_stage_0/vbiasp 0.44fF
C181 gm_c_stage_2/vcmn_tail1 gm_c_stage_2/vcmc 0.15fF
C182 ibiasn3 gm_c_stage_3/vcmc 0.11fF
C183 ibiasn4 gm_c_stage_2/vcmc 0.11fF
C184 vim gm_c_stage_0/vtail_diff 0.33fF
C185 gm_c_stage_1/vcmcn1 gm_c_stage_1/vcmc 2.37fF
C186 gm_c_stage_2/vcmcn1 vintm 0.12fF
C187 gm_c_stage_2/vcmcn2 gm_c_stage_2/vcmn_tail2 0.58fF
C188 gm_c_stage_1/vcmc gm_c_stage_1/vcmn_tail1 0.15fF
C189 gm_c_stage_3/vcmcn1 vintp 0.78fF
C190 gm_c_stage_3/vtail_diff gm_c_stage_3/vcmc 0.03fF
C191 gm_c_stage_0/vcmn_tail1 ibiasn1 0.07fF
C192 gm_c_stage_0/vcmcn vocm 2.07fF
C193 vfiltm gm_c_stage_3/vbiasp 0.44fF
C194 gm_c_stage_1/vcmcn1 gm_c_stage_1/vcmn_tail1 0.58fF
C195 gm_c_stage_2/vcmcn2 gm_c_stage_2/vbiasp 0.88fF
C196 gm_c_stage_2/vcmcn1 gm_c_stage_2/vcmcn 1.18fF
C197 gm_c_stage_0/vcmcn gm_c_stage_0/vbiasp 0.53fF
C198 gm_c_stage_0/vcmcn1 gm_c_stage_0/vcmn_tail1 0.58fF
C199 gm_c_stage_3/vbiasp VDD 3.04fF
C200 vfiltm gm_c_stage_2/vcmcn2 0.19fF
C201 gm_c_stage_2/vcmn_tail1 gm_c_stage_2/vcmcn1 0.58fF
C202 vocm gm_c_stage_2/vcmn_tail2 2.82fF
C203 gm_c_stage_0/vcmcn vintp 1.30fF
C204 gm_c_stage_0/vcmc gm_c_stage_0/vtail_diff 0.03fF
C205 gm_c_stage_0/vcmcn1 vintm 0.03fF
C206 gm_c_stage_2/vcmcn2 VDD 1.51fF
C207 ibiasn3 gm_c_stage_3/vbiasp 0.04fF
C208 gm_c_stage_1/vcmcn2 gm_c_stage_1/vbiasp 0.88fF
C209 gm_c_stage_3/vcmcn gm_c_stage_3/vcmcn2 1.28fF
C210 ibiasn2 gm_c_stage_1/vtail_diff 0.06fF
C211 gm_c_stage_1/vcmcn2 gm_c_stage_1/vcmn_tail2 0.58fF
C212 gm_c_stage_3/vcmcn vintm 0.19fF
C213 vintm gm_c_stage_1/vbiasp 0.61fF
C214 gm_c_stage_0/vcmcn2 vocm 0.28fF
C215 vfiltm gm_c_stage_2/vtail_diff 0.33fF
C216 vfiltm vocm 0.51fF
C217 gm_c_stage_3/vcmcn gm_c_stage_3/vcmn_tail2 0.58fF
C218 gm_c_stage_1/vcmcn gm_c_stage_1/vbiasp 0.53fF
C219 gm_c_stage_3/vcmcn2 VSS 3.23fF
C220 gm_c_stage_3/vcmcn1 VSS 3.18fF
C221 gm_c_stage_3/vcmcn VSS 10.01fF
C222 gm_c_stage_3/vbiasp VSS 5.02fF
C223 gm_c_stage_3/vtail_diff VSS 3.39fF
C224 gm_c_stage_3/vcmn_tail2 VSS 5.21fF
C225 gm_c_stage_3/vcmn_tail1 VSS 10.52fF
C226 ibiasn3 VSS 18.85fF
C227 gm_c_stage_3/vcmc VSS 6.85fF
C228 gm_c_stage_1/vcmcn2 VSS 3.23fF
C229 gm_c_stage_1/vcmcn1 VSS 3.18fF
C230 gm_c_stage_1/vcmcn VSS 10.01fF
C231 gm_c_stage_1/vbiasp VSS 5.02fF
C232 gm_c_stage_1/vtail_diff VSS 3.39fF
C233 gm_c_stage_1/vcmn_tail2 VSS 5.21fF
C234 gm_c_stage_1/vcmn_tail1 VSS 10.52fF
C235 ibiasn2 VSS 0.14fF
C236 gm_c_stage_1/vcmc VSS 6.85fF
C237 ibiasn4 VSS 18.85fF
C238 gm_c_stage_2/vcmn_tail2 VSS 5.21fF
C239 gm_c_stage_2/vtail_diff VSS 3.39fF
C240 gm_c_stage_2/vcmn_tail1 VSS 10.52fF
C241 vfiltm VSS 14.59fF
C242 vfiltp VSS 15.62fF
C243 ibiasn1 VSS 18.85fF
C244 gm_c_stage_0/vcmn_tail2 VSS 5.21fF
C245 gm_c_stage_0/vtail_diff VSS 3.39fF
C246 gm_c_stage_0/vcmn_tail1 VSS 10.52fF
C247 vim VSS 2.03fF
C248 vip VSS 2.50fF
C249 vocm VSS 38.83fF
C250 gm_c_stage_2/vcmc VSS 6.85fF
C251 gm_c_stage_2/vcmcn2 VSS 3.23fF
C252 gm_c_stage_2/vcmcn1 VSS 3.18fF
C253 gm_c_stage_2/vcmcn VSS 10.01fF
C254 gm_c_stage_2/vbiasp VSS 5.02fF
C255 gm_c_stage_0/vcmc VSS 6.85fF
C256 vintm VSS 37.79fF
C257 vintp VSS 37.02fF
C258 gm_c_stage_0/vcmcn2 VSS 3.23fF
C259 gm_c_stage_0/vcmcn1 VSS 3.18fF
C260 gm_c_stage_0/vcmcn VSS 10.01fF
C261 gm_c_stage_0/vbiasp VSS 5.02fF
C262 VDD VSS 436.63fF
.ends

