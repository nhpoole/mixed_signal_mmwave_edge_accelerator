* NGSPICE file created from metal_resistor_test_flat.ext - technology: sky130A

.subckt sky130_fd_pr__res_generic_m1_6PYWN2 VSUBS
R0 m1_n100_n87# m1_n100_30# sky130_fd_pr__res_generic_m1 w=1e+06u l=300000u
.ends


* Top level circuit metal_resistor_test_flat

Xsky130_fd_pr__res_generic_m1_6PYWN2_0 VSUBS sky130_fd_pr__res_generic_m1_6PYWN2
.end

