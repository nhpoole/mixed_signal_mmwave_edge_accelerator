magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect -1610 -2160 1504 2160
<< metal3 >>
rect -350 -900 244 900
<< mimcap >>
rect -250 752 150 800
rect -250 -752 -202 752
rect 102 -752 150 752
rect -250 -800 150 -752
<< mimcapcontact >>
rect -202 -752 102 752
<< metal4 >>
rect -211 752 111 761
rect -211 -752 -202 752
rect 102 -752 111 752
rect -211 -761 111 -752
<< properties >>
string FIXED_BBOX -350 -900 250 900
<< end >>
