magic
tech sky130A
timestamp 1624494425
<< error_p >>
rect 0 25 29 28
rect 0 8 6 25
rect 0 5 29 8
<< locali >>
rect 6 25 23 33
rect 6 0 23 8
<< viali >>
rect 6 8 23 25
<< metal1 >>
rect 0 25 29 28
rect 0 8 6 25
rect 23 8 29 25
rect 0 5 29 8
<< properties >>
string FIXED_BBOX 0 0 29 33
<< end >>
