magic
tech sky130A
magscale 1 2
timestamp 1626065694
<< checkpaint >>
rect -1302 -1260 1910 53400
<< metal1 >>
rect 78 0 114 52140
rect 150 0 186 52140
rect 222 51429 258 51770
rect 222 50639 258 51271
rect 222 49849 258 50481
rect 222 49059 258 49691
rect 222 48269 258 48901
rect 222 47479 258 48111
rect 222 46689 258 47321
rect 222 45899 258 46531
rect 222 45109 258 45741
rect 222 44319 258 44951
rect 222 43529 258 44161
rect 222 42739 258 43371
rect 222 41949 258 42581
rect 222 41159 258 41791
rect 222 40369 258 41001
rect 222 39579 258 40211
rect 222 38789 258 39421
rect 222 37999 258 38631
rect 222 37209 258 37841
rect 222 36419 258 37051
rect 222 35629 258 36261
rect 222 34839 258 35471
rect 222 34049 258 34681
rect 222 33259 258 33891
rect 222 32469 258 33101
rect 222 31679 258 32311
rect 222 30889 258 31521
rect 222 30099 258 30731
rect 222 29309 258 29941
rect 222 28519 258 29151
rect 222 27729 258 28361
rect 222 26939 258 27571
rect 222 26149 258 26781
rect 222 25359 258 25991
rect 222 24569 258 25201
rect 222 23779 258 24411
rect 222 22989 258 23621
rect 222 22199 258 22831
rect 222 21409 258 22041
rect 222 20619 258 21251
rect 222 19829 258 20461
rect 222 19039 258 19671
rect 222 18249 258 18881
rect 222 17459 258 18091
rect 222 16669 258 17301
rect 222 15879 258 16511
rect 222 15089 258 15721
rect 222 14299 258 14931
rect 222 13509 258 14141
rect 222 12719 258 13351
rect 222 11929 258 12561
rect 222 11139 258 11771
rect 222 10349 258 10981
rect 222 9559 258 10191
rect 222 8769 258 9401
rect 222 7979 258 8611
rect 222 7189 258 7821
rect 222 6399 258 7031
rect 222 5609 258 6241
rect 222 4819 258 5451
rect 222 4029 258 4661
rect 222 3239 258 3871
rect 222 2449 258 3081
rect 222 1659 258 2291
rect 222 869 258 1501
rect 222 370 258 711
rect 294 0 330 52140
rect 366 0 402 52140
<< metal2 >>
rect 0 51673 624 51721
rect 186 51549 294 51625
rect 0 51453 624 51501
rect 186 51295 294 51405
rect 0 51199 624 51247
rect 186 51075 294 51151
rect 0 50979 624 51027
rect 0 50883 624 50931
rect 186 50759 294 50835
rect 0 50663 624 50711
rect 186 50505 294 50615
rect 0 50409 624 50457
rect 186 50285 294 50361
rect 0 50189 624 50237
rect 0 50093 624 50141
rect 186 49969 294 50045
rect 0 49873 624 49921
rect 186 49715 294 49825
rect 0 49619 624 49667
rect 186 49495 294 49571
rect 0 49399 624 49447
rect 0 49303 624 49351
rect 186 49179 294 49255
rect 0 49083 624 49131
rect 186 48925 294 49035
rect 0 48829 624 48877
rect 186 48705 294 48781
rect 0 48609 624 48657
rect 0 48513 624 48561
rect 186 48389 294 48465
rect 0 48293 624 48341
rect 186 48135 294 48245
rect 0 48039 624 48087
rect 186 47915 294 47991
rect 0 47819 624 47867
rect 0 47723 624 47771
rect 186 47599 294 47675
rect 0 47503 624 47551
rect 186 47345 294 47455
rect 0 47249 624 47297
rect 186 47125 294 47201
rect 0 47029 624 47077
rect 0 46933 624 46981
rect 186 46809 294 46885
rect 0 46713 624 46761
rect 186 46555 294 46665
rect 0 46459 624 46507
rect 186 46335 294 46411
rect 0 46239 624 46287
rect 0 46143 624 46191
rect 186 46019 294 46095
rect 0 45923 624 45971
rect 186 45765 294 45875
rect 0 45669 624 45717
rect 186 45545 294 45621
rect 0 45449 624 45497
rect 0 45353 624 45401
rect 186 45229 294 45305
rect 0 45133 624 45181
rect 186 44975 294 45085
rect 0 44879 624 44927
rect 186 44755 294 44831
rect 0 44659 624 44707
rect 0 44563 624 44611
rect 186 44439 294 44515
rect 0 44343 624 44391
rect 186 44185 294 44295
rect 0 44089 624 44137
rect 186 43965 294 44041
rect 0 43869 624 43917
rect 0 43773 624 43821
rect 186 43649 294 43725
rect 0 43553 624 43601
rect 186 43395 294 43505
rect 0 43299 624 43347
rect 186 43175 294 43251
rect 0 43079 624 43127
rect 0 42983 624 43031
rect 186 42859 294 42935
rect 0 42763 624 42811
rect 186 42605 294 42715
rect 0 42509 624 42557
rect 186 42385 294 42461
rect 0 42289 624 42337
rect 0 42193 624 42241
rect 186 42069 294 42145
rect 0 41973 624 42021
rect 186 41815 294 41925
rect 0 41719 624 41767
rect 186 41595 294 41671
rect 0 41499 624 41547
rect 0 41403 624 41451
rect 186 41279 294 41355
rect 0 41183 624 41231
rect 186 41025 294 41135
rect 0 40929 624 40977
rect 186 40805 294 40881
rect 0 40709 624 40757
rect 0 40613 624 40661
rect 186 40489 294 40565
rect 0 40393 624 40441
rect 186 40235 294 40345
rect 0 40139 624 40187
rect 186 40015 294 40091
rect 0 39919 624 39967
rect 0 39823 624 39871
rect 186 39699 294 39775
rect 0 39603 624 39651
rect 186 39445 294 39555
rect 0 39349 624 39397
rect 186 39225 294 39301
rect 0 39129 624 39177
rect 0 39033 624 39081
rect 186 38909 294 38985
rect 0 38813 624 38861
rect 186 38655 294 38765
rect 0 38559 624 38607
rect 186 38435 294 38511
rect 0 38339 624 38387
rect 0 38243 624 38291
rect 186 38119 294 38195
rect 0 38023 624 38071
rect 186 37865 294 37975
rect 0 37769 624 37817
rect 186 37645 294 37721
rect 0 37549 624 37597
rect 0 37453 624 37501
rect 186 37329 294 37405
rect 0 37233 624 37281
rect 186 37075 294 37185
rect 0 36979 624 37027
rect 186 36855 294 36931
rect 0 36759 624 36807
rect 0 36663 624 36711
rect 186 36539 294 36615
rect 0 36443 624 36491
rect 186 36285 294 36395
rect 0 36189 624 36237
rect 186 36065 294 36141
rect 0 35969 624 36017
rect 0 35873 624 35921
rect 186 35749 294 35825
rect 0 35653 624 35701
rect 186 35495 294 35605
rect 0 35399 624 35447
rect 186 35275 294 35351
rect 0 35179 624 35227
rect 0 35083 624 35131
rect 186 34959 294 35035
rect 0 34863 624 34911
rect 186 34705 294 34815
rect 0 34609 624 34657
rect 186 34485 294 34561
rect 0 34389 624 34437
rect 0 34293 624 34341
rect 186 34169 294 34245
rect 0 34073 624 34121
rect 186 33915 294 34025
rect 0 33819 624 33867
rect 186 33695 294 33771
rect 0 33599 624 33647
rect 0 33503 624 33551
rect 186 33379 294 33455
rect 0 33283 624 33331
rect 186 33125 294 33235
rect 0 33029 624 33077
rect 186 32905 294 32981
rect 0 32809 624 32857
rect 0 32713 624 32761
rect 186 32589 294 32665
rect 0 32493 624 32541
rect 186 32335 294 32445
rect 0 32239 624 32287
rect 186 32115 294 32191
rect 0 32019 624 32067
rect 0 31923 624 31971
rect 186 31799 294 31875
rect 0 31703 624 31751
rect 186 31545 294 31655
rect 0 31449 624 31497
rect 186 31325 294 31401
rect 0 31229 624 31277
rect 0 31133 624 31181
rect 186 31009 294 31085
rect 0 30913 624 30961
rect 186 30755 294 30865
rect 0 30659 624 30707
rect 186 30535 294 30611
rect 0 30439 624 30487
rect 0 30343 624 30391
rect 186 30219 294 30295
rect 0 30123 624 30171
rect 186 29965 294 30075
rect 0 29869 624 29917
rect 186 29745 294 29821
rect 0 29649 624 29697
rect 0 29553 624 29601
rect 186 29429 294 29505
rect 0 29333 624 29381
rect 186 29175 294 29285
rect 0 29079 624 29127
rect 186 28955 294 29031
rect 0 28859 624 28907
rect 0 28763 624 28811
rect 186 28639 294 28715
rect 0 28543 624 28591
rect 186 28385 294 28495
rect 0 28289 624 28337
rect 186 28165 294 28241
rect 0 28069 624 28117
rect 0 27973 624 28021
rect 186 27849 294 27925
rect 0 27753 624 27801
rect 186 27595 294 27705
rect 0 27499 624 27547
rect 186 27375 294 27451
rect 0 27279 624 27327
rect 0 27183 624 27231
rect 186 27059 294 27135
rect 0 26963 624 27011
rect 186 26805 294 26915
rect 0 26709 624 26757
rect 186 26585 294 26661
rect 0 26489 624 26537
rect 0 26393 624 26441
rect 186 26269 294 26345
rect 0 26173 624 26221
rect 186 26015 294 26125
rect 0 25919 624 25967
rect 186 25795 294 25871
rect 0 25699 624 25747
rect 0 25603 624 25651
rect 186 25479 294 25555
rect 0 25383 624 25431
rect 186 25225 294 25335
rect 0 25129 624 25177
rect 186 25005 294 25081
rect 0 24909 624 24957
rect 0 24813 624 24861
rect 186 24689 294 24765
rect 0 24593 624 24641
rect 186 24435 294 24545
rect 0 24339 624 24387
rect 186 24215 294 24291
rect 0 24119 624 24167
rect 0 24023 624 24071
rect 186 23899 294 23975
rect 0 23803 624 23851
rect 186 23645 294 23755
rect 0 23549 624 23597
rect 186 23425 294 23501
rect 0 23329 624 23377
rect 0 23233 624 23281
rect 186 23109 294 23185
rect 0 23013 624 23061
rect 186 22855 294 22965
rect 0 22759 624 22807
rect 186 22635 294 22711
rect 0 22539 624 22587
rect 0 22443 624 22491
rect 186 22319 294 22395
rect 0 22223 624 22271
rect 186 22065 294 22175
rect 0 21969 624 22017
rect 186 21845 294 21921
rect 0 21749 624 21797
rect 0 21653 624 21701
rect 186 21529 294 21605
rect 0 21433 624 21481
rect 186 21275 294 21385
rect 0 21179 624 21227
rect 186 21055 294 21131
rect 0 20959 624 21007
rect 0 20863 624 20911
rect 186 20739 294 20815
rect 0 20643 624 20691
rect 186 20485 294 20595
rect 0 20389 624 20437
rect 186 20265 294 20341
rect 0 20169 624 20217
rect 0 20073 624 20121
rect 186 19949 294 20025
rect 0 19853 624 19901
rect 186 19695 294 19805
rect 0 19599 624 19647
rect 186 19475 294 19551
rect 0 19379 624 19427
rect 0 19283 624 19331
rect 186 19159 294 19235
rect 0 19063 624 19111
rect 186 18905 294 19015
rect 0 18809 624 18857
rect 186 18685 294 18761
rect 0 18589 624 18637
rect 0 18493 624 18541
rect 186 18369 294 18445
rect 0 18273 624 18321
rect 186 18115 294 18225
rect 0 18019 624 18067
rect 186 17895 294 17971
rect 0 17799 624 17847
rect 0 17703 624 17751
rect 186 17579 294 17655
rect 0 17483 624 17531
rect 186 17325 294 17435
rect 0 17229 624 17277
rect 186 17105 294 17181
rect 0 17009 624 17057
rect 0 16913 624 16961
rect 186 16789 294 16865
rect 0 16693 624 16741
rect 186 16535 294 16645
rect 0 16439 624 16487
rect 186 16315 294 16391
rect 0 16219 624 16267
rect 0 16123 624 16171
rect 186 15999 294 16075
rect 0 15903 624 15951
rect 186 15745 294 15855
rect 0 15649 624 15697
rect 186 15525 294 15601
rect 0 15429 624 15477
rect 0 15333 624 15381
rect 186 15209 294 15285
rect 0 15113 624 15161
rect 186 14955 294 15065
rect 0 14859 624 14907
rect 186 14735 294 14811
rect 0 14639 624 14687
rect 0 14543 624 14591
rect 186 14419 294 14495
rect 0 14323 624 14371
rect 186 14165 294 14275
rect 0 14069 624 14117
rect 186 13945 294 14021
rect 0 13849 624 13897
rect 0 13753 624 13801
rect 186 13629 294 13705
rect 0 13533 624 13581
rect 186 13375 294 13485
rect 0 13279 624 13327
rect 186 13155 294 13231
rect 0 13059 624 13107
rect 0 12963 624 13011
rect 186 12839 294 12915
rect 0 12743 624 12791
rect 186 12585 294 12695
rect 0 12489 624 12537
rect 186 12365 294 12441
rect 0 12269 624 12317
rect 0 12173 624 12221
rect 186 12049 294 12125
rect 0 11953 624 12001
rect 186 11795 294 11905
rect 0 11699 624 11747
rect 186 11575 294 11651
rect 0 11479 624 11527
rect 0 11383 624 11431
rect 186 11259 294 11335
rect 0 11163 624 11211
rect 186 11005 294 11115
rect 0 10909 624 10957
rect 186 10785 294 10861
rect 0 10689 624 10737
rect 0 10593 624 10641
rect 186 10469 294 10545
rect 0 10373 624 10421
rect 186 10215 294 10325
rect 0 10119 624 10167
rect 186 9995 294 10071
rect 0 9899 624 9947
rect 0 9803 624 9851
rect 186 9679 294 9755
rect 0 9583 624 9631
rect 186 9425 294 9535
rect 0 9329 624 9377
rect 186 9205 294 9281
rect 0 9109 624 9157
rect 0 9013 624 9061
rect 186 8889 294 8965
rect 0 8793 624 8841
rect 186 8635 294 8745
rect 0 8539 624 8587
rect 186 8415 294 8491
rect 0 8319 624 8367
rect 0 8223 624 8271
rect 186 8099 294 8175
rect 0 8003 624 8051
rect 186 7845 294 7955
rect 0 7749 624 7797
rect 186 7625 294 7701
rect 0 7529 624 7577
rect 0 7433 624 7481
rect 186 7309 294 7385
rect 0 7213 624 7261
rect 186 7055 294 7165
rect 0 6959 624 7007
rect 186 6835 294 6911
rect 0 6739 624 6787
rect 0 6643 624 6691
rect 186 6519 294 6595
rect 0 6423 624 6471
rect 186 6265 294 6375
rect 0 6169 624 6217
rect 186 6045 294 6121
rect 0 5949 624 5997
rect 0 5853 624 5901
rect 186 5729 294 5805
rect 0 5633 624 5681
rect 186 5475 294 5585
rect 0 5379 624 5427
rect 186 5255 294 5331
rect 0 5159 624 5207
rect 0 5063 624 5111
rect 186 4939 294 5015
rect 0 4843 624 4891
rect 186 4685 294 4795
rect 0 4589 624 4637
rect 186 4465 294 4541
rect 0 4369 624 4417
rect 0 4273 624 4321
rect 186 4149 294 4225
rect 0 4053 624 4101
rect 186 3895 294 4005
rect 0 3799 624 3847
rect 186 3675 294 3751
rect 0 3579 624 3627
rect 0 3483 624 3531
rect 186 3359 294 3435
rect 0 3263 624 3311
rect 186 3105 294 3215
rect 0 3009 624 3057
rect 186 2885 294 2961
rect 0 2789 624 2837
rect 0 2693 624 2741
rect 186 2569 294 2645
rect 0 2473 624 2521
rect 186 2315 294 2425
rect 0 2219 624 2267
rect 186 2095 294 2171
rect 0 1999 624 2047
rect 0 1903 624 1951
rect 186 1779 294 1855
rect 0 1683 624 1731
rect 186 1525 294 1635
rect 0 1429 624 1477
rect 186 1305 294 1381
rect 0 1209 624 1257
rect 0 1113 624 1161
rect 186 989 294 1065
rect 0 893 624 941
rect 186 735 294 845
rect 0 639 624 687
rect 186 515 294 591
rect 0 419 624 467
<< metal3 >>
rect 263 51862 361 51960
rect 263 180 361 278
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_1
timestamp 1626065694
transform 1 0 0 0 -1 52140
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_0
timestamp 1626065694
transform 1 0 0 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_0
timestamp 1626065694
transform 1 0 0 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_128
timestamp 1626065694
transform 1 0 0 0 -1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_127
timestamp 1626065694
transform 1 0 0 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_126
timestamp 1626065694
transform 1 0 0 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_125
timestamp 1626065694
transform 1 0 0 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_124
timestamp 1626065694
transform 1 0 0 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_123
timestamp 1626065694
transform 1 0 0 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_122
timestamp 1626065694
transform 1 0 0 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_121
timestamp 1626065694
transform 1 0 0 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_120
timestamp 1626065694
transform 1 0 0 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_119
timestamp 1626065694
transform 1 0 0 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_118
timestamp 1626065694
transform 1 0 0 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_117
timestamp 1626065694
transform 1 0 0 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_116
timestamp 1626065694
transform 1 0 0 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_115
timestamp 1626065694
transform 1 0 0 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_114
timestamp 1626065694
transform 1 0 0 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_113
timestamp 1626065694
transform 1 0 0 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_112
timestamp 1626065694
transform 1 0 0 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_111
timestamp 1626065694
transform 1 0 0 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_110
timestamp 1626065694
transform 1 0 0 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_109
timestamp 1626065694
transform 1 0 0 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_108
timestamp 1626065694
transform 1 0 0 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_107
timestamp 1626065694
transform 1 0 0 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_106
timestamp 1626065694
transform 1 0 0 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_105
timestamp 1626065694
transform 1 0 0 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_104
timestamp 1626065694
transform 1 0 0 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_103
timestamp 1626065694
transform 1 0 0 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_102
timestamp 1626065694
transform 1 0 0 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_101
timestamp 1626065694
transform 1 0 0 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_100
timestamp 1626065694
transform 1 0 0 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_99
timestamp 1626065694
transform 1 0 0 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_98
timestamp 1626065694
transform 1 0 0 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_97
timestamp 1626065694
transform 1 0 0 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_96
timestamp 1626065694
transform 1 0 0 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_95
timestamp 1626065694
transform 1 0 0 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_94
timestamp 1626065694
transform 1 0 0 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_93
timestamp 1626065694
transform 1 0 0 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_92
timestamp 1626065694
transform 1 0 0 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_91
timestamp 1626065694
transform 1 0 0 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_90
timestamp 1626065694
transform 1 0 0 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_89
timestamp 1626065694
transform 1 0 0 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_88
timestamp 1626065694
transform 1 0 0 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_87
timestamp 1626065694
transform 1 0 0 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_86
timestamp 1626065694
transform 1 0 0 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_85
timestamp 1626065694
transform 1 0 0 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_84
timestamp 1626065694
transform 1 0 0 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_83
timestamp 1626065694
transform 1 0 0 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_82
timestamp 1626065694
transform 1 0 0 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_81
timestamp 1626065694
transform 1 0 0 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_80
timestamp 1626065694
transform 1 0 0 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_79
timestamp 1626065694
transform 1 0 0 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_78
timestamp 1626065694
transform 1 0 0 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_77
timestamp 1626065694
transform 1 0 0 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_76
timestamp 1626065694
transform 1 0 0 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_75
timestamp 1626065694
transform 1 0 0 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_74
timestamp 1626065694
transform 1 0 0 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_73
timestamp 1626065694
transform 1 0 0 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_72
timestamp 1626065694
transform 1 0 0 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_71
timestamp 1626065694
transform 1 0 0 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_70
timestamp 1626065694
transform 1 0 0 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_69
timestamp 1626065694
transform 1 0 0 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_68
timestamp 1626065694
transform 1 0 0 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_67
timestamp 1626065694
transform 1 0 0 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_66
timestamp 1626065694
transform 1 0 0 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_65
timestamp 1626065694
transform 1 0 0 0 1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_64
timestamp 1626065694
transform 1 0 0 0 -1 51350
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_63
timestamp 1626065694
transform 1 0 0 0 1 51350
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_62
timestamp 1626065694
transform 1 0 0 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_61
timestamp 1626065694
transform 1 0 0 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_60
timestamp 1626065694
transform 1 0 0 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_59
timestamp 1626065694
transform 1 0 0 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_58
timestamp 1626065694
transform 1 0 0 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_57
timestamp 1626065694
transform 1 0 0 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_56
timestamp 1626065694
transform 1 0 0 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_55
timestamp 1626065694
transform 1 0 0 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_54
timestamp 1626065694
transform 1 0 0 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_53
timestamp 1626065694
transform 1 0 0 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_52
timestamp 1626065694
transform 1 0 0 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_51
timestamp 1626065694
transform 1 0 0 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_50
timestamp 1626065694
transform 1 0 0 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_49
timestamp 1626065694
transform 1 0 0 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_48
timestamp 1626065694
transform 1 0 0 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_47
timestamp 1626065694
transform 1 0 0 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_46
timestamp 1626065694
transform 1 0 0 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_45
timestamp 1626065694
transform 1 0 0 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_44
timestamp 1626065694
transform 1 0 0 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_43
timestamp 1626065694
transform 1 0 0 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_42
timestamp 1626065694
transform 1 0 0 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_41
timestamp 1626065694
transform 1 0 0 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_40
timestamp 1626065694
transform 1 0 0 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_39
timestamp 1626065694
transform 1 0 0 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_38
timestamp 1626065694
transform 1 0 0 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_37
timestamp 1626065694
transform 1 0 0 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_36
timestamp 1626065694
transform 1 0 0 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_35
timestamp 1626065694
transform 1 0 0 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_34
timestamp 1626065694
transform 1 0 0 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_33
timestamp 1626065694
transform 1 0 0 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_32
timestamp 1626065694
transform 1 0 0 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_31
timestamp 1626065694
transform 1 0 0 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_30
timestamp 1626065694
transform 1 0 0 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_29
timestamp 1626065694
transform 1 0 0 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_28
timestamp 1626065694
transform 1 0 0 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_27
timestamp 1626065694
transform 1 0 0 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_26
timestamp 1626065694
transform 1 0 0 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_25
timestamp 1626065694
transform 1 0 0 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_24
timestamp 1626065694
transform 1 0 0 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_23
timestamp 1626065694
transform 1 0 0 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_22
timestamp 1626065694
transform 1 0 0 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_21
timestamp 1626065694
transform 1 0 0 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_20
timestamp 1626065694
transform 1 0 0 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_19
timestamp 1626065694
transform 1 0 0 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_18
timestamp 1626065694
transform 1 0 0 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_17
timestamp 1626065694
transform 1 0 0 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_16
timestamp 1626065694
transform 1 0 0 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_15
timestamp 1626065694
transform 1 0 0 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_14
timestamp 1626065694
transform 1 0 0 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_13
timestamp 1626065694
transform 1 0 0 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_12
timestamp 1626065694
transform 1 0 0 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_11
timestamp 1626065694
transform 1 0 0 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_10
timestamp 1626065694
transform 1 0 0 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_9
timestamp 1626065694
transform 1 0 0 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_8
timestamp 1626065694
transform 1 0 0 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_7
timestamp 1626065694
transform 1 0 0 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_6
timestamp 1626065694
transform 1 0 0 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_5
timestamp 1626065694
transform 1 0 0 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_4
timestamp 1626065694
transform 1 0 0 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_3
timestamp 1626065694
transform 1 0 0 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_2
timestamp 1626065694
transform 1 0 0 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_1
timestamp 1626065694
transform 1 0 0 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_0
timestamp 1626065694
transform 1 0 0 0 1 790
box -42 -105 650 421
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_0
timestamp 1626065694
transform 1 0 279 0 1 192
box 0 0 66 74
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_1
timestamp 1626065694
transform 1 0 279 0 1 51874
box 0 0 66 74
<< labels >>
rlabel metal3 s 263 51862 361 51960 4 vdd
rlabel metal3 s 263 180 361 278 4 vdd
rlabel metal2 s 0 39033 624 39081 4 wl_0_97
rlabel metal2 s 0 39129 624 39177 4 wl_0_98
rlabel metal2 s 0 39823 624 39871 4 wl_0_99
rlabel metal2 s 0 39919 624 39967 4 wl_0_100
rlabel metal2 s 0 40613 624 40661 4 wl_0_101
rlabel metal2 s 0 40709 624 40757 4 wl_0_102
rlabel metal2 s 0 41403 624 41451 4 wl_0_103
rlabel metal2 s 0 41499 624 41547 4 wl_0_104
rlabel metal2 s 0 42193 624 42241 4 wl_0_105
rlabel metal2 s 0 42289 624 42337 4 wl_0_106
rlabel metal2 s 0 42983 624 43031 4 wl_0_107
rlabel metal2 s 0 43079 624 43127 4 wl_0_108
rlabel metal2 s 0 43773 624 43821 4 wl_0_109
rlabel metal2 s 0 43869 624 43917 4 wl_0_110
rlabel metal2 s 0 44563 624 44611 4 wl_0_111
rlabel metal2 s 0 44659 624 44707 4 wl_0_112
rlabel metal2 s 0 45353 624 45401 4 wl_0_113
rlabel metal2 s 0 45449 624 45497 4 wl_0_114
rlabel metal2 s 0 46143 624 46191 4 wl_0_115
rlabel metal2 s 0 46239 624 46287 4 wl_0_116
rlabel metal2 s 0 46933 624 46981 4 wl_0_117
rlabel metal2 s 0 47029 624 47077 4 wl_0_118
rlabel metal2 s 0 47723 624 47771 4 wl_0_119
rlabel metal2 s 0 47819 624 47867 4 wl_0_120
rlabel metal2 s 0 48513 624 48561 4 wl_0_121
rlabel metal2 s 0 48609 624 48657 4 wl_0_122
rlabel metal2 s 0 49303 624 49351 4 wl_0_123
rlabel metal2 s 0 49399 624 49447 4 wl_0_124
rlabel metal2 s 0 50093 624 50141 4 wl_0_125
rlabel metal2 s 0 50189 624 50237 4 wl_0_126
rlabel metal2 s 0 50883 624 50931 4 wl_0_127
rlabel metal2 s 0 50979 624 51027 4 wl_0_128
rlabel metal2 s 0 51673 624 51721 4 wl_0_129
rlabel metal2 s 0 39349 624 39397 4 wl_1_98
rlabel metal2 s 0 39603 624 39651 4 wl_1_99
rlabel metal2 s 0 40139 624 40187 4 wl_1_100
rlabel metal2 s 0 40393 624 40441 4 wl_1_101
rlabel metal2 s 0 40929 624 40977 4 wl_1_102
rlabel metal2 s 0 41183 624 41231 4 wl_1_103
rlabel metal2 s 0 41719 624 41767 4 wl_1_104
rlabel metal2 s 0 41973 624 42021 4 wl_1_105
rlabel metal2 s 0 42509 624 42557 4 wl_1_106
rlabel metal2 s 0 42763 624 42811 4 wl_1_107
rlabel metal2 s 0 43299 624 43347 4 wl_1_108
rlabel metal2 s 0 43553 624 43601 4 wl_1_109
rlabel metal2 s 0 44089 624 44137 4 wl_1_110
rlabel metal2 s 0 44343 624 44391 4 wl_1_111
rlabel metal2 s 0 44879 624 44927 4 wl_1_112
rlabel metal2 s 0 45133 624 45181 4 wl_1_113
rlabel metal2 s 0 45669 624 45717 4 wl_1_114
rlabel metal2 s 0 45923 624 45971 4 wl_1_115
rlabel metal2 s 0 46459 624 46507 4 wl_1_116
rlabel metal2 s 0 46713 624 46761 4 wl_1_117
rlabel metal2 s 0 47249 624 47297 4 wl_1_118
rlabel metal2 s 0 47503 624 47551 4 wl_1_119
rlabel metal2 s 0 48039 624 48087 4 wl_1_120
rlabel metal2 s 0 48293 624 48341 4 wl_1_121
rlabel metal2 s 0 48829 624 48877 4 wl_1_122
rlabel metal2 s 0 49083 624 49131 4 wl_1_123
rlabel metal2 s 0 49619 624 49667 4 wl_1_124
rlabel metal2 s 0 49873 624 49921 4 wl_1_125
rlabel metal2 s 0 50409 624 50457 4 wl_1_126
rlabel metal2 s 0 50663 624 50711 4 wl_1_127
rlabel metal2 s 0 51199 624 51247 4 wl_1_128
rlabel metal2 s 0 51453 624 51501 4 wl_1_129
rlabel metal2 s 0 26173 624 26221 4 wl_1_65
rlabel metal2 s 0 26709 624 26757 4 wl_1_66
rlabel metal2 s 0 26963 624 27011 4 wl_1_67
rlabel metal2 s 0 27499 624 27547 4 wl_1_68
rlabel metal2 s 0 27753 624 27801 4 wl_1_69
rlabel metal2 s 0 28289 624 28337 4 wl_1_70
rlabel metal2 s 0 28543 624 28591 4 wl_1_71
rlabel metal2 s 0 29079 624 29127 4 wl_1_72
rlabel metal2 s 0 29333 624 29381 4 wl_1_73
rlabel metal2 s 0 29869 624 29917 4 wl_1_74
rlabel metal2 s 0 30123 624 30171 4 wl_1_75
rlabel metal2 s 0 30659 624 30707 4 wl_1_76
rlabel metal2 s 0 30913 624 30961 4 wl_1_77
rlabel metal2 s 0 31449 624 31497 4 wl_1_78
rlabel metal2 s 0 31703 624 31751 4 wl_1_79
rlabel metal2 s 0 32239 624 32287 4 wl_1_80
rlabel metal2 s 0 32493 624 32541 4 wl_1_81
rlabel metal2 s 0 33029 624 33077 4 wl_1_82
rlabel metal2 s 0 33283 624 33331 4 wl_1_83
rlabel metal2 s 0 33819 624 33867 4 wl_1_84
rlabel metal2 s 0 34073 624 34121 4 wl_1_85
rlabel metal2 s 0 34609 624 34657 4 wl_1_86
rlabel metal2 s 0 34863 624 34911 4 wl_1_87
rlabel metal2 s 0 35399 624 35447 4 wl_1_88
rlabel metal2 s 0 35653 624 35701 4 wl_1_89
rlabel metal2 s 0 36189 624 36237 4 wl_1_90
rlabel metal2 s 0 36443 624 36491 4 wl_1_91
rlabel metal2 s 0 36979 624 37027 4 wl_1_92
rlabel metal2 s 0 37233 624 37281 4 wl_1_93
rlabel metal2 s 0 37769 624 37817 4 wl_1_94
rlabel metal2 s 0 38023 624 38071 4 wl_1_95
rlabel metal2 s 0 38559 624 38607 4 wl_1_96
rlabel metal2 s 0 38813 624 38861 4 wl_1_97
rlabel metal2 s 0 26489 624 26537 4 wl_0_66
rlabel metal2 s 0 27183 624 27231 4 wl_0_67
rlabel metal2 s 0 27279 624 27327 4 wl_0_68
rlabel metal2 s 0 27973 624 28021 4 wl_0_69
rlabel metal2 s 0 28069 624 28117 4 wl_0_70
rlabel metal2 s 0 28763 624 28811 4 wl_0_71
rlabel metal2 s 0 28859 624 28907 4 wl_0_72
rlabel metal2 s 0 29553 624 29601 4 wl_0_73
rlabel metal2 s 0 29649 624 29697 4 wl_0_74
rlabel metal2 s 0 30343 624 30391 4 wl_0_75
rlabel metal2 s 0 30439 624 30487 4 wl_0_76
rlabel metal2 s 0 31133 624 31181 4 wl_0_77
rlabel metal2 s 0 31229 624 31277 4 wl_0_78
rlabel metal2 s 0 31923 624 31971 4 wl_0_79
rlabel metal2 s 0 32019 624 32067 4 wl_0_80
rlabel metal2 s 0 32713 624 32761 4 wl_0_81
rlabel metal2 s 0 32809 624 32857 4 wl_0_82
rlabel metal2 s 0 33503 624 33551 4 wl_0_83
rlabel metal2 s 0 33599 624 33647 4 wl_0_84
rlabel metal2 s 0 34293 624 34341 4 wl_0_85
rlabel metal2 s 0 34389 624 34437 4 wl_0_86
rlabel metal2 s 0 35083 624 35131 4 wl_0_87
rlabel metal2 s 0 35179 624 35227 4 wl_0_88
rlabel metal2 s 0 35873 624 35921 4 wl_0_89
rlabel metal2 s 0 35969 624 36017 4 wl_0_90
rlabel metal2 s 0 36663 624 36711 4 wl_0_91
rlabel metal2 s 0 36759 624 36807 4 wl_0_92
rlabel metal2 s 0 37453 624 37501 4 wl_0_93
rlabel metal2 s 0 37549 624 37597 4 wl_0_94
rlabel metal2 s 0 38243 624 38291 4 wl_0_95
rlabel metal2 s 0 38339 624 38387 4 wl_0_96
rlabel metal2 s 0 26393 624 26441 4 wl_0_65
rlabel metal2 s 186 47599 294 47675 4 gnd
rlabel metal2 s 186 29175 294 29285 4 gnd
rlabel metal2 s 186 27375 294 27451 4 gnd
rlabel metal2 s 186 49495 294 49571 4 gnd
rlabel metal2 s 186 27849 294 27925 4 gnd
rlabel metal2 s 186 42069 294 42145 4 gnd
rlabel metal2 s 186 44755 294 44831 4 gnd
rlabel metal2 s 186 46019 294 46095 4 gnd
rlabel metal2 s 186 32589 294 32665 4 gnd
rlabel metal2 s 186 33695 294 33771 4 gnd
rlabel metal2 s 186 41025 294 41135 4 gnd
rlabel metal2 s 186 31009 294 31085 4 gnd
rlabel metal2 s 186 30219 294 30295 4 gnd
rlabel metal2 s 186 29745 294 29821 4 gnd
rlabel metal2 s 186 38435 294 38511 4 gnd
rlabel metal2 s 186 40805 294 40881 4 gnd
rlabel metal2 s 186 42859 294 42935 4 gnd
rlabel metal2 s 186 48705 294 48781 4 gnd
rlabel metal2 s 186 36539 294 36615 4 gnd
rlabel metal2 s 186 33379 294 33455 4 gnd
rlabel metal2 s 186 45545 294 45621 4 gnd
rlabel metal2 s 186 43395 294 43505 4 gnd
rlabel metal2 s 186 51075 294 51151 4 gnd
rlabel metal2 s 186 34959 294 35035 4 gnd
rlabel metal2 s 186 31545 294 31655 4 gnd
rlabel metal2 s 186 44185 294 44295 4 gnd
rlabel metal2 s 186 35749 294 35825 4 gnd
rlabel metal2 s 186 34169 294 34245 4 gnd
rlabel metal2 s 186 45229 294 45305 4 gnd
rlabel metal2 s 186 43649 294 43725 4 gnd
rlabel metal2 s 186 31325 294 31401 4 gnd
rlabel metal2 s 186 36065 294 36141 4 gnd
rlabel metal2 s 186 30535 294 30611 4 gnd
rlabel metal2 s 186 40489 294 40565 4 gnd
rlabel metal2 s 186 28165 294 28241 4 gnd
rlabel metal2 s 186 36855 294 36931 4 gnd
rlabel metal2 s 186 33125 294 33235 4 gnd
rlabel metal2 s 186 51549 294 51625 4 gnd
rlabel metal2 s 186 26805 294 26915 4 gnd
rlabel metal2 s 186 41595 294 41671 4 gnd
rlabel metal2 s 186 44439 294 44515 4 gnd
rlabel metal2 s 186 39699 294 39775 4 gnd
rlabel metal2 s 186 34705 294 34815 4 gnd
rlabel metal2 s 186 37645 294 37721 4 gnd
rlabel metal2 s 186 26585 294 26661 4 gnd
rlabel metal2 s 186 48135 294 48245 4 gnd
rlabel metal2 s 186 36285 294 36395 4 gnd
rlabel metal2 s 186 26269 294 26345 4 gnd
rlabel metal2 s 186 32905 294 32981 4 gnd
rlabel metal2 s 186 49179 294 49255 4 gnd
rlabel metal2 s 186 32335 294 32445 4 gnd
rlabel metal2 s 186 37329 294 37405 4 gnd
rlabel metal2 s 186 31799 294 31875 4 gnd
rlabel metal2 s 186 38655 294 38765 4 gnd
rlabel metal2 s 186 38119 294 38195 4 gnd
rlabel metal2 s 186 41279 294 41355 4 gnd
rlabel metal2 s 186 45765 294 45875 4 gnd
rlabel metal2 s 186 49715 294 49825 4 gnd
rlabel metal2 s 186 44975 294 45085 4 gnd
rlabel metal2 s 186 28385 294 28495 4 gnd
rlabel metal2 s 186 42605 294 42715 4 gnd
rlabel metal2 s 186 46335 294 46411 4 gnd
rlabel metal2 s 186 47915 294 47991 4 gnd
rlabel metal2 s 186 40015 294 40091 4 gnd
rlabel metal2 s 186 48925 294 49035 4 gnd
rlabel metal2 s 186 47125 294 47201 4 gnd
rlabel metal2 s 186 50285 294 50361 4 gnd
rlabel metal2 s 186 49969 294 50045 4 gnd
rlabel metal2 s 186 39445 294 39555 4 gnd
rlabel metal2 s 186 28639 294 28715 4 gnd
rlabel metal2 s 186 50505 294 50615 4 gnd
rlabel metal2 s 186 37075 294 37185 4 gnd
rlabel metal2 s 186 29429 294 29505 4 gnd
rlabel metal2 s 186 48389 294 48465 4 gnd
rlabel metal2 s 186 35275 294 35351 4 gnd
rlabel metal2 s 186 43175 294 43251 4 gnd
rlabel metal2 s 186 27059 294 27135 4 gnd
rlabel metal2 s 186 50759 294 50835 4 gnd
rlabel metal2 s 186 38909 294 38985 4 gnd
rlabel metal2 s 186 28955 294 29031 4 gnd
rlabel metal2 s 186 47345 294 47455 4 gnd
rlabel metal2 s 186 33915 294 34025 4 gnd
rlabel metal2 s 186 29965 294 30075 4 gnd
rlabel metal2 s 186 41815 294 41925 4 gnd
rlabel metal2 s 186 43965 294 44041 4 gnd
rlabel metal2 s 186 27595 294 27705 4 gnd
rlabel metal2 s 186 39225 294 39301 4 gnd
rlabel metal2 s 186 46555 294 46665 4 gnd
rlabel metal2 s 186 42385 294 42461 4 gnd
rlabel metal2 s 186 30755 294 30865 4 gnd
rlabel metal2 s 186 51295 294 51405 4 gnd
rlabel metal2 s 186 46809 294 46885 4 gnd
rlabel metal2 s 186 37865 294 37975 4 gnd
rlabel metal2 s 186 34485 294 34561 4 gnd
rlabel metal2 s 186 32115 294 32191 4 gnd
rlabel metal2 s 186 35495 294 35605 4 gnd
rlabel metal2 s 186 40235 294 40345 4 gnd
rlabel metal2 s 186 16535 294 16645 4 gnd
rlabel metal2 s 186 17579 294 17655 4 gnd
rlabel metal2 s 186 22855 294 22965 4 gnd
rlabel metal2 s 186 16315 294 16391 4 gnd
rlabel metal2 s 186 7845 294 7955 4 gnd
rlabel metal2 s 186 8635 294 8745 4 gnd
rlabel metal2 s 186 8099 294 8175 4 gnd
rlabel metal2 s 186 9425 294 9535 4 gnd
rlabel metal2 s 186 2095 294 2171 4 gnd
rlabel metal2 s 186 9679 294 9755 4 gnd
rlabel metal2 s 186 23425 294 23501 4 gnd
rlabel metal2 s 186 5729 294 5805 4 gnd
rlabel metal2 s 186 1779 294 1855 4 gnd
rlabel metal2 s 186 25225 294 25335 4 gnd
rlabel metal2 s 186 18115 294 18225 4 gnd
rlabel metal2 s 186 20485 294 20595 4 gnd
rlabel metal2 s 186 2315 294 2425 4 gnd
rlabel metal2 s 186 15745 294 15855 4 gnd
rlabel metal2 s 186 23109 294 23185 4 gnd
rlabel metal2 s 186 4939 294 5015 4 gnd
rlabel metal2 s 186 15525 294 15601 4 gnd
rlabel metal2 s 186 21529 294 21605 4 gnd
rlabel metal2 s 186 4465 294 4541 4 gnd
rlabel metal2 s 186 6265 294 6375 4 gnd
rlabel metal2 s 186 23645 294 23755 4 gnd
rlabel metal2 s 186 13629 294 13705 4 gnd
rlabel metal2 s 186 21055 294 21131 4 gnd
rlabel metal2 s 186 14735 294 14811 4 gnd
rlabel metal2 s 186 15999 294 16075 4 gnd
rlabel metal2 s 186 3675 294 3751 4 gnd
rlabel metal2 s 186 18685 294 18761 4 gnd
rlabel metal2 s 186 26015 294 26125 4 gnd
rlabel metal2 s 186 2885 294 2961 4 gnd
rlabel metal2 s 186 12839 294 12915 4 gnd
rlabel metal2 s 186 12049 294 12125 4 gnd
rlabel metal2 s 186 25795 294 25871 4 gnd
rlabel metal2 s 186 4685 294 4795 4 gnd
rlabel metal2 s 186 21845 294 21921 4 gnd
rlabel metal2 s 186 17105 294 17181 4 gnd
rlabel metal2 s 186 12365 294 12441 4 gnd
rlabel metal2 s 186 14955 294 15065 4 gnd
rlabel metal2 s 186 1305 294 1381 4 gnd
rlabel metal2 s 186 5475 294 5585 4 gnd
rlabel metal2 s 186 10469 294 10545 4 gnd
rlabel metal2 s 186 7309 294 7385 4 gnd
rlabel metal2 s 186 12585 294 12695 4 gnd
rlabel metal2 s 186 8889 294 8965 4 gnd
rlabel metal2 s 186 18905 294 19015 4 gnd
rlabel metal2 s 186 24435 294 24545 4 gnd
rlabel metal2 s 186 735 294 845 4 gnd
rlabel metal2 s 186 13375 294 13485 4 gnd
rlabel metal2 s 186 515 294 591 4 gnd
rlabel metal2 s 186 17895 294 17971 4 gnd
rlabel metal2 s 186 13155 294 13231 4 gnd
rlabel metal2 s 186 6835 294 6911 4 gnd
rlabel metal2 s 186 24215 294 24291 4 gnd
rlabel metal2 s 186 14165 294 14275 4 gnd
rlabel metal2 s 186 7625 294 7701 4 gnd
rlabel metal2 s 186 21275 294 21385 4 gnd
rlabel metal2 s 186 19695 294 19805 4 gnd
rlabel metal2 s 186 24689 294 24765 4 gnd
rlabel metal2 s 186 19159 294 19235 4 gnd
rlabel metal2 s 186 11575 294 11651 4 gnd
rlabel metal2 s 186 11005 294 11115 4 gnd
rlabel metal2 s 186 11259 294 11335 4 gnd
rlabel metal2 s 186 3895 294 4005 4 gnd
rlabel metal2 s 186 19949 294 20025 4 gnd
rlabel metal2 s 186 17325 294 17435 4 gnd
rlabel metal2 s 186 20739 294 20815 4 gnd
rlabel metal2 s 186 22065 294 22175 4 gnd
rlabel metal2 s 186 25005 294 25081 4 gnd
rlabel metal2 s 186 16789 294 16865 4 gnd
rlabel metal2 s 186 2569 294 2645 4 gnd
rlabel metal2 s 186 3359 294 3435 4 gnd
rlabel metal2 s 186 1525 294 1635 4 gnd
rlabel metal2 s 186 4149 294 4225 4 gnd
rlabel metal2 s 186 989 294 1065 4 gnd
rlabel metal2 s 186 3105 294 3215 4 gnd
rlabel metal2 s 186 14419 294 14495 4 gnd
rlabel metal2 s 186 13945 294 14021 4 gnd
rlabel metal2 s 186 25479 294 25555 4 gnd
rlabel metal2 s 186 18369 294 18445 4 gnd
rlabel metal2 s 186 7055 294 7165 4 gnd
rlabel metal2 s 186 22319 294 22395 4 gnd
rlabel metal2 s 186 19475 294 19551 4 gnd
rlabel metal2 s 186 15209 294 15285 4 gnd
rlabel metal2 s 186 11795 294 11905 4 gnd
rlabel metal2 s 186 9205 294 9281 4 gnd
rlabel metal2 s 186 20265 294 20341 4 gnd
rlabel metal2 s 186 10215 294 10325 4 gnd
rlabel metal2 s 186 6519 294 6595 4 gnd
rlabel metal2 s 186 8415 294 8491 4 gnd
rlabel metal2 s 186 9995 294 10071 4 gnd
rlabel metal2 s 186 22635 294 22711 4 gnd
rlabel metal2 s 186 23899 294 23975 4 gnd
rlabel metal2 s 186 6045 294 6121 4 gnd
rlabel metal2 s 186 5255 294 5331 4 gnd
rlabel metal2 s 186 10785 294 10861 4 gnd
rlabel metal2 s 0 13753 624 13801 4 wl_0_33
rlabel metal2 s 0 13849 624 13897 4 wl_0_34
rlabel metal2 s 0 14543 624 14591 4 wl_0_35
rlabel metal2 s 0 14639 624 14687 4 wl_0_36
rlabel metal2 s 0 15333 624 15381 4 wl_0_37
rlabel metal2 s 0 15429 624 15477 4 wl_0_38
rlabel metal2 s 0 16123 624 16171 4 wl_0_39
rlabel metal2 s 0 16219 624 16267 4 wl_0_40
rlabel metal2 s 0 16913 624 16961 4 wl_0_41
rlabel metal2 s 0 17009 624 17057 4 wl_0_42
rlabel metal2 s 0 17703 624 17751 4 wl_0_43
rlabel metal2 s 0 17799 624 17847 4 wl_0_44
rlabel metal2 s 0 18493 624 18541 4 wl_0_45
rlabel metal2 s 0 18589 624 18637 4 wl_0_46
rlabel metal2 s 0 19283 624 19331 4 wl_0_47
rlabel metal2 s 0 19379 624 19427 4 wl_0_48
rlabel metal2 s 0 20073 624 20121 4 wl_0_49
rlabel metal2 s 0 20169 624 20217 4 wl_0_50
rlabel metal2 s 0 20863 624 20911 4 wl_0_51
rlabel metal2 s 0 20959 624 21007 4 wl_0_52
rlabel metal2 s 0 21653 624 21701 4 wl_0_53
rlabel metal2 s 0 21749 624 21797 4 wl_0_54
rlabel metal2 s 0 22443 624 22491 4 wl_0_55
rlabel metal2 s 0 22539 624 22587 4 wl_0_56
rlabel metal2 s 0 23233 624 23281 4 wl_0_57
rlabel metal2 s 0 23329 624 23377 4 wl_0_58
rlabel metal2 s 0 24023 624 24071 4 wl_0_59
rlabel metal2 s 0 24119 624 24167 4 wl_0_60
rlabel metal2 s 0 24813 624 24861 4 wl_0_61
rlabel metal2 s 0 24909 624 24957 4 wl_0_62
rlabel metal2 s 0 25603 624 25651 4 wl_0_63
rlabel metal2 s 0 25699 624 25747 4 wl_0_64
rlabel metal2 s 0 13279 624 13327 4 wl_1_32
rlabel metal2 s 0 13533 624 13581 4 wl_1_33
rlabel metal2 s 0 14069 624 14117 4 wl_1_34
rlabel metal2 s 0 14323 624 14371 4 wl_1_35
rlabel metal2 s 0 14859 624 14907 4 wl_1_36
rlabel metal2 s 0 15113 624 15161 4 wl_1_37
rlabel metal2 s 0 15649 624 15697 4 wl_1_38
rlabel metal2 s 0 15903 624 15951 4 wl_1_39
rlabel metal2 s 0 16439 624 16487 4 wl_1_40
rlabel metal2 s 0 16693 624 16741 4 wl_1_41
rlabel metal2 s 0 17229 624 17277 4 wl_1_42
rlabel metal2 s 0 17483 624 17531 4 wl_1_43
rlabel metal2 s 0 18019 624 18067 4 wl_1_44
rlabel metal2 s 0 18273 624 18321 4 wl_1_45
rlabel metal2 s 0 18809 624 18857 4 wl_1_46
rlabel metal2 s 0 19063 624 19111 4 wl_1_47
rlabel metal2 s 0 19599 624 19647 4 wl_1_48
rlabel metal2 s 0 19853 624 19901 4 wl_1_49
rlabel metal2 s 0 20389 624 20437 4 wl_1_50
rlabel metal2 s 0 20643 624 20691 4 wl_1_51
rlabel metal2 s 0 21179 624 21227 4 wl_1_52
rlabel metal2 s 0 21433 624 21481 4 wl_1_53
rlabel metal2 s 0 21969 624 22017 4 wl_1_54
rlabel metal2 s 0 22223 624 22271 4 wl_1_55
rlabel metal2 s 0 22759 624 22807 4 wl_1_56
rlabel metal2 s 0 23013 624 23061 4 wl_1_57
rlabel metal2 s 0 23549 624 23597 4 wl_1_58
rlabel metal2 s 0 23803 624 23851 4 wl_1_59
rlabel metal2 s 0 24339 624 24387 4 wl_1_60
rlabel metal2 s 0 24593 624 24641 4 wl_1_61
rlabel metal2 s 0 25129 624 25177 4 wl_1_62
rlabel metal2 s 0 25383 624 25431 4 wl_1_63
rlabel metal2 s 0 25919 624 25967 4 wl_1_64
rlabel metal2 s 0 639 624 687 4 wl_1_0
rlabel metal2 s 0 893 624 941 4 wl_1_1
rlabel metal2 s 0 1429 624 1477 4 wl_1_2
rlabel metal2 s 0 1683 624 1731 4 wl_1_3
rlabel metal2 s 0 2219 624 2267 4 wl_1_4
rlabel metal2 s 0 2473 624 2521 4 wl_1_5
rlabel metal2 s 0 3009 624 3057 4 wl_1_6
rlabel metal2 s 0 3263 624 3311 4 wl_1_7
rlabel metal2 s 0 3799 624 3847 4 wl_1_8
rlabel metal2 s 0 4053 624 4101 4 wl_1_9
rlabel metal2 s 0 4589 624 4637 4 wl_1_10
rlabel metal2 s 0 4843 624 4891 4 wl_1_11
rlabel metal2 s 0 5379 624 5427 4 wl_1_12
rlabel metal2 s 0 5633 624 5681 4 wl_1_13
rlabel metal2 s 0 6169 624 6217 4 wl_1_14
rlabel metal2 s 0 6423 624 6471 4 wl_1_15
rlabel metal2 s 0 6959 624 7007 4 wl_1_16
rlabel metal2 s 0 7213 624 7261 4 wl_1_17
rlabel metal2 s 0 7749 624 7797 4 wl_1_18
rlabel metal2 s 0 8003 624 8051 4 wl_1_19
rlabel metal2 s 0 8539 624 8587 4 wl_1_20
rlabel metal2 s 0 8793 624 8841 4 wl_1_21
rlabel metal2 s 0 9329 624 9377 4 wl_1_22
rlabel metal2 s 0 9583 624 9631 4 wl_1_23
rlabel metal2 s 0 10119 624 10167 4 wl_1_24
rlabel metal2 s 0 10373 624 10421 4 wl_1_25
rlabel metal2 s 0 10909 624 10957 4 wl_1_26
rlabel metal2 s 0 11163 624 11211 4 wl_1_27
rlabel metal2 s 0 11699 624 11747 4 wl_1_28
rlabel metal2 s 0 11953 624 12001 4 wl_1_29
rlabel metal2 s 0 12489 624 12537 4 wl_1_30
rlabel metal2 s 0 12743 624 12791 4 wl_1_31
rlabel metal2 s 0 13059 624 13107 4 wl_0_32
rlabel metal2 s 0 419 624 467 4 wl_0_0
rlabel metal2 s 0 1113 624 1161 4 wl_0_1
rlabel metal2 s 0 1209 624 1257 4 wl_0_2
rlabel metal2 s 0 1903 624 1951 4 wl_0_3
rlabel metal2 s 0 1999 624 2047 4 wl_0_4
rlabel metal2 s 0 2693 624 2741 4 wl_0_5
rlabel metal2 s 0 2789 624 2837 4 wl_0_6
rlabel metal2 s 0 3483 624 3531 4 wl_0_7
rlabel metal2 s 0 3579 624 3627 4 wl_0_8
rlabel metal2 s 0 4273 624 4321 4 wl_0_9
rlabel metal2 s 0 4369 624 4417 4 wl_0_10
rlabel metal2 s 0 5063 624 5111 4 wl_0_11
rlabel metal2 s 0 5159 624 5207 4 wl_0_12
rlabel metal2 s 0 5853 624 5901 4 wl_0_13
rlabel metal2 s 0 5949 624 5997 4 wl_0_14
rlabel metal2 s 0 6643 624 6691 4 wl_0_15
rlabel metal2 s 0 6739 624 6787 4 wl_0_16
rlabel metal2 s 0 7433 624 7481 4 wl_0_17
rlabel metal2 s 0 7529 624 7577 4 wl_0_18
rlabel metal2 s 0 8223 624 8271 4 wl_0_19
rlabel metal2 s 0 8319 624 8367 4 wl_0_20
rlabel metal2 s 0 9013 624 9061 4 wl_0_21
rlabel metal2 s 0 9109 624 9157 4 wl_0_22
rlabel metal2 s 0 9803 624 9851 4 wl_0_23
rlabel metal2 s 0 9899 624 9947 4 wl_0_24
rlabel metal2 s 0 10593 624 10641 4 wl_0_25
rlabel metal2 s 0 10689 624 10737 4 wl_0_26
rlabel metal2 s 0 11383 624 11431 4 wl_0_27
rlabel metal2 s 0 11479 624 11527 4 wl_0_28
rlabel metal2 s 0 12173 624 12221 4 wl_0_29
rlabel metal2 s 0 12269 624 12317 4 wl_0_30
rlabel metal2 s 0 12963 624 13011 4 wl_0_31
rlabel metal1 s 222 35629 258 35970 4 vdd
rlabel metal1 s 222 45899 258 46240 4 vdd
rlabel metal1 s 222 46980 258 47321 4 vdd
rlabel metal1 s 222 34049 258 34390 4 vdd
rlabel metal1 s 222 38290 258 38631 4 vdd
rlabel metal1 s 222 46190 258 46531 4 vdd
rlabel metal1 s 222 27230 258 27571 4 vdd
rlabel metal1 s 222 30889 258 31230 4 vdd
rlabel metal1 s 222 45400 258 45741 4 vdd
rlabel metal1 s 222 26939 258 27280 4 vdd
rlabel metal1 s 222 36710 258 37051 4 vdd
rlabel metal1 s 222 35130 258 35471 4 vdd
rlabel metal1 s 222 39579 258 39920 4 vdd
rlabel metal1 s 222 50639 258 50980 4 vdd
rlabel metal1 s 222 31679 258 32020 4 vdd
rlabel metal1 s 222 33550 258 33891 4 vdd
rlabel metal1 s 222 51429 258 51770 4 vdd
rlabel metal1 s 222 43030 258 43371 4 vdd
rlabel metal1 s 222 30390 258 30731 4 vdd
rlabel metal1 s 222 39870 258 40211 4 vdd
rlabel metal1 s 222 42739 258 43080 4 vdd
rlabel metal1 s 222 37500 258 37841 4 vdd
rlabel metal1 s 222 29309 258 29650 4 vdd
rlabel metal1 s 222 50140 258 50481 4 vdd
rlabel metal1 s 222 31180 258 31521 4 vdd
rlabel metal1 s 222 47770 258 48111 4 vdd
rlabel metal1 s 222 31970 258 32311 4 vdd
rlabel metal1 s 222 32469 258 32810 4 vdd
rlabel metal1 s 222 43820 258 44161 4 vdd
rlabel metal1 s 222 26149 258 26490 4 vdd
rlabel metal1 s 222 48560 258 48901 4 vdd
rlabel metal1 s 222 50930 258 51271 4 vdd
rlabel metal1 s 222 30099 258 30440 4 vdd
rlabel metal1 s 222 37209 258 37550 4 vdd
rlabel metal1 s 222 41159 258 41500 4 vdd
rlabel metal1 s 222 40660 258 41001 4 vdd
rlabel metal1 s 222 46689 258 47030 4 vdd
rlabel metal1 s 222 28810 258 29151 4 vdd
rlabel metal1 s 222 28519 258 28860 4 vdd
rlabel metal1 s 222 29600 258 29941 4 vdd
rlabel metal1 s 222 41450 258 41791 4 vdd
rlabel metal1 s 222 36419 258 36760 4 vdd
rlabel metal1 s 222 45109 258 45450 4 vdd
rlabel metal1 s 222 48269 258 48610 4 vdd
rlabel metal1 s 222 37999 258 38340 4 vdd
rlabel metal1 s 222 44610 258 44951 4 vdd
rlabel metal1 s 222 35920 258 36261 4 vdd
rlabel metal1 s 222 41949 258 42290 4 vdd
rlabel metal1 s 222 34340 258 34681 4 vdd
rlabel metal1 s 222 40369 258 40710 4 vdd
rlabel metal1 s 222 42240 258 42581 4 vdd
rlabel metal1 s 222 49350 258 49691 4 vdd
rlabel metal1 s 222 39080 258 39421 4 vdd
rlabel metal1 s 222 47479 258 47820 4 vdd
rlabel metal1 s 222 27729 258 28070 4 vdd
rlabel metal1 s 222 38789 258 39130 4 vdd
rlabel metal1 s 222 34839 258 35180 4 vdd
rlabel metal1 s 222 26440 258 26781 4 vdd
rlabel metal1 s 222 28020 258 28361 4 vdd
rlabel metal1 s 222 33259 258 33600 4 vdd
rlabel metal1 s 222 43529 258 43870 4 vdd
rlabel metal1 s 222 32760 258 33101 4 vdd
rlabel metal1 s 222 49849 258 50190 4 vdd
rlabel metal1 s 222 44319 258 44660 4 vdd
rlabel metal1 s 222 49059 258 49400 4 vdd
rlabel metal1 s 78 0 114 52140 4 bl_0_0
rlabel metal1 s 222 4819 258 5160 4 vdd
rlabel metal1 s 222 20120 258 20461 4 vdd
rlabel metal1 s 222 14299 258 14640 4 vdd
rlabel metal1 s 222 22199 258 22540 4 vdd
rlabel metal1 s 222 11430 258 11771 4 vdd
rlabel metal1 s 222 9559 258 9900 4 vdd
rlabel metal1 s 222 8769 258 9110 4 vdd
rlabel metal1 s 222 9060 258 9401 4 vdd
rlabel metal1 s 222 1950 258 2291 4 vdd
rlabel metal1 s 222 11139 258 11480 4 vdd
rlabel metal1 s 222 17750 258 18091 4 vdd
rlabel metal1 s 222 13010 258 13351 4 vdd
rlabel metal1 s 222 2740 258 3081 4 vdd
rlabel metal1 s 222 12719 258 13060 4 vdd
rlabel metal1 s 222 25650 258 25991 4 vdd
rlabel metal1 s 222 7480 258 7821 4 vdd
rlabel metal1 s 222 869 258 1210 4 vdd
rlabel metal1 s 222 5900 258 6241 4 vdd
rlabel metal1 s 222 11929 258 12270 4 vdd
rlabel metal1 s 222 16669 258 17010 4 vdd
rlabel metal1 s 222 19039 258 19380 4 vdd
rlabel metal1 s 222 23280 258 23621 4 vdd
rlabel metal1 s 222 19330 258 19671 4 vdd
rlabel metal1 s 222 15380 258 15721 4 vdd
rlabel metal1 s 222 4029 258 4370 4 vdd
rlabel metal1 s 222 15879 258 16220 4 vdd
rlabel metal1 s 222 20910 258 21251 4 vdd
rlabel metal1 s 222 3530 258 3871 4 vdd
rlabel metal1 s 222 14590 258 14931 4 vdd
rlabel metal1 s 222 12220 258 12561 4 vdd
rlabel metal1 s 222 4320 258 4661 4 vdd
rlabel metal1 s 222 24070 258 24411 4 vdd
rlabel metal1 s 150 0 186 52140 4 br_0_0
rlabel metal1 s 222 18540 258 18881 4 vdd
rlabel metal1 s 222 24569 258 24910 4 vdd
rlabel metal1 s 222 10640 258 10981 4 vdd
rlabel metal1 s 222 21700 258 22041 4 vdd
rlabel metal1 s 222 3239 258 3580 4 vdd
rlabel metal1 s 222 20619 258 20960 4 vdd
rlabel metal1 s 222 23779 258 24120 4 vdd
rlabel metal1 s 294 0 330 52140 4 bl_1_0
rlabel metal1 s 222 6690 258 7031 4 vdd
rlabel metal1 s 222 25359 258 25700 4 vdd
rlabel metal1 s 222 22989 258 23330 4 vdd
rlabel metal1 s 222 16170 258 16511 4 vdd
rlabel metal1 s 366 0 402 52140 4 br_1_0
rlabel metal1 s 222 9850 258 10191 4 vdd
rlabel metal1 s 222 18249 258 18590 4 vdd
rlabel metal1 s 222 13509 258 13850 4 vdd
rlabel metal1 s 222 24860 258 25201 4 vdd
rlabel metal1 s 222 6399 258 6740 4 vdd
rlabel metal1 s 222 7979 258 8320 4 vdd
rlabel metal1 s 222 370 258 711 4 vdd
rlabel metal1 s 222 22490 258 22831 4 vdd
rlabel metal1 s 222 8270 258 8611 4 vdd
rlabel metal1 s 222 15089 258 15430 4 vdd
rlabel metal1 s 222 16960 258 17301 4 vdd
rlabel metal1 s 222 1160 258 1501 4 vdd
rlabel metal1 s 222 19829 258 20170 4 vdd
rlabel metal1 s 222 10349 258 10690 4 vdd
rlabel metal1 s 222 7189 258 7530 4 vdd
rlabel metal1 s 222 21409 258 21750 4 vdd
rlabel metal1 s 222 1659 258 2000 4 vdd
rlabel metal1 s 222 2449 258 2790 4 vdd
rlabel metal1 s 222 17459 258 17800 4 vdd
rlabel metal1 s 222 5609 258 5950 4 vdd
rlabel metal1 s 222 5110 258 5451 4 vdd
rlabel metal1 s 222 13800 258 14141 4 vdd
<< properties >>
string FIXED_BBOX 0 0 624 52140
<< end >>
