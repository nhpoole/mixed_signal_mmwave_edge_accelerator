magic
tech sky130A
timestamp 1626486988
<< checkpaint >>
rect -677 -654 677 654
<< metal3 >>
rect -47 16 47 24
rect -47 -16 -36 16
rect -4 -16 4 16
rect 36 -16 47 16
rect -47 -24 47 -16
<< via3 >>
rect -36 -16 -4 16
rect 4 -16 36 16
<< metal4 >>
rect -47 16 47 24
rect -47 -16 -36 16
rect -4 -16 4 16
rect 36 -16 47 16
rect -47 -24 47 -16
<< end >>
