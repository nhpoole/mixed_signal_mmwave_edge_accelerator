magic
tech sky130A
magscale 1 2
timestamp 1624180728
<< nwell >>
rect 342 -10384 24858 4358
<< pwell >>
rect -12358 -27258 24958 -11142
<< nmos >>
rect 2628 -12636 3588 -12036
rect 3646 -12636 4606 -12036
rect 4664 -12636 5624 -12036
rect 5682 -12636 6642 -12036
rect 6700 -12636 7660 -12036
rect 7718 -12636 8678 -12036
rect 8736 -12636 9696 -12036
rect 9754 -12636 10714 -12036
rect 10772 -12636 11732 -12036
rect 11790 -12636 12750 -12036
rect 12808 -12636 13768 -12036
rect 13826 -12636 14786 -12036
rect 14844 -12636 15804 -12036
rect 15862 -12636 16822 -12036
rect 16880 -12636 17840 -12036
rect 17898 -12636 18858 -12036
rect 18916 -12636 19876 -12036
rect 19934 -12636 20894 -12036
rect 20952 -12636 21912 -12036
rect 21970 -12636 22930 -12036
rect 2628 -13454 3588 -12854
rect 3646 -13454 4606 -12854
rect 4664 -13454 5624 -12854
rect 5682 -13454 6642 -12854
rect 6700 -13454 7660 -12854
rect 7718 -13454 8678 -12854
rect 8736 -13454 9696 -12854
rect 9754 -13454 10714 -12854
rect 10772 -13454 11732 -12854
rect 11790 -13454 12750 -12854
rect 12808 -13454 13768 -12854
rect 13826 -13454 14786 -12854
rect 14844 -13454 15804 -12854
rect 15862 -13454 16822 -12854
rect 16880 -13454 17840 -12854
rect 17898 -13454 18858 -12854
rect 18916 -13454 19876 -12854
rect 19934 -13454 20894 -12854
rect 20952 -13454 21912 -12854
rect 21970 -13454 22930 -12854
rect 2628 -14832 3588 -14232
rect 3646 -14832 4606 -14232
rect 4664 -14832 5624 -14232
rect 5682 -14832 6642 -14232
rect 6700 -14832 7660 -14232
rect 7718 -14832 8678 -14232
rect 8736 -14832 9696 -14232
rect 9754 -14832 10714 -14232
rect 10772 -14832 11732 -14232
rect 11790 -14832 12750 -14232
rect 12808 -14832 13768 -14232
rect 13826 -14832 14786 -14232
rect 14844 -14832 15804 -14232
rect 15862 -14832 16822 -14232
rect 16880 -14832 17840 -14232
rect 17898 -14832 18858 -14232
rect 18916 -14832 19876 -14232
rect 19934 -14832 20894 -14232
rect 20952 -14832 21912 -14232
rect 21970 -14832 22930 -14232
rect 2628 -16064 3588 -15464
rect 3646 -16064 4606 -15464
rect 4664 -16064 5624 -15464
rect 5682 -16064 6642 -15464
rect 6700 -16064 7660 -15464
rect 7718 -16064 8678 -15464
rect 8736 -16064 9696 -15464
rect 9754 -16064 10714 -15464
rect 10772 -16064 11732 -15464
rect 11790 -16064 12750 -15464
rect 12808 -16064 13768 -15464
rect 13826 -16064 14786 -15464
rect 14844 -16064 15804 -15464
rect 15862 -16064 16822 -15464
rect 16880 -16064 17840 -15464
rect 17898 -16064 18858 -15464
rect 18916 -16064 19876 -15464
rect 19934 -16064 20894 -15464
rect 20952 -16064 21912 -15464
rect 21970 -16064 22930 -15464
rect 2626 -17298 3586 -16698
rect 3644 -17298 4604 -16698
rect 4662 -17298 5622 -16698
rect 5680 -17298 6640 -16698
rect 6698 -17298 7658 -16698
rect 7716 -17298 8676 -16698
rect 8734 -17298 9694 -16698
rect 9752 -17298 10712 -16698
rect 10770 -17298 11730 -16698
rect 11788 -17298 12748 -16698
rect 12806 -17298 13766 -16698
rect 13824 -17298 14784 -16698
rect 14842 -17298 15802 -16698
rect 15860 -17298 16820 -16698
rect 16878 -17298 17838 -16698
rect 17896 -17298 18856 -16698
rect 18914 -17298 19874 -16698
rect 19932 -17298 20892 -16698
rect 20950 -17298 21910 -16698
rect 21968 -17298 22928 -16698
rect 2626 -18532 3586 -17932
rect 3644 -18532 4604 -17932
rect 4662 -18532 5622 -17932
rect 5680 -18532 6640 -17932
rect 6698 -18532 7658 -17932
rect 7716 -18532 8676 -17932
rect 8734 -18532 9694 -17932
rect 9752 -18532 10712 -17932
rect 10770 -18532 11730 -17932
rect 11788 -18532 12748 -17932
rect 12806 -18532 13766 -17932
rect 13824 -18532 14784 -17932
rect 14842 -18532 15802 -17932
rect 15860 -18532 16820 -17932
rect 16878 -18532 17838 -17932
rect 17896 -18532 18856 -17932
rect 18914 -18532 19874 -17932
rect 19932 -18532 20892 -17932
rect 20950 -18532 21910 -17932
rect 21968 -18532 22928 -17932
rect 2626 -19764 3586 -19164
rect 3644 -19764 4604 -19164
rect 4662 -19764 5622 -19164
rect 5680 -19764 6640 -19164
rect 6698 -19764 7658 -19164
rect 7716 -19764 8676 -19164
rect 8734 -19764 9694 -19164
rect 9752 -19764 10712 -19164
rect 10770 -19764 11730 -19164
rect 11788 -19764 12748 -19164
rect 12806 -19764 13766 -19164
rect 13824 -19764 14784 -19164
rect 14842 -19764 15802 -19164
rect 15860 -19764 16820 -19164
rect 16878 -19764 17838 -19164
rect 17896 -19764 18856 -19164
rect 18914 -19764 19874 -19164
rect 19932 -19764 20892 -19164
rect 20950 -19764 21910 -19164
rect 21968 -19764 22928 -19164
rect 2626 -20998 3586 -20398
rect 3644 -20998 4604 -20398
rect 4662 -20998 5622 -20398
rect 5680 -20998 6640 -20398
rect 6698 -20998 7658 -20398
rect 7716 -20998 8676 -20398
rect 8734 -20998 9694 -20398
rect 9752 -20998 10712 -20398
rect 10770 -20998 11730 -20398
rect 11788 -20998 12748 -20398
rect 12806 -20998 13766 -20398
rect 13824 -20998 14784 -20398
rect 14842 -20998 15802 -20398
rect 15860 -20998 16820 -20398
rect 16878 -20998 17838 -20398
rect 17896 -20998 18856 -20398
rect 18914 -20998 19874 -20398
rect 19932 -20998 20892 -20398
rect 20950 -20998 21910 -20398
rect 21968 -20998 22928 -20398
rect 2626 -22232 3586 -21632
rect 3644 -22232 4604 -21632
rect 4662 -22232 5622 -21632
rect 5680 -22232 6640 -21632
rect 6698 -22232 7658 -21632
rect 7716 -22232 8676 -21632
rect 8734 -22232 9694 -21632
rect 9752 -22232 10712 -21632
rect 10770 -22232 11730 -21632
rect 11788 -22232 12748 -21632
rect 12806 -22232 13766 -21632
rect 13824 -22232 14784 -21632
rect 14842 -22232 15802 -21632
rect 15860 -22232 16820 -21632
rect 16878 -22232 17838 -21632
rect 17896 -22232 18856 -21632
rect 18914 -22232 19874 -21632
rect 19932 -22232 20892 -21632
rect 20950 -22232 21910 -21632
rect 21968 -22232 22928 -21632
rect 2626 -23464 3586 -22864
rect 3644 -23464 4604 -22864
rect 4662 -23464 5622 -22864
rect 5680 -23464 6640 -22864
rect 6698 -23464 7658 -22864
rect 7716 -23464 8676 -22864
rect 8734 -23464 9694 -22864
rect 9752 -23464 10712 -22864
rect 10770 -23464 11730 -22864
rect 11788 -23464 12748 -22864
rect 12806 -23464 13766 -22864
rect 13824 -23464 14784 -22864
rect 14842 -23464 15802 -22864
rect 15860 -23464 16820 -22864
rect 16878 -23464 17838 -22864
rect 17896 -23464 18856 -22864
rect 18914 -23464 19874 -22864
rect 19932 -23464 20892 -22864
rect 20950 -23464 21910 -22864
rect 21968 -23464 22928 -22864
rect 2626 -24698 3586 -24098
rect 3644 -24698 4604 -24098
rect 4662 -24698 5622 -24098
rect 5680 -24698 6640 -24098
rect 6698 -24698 7658 -24098
rect 7716 -24698 8676 -24098
rect 8734 -24698 9694 -24098
rect 9752 -24698 10712 -24098
rect 10770 -24698 11730 -24098
rect 11788 -24698 12748 -24098
rect 12806 -24698 13766 -24098
rect 13824 -24698 14784 -24098
rect 14842 -24698 15802 -24098
rect 15860 -24698 16820 -24098
rect 16878 -24698 17838 -24098
rect 17896 -24698 18856 -24098
rect 18914 -24698 19874 -24098
rect 19932 -24698 20892 -24098
rect 20950 -24698 21910 -24098
rect 21968 -24698 22928 -24098
rect -10004 -25740 -9044 -25140
rect -8986 -25740 -8026 -25140
rect -7968 -25740 -7008 -25140
rect -6950 -25740 -5990 -25140
rect -5932 -25740 -4972 -25140
rect -4914 -25740 -3954 -25140
rect -3896 -25740 -2936 -25140
rect -2878 -25740 -1918 -25140
rect -1860 -25740 -900 -25140
rect -842 -25740 118 -25140
rect 2626 -25930 3586 -25330
rect 3644 -25930 4604 -25330
rect 4662 -25930 5622 -25330
rect 5680 -25930 6640 -25330
rect 6698 -25930 7658 -25330
rect 7716 -25930 8676 -25330
rect 8734 -25930 9694 -25330
rect 9752 -25930 10712 -25330
rect 10770 -25930 11730 -25330
rect 11788 -25930 12748 -25330
rect 12806 -25930 13766 -25330
rect 13824 -25930 14784 -25330
rect 14842 -25930 15802 -25330
rect 15860 -25930 16820 -25330
rect 16878 -25930 17838 -25330
rect 17896 -25930 18856 -25330
rect 18914 -25930 19874 -25330
rect 19932 -25930 20892 -25330
rect 20950 -25930 21910 -25330
rect 21968 -25930 22928 -25330
<< pmos >>
rect 7520 -5672 8480 -5072
rect 8538 -5672 9498 -5072
rect 9556 -5672 10516 -5072
rect 10574 -5672 11534 -5072
rect 11592 -5672 12552 -5072
rect 12610 -5672 13570 -5072
rect 13628 -5672 14588 -5072
rect 14646 -5672 15606 -5072
rect 15664 -5672 16624 -5072
rect 16682 -5672 17642 -5072
rect 17700 -5672 18660 -5072
rect 18718 -5672 19678 -5072
rect 19736 -5672 20696 -5072
rect 20754 -5672 21714 -5072
rect 21772 -5672 22732 -5072
rect 7520 -6928 8480 -6328
rect 8538 -6928 9498 -6328
rect 9556 -6928 10516 -6328
rect 10574 -6928 11534 -6328
rect 11592 -6928 12552 -6328
rect 12610 -6928 13570 -6328
rect 13628 -6928 14588 -6328
rect 14646 -6928 15606 -6328
rect 15664 -6928 16624 -6328
rect 16682 -6928 17642 -6328
rect 17700 -6928 18660 -6328
rect 18718 -6928 19678 -6328
rect 19736 -6928 20696 -6328
rect 20754 -6928 21714 -6328
rect 21772 -6928 22732 -6328
rect 7520 -8184 8480 -7584
rect 8538 -8184 9498 -7584
rect 9556 -8184 10516 -7584
rect 10574 -8184 11534 -7584
rect 11592 -8184 12552 -7584
rect 12610 -8184 13570 -7584
rect 13628 -8184 14588 -7584
rect 14646 -8184 15606 -7584
rect 15664 -8184 16624 -7584
rect 16682 -8184 17642 -7584
rect 17700 -8184 18660 -7584
rect 18718 -8184 19678 -7584
rect 19736 -8184 20696 -7584
rect 20754 -8184 21714 -7584
rect 21772 -8184 22732 -7584
rect 7520 -9440 8480 -8840
rect 8538 -9440 9498 -8840
rect 9556 -9440 10516 -8840
rect 10574 -9440 11534 -8840
rect 11592 -9440 12552 -8840
rect 12610 -9440 13570 -8840
rect 13628 -9440 14588 -8840
rect 14646 -9440 15606 -8840
rect 15664 -9440 16624 -8840
rect 16682 -9440 17642 -8840
rect 17700 -9440 18660 -8840
rect 18718 -9440 19678 -8840
rect 19736 -9440 20696 -8840
rect 20754 -9440 21714 -8840
rect 21772 -9440 22732 -8840
<< pmoslvt >>
rect 6534 874 7494 1474
rect 7552 874 8512 1474
rect 8570 874 9530 1474
rect 9588 874 10548 1474
rect 10606 874 11566 1474
rect 11624 874 12584 1474
rect 12642 874 13602 1474
rect 13660 874 14620 1474
rect 14678 874 15638 1474
rect 15696 874 16656 1474
rect 16714 874 17674 1474
rect 17732 874 18692 1474
rect 18750 874 19710 1474
rect 19768 874 20728 1474
rect 20786 874 21746 1474
rect 21804 874 22764 1474
rect 6534 -262 7494 338
rect 7552 -262 8512 338
rect 8570 -262 9530 338
rect 9588 -262 10548 338
rect 10606 -262 11566 338
rect 11624 -262 12584 338
rect 12642 -262 13602 338
rect 13660 -262 14620 338
rect 14678 -262 15638 338
rect 15696 -262 16656 338
rect 16714 -262 17674 338
rect 17732 -262 18692 338
rect 18750 -262 19710 338
rect 19768 -262 20728 338
rect 20786 -262 21746 338
rect 21804 -262 22764 338
rect 6534 -1398 7494 -798
rect 7552 -1398 8512 -798
rect 8570 -1398 9530 -798
rect 9588 -1398 10548 -798
rect 10606 -1398 11566 -798
rect 11624 -1398 12584 -798
rect 12642 -1398 13602 -798
rect 13660 -1398 14620 -798
rect 14678 -1398 15638 -798
rect 15696 -1398 16656 -798
rect 16714 -1398 17674 -798
rect 17732 -1398 18692 -798
rect 18750 -1398 19710 -798
rect 19768 -1398 20728 -798
rect 20786 -1398 21746 -798
rect 21804 -1398 22764 -798
rect 7728 -3036 8688 -2436
rect 8746 -3036 9706 -2436
rect 9764 -3036 10724 -2436
rect 10782 -3036 11742 -2436
rect 11800 -3036 12760 -2436
rect 12818 -3036 13778 -2436
rect 13836 -3036 14796 -2436
rect 14854 -3036 15814 -2436
rect 15872 -3036 16832 -2436
rect 16890 -3036 17850 -2436
rect 17908 -3036 18868 -2436
rect 18926 -3036 19886 -2436
rect 19944 -3036 20904 -2436
rect 20962 -3036 21922 -2436
rect 7728 -4068 8688 -3468
rect 8746 -4068 9706 -3468
rect 9764 -4068 10724 -3468
rect 10782 -4068 11742 -3468
rect 11800 -4068 12760 -3468
rect 12818 -4068 13778 -3468
rect 13836 -4068 14796 -3468
rect 14854 -4068 15814 -3468
rect 15872 -4068 16832 -3468
rect 16890 -4068 17850 -3468
rect 17908 -4068 18868 -3468
rect 18926 -4068 19886 -3468
rect 19944 -4068 20904 -3468
rect 20962 -4068 21922 -3468
rect 2216 -5776 3176 -5176
rect 3234 -5776 4194 -5176
rect 4252 -5776 5212 -5176
rect 5270 -5776 6230 -5176
rect 2216 -6808 3176 -6208
rect 3234 -6808 4194 -6208
rect 4252 -6808 5212 -6208
rect 5270 -6808 6230 -6208
rect 2216 -7840 3176 -7240
rect 3234 -7840 4194 -7240
rect 4252 -7840 5212 -7240
rect 5270 -7840 6230 -7240
rect 2216 -8872 3176 -8272
rect 3234 -8872 4194 -8272
rect 4252 -8872 5212 -8272
rect 5270 -8872 6230 -8272
<< nmoslvt >>
rect -9138 -13112 -8178 -12512
rect -8120 -13112 -7160 -12512
rect -7102 -13112 -6142 -12512
rect -6084 -13112 -5124 -12512
rect -5066 -13112 -4106 -12512
rect -4048 -13112 -3088 -12512
rect -3030 -13112 -2070 -12512
rect -2012 -13112 -1052 -12512
rect -994 -13112 -34 -12512
rect -9138 -13930 -8178 -13330
rect -8120 -13930 -7160 -13330
rect -7102 -13930 -6142 -13330
rect -6084 -13930 -5124 -13330
rect -5066 -13930 -4106 -13330
rect -4048 -13930 -3088 -13330
rect -3030 -13930 -2070 -13330
rect -2012 -13930 -1052 -13330
rect -994 -13930 -34 -13330
rect -9138 -14748 -8178 -14148
rect -8120 -14748 -7160 -14148
rect -7102 -14748 -6142 -14148
rect -6084 -14748 -5124 -14148
rect -5066 -14748 -4106 -14148
rect -4048 -14748 -3088 -14148
rect -3030 -14748 -2070 -14148
rect -2012 -14748 -1052 -14148
rect -994 -14748 -34 -14148
rect -9138 -15566 -8178 -14966
rect -8120 -15566 -7160 -14966
rect -7102 -15566 -6142 -14966
rect -6084 -15566 -5124 -14966
rect -5066 -15566 -4106 -14966
rect -4048 -15566 -3088 -14966
rect -3030 -15566 -2070 -14966
rect -2012 -15566 -1052 -14966
rect -994 -15566 -34 -14966
rect -9138 -16384 -8178 -15784
rect -8120 -16384 -7160 -15784
rect -7102 -16384 -6142 -15784
rect -6084 -16384 -5124 -15784
rect -5066 -16384 -4106 -15784
rect -4048 -16384 -3088 -15784
rect -3030 -16384 -2070 -15784
rect -2012 -16384 -1052 -15784
rect -994 -16384 -34 -15784
rect -9138 -17202 -8178 -16602
rect -8120 -17202 -7160 -16602
rect -7102 -17202 -6142 -16602
rect -6084 -17202 -5124 -16602
rect -5066 -17202 -4106 -16602
rect -4048 -17202 -3088 -16602
rect -3030 -17202 -2070 -16602
rect -2012 -17202 -1052 -16602
rect -994 -17202 -34 -16602
rect -9138 -18020 -8178 -17420
rect -8120 -18020 -7160 -17420
rect -7102 -18020 -6142 -17420
rect -6084 -18020 -5124 -17420
rect -5066 -18020 -4106 -17420
rect -4048 -18020 -3088 -17420
rect -3030 -18020 -2070 -17420
rect -2012 -18020 -1052 -17420
rect -994 -18020 -34 -17420
rect -9138 -18838 -8178 -18238
rect -8120 -18838 -7160 -18238
rect -7102 -18838 -6142 -18238
rect -6084 -18838 -5124 -18238
rect -5066 -18838 -4106 -18238
rect -4048 -18838 -3088 -18238
rect -3030 -18838 -2070 -18238
rect -2012 -18838 -1052 -18238
rect -994 -18838 -34 -18238
rect -10462 -20862 -9502 -20262
rect -9444 -20862 -8484 -20262
rect -8426 -20862 -7466 -20262
rect -7408 -20862 -6448 -20262
rect -6390 -20862 -5430 -20262
rect -5372 -20862 -4412 -20262
rect -4354 -20862 -3394 -20262
rect -3336 -20862 -2376 -20262
rect -2318 -20862 -1358 -20262
rect -1300 -20862 -340 -20262
rect -282 -20862 678 -20262
rect -10462 -21974 -9502 -21374
rect -9444 -21974 -8484 -21374
rect -8426 -21974 -7466 -21374
rect -7408 -21974 -6448 -21374
rect -6390 -21974 -5430 -21374
rect -5372 -21974 -4412 -21374
rect -4354 -21974 -3394 -21374
rect -3336 -21974 -2376 -21374
rect -2318 -21974 -1358 -21374
rect -1300 -21974 -340 -21374
rect -282 -21974 678 -21374
rect -10462 -23086 -9502 -22486
rect -9444 -23086 -8484 -22486
rect -8426 -23086 -7466 -22486
rect -7408 -23086 -6448 -22486
rect -6390 -23086 -5430 -22486
rect -5372 -23086 -4412 -22486
rect -4354 -23086 -3394 -22486
rect -3336 -23086 -2376 -22486
rect -2318 -23086 -1358 -22486
rect -1300 -23086 -340 -22486
rect -282 -23086 678 -22486
rect -10462 -24198 -9502 -23598
rect -9444 -24198 -8484 -23598
rect -8426 -24198 -7466 -23598
rect -7408 -24198 -6448 -23598
rect -6390 -24198 -5430 -23598
rect -5372 -24198 -4412 -23598
rect -4354 -24198 -3394 -23598
rect -3336 -24198 -2376 -23598
rect -2318 -24198 -1358 -23598
rect -1300 -24198 -340 -23598
rect -282 -24198 678 -23598
<< ndiff >>
rect 2570 -12048 2628 -12036
rect -9196 -12524 -9138 -12512
rect -9196 -13100 -9184 -12524
rect -9150 -13100 -9138 -12524
rect -9196 -13112 -9138 -13100
rect -8178 -12524 -8120 -12512
rect -8178 -13100 -8166 -12524
rect -8132 -13100 -8120 -12524
rect -8178 -13112 -8120 -13100
rect -7160 -12524 -7102 -12512
rect -7160 -13100 -7148 -12524
rect -7114 -13100 -7102 -12524
rect -7160 -13112 -7102 -13100
rect -6142 -12524 -6084 -12512
rect -6142 -13100 -6130 -12524
rect -6096 -13100 -6084 -12524
rect -6142 -13112 -6084 -13100
rect -5124 -12524 -5066 -12512
rect -5124 -13100 -5112 -12524
rect -5078 -13100 -5066 -12524
rect -5124 -13112 -5066 -13100
rect -4106 -12524 -4048 -12512
rect -4106 -13100 -4094 -12524
rect -4060 -13100 -4048 -12524
rect -4106 -13112 -4048 -13100
rect -3088 -12524 -3030 -12512
rect -3088 -13100 -3076 -12524
rect -3042 -13100 -3030 -12524
rect -3088 -13112 -3030 -13100
rect -2070 -12524 -2012 -12512
rect -2070 -13100 -2058 -12524
rect -2024 -13100 -2012 -12524
rect -2070 -13112 -2012 -13100
rect -1052 -12524 -994 -12512
rect -1052 -13100 -1040 -12524
rect -1006 -13100 -994 -12524
rect -1052 -13112 -994 -13100
rect -34 -12524 24 -12512
rect -34 -13100 -22 -12524
rect 12 -13100 24 -12524
rect 2570 -12624 2582 -12048
rect 2616 -12624 2628 -12048
rect 2570 -12636 2628 -12624
rect 3588 -12048 3646 -12036
rect 3588 -12624 3600 -12048
rect 3634 -12624 3646 -12048
rect 3588 -12636 3646 -12624
rect 4606 -12048 4664 -12036
rect 4606 -12624 4618 -12048
rect 4652 -12624 4664 -12048
rect 4606 -12636 4664 -12624
rect 5624 -12048 5682 -12036
rect 5624 -12624 5636 -12048
rect 5670 -12624 5682 -12048
rect 5624 -12636 5682 -12624
rect 6642 -12048 6700 -12036
rect 6642 -12624 6654 -12048
rect 6688 -12624 6700 -12048
rect 6642 -12636 6700 -12624
rect 7660 -12048 7718 -12036
rect 7660 -12624 7672 -12048
rect 7706 -12624 7718 -12048
rect 7660 -12636 7718 -12624
rect 8678 -12048 8736 -12036
rect 8678 -12624 8690 -12048
rect 8724 -12624 8736 -12048
rect 8678 -12636 8736 -12624
rect 9696 -12048 9754 -12036
rect 9696 -12624 9708 -12048
rect 9742 -12624 9754 -12048
rect 9696 -12636 9754 -12624
rect 10714 -12048 10772 -12036
rect 10714 -12624 10726 -12048
rect 10760 -12624 10772 -12048
rect 10714 -12636 10772 -12624
rect 11732 -12048 11790 -12036
rect 11732 -12624 11744 -12048
rect 11778 -12624 11790 -12048
rect 11732 -12636 11790 -12624
rect 12750 -12048 12808 -12036
rect 12750 -12624 12762 -12048
rect 12796 -12624 12808 -12048
rect 12750 -12636 12808 -12624
rect 13768 -12048 13826 -12036
rect 13768 -12624 13780 -12048
rect 13814 -12624 13826 -12048
rect 13768 -12636 13826 -12624
rect 14786 -12048 14844 -12036
rect 14786 -12624 14798 -12048
rect 14832 -12624 14844 -12048
rect 14786 -12636 14844 -12624
rect 15804 -12048 15862 -12036
rect 15804 -12624 15816 -12048
rect 15850 -12624 15862 -12048
rect 15804 -12636 15862 -12624
rect 16822 -12048 16880 -12036
rect 16822 -12624 16834 -12048
rect 16868 -12624 16880 -12048
rect 16822 -12636 16880 -12624
rect 17840 -12048 17898 -12036
rect 17840 -12624 17852 -12048
rect 17886 -12624 17898 -12048
rect 17840 -12636 17898 -12624
rect 18858 -12048 18916 -12036
rect 18858 -12624 18870 -12048
rect 18904 -12624 18916 -12048
rect 18858 -12636 18916 -12624
rect 19876 -12048 19934 -12036
rect 19876 -12624 19888 -12048
rect 19922 -12624 19934 -12048
rect 19876 -12636 19934 -12624
rect 20894 -12048 20952 -12036
rect 20894 -12624 20906 -12048
rect 20940 -12624 20952 -12048
rect 20894 -12636 20952 -12624
rect 21912 -12048 21970 -12036
rect 21912 -12624 21924 -12048
rect 21958 -12624 21970 -12048
rect 21912 -12636 21970 -12624
rect 22930 -12048 22988 -12036
rect 22930 -12624 22942 -12048
rect 22976 -12624 22988 -12048
rect 22930 -12636 22988 -12624
rect -34 -13112 24 -13100
rect 2570 -12866 2628 -12854
rect -9196 -13342 -9138 -13330
rect -9196 -13918 -9184 -13342
rect -9150 -13918 -9138 -13342
rect -9196 -13930 -9138 -13918
rect -8178 -13342 -8120 -13330
rect -8178 -13918 -8166 -13342
rect -8132 -13918 -8120 -13342
rect -8178 -13930 -8120 -13918
rect -7160 -13342 -7102 -13330
rect -7160 -13918 -7148 -13342
rect -7114 -13918 -7102 -13342
rect -7160 -13930 -7102 -13918
rect -6142 -13342 -6084 -13330
rect -6142 -13918 -6130 -13342
rect -6096 -13918 -6084 -13342
rect -6142 -13930 -6084 -13918
rect -5124 -13342 -5066 -13330
rect -5124 -13918 -5112 -13342
rect -5078 -13918 -5066 -13342
rect -5124 -13930 -5066 -13918
rect -4106 -13342 -4048 -13330
rect -4106 -13918 -4094 -13342
rect -4060 -13918 -4048 -13342
rect -4106 -13930 -4048 -13918
rect -3088 -13342 -3030 -13330
rect -3088 -13918 -3076 -13342
rect -3042 -13918 -3030 -13342
rect -3088 -13930 -3030 -13918
rect -2070 -13342 -2012 -13330
rect -2070 -13918 -2058 -13342
rect -2024 -13918 -2012 -13342
rect -2070 -13930 -2012 -13918
rect -1052 -13342 -994 -13330
rect -1052 -13918 -1040 -13342
rect -1006 -13918 -994 -13342
rect -1052 -13930 -994 -13918
rect -34 -13342 24 -13330
rect -34 -13918 -22 -13342
rect 12 -13918 24 -13342
rect 2570 -13442 2582 -12866
rect 2616 -13442 2628 -12866
rect 2570 -13454 2628 -13442
rect 3588 -12866 3646 -12854
rect 3588 -13442 3600 -12866
rect 3634 -13442 3646 -12866
rect 3588 -13454 3646 -13442
rect 4606 -12866 4664 -12854
rect 4606 -13442 4618 -12866
rect 4652 -13442 4664 -12866
rect 4606 -13454 4664 -13442
rect 5624 -12866 5682 -12854
rect 5624 -13442 5636 -12866
rect 5670 -13442 5682 -12866
rect 5624 -13454 5682 -13442
rect 6642 -12866 6700 -12854
rect 6642 -13442 6654 -12866
rect 6688 -13442 6700 -12866
rect 6642 -13454 6700 -13442
rect 7660 -12866 7718 -12854
rect 7660 -13442 7672 -12866
rect 7706 -13442 7718 -12866
rect 7660 -13454 7718 -13442
rect 8678 -12866 8736 -12854
rect 8678 -13442 8690 -12866
rect 8724 -13442 8736 -12866
rect 8678 -13454 8736 -13442
rect 9696 -12866 9754 -12854
rect 9696 -13442 9708 -12866
rect 9742 -13442 9754 -12866
rect 9696 -13454 9754 -13442
rect 10714 -12866 10772 -12854
rect 10714 -13442 10726 -12866
rect 10760 -13442 10772 -12866
rect 10714 -13454 10772 -13442
rect 11732 -12866 11790 -12854
rect 11732 -13442 11744 -12866
rect 11778 -13442 11790 -12866
rect 11732 -13454 11790 -13442
rect 12750 -12866 12808 -12854
rect 12750 -13442 12762 -12866
rect 12796 -13442 12808 -12866
rect 12750 -13454 12808 -13442
rect 13768 -12866 13826 -12854
rect 13768 -13442 13780 -12866
rect 13814 -13442 13826 -12866
rect 13768 -13454 13826 -13442
rect 14786 -12866 14844 -12854
rect 14786 -13442 14798 -12866
rect 14832 -13442 14844 -12866
rect 14786 -13454 14844 -13442
rect 15804 -12866 15862 -12854
rect 15804 -13442 15816 -12866
rect 15850 -13442 15862 -12866
rect 15804 -13454 15862 -13442
rect 16822 -12866 16880 -12854
rect 16822 -13442 16834 -12866
rect 16868 -13442 16880 -12866
rect 16822 -13454 16880 -13442
rect 17840 -12866 17898 -12854
rect 17840 -13442 17852 -12866
rect 17886 -13442 17898 -12866
rect 17840 -13454 17898 -13442
rect 18858 -12866 18916 -12854
rect 18858 -13442 18870 -12866
rect 18904 -13442 18916 -12866
rect 18858 -13454 18916 -13442
rect 19876 -12866 19934 -12854
rect 19876 -13442 19888 -12866
rect 19922 -13442 19934 -12866
rect 19876 -13454 19934 -13442
rect 20894 -12866 20952 -12854
rect 20894 -13442 20906 -12866
rect 20940 -13442 20952 -12866
rect 20894 -13454 20952 -13442
rect 21912 -12866 21970 -12854
rect 21912 -13442 21924 -12866
rect 21958 -13442 21970 -12866
rect 21912 -13454 21970 -13442
rect 22930 -12866 22988 -12854
rect 22930 -13442 22942 -12866
rect 22976 -13442 22988 -12866
rect 22930 -13454 22988 -13442
rect -34 -13930 24 -13918
rect -9196 -14160 -9138 -14148
rect -9196 -14736 -9184 -14160
rect -9150 -14736 -9138 -14160
rect -9196 -14748 -9138 -14736
rect -8178 -14160 -8120 -14148
rect -8178 -14736 -8166 -14160
rect -8132 -14736 -8120 -14160
rect -8178 -14748 -8120 -14736
rect -7160 -14160 -7102 -14148
rect -7160 -14736 -7148 -14160
rect -7114 -14736 -7102 -14160
rect -7160 -14748 -7102 -14736
rect -6142 -14160 -6084 -14148
rect -6142 -14736 -6130 -14160
rect -6096 -14736 -6084 -14160
rect -6142 -14748 -6084 -14736
rect -5124 -14160 -5066 -14148
rect -5124 -14736 -5112 -14160
rect -5078 -14736 -5066 -14160
rect -5124 -14748 -5066 -14736
rect -4106 -14160 -4048 -14148
rect -4106 -14736 -4094 -14160
rect -4060 -14736 -4048 -14160
rect -4106 -14748 -4048 -14736
rect -3088 -14160 -3030 -14148
rect -3088 -14736 -3076 -14160
rect -3042 -14736 -3030 -14160
rect -3088 -14748 -3030 -14736
rect -2070 -14160 -2012 -14148
rect -2070 -14736 -2058 -14160
rect -2024 -14736 -2012 -14160
rect -2070 -14748 -2012 -14736
rect -1052 -14160 -994 -14148
rect -1052 -14736 -1040 -14160
rect -1006 -14736 -994 -14160
rect -1052 -14748 -994 -14736
rect -34 -14160 24 -14148
rect -34 -14736 -22 -14160
rect 12 -14736 24 -14160
rect -34 -14748 24 -14736
rect 2570 -14244 2628 -14232
rect 2570 -14820 2582 -14244
rect 2616 -14820 2628 -14244
rect 2570 -14832 2628 -14820
rect 3588 -14244 3646 -14232
rect 3588 -14820 3600 -14244
rect 3634 -14820 3646 -14244
rect 3588 -14832 3646 -14820
rect 4606 -14244 4664 -14232
rect 4606 -14820 4618 -14244
rect 4652 -14820 4664 -14244
rect 4606 -14832 4664 -14820
rect 5624 -14244 5682 -14232
rect 5624 -14820 5636 -14244
rect 5670 -14820 5682 -14244
rect 5624 -14832 5682 -14820
rect 6642 -14244 6700 -14232
rect 6642 -14820 6654 -14244
rect 6688 -14820 6700 -14244
rect 6642 -14832 6700 -14820
rect 7660 -14244 7718 -14232
rect 7660 -14820 7672 -14244
rect 7706 -14820 7718 -14244
rect 7660 -14832 7718 -14820
rect 8678 -14244 8736 -14232
rect 8678 -14820 8690 -14244
rect 8724 -14820 8736 -14244
rect 8678 -14832 8736 -14820
rect 9696 -14244 9754 -14232
rect 9696 -14820 9708 -14244
rect 9742 -14820 9754 -14244
rect 9696 -14832 9754 -14820
rect 10714 -14244 10772 -14232
rect 10714 -14820 10726 -14244
rect 10760 -14820 10772 -14244
rect 10714 -14832 10772 -14820
rect 11732 -14244 11790 -14232
rect 11732 -14820 11744 -14244
rect 11778 -14820 11790 -14244
rect 11732 -14832 11790 -14820
rect 12750 -14244 12808 -14232
rect 12750 -14820 12762 -14244
rect 12796 -14820 12808 -14244
rect 12750 -14832 12808 -14820
rect 13768 -14244 13826 -14232
rect 13768 -14820 13780 -14244
rect 13814 -14820 13826 -14244
rect 13768 -14832 13826 -14820
rect 14786 -14244 14844 -14232
rect 14786 -14820 14798 -14244
rect 14832 -14820 14844 -14244
rect 14786 -14832 14844 -14820
rect 15804 -14244 15862 -14232
rect 15804 -14820 15816 -14244
rect 15850 -14820 15862 -14244
rect 15804 -14832 15862 -14820
rect 16822 -14244 16880 -14232
rect 16822 -14820 16834 -14244
rect 16868 -14820 16880 -14244
rect 16822 -14832 16880 -14820
rect 17840 -14244 17898 -14232
rect 17840 -14820 17852 -14244
rect 17886 -14820 17898 -14244
rect 17840 -14832 17898 -14820
rect 18858 -14244 18916 -14232
rect 18858 -14820 18870 -14244
rect 18904 -14820 18916 -14244
rect 18858 -14832 18916 -14820
rect 19876 -14244 19934 -14232
rect 19876 -14820 19888 -14244
rect 19922 -14820 19934 -14244
rect 19876 -14832 19934 -14820
rect 20894 -14244 20952 -14232
rect 20894 -14820 20906 -14244
rect 20940 -14820 20952 -14244
rect 20894 -14832 20952 -14820
rect 21912 -14244 21970 -14232
rect 21912 -14820 21924 -14244
rect 21958 -14820 21970 -14244
rect 21912 -14832 21970 -14820
rect 22930 -14244 22988 -14232
rect 22930 -14820 22942 -14244
rect 22976 -14820 22988 -14244
rect 22930 -14832 22988 -14820
rect -9196 -14978 -9138 -14966
rect -9196 -15554 -9184 -14978
rect -9150 -15554 -9138 -14978
rect -9196 -15566 -9138 -15554
rect -8178 -14978 -8120 -14966
rect -8178 -15554 -8166 -14978
rect -8132 -15554 -8120 -14978
rect -8178 -15566 -8120 -15554
rect -7160 -14978 -7102 -14966
rect -7160 -15554 -7148 -14978
rect -7114 -15554 -7102 -14978
rect -7160 -15566 -7102 -15554
rect -6142 -14978 -6084 -14966
rect -6142 -15554 -6130 -14978
rect -6096 -15554 -6084 -14978
rect -6142 -15566 -6084 -15554
rect -5124 -14978 -5066 -14966
rect -5124 -15554 -5112 -14978
rect -5078 -15554 -5066 -14978
rect -5124 -15566 -5066 -15554
rect -4106 -14978 -4048 -14966
rect -4106 -15554 -4094 -14978
rect -4060 -15554 -4048 -14978
rect -4106 -15566 -4048 -15554
rect -3088 -14978 -3030 -14966
rect -3088 -15554 -3076 -14978
rect -3042 -15554 -3030 -14978
rect -3088 -15566 -3030 -15554
rect -2070 -14978 -2012 -14966
rect -2070 -15554 -2058 -14978
rect -2024 -15554 -2012 -14978
rect -2070 -15566 -2012 -15554
rect -1052 -14978 -994 -14966
rect -1052 -15554 -1040 -14978
rect -1006 -15554 -994 -14978
rect -1052 -15566 -994 -15554
rect -34 -14978 24 -14966
rect -34 -15554 -22 -14978
rect 12 -15554 24 -14978
rect -34 -15566 24 -15554
rect 2570 -15476 2628 -15464
rect -9196 -15796 -9138 -15784
rect -9196 -16372 -9184 -15796
rect -9150 -16372 -9138 -15796
rect -9196 -16384 -9138 -16372
rect -8178 -15796 -8120 -15784
rect -8178 -16372 -8166 -15796
rect -8132 -16372 -8120 -15796
rect -8178 -16384 -8120 -16372
rect -7160 -15796 -7102 -15784
rect -7160 -16372 -7148 -15796
rect -7114 -16372 -7102 -15796
rect -7160 -16384 -7102 -16372
rect -6142 -15796 -6084 -15784
rect -6142 -16372 -6130 -15796
rect -6096 -16372 -6084 -15796
rect -6142 -16384 -6084 -16372
rect -5124 -15796 -5066 -15784
rect -5124 -16372 -5112 -15796
rect -5078 -16372 -5066 -15796
rect -5124 -16384 -5066 -16372
rect -4106 -15796 -4048 -15784
rect -4106 -16372 -4094 -15796
rect -4060 -16372 -4048 -15796
rect -4106 -16384 -4048 -16372
rect -3088 -15796 -3030 -15784
rect -3088 -16372 -3076 -15796
rect -3042 -16372 -3030 -15796
rect -3088 -16384 -3030 -16372
rect -2070 -15796 -2012 -15784
rect -2070 -16372 -2058 -15796
rect -2024 -16372 -2012 -15796
rect -2070 -16384 -2012 -16372
rect -1052 -15796 -994 -15784
rect -1052 -16372 -1040 -15796
rect -1006 -16372 -994 -15796
rect -1052 -16384 -994 -16372
rect -34 -15796 24 -15784
rect -34 -16372 -22 -15796
rect 12 -16372 24 -15796
rect 2570 -16052 2582 -15476
rect 2616 -16052 2628 -15476
rect 2570 -16064 2628 -16052
rect 3588 -15476 3646 -15464
rect 3588 -16052 3600 -15476
rect 3634 -16052 3646 -15476
rect 3588 -16064 3646 -16052
rect 4606 -15476 4664 -15464
rect 4606 -16052 4618 -15476
rect 4652 -16052 4664 -15476
rect 4606 -16064 4664 -16052
rect 5624 -15476 5682 -15464
rect 5624 -16052 5636 -15476
rect 5670 -16052 5682 -15476
rect 5624 -16064 5682 -16052
rect 6642 -15476 6700 -15464
rect 6642 -16052 6654 -15476
rect 6688 -16052 6700 -15476
rect 6642 -16064 6700 -16052
rect 7660 -15476 7718 -15464
rect 7660 -16052 7672 -15476
rect 7706 -16052 7718 -15476
rect 7660 -16064 7718 -16052
rect 8678 -15476 8736 -15464
rect 8678 -16052 8690 -15476
rect 8724 -16052 8736 -15476
rect 8678 -16064 8736 -16052
rect 9696 -15476 9754 -15464
rect 9696 -16052 9708 -15476
rect 9742 -16052 9754 -15476
rect 9696 -16064 9754 -16052
rect 10714 -15476 10772 -15464
rect 10714 -16052 10726 -15476
rect 10760 -16052 10772 -15476
rect 10714 -16064 10772 -16052
rect 11732 -15476 11790 -15464
rect 11732 -16052 11744 -15476
rect 11778 -16052 11790 -15476
rect 11732 -16064 11790 -16052
rect 12750 -15476 12808 -15464
rect 12750 -16052 12762 -15476
rect 12796 -16052 12808 -15476
rect 12750 -16064 12808 -16052
rect 13768 -15476 13826 -15464
rect 13768 -16052 13780 -15476
rect 13814 -16052 13826 -15476
rect 13768 -16064 13826 -16052
rect 14786 -15476 14844 -15464
rect 14786 -16052 14798 -15476
rect 14832 -16052 14844 -15476
rect 14786 -16064 14844 -16052
rect 15804 -15476 15862 -15464
rect 15804 -16052 15816 -15476
rect 15850 -16052 15862 -15476
rect 15804 -16064 15862 -16052
rect 16822 -15476 16880 -15464
rect 16822 -16052 16834 -15476
rect 16868 -16052 16880 -15476
rect 16822 -16064 16880 -16052
rect 17840 -15476 17898 -15464
rect 17840 -16052 17852 -15476
rect 17886 -16052 17898 -15476
rect 17840 -16064 17898 -16052
rect 18858 -15476 18916 -15464
rect 18858 -16052 18870 -15476
rect 18904 -16052 18916 -15476
rect 18858 -16064 18916 -16052
rect 19876 -15476 19934 -15464
rect 19876 -16052 19888 -15476
rect 19922 -16052 19934 -15476
rect 19876 -16064 19934 -16052
rect 20894 -15476 20952 -15464
rect 20894 -16052 20906 -15476
rect 20940 -16052 20952 -15476
rect 20894 -16064 20952 -16052
rect 21912 -15476 21970 -15464
rect 21912 -16052 21924 -15476
rect 21958 -16052 21970 -15476
rect 21912 -16064 21970 -16052
rect 22930 -15476 22988 -15464
rect 22930 -16052 22942 -15476
rect 22976 -16052 22988 -15476
rect 22930 -16064 22988 -16052
rect -34 -16384 24 -16372
rect -9196 -16614 -9138 -16602
rect -9196 -17190 -9184 -16614
rect -9150 -17190 -9138 -16614
rect -9196 -17202 -9138 -17190
rect -8178 -16614 -8120 -16602
rect -8178 -17190 -8166 -16614
rect -8132 -17190 -8120 -16614
rect -8178 -17202 -8120 -17190
rect -7160 -16614 -7102 -16602
rect -7160 -17190 -7148 -16614
rect -7114 -17190 -7102 -16614
rect -7160 -17202 -7102 -17190
rect -6142 -16614 -6084 -16602
rect -6142 -17190 -6130 -16614
rect -6096 -17190 -6084 -16614
rect -6142 -17202 -6084 -17190
rect -5124 -16614 -5066 -16602
rect -5124 -17190 -5112 -16614
rect -5078 -17190 -5066 -16614
rect -5124 -17202 -5066 -17190
rect -4106 -16614 -4048 -16602
rect -4106 -17190 -4094 -16614
rect -4060 -17190 -4048 -16614
rect -4106 -17202 -4048 -17190
rect -3088 -16614 -3030 -16602
rect -3088 -17190 -3076 -16614
rect -3042 -17190 -3030 -16614
rect -3088 -17202 -3030 -17190
rect -2070 -16614 -2012 -16602
rect -2070 -17190 -2058 -16614
rect -2024 -17190 -2012 -16614
rect -2070 -17202 -2012 -17190
rect -1052 -16614 -994 -16602
rect -1052 -17190 -1040 -16614
rect -1006 -17190 -994 -16614
rect -1052 -17202 -994 -17190
rect -34 -16614 24 -16602
rect -34 -17190 -22 -16614
rect 12 -17190 24 -16614
rect -34 -17202 24 -17190
rect 2568 -16710 2626 -16698
rect 2568 -17286 2580 -16710
rect 2614 -17286 2626 -16710
rect 2568 -17298 2626 -17286
rect 3586 -16710 3644 -16698
rect 3586 -17286 3598 -16710
rect 3632 -17286 3644 -16710
rect 3586 -17298 3644 -17286
rect 4604 -16710 4662 -16698
rect 4604 -17286 4616 -16710
rect 4650 -17286 4662 -16710
rect 4604 -17298 4662 -17286
rect 5622 -16710 5680 -16698
rect 5622 -17286 5634 -16710
rect 5668 -17286 5680 -16710
rect 5622 -17298 5680 -17286
rect 6640 -16710 6698 -16698
rect 6640 -17286 6652 -16710
rect 6686 -17286 6698 -16710
rect 6640 -17298 6698 -17286
rect 7658 -16710 7716 -16698
rect 7658 -17286 7670 -16710
rect 7704 -17286 7716 -16710
rect 7658 -17298 7716 -17286
rect 8676 -16710 8734 -16698
rect 8676 -17286 8688 -16710
rect 8722 -17286 8734 -16710
rect 8676 -17298 8734 -17286
rect 9694 -16710 9752 -16698
rect 9694 -17286 9706 -16710
rect 9740 -17286 9752 -16710
rect 9694 -17298 9752 -17286
rect 10712 -16710 10770 -16698
rect 10712 -17286 10724 -16710
rect 10758 -17286 10770 -16710
rect 10712 -17298 10770 -17286
rect 11730 -16710 11788 -16698
rect 11730 -17286 11742 -16710
rect 11776 -17286 11788 -16710
rect 11730 -17298 11788 -17286
rect 12748 -16710 12806 -16698
rect 12748 -17286 12760 -16710
rect 12794 -17286 12806 -16710
rect 12748 -17298 12806 -17286
rect 13766 -16710 13824 -16698
rect 13766 -17286 13778 -16710
rect 13812 -17286 13824 -16710
rect 13766 -17298 13824 -17286
rect 14784 -16710 14842 -16698
rect 14784 -17286 14796 -16710
rect 14830 -17286 14842 -16710
rect 14784 -17298 14842 -17286
rect 15802 -16710 15860 -16698
rect 15802 -17286 15814 -16710
rect 15848 -17286 15860 -16710
rect 15802 -17298 15860 -17286
rect 16820 -16710 16878 -16698
rect 16820 -17286 16832 -16710
rect 16866 -17286 16878 -16710
rect 16820 -17298 16878 -17286
rect 17838 -16710 17896 -16698
rect 17838 -17286 17850 -16710
rect 17884 -17286 17896 -16710
rect 17838 -17298 17896 -17286
rect 18856 -16710 18914 -16698
rect 18856 -17286 18868 -16710
rect 18902 -17286 18914 -16710
rect 18856 -17298 18914 -17286
rect 19874 -16710 19932 -16698
rect 19874 -17286 19886 -16710
rect 19920 -17286 19932 -16710
rect 19874 -17298 19932 -17286
rect 20892 -16710 20950 -16698
rect 20892 -17286 20904 -16710
rect 20938 -17286 20950 -16710
rect 20892 -17298 20950 -17286
rect 21910 -16710 21968 -16698
rect 21910 -17286 21922 -16710
rect 21956 -17286 21968 -16710
rect 21910 -17298 21968 -17286
rect 22928 -16710 22986 -16698
rect 22928 -17286 22940 -16710
rect 22974 -17286 22986 -16710
rect 22928 -17298 22986 -17286
rect -9196 -17432 -9138 -17420
rect -9196 -18008 -9184 -17432
rect -9150 -18008 -9138 -17432
rect -9196 -18020 -9138 -18008
rect -8178 -17432 -8120 -17420
rect -8178 -18008 -8166 -17432
rect -8132 -18008 -8120 -17432
rect -8178 -18020 -8120 -18008
rect -7160 -17432 -7102 -17420
rect -7160 -18008 -7148 -17432
rect -7114 -18008 -7102 -17432
rect -7160 -18020 -7102 -18008
rect -6142 -17432 -6084 -17420
rect -6142 -18008 -6130 -17432
rect -6096 -18008 -6084 -17432
rect -6142 -18020 -6084 -18008
rect -5124 -17432 -5066 -17420
rect -5124 -18008 -5112 -17432
rect -5078 -18008 -5066 -17432
rect -5124 -18020 -5066 -18008
rect -4106 -17432 -4048 -17420
rect -4106 -18008 -4094 -17432
rect -4060 -18008 -4048 -17432
rect -4106 -18020 -4048 -18008
rect -3088 -17432 -3030 -17420
rect -3088 -18008 -3076 -17432
rect -3042 -18008 -3030 -17432
rect -3088 -18020 -3030 -18008
rect -2070 -17432 -2012 -17420
rect -2070 -18008 -2058 -17432
rect -2024 -18008 -2012 -17432
rect -2070 -18020 -2012 -18008
rect -1052 -17432 -994 -17420
rect -1052 -18008 -1040 -17432
rect -1006 -18008 -994 -17432
rect -1052 -18020 -994 -18008
rect -34 -17432 24 -17420
rect -34 -18008 -22 -17432
rect 12 -18008 24 -17432
rect -34 -18020 24 -18008
rect 2568 -17944 2626 -17932
rect -9196 -18250 -9138 -18238
rect -9196 -18826 -9184 -18250
rect -9150 -18826 -9138 -18250
rect -9196 -18838 -9138 -18826
rect -8178 -18250 -8120 -18238
rect -8178 -18826 -8166 -18250
rect -8132 -18826 -8120 -18250
rect -8178 -18838 -8120 -18826
rect -7160 -18250 -7102 -18238
rect -7160 -18826 -7148 -18250
rect -7114 -18826 -7102 -18250
rect -7160 -18838 -7102 -18826
rect -6142 -18250 -6084 -18238
rect -6142 -18826 -6130 -18250
rect -6096 -18826 -6084 -18250
rect -6142 -18838 -6084 -18826
rect -5124 -18250 -5066 -18238
rect -5124 -18826 -5112 -18250
rect -5078 -18826 -5066 -18250
rect -5124 -18838 -5066 -18826
rect -4106 -18250 -4048 -18238
rect -4106 -18826 -4094 -18250
rect -4060 -18826 -4048 -18250
rect -4106 -18838 -4048 -18826
rect -3088 -18250 -3030 -18238
rect -3088 -18826 -3076 -18250
rect -3042 -18826 -3030 -18250
rect -3088 -18838 -3030 -18826
rect -2070 -18250 -2012 -18238
rect -2070 -18826 -2058 -18250
rect -2024 -18826 -2012 -18250
rect -2070 -18838 -2012 -18826
rect -1052 -18250 -994 -18238
rect -1052 -18826 -1040 -18250
rect -1006 -18826 -994 -18250
rect -1052 -18838 -994 -18826
rect -34 -18250 24 -18238
rect -34 -18826 -22 -18250
rect 12 -18826 24 -18250
rect 2568 -18520 2580 -17944
rect 2614 -18520 2626 -17944
rect 2568 -18532 2626 -18520
rect 3586 -17944 3644 -17932
rect 3586 -18520 3598 -17944
rect 3632 -18520 3644 -17944
rect 3586 -18532 3644 -18520
rect 4604 -17944 4662 -17932
rect 4604 -18520 4616 -17944
rect 4650 -18520 4662 -17944
rect 4604 -18532 4662 -18520
rect 5622 -17944 5680 -17932
rect 5622 -18520 5634 -17944
rect 5668 -18520 5680 -17944
rect 5622 -18532 5680 -18520
rect 6640 -17944 6698 -17932
rect 6640 -18520 6652 -17944
rect 6686 -18520 6698 -17944
rect 6640 -18532 6698 -18520
rect 7658 -17944 7716 -17932
rect 7658 -18520 7670 -17944
rect 7704 -18520 7716 -17944
rect 7658 -18532 7716 -18520
rect 8676 -17944 8734 -17932
rect 8676 -18520 8688 -17944
rect 8722 -18520 8734 -17944
rect 8676 -18532 8734 -18520
rect 9694 -17944 9752 -17932
rect 9694 -18520 9706 -17944
rect 9740 -18520 9752 -17944
rect 9694 -18532 9752 -18520
rect 10712 -17944 10770 -17932
rect 10712 -18520 10724 -17944
rect 10758 -18520 10770 -17944
rect 10712 -18532 10770 -18520
rect 11730 -17944 11788 -17932
rect 11730 -18520 11742 -17944
rect 11776 -18520 11788 -17944
rect 11730 -18532 11788 -18520
rect 12748 -17944 12806 -17932
rect 12748 -18520 12760 -17944
rect 12794 -18520 12806 -17944
rect 12748 -18532 12806 -18520
rect 13766 -17944 13824 -17932
rect 13766 -18520 13778 -17944
rect 13812 -18520 13824 -17944
rect 13766 -18532 13824 -18520
rect 14784 -17944 14842 -17932
rect 14784 -18520 14796 -17944
rect 14830 -18520 14842 -17944
rect 14784 -18532 14842 -18520
rect 15802 -17944 15860 -17932
rect 15802 -18520 15814 -17944
rect 15848 -18520 15860 -17944
rect 15802 -18532 15860 -18520
rect 16820 -17944 16878 -17932
rect 16820 -18520 16832 -17944
rect 16866 -18520 16878 -17944
rect 16820 -18532 16878 -18520
rect 17838 -17944 17896 -17932
rect 17838 -18520 17850 -17944
rect 17884 -18520 17896 -17944
rect 17838 -18532 17896 -18520
rect 18856 -17944 18914 -17932
rect 18856 -18520 18868 -17944
rect 18902 -18520 18914 -17944
rect 18856 -18532 18914 -18520
rect 19874 -17944 19932 -17932
rect 19874 -18520 19886 -17944
rect 19920 -18520 19932 -17944
rect 19874 -18532 19932 -18520
rect 20892 -17944 20950 -17932
rect 20892 -18520 20904 -17944
rect 20938 -18520 20950 -17944
rect 20892 -18532 20950 -18520
rect 21910 -17944 21968 -17932
rect 21910 -18520 21922 -17944
rect 21956 -18520 21968 -17944
rect 21910 -18532 21968 -18520
rect 22928 -17944 22986 -17932
rect 22928 -18520 22940 -17944
rect 22974 -18520 22986 -17944
rect 22928 -18532 22986 -18520
rect -34 -18838 24 -18826
rect 2568 -19176 2626 -19164
rect 2568 -19752 2580 -19176
rect 2614 -19752 2626 -19176
rect 2568 -19764 2626 -19752
rect 3586 -19176 3644 -19164
rect 3586 -19752 3598 -19176
rect 3632 -19752 3644 -19176
rect 3586 -19764 3644 -19752
rect 4604 -19176 4662 -19164
rect 4604 -19752 4616 -19176
rect 4650 -19752 4662 -19176
rect 4604 -19764 4662 -19752
rect 5622 -19176 5680 -19164
rect 5622 -19752 5634 -19176
rect 5668 -19752 5680 -19176
rect 5622 -19764 5680 -19752
rect 6640 -19176 6698 -19164
rect 6640 -19752 6652 -19176
rect 6686 -19752 6698 -19176
rect 6640 -19764 6698 -19752
rect 7658 -19176 7716 -19164
rect 7658 -19752 7670 -19176
rect 7704 -19752 7716 -19176
rect 7658 -19764 7716 -19752
rect 8676 -19176 8734 -19164
rect 8676 -19752 8688 -19176
rect 8722 -19752 8734 -19176
rect 8676 -19764 8734 -19752
rect 9694 -19176 9752 -19164
rect 9694 -19752 9706 -19176
rect 9740 -19752 9752 -19176
rect 9694 -19764 9752 -19752
rect 10712 -19176 10770 -19164
rect 10712 -19752 10724 -19176
rect 10758 -19752 10770 -19176
rect 10712 -19764 10770 -19752
rect 11730 -19176 11788 -19164
rect 11730 -19752 11742 -19176
rect 11776 -19752 11788 -19176
rect 11730 -19764 11788 -19752
rect 12748 -19176 12806 -19164
rect 12748 -19752 12760 -19176
rect 12794 -19752 12806 -19176
rect 12748 -19764 12806 -19752
rect 13766 -19176 13824 -19164
rect 13766 -19752 13778 -19176
rect 13812 -19752 13824 -19176
rect 13766 -19764 13824 -19752
rect 14784 -19176 14842 -19164
rect 14784 -19752 14796 -19176
rect 14830 -19752 14842 -19176
rect 14784 -19764 14842 -19752
rect 15802 -19176 15860 -19164
rect 15802 -19752 15814 -19176
rect 15848 -19752 15860 -19176
rect 15802 -19764 15860 -19752
rect 16820 -19176 16878 -19164
rect 16820 -19752 16832 -19176
rect 16866 -19752 16878 -19176
rect 16820 -19764 16878 -19752
rect 17838 -19176 17896 -19164
rect 17838 -19752 17850 -19176
rect 17884 -19752 17896 -19176
rect 17838 -19764 17896 -19752
rect 18856 -19176 18914 -19164
rect 18856 -19752 18868 -19176
rect 18902 -19752 18914 -19176
rect 18856 -19764 18914 -19752
rect 19874 -19176 19932 -19164
rect 19874 -19752 19886 -19176
rect 19920 -19752 19932 -19176
rect 19874 -19764 19932 -19752
rect 20892 -19176 20950 -19164
rect 20892 -19752 20904 -19176
rect 20938 -19752 20950 -19176
rect 20892 -19764 20950 -19752
rect 21910 -19176 21968 -19164
rect 21910 -19752 21922 -19176
rect 21956 -19752 21968 -19176
rect 21910 -19764 21968 -19752
rect 22928 -19176 22986 -19164
rect 22928 -19752 22940 -19176
rect 22974 -19752 22986 -19176
rect 22928 -19764 22986 -19752
rect -10520 -20274 -10462 -20262
rect -10520 -20850 -10508 -20274
rect -10474 -20850 -10462 -20274
rect -10520 -20862 -10462 -20850
rect -9502 -20274 -9444 -20262
rect -9502 -20850 -9490 -20274
rect -9456 -20850 -9444 -20274
rect -9502 -20862 -9444 -20850
rect -8484 -20274 -8426 -20262
rect -8484 -20850 -8472 -20274
rect -8438 -20850 -8426 -20274
rect -8484 -20862 -8426 -20850
rect -7466 -20274 -7408 -20262
rect -7466 -20850 -7454 -20274
rect -7420 -20850 -7408 -20274
rect -7466 -20862 -7408 -20850
rect -6448 -20274 -6390 -20262
rect -6448 -20850 -6436 -20274
rect -6402 -20850 -6390 -20274
rect -6448 -20862 -6390 -20850
rect -5430 -20274 -5372 -20262
rect -5430 -20850 -5418 -20274
rect -5384 -20850 -5372 -20274
rect -5430 -20862 -5372 -20850
rect -4412 -20274 -4354 -20262
rect -4412 -20850 -4400 -20274
rect -4366 -20850 -4354 -20274
rect -4412 -20862 -4354 -20850
rect -3394 -20274 -3336 -20262
rect -3394 -20850 -3382 -20274
rect -3348 -20850 -3336 -20274
rect -3394 -20862 -3336 -20850
rect -2376 -20274 -2318 -20262
rect -2376 -20850 -2364 -20274
rect -2330 -20850 -2318 -20274
rect -2376 -20862 -2318 -20850
rect -1358 -20274 -1300 -20262
rect -1358 -20850 -1346 -20274
rect -1312 -20850 -1300 -20274
rect -1358 -20862 -1300 -20850
rect -340 -20274 -282 -20262
rect -340 -20850 -328 -20274
rect -294 -20850 -282 -20274
rect -340 -20862 -282 -20850
rect 678 -20274 736 -20262
rect 678 -20850 690 -20274
rect 724 -20850 736 -20274
rect 678 -20862 736 -20850
rect 2568 -20410 2626 -20398
rect 2568 -20986 2580 -20410
rect 2614 -20986 2626 -20410
rect 2568 -20998 2626 -20986
rect 3586 -20410 3644 -20398
rect 3586 -20986 3598 -20410
rect 3632 -20986 3644 -20410
rect 3586 -20998 3644 -20986
rect 4604 -20410 4662 -20398
rect 4604 -20986 4616 -20410
rect 4650 -20986 4662 -20410
rect 4604 -20998 4662 -20986
rect 5622 -20410 5680 -20398
rect 5622 -20986 5634 -20410
rect 5668 -20986 5680 -20410
rect 5622 -20998 5680 -20986
rect 6640 -20410 6698 -20398
rect 6640 -20986 6652 -20410
rect 6686 -20986 6698 -20410
rect 6640 -20998 6698 -20986
rect 7658 -20410 7716 -20398
rect 7658 -20986 7670 -20410
rect 7704 -20986 7716 -20410
rect 7658 -20998 7716 -20986
rect 8676 -20410 8734 -20398
rect 8676 -20986 8688 -20410
rect 8722 -20986 8734 -20410
rect 8676 -20998 8734 -20986
rect 9694 -20410 9752 -20398
rect 9694 -20986 9706 -20410
rect 9740 -20986 9752 -20410
rect 9694 -20998 9752 -20986
rect 10712 -20410 10770 -20398
rect 10712 -20986 10724 -20410
rect 10758 -20986 10770 -20410
rect 10712 -20998 10770 -20986
rect 11730 -20410 11788 -20398
rect 11730 -20986 11742 -20410
rect 11776 -20986 11788 -20410
rect 11730 -20998 11788 -20986
rect 12748 -20410 12806 -20398
rect 12748 -20986 12760 -20410
rect 12794 -20986 12806 -20410
rect 12748 -20998 12806 -20986
rect 13766 -20410 13824 -20398
rect 13766 -20986 13778 -20410
rect 13812 -20986 13824 -20410
rect 13766 -20998 13824 -20986
rect 14784 -20410 14842 -20398
rect 14784 -20986 14796 -20410
rect 14830 -20986 14842 -20410
rect 14784 -20998 14842 -20986
rect 15802 -20410 15860 -20398
rect 15802 -20986 15814 -20410
rect 15848 -20986 15860 -20410
rect 15802 -20998 15860 -20986
rect 16820 -20410 16878 -20398
rect 16820 -20986 16832 -20410
rect 16866 -20986 16878 -20410
rect 16820 -20998 16878 -20986
rect 17838 -20410 17896 -20398
rect 17838 -20986 17850 -20410
rect 17884 -20986 17896 -20410
rect 17838 -20998 17896 -20986
rect 18856 -20410 18914 -20398
rect 18856 -20986 18868 -20410
rect 18902 -20986 18914 -20410
rect 18856 -20998 18914 -20986
rect 19874 -20410 19932 -20398
rect 19874 -20986 19886 -20410
rect 19920 -20986 19932 -20410
rect 19874 -20998 19932 -20986
rect 20892 -20410 20950 -20398
rect 20892 -20986 20904 -20410
rect 20938 -20986 20950 -20410
rect 20892 -20998 20950 -20986
rect 21910 -20410 21968 -20398
rect 21910 -20986 21922 -20410
rect 21956 -20986 21968 -20410
rect 21910 -20998 21968 -20986
rect 22928 -20410 22986 -20398
rect 22928 -20986 22940 -20410
rect 22974 -20986 22986 -20410
rect 22928 -20998 22986 -20986
rect -10520 -21386 -10462 -21374
rect -10520 -21962 -10508 -21386
rect -10474 -21962 -10462 -21386
rect -10520 -21974 -10462 -21962
rect -9502 -21386 -9444 -21374
rect -9502 -21962 -9490 -21386
rect -9456 -21962 -9444 -21386
rect -9502 -21974 -9444 -21962
rect -8484 -21386 -8426 -21374
rect -8484 -21962 -8472 -21386
rect -8438 -21962 -8426 -21386
rect -8484 -21974 -8426 -21962
rect -7466 -21386 -7408 -21374
rect -7466 -21962 -7454 -21386
rect -7420 -21962 -7408 -21386
rect -7466 -21974 -7408 -21962
rect -6448 -21386 -6390 -21374
rect -6448 -21962 -6436 -21386
rect -6402 -21962 -6390 -21386
rect -6448 -21974 -6390 -21962
rect -5430 -21386 -5372 -21374
rect -5430 -21962 -5418 -21386
rect -5384 -21962 -5372 -21386
rect -5430 -21974 -5372 -21962
rect -4412 -21386 -4354 -21374
rect -4412 -21962 -4400 -21386
rect -4366 -21962 -4354 -21386
rect -4412 -21974 -4354 -21962
rect -3394 -21386 -3336 -21374
rect -3394 -21962 -3382 -21386
rect -3348 -21962 -3336 -21386
rect -3394 -21974 -3336 -21962
rect -2376 -21386 -2318 -21374
rect -2376 -21962 -2364 -21386
rect -2330 -21962 -2318 -21386
rect -2376 -21974 -2318 -21962
rect -1358 -21386 -1300 -21374
rect -1358 -21962 -1346 -21386
rect -1312 -21962 -1300 -21386
rect -1358 -21974 -1300 -21962
rect -340 -21386 -282 -21374
rect -340 -21962 -328 -21386
rect -294 -21962 -282 -21386
rect -340 -21974 -282 -21962
rect 678 -21386 736 -21374
rect 678 -21962 690 -21386
rect 724 -21962 736 -21386
rect 678 -21974 736 -21962
rect 2568 -21644 2626 -21632
rect 2568 -22220 2580 -21644
rect 2614 -22220 2626 -21644
rect 2568 -22232 2626 -22220
rect 3586 -21644 3644 -21632
rect 3586 -22220 3598 -21644
rect 3632 -22220 3644 -21644
rect 3586 -22232 3644 -22220
rect 4604 -21644 4662 -21632
rect 4604 -22220 4616 -21644
rect 4650 -22220 4662 -21644
rect 4604 -22232 4662 -22220
rect 5622 -21644 5680 -21632
rect 5622 -22220 5634 -21644
rect 5668 -22220 5680 -21644
rect 5622 -22232 5680 -22220
rect 6640 -21644 6698 -21632
rect 6640 -22220 6652 -21644
rect 6686 -22220 6698 -21644
rect 6640 -22232 6698 -22220
rect 7658 -21644 7716 -21632
rect 7658 -22220 7670 -21644
rect 7704 -22220 7716 -21644
rect 7658 -22232 7716 -22220
rect 8676 -21644 8734 -21632
rect 8676 -22220 8688 -21644
rect 8722 -22220 8734 -21644
rect 8676 -22232 8734 -22220
rect 9694 -21644 9752 -21632
rect 9694 -22220 9706 -21644
rect 9740 -22220 9752 -21644
rect 9694 -22232 9752 -22220
rect 10712 -21644 10770 -21632
rect 10712 -22220 10724 -21644
rect 10758 -22220 10770 -21644
rect 10712 -22232 10770 -22220
rect 11730 -21644 11788 -21632
rect 11730 -22220 11742 -21644
rect 11776 -22220 11788 -21644
rect 11730 -22232 11788 -22220
rect 12748 -21644 12806 -21632
rect 12748 -22220 12760 -21644
rect 12794 -22220 12806 -21644
rect 12748 -22232 12806 -22220
rect 13766 -21644 13824 -21632
rect 13766 -22220 13778 -21644
rect 13812 -22220 13824 -21644
rect 13766 -22232 13824 -22220
rect 14784 -21644 14842 -21632
rect 14784 -22220 14796 -21644
rect 14830 -22220 14842 -21644
rect 14784 -22232 14842 -22220
rect 15802 -21644 15860 -21632
rect 15802 -22220 15814 -21644
rect 15848 -22220 15860 -21644
rect 15802 -22232 15860 -22220
rect 16820 -21644 16878 -21632
rect 16820 -22220 16832 -21644
rect 16866 -22220 16878 -21644
rect 16820 -22232 16878 -22220
rect 17838 -21644 17896 -21632
rect 17838 -22220 17850 -21644
rect 17884 -22220 17896 -21644
rect 17838 -22232 17896 -22220
rect 18856 -21644 18914 -21632
rect 18856 -22220 18868 -21644
rect 18902 -22220 18914 -21644
rect 18856 -22232 18914 -22220
rect 19874 -21644 19932 -21632
rect 19874 -22220 19886 -21644
rect 19920 -22220 19932 -21644
rect 19874 -22232 19932 -22220
rect 20892 -21644 20950 -21632
rect 20892 -22220 20904 -21644
rect 20938 -22220 20950 -21644
rect 20892 -22232 20950 -22220
rect 21910 -21644 21968 -21632
rect 21910 -22220 21922 -21644
rect 21956 -22220 21968 -21644
rect 21910 -22232 21968 -22220
rect 22928 -21644 22986 -21632
rect 22928 -22220 22940 -21644
rect 22974 -22220 22986 -21644
rect 22928 -22232 22986 -22220
rect -10520 -22498 -10462 -22486
rect -10520 -23074 -10508 -22498
rect -10474 -23074 -10462 -22498
rect -10520 -23086 -10462 -23074
rect -9502 -22498 -9444 -22486
rect -9502 -23074 -9490 -22498
rect -9456 -23074 -9444 -22498
rect -9502 -23086 -9444 -23074
rect -8484 -22498 -8426 -22486
rect -8484 -23074 -8472 -22498
rect -8438 -23074 -8426 -22498
rect -8484 -23086 -8426 -23074
rect -7466 -22498 -7408 -22486
rect -7466 -23074 -7454 -22498
rect -7420 -23074 -7408 -22498
rect -7466 -23086 -7408 -23074
rect -6448 -22498 -6390 -22486
rect -6448 -23074 -6436 -22498
rect -6402 -23074 -6390 -22498
rect -6448 -23086 -6390 -23074
rect -5430 -22498 -5372 -22486
rect -5430 -23074 -5418 -22498
rect -5384 -23074 -5372 -22498
rect -5430 -23086 -5372 -23074
rect -4412 -22498 -4354 -22486
rect -4412 -23074 -4400 -22498
rect -4366 -23074 -4354 -22498
rect -4412 -23086 -4354 -23074
rect -3394 -22498 -3336 -22486
rect -3394 -23074 -3382 -22498
rect -3348 -23074 -3336 -22498
rect -3394 -23086 -3336 -23074
rect -2376 -22498 -2318 -22486
rect -2376 -23074 -2364 -22498
rect -2330 -23074 -2318 -22498
rect -2376 -23086 -2318 -23074
rect -1358 -22498 -1300 -22486
rect -1358 -23074 -1346 -22498
rect -1312 -23074 -1300 -22498
rect -1358 -23086 -1300 -23074
rect -340 -22498 -282 -22486
rect -340 -23074 -328 -22498
rect -294 -23074 -282 -22498
rect -340 -23086 -282 -23074
rect 678 -22498 736 -22486
rect 678 -23074 690 -22498
rect 724 -23074 736 -22498
rect 678 -23086 736 -23074
rect 2568 -22876 2626 -22864
rect 2568 -23452 2580 -22876
rect 2614 -23452 2626 -22876
rect 2568 -23464 2626 -23452
rect 3586 -22876 3644 -22864
rect 3586 -23452 3598 -22876
rect 3632 -23452 3644 -22876
rect 3586 -23464 3644 -23452
rect 4604 -22876 4662 -22864
rect 4604 -23452 4616 -22876
rect 4650 -23452 4662 -22876
rect 4604 -23464 4662 -23452
rect 5622 -22876 5680 -22864
rect 5622 -23452 5634 -22876
rect 5668 -23452 5680 -22876
rect 5622 -23464 5680 -23452
rect 6640 -22876 6698 -22864
rect 6640 -23452 6652 -22876
rect 6686 -23452 6698 -22876
rect 6640 -23464 6698 -23452
rect 7658 -22876 7716 -22864
rect 7658 -23452 7670 -22876
rect 7704 -23452 7716 -22876
rect 7658 -23464 7716 -23452
rect 8676 -22876 8734 -22864
rect 8676 -23452 8688 -22876
rect 8722 -23452 8734 -22876
rect 8676 -23464 8734 -23452
rect 9694 -22876 9752 -22864
rect 9694 -23452 9706 -22876
rect 9740 -23452 9752 -22876
rect 9694 -23464 9752 -23452
rect 10712 -22876 10770 -22864
rect 10712 -23452 10724 -22876
rect 10758 -23452 10770 -22876
rect 10712 -23464 10770 -23452
rect 11730 -22876 11788 -22864
rect 11730 -23452 11742 -22876
rect 11776 -23452 11788 -22876
rect 11730 -23464 11788 -23452
rect 12748 -22876 12806 -22864
rect 12748 -23452 12760 -22876
rect 12794 -23452 12806 -22876
rect 12748 -23464 12806 -23452
rect 13766 -22876 13824 -22864
rect 13766 -23452 13778 -22876
rect 13812 -23452 13824 -22876
rect 13766 -23464 13824 -23452
rect 14784 -22876 14842 -22864
rect 14784 -23452 14796 -22876
rect 14830 -23452 14842 -22876
rect 14784 -23464 14842 -23452
rect 15802 -22876 15860 -22864
rect 15802 -23452 15814 -22876
rect 15848 -23452 15860 -22876
rect 15802 -23464 15860 -23452
rect 16820 -22876 16878 -22864
rect 16820 -23452 16832 -22876
rect 16866 -23452 16878 -22876
rect 16820 -23464 16878 -23452
rect 17838 -22876 17896 -22864
rect 17838 -23452 17850 -22876
rect 17884 -23452 17896 -22876
rect 17838 -23464 17896 -23452
rect 18856 -22876 18914 -22864
rect 18856 -23452 18868 -22876
rect 18902 -23452 18914 -22876
rect 18856 -23464 18914 -23452
rect 19874 -22876 19932 -22864
rect 19874 -23452 19886 -22876
rect 19920 -23452 19932 -22876
rect 19874 -23464 19932 -23452
rect 20892 -22876 20950 -22864
rect 20892 -23452 20904 -22876
rect 20938 -23452 20950 -22876
rect 20892 -23464 20950 -23452
rect 21910 -22876 21968 -22864
rect 21910 -23452 21922 -22876
rect 21956 -23452 21968 -22876
rect 21910 -23464 21968 -23452
rect 22928 -22876 22986 -22864
rect 22928 -23452 22940 -22876
rect 22974 -23452 22986 -22876
rect 22928 -23464 22986 -23452
rect -10520 -23610 -10462 -23598
rect -10520 -24186 -10508 -23610
rect -10474 -24186 -10462 -23610
rect -10520 -24198 -10462 -24186
rect -9502 -23610 -9444 -23598
rect -9502 -24186 -9490 -23610
rect -9456 -24186 -9444 -23610
rect -9502 -24198 -9444 -24186
rect -8484 -23610 -8426 -23598
rect -8484 -24186 -8472 -23610
rect -8438 -24186 -8426 -23610
rect -8484 -24198 -8426 -24186
rect -7466 -23610 -7408 -23598
rect -7466 -24186 -7454 -23610
rect -7420 -24186 -7408 -23610
rect -7466 -24198 -7408 -24186
rect -6448 -23610 -6390 -23598
rect -6448 -24186 -6436 -23610
rect -6402 -24186 -6390 -23610
rect -6448 -24198 -6390 -24186
rect -5430 -23610 -5372 -23598
rect -5430 -24186 -5418 -23610
rect -5384 -24186 -5372 -23610
rect -5430 -24198 -5372 -24186
rect -4412 -23610 -4354 -23598
rect -4412 -24186 -4400 -23610
rect -4366 -24186 -4354 -23610
rect -4412 -24198 -4354 -24186
rect -3394 -23610 -3336 -23598
rect -3394 -24186 -3382 -23610
rect -3348 -24186 -3336 -23610
rect -3394 -24198 -3336 -24186
rect -2376 -23610 -2318 -23598
rect -2376 -24186 -2364 -23610
rect -2330 -24186 -2318 -23610
rect -2376 -24198 -2318 -24186
rect -1358 -23610 -1300 -23598
rect -1358 -24186 -1346 -23610
rect -1312 -24186 -1300 -23610
rect -1358 -24198 -1300 -24186
rect -340 -23610 -282 -23598
rect -340 -24186 -328 -23610
rect -294 -24186 -282 -23610
rect -340 -24198 -282 -24186
rect 678 -23610 736 -23598
rect 678 -24186 690 -23610
rect 724 -24186 736 -23610
rect 678 -24198 736 -24186
rect 2568 -24110 2626 -24098
rect 2568 -24686 2580 -24110
rect 2614 -24686 2626 -24110
rect 2568 -24698 2626 -24686
rect 3586 -24110 3644 -24098
rect 3586 -24686 3598 -24110
rect 3632 -24686 3644 -24110
rect 3586 -24698 3644 -24686
rect 4604 -24110 4662 -24098
rect 4604 -24686 4616 -24110
rect 4650 -24686 4662 -24110
rect 4604 -24698 4662 -24686
rect 5622 -24110 5680 -24098
rect 5622 -24686 5634 -24110
rect 5668 -24686 5680 -24110
rect 5622 -24698 5680 -24686
rect 6640 -24110 6698 -24098
rect 6640 -24686 6652 -24110
rect 6686 -24686 6698 -24110
rect 6640 -24698 6698 -24686
rect 7658 -24110 7716 -24098
rect 7658 -24686 7670 -24110
rect 7704 -24686 7716 -24110
rect 7658 -24698 7716 -24686
rect 8676 -24110 8734 -24098
rect 8676 -24686 8688 -24110
rect 8722 -24686 8734 -24110
rect 8676 -24698 8734 -24686
rect 9694 -24110 9752 -24098
rect 9694 -24686 9706 -24110
rect 9740 -24686 9752 -24110
rect 9694 -24698 9752 -24686
rect 10712 -24110 10770 -24098
rect 10712 -24686 10724 -24110
rect 10758 -24686 10770 -24110
rect 10712 -24698 10770 -24686
rect 11730 -24110 11788 -24098
rect 11730 -24686 11742 -24110
rect 11776 -24686 11788 -24110
rect 11730 -24698 11788 -24686
rect 12748 -24110 12806 -24098
rect 12748 -24686 12760 -24110
rect 12794 -24686 12806 -24110
rect 12748 -24698 12806 -24686
rect 13766 -24110 13824 -24098
rect 13766 -24686 13778 -24110
rect 13812 -24686 13824 -24110
rect 13766 -24698 13824 -24686
rect 14784 -24110 14842 -24098
rect 14784 -24686 14796 -24110
rect 14830 -24686 14842 -24110
rect 14784 -24698 14842 -24686
rect 15802 -24110 15860 -24098
rect 15802 -24686 15814 -24110
rect 15848 -24686 15860 -24110
rect 15802 -24698 15860 -24686
rect 16820 -24110 16878 -24098
rect 16820 -24686 16832 -24110
rect 16866 -24686 16878 -24110
rect 16820 -24698 16878 -24686
rect 17838 -24110 17896 -24098
rect 17838 -24686 17850 -24110
rect 17884 -24686 17896 -24110
rect 17838 -24698 17896 -24686
rect 18856 -24110 18914 -24098
rect 18856 -24686 18868 -24110
rect 18902 -24686 18914 -24110
rect 18856 -24698 18914 -24686
rect 19874 -24110 19932 -24098
rect 19874 -24686 19886 -24110
rect 19920 -24686 19932 -24110
rect 19874 -24698 19932 -24686
rect 20892 -24110 20950 -24098
rect 20892 -24686 20904 -24110
rect 20938 -24686 20950 -24110
rect 20892 -24698 20950 -24686
rect 21910 -24110 21968 -24098
rect 21910 -24686 21922 -24110
rect 21956 -24686 21968 -24110
rect 21910 -24698 21968 -24686
rect 22928 -24110 22986 -24098
rect 22928 -24686 22940 -24110
rect 22974 -24686 22986 -24110
rect 22928 -24698 22986 -24686
rect -10062 -25152 -10004 -25140
rect -10062 -25728 -10050 -25152
rect -10016 -25728 -10004 -25152
rect -10062 -25740 -10004 -25728
rect -9044 -25152 -8986 -25140
rect -9044 -25728 -9032 -25152
rect -8998 -25728 -8986 -25152
rect -9044 -25740 -8986 -25728
rect -8026 -25152 -7968 -25140
rect -8026 -25728 -8014 -25152
rect -7980 -25728 -7968 -25152
rect -8026 -25740 -7968 -25728
rect -7008 -25152 -6950 -25140
rect -7008 -25728 -6996 -25152
rect -6962 -25728 -6950 -25152
rect -7008 -25740 -6950 -25728
rect -5990 -25152 -5932 -25140
rect -5990 -25728 -5978 -25152
rect -5944 -25728 -5932 -25152
rect -5990 -25740 -5932 -25728
rect -4972 -25152 -4914 -25140
rect -4972 -25728 -4960 -25152
rect -4926 -25728 -4914 -25152
rect -4972 -25740 -4914 -25728
rect -3954 -25152 -3896 -25140
rect -3954 -25728 -3942 -25152
rect -3908 -25728 -3896 -25152
rect -3954 -25740 -3896 -25728
rect -2936 -25152 -2878 -25140
rect -2936 -25728 -2924 -25152
rect -2890 -25728 -2878 -25152
rect -2936 -25740 -2878 -25728
rect -1918 -25152 -1860 -25140
rect -1918 -25728 -1906 -25152
rect -1872 -25728 -1860 -25152
rect -1918 -25740 -1860 -25728
rect -900 -25152 -842 -25140
rect -900 -25728 -888 -25152
rect -854 -25728 -842 -25152
rect -900 -25740 -842 -25728
rect 118 -25152 176 -25140
rect 118 -25728 130 -25152
rect 164 -25728 176 -25152
rect 118 -25740 176 -25728
rect 2568 -25342 2626 -25330
rect 2568 -25918 2580 -25342
rect 2614 -25918 2626 -25342
rect 2568 -25930 2626 -25918
rect 3586 -25342 3644 -25330
rect 3586 -25918 3598 -25342
rect 3632 -25918 3644 -25342
rect 3586 -25930 3644 -25918
rect 4604 -25342 4662 -25330
rect 4604 -25918 4616 -25342
rect 4650 -25918 4662 -25342
rect 4604 -25930 4662 -25918
rect 5622 -25342 5680 -25330
rect 5622 -25918 5634 -25342
rect 5668 -25918 5680 -25342
rect 5622 -25930 5680 -25918
rect 6640 -25342 6698 -25330
rect 6640 -25918 6652 -25342
rect 6686 -25918 6698 -25342
rect 6640 -25930 6698 -25918
rect 7658 -25342 7716 -25330
rect 7658 -25918 7670 -25342
rect 7704 -25918 7716 -25342
rect 7658 -25930 7716 -25918
rect 8676 -25342 8734 -25330
rect 8676 -25918 8688 -25342
rect 8722 -25918 8734 -25342
rect 8676 -25930 8734 -25918
rect 9694 -25342 9752 -25330
rect 9694 -25918 9706 -25342
rect 9740 -25918 9752 -25342
rect 9694 -25930 9752 -25918
rect 10712 -25342 10770 -25330
rect 10712 -25918 10724 -25342
rect 10758 -25918 10770 -25342
rect 10712 -25930 10770 -25918
rect 11730 -25342 11788 -25330
rect 11730 -25918 11742 -25342
rect 11776 -25918 11788 -25342
rect 11730 -25930 11788 -25918
rect 12748 -25342 12806 -25330
rect 12748 -25918 12760 -25342
rect 12794 -25918 12806 -25342
rect 12748 -25930 12806 -25918
rect 13766 -25342 13824 -25330
rect 13766 -25918 13778 -25342
rect 13812 -25918 13824 -25342
rect 13766 -25930 13824 -25918
rect 14784 -25342 14842 -25330
rect 14784 -25918 14796 -25342
rect 14830 -25918 14842 -25342
rect 14784 -25930 14842 -25918
rect 15802 -25342 15860 -25330
rect 15802 -25918 15814 -25342
rect 15848 -25918 15860 -25342
rect 15802 -25930 15860 -25918
rect 16820 -25342 16878 -25330
rect 16820 -25918 16832 -25342
rect 16866 -25918 16878 -25342
rect 16820 -25930 16878 -25918
rect 17838 -25342 17896 -25330
rect 17838 -25918 17850 -25342
rect 17884 -25918 17896 -25342
rect 17838 -25930 17896 -25918
rect 18856 -25342 18914 -25330
rect 18856 -25918 18868 -25342
rect 18902 -25918 18914 -25342
rect 18856 -25930 18914 -25918
rect 19874 -25342 19932 -25330
rect 19874 -25918 19886 -25342
rect 19920 -25918 19932 -25342
rect 19874 -25930 19932 -25918
rect 20892 -25342 20950 -25330
rect 20892 -25918 20904 -25342
rect 20938 -25918 20950 -25342
rect 20892 -25930 20950 -25918
rect 21910 -25342 21968 -25330
rect 21910 -25918 21922 -25342
rect 21956 -25918 21968 -25342
rect 21910 -25930 21968 -25918
rect 22928 -25342 22986 -25330
rect 22928 -25918 22940 -25342
rect 22974 -25918 22986 -25342
rect 22928 -25930 22986 -25918
<< pdiff >>
rect 6476 1462 6534 1474
rect 6476 886 6488 1462
rect 6522 886 6534 1462
rect 6476 874 6534 886
rect 7494 1462 7552 1474
rect 7494 886 7506 1462
rect 7540 886 7552 1462
rect 7494 874 7552 886
rect 8512 1462 8570 1474
rect 8512 886 8524 1462
rect 8558 886 8570 1462
rect 8512 874 8570 886
rect 9530 1462 9588 1474
rect 9530 886 9542 1462
rect 9576 886 9588 1462
rect 9530 874 9588 886
rect 10548 1462 10606 1474
rect 10548 886 10560 1462
rect 10594 886 10606 1462
rect 10548 874 10606 886
rect 11566 1462 11624 1474
rect 11566 886 11578 1462
rect 11612 886 11624 1462
rect 11566 874 11624 886
rect 12584 1462 12642 1474
rect 12584 886 12596 1462
rect 12630 886 12642 1462
rect 12584 874 12642 886
rect 13602 1462 13660 1474
rect 13602 886 13614 1462
rect 13648 886 13660 1462
rect 13602 874 13660 886
rect 14620 1462 14678 1474
rect 14620 886 14632 1462
rect 14666 886 14678 1462
rect 14620 874 14678 886
rect 15638 1462 15696 1474
rect 15638 886 15650 1462
rect 15684 886 15696 1462
rect 15638 874 15696 886
rect 16656 1462 16714 1474
rect 16656 886 16668 1462
rect 16702 886 16714 1462
rect 16656 874 16714 886
rect 17674 1462 17732 1474
rect 17674 886 17686 1462
rect 17720 886 17732 1462
rect 17674 874 17732 886
rect 18692 1462 18750 1474
rect 18692 886 18704 1462
rect 18738 886 18750 1462
rect 18692 874 18750 886
rect 19710 1462 19768 1474
rect 19710 886 19722 1462
rect 19756 886 19768 1462
rect 19710 874 19768 886
rect 20728 1462 20786 1474
rect 20728 886 20740 1462
rect 20774 886 20786 1462
rect 20728 874 20786 886
rect 21746 1462 21804 1474
rect 21746 886 21758 1462
rect 21792 886 21804 1462
rect 21746 874 21804 886
rect 22764 1462 22822 1474
rect 22764 886 22776 1462
rect 22810 886 22822 1462
rect 22764 874 22822 886
rect 6476 326 6534 338
rect 6476 -250 6488 326
rect 6522 -250 6534 326
rect 6476 -262 6534 -250
rect 7494 326 7552 338
rect 7494 -250 7506 326
rect 7540 -250 7552 326
rect 7494 -262 7552 -250
rect 8512 326 8570 338
rect 8512 -250 8524 326
rect 8558 -250 8570 326
rect 8512 -262 8570 -250
rect 9530 326 9588 338
rect 9530 -250 9542 326
rect 9576 -250 9588 326
rect 9530 -262 9588 -250
rect 10548 326 10606 338
rect 10548 -250 10560 326
rect 10594 -250 10606 326
rect 10548 -262 10606 -250
rect 11566 326 11624 338
rect 11566 -250 11578 326
rect 11612 -250 11624 326
rect 11566 -262 11624 -250
rect 12584 326 12642 338
rect 12584 -250 12596 326
rect 12630 -250 12642 326
rect 12584 -262 12642 -250
rect 13602 326 13660 338
rect 13602 -250 13614 326
rect 13648 -250 13660 326
rect 13602 -262 13660 -250
rect 14620 326 14678 338
rect 14620 -250 14632 326
rect 14666 -250 14678 326
rect 14620 -262 14678 -250
rect 15638 326 15696 338
rect 15638 -250 15650 326
rect 15684 -250 15696 326
rect 15638 -262 15696 -250
rect 16656 326 16714 338
rect 16656 -250 16668 326
rect 16702 -250 16714 326
rect 16656 -262 16714 -250
rect 17674 326 17732 338
rect 17674 -250 17686 326
rect 17720 -250 17732 326
rect 17674 -262 17732 -250
rect 18692 326 18750 338
rect 18692 -250 18704 326
rect 18738 -250 18750 326
rect 18692 -262 18750 -250
rect 19710 326 19768 338
rect 19710 -250 19722 326
rect 19756 -250 19768 326
rect 19710 -262 19768 -250
rect 20728 326 20786 338
rect 20728 -250 20740 326
rect 20774 -250 20786 326
rect 20728 -262 20786 -250
rect 21746 326 21804 338
rect 21746 -250 21758 326
rect 21792 -250 21804 326
rect 21746 -262 21804 -250
rect 22764 326 22822 338
rect 22764 -250 22776 326
rect 22810 -250 22822 326
rect 22764 -262 22822 -250
rect 6476 -810 6534 -798
rect 6476 -1386 6488 -810
rect 6522 -1386 6534 -810
rect 6476 -1398 6534 -1386
rect 7494 -810 7552 -798
rect 7494 -1386 7506 -810
rect 7540 -1386 7552 -810
rect 7494 -1398 7552 -1386
rect 8512 -810 8570 -798
rect 8512 -1386 8524 -810
rect 8558 -1386 8570 -810
rect 8512 -1398 8570 -1386
rect 9530 -810 9588 -798
rect 9530 -1386 9542 -810
rect 9576 -1386 9588 -810
rect 9530 -1398 9588 -1386
rect 10548 -810 10606 -798
rect 10548 -1386 10560 -810
rect 10594 -1386 10606 -810
rect 10548 -1398 10606 -1386
rect 11566 -810 11624 -798
rect 11566 -1386 11578 -810
rect 11612 -1386 11624 -810
rect 11566 -1398 11624 -1386
rect 12584 -810 12642 -798
rect 12584 -1386 12596 -810
rect 12630 -1386 12642 -810
rect 12584 -1398 12642 -1386
rect 13602 -810 13660 -798
rect 13602 -1386 13614 -810
rect 13648 -1386 13660 -810
rect 13602 -1398 13660 -1386
rect 14620 -810 14678 -798
rect 14620 -1386 14632 -810
rect 14666 -1386 14678 -810
rect 14620 -1398 14678 -1386
rect 15638 -810 15696 -798
rect 15638 -1386 15650 -810
rect 15684 -1386 15696 -810
rect 15638 -1398 15696 -1386
rect 16656 -810 16714 -798
rect 16656 -1386 16668 -810
rect 16702 -1386 16714 -810
rect 16656 -1398 16714 -1386
rect 17674 -810 17732 -798
rect 17674 -1386 17686 -810
rect 17720 -1386 17732 -810
rect 17674 -1398 17732 -1386
rect 18692 -810 18750 -798
rect 18692 -1386 18704 -810
rect 18738 -1386 18750 -810
rect 18692 -1398 18750 -1386
rect 19710 -810 19768 -798
rect 19710 -1386 19722 -810
rect 19756 -1386 19768 -810
rect 19710 -1398 19768 -1386
rect 20728 -810 20786 -798
rect 20728 -1386 20740 -810
rect 20774 -1386 20786 -810
rect 20728 -1398 20786 -1386
rect 21746 -810 21804 -798
rect 21746 -1386 21758 -810
rect 21792 -1386 21804 -810
rect 21746 -1398 21804 -1386
rect 22764 -810 22822 -798
rect 22764 -1386 22776 -810
rect 22810 -1386 22822 -810
rect 22764 -1398 22822 -1386
rect 7670 -2448 7728 -2436
rect 7670 -3024 7682 -2448
rect 7716 -3024 7728 -2448
rect 7670 -3036 7728 -3024
rect 8688 -2448 8746 -2436
rect 8688 -3024 8700 -2448
rect 8734 -3024 8746 -2448
rect 8688 -3036 8746 -3024
rect 9706 -2448 9764 -2436
rect 9706 -3024 9718 -2448
rect 9752 -3024 9764 -2448
rect 9706 -3036 9764 -3024
rect 10724 -2448 10782 -2436
rect 10724 -3024 10736 -2448
rect 10770 -3024 10782 -2448
rect 10724 -3036 10782 -3024
rect 11742 -2448 11800 -2436
rect 11742 -3024 11754 -2448
rect 11788 -3024 11800 -2448
rect 11742 -3036 11800 -3024
rect 12760 -2448 12818 -2436
rect 12760 -3024 12772 -2448
rect 12806 -3024 12818 -2448
rect 12760 -3036 12818 -3024
rect 13778 -2448 13836 -2436
rect 13778 -3024 13790 -2448
rect 13824 -3024 13836 -2448
rect 13778 -3036 13836 -3024
rect 14796 -2448 14854 -2436
rect 14796 -3024 14808 -2448
rect 14842 -3024 14854 -2448
rect 14796 -3036 14854 -3024
rect 15814 -2448 15872 -2436
rect 15814 -3024 15826 -2448
rect 15860 -3024 15872 -2448
rect 15814 -3036 15872 -3024
rect 16832 -2448 16890 -2436
rect 16832 -3024 16844 -2448
rect 16878 -3024 16890 -2448
rect 16832 -3036 16890 -3024
rect 17850 -2448 17908 -2436
rect 17850 -3024 17862 -2448
rect 17896 -3024 17908 -2448
rect 17850 -3036 17908 -3024
rect 18868 -2448 18926 -2436
rect 18868 -3024 18880 -2448
rect 18914 -3024 18926 -2448
rect 18868 -3036 18926 -3024
rect 19886 -2448 19944 -2436
rect 19886 -3024 19898 -2448
rect 19932 -3024 19944 -2448
rect 19886 -3036 19944 -3024
rect 20904 -2448 20962 -2436
rect 20904 -3024 20916 -2448
rect 20950 -3024 20962 -2448
rect 20904 -3036 20962 -3024
rect 21922 -2448 21980 -2436
rect 21922 -3024 21934 -2448
rect 21968 -3024 21980 -2448
rect 21922 -3036 21980 -3024
rect 7670 -3480 7728 -3468
rect 7670 -4056 7682 -3480
rect 7716 -4056 7728 -3480
rect 7670 -4068 7728 -4056
rect 8688 -3480 8746 -3468
rect 8688 -4056 8700 -3480
rect 8734 -4056 8746 -3480
rect 8688 -4068 8746 -4056
rect 9706 -3480 9764 -3468
rect 9706 -4056 9718 -3480
rect 9752 -4056 9764 -3480
rect 9706 -4068 9764 -4056
rect 10724 -3480 10782 -3468
rect 10724 -4056 10736 -3480
rect 10770 -4056 10782 -3480
rect 10724 -4068 10782 -4056
rect 11742 -3480 11800 -3468
rect 11742 -4056 11754 -3480
rect 11788 -4056 11800 -3480
rect 11742 -4068 11800 -4056
rect 12760 -3480 12818 -3468
rect 12760 -4056 12772 -3480
rect 12806 -4056 12818 -3480
rect 12760 -4068 12818 -4056
rect 13778 -3480 13836 -3468
rect 13778 -4056 13790 -3480
rect 13824 -4056 13836 -3480
rect 13778 -4068 13836 -4056
rect 14796 -3480 14854 -3468
rect 14796 -4056 14808 -3480
rect 14842 -4056 14854 -3480
rect 14796 -4068 14854 -4056
rect 15814 -3480 15872 -3468
rect 15814 -4056 15826 -3480
rect 15860 -4056 15872 -3480
rect 15814 -4068 15872 -4056
rect 16832 -3480 16890 -3468
rect 16832 -4056 16844 -3480
rect 16878 -4056 16890 -3480
rect 16832 -4068 16890 -4056
rect 17850 -3480 17908 -3468
rect 17850 -4056 17862 -3480
rect 17896 -4056 17908 -3480
rect 17850 -4068 17908 -4056
rect 18868 -3480 18926 -3468
rect 18868 -4056 18880 -3480
rect 18914 -4056 18926 -3480
rect 18868 -4068 18926 -4056
rect 19886 -3480 19944 -3468
rect 19886 -4056 19898 -3480
rect 19932 -4056 19944 -3480
rect 19886 -4068 19944 -4056
rect 20904 -3480 20962 -3468
rect 20904 -4056 20916 -3480
rect 20950 -4056 20962 -3480
rect 20904 -4068 20962 -4056
rect 21922 -3480 21980 -3468
rect 21922 -4056 21934 -3480
rect 21968 -4056 21980 -3480
rect 21922 -4068 21980 -4056
rect 7462 -5084 7520 -5072
rect 2158 -5188 2216 -5176
rect 2158 -5764 2170 -5188
rect 2204 -5764 2216 -5188
rect 2158 -5776 2216 -5764
rect 3176 -5188 3234 -5176
rect 3176 -5764 3188 -5188
rect 3222 -5764 3234 -5188
rect 3176 -5776 3234 -5764
rect 4194 -5188 4252 -5176
rect 4194 -5764 4206 -5188
rect 4240 -5764 4252 -5188
rect 4194 -5776 4252 -5764
rect 5212 -5188 5270 -5176
rect 5212 -5764 5224 -5188
rect 5258 -5764 5270 -5188
rect 5212 -5776 5270 -5764
rect 6230 -5188 6288 -5176
rect 6230 -5764 6242 -5188
rect 6276 -5764 6288 -5188
rect 7462 -5660 7474 -5084
rect 7508 -5660 7520 -5084
rect 7462 -5672 7520 -5660
rect 8480 -5084 8538 -5072
rect 8480 -5660 8492 -5084
rect 8526 -5660 8538 -5084
rect 8480 -5672 8538 -5660
rect 9498 -5084 9556 -5072
rect 9498 -5660 9510 -5084
rect 9544 -5660 9556 -5084
rect 9498 -5672 9556 -5660
rect 10516 -5084 10574 -5072
rect 10516 -5660 10528 -5084
rect 10562 -5660 10574 -5084
rect 10516 -5672 10574 -5660
rect 11534 -5084 11592 -5072
rect 11534 -5660 11546 -5084
rect 11580 -5660 11592 -5084
rect 11534 -5672 11592 -5660
rect 12552 -5084 12610 -5072
rect 12552 -5660 12564 -5084
rect 12598 -5660 12610 -5084
rect 12552 -5672 12610 -5660
rect 13570 -5084 13628 -5072
rect 13570 -5660 13582 -5084
rect 13616 -5660 13628 -5084
rect 13570 -5672 13628 -5660
rect 14588 -5084 14646 -5072
rect 14588 -5660 14600 -5084
rect 14634 -5660 14646 -5084
rect 14588 -5672 14646 -5660
rect 15606 -5084 15664 -5072
rect 15606 -5660 15618 -5084
rect 15652 -5660 15664 -5084
rect 15606 -5672 15664 -5660
rect 16624 -5084 16682 -5072
rect 16624 -5660 16636 -5084
rect 16670 -5660 16682 -5084
rect 16624 -5672 16682 -5660
rect 17642 -5084 17700 -5072
rect 17642 -5660 17654 -5084
rect 17688 -5660 17700 -5084
rect 17642 -5672 17700 -5660
rect 18660 -5084 18718 -5072
rect 18660 -5660 18672 -5084
rect 18706 -5660 18718 -5084
rect 18660 -5672 18718 -5660
rect 19678 -5084 19736 -5072
rect 19678 -5660 19690 -5084
rect 19724 -5660 19736 -5084
rect 19678 -5672 19736 -5660
rect 20696 -5084 20754 -5072
rect 20696 -5660 20708 -5084
rect 20742 -5660 20754 -5084
rect 20696 -5672 20754 -5660
rect 21714 -5084 21772 -5072
rect 21714 -5660 21726 -5084
rect 21760 -5660 21772 -5084
rect 21714 -5672 21772 -5660
rect 22732 -5084 22790 -5072
rect 22732 -5660 22744 -5084
rect 22778 -5660 22790 -5084
rect 22732 -5672 22790 -5660
rect 6230 -5776 6288 -5764
rect 2158 -6220 2216 -6208
rect 2158 -6796 2170 -6220
rect 2204 -6796 2216 -6220
rect 2158 -6808 2216 -6796
rect 3176 -6220 3234 -6208
rect 3176 -6796 3188 -6220
rect 3222 -6796 3234 -6220
rect 3176 -6808 3234 -6796
rect 4194 -6220 4252 -6208
rect 4194 -6796 4206 -6220
rect 4240 -6796 4252 -6220
rect 4194 -6808 4252 -6796
rect 5212 -6220 5270 -6208
rect 5212 -6796 5224 -6220
rect 5258 -6796 5270 -6220
rect 5212 -6808 5270 -6796
rect 6230 -6220 6288 -6208
rect 6230 -6796 6242 -6220
rect 6276 -6796 6288 -6220
rect 6230 -6808 6288 -6796
rect 7462 -6340 7520 -6328
rect 7462 -6916 7474 -6340
rect 7508 -6916 7520 -6340
rect 7462 -6928 7520 -6916
rect 8480 -6340 8538 -6328
rect 8480 -6916 8492 -6340
rect 8526 -6916 8538 -6340
rect 8480 -6928 8538 -6916
rect 9498 -6340 9556 -6328
rect 9498 -6916 9510 -6340
rect 9544 -6916 9556 -6340
rect 9498 -6928 9556 -6916
rect 10516 -6340 10574 -6328
rect 10516 -6916 10528 -6340
rect 10562 -6916 10574 -6340
rect 10516 -6928 10574 -6916
rect 11534 -6340 11592 -6328
rect 11534 -6916 11546 -6340
rect 11580 -6916 11592 -6340
rect 11534 -6928 11592 -6916
rect 12552 -6340 12610 -6328
rect 12552 -6916 12564 -6340
rect 12598 -6916 12610 -6340
rect 12552 -6928 12610 -6916
rect 13570 -6340 13628 -6328
rect 13570 -6916 13582 -6340
rect 13616 -6916 13628 -6340
rect 13570 -6928 13628 -6916
rect 14588 -6340 14646 -6328
rect 14588 -6916 14600 -6340
rect 14634 -6916 14646 -6340
rect 14588 -6928 14646 -6916
rect 15606 -6340 15664 -6328
rect 15606 -6916 15618 -6340
rect 15652 -6916 15664 -6340
rect 15606 -6928 15664 -6916
rect 16624 -6340 16682 -6328
rect 16624 -6916 16636 -6340
rect 16670 -6916 16682 -6340
rect 16624 -6928 16682 -6916
rect 17642 -6340 17700 -6328
rect 17642 -6916 17654 -6340
rect 17688 -6916 17700 -6340
rect 17642 -6928 17700 -6916
rect 18660 -6340 18718 -6328
rect 18660 -6916 18672 -6340
rect 18706 -6916 18718 -6340
rect 18660 -6928 18718 -6916
rect 19678 -6340 19736 -6328
rect 19678 -6916 19690 -6340
rect 19724 -6916 19736 -6340
rect 19678 -6928 19736 -6916
rect 20696 -6340 20754 -6328
rect 20696 -6916 20708 -6340
rect 20742 -6916 20754 -6340
rect 20696 -6928 20754 -6916
rect 21714 -6340 21772 -6328
rect 21714 -6916 21726 -6340
rect 21760 -6916 21772 -6340
rect 21714 -6928 21772 -6916
rect 22732 -6340 22790 -6328
rect 22732 -6916 22744 -6340
rect 22778 -6916 22790 -6340
rect 22732 -6928 22790 -6916
rect 2158 -7252 2216 -7240
rect 2158 -7828 2170 -7252
rect 2204 -7828 2216 -7252
rect 2158 -7840 2216 -7828
rect 3176 -7252 3234 -7240
rect 3176 -7828 3188 -7252
rect 3222 -7828 3234 -7252
rect 3176 -7840 3234 -7828
rect 4194 -7252 4252 -7240
rect 4194 -7828 4206 -7252
rect 4240 -7828 4252 -7252
rect 4194 -7840 4252 -7828
rect 5212 -7252 5270 -7240
rect 5212 -7828 5224 -7252
rect 5258 -7828 5270 -7252
rect 5212 -7840 5270 -7828
rect 6230 -7252 6288 -7240
rect 6230 -7828 6242 -7252
rect 6276 -7828 6288 -7252
rect 6230 -7840 6288 -7828
rect 7462 -7596 7520 -7584
rect 7462 -8172 7474 -7596
rect 7508 -8172 7520 -7596
rect 7462 -8184 7520 -8172
rect 8480 -7596 8538 -7584
rect 8480 -8172 8492 -7596
rect 8526 -8172 8538 -7596
rect 8480 -8184 8538 -8172
rect 9498 -7596 9556 -7584
rect 9498 -8172 9510 -7596
rect 9544 -8172 9556 -7596
rect 9498 -8184 9556 -8172
rect 10516 -7596 10574 -7584
rect 10516 -8172 10528 -7596
rect 10562 -8172 10574 -7596
rect 10516 -8184 10574 -8172
rect 11534 -7596 11592 -7584
rect 11534 -8172 11546 -7596
rect 11580 -8172 11592 -7596
rect 11534 -8184 11592 -8172
rect 12552 -7596 12610 -7584
rect 12552 -8172 12564 -7596
rect 12598 -8172 12610 -7596
rect 12552 -8184 12610 -8172
rect 13570 -7596 13628 -7584
rect 13570 -8172 13582 -7596
rect 13616 -8172 13628 -7596
rect 13570 -8184 13628 -8172
rect 14588 -7596 14646 -7584
rect 14588 -8172 14600 -7596
rect 14634 -8172 14646 -7596
rect 14588 -8184 14646 -8172
rect 15606 -7596 15664 -7584
rect 15606 -8172 15618 -7596
rect 15652 -8172 15664 -7596
rect 15606 -8184 15664 -8172
rect 16624 -7596 16682 -7584
rect 16624 -8172 16636 -7596
rect 16670 -8172 16682 -7596
rect 16624 -8184 16682 -8172
rect 17642 -7596 17700 -7584
rect 17642 -8172 17654 -7596
rect 17688 -8172 17700 -7596
rect 17642 -8184 17700 -8172
rect 18660 -7596 18718 -7584
rect 18660 -8172 18672 -7596
rect 18706 -8172 18718 -7596
rect 18660 -8184 18718 -8172
rect 19678 -7596 19736 -7584
rect 19678 -8172 19690 -7596
rect 19724 -8172 19736 -7596
rect 19678 -8184 19736 -8172
rect 20696 -7596 20754 -7584
rect 20696 -8172 20708 -7596
rect 20742 -8172 20754 -7596
rect 20696 -8184 20754 -8172
rect 21714 -7596 21772 -7584
rect 21714 -8172 21726 -7596
rect 21760 -8172 21772 -7596
rect 21714 -8184 21772 -8172
rect 22732 -7596 22790 -7584
rect 22732 -8172 22744 -7596
rect 22778 -8172 22790 -7596
rect 22732 -8184 22790 -8172
rect 2158 -8284 2216 -8272
rect 2158 -8860 2170 -8284
rect 2204 -8860 2216 -8284
rect 2158 -8872 2216 -8860
rect 3176 -8284 3234 -8272
rect 3176 -8860 3188 -8284
rect 3222 -8860 3234 -8284
rect 3176 -8872 3234 -8860
rect 4194 -8284 4252 -8272
rect 4194 -8860 4206 -8284
rect 4240 -8860 4252 -8284
rect 4194 -8872 4252 -8860
rect 5212 -8284 5270 -8272
rect 5212 -8860 5224 -8284
rect 5258 -8860 5270 -8284
rect 5212 -8872 5270 -8860
rect 6230 -8284 6288 -8272
rect 6230 -8860 6242 -8284
rect 6276 -8860 6288 -8284
rect 6230 -8872 6288 -8860
rect 7462 -8852 7520 -8840
rect 7462 -9428 7474 -8852
rect 7508 -9428 7520 -8852
rect 7462 -9440 7520 -9428
rect 8480 -8852 8538 -8840
rect 8480 -9428 8492 -8852
rect 8526 -9428 8538 -8852
rect 8480 -9440 8538 -9428
rect 9498 -8852 9556 -8840
rect 9498 -9428 9510 -8852
rect 9544 -9428 9556 -8852
rect 9498 -9440 9556 -9428
rect 10516 -8852 10574 -8840
rect 10516 -9428 10528 -8852
rect 10562 -9428 10574 -8852
rect 10516 -9440 10574 -9428
rect 11534 -8852 11592 -8840
rect 11534 -9428 11546 -8852
rect 11580 -9428 11592 -8852
rect 11534 -9440 11592 -9428
rect 12552 -8852 12610 -8840
rect 12552 -9428 12564 -8852
rect 12598 -9428 12610 -8852
rect 12552 -9440 12610 -9428
rect 13570 -8852 13628 -8840
rect 13570 -9428 13582 -8852
rect 13616 -9428 13628 -8852
rect 13570 -9440 13628 -9428
rect 14588 -8852 14646 -8840
rect 14588 -9428 14600 -8852
rect 14634 -9428 14646 -8852
rect 14588 -9440 14646 -9428
rect 15606 -8852 15664 -8840
rect 15606 -9428 15618 -8852
rect 15652 -9428 15664 -8852
rect 15606 -9440 15664 -9428
rect 16624 -8852 16682 -8840
rect 16624 -9428 16636 -8852
rect 16670 -9428 16682 -8852
rect 16624 -9440 16682 -9428
rect 17642 -8852 17700 -8840
rect 17642 -9428 17654 -8852
rect 17688 -9428 17700 -8852
rect 17642 -9440 17700 -9428
rect 18660 -8852 18718 -8840
rect 18660 -9428 18672 -8852
rect 18706 -9428 18718 -8852
rect 18660 -9440 18718 -9428
rect 19678 -8852 19736 -8840
rect 19678 -9428 19690 -8852
rect 19724 -9428 19736 -8852
rect 19678 -9440 19736 -9428
rect 20696 -8852 20754 -8840
rect 20696 -9428 20708 -8852
rect 20742 -9428 20754 -8852
rect 20696 -9440 20754 -9428
rect 21714 -8852 21772 -8840
rect 21714 -9428 21726 -8852
rect 21760 -9428 21772 -8852
rect 21714 -9440 21772 -9428
rect 22732 -8852 22790 -8840
rect 22732 -9428 22744 -8852
rect 22778 -9428 22790 -8852
rect 22732 -9440 22790 -9428
<< ndiffc >>
rect -9184 -13100 -9150 -12524
rect -8166 -13100 -8132 -12524
rect -7148 -13100 -7114 -12524
rect -6130 -13100 -6096 -12524
rect -5112 -13100 -5078 -12524
rect -4094 -13100 -4060 -12524
rect -3076 -13100 -3042 -12524
rect -2058 -13100 -2024 -12524
rect -1040 -13100 -1006 -12524
rect -22 -13100 12 -12524
rect 2582 -12624 2616 -12048
rect 3600 -12624 3634 -12048
rect 4618 -12624 4652 -12048
rect 5636 -12624 5670 -12048
rect 6654 -12624 6688 -12048
rect 7672 -12624 7706 -12048
rect 8690 -12624 8724 -12048
rect 9708 -12624 9742 -12048
rect 10726 -12624 10760 -12048
rect 11744 -12624 11778 -12048
rect 12762 -12624 12796 -12048
rect 13780 -12624 13814 -12048
rect 14798 -12624 14832 -12048
rect 15816 -12624 15850 -12048
rect 16834 -12624 16868 -12048
rect 17852 -12624 17886 -12048
rect 18870 -12624 18904 -12048
rect 19888 -12624 19922 -12048
rect 20906 -12624 20940 -12048
rect 21924 -12624 21958 -12048
rect 22942 -12624 22976 -12048
rect -9184 -13918 -9150 -13342
rect -8166 -13918 -8132 -13342
rect -7148 -13918 -7114 -13342
rect -6130 -13918 -6096 -13342
rect -5112 -13918 -5078 -13342
rect -4094 -13918 -4060 -13342
rect -3076 -13918 -3042 -13342
rect -2058 -13918 -2024 -13342
rect -1040 -13918 -1006 -13342
rect -22 -13918 12 -13342
rect 2582 -13442 2616 -12866
rect 3600 -13442 3634 -12866
rect 4618 -13442 4652 -12866
rect 5636 -13442 5670 -12866
rect 6654 -13442 6688 -12866
rect 7672 -13442 7706 -12866
rect 8690 -13442 8724 -12866
rect 9708 -13442 9742 -12866
rect 10726 -13442 10760 -12866
rect 11744 -13442 11778 -12866
rect 12762 -13442 12796 -12866
rect 13780 -13442 13814 -12866
rect 14798 -13442 14832 -12866
rect 15816 -13442 15850 -12866
rect 16834 -13442 16868 -12866
rect 17852 -13442 17886 -12866
rect 18870 -13442 18904 -12866
rect 19888 -13442 19922 -12866
rect 20906 -13442 20940 -12866
rect 21924 -13442 21958 -12866
rect 22942 -13442 22976 -12866
rect -9184 -14736 -9150 -14160
rect -8166 -14736 -8132 -14160
rect -7148 -14736 -7114 -14160
rect -6130 -14736 -6096 -14160
rect -5112 -14736 -5078 -14160
rect -4094 -14736 -4060 -14160
rect -3076 -14736 -3042 -14160
rect -2058 -14736 -2024 -14160
rect -1040 -14736 -1006 -14160
rect -22 -14736 12 -14160
rect 2582 -14820 2616 -14244
rect 3600 -14820 3634 -14244
rect 4618 -14820 4652 -14244
rect 5636 -14820 5670 -14244
rect 6654 -14820 6688 -14244
rect 7672 -14820 7706 -14244
rect 8690 -14820 8724 -14244
rect 9708 -14820 9742 -14244
rect 10726 -14820 10760 -14244
rect 11744 -14820 11778 -14244
rect 12762 -14820 12796 -14244
rect 13780 -14820 13814 -14244
rect 14798 -14820 14832 -14244
rect 15816 -14820 15850 -14244
rect 16834 -14820 16868 -14244
rect 17852 -14820 17886 -14244
rect 18870 -14820 18904 -14244
rect 19888 -14820 19922 -14244
rect 20906 -14820 20940 -14244
rect 21924 -14820 21958 -14244
rect 22942 -14820 22976 -14244
rect -9184 -15554 -9150 -14978
rect -8166 -15554 -8132 -14978
rect -7148 -15554 -7114 -14978
rect -6130 -15554 -6096 -14978
rect -5112 -15554 -5078 -14978
rect -4094 -15554 -4060 -14978
rect -3076 -15554 -3042 -14978
rect -2058 -15554 -2024 -14978
rect -1040 -15554 -1006 -14978
rect -22 -15554 12 -14978
rect -9184 -16372 -9150 -15796
rect -8166 -16372 -8132 -15796
rect -7148 -16372 -7114 -15796
rect -6130 -16372 -6096 -15796
rect -5112 -16372 -5078 -15796
rect -4094 -16372 -4060 -15796
rect -3076 -16372 -3042 -15796
rect -2058 -16372 -2024 -15796
rect -1040 -16372 -1006 -15796
rect -22 -16372 12 -15796
rect 2582 -16052 2616 -15476
rect 3600 -16052 3634 -15476
rect 4618 -16052 4652 -15476
rect 5636 -16052 5670 -15476
rect 6654 -16052 6688 -15476
rect 7672 -16052 7706 -15476
rect 8690 -16052 8724 -15476
rect 9708 -16052 9742 -15476
rect 10726 -16052 10760 -15476
rect 11744 -16052 11778 -15476
rect 12762 -16052 12796 -15476
rect 13780 -16052 13814 -15476
rect 14798 -16052 14832 -15476
rect 15816 -16052 15850 -15476
rect 16834 -16052 16868 -15476
rect 17852 -16052 17886 -15476
rect 18870 -16052 18904 -15476
rect 19888 -16052 19922 -15476
rect 20906 -16052 20940 -15476
rect 21924 -16052 21958 -15476
rect 22942 -16052 22976 -15476
rect -9184 -17190 -9150 -16614
rect -8166 -17190 -8132 -16614
rect -7148 -17190 -7114 -16614
rect -6130 -17190 -6096 -16614
rect -5112 -17190 -5078 -16614
rect -4094 -17190 -4060 -16614
rect -3076 -17190 -3042 -16614
rect -2058 -17190 -2024 -16614
rect -1040 -17190 -1006 -16614
rect -22 -17190 12 -16614
rect 2580 -17286 2614 -16710
rect 3598 -17286 3632 -16710
rect 4616 -17286 4650 -16710
rect 5634 -17286 5668 -16710
rect 6652 -17286 6686 -16710
rect 7670 -17286 7704 -16710
rect 8688 -17286 8722 -16710
rect 9706 -17286 9740 -16710
rect 10724 -17286 10758 -16710
rect 11742 -17286 11776 -16710
rect 12760 -17286 12794 -16710
rect 13778 -17286 13812 -16710
rect 14796 -17286 14830 -16710
rect 15814 -17286 15848 -16710
rect 16832 -17286 16866 -16710
rect 17850 -17286 17884 -16710
rect 18868 -17286 18902 -16710
rect 19886 -17286 19920 -16710
rect 20904 -17286 20938 -16710
rect 21922 -17286 21956 -16710
rect 22940 -17286 22974 -16710
rect -9184 -18008 -9150 -17432
rect -8166 -18008 -8132 -17432
rect -7148 -18008 -7114 -17432
rect -6130 -18008 -6096 -17432
rect -5112 -18008 -5078 -17432
rect -4094 -18008 -4060 -17432
rect -3076 -18008 -3042 -17432
rect -2058 -18008 -2024 -17432
rect -1040 -18008 -1006 -17432
rect -22 -18008 12 -17432
rect -9184 -18826 -9150 -18250
rect -8166 -18826 -8132 -18250
rect -7148 -18826 -7114 -18250
rect -6130 -18826 -6096 -18250
rect -5112 -18826 -5078 -18250
rect -4094 -18826 -4060 -18250
rect -3076 -18826 -3042 -18250
rect -2058 -18826 -2024 -18250
rect -1040 -18826 -1006 -18250
rect -22 -18826 12 -18250
rect 2580 -18520 2614 -17944
rect 3598 -18520 3632 -17944
rect 4616 -18520 4650 -17944
rect 5634 -18520 5668 -17944
rect 6652 -18520 6686 -17944
rect 7670 -18520 7704 -17944
rect 8688 -18520 8722 -17944
rect 9706 -18520 9740 -17944
rect 10724 -18520 10758 -17944
rect 11742 -18520 11776 -17944
rect 12760 -18520 12794 -17944
rect 13778 -18520 13812 -17944
rect 14796 -18520 14830 -17944
rect 15814 -18520 15848 -17944
rect 16832 -18520 16866 -17944
rect 17850 -18520 17884 -17944
rect 18868 -18520 18902 -17944
rect 19886 -18520 19920 -17944
rect 20904 -18520 20938 -17944
rect 21922 -18520 21956 -17944
rect 22940 -18520 22974 -17944
rect 2580 -19752 2614 -19176
rect 3598 -19752 3632 -19176
rect 4616 -19752 4650 -19176
rect 5634 -19752 5668 -19176
rect 6652 -19752 6686 -19176
rect 7670 -19752 7704 -19176
rect 8688 -19752 8722 -19176
rect 9706 -19752 9740 -19176
rect 10724 -19752 10758 -19176
rect 11742 -19752 11776 -19176
rect 12760 -19752 12794 -19176
rect 13778 -19752 13812 -19176
rect 14796 -19752 14830 -19176
rect 15814 -19752 15848 -19176
rect 16832 -19752 16866 -19176
rect 17850 -19752 17884 -19176
rect 18868 -19752 18902 -19176
rect 19886 -19752 19920 -19176
rect 20904 -19752 20938 -19176
rect 21922 -19752 21956 -19176
rect 22940 -19752 22974 -19176
rect -10508 -20850 -10474 -20274
rect -9490 -20850 -9456 -20274
rect -8472 -20850 -8438 -20274
rect -7454 -20850 -7420 -20274
rect -6436 -20850 -6402 -20274
rect -5418 -20850 -5384 -20274
rect -4400 -20850 -4366 -20274
rect -3382 -20850 -3348 -20274
rect -2364 -20850 -2330 -20274
rect -1346 -20850 -1312 -20274
rect -328 -20850 -294 -20274
rect 690 -20850 724 -20274
rect 2580 -20986 2614 -20410
rect 3598 -20986 3632 -20410
rect 4616 -20986 4650 -20410
rect 5634 -20986 5668 -20410
rect 6652 -20986 6686 -20410
rect 7670 -20986 7704 -20410
rect 8688 -20986 8722 -20410
rect 9706 -20986 9740 -20410
rect 10724 -20986 10758 -20410
rect 11742 -20986 11776 -20410
rect 12760 -20986 12794 -20410
rect 13778 -20986 13812 -20410
rect 14796 -20986 14830 -20410
rect 15814 -20986 15848 -20410
rect 16832 -20986 16866 -20410
rect 17850 -20986 17884 -20410
rect 18868 -20986 18902 -20410
rect 19886 -20986 19920 -20410
rect 20904 -20986 20938 -20410
rect 21922 -20986 21956 -20410
rect 22940 -20986 22974 -20410
rect -10508 -21962 -10474 -21386
rect -9490 -21962 -9456 -21386
rect -8472 -21962 -8438 -21386
rect -7454 -21962 -7420 -21386
rect -6436 -21962 -6402 -21386
rect -5418 -21962 -5384 -21386
rect -4400 -21962 -4366 -21386
rect -3382 -21962 -3348 -21386
rect -2364 -21962 -2330 -21386
rect -1346 -21962 -1312 -21386
rect -328 -21962 -294 -21386
rect 690 -21962 724 -21386
rect 2580 -22220 2614 -21644
rect 3598 -22220 3632 -21644
rect 4616 -22220 4650 -21644
rect 5634 -22220 5668 -21644
rect 6652 -22220 6686 -21644
rect 7670 -22220 7704 -21644
rect 8688 -22220 8722 -21644
rect 9706 -22220 9740 -21644
rect 10724 -22220 10758 -21644
rect 11742 -22220 11776 -21644
rect 12760 -22220 12794 -21644
rect 13778 -22220 13812 -21644
rect 14796 -22220 14830 -21644
rect 15814 -22220 15848 -21644
rect 16832 -22220 16866 -21644
rect 17850 -22220 17884 -21644
rect 18868 -22220 18902 -21644
rect 19886 -22220 19920 -21644
rect 20904 -22220 20938 -21644
rect 21922 -22220 21956 -21644
rect 22940 -22220 22974 -21644
rect -10508 -23074 -10474 -22498
rect -9490 -23074 -9456 -22498
rect -8472 -23074 -8438 -22498
rect -7454 -23074 -7420 -22498
rect -6436 -23074 -6402 -22498
rect -5418 -23074 -5384 -22498
rect -4400 -23074 -4366 -22498
rect -3382 -23074 -3348 -22498
rect -2364 -23074 -2330 -22498
rect -1346 -23074 -1312 -22498
rect -328 -23074 -294 -22498
rect 690 -23074 724 -22498
rect 2580 -23452 2614 -22876
rect 3598 -23452 3632 -22876
rect 4616 -23452 4650 -22876
rect 5634 -23452 5668 -22876
rect 6652 -23452 6686 -22876
rect 7670 -23452 7704 -22876
rect 8688 -23452 8722 -22876
rect 9706 -23452 9740 -22876
rect 10724 -23452 10758 -22876
rect 11742 -23452 11776 -22876
rect 12760 -23452 12794 -22876
rect 13778 -23452 13812 -22876
rect 14796 -23452 14830 -22876
rect 15814 -23452 15848 -22876
rect 16832 -23452 16866 -22876
rect 17850 -23452 17884 -22876
rect 18868 -23452 18902 -22876
rect 19886 -23452 19920 -22876
rect 20904 -23452 20938 -22876
rect 21922 -23452 21956 -22876
rect 22940 -23452 22974 -22876
rect -10508 -24186 -10474 -23610
rect -9490 -24186 -9456 -23610
rect -8472 -24186 -8438 -23610
rect -7454 -24186 -7420 -23610
rect -6436 -24186 -6402 -23610
rect -5418 -24186 -5384 -23610
rect -4400 -24186 -4366 -23610
rect -3382 -24186 -3348 -23610
rect -2364 -24186 -2330 -23610
rect -1346 -24186 -1312 -23610
rect -328 -24186 -294 -23610
rect 690 -24186 724 -23610
rect 2580 -24686 2614 -24110
rect 3598 -24686 3632 -24110
rect 4616 -24686 4650 -24110
rect 5634 -24686 5668 -24110
rect 6652 -24686 6686 -24110
rect 7670 -24686 7704 -24110
rect 8688 -24686 8722 -24110
rect 9706 -24686 9740 -24110
rect 10724 -24686 10758 -24110
rect 11742 -24686 11776 -24110
rect 12760 -24686 12794 -24110
rect 13778 -24686 13812 -24110
rect 14796 -24686 14830 -24110
rect 15814 -24686 15848 -24110
rect 16832 -24686 16866 -24110
rect 17850 -24686 17884 -24110
rect 18868 -24686 18902 -24110
rect 19886 -24686 19920 -24110
rect 20904 -24686 20938 -24110
rect 21922 -24686 21956 -24110
rect 22940 -24686 22974 -24110
rect -10050 -25728 -10016 -25152
rect -9032 -25728 -8998 -25152
rect -8014 -25728 -7980 -25152
rect -6996 -25728 -6962 -25152
rect -5978 -25728 -5944 -25152
rect -4960 -25728 -4926 -25152
rect -3942 -25728 -3908 -25152
rect -2924 -25728 -2890 -25152
rect -1906 -25728 -1872 -25152
rect -888 -25728 -854 -25152
rect 130 -25728 164 -25152
rect 2580 -25918 2614 -25342
rect 3598 -25918 3632 -25342
rect 4616 -25918 4650 -25342
rect 5634 -25918 5668 -25342
rect 6652 -25918 6686 -25342
rect 7670 -25918 7704 -25342
rect 8688 -25918 8722 -25342
rect 9706 -25918 9740 -25342
rect 10724 -25918 10758 -25342
rect 11742 -25918 11776 -25342
rect 12760 -25918 12794 -25342
rect 13778 -25918 13812 -25342
rect 14796 -25918 14830 -25342
rect 15814 -25918 15848 -25342
rect 16832 -25918 16866 -25342
rect 17850 -25918 17884 -25342
rect 18868 -25918 18902 -25342
rect 19886 -25918 19920 -25342
rect 20904 -25918 20938 -25342
rect 21922 -25918 21956 -25342
rect 22940 -25918 22974 -25342
<< pdiffc >>
rect 6488 886 6522 1462
rect 7506 886 7540 1462
rect 8524 886 8558 1462
rect 9542 886 9576 1462
rect 10560 886 10594 1462
rect 11578 886 11612 1462
rect 12596 886 12630 1462
rect 13614 886 13648 1462
rect 14632 886 14666 1462
rect 15650 886 15684 1462
rect 16668 886 16702 1462
rect 17686 886 17720 1462
rect 18704 886 18738 1462
rect 19722 886 19756 1462
rect 20740 886 20774 1462
rect 21758 886 21792 1462
rect 22776 886 22810 1462
rect 6488 -250 6522 326
rect 7506 -250 7540 326
rect 8524 -250 8558 326
rect 9542 -250 9576 326
rect 10560 -250 10594 326
rect 11578 -250 11612 326
rect 12596 -250 12630 326
rect 13614 -250 13648 326
rect 14632 -250 14666 326
rect 15650 -250 15684 326
rect 16668 -250 16702 326
rect 17686 -250 17720 326
rect 18704 -250 18738 326
rect 19722 -250 19756 326
rect 20740 -250 20774 326
rect 21758 -250 21792 326
rect 22776 -250 22810 326
rect 6488 -1386 6522 -810
rect 7506 -1386 7540 -810
rect 8524 -1386 8558 -810
rect 9542 -1386 9576 -810
rect 10560 -1386 10594 -810
rect 11578 -1386 11612 -810
rect 12596 -1386 12630 -810
rect 13614 -1386 13648 -810
rect 14632 -1386 14666 -810
rect 15650 -1386 15684 -810
rect 16668 -1386 16702 -810
rect 17686 -1386 17720 -810
rect 18704 -1386 18738 -810
rect 19722 -1386 19756 -810
rect 20740 -1386 20774 -810
rect 21758 -1386 21792 -810
rect 22776 -1386 22810 -810
rect 7682 -3024 7716 -2448
rect 8700 -3024 8734 -2448
rect 9718 -3024 9752 -2448
rect 10736 -3024 10770 -2448
rect 11754 -3024 11788 -2448
rect 12772 -3024 12806 -2448
rect 13790 -3024 13824 -2448
rect 14808 -3024 14842 -2448
rect 15826 -3024 15860 -2448
rect 16844 -3024 16878 -2448
rect 17862 -3024 17896 -2448
rect 18880 -3024 18914 -2448
rect 19898 -3024 19932 -2448
rect 20916 -3024 20950 -2448
rect 21934 -3024 21968 -2448
rect 7682 -4056 7716 -3480
rect 8700 -4056 8734 -3480
rect 9718 -4056 9752 -3480
rect 10736 -4056 10770 -3480
rect 11754 -4056 11788 -3480
rect 12772 -4056 12806 -3480
rect 13790 -4056 13824 -3480
rect 14808 -4056 14842 -3480
rect 15826 -4056 15860 -3480
rect 16844 -4056 16878 -3480
rect 17862 -4056 17896 -3480
rect 18880 -4056 18914 -3480
rect 19898 -4056 19932 -3480
rect 20916 -4056 20950 -3480
rect 21934 -4056 21968 -3480
rect 2170 -5764 2204 -5188
rect 3188 -5764 3222 -5188
rect 4206 -5764 4240 -5188
rect 5224 -5764 5258 -5188
rect 6242 -5764 6276 -5188
rect 7474 -5660 7508 -5084
rect 8492 -5660 8526 -5084
rect 9510 -5660 9544 -5084
rect 10528 -5660 10562 -5084
rect 11546 -5660 11580 -5084
rect 12564 -5660 12598 -5084
rect 13582 -5660 13616 -5084
rect 14600 -5660 14634 -5084
rect 15618 -5660 15652 -5084
rect 16636 -5660 16670 -5084
rect 17654 -5660 17688 -5084
rect 18672 -5660 18706 -5084
rect 19690 -5660 19724 -5084
rect 20708 -5660 20742 -5084
rect 21726 -5660 21760 -5084
rect 22744 -5660 22778 -5084
rect 2170 -6796 2204 -6220
rect 3188 -6796 3222 -6220
rect 4206 -6796 4240 -6220
rect 5224 -6796 5258 -6220
rect 6242 -6796 6276 -6220
rect 7474 -6916 7508 -6340
rect 8492 -6916 8526 -6340
rect 9510 -6916 9544 -6340
rect 10528 -6916 10562 -6340
rect 11546 -6916 11580 -6340
rect 12564 -6916 12598 -6340
rect 13582 -6916 13616 -6340
rect 14600 -6916 14634 -6340
rect 15618 -6916 15652 -6340
rect 16636 -6916 16670 -6340
rect 17654 -6916 17688 -6340
rect 18672 -6916 18706 -6340
rect 19690 -6916 19724 -6340
rect 20708 -6916 20742 -6340
rect 21726 -6916 21760 -6340
rect 22744 -6916 22778 -6340
rect 2170 -7828 2204 -7252
rect 3188 -7828 3222 -7252
rect 4206 -7828 4240 -7252
rect 5224 -7828 5258 -7252
rect 6242 -7828 6276 -7252
rect 7474 -8172 7508 -7596
rect 8492 -8172 8526 -7596
rect 9510 -8172 9544 -7596
rect 10528 -8172 10562 -7596
rect 11546 -8172 11580 -7596
rect 12564 -8172 12598 -7596
rect 13582 -8172 13616 -7596
rect 14600 -8172 14634 -7596
rect 15618 -8172 15652 -7596
rect 16636 -8172 16670 -7596
rect 17654 -8172 17688 -7596
rect 18672 -8172 18706 -7596
rect 19690 -8172 19724 -7596
rect 20708 -8172 20742 -7596
rect 21726 -8172 21760 -7596
rect 22744 -8172 22778 -7596
rect 2170 -8860 2204 -8284
rect 3188 -8860 3222 -8284
rect 4206 -8860 4240 -8284
rect 5224 -8860 5258 -8284
rect 6242 -8860 6276 -8284
rect 7474 -9428 7508 -8852
rect 8492 -9428 8526 -8852
rect 9510 -9428 9544 -8852
rect 10528 -9428 10562 -8852
rect 11546 -9428 11580 -8852
rect 12564 -9428 12598 -8852
rect 13582 -9428 13616 -8852
rect 14600 -9428 14634 -8852
rect 15618 -9428 15652 -8852
rect 16636 -9428 16670 -8852
rect 17654 -9428 17688 -8852
rect 18672 -9428 18706 -8852
rect 19690 -9428 19724 -8852
rect 20708 -9428 20742 -8852
rect 21726 -9428 21760 -8852
rect 22744 -9428 22778 -8852
<< psubdiff >>
rect -12322 -11278 -12160 -11178
rect 24760 -11278 24922 -11178
rect -12322 -11340 -12222 -11278
rect 24822 -11340 24922 -11278
rect 3086 -11784 3168 -11760
rect 3086 -11818 3110 -11784
rect 3144 -11818 3168 -11784
rect 3086 -11842 3168 -11818
rect 4104 -11784 4186 -11760
rect 4104 -11818 4128 -11784
rect 4162 -11818 4186 -11784
rect 4104 -11842 4186 -11818
rect 5122 -11784 5204 -11760
rect 5122 -11818 5146 -11784
rect 5180 -11818 5204 -11784
rect 5122 -11842 5204 -11818
rect 6140 -11784 6222 -11760
rect 6140 -11818 6164 -11784
rect 6198 -11818 6222 -11784
rect 6140 -11842 6222 -11818
rect 7158 -11784 7240 -11760
rect 7158 -11818 7182 -11784
rect 7216 -11818 7240 -11784
rect 7158 -11842 7240 -11818
rect 8176 -11784 8258 -11760
rect 8176 -11818 8200 -11784
rect 8234 -11818 8258 -11784
rect 8176 -11842 8258 -11818
rect 9194 -11784 9276 -11760
rect 9194 -11818 9218 -11784
rect 9252 -11818 9276 -11784
rect 9194 -11842 9276 -11818
rect 10212 -11784 10294 -11760
rect 10212 -11818 10236 -11784
rect 10270 -11818 10294 -11784
rect 10212 -11842 10294 -11818
rect 11230 -11784 11312 -11760
rect 11230 -11818 11254 -11784
rect 11288 -11818 11312 -11784
rect 11230 -11842 11312 -11818
rect 12248 -11784 12330 -11760
rect 12248 -11818 12272 -11784
rect 12306 -11818 12330 -11784
rect 12248 -11842 12330 -11818
rect 13266 -11784 13348 -11760
rect 13266 -11818 13290 -11784
rect 13324 -11818 13348 -11784
rect 13266 -11842 13348 -11818
rect 14284 -11784 14366 -11760
rect 14284 -11818 14308 -11784
rect 14342 -11818 14366 -11784
rect 14284 -11842 14366 -11818
rect 15302 -11784 15384 -11760
rect 15302 -11818 15326 -11784
rect 15360 -11818 15384 -11784
rect 15302 -11842 15384 -11818
rect 16320 -11784 16402 -11760
rect 16320 -11818 16344 -11784
rect 16378 -11818 16402 -11784
rect 16320 -11842 16402 -11818
rect 17338 -11784 17420 -11760
rect 17338 -11818 17362 -11784
rect 17396 -11818 17420 -11784
rect 17338 -11842 17420 -11818
rect 18356 -11784 18438 -11760
rect 18356 -11818 18380 -11784
rect 18414 -11818 18438 -11784
rect 18356 -11842 18438 -11818
rect 19374 -11784 19456 -11760
rect 19374 -11818 19398 -11784
rect 19432 -11818 19456 -11784
rect 19374 -11842 19456 -11818
rect 20392 -11784 20474 -11760
rect 20392 -11818 20416 -11784
rect 20450 -11818 20474 -11784
rect 20392 -11842 20474 -11818
rect 21410 -11784 21492 -11760
rect 21410 -11818 21434 -11784
rect 21468 -11818 21492 -11784
rect 21410 -11842 21492 -11818
rect 22428 -11784 22510 -11760
rect 22428 -11818 22452 -11784
rect 22486 -11818 22510 -11784
rect 22428 -11842 22510 -11818
rect -9208 -12386 -9126 -12362
rect -9208 -12420 -9184 -12386
rect -9150 -12420 -9126 -12386
rect -9208 -12444 -9126 -12420
rect -8190 -12386 -8108 -12362
rect -8190 -12420 -8166 -12386
rect -8132 -12420 -8108 -12386
rect -8190 -12444 -8108 -12420
rect -7172 -12386 -7090 -12362
rect -7172 -12420 -7148 -12386
rect -7114 -12420 -7090 -12386
rect -7172 -12444 -7090 -12420
rect -6154 -12386 -6072 -12362
rect -6154 -12420 -6130 -12386
rect -6096 -12420 -6072 -12386
rect -6154 -12444 -6072 -12420
rect -5136 -12386 -5054 -12362
rect -5136 -12420 -5112 -12386
rect -5078 -12420 -5054 -12386
rect -5136 -12444 -5054 -12420
rect -4118 -12386 -4036 -12362
rect -4118 -12420 -4094 -12386
rect -4060 -12420 -4036 -12386
rect -4118 -12444 -4036 -12420
rect -3100 -12386 -3018 -12362
rect -3100 -12420 -3076 -12386
rect -3042 -12420 -3018 -12386
rect -3100 -12444 -3018 -12420
rect -2082 -12386 -2000 -12362
rect -2082 -12420 -2058 -12386
rect -2024 -12420 -2000 -12386
rect -2082 -12444 -2000 -12420
rect -1064 -12386 -982 -12362
rect -1064 -12420 -1040 -12386
rect -1006 -12420 -982 -12386
rect -1064 -12444 -982 -12420
rect -36 -12386 46 -12362
rect -36 -12420 -12 -12386
rect 22 -12420 46 -12386
rect -36 -12444 46 -12420
rect -9208 -13204 -9126 -13180
rect -9208 -13238 -9184 -13204
rect -9150 -13238 -9126 -13204
rect -9208 -13262 -9126 -13238
rect -8190 -13204 -8108 -13180
rect -8190 -13238 -8166 -13204
rect -8132 -13238 -8108 -13204
rect -8190 -13262 -8108 -13238
rect -7172 -13204 -7090 -13180
rect -7172 -13238 -7148 -13204
rect -7114 -13238 -7090 -13204
rect -7172 -13262 -7090 -13238
rect -6154 -13204 -6072 -13180
rect -6154 -13238 -6130 -13204
rect -6096 -13238 -6072 -13204
rect -6154 -13262 -6072 -13238
rect -5136 -13204 -5054 -13180
rect -5136 -13238 -5112 -13204
rect -5078 -13238 -5054 -13204
rect -5136 -13262 -5054 -13238
rect -4118 -13204 -4036 -13180
rect -4118 -13238 -4094 -13204
rect -4060 -13238 -4036 -13204
rect -4118 -13262 -4036 -13238
rect -3100 -13204 -3018 -13180
rect -3100 -13238 -3076 -13204
rect -3042 -13238 -3018 -13204
rect -3100 -13262 -3018 -13238
rect -2082 -13204 -2000 -13180
rect -2082 -13238 -2058 -13204
rect -2024 -13238 -2000 -13204
rect -2082 -13262 -2000 -13238
rect -1064 -13204 -982 -13180
rect -1064 -13238 -1040 -13204
rect -1006 -13238 -982 -13204
rect -1064 -13262 -982 -13238
rect -36 -13204 46 -13180
rect -36 -13238 -12 -13204
rect 22 -13238 46 -13204
rect -36 -13262 46 -13238
rect 3098 -13810 3180 -13786
rect 3098 -13844 3122 -13810
rect 3156 -13844 3180 -13810
rect 3098 -13868 3180 -13844
rect 4116 -13810 4198 -13786
rect 4116 -13844 4140 -13810
rect 4174 -13844 4198 -13810
rect 4116 -13868 4198 -13844
rect 5134 -13810 5216 -13786
rect 5134 -13844 5158 -13810
rect 5192 -13844 5216 -13810
rect 5134 -13868 5216 -13844
rect 6152 -13810 6234 -13786
rect 6152 -13844 6176 -13810
rect 6210 -13844 6234 -13810
rect 6152 -13868 6234 -13844
rect 7170 -13810 7252 -13786
rect 7170 -13844 7194 -13810
rect 7228 -13844 7252 -13810
rect 7170 -13868 7252 -13844
rect 8188 -13810 8270 -13786
rect 8188 -13844 8212 -13810
rect 8246 -13844 8270 -13810
rect 8188 -13868 8270 -13844
rect 9206 -13810 9288 -13786
rect 9206 -13844 9230 -13810
rect 9264 -13844 9288 -13810
rect 9206 -13868 9288 -13844
rect 10224 -13810 10306 -13786
rect 10224 -13844 10248 -13810
rect 10282 -13844 10306 -13810
rect 10224 -13868 10306 -13844
rect 11242 -13810 11324 -13786
rect 11242 -13844 11266 -13810
rect 11300 -13844 11324 -13810
rect 11242 -13868 11324 -13844
rect 12260 -13810 12342 -13786
rect 12260 -13844 12284 -13810
rect 12318 -13844 12342 -13810
rect 12260 -13868 12342 -13844
rect 13278 -13810 13360 -13786
rect 13278 -13844 13302 -13810
rect 13336 -13844 13360 -13810
rect 13278 -13868 13360 -13844
rect 14296 -13810 14378 -13786
rect 14296 -13844 14320 -13810
rect 14354 -13844 14378 -13810
rect 14296 -13868 14378 -13844
rect 15314 -13810 15396 -13786
rect 15314 -13844 15338 -13810
rect 15372 -13844 15396 -13810
rect 15314 -13868 15396 -13844
rect 16332 -13810 16414 -13786
rect 16332 -13844 16356 -13810
rect 16390 -13844 16414 -13810
rect 16332 -13868 16414 -13844
rect 17350 -13810 17432 -13786
rect 17350 -13844 17374 -13810
rect 17408 -13844 17432 -13810
rect 17350 -13868 17432 -13844
rect 18368 -13810 18450 -13786
rect 18368 -13844 18392 -13810
rect 18426 -13844 18450 -13810
rect 18368 -13868 18450 -13844
rect 19386 -13810 19468 -13786
rect 19386 -13844 19410 -13810
rect 19444 -13844 19468 -13810
rect 19386 -13868 19468 -13844
rect 20404 -13810 20486 -13786
rect 20404 -13844 20428 -13810
rect 20462 -13844 20486 -13810
rect 20404 -13868 20486 -13844
rect 21422 -13810 21504 -13786
rect 21422 -13844 21446 -13810
rect 21480 -13844 21504 -13810
rect 21422 -13868 21504 -13844
rect 22440 -13810 22522 -13786
rect 22440 -13844 22464 -13810
rect 22498 -13844 22522 -13810
rect 22440 -13868 22522 -13844
rect -9208 -14022 -9126 -13998
rect -9208 -14056 -9184 -14022
rect -9150 -14056 -9126 -14022
rect -9208 -14080 -9126 -14056
rect -8190 -14022 -8108 -13998
rect -8190 -14056 -8166 -14022
rect -8132 -14056 -8108 -14022
rect -8190 -14080 -8108 -14056
rect -7172 -14022 -7090 -13998
rect -7172 -14056 -7148 -14022
rect -7114 -14056 -7090 -14022
rect -7172 -14080 -7090 -14056
rect -6154 -14022 -6072 -13998
rect -6154 -14056 -6130 -14022
rect -6096 -14056 -6072 -14022
rect -6154 -14080 -6072 -14056
rect -5136 -14022 -5054 -13998
rect -5136 -14056 -5112 -14022
rect -5078 -14056 -5054 -14022
rect -5136 -14080 -5054 -14056
rect -4118 -14022 -4036 -13998
rect -4118 -14056 -4094 -14022
rect -4060 -14056 -4036 -14022
rect -4118 -14080 -4036 -14056
rect -3100 -14022 -3018 -13998
rect -3100 -14056 -3076 -14022
rect -3042 -14056 -3018 -14022
rect -3100 -14080 -3018 -14056
rect -2082 -14022 -2000 -13998
rect -2082 -14056 -2058 -14022
rect -2024 -14056 -2000 -14022
rect -2082 -14080 -2000 -14056
rect -1064 -14022 -982 -13998
rect -1064 -14056 -1040 -14022
rect -1006 -14056 -982 -14022
rect -1064 -14080 -982 -14056
rect -36 -14022 46 -13998
rect -36 -14056 -12 -14022
rect 22 -14056 46 -14022
rect -36 -14080 46 -14056
rect -9208 -14840 -9126 -14816
rect -9208 -14874 -9184 -14840
rect -9150 -14874 -9126 -14840
rect -9208 -14898 -9126 -14874
rect -8190 -14840 -8108 -14816
rect -8190 -14874 -8166 -14840
rect -8132 -14874 -8108 -14840
rect -8190 -14898 -8108 -14874
rect -7172 -14840 -7090 -14816
rect -7172 -14874 -7148 -14840
rect -7114 -14874 -7090 -14840
rect -7172 -14898 -7090 -14874
rect -6154 -14840 -6072 -14816
rect -6154 -14874 -6130 -14840
rect -6096 -14874 -6072 -14840
rect -6154 -14898 -6072 -14874
rect -5136 -14840 -5054 -14816
rect -5136 -14874 -5112 -14840
rect -5078 -14874 -5054 -14840
rect -5136 -14898 -5054 -14874
rect -4118 -14840 -4036 -14816
rect -4118 -14874 -4094 -14840
rect -4060 -14874 -4036 -14840
rect -4118 -14898 -4036 -14874
rect -3100 -14840 -3018 -14816
rect -3100 -14874 -3076 -14840
rect -3042 -14874 -3018 -14840
rect -3100 -14898 -3018 -14874
rect -2082 -14840 -2000 -14816
rect -2082 -14874 -2058 -14840
rect -2024 -14874 -2000 -14840
rect -2082 -14898 -2000 -14874
rect -1064 -14840 -982 -14816
rect -1064 -14874 -1040 -14840
rect -1006 -14874 -982 -14840
rect -1064 -14898 -982 -14874
rect -36 -14840 46 -14816
rect -36 -14874 -12 -14840
rect 22 -14874 46 -14840
rect -36 -14898 46 -14874
rect 3086 -15116 3168 -15092
rect 3086 -15150 3110 -15116
rect 3144 -15150 3168 -15116
rect 3086 -15174 3168 -15150
rect 4104 -15116 4186 -15092
rect 4104 -15150 4128 -15116
rect 4162 -15150 4186 -15116
rect 4104 -15174 4186 -15150
rect 5122 -15116 5204 -15092
rect 5122 -15150 5146 -15116
rect 5180 -15150 5204 -15116
rect 5122 -15174 5204 -15150
rect 6140 -15116 6222 -15092
rect 6140 -15150 6164 -15116
rect 6198 -15150 6222 -15116
rect 6140 -15174 6222 -15150
rect 7158 -15116 7240 -15092
rect 7158 -15150 7182 -15116
rect 7216 -15150 7240 -15116
rect 7158 -15174 7240 -15150
rect 8176 -15116 8258 -15092
rect 8176 -15150 8200 -15116
rect 8234 -15150 8258 -15116
rect 8176 -15174 8258 -15150
rect 9194 -15116 9276 -15092
rect 9194 -15150 9218 -15116
rect 9252 -15150 9276 -15116
rect 9194 -15174 9276 -15150
rect 10212 -15116 10294 -15092
rect 10212 -15150 10236 -15116
rect 10270 -15150 10294 -15116
rect 10212 -15174 10294 -15150
rect 11230 -15116 11312 -15092
rect 11230 -15150 11254 -15116
rect 11288 -15150 11312 -15116
rect 11230 -15174 11312 -15150
rect 12248 -15116 12330 -15092
rect 12248 -15150 12272 -15116
rect 12306 -15150 12330 -15116
rect 12248 -15174 12330 -15150
rect 13266 -15116 13348 -15092
rect 13266 -15150 13290 -15116
rect 13324 -15150 13348 -15116
rect 13266 -15174 13348 -15150
rect 14284 -15116 14366 -15092
rect 14284 -15150 14308 -15116
rect 14342 -15150 14366 -15116
rect 14284 -15174 14366 -15150
rect 15302 -15116 15384 -15092
rect 15302 -15150 15326 -15116
rect 15360 -15150 15384 -15116
rect 15302 -15174 15384 -15150
rect 16320 -15116 16402 -15092
rect 16320 -15150 16344 -15116
rect 16378 -15150 16402 -15116
rect 16320 -15174 16402 -15150
rect 17338 -15116 17420 -15092
rect 17338 -15150 17362 -15116
rect 17396 -15150 17420 -15116
rect 17338 -15174 17420 -15150
rect 18356 -15116 18438 -15092
rect 18356 -15150 18380 -15116
rect 18414 -15150 18438 -15116
rect 18356 -15174 18438 -15150
rect 19374 -15116 19456 -15092
rect 19374 -15150 19398 -15116
rect 19432 -15150 19456 -15116
rect 19374 -15174 19456 -15150
rect 20392 -15116 20474 -15092
rect 20392 -15150 20416 -15116
rect 20450 -15150 20474 -15116
rect 20392 -15174 20474 -15150
rect 21410 -15116 21492 -15092
rect 21410 -15150 21434 -15116
rect 21468 -15150 21492 -15116
rect 21410 -15174 21492 -15150
rect 22428 -15116 22510 -15092
rect 22428 -15150 22452 -15116
rect 22486 -15150 22510 -15116
rect 22428 -15174 22510 -15150
rect -9208 -15658 -9126 -15634
rect -9208 -15692 -9184 -15658
rect -9150 -15692 -9126 -15658
rect -9208 -15716 -9126 -15692
rect -8190 -15658 -8108 -15634
rect -8190 -15692 -8166 -15658
rect -8132 -15692 -8108 -15658
rect -8190 -15716 -8108 -15692
rect -7172 -15658 -7090 -15634
rect -7172 -15692 -7148 -15658
rect -7114 -15692 -7090 -15658
rect -7172 -15716 -7090 -15692
rect -6154 -15658 -6072 -15634
rect -6154 -15692 -6130 -15658
rect -6096 -15692 -6072 -15658
rect -6154 -15716 -6072 -15692
rect -5136 -15658 -5054 -15634
rect -5136 -15692 -5112 -15658
rect -5078 -15692 -5054 -15658
rect -5136 -15716 -5054 -15692
rect -4118 -15658 -4036 -15634
rect -4118 -15692 -4094 -15658
rect -4060 -15692 -4036 -15658
rect -4118 -15716 -4036 -15692
rect -3100 -15658 -3018 -15634
rect -3100 -15692 -3076 -15658
rect -3042 -15692 -3018 -15658
rect -3100 -15716 -3018 -15692
rect -2082 -15658 -2000 -15634
rect -2082 -15692 -2058 -15658
rect -2024 -15692 -2000 -15658
rect -2082 -15716 -2000 -15692
rect -1064 -15658 -982 -15634
rect -1064 -15692 -1040 -15658
rect -1006 -15692 -982 -15658
rect -1064 -15716 -982 -15692
rect -36 -15658 46 -15634
rect -36 -15692 -12 -15658
rect 22 -15692 46 -15658
rect -36 -15716 46 -15692
rect 3074 -16352 3156 -16328
rect -9208 -16476 -9126 -16452
rect -9208 -16510 -9184 -16476
rect -9150 -16510 -9126 -16476
rect -9208 -16534 -9126 -16510
rect -8190 -16476 -8108 -16452
rect -8190 -16510 -8166 -16476
rect -8132 -16510 -8108 -16476
rect -8190 -16534 -8108 -16510
rect -7172 -16476 -7090 -16452
rect -7172 -16510 -7148 -16476
rect -7114 -16510 -7090 -16476
rect -7172 -16534 -7090 -16510
rect -6154 -16476 -6072 -16452
rect -6154 -16510 -6130 -16476
rect -6096 -16510 -6072 -16476
rect -6154 -16534 -6072 -16510
rect -5136 -16476 -5054 -16452
rect -5136 -16510 -5112 -16476
rect -5078 -16510 -5054 -16476
rect -5136 -16534 -5054 -16510
rect -4118 -16476 -4036 -16452
rect -4118 -16510 -4094 -16476
rect -4060 -16510 -4036 -16476
rect -4118 -16534 -4036 -16510
rect -3100 -16476 -3018 -16452
rect -3100 -16510 -3076 -16476
rect -3042 -16510 -3018 -16476
rect -3100 -16534 -3018 -16510
rect -2082 -16476 -2000 -16452
rect 3074 -16386 3098 -16352
rect 3132 -16386 3156 -16352
rect 3074 -16410 3156 -16386
rect 4092 -16352 4174 -16328
rect 4092 -16386 4116 -16352
rect 4150 -16386 4174 -16352
rect 4092 -16410 4174 -16386
rect 5110 -16352 5192 -16328
rect 5110 -16386 5134 -16352
rect 5168 -16386 5192 -16352
rect 5110 -16410 5192 -16386
rect 6128 -16352 6210 -16328
rect 6128 -16386 6152 -16352
rect 6186 -16386 6210 -16352
rect 6128 -16410 6210 -16386
rect 7146 -16352 7228 -16328
rect 7146 -16386 7170 -16352
rect 7204 -16386 7228 -16352
rect 7146 -16410 7228 -16386
rect 8164 -16352 8246 -16328
rect 8164 -16386 8188 -16352
rect 8222 -16386 8246 -16352
rect 8164 -16410 8246 -16386
rect 9182 -16352 9264 -16328
rect 9182 -16386 9206 -16352
rect 9240 -16386 9264 -16352
rect 9182 -16410 9264 -16386
rect 10200 -16352 10282 -16328
rect 10200 -16386 10224 -16352
rect 10258 -16386 10282 -16352
rect 10200 -16410 10282 -16386
rect 11218 -16352 11300 -16328
rect 11218 -16386 11242 -16352
rect 11276 -16386 11300 -16352
rect 11218 -16410 11300 -16386
rect 12236 -16352 12318 -16328
rect 12236 -16386 12260 -16352
rect 12294 -16386 12318 -16352
rect 12236 -16410 12318 -16386
rect 13254 -16352 13336 -16328
rect 13254 -16386 13278 -16352
rect 13312 -16386 13336 -16352
rect 13254 -16410 13336 -16386
rect 14272 -16352 14354 -16328
rect 14272 -16386 14296 -16352
rect 14330 -16386 14354 -16352
rect 14272 -16410 14354 -16386
rect 15290 -16352 15372 -16328
rect 15290 -16386 15314 -16352
rect 15348 -16386 15372 -16352
rect 15290 -16410 15372 -16386
rect 16308 -16352 16390 -16328
rect 16308 -16386 16332 -16352
rect 16366 -16386 16390 -16352
rect 16308 -16410 16390 -16386
rect 17326 -16352 17408 -16328
rect 17326 -16386 17350 -16352
rect 17384 -16386 17408 -16352
rect 17326 -16410 17408 -16386
rect 18344 -16352 18426 -16328
rect 18344 -16386 18368 -16352
rect 18402 -16386 18426 -16352
rect 18344 -16410 18426 -16386
rect 19362 -16352 19444 -16328
rect 19362 -16386 19386 -16352
rect 19420 -16386 19444 -16352
rect 19362 -16410 19444 -16386
rect 20380 -16352 20462 -16328
rect 20380 -16386 20404 -16352
rect 20438 -16386 20462 -16352
rect 20380 -16410 20462 -16386
rect 21398 -16352 21480 -16328
rect 21398 -16386 21422 -16352
rect 21456 -16386 21480 -16352
rect 21398 -16410 21480 -16386
rect 22416 -16352 22498 -16328
rect 22416 -16386 22440 -16352
rect 22474 -16386 22498 -16352
rect 22416 -16410 22498 -16386
rect -2082 -16510 -2058 -16476
rect -2024 -16510 -2000 -16476
rect -2082 -16534 -2000 -16510
rect -1064 -16476 -982 -16452
rect -1064 -16510 -1040 -16476
rect -1006 -16510 -982 -16476
rect -1064 -16534 -982 -16510
rect -36 -16476 46 -16452
rect -36 -16510 -12 -16476
rect 22 -16510 46 -16476
rect -36 -16534 46 -16510
rect -9208 -17294 -9126 -17270
rect -9208 -17328 -9184 -17294
rect -9150 -17328 -9126 -17294
rect -9208 -17352 -9126 -17328
rect -8190 -17294 -8108 -17270
rect -8190 -17328 -8166 -17294
rect -8132 -17328 -8108 -17294
rect -8190 -17352 -8108 -17328
rect -7172 -17294 -7090 -17270
rect -7172 -17328 -7148 -17294
rect -7114 -17328 -7090 -17294
rect -7172 -17352 -7090 -17328
rect -6154 -17294 -6072 -17270
rect -6154 -17328 -6130 -17294
rect -6096 -17328 -6072 -17294
rect -6154 -17352 -6072 -17328
rect -5136 -17294 -5054 -17270
rect -5136 -17328 -5112 -17294
rect -5078 -17328 -5054 -17294
rect -5136 -17352 -5054 -17328
rect -4118 -17294 -4036 -17270
rect -4118 -17328 -4094 -17294
rect -4060 -17328 -4036 -17294
rect -4118 -17352 -4036 -17328
rect -3100 -17294 -3018 -17270
rect -3100 -17328 -3076 -17294
rect -3042 -17328 -3018 -17294
rect -3100 -17352 -3018 -17328
rect -2082 -17294 -2000 -17270
rect -2082 -17328 -2058 -17294
rect -2024 -17328 -2000 -17294
rect -2082 -17352 -2000 -17328
rect -1064 -17294 -982 -17270
rect -1064 -17328 -1040 -17294
rect -1006 -17328 -982 -17294
rect -1064 -17352 -982 -17328
rect -36 -17294 46 -17270
rect -36 -17328 -12 -17294
rect 22 -17328 46 -17294
rect -36 -17352 46 -17328
rect 3074 -17576 3156 -17552
rect 3074 -17610 3098 -17576
rect 3132 -17610 3156 -17576
rect 3074 -17634 3156 -17610
rect 4092 -17576 4174 -17552
rect 4092 -17610 4116 -17576
rect 4150 -17610 4174 -17576
rect 4092 -17634 4174 -17610
rect 5110 -17576 5192 -17552
rect 5110 -17610 5134 -17576
rect 5168 -17610 5192 -17576
rect 5110 -17634 5192 -17610
rect 6128 -17576 6210 -17552
rect 6128 -17610 6152 -17576
rect 6186 -17610 6210 -17576
rect 6128 -17634 6210 -17610
rect 7146 -17576 7228 -17552
rect 7146 -17610 7170 -17576
rect 7204 -17610 7228 -17576
rect 7146 -17634 7228 -17610
rect 8164 -17576 8246 -17552
rect 8164 -17610 8188 -17576
rect 8222 -17610 8246 -17576
rect 8164 -17634 8246 -17610
rect 9182 -17576 9264 -17552
rect 9182 -17610 9206 -17576
rect 9240 -17610 9264 -17576
rect 9182 -17634 9264 -17610
rect 10200 -17576 10282 -17552
rect 10200 -17610 10224 -17576
rect 10258 -17610 10282 -17576
rect 10200 -17634 10282 -17610
rect 11218 -17576 11300 -17552
rect 11218 -17610 11242 -17576
rect 11276 -17610 11300 -17576
rect 11218 -17634 11300 -17610
rect 12236 -17576 12318 -17552
rect 12236 -17610 12260 -17576
rect 12294 -17610 12318 -17576
rect 12236 -17634 12318 -17610
rect 13254 -17576 13336 -17552
rect 13254 -17610 13278 -17576
rect 13312 -17610 13336 -17576
rect 13254 -17634 13336 -17610
rect 14272 -17576 14354 -17552
rect 14272 -17610 14296 -17576
rect 14330 -17610 14354 -17576
rect 14272 -17634 14354 -17610
rect 15290 -17576 15372 -17552
rect 15290 -17610 15314 -17576
rect 15348 -17610 15372 -17576
rect 15290 -17634 15372 -17610
rect 16308 -17576 16390 -17552
rect 16308 -17610 16332 -17576
rect 16366 -17610 16390 -17576
rect 16308 -17634 16390 -17610
rect 17326 -17576 17408 -17552
rect 17326 -17610 17350 -17576
rect 17384 -17610 17408 -17576
rect 17326 -17634 17408 -17610
rect 18344 -17576 18426 -17552
rect 18344 -17610 18368 -17576
rect 18402 -17610 18426 -17576
rect 18344 -17634 18426 -17610
rect 19362 -17576 19444 -17552
rect 19362 -17610 19386 -17576
rect 19420 -17610 19444 -17576
rect 19362 -17634 19444 -17610
rect 20380 -17576 20462 -17552
rect 20380 -17610 20404 -17576
rect 20438 -17610 20462 -17576
rect 20380 -17634 20462 -17610
rect 21398 -17576 21480 -17552
rect 21398 -17610 21422 -17576
rect 21456 -17610 21480 -17576
rect 21398 -17634 21480 -17610
rect 22416 -17576 22498 -17552
rect 22416 -17610 22440 -17576
rect 22474 -17610 22498 -17576
rect 22416 -17634 22498 -17610
rect -9208 -18112 -9126 -18088
rect -9208 -18146 -9184 -18112
rect -9150 -18146 -9126 -18112
rect -9208 -18170 -9126 -18146
rect -8190 -18112 -8108 -18088
rect -8190 -18146 -8166 -18112
rect -8132 -18146 -8108 -18112
rect -8190 -18170 -8108 -18146
rect -7172 -18112 -7090 -18088
rect -7172 -18146 -7148 -18112
rect -7114 -18146 -7090 -18112
rect -7172 -18170 -7090 -18146
rect -6154 -18112 -6072 -18088
rect -6154 -18146 -6130 -18112
rect -6096 -18146 -6072 -18112
rect -6154 -18170 -6072 -18146
rect -5136 -18112 -5054 -18088
rect -5136 -18146 -5112 -18112
rect -5078 -18146 -5054 -18112
rect -5136 -18170 -5054 -18146
rect -4118 -18112 -4036 -18088
rect -4118 -18146 -4094 -18112
rect -4060 -18146 -4036 -18112
rect -4118 -18170 -4036 -18146
rect -3100 -18112 -3018 -18088
rect -3100 -18146 -3076 -18112
rect -3042 -18146 -3018 -18112
rect -3100 -18170 -3018 -18146
rect -2082 -18112 -2000 -18088
rect -2082 -18146 -2058 -18112
rect -2024 -18146 -2000 -18112
rect -2082 -18170 -2000 -18146
rect -1064 -18112 -982 -18088
rect -1064 -18146 -1040 -18112
rect -1006 -18146 -982 -18112
rect -1064 -18170 -982 -18146
rect -36 -18112 46 -18088
rect -36 -18146 -12 -18112
rect 22 -18146 46 -18112
rect -36 -18170 46 -18146
rect 3086 -18812 3168 -18788
rect 3086 -18846 3110 -18812
rect 3144 -18846 3168 -18812
rect 3086 -18870 3168 -18846
rect 4104 -18812 4186 -18788
rect 4104 -18846 4128 -18812
rect 4162 -18846 4186 -18812
rect 4104 -18870 4186 -18846
rect 5122 -18812 5204 -18788
rect 5122 -18846 5146 -18812
rect 5180 -18846 5204 -18812
rect 5122 -18870 5204 -18846
rect 6140 -18812 6222 -18788
rect 6140 -18846 6164 -18812
rect 6198 -18846 6222 -18812
rect 6140 -18870 6222 -18846
rect 7158 -18812 7240 -18788
rect 7158 -18846 7182 -18812
rect 7216 -18846 7240 -18812
rect 7158 -18870 7240 -18846
rect 8176 -18812 8258 -18788
rect 8176 -18846 8200 -18812
rect 8234 -18846 8258 -18812
rect 8176 -18870 8258 -18846
rect 9194 -18812 9276 -18788
rect 9194 -18846 9218 -18812
rect 9252 -18846 9276 -18812
rect 9194 -18870 9276 -18846
rect 10212 -18812 10294 -18788
rect 10212 -18846 10236 -18812
rect 10270 -18846 10294 -18812
rect 10212 -18870 10294 -18846
rect 11230 -18812 11312 -18788
rect 11230 -18846 11254 -18812
rect 11288 -18846 11312 -18812
rect 11230 -18870 11312 -18846
rect 12248 -18812 12330 -18788
rect 12248 -18846 12272 -18812
rect 12306 -18846 12330 -18812
rect 12248 -18870 12330 -18846
rect 13266 -18812 13348 -18788
rect 13266 -18846 13290 -18812
rect 13324 -18846 13348 -18812
rect 13266 -18870 13348 -18846
rect 14284 -18812 14366 -18788
rect 14284 -18846 14308 -18812
rect 14342 -18846 14366 -18812
rect 14284 -18870 14366 -18846
rect 15302 -18812 15384 -18788
rect 15302 -18846 15326 -18812
rect 15360 -18846 15384 -18812
rect 15302 -18870 15384 -18846
rect 16320 -18812 16402 -18788
rect 16320 -18846 16344 -18812
rect 16378 -18846 16402 -18812
rect 16320 -18870 16402 -18846
rect 17338 -18812 17420 -18788
rect 17338 -18846 17362 -18812
rect 17396 -18846 17420 -18812
rect 17338 -18870 17420 -18846
rect 18356 -18812 18438 -18788
rect 18356 -18846 18380 -18812
rect 18414 -18846 18438 -18812
rect 18356 -18870 18438 -18846
rect 19374 -18812 19456 -18788
rect 19374 -18846 19398 -18812
rect 19432 -18846 19456 -18812
rect 19374 -18870 19456 -18846
rect 20392 -18812 20474 -18788
rect 20392 -18846 20416 -18812
rect 20450 -18846 20474 -18812
rect 20392 -18870 20474 -18846
rect 21410 -18812 21492 -18788
rect 21410 -18846 21434 -18812
rect 21468 -18846 21492 -18812
rect 21410 -18870 21492 -18846
rect 22428 -18812 22510 -18788
rect 22428 -18846 22452 -18812
rect 22486 -18846 22510 -18812
rect 22428 -18870 22510 -18846
rect -9220 -19006 -9138 -18982
rect -9220 -19040 -9196 -19006
rect -9162 -19040 -9138 -19006
rect -9220 -19064 -9138 -19040
rect -8202 -19006 -8120 -18982
rect -8202 -19040 -8178 -19006
rect -8144 -19040 -8120 -19006
rect -8202 -19064 -8120 -19040
rect -7184 -19006 -7102 -18982
rect -7184 -19040 -7160 -19006
rect -7126 -19040 -7102 -19006
rect -7184 -19064 -7102 -19040
rect -6166 -19006 -6084 -18982
rect -6166 -19040 -6142 -19006
rect -6108 -19040 -6084 -19006
rect -6166 -19064 -6084 -19040
rect -5148 -19006 -5066 -18982
rect -5148 -19040 -5124 -19006
rect -5090 -19040 -5066 -19006
rect -5148 -19064 -5066 -19040
rect -4130 -19006 -4048 -18982
rect -4130 -19040 -4106 -19006
rect -4072 -19040 -4048 -19006
rect -4130 -19064 -4048 -19040
rect -3112 -19006 -3030 -18982
rect -3112 -19040 -3088 -19006
rect -3054 -19040 -3030 -19006
rect -3112 -19064 -3030 -19040
rect -2094 -19006 -2012 -18982
rect -2094 -19040 -2070 -19006
rect -2036 -19040 -2012 -19006
rect -2094 -19064 -2012 -19040
rect -1076 -19006 -994 -18982
rect -1076 -19040 -1052 -19006
rect -1018 -19040 -994 -19006
rect -1076 -19064 -994 -19040
rect -48 -19006 34 -18982
rect -48 -19040 -24 -19006
rect 10 -19040 34 -19006
rect -48 -19064 34 -19040
rect -10016 -19954 -9934 -19930
rect -10016 -19988 -9992 -19954
rect -9958 -19988 -9934 -19954
rect -10016 -20012 -9934 -19988
rect -8998 -19954 -8916 -19930
rect -8998 -19988 -8974 -19954
rect -8940 -19988 -8916 -19954
rect -8998 -20012 -8916 -19988
rect -7980 -19954 -7898 -19930
rect -7980 -19988 -7956 -19954
rect -7922 -19988 -7898 -19954
rect -7980 -20012 -7898 -19988
rect -6962 -19954 -6880 -19930
rect -6962 -19988 -6938 -19954
rect -6904 -19988 -6880 -19954
rect -6962 -20012 -6880 -19988
rect -5944 -19954 -5862 -19930
rect -5944 -19988 -5920 -19954
rect -5886 -19988 -5862 -19954
rect -5944 -20012 -5862 -19988
rect -4926 -19954 -4844 -19930
rect -4926 -19988 -4902 -19954
rect -4868 -19988 -4844 -19954
rect -4926 -20012 -4844 -19988
rect -3908 -19954 -3826 -19930
rect -3908 -19988 -3884 -19954
rect -3850 -19988 -3826 -19954
rect -3908 -20012 -3826 -19988
rect -2890 -19954 -2808 -19930
rect -2890 -19988 -2866 -19954
rect -2832 -19988 -2808 -19954
rect -2890 -20012 -2808 -19988
rect -1872 -19954 -1790 -19930
rect -1872 -19988 -1848 -19954
rect -1814 -19988 -1790 -19954
rect -1872 -20012 -1790 -19988
rect -854 -19954 -772 -19930
rect -854 -19988 -830 -19954
rect -796 -19988 -772 -19954
rect -854 -20012 -772 -19988
rect 164 -19954 246 -19930
rect 164 -19988 188 -19954
rect 222 -19988 246 -19954
rect 164 -20012 246 -19988
rect 3086 -20060 3168 -20036
rect 3086 -20094 3110 -20060
rect 3144 -20094 3168 -20060
rect 3086 -20118 3168 -20094
rect 4104 -20060 4186 -20036
rect 4104 -20094 4128 -20060
rect 4162 -20094 4186 -20060
rect 4104 -20118 4186 -20094
rect 5122 -20060 5204 -20036
rect 5122 -20094 5146 -20060
rect 5180 -20094 5204 -20060
rect 5122 -20118 5204 -20094
rect 6140 -20060 6222 -20036
rect 6140 -20094 6164 -20060
rect 6198 -20094 6222 -20060
rect 6140 -20118 6222 -20094
rect 7158 -20060 7240 -20036
rect 7158 -20094 7182 -20060
rect 7216 -20094 7240 -20060
rect 7158 -20118 7240 -20094
rect 8176 -20060 8258 -20036
rect 8176 -20094 8200 -20060
rect 8234 -20094 8258 -20060
rect 8176 -20118 8258 -20094
rect 9194 -20060 9276 -20036
rect 9194 -20094 9218 -20060
rect 9252 -20094 9276 -20060
rect 9194 -20118 9276 -20094
rect 10212 -20060 10294 -20036
rect 10212 -20094 10236 -20060
rect 10270 -20094 10294 -20060
rect 10212 -20118 10294 -20094
rect 11230 -20060 11312 -20036
rect 11230 -20094 11254 -20060
rect 11288 -20094 11312 -20060
rect 11230 -20118 11312 -20094
rect 12248 -20060 12330 -20036
rect 12248 -20094 12272 -20060
rect 12306 -20094 12330 -20060
rect 12248 -20118 12330 -20094
rect 13266 -20060 13348 -20036
rect 13266 -20094 13290 -20060
rect 13324 -20094 13348 -20060
rect 13266 -20118 13348 -20094
rect 14284 -20060 14366 -20036
rect 14284 -20094 14308 -20060
rect 14342 -20094 14366 -20060
rect 14284 -20118 14366 -20094
rect 15302 -20060 15384 -20036
rect 15302 -20094 15326 -20060
rect 15360 -20094 15384 -20060
rect 15302 -20118 15384 -20094
rect 16320 -20060 16402 -20036
rect 16320 -20094 16344 -20060
rect 16378 -20094 16402 -20060
rect 16320 -20118 16402 -20094
rect 17338 -20060 17420 -20036
rect 17338 -20094 17362 -20060
rect 17396 -20094 17420 -20060
rect 17338 -20118 17420 -20094
rect 18356 -20060 18438 -20036
rect 18356 -20094 18380 -20060
rect 18414 -20094 18438 -20060
rect 18356 -20118 18438 -20094
rect 19374 -20060 19456 -20036
rect 19374 -20094 19398 -20060
rect 19432 -20094 19456 -20060
rect 19374 -20118 19456 -20094
rect 20392 -20060 20474 -20036
rect 20392 -20094 20416 -20060
rect 20450 -20094 20474 -20060
rect 20392 -20118 20474 -20094
rect 21410 -20060 21492 -20036
rect 21410 -20094 21434 -20060
rect 21468 -20094 21492 -20060
rect 21410 -20118 21492 -20094
rect 22428 -20060 22510 -20036
rect 22428 -20094 22452 -20060
rect 22486 -20094 22510 -20060
rect 22428 -20118 22510 -20094
rect -10004 -21096 -9922 -21072
rect -10004 -21130 -9980 -21096
rect -9946 -21130 -9922 -21096
rect -10004 -21154 -9922 -21130
rect -8986 -21096 -8904 -21072
rect -8986 -21130 -8962 -21096
rect -8928 -21130 -8904 -21096
rect -8986 -21154 -8904 -21130
rect -7968 -21096 -7886 -21072
rect -7968 -21130 -7944 -21096
rect -7910 -21130 -7886 -21096
rect -7968 -21154 -7886 -21130
rect -6950 -21096 -6868 -21072
rect -6950 -21130 -6926 -21096
rect -6892 -21130 -6868 -21096
rect -6950 -21154 -6868 -21130
rect -5932 -21096 -5850 -21072
rect -5932 -21130 -5908 -21096
rect -5874 -21130 -5850 -21096
rect -5932 -21154 -5850 -21130
rect -4914 -21096 -4832 -21072
rect -4914 -21130 -4890 -21096
rect -4856 -21130 -4832 -21096
rect -4914 -21154 -4832 -21130
rect -3896 -21096 -3814 -21072
rect -3896 -21130 -3872 -21096
rect -3838 -21130 -3814 -21096
rect -3896 -21154 -3814 -21130
rect -2878 -21096 -2796 -21072
rect -2878 -21130 -2854 -21096
rect -2820 -21130 -2796 -21096
rect -2878 -21154 -2796 -21130
rect -1860 -21096 -1778 -21072
rect -1860 -21130 -1836 -21096
rect -1802 -21130 -1778 -21096
rect -1860 -21154 -1778 -21130
rect -842 -21096 -760 -21072
rect -842 -21130 -818 -21096
rect -784 -21130 -760 -21096
rect -842 -21154 -760 -21130
rect 176 -21096 258 -21072
rect 176 -21130 200 -21096
rect 234 -21130 258 -21096
rect 176 -21154 258 -21130
rect 3062 -21296 3144 -21272
rect 3062 -21330 3086 -21296
rect 3120 -21330 3144 -21296
rect 3062 -21354 3144 -21330
rect 4080 -21296 4162 -21272
rect 4080 -21330 4104 -21296
rect 4138 -21330 4162 -21296
rect 4080 -21354 4162 -21330
rect 5098 -21296 5180 -21272
rect 5098 -21330 5122 -21296
rect 5156 -21330 5180 -21296
rect 5098 -21354 5180 -21330
rect 6116 -21296 6198 -21272
rect 6116 -21330 6140 -21296
rect 6174 -21330 6198 -21296
rect 6116 -21354 6198 -21330
rect 7134 -21296 7216 -21272
rect 7134 -21330 7158 -21296
rect 7192 -21330 7216 -21296
rect 7134 -21354 7216 -21330
rect 8152 -21296 8234 -21272
rect 8152 -21330 8176 -21296
rect 8210 -21330 8234 -21296
rect 8152 -21354 8234 -21330
rect 9170 -21296 9252 -21272
rect 9170 -21330 9194 -21296
rect 9228 -21330 9252 -21296
rect 9170 -21354 9252 -21330
rect 10188 -21296 10270 -21272
rect 10188 -21330 10212 -21296
rect 10246 -21330 10270 -21296
rect 10188 -21354 10270 -21330
rect 11206 -21296 11288 -21272
rect 11206 -21330 11230 -21296
rect 11264 -21330 11288 -21296
rect 11206 -21354 11288 -21330
rect 12224 -21296 12306 -21272
rect 12224 -21330 12248 -21296
rect 12282 -21330 12306 -21296
rect 12224 -21354 12306 -21330
rect 13242 -21296 13324 -21272
rect 13242 -21330 13266 -21296
rect 13300 -21330 13324 -21296
rect 13242 -21354 13324 -21330
rect 14260 -21296 14342 -21272
rect 14260 -21330 14284 -21296
rect 14318 -21330 14342 -21296
rect 14260 -21354 14342 -21330
rect 15278 -21296 15360 -21272
rect 15278 -21330 15302 -21296
rect 15336 -21330 15360 -21296
rect 15278 -21354 15360 -21330
rect 16296 -21296 16378 -21272
rect 16296 -21330 16320 -21296
rect 16354 -21330 16378 -21296
rect 16296 -21354 16378 -21330
rect 17314 -21296 17396 -21272
rect 17314 -21330 17338 -21296
rect 17372 -21330 17396 -21296
rect 17314 -21354 17396 -21330
rect 18332 -21296 18414 -21272
rect 18332 -21330 18356 -21296
rect 18390 -21330 18414 -21296
rect 18332 -21354 18414 -21330
rect 19350 -21296 19432 -21272
rect 19350 -21330 19374 -21296
rect 19408 -21330 19432 -21296
rect 19350 -21354 19432 -21330
rect 20368 -21296 20450 -21272
rect 20368 -21330 20392 -21296
rect 20426 -21330 20450 -21296
rect 20368 -21354 20450 -21330
rect 21386 -21296 21468 -21272
rect 21386 -21330 21410 -21296
rect 21444 -21330 21468 -21296
rect 21386 -21354 21468 -21330
rect 22404 -21296 22486 -21272
rect 22404 -21330 22428 -21296
rect 22462 -21330 22486 -21296
rect 22404 -21354 22486 -21330
rect -10026 -22204 -9944 -22180
rect -10026 -22238 -10002 -22204
rect -9968 -22238 -9944 -22204
rect -10026 -22262 -9944 -22238
rect -9008 -22204 -8926 -22180
rect -9008 -22238 -8984 -22204
rect -8950 -22238 -8926 -22204
rect -9008 -22262 -8926 -22238
rect -7990 -22204 -7908 -22180
rect -7990 -22238 -7966 -22204
rect -7932 -22238 -7908 -22204
rect -7990 -22262 -7908 -22238
rect -6972 -22204 -6890 -22180
rect -6972 -22238 -6948 -22204
rect -6914 -22238 -6890 -22204
rect -6972 -22262 -6890 -22238
rect -5954 -22204 -5872 -22180
rect -5954 -22238 -5930 -22204
rect -5896 -22238 -5872 -22204
rect -5954 -22262 -5872 -22238
rect -4936 -22204 -4854 -22180
rect -4936 -22238 -4912 -22204
rect -4878 -22238 -4854 -22204
rect -4936 -22262 -4854 -22238
rect -3918 -22204 -3836 -22180
rect -3918 -22238 -3894 -22204
rect -3860 -22238 -3836 -22204
rect -3918 -22262 -3836 -22238
rect -2900 -22204 -2818 -22180
rect -2900 -22238 -2876 -22204
rect -2842 -22238 -2818 -22204
rect -2900 -22262 -2818 -22238
rect -1882 -22204 -1800 -22180
rect -1882 -22238 -1858 -22204
rect -1824 -22238 -1800 -22204
rect -1882 -22262 -1800 -22238
rect -864 -22204 -782 -22180
rect -864 -22238 -840 -22204
rect -806 -22238 -782 -22204
rect -864 -22262 -782 -22238
rect 154 -22204 236 -22180
rect 154 -22238 178 -22204
rect 212 -22238 236 -22204
rect 154 -22262 236 -22238
rect 3074 -22520 3156 -22496
rect 3074 -22554 3098 -22520
rect 3132 -22554 3156 -22520
rect 3074 -22578 3156 -22554
rect 4092 -22520 4174 -22496
rect 4092 -22554 4116 -22520
rect 4150 -22554 4174 -22520
rect 4092 -22578 4174 -22554
rect 5110 -22520 5192 -22496
rect 5110 -22554 5134 -22520
rect 5168 -22554 5192 -22520
rect 5110 -22578 5192 -22554
rect 6128 -22520 6210 -22496
rect 6128 -22554 6152 -22520
rect 6186 -22554 6210 -22520
rect 6128 -22578 6210 -22554
rect 7146 -22520 7228 -22496
rect 7146 -22554 7170 -22520
rect 7204 -22554 7228 -22520
rect 7146 -22578 7228 -22554
rect 8164 -22520 8246 -22496
rect 8164 -22554 8188 -22520
rect 8222 -22554 8246 -22520
rect 8164 -22578 8246 -22554
rect 9182 -22520 9264 -22496
rect 9182 -22554 9206 -22520
rect 9240 -22554 9264 -22520
rect 9182 -22578 9264 -22554
rect 10200 -22520 10282 -22496
rect 10200 -22554 10224 -22520
rect 10258 -22554 10282 -22520
rect 10200 -22578 10282 -22554
rect 11218 -22520 11300 -22496
rect 11218 -22554 11242 -22520
rect 11276 -22554 11300 -22520
rect 11218 -22578 11300 -22554
rect 12236 -22520 12318 -22496
rect 12236 -22554 12260 -22520
rect 12294 -22554 12318 -22520
rect 12236 -22578 12318 -22554
rect 13254 -22520 13336 -22496
rect 13254 -22554 13278 -22520
rect 13312 -22554 13336 -22520
rect 13254 -22578 13336 -22554
rect 14272 -22520 14354 -22496
rect 14272 -22554 14296 -22520
rect 14330 -22554 14354 -22520
rect 14272 -22578 14354 -22554
rect 15290 -22520 15372 -22496
rect 15290 -22554 15314 -22520
rect 15348 -22554 15372 -22520
rect 15290 -22578 15372 -22554
rect 16308 -22520 16390 -22496
rect 16308 -22554 16332 -22520
rect 16366 -22554 16390 -22520
rect 16308 -22578 16390 -22554
rect 17326 -22520 17408 -22496
rect 17326 -22554 17350 -22520
rect 17384 -22554 17408 -22520
rect 17326 -22578 17408 -22554
rect 18344 -22520 18426 -22496
rect 18344 -22554 18368 -22520
rect 18402 -22554 18426 -22520
rect 18344 -22578 18426 -22554
rect 19362 -22520 19444 -22496
rect 19362 -22554 19386 -22520
rect 19420 -22554 19444 -22520
rect 19362 -22578 19444 -22554
rect 20380 -22520 20462 -22496
rect 20380 -22554 20404 -22520
rect 20438 -22554 20462 -22520
rect 20380 -22578 20462 -22554
rect 21398 -22520 21480 -22496
rect 21398 -22554 21422 -22520
rect 21456 -22554 21480 -22520
rect 21398 -22578 21480 -22554
rect 22416 -22520 22498 -22496
rect 22416 -22554 22440 -22520
rect 22474 -22554 22498 -22520
rect 22416 -22578 22498 -22554
rect -10026 -23310 -9944 -23286
rect -10026 -23344 -10002 -23310
rect -9968 -23344 -9944 -23310
rect -10026 -23368 -9944 -23344
rect -9008 -23310 -8926 -23286
rect -9008 -23344 -8984 -23310
rect -8950 -23344 -8926 -23310
rect -9008 -23368 -8926 -23344
rect -7990 -23310 -7908 -23286
rect -7990 -23344 -7966 -23310
rect -7932 -23344 -7908 -23310
rect -7990 -23368 -7908 -23344
rect -6972 -23310 -6890 -23286
rect -6972 -23344 -6948 -23310
rect -6914 -23344 -6890 -23310
rect -6972 -23368 -6890 -23344
rect -5954 -23310 -5872 -23286
rect -5954 -23344 -5930 -23310
rect -5896 -23344 -5872 -23310
rect -5954 -23368 -5872 -23344
rect -4936 -23310 -4854 -23286
rect -4936 -23344 -4912 -23310
rect -4878 -23344 -4854 -23310
rect -4936 -23368 -4854 -23344
rect -3918 -23310 -3836 -23286
rect -3918 -23344 -3894 -23310
rect -3860 -23344 -3836 -23310
rect -3918 -23368 -3836 -23344
rect -2900 -23310 -2818 -23286
rect -2900 -23344 -2876 -23310
rect -2842 -23344 -2818 -23310
rect -2900 -23368 -2818 -23344
rect -1882 -23310 -1800 -23286
rect -1882 -23344 -1858 -23310
rect -1824 -23344 -1800 -23310
rect -1882 -23368 -1800 -23344
rect -864 -23310 -782 -23286
rect -864 -23344 -840 -23310
rect -806 -23344 -782 -23310
rect -864 -23368 -782 -23344
rect 154 -23310 236 -23286
rect 154 -23344 178 -23310
rect 212 -23344 236 -23310
rect 154 -23368 236 -23344
rect 3074 -23756 3156 -23732
rect 3074 -23790 3098 -23756
rect 3132 -23790 3156 -23756
rect 3074 -23814 3156 -23790
rect 4092 -23756 4174 -23732
rect 4092 -23790 4116 -23756
rect 4150 -23790 4174 -23756
rect 4092 -23814 4174 -23790
rect 5110 -23756 5192 -23732
rect 5110 -23790 5134 -23756
rect 5168 -23790 5192 -23756
rect 5110 -23814 5192 -23790
rect 6128 -23756 6210 -23732
rect 6128 -23790 6152 -23756
rect 6186 -23790 6210 -23756
rect 6128 -23814 6210 -23790
rect 7146 -23756 7228 -23732
rect 7146 -23790 7170 -23756
rect 7204 -23790 7228 -23756
rect 7146 -23814 7228 -23790
rect 8164 -23756 8246 -23732
rect 8164 -23790 8188 -23756
rect 8222 -23790 8246 -23756
rect 8164 -23814 8246 -23790
rect 9182 -23756 9264 -23732
rect 9182 -23790 9206 -23756
rect 9240 -23790 9264 -23756
rect 9182 -23814 9264 -23790
rect 10200 -23756 10282 -23732
rect 10200 -23790 10224 -23756
rect 10258 -23790 10282 -23756
rect 10200 -23814 10282 -23790
rect 11218 -23756 11300 -23732
rect 11218 -23790 11242 -23756
rect 11276 -23790 11300 -23756
rect 11218 -23814 11300 -23790
rect 12236 -23756 12318 -23732
rect 12236 -23790 12260 -23756
rect 12294 -23790 12318 -23756
rect 12236 -23814 12318 -23790
rect 13254 -23756 13336 -23732
rect 13254 -23790 13278 -23756
rect 13312 -23790 13336 -23756
rect 13254 -23814 13336 -23790
rect 14272 -23756 14354 -23732
rect 14272 -23790 14296 -23756
rect 14330 -23790 14354 -23756
rect 14272 -23814 14354 -23790
rect 15290 -23756 15372 -23732
rect 15290 -23790 15314 -23756
rect 15348 -23790 15372 -23756
rect 15290 -23814 15372 -23790
rect 16308 -23756 16390 -23732
rect 16308 -23790 16332 -23756
rect 16366 -23790 16390 -23756
rect 16308 -23814 16390 -23790
rect 17326 -23756 17408 -23732
rect 17326 -23790 17350 -23756
rect 17384 -23790 17408 -23756
rect 17326 -23814 17408 -23790
rect 18344 -23756 18426 -23732
rect 18344 -23790 18368 -23756
rect 18402 -23790 18426 -23756
rect 18344 -23814 18426 -23790
rect 19362 -23756 19444 -23732
rect 19362 -23790 19386 -23756
rect 19420 -23790 19444 -23756
rect 19362 -23814 19444 -23790
rect 20380 -23756 20462 -23732
rect 20380 -23790 20404 -23756
rect 20438 -23790 20462 -23756
rect 20380 -23814 20462 -23790
rect 21398 -23756 21480 -23732
rect 21398 -23790 21422 -23756
rect 21456 -23790 21480 -23756
rect 21398 -23814 21480 -23790
rect 22416 -23756 22498 -23732
rect 22416 -23790 22440 -23756
rect 22474 -23790 22498 -23756
rect 22416 -23814 22498 -23790
rect -10026 -24652 -9944 -24628
rect -10026 -24686 -10002 -24652
rect -9968 -24686 -9944 -24652
rect -10026 -24710 -9944 -24686
rect -9008 -24652 -8926 -24628
rect -9008 -24686 -8984 -24652
rect -8950 -24686 -8926 -24652
rect -9008 -24710 -8926 -24686
rect -7990 -24652 -7908 -24628
rect -7990 -24686 -7966 -24652
rect -7932 -24686 -7908 -24652
rect -7990 -24710 -7908 -24686
rect -6972 -24652 -6890 -24628
rect -6972 -24686 -6948 -24652
rect -6914 -24686 -6890 -24652
rect -6972 -24710 -6890 -24686
rect -5954 -24652 -5872 -24628
rect -5954 -24686 -5930 -24652
rect -5896 -24686 -5872 -24652
rect -5954 -24710 -5872 -24686
rect -4936 -24652 -4854 -24628
rect -4936 -24686 -4912 -24652
rect -4878 -24686 -4854 -24652
rect -4936 -24710 -4854 -24686
rect -3918 -24652 -3836 -24628
rect -3918 -24686 -3894 -24652
rect -3860 -24686 -3836 -24652
rect -3918 -24710 -3836 -24686
rect -2900 -24652 -2818 -24628
rect -2900 -24686 -2876 -24652
rect -2842 -24686 -2818 -24652
rect -2900 -24710 -2818 -24686
rect -1882 -24652 -1800 -24628
rect -1882 -24686 -1858 -24652
rect -1824 -24686 -1800 -24652
rect -1882 -24710 -1800 -24686
rect -864 -24652 -782 -24628
rect -864 -24686 -840 -24652
rect -806 -24686 -782 -24652
rect -864 -24710 -782 -24686
rect 154 -24652 236 -24628
rect 154 -24686 178 -24652
rect 212 -24686 236 -24652
rect 154 -24710 236 -24686
rect 3086 -25002 3168 -24978
rect 3086 -25036 3110 -25002
rect 3144 -25036 3168 -25002
rect 3086 -25060 3168 -25036
rect 4104 -25002 4186 -24978
rect 4104 -25036 4128 -25002
rect 4162 -25036 4186 -25002
rect 4104 -25060 4186 -25036
rect 5122 -25002 5204 -24978
rect 5122 -25036 5146 -25002
rect 5180 -25036 5204 -25002
rect 5122 -25060 5204 -25036
rect 6140 -25002 6222 -24978
rect 6140 -25036 6164 -25002
rect 6198 -25036 6222 -25002
rect 6140 -25060 6222 -25036
rect 7158 -25002 7240 -24978
rect 7158 -25036 7182 -25002
rect 7216 -25036 7240 -25002
rect 7158 -25060 7240 -25036
rect 8176 -25002 8258 -24978
rect 8176 -25036 8200 -25002
rect 8234 -25036 8258 -25002
rect 8176 -25060 8258 -25036
rect 9194 -25002 9276 -24978
rect 9194 -25036 9218 -25002
rect 9252 -25036 9276 -25002
rect 9194 -25060 9276 -25036
rect 10212 -25002 10294 -24978
rect 10212 -25036 10236 -25002
rect 10270 -25036 10294 -25002
rect 10212 -25060 10294 -25036
rect 11230 -25002 11312 -24978
rect 11230 -25036 11254 -25002
rect 11288 -25036 11312 -25002
rect 11230 -25060 11312 -25036
rect 12248 -25002 12330 -24978
rect 12248 -25036 12272 -25002
rect 12306 -25036 12330 -25002
rect 12248 -25060 12330 -25036
rect 13266 -25002 13348 -24978
rect 13266 -25036 13290 -25002
rect 13324 -25036 13348 -25002
rect 13266 -25060 13348 -25036
rect 14284 -25002 14366 -24978
rect 14284 -25036 14308 -25002
rect 14342 -25036 14366 -25002
rect 14284 -25060 14366 -25036
rect 15302 -25002 15384 -24978
rect 15302 -25036 15326 -25002
rect 15360 -25036 15384 -25002
rect 15302 -25060 15384 -25036
rect 16320 -25002 16402 -24978
rect 16320 -25036 16344 -25002
rect 16378 -25036 16402 -25002
rect 16320 -25060 16402 -25036
rect 17338 -25002 17420 -24978
rect 17338 -25036 17362 -25002
rect 17396 -25036 17420 -25002
rect 17338 -25060 17420 -25036
rect 18356 -25002 18438 -24978
rect 18356 -25036 18380 -25002
rect 18414 -25036 18438 -25002
rect 18356 -25060 18438 -25036
rect 19374 -25002 19456 -24978
rect 19374 -25036 19398 -25002
rect 19432 -25036 19456 -25002
rect 19374 -25060 19456 -25036
rect 20392 -25002 20474 -24978
rect 20392 -25036 20416 -25002
rect 20450 -25036 20474 -25002
rect 20392 -25060 20474 -25036
rect 21410 -25002 21492 -24978
rect 21410 -25036 21434 -25002
rect 21468 -25036 21492 -25002
rect 21410 -25060 21492 -25036
rect 22428 -25002 22510 -24978
rect 22428 -25036 22452 -25002
rect 22486 -25036 22510 -25002
rect 22428 -25060 22510 -25036
rect -10216 -26098 -10134 -26074
rect -10216 -26132 -10192 -26098
rect -10158 -26132 -10134 -26098
rect -10216 -26156 -10134 -26132
rect -9198 -26098 -9116 -26074
rect -9198 -26132 -9174 -26098
rect -9140 -26132 -9116 -26098
rect -9198 -26156 -9116 -26132
rect -8180 -26098 -8098 -26074
rect -8180 -26132 -8156 -26098
rect -8122 -26132 -8098 -26098
rect -8180 -26156 -8098 -26132
rect -7162 -26098 -7080 -26074
rect -7162 -26132 -7138 -26098
rect -7104 -26132 -7080 -26098
rect -7162 -26156 -7080 -26132
rect -6144 -26098 -6062 -26074
rect -6144 -26132 -6120 -26098
rect -6086 -26132 -6062 -26098
rect -6144 -26156 -6062 -26132
rect -5126 -26098 -5044 -26074
rect -5126 -26132 -5102 -26098
rect -5068 -26132 -5044 -26098
rect -5126 -26156 -5044 -26132
rect -4108 -26098 -4026 -26074
rect -4108 -26132 -4084 -26098
rect -4050 -26132 -4026 -26098
rect -4108 -26156 -4026 -26132
rect -3090 -26098 -3008 -26074
rect -3090 -26132 -3066 -26098
rect -3032 -26132 -3008 -26098
rect -3090 -26156 -3008 -26132
rect -2072 -26098 -1990 -26074
rect -2072 -26132 -2048 -26098
rect -2014 -26132 -1990 -26098
rect -2072 -26156 -1990 -26132
rect -1054 -26098 -972 -26074
rect -1054 -26132 -1030 -26098
rect -996 -26132 -972 -26098
rect -1054 -26156 -972 -26132
rect -36 -26098 46 -26074
rect -36 -26132 -12 -26098
rect 22 -26132 46 -26098
rect -36 -26156 46 -26132
rect 3074 -26180 3156 -26156
rect 3074 -26214 3098 -26180
rect 3132 -26214 3156 -26180
rect 3074 -26238 3156 -26214
rect 4092 -26180 4174 -26156
rect 4092 -26214 4116 -26180
rect 4150 -26214 4174 -26180
rect 4092 -26238 4174 -26214
rect 5110 -26180 5192 -26156
rect 5110 -26214 5134 -26180
rect 5168 -26214 5192 -26180
rect 5110 -26238 5192 -26214
rect 6128 -26180 6210 -26156
rect 6128 -26214 6152 -26180
rect 6186 -26214 6210 -26180
rect 6128 -26238 6210 -26214
rect 7146 -26180 7228 -26156
rect 7146 -26214 7170 -26180
rect 7204 -26214 7228 -26180
rect 7146 -26238 7228 -26214
rect 8164 -26180 8246 -26156
rect 8164 -26214 8188 -26180
rect 8222 -26214 8246 -26180
rect 8164 -26238 8246 -26214
rect 9182 -26180 9264 -26156
rect 9182 -26214 9206 -26180
rect 9240 -26214 9264 -26180
rect 9182 -26238 9264 -26214
rect 10200 -26180 10282 -26156
rect 10200 -26214 10224 -26180
rect 10258 -26214 10282 -26180
rect 10200 -26238 10282 -26214
rect 11218 -26180 11300 -26156
rect 11218 -26214 11242 -26180
rect 11276 -26214 11300 -26180
rect 11218 -26238 11300 -26214
rect 12236 -26180 12318 -26156
rect 12236 -26214 12260 -26180
rect 12294 -26214 12318 -26180
rect 12236 -26238 12318 -26214
rect 13254 -26180 13336 -26156
rect 13254 -26214 13278 -26180
rect 13312 -26214 13336 -26180
rect 13254 -26238 13336 -26214
rect 14272 -26180 14354 -26156
rect 14272 -26214 14296 -26180
rect 14330 -26214 14354 -26180
rect 14272 -26238 14354 -26214
rect 15290 -26180 15372 -26156
rect 15290 -26214 15314 -26180
rect 15348 -26214 15372 -26180
rect 15290 -26238 15372 -26214
rect 16308 -26180 16390 -26156
rect 16308 -26214 16332 -26180
rect 16366 -26214 16390 -26180
rect 16308 -26238 16390 -26214
rect 17326 -26180 17408 -26156
rect 17326 -26214 17350 -26180
rect 17384 -26214 17408 -26180
rect 17326 -26238 17408 -26214
rect 18344 -26180 18426 -26156
rect 18344 -26214 18368 -26180
rect 18402 -26214 18426 -26180
rect 18344 -26238 18426 -26214
rect 19362 -26180 19444 -26156
rect 19362 -26214 19386 -26180
rect 19420 -26214 19444 -26180
rect 19362 -26238 19444 -26214
rect 20380 -26180 20462 -26156
rect 20380 -26214 20404 -26180
rect 20438 -26214 20462 -26180
rect 20380 -26238 20462 -26214
rect 21398 -26180 21480 -26156
rect 21398 -26214 21422 -26180
rect 21456 -26214 21480 -26180
rect 21398 -26238 21480 -26214
rect 22416 -26180 22498 -26156
rect 22416 -26214 22440 -26180
rect 22474 -26214 22498 -26180
rect 22416 -26238 22498 -26214
rect -12322 -27122 -12222 -27060
rect 24822 -27122 24922 -27060
rect -12322 -27222 -12160 -27122
rect 24760 -27222 24922 -27122
<< nsubdiff >>
rect 378 4222 540 4322
rect 24660 4222 24822 4322
rect 378 4160 478 4222
rect 24722 4160 24822 4222
rect 6972 1778 7054 1804
rect 6972 1744 6996 1778
rect 7030 1744 7054 1778
rect 6972 1720 7054 1744
rect 7990 1778 8072 1804
rect 7990 1744 8014 1778
rect 8048 1744 8072 1778
rect 7990 1720 8072 1744
rect 9008 1778 9090 1804
rect 9008 1744 9032 1778
rect 9066 1744 9090 1778
rect 9008 1720 9090 1744
rect 10026 1778 10108 1804
rect 10026 1744 10050 1778
rect 10084 1744 10108 1778
rect 10026 1720 10108 1744
rect 11044 1778 11126 1804
rect 11044 1744 11068 1778
rect 11102 1744 11126 1778
rect 11044 1720 11126 1744
rect 12062 1778 12144 1804
rect 12062 1744 12086 1778
rect 12120 1744 12144 1778
rect 12062 1720 12144 1744
rect 13080 1778 13162 1804
rect 13080 1744 13104 1778
rect 13138 1744 13162 1778
rect 13080 1720 13162 1744
rect 14098 1778 14180 1804
rect 14098 1744 14122 1778
rect 14156 1744 14180 1778
rect 14098 1720 14180 1744
rect 15116 1778 15198 1804
rect 15116 1744 15140 1778
rect 15174 1744 15198 1778
rect 15116 1720 15198 1744
rect 16134 1778 16216 1804
rect 16134 1744 16158 1778
rect 16192 1744 16216 1778
rect 16134 1720 16216 1744
rect 17152 1778 17234 1804
rect 17152 1744 17176 1778
rect 17210 1744 17234 1778
rect 17152 1720 17234 1744
rect 18170 1778 18252 1804
rect 18170 1744 18194 1778
rect 18228 1744 18252 1778
rect 18170 1720 18252 1744
rect 19188 1778 19270 1804
rect 19188 1744 19212 1778
rect 19246 1744 19270 1778
rect 19188 1720 19270 1744
rect 20206 1778 20288 1804
rect 20206 1744 20230 1778
rect 20264 1744 20288 1778
rect 20206 1720 20288 1744
rect 21224 1778 21306 1804
rect 21224 1744 21248 1778
rect 21282 1744 21306 1778
rect 21224 1720 21306 1744
rect 22242 1778 22324 1804
rect 22242 1744 22266 1778
rect 22300 1744 22324 1778
rect 22242 1720 22324 1744
rect 6994 624 7076 650
rect 6994 590 7018 624
rect 7052 590 7076 624
rect 6994 566 7076 590
rect 8012 624 8094 650
rect 8012 590 8036 624
rect 8070 590 8094 624
rect 8012 566 8094 590
rect 9030 624 9112 650
rect 9030 590 9054 624
rect 9088 590 9112 624
rect 9030 566 9112 590
rect 10048 624 10130 650
rect 10048 590 10072 624
rect 10106 590 10130 624
rect 10048 566 10130 590
rect 11066 624 11148 650
rect 11066 590 11090 624
rect 11124 590 11148 624
rect 11066 566 11148 590
rect 12084 624 12166 650
rect 12084 590 12108 624
rect 12142 590 12166 624
rect 12084 566 12166 590
rect 13102 624 13184 650
rect 13102 590 13126 624
rect 13160 590 13184 624
rect 13102 566 13184 590
rect 14120 624 14202 650
rect 14120 590 14144 624
rect 14178 590 14202 624
rect 14120 566 14202 590
rect 15138 624 15220 650
rect 15138 590 15162 624
rect 15196 590 15220 624
rect 15138 566 15220 590
rect 16156 624 16238 650
rect 16156 590 16180 624
rect 16214 590 16238 624
rect 16156 566 16238 590
rect 17174 624 17256 650
rect 17174 590 17198 624
rect 17232 590 17256 624
rect 17174 566 17256 590
rect 18192 624 18274 650
rect 18192 590 18216 624
rect 18250 590 18274 624
rect 18192 566 18274 590
rect 19210 624 19292 650
rect 19210 590 19234 624
rect 19268 590 19292 624
rect 19210 566 19292 590
rect 20228 624 20310 650
rect 20228 590 20252 624
rect 20286 590 20310 624
rect 20228 566 20310 590
rect 21246 624 21328 650
rect 21246 590 21270 624
rect 21304 590 21328 624
rect 21246 566 21328 590
rect 22264 624 22346 650
rect 22264 590 22288 624
rect 22322 590 22346 624
rect 22264 566 22346 590
rect 6972 -508 7054 -482
rect 6972 -542 6996 -508
rect 7030 -542 7054 -508
rect 6972 -566 7054 -542
rect 7990 -508 8072 -482
rect 7990 -542 8014 -508
rect 8048 -542 8072 -508
rect 7990 -566 8072 -542
rect 9008 -508 9090 -482
rect 9008 -542 9032 -508
rect 9066 -542 9090 -508
rect 9008 -566 9090 -542
rect 10026 -508 10108 -482
rect 10026 -542 10050 -508
rect 10084 -542 10108 -508
rect 10026 -566 10108 -542
rect 11044 -508 11126 -482
rect 11044 -542 11068 -508
rect 11102 -542 11126 -508
rect 11044 -566 11126 -542
rect 12062 -508 12144 -482
rect 12062 -542 12086 -508
rect 12120 -542 12144 -508
rect 12062 -566 12144 -542
rect 13080 -508 13162 -482
rect 13080 -542 13104 -508
rect 13138 -542 13162 -508
rect 13080 -566 13162 -542
rect 14098 -508 14180 -482
rect 14098 -542 14122 -508
rect 14156 -542 14180 -508
rect 14098 -566 14180 -542
rect 15116 -508 15198 -482
rect 15116 -542 15140 -508
rect 15174 -542 15198 -508
rect 15116 -566 15198 -542
rect 16134 -508 16216 -482
rect 16134 -542 16158 -508
rect 16192 -542 16216 -508
rect 16134 -566 16216 -542
rect 17152 -508 17234 -482
rect 17152 -542 17176 -508
rect 17210 -542 17234 -508
rect 17152 -566 17234 -542
rect 18170 -508 18252 -482
rect 18170 -542 18194 -508
rect 18228 -542 18252 -508
rect 18170 -566 18252 -542
rect 19188 -508 19270 -482
rect 19188 -542 19212 -508
rect 19246 -542 19270 -508
rect 19188 -566 19270 -542
rect 20206 -508 20288 -482
rect 20206 -542 20230 -508
rect 20264 -542 20288 -508
rect 20206 -566 20288 -542
rect 21224 -508 21306 -482
rect 21224 -542 21248 -508
rect 21282 -542 21306 -508
rect 21224 -566 21306 -542
rect 22242 -508 22324 -482
rect 22242 -542 22266 -508
rect 22300 -542 22324 -508
rect 22242 -566 22324 -542
rect 6972 -1890 7054 -1864
rect 6972 -1924 6996 -1890
rect 7030 -1924 7054 -1890
rect 6972 -1948 7054 -1924
rect 7990 -1890 8072 -1864
rect 7990 -1924 8014 -1890
rect 8048 -1924 8072 -1890
rect 7990 -1948 8072 -1924
rect 9008 -1890 9090 -1864
rect 9008 -1924 9032 -1890
rect 9066 -1924 9090 -1890
rect 9008 -1948 9090 -1924
rect 10026 -1890 10108 -1864
rect 10026 -1924 10050 -1890
rect 10084 -1924 10108 -1890
rect 10026 -1948 10108 -1924
rect 11044 -1890 11126 -1864
rect 11044 -1924 11068 -1890
rect 11102 -1924 11126 -1890
rect 11044 -1948 11126 -1924
rect 12062 -1890 12144 -1864
rect 12062 -1924 12086 -1890
rect 12120 -1924 12144 -1890
rect 12062 -1948 12144 -1924
rect 13080 -1890 13162 -1864
rect 13080 -1924 13104 -1890
rect 13138 -1924 13162 -1890
rect 13080 -1948 13162 -1924
rect 14098 -1890 14180 -1864
rect 14098 -1924 14122 -1890
rect 14156 -1924 14180 -1890
rect 14098 -1948 14180 -1924
rect 15116 -1890 15198 -1864
rect 15116 -1924 15140 -1890
rect 15174 -1924 15198 -1890
rect 15116 -1948 15198 -1924
rect 16134 -1890 16216 -1864
rect 16134 -1924 16158 -1890
rect 16192 -1924 16216 -1890
rect 16134 -1948 16216 -1924
rect 17152 -1890 17234 -1864
rect 17152 -1924 17176 -1890
rect 17210 -1924 17234 -1890
rect 17152 -1948 17234 -1924
rect 18170 -1890 18252 -1864
rect 18170 -1924 18194 -1890
rect 18228 -1924 18252 -1890
rect 18170 -1948 18252 -1924
rect 19188 -1890 19270 -1864
rect 19188 -1924 19212 -1890
rect 19246 -1924 19270 -1890
rect 19188 -1948 19270 -1924
rect 20206 -1890 20288 -1864
rect 20206 -1924 20230 -1890
rect 20264 -1924 20288 -1890
rect 20206 -1948 20288 -1924
rect 21224 -1890 21306 -1864
rect 21224 -1924 21248 -1890
rect 21282 -1924 21306 -1890
rect 21224 -1948 21306 -1924
rect 22242 -1890 22324 -1864
rect 22242 -1924 22266 -1890
rect 22300 -1924 22324 -1890
rect 22242 -1948 22324 -1924
rect 7660 -3238 7742 -3212
rect 7660 -3272 7684 -3238
rect 7718 -3272 7742 -3238
rect 7660 -3296 7742 -3272
rect 8678 -3238 8760 -3212
rect 8678 -3272 8702 -3238
rect 8736 -3272 8760 -3238
rect 8678 -3296 8760 -3272
rect 9696 -3238 9778 -3212
rect 9696 -3272 9720 -3238
rect 9754 -3272 9778 -3238
rect 9696 -3296 9778 -3272
rect 10714 -3238 10796 -3212
rect 10714 -3272 10738 -3238
rect 10772 -3272 10796 -3238
rect 10714 -3296 10796 -3272
rect 11732 -3238 11814 -3212
rect 11732 -3272 11756 -3238
rect 11790 -3272 11814 -3238
rect 11732 -3296 11814 -3272
rect 12750 -3238 12832 -3212
rect 12750 -3272 12774 -3238
rect 12808 -3272 12832 -3238
rect 12750 -3296 12832 -3272
rect 13768 -3238 13850 -3212
rect 13768 -3272 13792 -3238
rect 13826 -3272 13850 -3238
rect 13768 -3296 13850 -3272
rect 14786 -3238 14868 -3212
rect 14786 -3272 14810 -3238
rect 14844 -3272 14868 -3238
rect 14786 -3296 14868 -3272
rect 15804 -3238 15886 -3212
rect 15804 -3272 15828 -3238
rect 15862 -3272 15886 -3238
rect 15804 -3296 15886 -3272
rect 16822 -3238 16904 -3212
rect 16822 -3272 16846 -3238
rect 16880 -3272 16904 -3238
rect 16822 -3296 16904 -3272
rect 17840 -3238 17922 -3212
rect 17840 -3272 17864 -3238
rect 17898 -3272 17922 -3238
rect 17840 -3296 17922 -3272
rect 18858 -3238 18940 -3212
rect 18858 -3272 18882 -3238
rect 18916 -3272 18940 -3238
rect 18858 -3296 18940 -3272
rect 19876 -3238 19958 -3212
rect 19876 -3272 19900 -3238
rect 19934 -3272 19958 -3238
rect 19876 -3296 19958 -3272
rect 20894 -3238 20976 -3212
rect 20894 -3272 20918 -3238
rect 20952 -3272 20976 -3238
rect 20894 -3296 20976 -3272
rect 21912 -3238 21994 -3212
rect 21912 -3272 21936 -3238
rect 21970 -3272 21994 -3238
rect 21912 -3296 21994 -3272
rect 7266 -4516 7348 -4490
rect 7266 -4550 7290 -4516
rect 7324 -4550 7348 -4516
rect 7266 -4574 7348 -4550
rect 8284 -4516 8366 -4490
rect 8284 -4550 8308 -4516
rect 8342 -4550 8366 -4516
rect 8284 -4574 8366 -4550
rect 9302 -4516 9384 -4490
rect 9302 -4550 9326 -4516
rect 9360 -4550 9384 -4516
rect 9302 -4574 9384 -4550
rect 10320 -4516 10402 -4490
rect 10320 -4550 10344 -4516
rect 10378 -4550 10402 -4516
rect 10320 -4574 10402 -4550
rect 11338 -4516 11420 -4490
rect 11338 -4550 11362 -4516
rect 11396 -4550 11420 -4516
rect 11338 -4574 11420 -4550
rect 12356 -4516 12438 -4490
rect 12356 -4550 12380 -4516
rect 12414 -4550 12438 -4516
rect 12356 -4574 12438 -4550
rect 13374 -4516 13456 -4490
rect 13374 -4550 13398 -4516
rect 13432 -4550 13456 -4516
rect 13374 -4574 13456 -4550
rect 14392 -4516 14474 -4490
rect 14392 -4550 14416 -4516
rect 14450 -4550 14474 -4516
rect 14392 -4574 14474 -4550
rect 15410 -4516 15492 -4490
rect 15410 -4550 15434 -4516
rect 15468 -4550 15492 -4516
rect 15410 -4574 15492 -4550
rect 16428 -4516 16510 -4490
rect 16428 -4550 16452 -4516
rect 16486 -4550 16510 -4516
rect 16428 -4574 16510 -4550
rect 17446 -4516 17528 -4490
rect 17446 -4550 17470 -4516
rect 17504 -4550 17528 -4516
rect 17446 -4574 17528 -4550
rect 18464 -4516 18546 -4490
rect 18464 -4550 18488 -4516
rect 18522 -4550 18546 -4516
rect 18464 -4574 18546 -4550
rect 19482 -4516 19564 -4490
rect 19482 -4550 19506 -4516
rect 19540 -4550 19564 -4516
rect 19482 -4574 19564 -4550
rect 20500 -4516 20582 -4490
rect 20500 -4550 20524 -4516
rect 20558 -4550 20582 -4516
rect 20500 -4574 20582 -4550
rect 21518 -4516 21600 -4490
rect 21518 -4550 21542 -4516
rect 21576 -4550 21600 -4516
rect 21518 -4574 21600 -4550
rect 22536 -4516 22618 -4490
rect 22536 -4550 22560 -4516
rect 22594 -4550 22618 -4516
rect 22536 -4574 22618 -4550
rect 2668 -4826 2750 -4800
rect 2668 -4860 2692 -4826
rect 2726 -4860 2750 -4826
rect 2668 -4884 2750 -4860
rect 3686 -4826 3768 -4800
rect 3686 -4860 3710 -4826
rect 3744 -4860 3768 -4826
rect 3686 -4884 3768 -4860
rect 4704 -4826 4786 -4800
rect 4704 -4860 4728 -4826
rect 4762 -4860 4786 -4826
rect 4704 -4884 4786 -4860
rect 5722 -4826 5804 -4800
rect 5722 -4860 5746 -4826
rect 5780 -4860 5804 -4826
rect 5722 -4884 5804 -4860
rect 2144 -5980 2226 -5954
rect 2144 -6014 2168 -5980
rect 2202 -6014 2226 -5980
rect 2144 -6038 2226 -6014
rect 3162 -5980 3244 -5954
rect 3162 -6014 3186 -5980
rect 3220 -6014 3244 -5980
rect 3162 -6038 3244 -6014
rect 4180 -5980 4262 -5954
rect 4180 -6014 4204 -5980
rect 4238 -6014 4262 -5980
rect 4180 -6038 4262 -6014
rect 5198 -5980 5280 -5954
rect 5198 -6014 5222 -5980
rect 5256 -6014 5280 -5980
rect 5198 -6038 5280 -6014
rect 7356 -5964 7438 -5938
rect 7356 -5998 7380 -5964
rect 7414 -5998 7438 -5964
rect 7356 -6022 7438 -5998
rect 8374 -5964 8456 -5938
rect 8374 -5998 8398 -5964
rect 8432 -5998 8456 -5964
rect 8374 -6022 8456 -5998
rect 9392 -5964 9474 -5938
rect 9392 -5998 9416 -5964
rect 9450 -5998 9474 -5964
rect 9392 -6022 9474 -5998
rect 10410 -5964 10492 -5938
rect 10410 -5998 10434 -5964
rect 10468 -5998 10492 -5964
rect 10410 -6022 10492 -5998
rect 11428 -5964 11510 -5938
rect 11428 -5998 11452 -5964
rect 11486 -5998 11510 -5964
rect 11428 -6022 11510 -5998
rect 12446 -5964 12528 -5938
rect 12446 -5998 12470 -5964
rect 12504 -5998 12528 -5964
rect 12446 -6022 12528 -5998
rect 13464 -5964 13546 -5938
rect 13464 -5998 13488 -5964
rect 13522 -5998 13546 -5964
rect 13464 -6022 13546 -5998
rect 14482 -5964 14564 -5938
rect 14482 -5998 14506 -5964
rect 14540 -5998 14564 -5964
rect 14482 -6022 14564 -5998
rect 15500 -5964 15582 -5938
rect 15500 -5998 15524 -5964
rect 15558 -5998 15582 -5964
rect 15500 -6022 15582 -5998
rect 16518 -5964 16600 -5938
rect 16518 -5998 16542 -5964
rect 16576 -5998 16600 -5964
rect 16518 -6022 16600 -5998
rect 17536 -5964 17618 -5938
rect 17536 -5998 17560 -5964
rect 17594 -5998 17618 -5964
rect 17536 -6022 17618 -5998
rect 18554 -5964 18636 -5938
rect 18554 -5998 18578 -5964
rect 18612 -5998 18636 -5964
rect 18554 -6022 18636 -5998
rect 19572 -5964 19654 -5938
rect 19572 -5998 19596 -5964
rect 19630 -5998 19654 -5964
rect 19572 -6022 19654 -5998
rect 20590 -5964 20672 -5938
rect 20590 -5998 20614 -5964
rect 20648 -5998 20672 -5964
rect 20590 -6022 20672 -5998
rect 21608 -5964 21690 -5938
rect 21608 -5998 21632 -5964
rect 21666 -5998 21690 -5964
rect 21608 -6022 21690 -5998
rect 22626 -5964 22708 -5938
rect 22626 -5998 22650 -5964
rect 22684 -5998 22708 -5964
rect 22626 -6022 22708 -5998
rect 2154 -7008 2236 -6982
rect 2154 -7042 2178 -7008
rect 2212 -7042 2236 -7008
rect 2154 -7066 2236 -7042
rect 3172 -7008 3254 -6982
rect 3172 -7042 3196 -7008
rect 3230 -7042 3254 -7008
rect 3172 -7066 3254 -7042
rect 4190 -7008 4272 -6982
rect 4190 -7042 4214 -7008
rect 4248 -7042 4272 -7008
rect 4190 -7066 4272 -7042
rect 5208 -7008 5290 -6982
rect 5208 -7042 5232 -7008
rect 5266 -7042 5290 -7008
rect 5208 -7066 5290 -7042
rect 7380 -7232 7462 -7206
rect 7380 -7266 7404 -7232
rect 7438 -7266 7462 -7232
rect 7380 -7290 7462 -7266
rect 8398 -7232 8480 -7206
rect 8398 -7266 8422 -7232
rect 8456 -7266 8480 -7232
rect 8398 -7290 8480 -7266
rect 9416 -7232 9498 -7206
rect 9416 -7266 9440 -7232
rect 9474 -7266 9498 -7232
rect 9416 -7290 9498 -7266
rect 10434 -7232 10516 -7206
rect 10434 -7266 10458 -7232
rect 10492 -7266 10516 -7232
rect 10434 -7290 10516 -7266
rect 11452 -7232 11534 -7206
rect 11452 -7266 11476 -7232
rect 11510 -7266 11534 -7232
rect 11452 -7290 11534 -7266
rect 12470 -7232 12552 -7206
rect 12470 -7266 12494 -7232
rect 12528 -7266 12552 -7232
rect 12470 -7290 12552 -7266
rect 13488 -7232 13570 -7206
rect 13488 -7266 13512 -7232
rect 13546 -7266 13570 -7232
rect 13488 -7290 13570 -7266
rect 14506 -7232 14588 -7206
rect 14506 -7266 14530 -7232
rect 14564 -7266 14588 -7232
rect 14506 -7290 14588 -7266
rect 15524 -7232 15606 -7206
rect 15524 -7266 15548 -7232
rect 15582 -7266 15606 -7232
rect 15524 -7290 15606 -7266
rect 16542 -7232 16624 -7206
rect 16542 -7266 16566 -7232
rect 16600 -7266 16624 -7232
rect 16542 -7290 16624 -7266
rect 17560 -7232 17642 -7206
rect 17560 -7266 17584 -7232
rect 17618 -7266 17642 -7232
rect 17560 -7290 17642 -7266
rect 18578 -7232 18660 -7206
rect 18578 -7266 18602 -7232
rect 18636 -7266 18660 -7232
rect 18578 -7290 18660 -7266
rect 19596 -7232 19678 -7206
rect 19596 -7266 19620 -7232
rect 19654 -7266 19678 -7232
rect 19596 -7290 19678 -7266
rect 20614 -7232 20696 -7206
rect 20614 -7266 20638 -7232
rect 20672 -7266 20696 -7232
rect 20614 -7290 20696 -7266
rect 21632 -7232 21714 -7206
rect 21632 -7266 21656 -7232
rect 21690 -7266 21714 -7232
rect 21632 -7290 21714 -7266
rect 22650 -7232 22732 -7206
rect 22650 -7266 22674 -7232
rect 22708 -7266 22732 -7232
rect 22650 -7290 22732 -7266
rect 2144 -8036 2226 -8010
rect 2144 -8070 2168 -8036
rect 2202 -8070 2226 -8036
rect 2144 -8094 2226 -8070
rect 3162 -8036 3244 -8010
rect 3162 -8070 3186 -8036
rect 3220 -8070 3244 -8036
rect 3162 -8094 3244 -8070
rect 4180 -8036 4262 -8010
rect 4180 -8070 4204 -8036
rect 4238 -8070 4262 -8036
rect 4180 -8094 4262 -8070
rect 5198 -8036 5280 -8010
rect 5198 -8070 5222 -8036
rect 5256 -8070 5280 -8036
rect 5198 -8094 5280 -8070
rect 7244 -8476 7326 -8450
rect 7244 -8510 7268 -8476
rect 7302 -8510 7326 -8476
rect 7244 -8534 7326 -8510
rect 8262 -8476 8344 -8450
rect 8262 -8510 8286 -8476
rect 8320 -8510 8344 -8476
rect 8262 -8534 8344 -8510
rect 9280 -8476 9362 -8450
rect 9280 -8510 9304 -8476
rect 9338 -8510 9362 -8476
rect 9280 -8534 9362 -8510
rect 10298 -8476 10380 -8450
rect 10298 -8510 10322 -8476
rect 10356 -8510 10380 -8476
rect 10298 -8534 10380 -8510
rect 11316 -8476 11398 -8450
rect 11316 -8510 11340 -8476
rect 11374 -8510 11398 -8476
rect 11316 -8534 11398 -8510
rect 12334 -8476 12416 -8450
rect 12334 -8510 12358 -8476
rect 12392 -8510 12416 -8476
rect 12334 -8534 12416 -8510
rect 13352 -8476 13434 -8450
rect 13352 -8510 13376 -8476
rect 13410 -8510 13434 -8476
rect 13352 -8534 13434 -8510
rect 14370 -8476 14452 -8450
rect 14370 -8510 14394 -8476
rect 14428 -8510 14452 -8476
rect 14370 -8534 14452 -8510
rect 15388 -8476 15470 -8450
rect 15388 -8510 15412 -8476
rect 15446 -8510 15470 -8476
rect 15388 -8534 15470 -8510
rect 16406 -8476 16488 -8450
rect 16406 -8510 16430 -8476
rect 16464 -8510 16488 -8476
rect 16406 -8534 16488 -8510
rect 17424 -8476 17506 -8450
rect 17424 -8510 17448 -8476
rect 17482 -8510 17506 -8476
rect 17424 -8534 17506 -8510
rect 18442 -8476 18524 -8450
rect 18442 -8510 18466 -8476
rect 18500 -8510 18524 -8476
rect 18442 -8534 18524 -8510
rect 19460 -8476 19542 -8450
rect 19460 -8510 19484 -8476
rect 19518 -8510 19542 -8476
rect 19460 -8534 19542 -8510
rect 20478 -8476 20560 -8450
rect 20478 -8510 20502 -8476
rect 20536 -8510 20560 -8476
rect 20478 -8534 20560 -8510
rect 21496 -8476 21578 -8450
rect 21496 -8510 21520 -8476
rect 21554 -8510 21578 -8476
rect 21496 -8534 21578 -8510
rect 22514 -8476 22596 -8450
rect 22514 -8510 22538 -8476
rect 22572 -8510 22596 -8476
rect 22514 -8534 22596 -8510
rect 2668 -9188 2750 -9162
rect 2668 -9222 2692 -9188
rect 2726 -9222 2750 -9188
rect 2668 -9246 2750 -9222
rect 3686 -9188 3768 -9162
rect 3686 -9222 3710 -9188
rect 3744 -9222 3768 -9188
rect 3686 -9246 3768 -9222
rect 4704 -9188 4786 -9162
rect 4704 -9222 4728 -9188
rect 4762 -9222 4786 -9188
rect 4704 -9246 4786 -9222
rect 5722 -9188 5804 -9162
rect 5722 -9222 5746 -9188
rect 5780 -9222 5804 -9188
rect 5722 -9246 5804 -9222
rect 378 -10248 478 -10186
rect 24722 -10248 24822 -10186
rect 378 -10348 540 -10248
rect 24660 -10348 24822 -10248
<< psubdiffcont >>
rect -12160 -11278 24760 -11178
rect -12322 -27060 -12222 -11340
rect 3110 -11818 3144 -11784
rect 4128 -11818 4162 -11784
rect 5146 -11818 5180 -11784
rect 6164 -11818 6198 -11784
rect 7182 -11818 7216 -11784
rect 8200 -11818 8234 -11784
rect 9218 -11818 9252 -11784
rect 10236 -11818 10270 -11784
rect 11254 -11818 11288 -11784
rect 12272 -11818 12306 -11784
rect 13290 -11818 13324 -11784
rect 14308 -11818 14342 -11784
rect 15326 -11818 15360 -11784
rect 16344 -11818 16378 -11784
rect 17362 -11818 17396 -11784
rect 18380 -11818 18414 -11784
rect 19398 -11818 19432 -11784
rect 20416 -11818 20450 -11784
rect 21434 -11818 21468 -11784
rect 22452 -11818 22486 -11784
rect -9184 -12420 -9150 -12386
rect -8166 -12420 -8132 -12386
rect -7148 -12420 -7114 -12386
rect -6130 -12420 -6096 -12386
rect -5112 -12420 -5078 -12386
rect -4094 -12420 -4060 -12386
rect -3076 -12420 -3042 -12386
rect -2058 -12420 -2024 -12386
rect -1040 -12420 -1006 -12386
rect -12 -12420 22 -12386
rect -9184 -13238 -9150 -13204
rect -8166 -13238 -8132 -13204
rect -7148 -13238 -7114 -13204
rect -6130 -13238 -6096 -13204
rect -5112 -13238 -5078 -13204
rect -4094 -13238 -4060 -13204
rect -3076 -13238 -3042 -13204
rect -2058 -13238 -2024 -13204
rect -1040 -13238 -1006 -13204
rect -12 -13238 22 -13204
rect 3122 -13844 3156 -13810
rect 4140 -13844 4174 -13810
rect 5158 -13844 5192 -13810
rect 6176 -13844 6210 -13810
rect 7194 -13844 7228 -13810
rect 8212 -13844 8246 -13810
rect 9230 -13844 9264 -13810
rect 10248 -13844 10282 -13810
rect 11266 -13844 11300 -13810
rect 12284 -13844 12318 -13810
rect 13302 -13844 13336 -13810
rect 14320 -13844 14354 -13810
rect 15338 -13844 15372 -13810
rect 16356 -13844 16390 -13810
rect 17374 -13844 17408 -13810
rect 18392 -13844 18426 -13810
rect 19410 -13844 19444 -13810
rect 20428 -13844 20462 -13810
rect 21446 -13844 21480 -13810
rect 22464 -13844 22498 -13810
rect -9184 -14056 -9150 -14022
rect -8166 -14056 -8132 -14022
rect -7148 -14056 -7114 -14022
rect -6130 -14056 -6096 -14022
rect -5112 -14056 -5078 -14022
rect -4094 -14056 -4060 -14022
rect -3076 -14056 -3042 -14022
rect -2058 -14056 -2024 -14022
rect -1040 -14056 -1006 -14022
rect -12 -14056 22 -14022
rect -9184 -14874 -9150 -14840
rect -8166 -14874 -8132 -14840
rect -7148 -14874 -7114 -14840
rect -6130 -14874 -6096 -14840
rect -5112 -14874 -5078 -14840
rect -4094 -14874 -4060 -14840
rect -3076 -14874 -3042 -14840
rect -2058 -14874 -2024 -14840
rect -1040 -14874 -1006 -14840
rect -12 -14874 22 -14840
rect 3110 -15150 3144 -15116
rect 4128 -15150 4162 -15116
rect 5146 -15150 5180 -15116
rect 6164 -15150 6198 -15116
rect 7182 -15150 7216 -15116
rect 8200 -15150 8234 -15116
rect 9218 -15150 9252 -15116
rect 10236 -15150 10270 -15116
rect 11254 -15150 11288 -15116
rect 12272 -15150 12306 -15116
rect 13290 -15150 13324 -15116
rect 14308 -15150 14342 -15116
rect 15326 -15150 15360 -15116
rect 16344 -15150 16378 -15116
rect 17362 -15150 17396 -15116
rect 18380 -15150 18414 -15116
rect 19398 -15150 19432 -15116
rect 20416 -15150 20450 -15116
rect 21434 -15150 21468 -15116
rect 22452 -15150 22486 -15116
rect -9184 -15692 -9150 -15658
rect -8166 -15692 -8132 -15658
rect -7148 -15692 -7114 -15658
rect -6130 -15692 -6096 -15658
rect -5112 -15692 -5078 -15658
rect -4094 -15692 -4060 -15658
rect -3076 -15692 -3042 -15658
rect -2058 -15692 -2024 -15658
rect -1040 -15692 -1006 -15658
rect -12 -15692 22 -15658
rect -9184 -16510 -9150 -16476
rect -8166 -16510 -8132 -16476
rect -7148 -16510 -7114 -16476
rect -6130 -16510 -6096 -16476
rect -5112 -16510 -5078 -16476
rect -4094 -16510 -4060 -16476
rect -3076 -16510 -3042 -16476
rect 3098 -16386 3132 -16352
rect 4116 -16386 4150 -16352
rect 5134 -16386 5168 -16352
rect 6152 -16386 6186 -16352
rect 7170 -16386 7204 -16352
rect 8188 -16386 8222 -16352
rect 9206 -16386 9240 -16352
rect 10224 -16386 10258 -16352
rect 11242 -16386 11276 -16352
rect 12260 -16386 12294 -16352
rect 13278 -16386 13312 -16352
rect 14296 -16386 14330 -16352
rect 15314 -16386 15348 -16352
rect 16332 -16386 16366 -16352
rect 17350 -16386 17384 -16352
rect 18368 -16386 18402 -16352
rect 19386 -16386 19420 -16352
rect 20404 -16386 20438 -16352
rect 21422 -16386 21456 -16352
rect 22440 -16386 22474 -16352
rect -2058 -16510 -2024 -16476
rect -1040 -16510 -1006 -16476
rect -12 -16510 22 -16476
rect -9184 -17328 -9150 -17294
rect -8166 -17328 -8132 -17294
rect -7148 -17328 -7114 -17294
rect -6130 -17328 -6096 -17294
rect -5112 -17328 -5078 -17294
rect -4094 -17328 -4060 -17294
rect -3076 -17328 -3042 -17294
rect -2058 -17328 -2024 -17294
rect -1040 -17328 -1006 -17294
rect -12 -17328 22 -17294
rect 3098 -17610 3132 -17576
rect 4116 -17610 4150 -17576
rect 5134 -17610 5168 -17576
rect 6152 -17610 6186 -17576
rect 7170 -17610 7204 -17576
rect 8188 -17610 8222 -17576
rect 9206 -17610 9240 -17576
rect 10224 -17610 10258 -17576
rect 11242 -17610 11276 -17576
rect 12260 -17610 12294 -17576
rect 13278 -17610 13312 -17576
rect 14296 -17610 14330 -17576
rect 15314 -17610 15348 -17576
rect 16332 -17610 16366 -17576
rect 17350 -17610 17384 -17576
rect 18368 -17610 18402 -17576
rect 19386 -17610 19420 -17576
rect 20404 -17610 20438 -17576
rect 21422 -17610 21456 -17576
rect 22440 -17610 22474 -17576
rect -9184 -18146 -9150 -18112
rect -8166 -18146 -8132 -18112
rect -7148 -18146 -7114 -18112
rect -6130 -18146 -6096 -18112
rect -5112 -18146 -5078 -18112
rect -4094 -18146 -4060 -18112
rect -3076 -18146 -3042 -18112
rect -2058 -18146 -2024 -18112
rect -1040 -18146 -1006 -18112
rect -12 -18146 22 -18112
rect 3110 -18846 3144 -18812
rect 4128 -18846 4162 -18812
rect 5146 -18846 5180 -18812
rect 6164 -18846 6198 -18812
rect 7182 -18846 7216 -18812
rect 8200 -18846 8234 -18812
rect 9218 -18846 9252 -18812
rect 10236 -18846 10270 -18812
rect 11254 -18846 11288 -18812
rect 12272 -18846 12306 -18812
rect 13290 -18846 13324 -18812
rect 14308 -18846 14342 -18812
rect 15326 -18846 15360 -18812
rect 16344 -18846 16378 -18812
rect 17362 -18846 17396 -18812
rect 18380 -18846 18414 -18812
rect 19398 -18846 19432 -18812
rect 20416 -18846 20450 -18812
rect 21434 -18846 21468 -18812
rect 22452 -18846 22486 -18812
rect -9196 -19040 -9162 -19006
rect -8178 -19040 -8144 -19006
rect -7160 -19040 -7126 -19006
rect -6142 -19040 -6108 -19006
rect -5124 -19040 -5090 -19006
rect -4106 -19040 -4072 -19006
rect -3088 -19040 -3054 -19006
rect -2070 -19040 -2036 -19006
rect -1052 -19040 -1018 -19006
rect -24 -19040 10 -19006
rect -9992 -19988 -9958 -19954
rect -8974 -19988 -8940 -19954
rect -7956 -19988 -7922 -19954
rect -6938 -19988 -6904 -19954
rect -5920 -19988 -5886 -19954
rect -4902 -19988 -4868 -19954
rect -3884 -19988 -3850 -19954
rect -2866 -19988 -2832 -19954
rect -1848 -19988 -1814 -19954
rect -830 -19988 -796 -19954
rect 188 -19988 222 -19954
rect 3110 -20094 3144 -20060
rect 4128 -20094 4162 -20060
rect 5146 -20094 5180 -20060
rect 6164 -20094 6198 -20060
rect 7182 -20094 7216 -20060
rect 8200 -20094 8234 -20060
rect 9218 -20094 9252 -20060
rect 10236 -20094 10270 -20060
rect 11254 -20094 11288 -20060
rect 12272 -20094 12306 -20060
rect 13290 -20094 13324 -20060
rect 14308 -20094 14342 -20060
rect 15326 -20094 15360 -20060
rect 16344 -20094 16378 -20060
rect 17362 -20094 17396 -20060
rect 18380 -20094 18414 -20060
rect 19398 -20094 19432 -20060
rect 20416 -20094 20450 -20060
rect 21434 -20094 21468 -20060
rect 22452 -20094 22486 -20060
rect -9980 -21130 -9946 -21096
rect -8962 -21130 -8928 -21096
rect -7944 -21130 -7910 -21096
rect -6926 -21130 -6892 -21096
rect -5908 -21130 -5874 -21096
rect -4890 -21130 -4856 -21096
rect -3872 -21130 -3838 -21096
rect -2854 -21130 -2820 -21096
rect -1836 -21130 -1802 -21096
rect -818 -21130 -784 -21096
rect 200 -21130 234 -21096
rect 3086 -21330 3120 -21296
rect 4104 -21330 4138 -21296
rect 5122 -21330 5156 -21296
rect 6140 -21330 6174 -21296
rect 7158 -21330 7192 -21296
rect 8176 -21330 8210 -21296
rect 9194 -21330 9228 -21296
rect 10212 -21330 10246 -21296
rect 11230 -21330 11264 -21296
rect 12248 -21330 12282 -21296
rect 13266 -21330 13300 -21296
rect 14284 -21330 14318 -21296
rect 15302 -21330 15336 -21296
rect 16320 -21330 16354 -21296
rect 17338 -21330 17372 -21296
rect 18356 -21330 18390 -21296
rect 19374 -21330 19408 -21296
rect 20392 -21330 20426 -21296
rect 21410 -21330 21444 -21296
rect 22428 -21330 22462 -21296
rect -10002 -22238 -9968 -22204
rect -8984 -22238 -8950 -22204
rect -7966 -22238 -7932 -22204
rect -6948 -22238 -6914 -22204
rect -5930 -22238 -5896 -22204
rect -4912 -22238 -4878 -22204
rect -3894 -22238 -3860 -22204
rect -2876 -22238 -2842 -22204
rect -1858 -22238 -1824 -22204
rect -840 -22238 -806 -22204
rect 178 -22238 212 -22204
rect 3098 -22554 3132 -22520
rect 4116 -22554 4150 -22520
rect 5134 -22554 5168 -22520
rect 6152 -22554 6186 -22520
rect 7170 -22554 7204 -22520
rect 8188 -22554 8222 -22520
rect 9206 -22554 9240 -22520
rect 10224 -22554 10258 -22520
rect 11242 -22554 11276 -22520
rect 12260 -22554 12294 -22520
rect 13278 -22554 13312 -22520
rect 14296 -22554 14330 -22520
rect 15314 -22554 15348 -22520
rect 16332 -22554 16366 -22520
rect 17350 -22554 17384 -22520
rect 18368 -22554 18402 -22520
rect 19386 -22554 19420 -22520
rect 20404 -22554 20438 -22520
rect 21422 -22554 21456 -22520
rect 22440 -22554 22474 -22520
rect -10002 -23344 -9968 -23310
rect -8984 -23344 -8950 -23310
rect -7966 -23344 -7932 -23310
rect -6948 -23344 -6914 -23310
rect -5930 -23344 -5896 -23310
rect -4912 -23344 -4878 -23310
rect -3894 -23344 -3860 -23310
rect -2876 -23344 -2842 -23310
rect -1858 -23344 -1824 -23310
rect -840 -23344 -806 -23310
rect 178 -23344 212 -23310
rect 3098 -23790 3132 -23756
rect 4116 -23790 4150 -23756
rect 5134 -23790 5168 -23756
rect 6152 -23790 6186 -23756
rect 7170 -23790 7204 -23756
rect 8188 -23790 8222 -23756
rect 9206 -23790 9240 -23756
rect 10224 -23790 10258 -23756
rect 11242 -23790 11276 -23756
rect 12260 -23790 12294 -23756
rect 13278 -23790 13312 -23756
rect 14296 -23790 14330 -23756
rect 15314 -23790 15348 -23756
rect 16332 -23790 16366 -23756
rect 17350 -23790 17384 -23756
rect 18368 -23790 18402 -23756
rect 19386 -23790 19420 -23756
rect 20404 -23790 20438 -23756
rect 21422 -23790 21456 -23756
rect 22440 -23790 22474 -23756
rect -10002 -24686 -9968 -24652
rect -8984 -24686 -8950 -24652
rect -7966 -24686 -7932 -24652
rect -6948 -24686 -6914 -24652
rect -5930 -24686 -5896 -24652
rect -4912 -24686 -4878 -24652
rect -3894 -24686 -3860 -24652
rect -2876 -24686 -2842 -24652
rect -1858 -24686 -1824 -24652
rect -840 -24686 -806 -24652
rect 178 -24686 212 -24652
rect 3110 -25036 3144 -25002
rect 4128 -25036 4162 -25002
rect 5146 -25036 5180 -25002
rect 6164 -25036 6198 -25002
rect 7182 -25036 7216 -25002
rect 8200 -25036 8234 -25002
rect 9218 -25036 9252 -25002
rect 10236 -25036 10270 -25002
rect 11254 -25036 11288 -25002
rect 12272 -25036 12306 -25002
rect 13290 -25036 13324 -25002
rect 14308 -25036 14342 -25002
rect 15326 -25036 15360 -25002
rect 16344 -25036 16378 -25002
rect 17362 -25036 17396 -25002
rect 18380 -25036 18414 -25002
rect 19398 -25036 19432 -25002
rect 20416 -25036 20450 -25002
rect 21434 -25036 21468 -25002
rect 22452 -25036 22486 -25002
rect -10192 -26132 -10158 -26098
rect -9174 -26132 -9140 -26098
rect -8156 -26132 -8122 -26098
rect -7138 -26132 -7104 -26098
rect -6120 -26132 -6086 -26098
rect -5102 -26132 -5068 -26098
rect -4084 -26132 -4050 -26098
rect -3066 -26132 -3032 -26098
rect -2048 -26132 -2014 -26098
rect -1030 -26132 -996 -26098
rect -12 -26132 22 -26098
rect 3098 -26214 3132 -26180
rect 4116 -26214 4150 -26180
rect 5134 -26214 5168 -26180
rect 6152 -26214 6186 -26180
rect 7170 -26214 7204 -26180
rect 8188 -26214 8222 -26180
rect 9206 -26214 9240 -26180
rect 10224 -26214 10258 -26180
rect 11242 -26214 11276 -26180
rect 12260 -26214 12294 -26180
rect 13278 -26214 13312 -26180
rect 14296 -26214 14330 -26180
rect 15314 -26214 15348 -26180
rect 16332 -26214 16366 -26180
rect 17350 -26214 17384 -26180
rect 18368 -26214 18402 -26180
rect 19386 -26214 19420 -26180
rect 20404 -26214 20438 -26180
rect 21422 -26214 21456 -26180
rect 22440 -26214 22474 -26180
rect 24822 -27060 24922 -11340
rect -12160 -27222 24760 -27122
<< nsubdiffcont >>
rect 540 4222 24660 4322
rect 378 -10186 478 4160
rect 6996 1744 7030 1778
rect 8014 1744 8048 1778
rect 9032 1744 9066 1778
rect 10050 1744 10084 1778
rect 11068 1744 11102 1778
rect 12086 1744 12120 1778
rect 13104 1744 13138 1778
rect 14122 1744 14156 1778
rect 15140 1744 15174 1778
rect 16158 1744 16192 1778
rect 17176 1744 17210 1778
rect 18194 1744 18228 1778
rect 19212 1744 19246 1778
rect 20230 1744 20264 1778
rect 21248 1744 21282 1778
rect 22266 1744 22300 1778
rect 7018 590 7052 624
rect 8036 590 8070 624
rect 9054 590 9088 624
rect 10072 590 10106 624
rect 11090 590 11124 624
rect 12108 590 12142 624
rect 13126 590 13160 624
rect 14144 590 14178 624
rect 15162 590 15196 624
rect 16180 590 16214 624
rect 17198 590 17232 624
rect 18216 590 18250 624
rect 19234 590 19268 624
rect 20252 590 20286 624
rect 21270 590 21304 624
rect 22288 590 22322 624
rect 6996 -542 7030 -508
rect 8014 -542 8048 -508
rect 9032 -542 9066 -508
rect 10050 -542 10084 -508
rect 11068 -542 11102 -508
rect 12086 -542 12120 -508
rect 13104 -542 13138 -508
rect 14122 -542 14156 -508
rect 15140 -542 15174 -508
rect 16158 -542 16192 -508
rect 17176 -542 17210 -508
rect 18194 -542 18228 -508
rect 19212 -542 19246 -508
rect 20230 -542 20264 -508
rect 21248 -542 21282 -508
rect 22266 -542 22300 -508
rect 6996 -1924 7030 -1890
rect 8014 -1924 8048 -1890
rect 9032 -1924 9066 -1890
rect 10050 -1924 10084 -1890
rect 11068 -1924 11102 -1890
rect 12086 -1924 12120 -1890
rect 13104 -1924 13138 -1890
rect 14122 -1924 14156 -1890
rect 15140 -1924 15174 -1890
rect 16158 -1924 16192 -1890
rect 17176 -1924 17210 -1890
rect 18194 -1924 18228 -1890
rect 19212 -1924 19246 -1890
rect 20230 -1924 20264 -1890
rect 21248 -1924 21282 -1890
rect 22266 -1924 22300 -1890
rect 7684 -3272 7718 -3238
rect 8702 -3272 8736 -3238
rect 9720 -3272 9754 -3238
rect 10738 -3272 10772 -3238
rect 11756 -3272 11790 -3238
rect 12774 -3272 12808 -3238
rect 13792 -3272 13826 -3238
rect 14810 -3272 14844 -3238
rect 15828 -3272 15862 -3238
rect 16846 -3272 16880 -3238
rect 17864 -3272 17898 -3238
rect 18882 -3272 18916 -3238
rect 19900 -3272 19934 -3238
rect 20918 -3272 20952 -3238
rect 21936 -3272 21970 -3238
rect 7290 -4550 7324 -4516
rect 8308 -4550 8342 -4516
rect 9326 -4550 9360 -4516
rect 10344 -4550 10378 -4516
rect 11362 -4550 11396 -4516
rect 12380 -4550 12414 -4516
rect 13398 -4550 13432 -4516
rect 14416 -4550 14450 -4516
rect 15434 -4550 15468 -4516
rect 16452 -4550 16486 -4516
rect 17470 -4550 17504 -4516
rect 18488 -4550 18522 -4516
rect 19506 -4550 19540 -4516
rect 20524 -4550 20558 -4516
rect 21542 -4550 21576 -4516
rect 22560 -4550 22594 -4516
rect 2692 -4860 2726 -4826
rect 3710 -4860 3744 -4826
rect 4728 -4860 4762 -4826
rect 5746 -4860 5780 -4826
rect 2168 -6014 2202 -5980
rect 3186 -6014 3220 -5980
rect 4204 -6014 4238 -5980
rect 5222 -6014 5256 -5980
rect 7380 -5998 7414 -5964
rect 8398 -5998 8432 -5964
rect 9416 -5998 9450 -5964
rect 10434 -5998 10468 -5964
rect 11452 -5998 11486 -5964
rect 12470 -5998 12504 -5964
rect 13488 -5998 13522 -5964
rect 14506 -5998 14540 -5964
rect 15524 -5998 15558 -5964
rect 16542 -5998 16576 -5964
rect 17560 -5998 17594 -5964
rect 18578 -5998 18612 -5964
rect 19596 -5998 19630 -5964
rect 20614 -5998 20648 -5964
rect 21632 -5998 21666 -5964
rect 22650 -5998 22684 -5964
rect 2178 -7042 2212 -7008
rect 3196 -7042 3230 -7008
rect 4214 -7042 4248 -7008
rect 5232 -7042 5266 -7008
rect 7404 -7266 7438 -7232
rect 8422 -7266 8456 -7232
rect 9440 -7266 9474 -7232
rect 10458 -7266 10492 -7232
rect 11476 -7266 11510 -7232
rect 12494 -7266 12528 -7232
rect 13512 -7266 13546 -7232
rect 14530 -7266 14564 -7232
rect 15548 -7266 15582 -7232
rect 16566 -7266 16600 -7232
rect 17584 -7266 17618 -7232
rect 18602 -7266 18636 -7232
rect 19620 -7266 19654 -7232
rect 20638 -7266 20672 -7232
rect 21656 -7266 21690 -7232
rect 22674 -7266 22708 -7232
rect 2168 -8070 2202 -8036
rect 3186 -8070 3220 -8036
rect 4204 -8070 4238 -8036
rect 5222 -8070 5256 -8036
rect 7268 -8510 7302 -8476
rect 8286 -8510 8320 -8476
rect 9304 -8510 9338 -8476
rect 10322 -8510 10356 -8476
rect 11340 -8510 11374 -8476
rect 12358 -8510 12392 -8476
rect 13376 -8510 13410 -8476
rect 14394 -8510 14428 -8476
rect 15412 -8510 15446 -8476
rect 16430 -8510 16464 -8476
rect 17448 -8510 17482 -8476
rect 18466 -8510 18500 -8476
rect 19484 -8510 19518 -8476
rect 20502 -8510 20536 -8476
rect 21520 -8510 21554 -8476
rect 22538 -8510 22572 -8476
rect 2692 -9222 2726 -9188
rect 3710 -9222 3744 -9188
rect 4728 -9222 4762 -9188
rect 5746 -9222 5780 -9188
rect 24722 -10186 24822 4160
rect 540 -10348 24660 -10248
<< poly >>
rect 6720 1555 7308 1571
rect 6720 1538 6736 1555
rect 6534 1521 6736 1538
rect 7292 1538 7308 1555
rect 7738 1555 8326 1571
rect 7738 1538 7754 1555
rect 7292 1521 7494 1538
rect 6534 1474 7494 1521
rect 7552 1521 7754 1538
rect 8310 1538 8326 1555
rect 8756 1555 9344 1571
rect 8756 1538 8772 1555
rect 8310 1521 8512 1538
rect 7552 1474 8512 1521
rect 8570 1521 8772 1538
rect 9328 1538 9344 1555
rect 9774 1555 10362 1571
rect 9774 1538 9790 1555
rect 9328 1521 9530 1538
rect 8570 1474 9530 1521
rect 9588 1521 9790 1538
rect 10346 1538 10362 1555
rect 10792 1555 11380 1571
rect 10792 1538 10808 1555
rect 10346 1521 10548 1538
rect 9588 1474 10548 1521
rect 10606 1521 10808 1538
rect 11364 1538 11380 1555
rect 11810 1555 12398 1571
rect 11810 1538 11826 1555
rect 11364 1521 11566 1538
rect 10606 1474 11566 1521
rect 11624 1521 11826 1538
rect 12382 1538 12398 1555
rect 12828 1555 13416 1571
rect 12828 1538 12844 1555
rect 12382 1521 12584 1538
rect 11624 1474 12584 1521
rect 12642 1521 12844 1538
rect 13400 1538 13416 1555
rect 13846 1555 14434 1571
rect 13846 1538 13862 1555
rect 13400 1521 13602 1538
rect 12642 1474 13602 1521
rect 13660 1521 13862 1538
rect 14418 1538 14434 1555
rect 14864 1555 15452 1571
rect 14864 1538 14880 1555
rect 14418 1521 14620 1538
rect 13660 1474 14620 1521
rect 14678 1521 14880 1538
rect 15436 1538 15452 1555
rect 15882 1555 16470 1571
rect 15882 1538 15898 1555
rect 15436 1521 15638 1538
rect 14678 1474 15638 1521
rect 15696 1521 15898 1538
rect 16454 1538 16470 1555
rect 16900 1555 17488 1571
rect 16900 1538 16916 1555
rect 16454 1521 16656 1538
rect 15696 1474 16656 1521
rect 16714 1521 16916 1538
rect 17472 1538 17488 1555
rect 17918 1555 18506 1571
rect 17918 1538 17934 1555
rect 17472 1521 17674 1538
rect 16714 1474 17674 1521
rect 17732 1521 17934 1538
rect 18490 1538 18506 1555
rect 18936 1555 19524 1571
rect 18936 1538 18952 1555
rect 18490 1521 18692 1538
rect 17732 1474 18692 1521
rect 18750 1521 18952 1538
rect 19508 1538 19524 1555
rect 19954 1555 20542 1571
rect 19954 1538 19970 1555
rect 19508 1521 19710 1538
rect 18750 1474 19710 1521
rect 19768 1521 19970 1538
rect 20526 1538 20542 1555
rect 20972 1555 21560 1571
rect 20972 1538 20988 1555
rect 20526 1521 20728 1538
rect 19768 1474 20728 1521
rect 20786 1521 20988 1538
rect 21544 1538 21560 1555
rect 21990 1555 22578 1571
rect 21990 1538 22006 1555
rect 21544 1521 21746 1538
rect 20786 1474 21746 1521
rect 21804 1521 22006 1538
rect 22562 1538 22578 1555
rect 22562 1521 22764 1538
rect 21804 1474 22764 1521
rect 6534 827 7494 874
rect 6534 810 6736 827
rect 6720 793 6736 810
rect 7292 810 7494 827
rect 7552 827 8512 874
rect 7552 810 7754 827
rect 7292 793 7308 810
rect 6720 777 7308 793
rect 7738 793 7754 810
rect 8310 810 8512 827
rect 8570 827 9530 874
rect 8570 810 8772 827
rect 8310 793 8326 810
rect 7738 777 8326 793
rect 8756 793 8772 810
rect 9328 810 9530 827
rect 9588 827 10548 874
rect 9588 810 9790 827
rect 9328 793 9344 810
rect 8756 777 9344 793
rect 9774 793 9790 810
rect 10346 810 10548 827
rect 10606 827 11566 874
rect 10606 810 10808 827
rect 10346 793 10362 810
rect 9774 777 10362 793
rect 10792 793 10808 810
rect 11364 810 11566 827
rect 11624 827 12584 874
rect 11624 810 11826 827
rect 11364 793 11380 810
rect 10792 777 11380 793
rect 11810 793 11826 810
rect 12382 810 12584 827
rect 12642 827 13602 874
rect 12642 810 12844 827
rect 12382 793 12398 810
rect 11810 777 12398 793
rect 12828 793 12844 810
rect 13400 810 13602 827
rect 13660 827 14620 874
rect 13660 810 13862 827
rect 13400 793 13416 810
rect 12828 777 13416 793
rect 13846 793 13862 810
rect 14418 810 14620 827
rect 14678 827 15638 874
rect 14678 810 14880 827
rect 14418 793 14434 810
rect 13846 777 14434 793
rect 14864 793 14880 810
rect 15436 810 15638 827
rect 15696 827 16656 874
rect 15696 810 15898 827
rect 15436 793 15452 810
rect 14864 777 15452 793
rect 15882 793 15898 810
rect 16454 810 16656 827
rect 16714 827 17674 874
rect 16714 810 16916 827
rect 16454 793 16470 810
rect 15882 777 16470 793
rect 16900 793 16916 810
rect 17472 810 17674 827
rect 17732 827 18692 874
rect 17732 810 17934 827
rect 17472 793 17488 810
rect 16900 777 17488 793
rect 17918 793 17934 810
rect 18490 810 18692 827
rect 18750 827 19710 874
rect 18750 810 18952 827
rect 18490 793 18506 810
rect 17918 777 18506 793
rect 18936 793 18952 810
rect 19508 810 19710 827
rect 19768 827 20728 874
rect 19768 810 19970 827
rect 19508 793 19524 810
rect 18936 777 19524 793
rect 19954 793 19970 810
rect 20526 810 20728 827
rect 20786 827 21746 874
rect 20786 810 20988 827
rect 20526 793 20542 810
rect 19954 777 20542 793
rect 20972 793 20988 810
rect 21544 810 21746 827
rect 21804 827 22764 874
rect 21804 810 22006 827
rect 21544 793 21560 810
rect 20972 777 21560 793
rect 21990 793 22006 810
rect 22562 810 22764 827
rect 22562 793 22578 810
rect 21990 777 22578 793
rect 6720 419 7308 435
rect 6720 402 6736 419
rect 6534 385 6736 402
rect 7292 402 7308 419
rect 7738 419 8326 435
rect 7738 402 7754 419
rect 7292 385 7494 402
rect 6534 338 7494 385
rect 7552 385 7754 402
rect 8310 402 8326 419
rect 8756 419 9344 435
rect 8756 402 8772 419
rect 8310 385 8512 402
rect 7552 338 8512 385
rect 8570 385 8772 402
rect 9328 402 9344 419
rect 9774 419 10362 435
rect 9774 402 9790 419
rect 9328 385 9530 402
rect 8570 338 9530 385
rect 9588 385 9790 402
rect 10346 402 10362 419
rect 10792 419 11380 435
rect 10792 402 10808 419
rect 10346 385 10548 402
rect 9588 338 10548 385
rect 10606 385 10808 402
rect 11364 402 11380 419
rect 11810 419 12398 435
rect 11810 402 11826 419
rect 11364 385 11566 402
rect 10606 338 11566 385
rect 11624 385 11826 402
rect 12382 402 12398 419
rect 12828 419 13416 435
rect 12828 402 12844 419
rect 12382 385 12584 402
rect 11624 338 12584 385
rect 12642 385 12844 402
rect 13400 402 13416 419
rect 13846 419 14434 435
rect 13846 402 13862 419
rect 13400 385 13602 402
rect 12642 338 13602 385
rect 13660 385 13862 402
rect 14418 402 14434 419
rect 14864 419 15452 435
rect 14864 402 14880 419
rect 14418 385 14620 402
rect 13660 338 14620 385
rect 14678 385 14880 402
rect 15436 402 15452 419
rect 15882 419 16470 435
rect 15882 402 15898 419
rect 15436 385 15638 402
rect 14678 338 15638 385
rect 15696 385 15898 402
rect 16454 402 16470 419
rect 16900 419 17488 435
rect 16900 402 16916 419
rect 16454 385 16656 402
rect 15696 338 16656 385
rect 16714 385 16916 402
rect 17472 402 17488 419
rect 17918 419 18506 435
rect 17918 402 17934 419
rect 17472 385 17674 402
rect 16714 338 17674 385
rect 17732 385 17934 402
rect 18490 402 18506 419
rect 18936 419 19524 435
rect 18936 402 18952 419
rect 18490 385 18692 402
rect 17732 338 18692 385
rect 18750 385 18952 402
rect 19508 402 19524 419
rect 19954 419 20542 435
rect 19954 402 19970 419
rect 19508 385 19710 402
rect 18750 338 19710 385
rect 19768 385 19970 402
rect 20526 402 20542 419
rect 20972 419 21560 435
rect 20972 402 20988 419
rect 20526 385 20728 402
rect 19768 338 20728 385
rect 20786 385 20988 402
rect 21544 402 21560 419
rect 21990 419 22578 435
rect 21990 402 22006 419
rect 21544 385 21746 402
rect 20786 338 21746 385
rect 21804 385 22006 402
rect 22562 402 22578 419
rect 22562 385 22764 402
rect 21804 338 22764 385
rect 6534 -309 7494 -262
rect 6534 -326 6736 -309
rect 6720 -343 6736 -326
rect 7292 -326 7494 -309
rect 7552 -309 8512 -262
rect 7552 -326 7754 -309
rect 7292 -343 7308 -326
rect 6720 -359 7308 -343
rect 7738 -343 7754 -326
rect 8310 -326 8512 -309
rect 8570 -309 9530 -262
rect 8570 -326 8772 -309
rect 8310 -343 8326 -326
rect 7738 -359 8326 -343
rect 8756 -343 8772 -326
rect 9328 -326 9530 -309
rect 9588 -309 10548 -262
rect 9588 -326 9790 -309
rect 9328 -343 9344 -326
rect 8756 -359 9344 -343
rect 9774 -343 9790 -326
rect 10346 -326 10548 -309
rect 10606 -309 11566 -262
rect 10606 -326 10808 -309
rect 10346 -343 10362 -326
rect 9774 -359 10362 -343
rect 10792 -343 10808 -326
rect 11364 -326 11566 -309
rect 11624 -309 12584 -262
rect 11624 -326 11826 -309
rect 11364 -343 11380 -326
rect 10792 -359 11380 -343
rect 11810 -343 11826 -326
rect 12382 -326 12584 -309
rect 12642 -309 13602 -262
rect 12642 -326 12844 -309
rect 12382 -343 12398 -326
rect 11810 -359 12398 -343
rect 12828 -343 12844 -326
rect 13400 -326 13602 -309
rect 13660 -309 14620 -262
rect 13660 -326 13862 -309
rect 13400 -343 13416 -326
rect 12828 -359 13416 -343
rect 13846 -343 13862 -326
rect 14418 -326 14620 -309
rect 14678 -309 15638 -262
rect 14678 -326 14880 -309
rect 14418 -343 14434 -326
rect 13846 -359 14434 -343
rect 14864 -343 14880 -326
rect 15436 -326 15638 -309
rect 15696 -309 16656 -262
rect 15696 -326 15898 -309
rect 15436 -343 15452 -326
rect 14864 -359 15452 -343
rect 15882 -343 15898 -326
rect 16454 -326 16656 -309
rect 16714 -309 17674 -262
rect 16714 -326 16916 -309
rect 16454 -343 16470 -326
rect 15882 -359 16470 -343
rect 16900 -343 16916 -326
rect 17472 -326 17674 -309
rect 17732 -309 18692 -262
rect 17732 -326 17934 -309
rect 17472 -343 17488 -326
rect 16900 -359 17488 -343
rect 17918 -343 17934 -326
rect 18490 -326 18692 -309
rect 18750 -309 19710 -262
rect 18750 -326 18952 -309
rect 18490 -343 18506 -326
rect 17918 -359 18506 -343
rect 18936 -343 18952 -326
rect 19508 -326 19710 -309
rect 19768 -309 20728 -262
rect 19768 -326 19970 -309
rect 19508 -343 19524 -326
rect 18936 -359 19524 -343
rect 19954 -343 19970 -326
rect 20526 -326 20728 -309
rect 20786 -309 21746 -262
rect 20786 -326 20988 -309
rect 20526 -343 20542 -326
rect 19954 -359 20542 -343
rect 20972 -343 20988 -326
rect 21544 -326 21746 -309
rect 21804 -309 22764 -262
rect 21804 -326 22006 -309
rect 21544 -343 21560 -326
rect 20972 -359 21560 -343
rect 21990 -343 22006 -326
rect 22562 -326 22764 -309
rect 22562 -343 22578 -326
rect 21990 -359 22578 -343
rect 6720 -717 7308 -701
rect 6720 -734 6736 -717
rect 6534 -751 6736 -734
rect 7292 -734 7308 -717
rect 7738 -717 8326 -701
rect 7738 -734 7754 -717
rect 7292 -751 7494 -734
rect 6534 -798 7494 -751
rect 7552 -751 7754 -734
rect 8310 -734 8326 -717
rect 8756 -717 9344 -701
rect 8756 -734 8772 -717
rect 8310 -751 8512 -734
rect 7552 -798 8512 -751
rect 8570 -751 8772 -734
rect 9328 -734 9344 -717
rect 9774 -717 10362 -701
rect 9774 -734 9790 -717
rect 9328 -751 9530 -734
rect 8570 -798 9530 -751
rect 9588 -751 9790 -734
rect 10346 -734 10362 -717
rect 10792 -717 11380 -701
rect 10792 -734 10808 -717
rect 10346 -751 10548 -734
rect 9588 -798 10548 -751
rect 10606 -751 10808 -734
rect 11364 -734 11380 -717
rect 11810 -717 12398 -701
rect 11810 -734 11826 -717
rect 11364 -751 11566 -734
rect 10606 -798 11566 -751
rect 11624 -751 11826 -734
rect 12382 -734 12398 -717
rect 12828 -717 13416 -701
rect 12828 -734 12844 -717
rect 12382 -751 12584 -734
rect 11624 -798 12584 -751
rect 12642 -751 12844 -734
rect 13400 -734 13416 -717
rect 13846 -717 14434 -701
rect 13846 -734 13862 -717
rect 13400 -751 13602 -734
rect 12642 -798 13602 -751
rect 13660 -751 13862 -734
rect 14418 -734 14434 -717
rect 14864 -717 15452 -701
rect 14864 -734 14880 -717
rect 14418 -751 14620 -734
rect 13660 -798 14620 -751
rect 14678 -751 14880 -734
rect 15436 -734 15452 -717
rect 15882 -717 16470 -701
rect 15882 -734 15898 -717
rect 15436 -751 15638 -734
rect 14678 -798 15638 -751
rect 15696 -751 15898 -734
rect 16454 -734 16470 -717
rect 16900 -717 17488 -701
rect 16900 -734 16916 -717
rect 16454 -751 16656 -734
rect 15696 -798 16656 -751
rect 16714 -751 16916 -734
rect 17472 -734 17488 -717
rect 17918 -717 18506 -701
rect 17918 -734 17934 -717
rect 17472 -751 17674 -734
rect 16714 -798 17674 -751
rect 17732 -751 17934 -734
rect 18490 -734 18506 -717
rect 18936 -717 19524 -701
rect 18936 -734 18952 -717
rect 18490 -751 18692 -734
rect 17732 -798 18692 -751
rect 18750 -751 18952 -734
rect 19508 -734 19524 -717
rect 19954 -717 20542 -701
rect 19954 -734 19970 -717
rect 19508 -751 19710 -734
rect 18750 -798 19710 -751
rect 19768 -751 19970 -734
rect 20526 -734 20542 -717
rect 20972 -717 21560 -701
rect 20972 -734 20988 -717
rect 20526 -751 20728 -734
rect 19768 -798 20728 -751
rect 20786 -751 20988 -734
rect 21544 -734 21560 -717
rect 21990 -717 22578 -701
rect 21990 -734 22006 -717
rect 21544 -751 21746 -734
rect 20786 -798 21746 -751
rect 21804 -751 22006 -734
rect 22562 -734 22578 -717
rect 22562 -751 22764 -734
rect 21804 -798 22764 -751
rect 6534 -1445 7494 -1398
rect 6534 -1462 6736 -1445
rect 6720 -1479 6736 -1462
rect 7292 -1462 7494 -1445
rect 7552 -1445 8512 -1398
rect 7552 -1462 7754 -1445
rect 7292 -1479 7308 -1462
rect 6720 -1495 7308 -1479
rect 7738 -1479 7754 -1462
rect 8310 -1462 8512 -1445
rect 8570 -1445 9530 -1398
rect 8570 -1462 8772 -1445
rect 8310 -1479 8326 -1462
rect 7738 -1495 8326 -1479
rect 8756 -1479 8772 -1462
rect 9328 -1462 9530 -1445
rect 9588 -1445 10548 -1398
rect 9588 -1462 9790 -1445
rect 9328 -1479 9344 -1462
rect 8756 -1495 9344 -1479
rect 9774 -1479 9790 -1462
rect 10346 -1462 10548 -1445
rect 10606 -1445 11566 -1398
rect 10606 -1462 10808 -1445
rect 10346 -1479 10362 -1462
rect 9774 -1495 10362 -1479
rect 10792 -1479 10808 -1462
rect 11364 -1462 11566 -1445
rect 11624 -1445 12584 -1398
rect 11624 -1462 11826 -1445
rect 11364 -1479 11380 -1462
rect 10792 -1495 11380 -1479
rect 11810 -1479 11826 -1462
rect 12382 -1462 12584 -1445
rect 12642 -1445 13602 -1398
rect 12642 -1462 12844 -1445
rect 12382 -1479 12398 -1462
rect 11810 -1495 12398 -1479
rect 12828 -1479 12844 -1462
rect 13400 -1462 13602 -1445
rect 13660 -1445 14620 -1398
rect 13660 -1462 13862 -1445
rect 13400 -1479 13416 -1462
rect 12828 -1495 13416 -1479
rect 13846 -1479 13862 -1462
rect 14418 -1462 14620 -1445
rect 14678 -1445 15638 -1398
rect 14678 -1462 14880 -1445
rect 14418 -1479 14434 -1462
rect 13846 -1495 14434 -1479
rect 14864 -1479 14880 -1462
rect 15436 -1462 15638 -1445
rect 15696 -1445 16656 -1398
rect 15696 -1462 15898 -1445
rect 15436 -1479 15452 -1462
rect 14864 -1495 15452 -1479
rect 15882 -1479 15898 -1462
rect 16454 -1462 16656 -1445
rect 16714 -1445 17674 -1398
rect 16714 -1462 16916 -1445
rect 16454 -1479 16470 -1462
rect 15882 -1495 16470 -1479
rect 16900 -1479 16916 -1462
rect 17472 -1462 17674 -1445
rect 17732 -1445 18692 -1398
rect 17732 -1462 17934 -1445
rect 17472 -1479 17488 -1462
rect 16900 -1495 17488 -1479
rect 17918 -1479 17934 -1462
rect 18490 -1462 18692 -1445
rect 18750 -1445 19710 -1398
rect 18750 -1462 18952 -1445
rect 18490 -1479 18506 -1462
rect 17918 -1495 18506 -1479
rect 18936 -1479 18952 -1462
rect 19508 -1462 19710 -1445
rect 19768 -1445 20728 -1398
rect 19768 -1462 19970 -1445
rect 19508 -1479 19524 -1462
rect 18936 -1495 19524 -1479
rect 19954 -1479 19970 -1462
rect 20526 -1462 20728 -1445
rect 20786 -1445 21746 -1398
rect 20786 -1462 20988 -1445
rect 20526 -1479 20542 -1462
rect 19954 -1495 20542 -1479
rect 20972 -1479 20988 -1462
rect 21544 -1462 21746 -1445
rect 21804 -1445 22764 -1398
rect 21804 -1462 22006 -1445
rect 21544 -1479 21560 -1462
rect 20972 -1495 21560 -1479
rect 21990 -1479 22006 -1462
rect 22562 -1462 22764 -1445
rect 22562 -1479 22578 -1462
rect 21990 -1495 22578 -1479
rect 7914 -2355 8502 -2339
rect 7914 -2372 7930 -2355
rect 7728 -2389 7930 -2372
rect 8486 -2372 8502 -2355
rect 8932 -2355 9520 -2339
rect 8932 -2372 8948 -2355
rect 8486 -2389 8688 -2372
rect 7728 -2436 8688 -2389
rect 8746 -2389 8948 -2372
rect 9504 -2372 9520 -2355
rect 9950 -2355 10538 -2339
rect 9950 -2372 9966 -2355
rect 9504 -2389 9706 -2372
rect 8746 -2436 9706 -2389
rect 9764 -2389 9966 -2372
rect 10522 -2372 10538 -2355
rect 10968 -2355 11556 -2339
rect 10968 -2372 10984 -2355
rect 10522 -2389 10724 -2372
rect 9764 -2436 10724 -2389
rect 10782 -2389 10984 -2372
rect 11540 -2372 11556 -2355
rect 11986 -2355 12574 -2339
rect 11986 -2372 12002 -2355
rect 11540 -2389 11742 -2372
rect 10782 -2436 11742 -2389
rect 11800 -2389 12002 -2372
rect 12558 -2372 12574 -2355
rect 13004 -2355 13592 -2339
rect 13004 -2372 13020 -2355
rect 12558 -2389 12760 -2372
rect 11800 -2436 12760 -2389
rect 12818 -2389 13020 -2372
rect 13576 -2372 13592 -2355
rect 14022 -2355 14610 -2339
rect 14022 -2372 14038 -2355
rect 13576 -2389 13778 -2372
rect 12818 -2436 13778 -2389
rect 13836 -2389 14038 -2372
rect 14594 -2372 14610 -2355
rect 15040 -2355 15628 -2339
rect 15040 -2372 15056 -2355
rect 14594 -2389 14796 -2372
rect 13836 -2436 14796 -2389
rect 14854 -2389 15056 -2372
rect 15612 -2372 15628 -2355
rect 16058 -2355 16646 -2339
rect 16058 -2372 16074 -2355
rect 15612 -2389 15814 -2372
rect 14854 -2436 15814 -2389
rect 15872 -2389 16074 -2372
rect 16630 -2372 16646 -2355
rect 17076 -2355 17664 -2339
rect 17076 -2372 17092 -2355
rect 16630 -2389 16832 -2372
rect 15872 -2436 16832 -2389
rect 16890 -2389 17092 -2372
rect 17648 -2372 17664 -2355
rect 18094 -2355 18682 -2339
rect 18094 -2372 18110 -2355
rect 17648 -2389 17850 -2372
rect 16890 -2436 17850 -2389
rect 17908 -2389 18110 -2372
rect 18666 -2372 18682 -2355
rect 19112 -2355 19700 -2339
rect 19112 -2372 19128 -2355
rect 18666 -2389 18868 -2372
rect 17908 -2436 18868 -2389
rect 18926 -2389 19128 -2372
rect 19684 -2372 19700 -2355
rect 20130 -2355 20718 -2339
rect 20130 -2372 20146 -2355
rect 19684 -2389 19886 -2372
rect 18926 -2436 19886 -2389
rect 19944 -2389 20146 -2372
rect 20702 -2372 20718 -2355
rect 21148 -2355 21736 -2339
rect 21148 -2372 21164 -2355
rect 20702 -2389 20904 -2372
rect 19944 -2436 20904 -2389
rect 20962 -2389 21164 -2372
rect 21720 -2372 21736 -2355
rect 21720 -2389 21922 -2372
rect 20962 -2436 21922 -2389
rect 7728 -3083 8688 -3036
rect 7728 -3100 7930 -3083
rect 7914 -3117 7930 -3100
rect 8486 -3100 8688 -3083
rect 8746 -3083 9706 -3036
rect 8746 -3100 8948 -3083
rect 8486 -3117 8502 -3100
rect 7914 -3133 8502 -3117
rect 8932 -3117 8948 -3100
rect 9504 -3100 9706 -3083
rect 9764 -3083 10724 -3036
rect 9764 -3100 9966 -3083
rect 9504 -3117 9520 -3100
rect 8932 -3133 9520 -3117
rect 9950 -3117 9966 -3100
rect 10522 -3100 10724 -3083
rect 10782 -3083 11742 -3036
rect 10782 -3100 10984 -3083
rect 10522 -3117 10538 -3100
rect 9950 -3133 10538 -3117
rect 10968 -3117 10984 -3100
rect 11540 -3100 11742 -3083
rect 11800 -3083 12760 -3036
rect 11800 -3100 12002 -3083
rect 11540 -3117 11556 -3100
rect 10968 -3133 11556 -3117
rect 11986 -3117 12002 -3100
rect 12558 -3100 12760 -3083
rect 12818 -3083 13778 -3036
rect 12818 -3100 13020 -3083
rect 12558 -3117 12574 -3100
rect 11986 -3133 12574 -3117
rect 13004 -3117 13020 -3100
rect 13576 -3100 13778 -3083
rect 13836 -3083 14796 -3036
rect 13836 -3100 14038 -3083
rect 13576 -3117 13592 -3100
rect 13004 -3133 13592 -3117
rect 14022 -3117 14038 -3100
rect 14594 -3100 14796 -3083
rect 14854 -3083 15814 -3036
rect 14854 -3100 15056 -3083
rect 14594 -3117 14610 -3100
rect 14022 -3133 14610 -3117
rect 15040 -3117 15056 -3100
rect 15612 -3100 15814 -3083
rect 15872 -3083 16832 -3036
rect 15872 -3100 16074 -3083
rect 15612 -3117 15628 -3100
rect 15040 -3133 15628 -3117
rect 16058 -3117 16074 -3100
rect 16630 -3100 16832 -3083
rect 16890 -3083 17850 -3036
rect 16890 -3100 17092 -3083
rect 16630 -3117 16646 -3100
rect 16058 -3133 16646 -3117
rect 17076 -3117 17092 -3100
rect 17648 -3100 17850 -3083
rect 17908 -3083 18868 -3036
rect 17908 -3100 18110 -3083
rect 17648 -3117 17664 -3100
rect 17076 -3133 17664 -3117
rect 18094 -3117 18110 -3100
rect 18666 -3100 18868 -3083
rect 18926 -3083 19886 -3036
rect 18926 -3100 19128 -3083
rect 18666 -3117 18682 -3100
rect 18094 -3133 18682 -3117
rect 19112 -3117 19128 -3100
rect 19684 -3100 19886 -3083
rect 19944 -3083 20904 -3036
rect 19944 -3100 20146 -3083
rect 19684 -3117 19700 -3100
rect 19112 -3133 19700 -3117
rect 20130 -3117 20146 -3100
rect 20702 -3100 20904 -3083
rect 20962 -3083 21922 -3036
rect 20962 -3100 21164 -3083
rect 20702 -3117 20718 -3100
rect 20130 -3133 20718 -3117
rect 21148 -3117 21164 -3100
rect 21720 -3100 21922 -3083
rect 21720 -3117 21736 -3100
rect 21148 -3133 21736 -3117
rect 7914 -3387 8502 -3371
rect 7914 -3404 7930 -3387
rect 7728 -3421 7930 -3404
rect 8486 -3404 8502 -3387
rect 8932 -3387 9520 -3371
rect 8932 -3404 8948 -3387
rect 8486 -3421 8688 -3404
rect 7728 -3468 8688 -3421
rect 8746 -3421 8948 -3404
rect 9504 -3404 9520 -3387
rect 9950 -3387 10538 -3371
rect 9950 -3404 9966 -3387
rect 9504 -3421 9706 -3404
rect 8746 -3468 9706 -3421
rect 9764 -3421 9966 -3404
rect 10522 -3404 10538 -3387
rect 10968 -3387 11556 -3371
rect 10968 -3404 10984 -3387
rect 10522 -3421 10724 -3404
rect 9764 -3468 10724 -3421
rect 10782 -3421 10984 -3404
rect 11540 -3404 11556 -3387
rect 11986 -3387 12574 -3371
rect 11986 -3404 12002 -3387
rect 11540 -3421 11742 -3404
rect 10782 -3468 11742 -3421
rect 11800 -3421 12002 -3404
rect 12558 -3404 12574 -3387
rect 13004 -3387 13592 -3371
rect 13004 -3404 13020 -3387
rect 12558 -3421 12760 -3404
rect 11800 -3468 12760 -3421
rect 12818 -3421 13020 -3404
rect 13576 -3404 13592 -3387
rect 14022 -3387 14610 -3371
rect 14022 -3404 14038 -3387
rect 13576 -3421 13778 -3404
rect 12818 -3468 13778 -3421
rect 13836 -3421 14038 -3404
rect 14594 -3404 14610 -3387
rect 15040 -3387 15628 -3371
rect 15040 -3404 15056 -3387
rect 14594 -3421 14796 -3404
rect 13836 -3468 14796 -3421
rect 14854 -3421 15056 -3404
rect 15612 -3404 15628 -3387
rect 16058 -3387 16646 -3371
rect 16058 -3404 16074 -3387
rect 15612 -3421 15814 -3404
rect 14854 -3468 15814 -3421
rect 15872 -3421 16074 -3404
rect 16630 -3404 16646 -3387
rect 17076 -3387 17664 -3371
rect 17076 -3404 17092 -3387
rect 16630 -3421 16832 -3404
rect 15872 -3468 16832 -3421
rect 16890 -3421 17092 -3404
rect 17648 -3404 17664 -3387
rect 18094 -3387 18682 -3371
rect 18094 -3404 18110 -3387
rect 17648 -3421 17850 -3404
rect 16890 -3468 17850 -3421
rect 17908 -3421 18110 -3404
rect 18666 -3404 18682 -3387
rect 19112 -3387 19700 -3371
rect 19112 -3404 19128 -3387
rect 18666 -3421 18868 -3404
rect 17908 -3468 18868 -3421
rect 18926 -3421 19128 -3404
rect 19684 -3404 19700 -3387
rect 20130 -3387 20718 -3371
rect 20130 -3404 20146 -3387
rect 19684 -3421 19886 -3404
rect 18926 -3468 19886 -3421
rect 19944 -3421 20146 -3404
rect 20702 -3404 20718 -3387
rect 21148 -3387 21736 -3371
rect 21148 -3404 21164 -3387
rect 20702 -3421 20904 -3404
rect 19944 -3468 20904 -3421
rect 20962 -3421 21164 -3404
rect 21720 -3404 21736 -3387
rect 21720 -3421 21922 -3404
rect 20962 -3468 21922 -3421
rect 7728 -4115 8688 -4068
rect 7728 -4132 7930 -4115
rect 7914 -4149 7930 -4132
rect 8486 -4132 8688 -4115
rect 8746 -4115 9706 -4068
rect 8746 -4132 8948 -4115
rect 8486 -4149 8502 -4132
rect 7914 -4165 8502 -4149
rect 8932 -4149 8948 -4132
rect 9504 -4132 9706 -4115
rect 9764 -4115 10724 -4068
rect 9764 -4132 9966 -4115
rect 9504 -4149 9520 -4132
rect 8932 -4165 9520 -4149
rect 9950 -4149 9966 -4132
rect 10522 -4132 10724 -4115
rect 10782 -4115 11742 -4068
rect 10782 -4132 10984 -4115
rect 10522 -4149 10538 -4132
rect 9950 -4165 10538 -4149
rect 10968 -4149 10984 -4132
rect 11540 -4132 11742 -4115
rect 11800 -4115 12760 -4068
rect 11800 -4132 12002 -4115
rect 11540 -4149 11556 -4132
rect 10968 -4165 11556 -4149
rect 11986 -4149 12002 -4132
rect 12558 -4132 12760 -4115
rect 12818 -4115 13778 -4068
rect 12818 -4132 13020 -4115
rect 12558 -4149 12574 -4132
rect 11986 -4165 12574 -4149
rect 13004 -4149 13020 -4132
rect 13576 -4132 13778 -4115
rect 13836 -4115 14796 -4068
rect 13836 -4132 14038 -4115
rect 13576 -4149 13592 -4132
rect 13004 -4165 13592 -4149
rect 14022 -4149 14038 -4132
rect 14594 -4132 14796 -4115
rect 14854 -4115 15814 -4068
rect 14854 -4132 15056 -4115
rect 14594 -4149 14610 -4132
rect 14022 -4165 14610 -4149
rect 15040 -4149 15056 -4132
rect 15612 -4132 15814 -4115
rect 15872 -4115 16832 -4068
rect 15872 -4132 16074 -4115
rect 15612 -4149 15628 -4132
rect 15040 -4165 15628 -4149
rect 16058 -4149 16074 -4132
rect 16630 -4132 16832 -4115
rect 16890 -4115 17850 -4068
rect 16890 -4132 17092 -4115
rect 16630 -4149 16646 -4132
rect 16058 -4165 16646 -4149
rect 17076 -4149 17092 -4132
rect 17648 -4132 17850 -4115
rect 17908 -4115 18868 -4068
rect 17908 -4132 18110 -4115
rect 17648 -4149 17664 -4132
rect 17076 -4165 17664 -4149
rect 18094 -4149 18110 -4132
rect 18666 -4132 18868 -4115
rect 18926 -4115 19886 -4068
rect 18926 -4132 19128 -4115
rect 18666 -4149 18682 -4132
rect 18094 -4165 18682 -4149
rect 19112 -4149 19128 -4132
rect 19684 -4132 19886 -4115
rect 19944 -4115 20904 -4068
rect 19944 -4132 20146 -4115
rect 19684 -4149 19700 -4132
rect 19112 -4165 19700 -4149
rect 20130 -4149 20146 -4132
rect 20702 -4132 20904 -4115
rect 20962 -4115 21922 -4068
rect 20962 -4132 21164 -4115
rect 20702 -4149 20718 -4132
rect 20130 -4165 20718 -4149
rect 21148 -4149 21164 -4132
rect 21720 -4132 21922 -4115
rect 21720 -4149 21736 -4132
rect 21148 -4165 21736 -4149
rect 7706 -4991 8294 -4975
rect 7706 -5008 7722 -4991
rect 7520 -5025 7722 -5008
rect 8278 -5008 8294 -4991
rect 8724 -4991 9312 -4975
rect 8724 -5008 8740 -4991
rect 8278 -5025 8480 -5008
rect 7520 -5072 8480 -5025
rect 8538 -5025 8740 -5008
rect 9296 -5008 9312 -4991
rect 9742 -4991 10330 -4975
rect 9742 -5008 9758 -4991
rect 9296 -5025 9498 -5008
rect 8538 -5072 9498 -5025
rect 9556 -5025 9758 -5008
rect 10314 -5008 10330 -4991
rect 10760 -4991 11348 -4975
rect 10760 -5008 10776 -4991
rect 10314 -5025 10516 -5008
rect 9556 -5072 10516 -5025
rect 10574 -5025 10776 -5008
rect 11332 -5008 11348 -4991
rect 11778 -4991 12366 -4975
rect 11778 -5008 11794 -4991
rect 11332 -5025 11534 -5008
rect 10574 -5072 11534 -5025
rect 11592 -5025 11794 -5008
rect 12350 -5008 12366 -4991
rect 12796 -4991 13384 -4975
rect 12796 -5008 12812 -4991
rect 12350 -5025 12552 -5008
rect 11592 -5072 12552 -5025
rect 12610 -5025 12812 -5008
rect 13368 -5008 13384 -4991
rect 13814 -4991 14402 -4975
rect 13814 -5008 13830 -4991
rect 13368 -5025 13570 -5008
rect 12610 -5072 13570 -5025
rect 13628 -5025 13830 -5008
rect 14386 -5008 14402 -4991
rect 14832 -4991 15420 -4975
rect 14832 -5008 14848 -4991
rect 14386 -5025 14588 -5008
rect 13628 -5072 14588 -5025
rect 14646 -5025 14848 -5008
rect 15404 -5008 15420 -4991
rect 15850 -4991 16438 -4975
rect 15850 -5008 15866 -4991
rect 15404 -5025 15606 -5008
rect 14646 -5072 15606 -5025
rect 15664 -5025 15866 -5008
rect 16422 -5008 16438 -4991
rect 16868 -4991 17456 -4975
rect 16868 -5008 16884 -4991
rect 16422 -5025 16624 -5008
rect 15664 -5072 16624 -5025
rect 16682 -5025 16884 -5008
rect 17440 -5008 17456 -4991
rect 17886 -4991 18474 -4975
rect 17886 -5008 17902 -4991
rect 17440 -5025 17642 -5008
rect 16682 -5072 17642 -5025
rect 17700 -5025 17902 -5008
rect 18458 -5008 18474 -4991
rect 18904 -4991 19492 -4975
rect 18904 -5008 18920 -4991
rect 18458 -5025 18660 -5008
rect 17700 -5072 18660 -5025
rect 18718 -5025 18920 -5008
rect 19476 -5008 19492 -4991
rect 19922 -4991 20510 -4975
rect 19922 -5008 19938 -4991
rect 19476 -5025 19678 -5008
rect 18718 -5072 19678 -5025
rect 19736 -5025 19938 -5008
rect 20494 -5008 20510 -4991
rect 20940 -4991 21528 -4975
rect 20940 -5008 20956 -4991
rect 20494 -5025 20696 -5008
rect 19736 -5072 20696 -5025
rect 20754 -5025 20956 -5008
rect 21512 -5008 21528 -4991
rect 21958 -4991 22546 -4975
rect 21958 -5008 21974 -4991
rect 21512 -5025 21714 -5008
rect 20754 -5072 21714 -5025
rect 21772 -5025 21974 -5008
rect 22530 -5008 22546 -4991
rect 22530 -5025 22732 -5008
rect 21772 -5072 22732 -5025
rect 2402 -5095 2990 -5079
rect 2402 -5112 2418 -5095
rect 2216 -5129 2418 -5112
rect 2974 -5112 2990 -5095
rect 3420 -5095 4008 -5079
rect 3420 -5112 3436 -5095
rect 2974 -5129 3176 -5112
rect 2216 -5176 3176 -5129
rect 3234 -5129 3436 -5112
rect 3992 -5112 4008 -5095
rect 4438 -5095 5026 -5079
rect 4438 -5112 4454 -5095
rect 3992 -5129 4194 -5112
rect 3234 -5176 4194 -5129
rect 4252 -5129 4454 -5112
rect 5010 -5112 5026 -5095
rect 5456 -5095 6044 -5079
rect 5456 -5112 5472 -5095
rect 5010 -5129 5212 -5112
rect 4252 -5176 5212 -5129
rect 5270 -5129 5472 -5112
rect 6028 -5112 6044 -5095
rect 6028 -5129 6230 -5112
rect 5270 -5176 6230 -5129
rect 7520 -5719 8480 -5672
rect 7520 -5736 7722 -5719
rect 7706 -5753 7722 -5736
rect 8278 -5736 8480 -5719
rect 8538 -5719 9498 -5672
rect 8538 -5736 8740 -5719
rect 8278 -5753 8294 -5736
rect 7706 -5769 8294 -5753
rect 8724 -5753 8740 -5736
rect 9296 -5736 9498 -5719
rect 9556 -5719 10516 -5672
rect 9556 -5736 9758 -5719
rect 9296 -5753 9312 -5736
rect 8724 -5769 9312 -5753
rect 9742 -5753 9758 -5736
rect 10314 -5736 10516 -5719
rect 10574 -5719 11534 -5672
rect 10574 -5736 10776 -5719
rect 10314 -5753 10330 -5736
rect 9742 -5769 10330 -5753
rect 10760 -5753 10776 -5736
rect 11332 -5736 11534 -5719
rect 11592 -5719 12552 -5672
rect 11592 -5736 11794 -5719
rect 11332 -5753 11348 -5736
rect 10760 -5769 11348 -5753
rect 11778 -5753 11794 -5736
rect 12350 -5736 12552 -5719
rect 12610 -5719 13570 -5672
rect 12610 -5736 12812 -5719
rect 12350 -5753 12366 -5736
rect 11778 -5769 12366 -5753
rect 12796 -5753 12812 -5736
rect 13368 -5736 13570 -5719
rect 13628 -5719 14588 -5672
rect 13628 -5736 13830 -5719
rect 13368 -5753 13384 -5736
rect 12796 -5769 13384 -5753
rect 13814 -5753 13830 -5736
rect 14386 -5736 14588 -5719
rect 14646 -5719 15606 -5672
rect 14646 -5736 14848 -5719
rect 14386 -5753 14402 -5736
rect 13814 -5769 14402 -5753
rect 14832 -5753 14848 -5736
rect 15404 -5736 15606 -5719
rect 15664 -5719 16624 -5672
rect 15664 -5736 15866 -5719
rect 15404 -5753 15420 -5736
rect 14832 -5769 15420 -5753
rect 15850 -5753 15866 -5736
rect 16422 -5736 16624 -5719
rect 16682 -5719 17642 -5672
rect 16682 -5736 16884 -5719
rect 16422 -5753 16438 -5736
rect 15850 -5769 16438 -5753
rect 16868 -5753 16884 -5736
rect 17440 -5736 17642 -5719
rect 17700 -5719 18660 -5672
rect 17700 -5736 17902 -5719
rect 17440 -5753 17456 -5736
rect 16868 -5769 17456 -5753
rect 17886 -5753 17902 -5736
rect 18458 -5736 18660 -5719
rect 18718 -5719 19678 -5672
rect 18718 -5736 18920 -5719
rect 18458 -5753 18474 -5736
rect 17886 -5769 18474 -5753
rect 18904 -5753 18920 -5736
rect 19476 -5736 19678 -5719
rect 19736 -5719 20696 -5672
rect 19736 -5736 19938 -5719
rect 19476 -5753 19492 -5736
rect 18904 -5769 19492 -5753
rect 19922 -5753 19938 -5736
rect 20494 -5736 20696 -5719
rect 20754 -5719 21714 -5672
rect 20754 -5736 20956 -5719
rect 20494 -5753 20510 -5736
rect 19922 -5769 20510 -5753
rect 20940 -5753 20956 -5736
rect 21512 -5736 21714 -5719
rect 21772 -5719 22732 -5672
rect 21772 -5736 21974 -5719
rect 21512 -5753 21528 -5736
rect 20940 -5769 21528 -5753
rect 21958 -5753 21974 -5736
rect 22530 -5736 22732 -5719
rect 22530 -5753 22546 -5736
rect 21958 -5769 22546 -5753
rect 2216 -5823 3176 -5776
rect 2216 -5840 2418 -5823
rect 2402 -5857 2418 -5840
rect 2974 -5840 3176 -5823
rect 3234 -5823 4194 -5776
rect 3234 -5840 3436 -5823
rect 2974 -5857 2990 -5840
rect 2402 -5873 2990 -5857
rect 3420 -5857 3436 -5840
rect 3992 -5840 4194 -5823
rect 4252 -5823 5212 -5776
rect 4252 -5840 4454 -5823
rect 3992 -5857 4008 -5840
rect 3420 -5873 4008 -5857
rect 4438 -5857 4454 -5840
rect 5010 -5840 5212 -5823
rect 5270 -5823 6230 -5776
rect 5270 -5840 5472 -5823
rect 5010 -5857 5026 -5840
rect 4438 -5873 5026 -5857
rect 5456 -5857 5472 -5840
rect 6028 -5840 6230 -5823
rect 6028 -5857 6044 -5840
rect 5456 -5873 6044 -5857
rect 2402 -6127 2990 -6111
rect 2402 -6144 2418 -6127
rect 2216 -6161 2418 -6144
rect 2974 -6144 2990 -6127
rect 3420 -6127 4008 -6111
rect 3420 -6144 3436 -6127
rect 2974 -6161 3176 -6144
rect 2216 -6208 3176 -6161
rect 3234 -6161 3436 -6144
rect 3992 -6144 4008 -6127
rect 4438 -6127 5026 -6111
rect 4438 -6144 4454 -6127
rect 3992 -6161 4194 -6144
rect 3234 -6208 4194 -6161
rect 4252 -6161 4454 -6144
rect 5010 -6144 5026 -6127
rect 5456 -6127 6044 -6111
rect 5456 -6144 5472 -6127
rect 5010 -6161 5212 -6144
rect 4252 -6208 5212 -6161
rect 5270 -6161 5472 -6144
rect 6028 -6144 6044 -6127
rect 6028 -6161 6230 -6144
rect 5270 -6208 6230 -6161
rect 7706 -6247 8294 -6231
rect 7706 -6264 7722 -6247
rect 7520 -6281 7722 -6264
rect 8278 -6264 8294 -6247
rect 8724 -6247 9312 -6231
rect 8724 -6264 8740 -6247
rect 8278 -6281 8480 -6264
rect 7520 -6328 8480 -6281
rect 8538 -6281 8740 -6264
rect 9296 -6264 9312 -6247
rect 9742 -6247 10330 -6231
rect 9742 -6264 9758 -6247
rect 9296 -6281 9498 -6264
rect 8538 -6328 9498 -6281
rect 9556 -6281 9758 -6264
rect 10314 -6264 10330 -6247
rect 10760 -6247 11348 -6231
rect 10760 -6264 10776 -6247
rect 10314 -6281 10516 -6264
rect 9556 -6328 10516 -6281
rect 10574 -6281 10776 -6264
rect 11332 -6264 11348 -6247
rect 11778 -6247 12366 -6231
rect 11778 -6264 11794 -6247
rect 11332 -6281 11534 -6264
rect 10574 -6328 11534 -6281
rect 11592 -6281 11794 -6264
rect 12350 -6264 12366 -6247
rect 12796 -6247 13384 -6231
rect 12796 -6264 12812 -6247
rect 12350 -6281 12552 -6264
rect 11592 -6328 12552 -6281
rect 12610 -6281 12812 -6264
rect 13368 -6264 13384 -6247
rect 13814 -6247 14402 -6231
rect 13814 -6264 13830 -6247
rect 13368 -6281 13570 -6264
rect 12610 -6328 13570 -6281
rect 13628 -6281 13830 -6264
rect 14386 -6264 14402 -6247
rect 14832 -6247 15420 -6231
rect 14832 -6264 14848 -6247
rect 14386 -6281 14588 -6264
rect 13628 -6328 14588 -6281
rect 14646 -6281 14848 -6264
rect 15404 -6264 15420 -6247
rect 15850 -6247 16438 -6231
rect 15850 -6264 15866 -6247
rect 15404 -6281 15606 -6264
rect 14646 -6328 15606 -6281
rect 15664 -6281 15866 -6264
rect 16422 -6264 16438 -6247
rect 16868 -6247 17456 -6231
rect 16868 -6264 16884 -6247
rect 16422 -6281 16624 -6264
rect 15664 -6328 16624 -6281
rect 16682 -6281 16884 -6264
rect 17440 -6264 17456 -6247
rect 17886 -6247 18474 -6231
rect 17886 -6264 17902 -6247
rect 17440 -6281 17642 -6264
rect 16682 -6328 17642 -6281
rect 17700 -6281 17902 -6264
rect 18458 -6264 18474 -6247
rect 18904 -6247 19492 -6231
rect 18904 -6264 18920 -6247
rect 18458 -6281 18660 -6264
rect 17700 -6328 18660 -6281
rect 18718 -6281 18920 -6264
rect 19476 -6264 19492 -6247
rect 19922 -6247 20510 -6231
rect 19922 -6264 19938 -6247
rect 19476 -6281 19678 -6264
rect 18718 -6328 19678 -6281
rect 19736 -6281 19938 -6264
rect 20494 -6264 20510 -6247
rect 20940 -6247 21528 -6231
rect 20940 -6264 20956 -6247
rect 20494 -6281 20696 -6264
rect 19736 -6328 20696 -6281
rect 20754 -6281 20956 -6264
rect 21512 -6264 21528 -6247
rect 21958 -6247 22546 -6231
rect 21958 -6264 21974 -6247
rect 21512 -6281 21714 -6264
rect 20754 -6328 21714 -6281
rect 21772 -6281 21974 -6264
rect 22530 -6264 22546 -6247
rect 22530 -6281 22732 -6264
rect 21772 -6328 22732 -6281
rect 2216 -6855 3176 -6808
rect 2216 -6872 2418 -6855
rect 2402 -6889 2418 -6872
rect 2974 -6872 3176 -6855
rect 3234 -6855 4194 -6808
rect 3234 -6872 3436 -6855
rect 2974 -6889 2990 -6872
rect 2402 -6905 2990 -6889
rect 3420 -6889 3436 -6872
rect 3992 -6872 4194 -6855
rect 4252 -6855 5212 -6808
rect 4252 -6872 4454 -6855
rect 3992 -6889 4008 -6872
rect 3420 -6905 4008 -6889
rect 4438 -6889 4454 -6872
rect 5010 -6872 5212 -6855
rect 5270 -6855 6230 -6808
rect 5270 -6872 5472 -6855
rect 5010 -6889 5026 -6872
rect 4438 -6905 5026 -6889
rect 5456 -6889 5472 -6872
rect 6028 -6872 6230 -6855
rect 6028 -6889 6044 -6872
rect 5456 -6905 6044 -6889
rect 7520 -6975 8480 -6928
rect 7520 -6992 7722 -6975
rect 7706 -7009 7722 -6992
rect 8278 -6992 8480 -6975
rect 8538 -6975 9498 -6928
rect 8538 -6992 8740 -6975
rect 8278 -7009 8294 -6992
rect 7706 -7025 8294 -7009
rect 8724 -7009 8740 -6992
rect 9296 -6992 9498 -6975
rect 9556 -6975 10516 -6928
rect 9556 -6992 9758 -6975
rect 9296 -7009 9312 -6992
rect 8724 -7025 9312 -7009
rect 9742 -7009 9758 -6992
rect 10314 -6992 10516 -6975
rect 10574 -6975 11534 -6928
rect 10574 -6992 10776 -6975
rect 10314 -7009 10330 -6992
rect 9742 -7025 10330 -7009
rect 10760 -7009 10776 -6992
rect 11332 -6992 11534 -6975
rect 11592 -6975 12552 -6928
rect 11592 -6992 11794 -6975
rect 11332 -7009 11348 -6992
rect 10760 -7025 11348 -7009
rect 11778 -7009 11794 -6992
rect 12350 -6992 12552 -6975
rect 12610 -6975 13570 -6928
rect 12610 -6992 12812 -6975
rect 12350 -7009 12366 -6992
rect 11778 -7025 12366 -7009
rect 12796 -7009 12812 -6992
rect 13368 -6992 13570 -6975
rect 13628 -6975 14588 -6928
rect 13628 -6992 13830 -6975
rect 13368 -7009 13384 -6992
rect 12796 -7025 13384 -7009
rect 13814 -7009 13830 -6992
rect 14386 -6992 14588 -6975
rect 14646 -6975 15606 -6928
rect 14646 -6992 14848 -6975
rect 14386 -7009 14402 -6992
rect 13814 -7025 14402 -7009
rect 14832 -7009 14848 -6992
rect 15404 -6992 15606 -6975
rect 15664 -6975 16624 -6928
rect 15664 -6992 15866 -6975
rect 15404 -7009 15420 -6992
rect 14832 -7025 15420 -7009
rect 15850 -7009 15866 -6992
rect 16422 -6992 16624 -6975
rect 16682 -6975 17642 -6928
rect 16682 -6992 16884 -6975
rect 16422 -7009 16438 -6992
rect 15850 -7025 16438 -7009
rect 16868 -7009 16884 -6992
rect 17440 -6992 17642 -6975
rect 17700 -6975 18660 -6928
rect 17700 -6992 17902 -6975
rect 17440 -7009 17456 -6992
rect 16868 -7025 17456 -7009
rect 17886 -7009 17902 -6992
rect 18458 -6992 18660 -6975
rect 18718 -6975 19678 -6928
rect 18718 -6992 18920 -6975
rect 18458 -7009 18474 -6992
rect 17886 -7025 18474 -7009
rect 18904 -7009 18920 -6992
rect 19476 -6992 19678 -6975
rect 19736 -6975 20696 -6928
rect 19736 -6992 19938 -6975
rect 19476 -7009 19492 -6992
rect 18904 -7025 19492 -7009
rect 19922 -7009 19938 -6992
rect 20494 -6992 20696 -6975
rect 20754 -6975 21714 -6928
rect 20754 -6992 20956 -6975
rect 20494 -7009 20510 -6992
rect 19922 -7025 20510 -7009
rect 20940 -7009 20956 -6992
rect 21512 -6992 21714 -6975
rect 21772 -6975 22732 -6928
rect 21772 -6992 21974 -6975
rect 21512 -7009 21528 -6992
rect 20940 -7025 21528 -7009
rect 21958 -7009 21974 -6992
rect 22530 -6992 22732 -6975
rect 22530 -7009 22546 -6992
rect 21958 -7025 22546 -7009
rect 2402 -7159 2990 -7143
rect 2402 -7176 2418 -7159
rect 2216 -7193 2418 -7176
rect 2974 -7176 2990 -7159
rect 3420 -7159 4008 -7143
rect 3420 -7176 3436 -7159
rect 2974 -7193 3176 -7176
rect 2216 -7240 3176 -7193
rect 3234 -7193 3436 -7176
rect 3992 -7176 4008 -7159
rect 4438 -7159 5026 -7143
rect 4438 -7176 4454 -7159
rect 3992 -7193 4194 -7176
rect 3234 -7240 4194 -7193
rect 4252 -7193 4454 -7176
rect 5010 -7176 5026 -7159
rect 5456 -7159 6044 -7143
rect 5456 -7176 5472 -7159
rect 5010 -7193 5212 -7176
rect 4252 -7240 5212 -7193
rect 5270 -7193 5472 -7176
rect 6028 -7176 6044 -7159
rect 6028 -7193 6230 -7176
rect 5270 -7240 6230 -7193
rect 7706 -7503 8294 -7487
rect 7706 -7520 7722 -7503
rect 7520 -7537 7722 -7520
rect 8278 -7520 8294 -7503
rect 8724 -7503 9312 -7487
rect 8724 -7520 8740 -7503
rect 8278 -7537 8480 -7520
rect 7520 -7584 8480 -7537
rect 8538 -7537 8740 -7520
rect 9296 -7520 9312 -7503
rect 9742 -7503 10330 -7487
rect 9742 -7520 9758 -7503
rect 9296 -7537 9498 -7520
rect 8538 -7584 9498 -7537
rect 9556 -7537 9758 -7520
rect 10314 -7520 10330 -7503
rect 10760 -7503 11348 -7487
rect 10760 -7520 10776 -7503
rect 10314 -7537 10516 -7520
rect 9556 -7584 10516 -7537
rect 10574 -7537 10776 -7520
rect 11332 -7520 11348 -7503
rect 11778 -7503 12366 -7487
rect 11778 -7520 11794 -7503
rect 11332 -7537 11534 -7520
rect 10574 -7584 11534 -7537
rect 11592 -7537 11794 -7520
rect 12350 -7520 12366 -7503
rect 12796 -7503 13384 -7487
rect 12796 -7520 12812 -7503
rect 12350 -7537 12552 -7520
rect 11592 -7584 12552 -7537
rect 12610 -7537 12812 -7520
rect 13368 -7520 13384 -7503
rect 13814 -7503 14402 -7487
rect 13814 -7520 13830 -7503
rect 13368 -7537 13570 -7520
rect 12610 -7584 13570 -7537
rect 13628 -7537 13830 -7520
rect 14386 -7520 14402 -7503
rect 14832 -7503 15420 -7487
rect 14832 -7520 14848 -7503
rect 14386 -7537 14588 -7520
rect 13628 -7584 14588 -7537
rect 14646 -7537 14848 -7520
rect 15404 -7520 15420 -7503
rect 15850 -7503 16438 -7487
rect 15850 -7520 15866 -7503
rect 15404 -7537 15606 -7520
rect 14646 -7584 15606 -7537
rect 15664 -7537 15866 -7520
rect 16422 -7520 16438 -7503
rect 16868 -7503 17456 -7487
rect 16868 -7520 16884 -7503
rect 16422 -7537 16624 -7520
rect 15664 -7584 16624 -7537
rect 16682 -7537 16884 -7520
rect 17440 -7520 17456 -7503
rect 17886 -7503 18474 -7487
rect 17886 -7520 17902 -7503
rect 17440 -7537 17642 -7520
rect 16682 -7584 17642 -7537
rect 17700 -7537 17902 -7520
rect 18458 -7520 18474 -7503
rect 18904 -7503 19492 -7487
rect 18904 -7520 18920 -7503
rect 18458 -7537 18660 -7520
rect 17700 -7584 18660 -7537
rect 18718 -7537 18920 -7520
rect 19476 -7520 19492 -7503
rect 19922 -7503 20510 -7487
rect 19922 -7520 19938 -7503
rect 19476 -7537 19678 -7520
rect 18718 -7584 19678 -7537
rect 19736 -7537 19938 -7520
rect 20494 -7520 20510 -7503
rect 20940 -7503 21528 -7487
rect 20940 -7520 20956 -7503
rect 20494 -7537 20696 -7520
rect 19736 -7584 20696 -7537
rect 20754 -7537 20956 -7520
rect 21512 -7520 21528 -7503
rect 21958 -7503 22546 -7487
rect 21958 -7520 21974 -7503
rect 21512 -7537 21714 -7520
rect 20754 -7584 21714 -7537
rect 21772 -7537 21974 -7520
rect 22530 -7520 22546 -7503
rect 22530 -7537 22732 -7520
rect 21772 -7584 22732 -7537
rect 2216 -7887 3176 -7840
rect 2216 -7904 2418 -7887
rect 2402 -7921 2418 -7904
rect 2974 -7904 3176 -7887
rect 3234 -7887 4194 -7840
rect 3234 -7904 3436 -7887
rect 2974 -7921 2990 -7904
rect 2402 -7937 2990 -7921
rect 3420 -7921 3436 -7904
rect 3992 -7904 4194 -7887
rect 4252 -7887 5212 -7840
rect 4252 -7904 4454 -7887
rect 3992 -7921 4008 -7904
rect 3420 -7937 4008 -7921
rect 4438 -7921 4454 -7904
rect 5010 -7904 5212 -7887
rect 5270 -7887 6230 -7840
rect 5270 -7904 5472 -7887
rect 5010 -7921 5026 -7904
rect 4438 -7937 5026 -7921
rect 5456 -7921 5472 -7904
rect 6028 -7904 6230 -7887
rect 6028 -7921 6044 -7904
rect 5456 -7937 6044 -7921
rect 2402 -8191 2990 -8175
rect 2402 -8208 2418 -8191
rect 2216 -8225 2418 -8208
rect 2974 -8208 2990 -8191
rect 3420 -8191 4008 -8175
rect 3420 -8208 3436 -8191
rect 2974 -8225 3176 -8208
rect 2216 -8272 3176 -8225
rect 3234 -8225 3436 -8208
rect 3992 -8208 4008 -8191
rect 4438 -8191 5026 -8175
rect 4438 -8208 4454 -8191
rect 3992 -8225 4194 -8208
rect 3234 -8272 4194 -8225
rect 4252 -8225 4454 -8208
rect 5010 -8208 5026 -8191
rect 5456 -8191 6044 -8175
rect 5456 -8208 5472 -8191
rect 5010 -8225 5212 -8208
rect 4252 -8272 5212 -8225
rect 5270 -8225 5472 -8208
rect 6028 -8208 6044 -8191
rect 6028 -8225 6230 -8208
rect 5270 -8272 6230 -8225
rect 7520 -8231 8480 -8184
rect 7520 -8248 7722 -8231
rect 7706 -8265 7722 -8248
rect 8278 -8248 8480 -8231
rect 8538 -8231 9498 -8184
rect 8538 -8248 8740 -8231
rect 8278 -8265 8294 -8248
rect 7706 -8281 8294 -8265
rect 8724 -8265 8740 -8248
rect 9296 -8248 9498 -8231
rect 9556 -8231 10516 -8184
rect 9556 -8248 9758 -8231
rect 9296 -8265 9312 -8248
rect 8724 -8281 9312 -8265
rect 9742 -8265 9758 -8248
rect 10314 -8248 10516 -8231
rect 10574 -8231 11534 -8184
rect 10574 -8248 10776 -8231
rect 10314 -8265 10330 -8248
rect 9742 -8281 10330 -8265
rect 10760 -8265 10776 -8248
rect 11332 -8248 11534 -8231
rect 11592 -8231 12552 -8184
rect 11592 -8248 11794 -8231
rect 11332 -8265 11348 -8248
rect 10760 -8281 11348 -8265
rect 11778 -8265 11794 -8248
rect 12350 -8248 12552 -8231
rect 12610 -8231 13570 -8184
rect 12610 -8248 12812 -8231
rect 12350 -8265 12366 -8248
rect 11778 -8281 12366 -8265
rect 12796 -8265 12812 -8248
rect 13368 -8248 13570 -8231
rect 13628 -8231 14588 -8184
rect 13628 -8248 13830 -8231
rect 13368 -8265 13384 -8248
rect 12796 -8281 13384 -8265
rect 13814 -8265 13830 -8248
rect 14386 -8248 14588 -8231
rect 14646 -8231 15606 -8184
rect 14646 -8248 14848 -8231
rect 14386 -8265 14402 -8248
rect 13814 -8281 14402 -8265
rect 14832 -8265 14848 -8248
rect 15404 -8248 15606 -8231
rect 15664 -8231 16624 -8184
rect 15664 -8248 15866 -8231
rect 15404 -8265 15420 -8248
rect 14832 -8281 15420 -8265
rect 15850 -8265 15866 -8248
rect 16422 -8248 16624 -8231
rect 16682 -8231 17642 -8184
rect 16682 -8248 16884 -8231
rect 16422 -8265 16438 -8248
rect 15850 -8281 16438 -8265
rect 16868 -8265 16884 -8248
rect 17440 -8248 17642 -8231
rect 17700 -8231 18660 -8184
rect 17700 -8248 17902 -8231
rect 17440 -8265 17456 -8248
rect 16868 -8281 17456 -8265
rect 17886 -8265 17902 -8248
rect 18458 -8248 18660 -8231
rect 18718 -8231 19678 -8184
rect 18718 -8248 18920 -8231
rect 18458 -8265 18474 -8248
rect 17886 -8281 18474 -8265
rect 18904 -8265 18920 -8248
rect 19476 -8248 19678 -8231
rect 19736 -8231 20696 -8184
rect 19736 -8248 19938 -8231
rect 19476 -8265 19492 -8248
rect 18904 -8281 19492 -8265
rect 19922 -8265 19938 -8248
rect 20494 -8248 20696 -8231
rect 20754 -8231 21714 -8184
rect 20754 -8248 20956 -8231
rect 20494 -8265 20510 -8248
rect 19922 -8281 20510 -8265
rect 20940 -8265 20956 -8248
rect 21512 -8248 21714 -8231
rect 21772 -8231 22732 -8184
rect 21772 -8248 21974 -8231
rect 21512 -8265 21528 -8248
rect 20940 -8281 21528 -8265
rect 21958 -8265 21974 -8248
rect 22530 -8248 22732 -8231
rect 22530 -8265 22546 -8248
rect 21958 -8281 22546 -8265
rect 7706 -8759 8294 -8743
rect 7706 -8776 7722 -8759
rect 7520 -8793 7722 -8776
rect 8278 -8776 8294 -8759
rect 8724 -8759 9312 -8743
rect 8724 -8776 8740 -8759
rect 8278 -8793 8480 -8776
rect 7520 -8840 8480 -8793
rect 8538 -8793 8740 -8776
rect 9296 -8776 9312 -8759
rect 9742 -8759 10330 -8743
rect 9742 -8776 9758 -8759
rect 9296 -8793 9498 -8776
rect 8538 -8840 9498 -8793
rect 9556 -8793 9758 -8776
rect 10314 -8776 10330 -8759
rect 10760 -8759 11348 -8743
rect 10760 -8776 10776 -8759
rect 10314 -8793 10516 -8776
rect 9556 -8840 10516 -8793
rect 10574 -8793 10776 -8776
rect 11332 -8776 11348 -8759
rect 11778 -8759 12366 -8743
rect 11778 -8776 11794 -8759
rect 11332 -8793 11534 -8776
rect 10574 -8840 11534 -8793
rect 11592 -8793 11794 -8776
rect 12350 -8776 12366 -8759
rect 12796 -8759 13384 -8743
rect 12796 -8776 12812 -8759
rect 12350 -8793 12552 -8776
rect 11592 -8840 12552 -8793
rect 12610 -8793 12812 -8776
rect 13368 -8776 13384 -8759
rect 13814 -8759 14402 -8743
rect 13814 -8776 13830 -8759
rect 13368 -8793 13570 -8776
rect 12610 -8840 13570 -8793
rect 13628 -8793 13830 -8776
rect 14386 -8776 14402 -8759
rect 14832 -8759 15420 -8743
rect 14832 -8776 14848 -8759
rect 14386 -8793 14588 -8776
rect 13628 -8840 14588 -8793
rect 14646 -8793 14848 -8776
rect 15404 -8776 15420 -8759
rect 15850 -8759 16438 -8743
rect 15850 -8776 15866 -8759
rect 15404 -8793 15606 -8776
rect 14646 -8840 15606 -8793
rect 15664 -8793 15866 -8776
rect 16422 -8776 16438 -8759
rect 16868 -8759 17456 -8743
rect 16868 -8776 16884 -8759
rect 16422 -8793 16624 -8776
rect 15664 -8840 16624 -8793
rect 16682 -8793 16884 -8776
rect 17440 -8776 17456 -8759
rect 17886 -8759 18474 -8743
rect 17886 -8776 17902 -8759
rect 17440 -8793 17642 -8776
rect 16682 -8840 17642 -8793
rect 17700 -8793 17902 -8776
rect 18458 -8776 18474 -8759
rect 18904 -8759 19492 -8743
rect 18904 -8776 18920 -8759
rect 18458 -8793 18660 -8776
rect 17700 -8840 18660 -8793
rect 18718 -8793 18920 -8776
rect 19476 -8776 19492 -8759
rect 19922 -8759 20510 -8743
rect 19922 -8776 19938 -8759
rect 19476 -8793 19678 -8776
rect 18718 -8840 19678 -8793
rect 19736 -8793 19938 -8776
rect 20494 -8776 20510 -8759
rect 20940 -8759 21528 -8743
rect 20940 -8776 20956 -8759
rect 20494 -8793 20696 -8776
rect 19736 -8840 20696 -8793
rect 20754 -8793 20956 -8776
rect 21512 -8776 21528 -8759
rect 21958 -8759 22546 -8743
rect 21958 -8776 21974 -8759
rect 21512 -8793 21714 -8776
rect 20754 -8840 21714 -8793
rect 21772 -8793 21974 -8776
rect 22530 -8776 22546 -8759
rect 22530 -8793 22732 -8776
rect 21772 -8840 22732 -8793
rect 2216 -8919 3176 -8872
rect 2216 -8936 2418 -8919
rect 2402 -8953 2418 -8936
rect 2974 -8936 3176 -8919
rect 3234 -8919 4194 -8872
rect 3234 -8936 3436 -8919
rect 2974 -8953 2990 -8936
rect 2402 -8969 2990 -8953
rect 3420 -8953 3436 -8936
rect 3992 -8936 4194 -8919
rect 4252 -8919 5212 -8872
rect 4252 -8936 4454 -8919
rect 3992 -8953 4008 -8936
rect 3420 -8969 4008 -8953
rect 4438 -8953 4454 -8936
rect 5010 -8936 5212 -8919
rect 5270 -8919 6230 -8872
rect 5270 -8936 5472 -8919
rect 5010 -8953 5026 -8936
rect 4438 -8969 5026 -8953
rect 5456 -8953 5472 -8936
rect 6028 -8936 6230 -8919
rect 6028 -8953 6044 -8936
rect 5456 -8969 6044 -8953
rect 7520 -9487 8480 -9440
rect 7520 -9504 7722 -9487
rect 7706 -9521 7722 -9504
rect 8278 -9504 8480 -9487
rect 8538 -9487 9498 -9440
rect 8538 -9504 8740 -9487
rect 8278 -9521 8294 -9504
rect 7706 -9537 8294 -9521
rect 8724 -9521 8740 -9504
rect 9296 -9504 9498 -9487
rect 9556 -9487 10516 -9440
rect 9556 -9504 9758 -9487
rect 9296 -9521 9312 -9504
rect 8724 -9537 9312 -9521
rect 9742 -9521 9758 -9504
rect 10314 -9504 10516 -9487
rect 10574 -9487 11534 -9440
rect 10574 -9504 10776 -9487
rect 10314 -9521 10330 -9504
rect 9742 -9537 10330 -9521
rect 10760 -9521 10776 -9504
rect 11332 -9504 11534 -9487
rect 11592 -9487 12552 -9440
rect 11592 -9504 11794 -9487
rect 11332 -9521 11348 -9504
rect 10760 -9537 11348 -9521
rect 11778 -9521 11794 -9504
rect 12350 -9504 12552 -9487
rect 12610 -9487 13570 -9440
rect 12610 -9504 12812 -9487
rect 12350 -9521 12366 -9504
rect 11778 -9537 12366 -9521
rect 12796 -9521 12812 -9504
rect 13368 -9504 13570 -9487
rect 13628 -9487 14588 -9440
rect 13628 -9504 13830 -9487
rect 13368 -9521 13384 -9504
rect 12796 -9537 13384 -9521
rect 13814 -9521 13830 -9504
rect 14386 -9504 14588 -9487
rect 14646 -9487 15606 -9440
rect 14646 -9504 14848 -9487
rect 14386 -9521 14402 -9504
rect 13814 -9537 14402 -9521
rect 14832 -9521 14848 -9504
rect 15404 -9504 15606 -9487
rect 15664 -9487 16624 -9440
rect 15664 -9504 15866 -9487
rect 15404 -9521 15420 -9504
rect 14832 -9537 15420 -9521
rect 15850 -9521 15866 -9504
rect 16422 -9504 16624 -9487
rect 16682 -9487 17642 -9440
rect 16682 -9504 16884 -9487
rect 16422 -9521 16438 -9504
rect 15850 -9537 16438 -9521
rect 16868 -9521 16884 -9504
rect 17440 -9504 17642 -9487
rect 17700 -9487 18660 -9440
rect 17700 -9504 17902 -9487
rect 17440 -9521 17456 -9504
rect 16868 -9537 17456 -9521
rect 17886 -9521 17902 -9504
rect 18458 -9504 18660 -9487
rect 18718 -9487 19678 -9440
rect 18718 -9504 18920 -9487
rect 18458 -9521 18474 -9504
rect 17886 -9537 18474 -9521
rect 18904 -9521 18920 -9504
rect 19476 -9504 19678 -9487
rect 19736 -9487 20696 -9440
rect 19736 -9504 19938 -9487
rect 19476 -9521 19492 -9504
rect 18904 -9537 19492 -9521
rect 19922 -9521 19938 -9504
rect 20494 -9504 20696 -9487
rect 20754 -9487 21714 -9440
rect 20754 -9504 20956 -9487
rect 20494 -9521 20510 -9504
rect 19922 -9537 20510 -9521
rect 20940 -9521 20956 -9504
rect 21512 -9504 21714 -9487
rect 21772 -9487 22732 -9440
rect 21772 -9504 21974 -9487
rect 21512 -9521 21528 -9504
rect 20940 -9537 21528 -9521
rect 21958 -9521 21974 -9504
rect 22530 -9504 22732 -9487
rect 22530 -9521 22546 -9504
rect 21958 -9537 22546 -9521
rect 2814 -11964 3402 -11948
rect 2814 -11981 2830 -11964
rect 2628 -11998 2830 -11981
rect 3386 -11981 3402 -11964
rect 3832 -11964 4420 -11948
rect 3832 -11981 3848 -11964
rect 3386 -11998 3588 -11981
rect 2628 -12036 3588 -11998
rect 3646 -11998 3848 -11981
rect 4404 -11981 4420 -11964
rect 4850 -11964 5438 -11948
rect 4850 -11981 4866 -11964
rect 4404 -11998 4606 -11981
rect 3646 -12036 4606 -11998
rect 4664 -11998 4866 -11981
rect 5422 -11981 5438 -11964
rect 5868 -11964 6456 -11948
rect 5868 -11981 5884 -11964
rect 5422 -11998 5624 -11981
rect 4664 -12036 5624 -11998
rect 5682 -11998 5884 -11981
rect 6440 -11981 6456 -11964
rect 6886 -11964 7474 -11948
rect 6886 -11981 6902 -11964
rect 6440 -11998 6642 -11981
rect 5682 -12036 6642 -11998
rect 6700 -11998 6902 -11981
rect 7458 -11981 7474 -11964
rect 7904 -11964 8492 -11948
rect 7904 -11981 7920 -11964
rect 7458 -11998 7660 -11981
rect 6700 -12036 7660 -11998
rect 7718 -11998 7920 -11981
rect 8476 -11981 8492 -11964
rect 8922 -11964 9510 -11948
rect 8922 -11981 8938 -11964
rect 8476 -11998 8678 -11981
rect 7718 -12036 8678 -11998
rect 8736 -11998 8938 -11981
rect 9494 -11981 9510 -11964
rect 9940 -11964 10528 -11948
rect 9940 -11981 9956 -11964
rect 9494 -11998 9696 -11981
rect 8736 -12036 9696 -11998
rect 9754 -11998 9956 -11981
rect 10512 -11981 10528 -11964
rect 10958 -11964 11546 -11948
rect 10958 -11981 10974 -11964
rect 10512 -11998 10714 -11981
rect 9754 -12036 10714 -11998
rect 10772 -11998 10974 -11981
rect 11530 -11981 11546 -11964
rect 11976 -11964 12564 -11948
rect 11976 -11981 11992 -11964
rect 11530 -11998 11732 -11981
rect 10772 -12036 11732 -11998
rect 11790 -11998 11992 -11981
rect 12548 -11981 12564 -11964
rect 12994 -11964 13582 -11948
rect 12994 -11981 13010 -11964
rect 12548 -11998 12750 -11981
rect 11790 -12036 12750 -11998
rect 12808 -11998 13010 -11981
rect 13566 -11981 13582 -11964
rect 14012 -11964 14600 -11948
rect 14012 -11981 14028 -11964
rect 13566 -11998 13768 -11981
rect 12808 -12036 13768 -11998
rect 13826 -11998 14028 -11981
rect 14584 -11981 14600 -11964
rect 15030 -11964 15618 -11948
rect 15030 -11981 15046 -11964
rect 14584 -11998 14786 -11981
rect 13826 -12036 14786 -11998
rect 14844 -11998 15046 -11981
rect 15602 -11981 15618 -11964
rect 16048 -11964 16636 -11948
rect 16048 -11981 16064 -11964
rect 15602 -11998 15804 -11981
rect 14844 -12036 15804 -11998
rect 15862 -11998 16064 -11981
rect 16620 -11981 16636 -11964
rect 17066 -11964 17654 -11948
rect 17066 -11981 17082 -11964
rect 16620 -11998 16822 -11981
rect 15862 -12036 16822 -11998
rect 16880 -11998 17082 -11981
rect 17638 -11981 17654 -11964
rect 18084 -11964 18672 -11948
rect 18084 -11981 18100 -11964
rect 17638 -11998 17840 -11981
rect 16880 -12036 17840 -11998
rect 17898 -11998 18100 -11981
rect 18656 -11981 18672 -11964
rect 19102 -11964 19690 -11948
rect 19102 -11981 19118 -11964
rect 18656 -11998 18858 -11981
rect 17898 -12036 18858 -11998
rect 18916 -11998 19118 -11981
rect 19674 -11981 19690 -11964
rect 20120 -11964 20708 -11948
rect 20120 -11981 20136 -11964
rect 19674 -11998 19876 -11981
rect 18916 -12036 19876 -11998
rect 19934 -11998 20136 -11981
rect 20692 -11981 20708 -11964
rect 21138 -11964 21726 -11948
rect 21138 -11981 21154 -11964
rect 20692 -11998 20894 -11981
rect 19934 -12036 20894 -11998
rect 20952 -11998 21154 -11981
rect 21710 -11981 21726 -11964
rect 22156 -11964 22744 -11948
rect 22156 -11981 22172 -11964
rect 21710 -11998 21912 -11981
rect 20952 -12036 21912 -11998
rect 21970 -11998 22172 -11981
rect 22728 -11981 22744 -11964
rect 22728 -11998 22930 -11981
rect 21970 -12036 22930 -11998
rect -8952 -12440 -8364 -12424
rect -8952 -12457 -8936 -12440
rect -9138 -12474 -8936 -12457
rect -8380 -12457 -8364 -12440
rect -7934 -12440 -7346 -12424
rect -7934 -12457 -7918 -12440
rect -8380 -12474 -8178 -12457
rect -9138 -12512 -8178 -12474
rect -8120 -12474 -7918 -12457
rect -7362 -12457 -7346 -12440
rect -6916 -12440 -6328 -12424
rect -6916 -12457 -6900 -12440
rect -7362 -12474 -7160 -12457
rect -8120 -12512 -7160 -12474
rect -7102 -12474 -6900 -12457
rect -6344 -12457 -6328 -12440
rect -5898 -12440 -5310 -12424
rect -5898 -12457 -5882 -12440
rect -6344 -12474 -6142 -12457
rect -7102 -12512 -6142 -12474
rect -6084 -12474 -5882 -12457
rect -5326 -12457 -5310 -12440
rect -4880 -12440 -4292 -12424
rect -4880 -12457 -4864 -12440
rect -5326 -12474 -5124 -12457
rect -6084 -12512 -5124 -12474
rect -5066 -12474 -4864 -12457
rect -4308 -12457 -4292 -12440
rect -3862 -12440 -3274 -12424
rect -3862 -12457 -3846 -12440
rect -4308 -12474 -4106 -12457
rect -5066 -12512 -4106 -12474
rect -4048 -12474 -3846 -12457
rect -3290 -12457 -3274 -12440
rect -2844 -12440 -2256 -12424
rect -2844 -12457 -2828 -12440
rect -3290 -12474 -3088 -12457
rect -4048 -12512 -3088 -12474
rect -3030 -12474 -2828 -12457
rect -2272 -12457 -2256 -12440
rect -1826 -12440 -1238 -12424
rect -1826 -12457 -1810 -12440
rect -2272 -12474 -2070 -12457
rect -3030 -12512 -2070 -12474
rect -2012 -12474 -1810 -12457
rect -1254 -12457 -1238 -12440
rect -808 -12440 -220 -12424
rect -808 -12457 -792 -12440
rect -1254 -12474 -1052 -12457
rect -2012 -12512 -1052 -12474
rect -994 -12474 -792 -12457
rect -236 -12457 -220 -12440
rect -236 -12474 -34 -12457
rect -994 -12512 -34 -12474
rect 2628 -12674 3588 -12636
rect 2628 -12691 2830 -12674
rect 2814 -12708 2830 -12691
rect 3386 -12691 3588 -12674
rect 3646 -12674 4606 -12636
rect 3646 -12691 3848 -12674
rect 3386 -12708 3402 -12691
rect 2814 -12724 3402 -12708
rect 3832 -12708 3848 -12691
rect 4404 -12691 4606 -12674
rect 4664 -12674 5624 -12636
rect 4664 -12691 4866 -12674
rect 4404 -12708 4420 -12691
rect 3832 -12724 4420 -12708
rect 4850 -12708 4866 -12691
rect 5422 -12691 5624 -12674
rect 5682 -12674 6642 -12636
rect 5682 -12691 5884 -12674
rect 5422 -12708 5438 -12691
rect 4850 -12724 5438 -12708
rect 5868 -12708 5884 -12691
rect 6440 -12691 6642 -12674
rect 6700 -12674 7660 -12636
rect 6700 -12691 6902 -12674
rect 6440 -12708 6456 -12691
rect 5868 -12724 6456 -12708
rect 6886 -12708 6902 -12691
rect 7458 -12691 7660 -12674
rect 7718 -12674 8678 -12636
rect 7718 -12691 7920 -12674
rect 7458 -12708 7474 -12691
rect 6886 -12724 7474 -12708
rect 7904 -12708 7920 -12691
rect 8476 -12691 8678 -12674
rect 8736 -12674 9696 -12636
rect 8736 -12691 8938 -12674
rect 8476 -12708 8492 -12691
rect 7904 -12724 8492 -12708
rect 8922 -12708 8938 -12691
rect 9494 -12691 9696 -12674
rect 9754 -12674 10714 -12636
rect 9754 -12691 9956 -12674
rect 9494 -12708 9510 -12691
rect 8922 -12724 9510 -12708
rect 9940 -12708 9956 -12691
rect 10512 -12691 10714 -12674
rect 10772 -12674 11732 -12636
rect 10772 -12691 10974 -12674
rect 10512 -12708 10528 -12691
rect 9940 -12724 10528 -12708
rect 10958 -12708 10974 -12691
rect 11530 -12691 11732 -12674
rect 11790 -12674 12750 -12636
rect 11790 -12691 11992 -12674
rect 11530 -12708 11546 -12691
rect 10958 -12724 11546 -12708
rect 11976 -12708 11992 -12691
rect 12548 -12691 12750 -12674
rect 12808 -12674 13768 -12636
rect 12808 -12691 13010 -12674
rect 12548 -12708 12564 -12691
rect 11976 -12724 12564 -12708
rect 12994 -12708 13010 -12691
rect 13566 -12691 13768 -12674
rect 13826 -12674 14786 -12636
rect 13826 -12691 14028 -12674
rect 13566 -12708 13582 -12691
rect 12994 -12724 13582 -12708
rect 14012 -12708 14028 -12691
rect 14584 -12691 14786 -12674
rect 14844 -12674 15804 -12636
rect 14844 -12691 15046 -12674
rect 14584 -12708 14600 -12691
rect 14012 -12724 14600 -12708
rect 15030 -12708 15046 -12691
rect 15602 -12691 15804 -12674
rect 15862 -12674 16822 -12636
rect 15862 -12691 16064 -12674
rect 15602 -12708 15618 -12691
rect 15030 -12724 15618 -12708
rect 16048 -12708 16064 -12691
rect 16620 -12691 16822 -12674
rect 16880 -12674 17840 -12636
rect 16880 -12691 17082 -12674
rect 16620 -12708 16636 -12691
rect 16048 -12724 16636 -12708
rect 17066 -12708 17082 -12691
rect 17638 -12691 17840 -12674
rect 17898 -12674 18858 -12636
rect 17898 -12691 18100 -12674
rect 17638 -12708 17654 -12691
rect 17066 -12724 17654 -12708
rect 18084 -12708 18100 -12691
rect 18656 -12691 18858 -12674
rect 18916 -12674 19876 -12636
rect 18916 -12691 19118 -12674
rect 18656 -12708 18672 -12691
rect 18084 -12724 18672 -12708
rect 19102 -12708 19118 -12691
rect 19674 -12691 19876 -12674
rect 19934 -12674 20894 -12636
rect 19934 -12691 20136 -12674
rect 19674 -12708 19690 -12691
rect 19102 -12724 19690 -12708
rect 20120 -12708 20136 -12691
rect 20692 -12691 20894 -12674
rect 20952 -12674 21912 -12636
rect 20952 -12691 21154 -12674
rect 20692 -12708 20708 -12691
rect 20120 -12724 20708 -12708
rect 21138 -12708 21154 -12691
rect 21710 -12691 21912 -12674
rect 21970 -12674 22930 -12636
rect 21970 -12691 22172 -12674
rect 21710 -12708 21726 -12691
rect 21138 -12724 21726 -12708
rect 22156 -12708 22172 -12691
rect 22728 -12691 22930 -12674
rect 22728 -12708 22744 -12691
rect 22156 -12724 22744 -12708
rect 2814 -12782 3402 -12766
rect 2814 -12799 2830 -12782
rect 2628 -12816 2830 -12799
rect 3386 -12799 3402 -12782
rect 3832 -12782 4420 -12766
rect 3832 -12799 3848 -12782
rect 3386 -12816 3588 -12799
rect 2628 -12854 3588 -12816
rect 3646 -12816 3848 -12799
rect 4404 -12799 4420 -12782
rect 4850 -12782 5438 -12766
rect 4850 -12799 4866 -12782
rect 4404 -12816 4606 -12799
rect 3646 -12854 4606 -12816
rect 4664 -12816 4866 -12799
rect 5422 -12799 5438 -12782
rect 5868 -12782 6456 -12766
rect 5868 -12799 5884 -12782
rect 5422 -12816 5624 -12799
rect 4664 -12854 5624 -12816
rect 5682 -12816 5884 -12799
rect 6440 -12799 6456 -12782
rect 6886 -12782 7474 -12766
rect 6886 -12799 6902 -12782
rect 6440 -12816 6642 -12799
rect 5682 -12854 6642 -12816
rect 6700 -12816 6902 -12799
rect 7458 -12799 7474 -12782
rect 7904 -12782 8492 -12766
rect 7904 -12799 7920 -12782
rect 7458 -12816 7660 -12799
rect 6700 -12854 7660 -12816
rect 7718 -12816 7920 -12799
rect 8476 -12799 8492 -12782
rect 8922 -12782 9510 -12766
rect 8922 -12799 8938 -12782
rect 8476 -12816 8678 -12799
rect 7718 -12854 8678 -12816
rect 8736 -12816 8938 -12799
rect 9494 -12799 9510 -12782
rect 9940 -12782 10528 -12766
rect 9940 -12799 9956 -12782
rect 9494 -12816 9696 -12799
rect 8736 -12854 9696 -12816
rect 9754 -12816 9956 -12799
rect 10512 -12799 10528 -12782
rect 10958 -12782 11546 -12766
rect 10958 -12799 10974 -12782
rect 10512 -12816 10714 -12799
rect 9754 -12854 10714 -12816
rect 10772 -12816 10974 -12799
rect 11530 -12799 11546 -12782
rect 11976 -12782 12564 -12766
rect 11976 -12799 11992 -12782
rect 11530 -12816 11732 -12799
rect 10772 -12854 11732 -12816
rect 11790 -12816 11992 -12799
rect 12548 -12799 12564 -12782
rect 12994 -12782 13582 -12766
rect 12994 -12799 13010 -12782
rect 12548 -12816 12750 -12799
rect 11790 -12854 12750 -12816
rect 12808 -12816 13010 -12799
rect 13566 -12799 13582 -12782
rect 14012 -12782 14600 -12766
rect 14012 -12799 14028 -12782
rect 13566 -12816 13768 -12799
rect 12808 -12854 13768 -12816
rect 13826 -12816 14028 -12799
rect 14584 -12799 14600 -12782
rect 15030 -12782 15618 -12766
rect 15030 -12799 15046 -12782
rect 14584 -12816 14786 -12799
rect 13826 -12854 14786 -12816
rect 14844 -12816 15046 -12799
rect 15602 -12799 15618 -12782
rect 16048 -12782 16636 -12766
rect 16048 -12799 16064 -12782
rect 15602 -12816 15804 -12799
rect 14844 -12854 15804 -12816
rect 15862 -12816 16064 -12799
rect 16620 -12799 16636 -12782
rect 17066 -12782 17654 -12766
rect 17066 -12799 17082 -12782
rect 16620 -12816 16822 -12799
rect 15862 -12854 16822 -12816
rect 16880 -12816 17082 -12799
rect 17638 -12799 17654 -12782
rect 18084 -12782 18672 -12766
rect 18084 -12799 18100 -12782
rect 17638 -12816 17840 -12799
rect 16880 -12854 17840 -12816
rect 17898 -12816 18100 -12799
rect 18656 -12799 18672 -12782
rect 19102 -12782 19690 -12766
rect 19102 -12799 19118 -12782
rect 18656 -12816 18858 -12799
rect 17898 -12854 18858 -12816
rect 18916 -12816 19118 -12799
rect 19674 -12799 19690 -12782
rect 20120 -12782 20708 -12766
rect 20120 -12799 20136 -12782
rect 19674 -12816 19876 -12799
rect 18916 -12854 19876 -12816
rect 19934 -12816 20136 -12799
rect 20692 -12799 20708 -12782
rect 21138 -12782 21726 -12766
rect 21138 -12799 21154 -12782
rect 20692 -12816 20894 -12799
rect 19934 -12854 20894 -12816
rect 20952 -12816 21154 -12799
rect 21710 -12799 21726 -12782
rect 22156 -12782 22744 -12766
rect 22156 -12799 22172 -12782
rect 21710 -12816 21912 -12799
rect 20952 -12854 21912 -12816
rect 21970 -12816 22172 -12799
rect 22728 -12799 22744 -12782
rect 22728 -12816 22930 -12799
rect 21970 -12854 22930 -12816
rect -9138 -13150 -8178 -13112
rect -9138 -13167 -8936 -13150
rect -8952 -13184 -8936 -13167
rect -8380 -13167 -8178 -13150
rect -8120 -13150 -7160 -13112
rect -8120 -13167 -7918 -13150
rect -8380 -13184 -8364 -13167
rect -8952 -13200 -8364 -13184
rect -7934 -13184 -7918 -13167
rect -7362 -13167 -7160 -13150
rect -7102 -13150 -6142 -13112
rect -7102 -13167 -6900 -13150
rect -7362 -13184 -7346 -13167
rect -7934 -13200 -7346 -13184
rect -8952 -13258 -8364 -13242
rect -8952 -13275 -8936 -13258
rect -9138 -13292 -8936 -13275
rect -8380 -13275 -8364 -13258
rect -6916 -13184 -6900 -13167
rect -6344 -13167 -6142 -13150
rect -6084 -13150 -5124 -13112
rect -6084 -13167 -5882 -13150
rect -6344 -13184 -6328 -13167
rect -6916 -13200 -6328 -13184
rect -7934 -13258 -7346 -13242
rect -7934 -13275 -7918 -13258
rect -8380 -13292 -8178 -13275
rect -9138 -13330 -8178 -13292
rect -8120 -13292 -7918 -13275
rect -7362 -13275 -7346 -13258
rect -5898 -13184 -5882 -13167
rect -5326 -13167 -5124 -13150
rect -5066 -13150 -4106 -13112
rect -5066 -13167 -4864 -13150
rect -5326 -13184 -5310 -13167
rect -5898 -13200 -5310 -13184
rect -6916 -13258 -6328 -13242
rect -6916 -13275 -6900 -13258
rect -7362 -13292 -7160 -13275
rect -8120 -13330 -7160 -13292
rect -7102 -13292 -6900 -13275
rect -6344 -13275 -6328 -13258
rect -4880 -13184 -4864 -13167
rect -4308 -13167 -4106 -13150
rect -4048 -13150 -3088 -13112
rect -4048 -13167 -3846 -13150
rect -4308 -13184 -4292 -13167
rect -4880 -13200 -4292 -13184
rect -5898 -13258 -5310 -13242
rect -5898 -13275 -5882 -13258
rect -6344 -13292 -6142 -13275
rect -7102 -13330 -6142 -13292
rect -6084 -13292 -5882 -13275
rect -5326 -13275 -5310 -13258
rect -3862 -13184 -3846 -13167
rect -3290 -13167 -3088 -13150
rect -3030 -13150 -2070 -13112
rect -3030 -13167 -2828 -13150
rect -3290 -13184 -3274 -13167
rect -3862 -13200 -3274 -13184
rect -4880 -13258 -4292 -13242
rect -4880 -13275 -4864 -13258
rect -5326 -13292 -5124 -13275
rect -6084 -13330 -5124 -13292
rect -5066 -13292 -4864 -13275
rect -4308 -13275 -4292 -13258
rect -2844 -13184 -2828 -13167
rect -2272 -13167 -2070 -13150
rect -2012 -13150 -1052 -13112
rect -2012 -13167 -1810 -13150
rect -2272 -13184 -2256 -13167
rect -2844 -13200 -2256 -13184
rect -3862 -13258 -3274 -13242
rect -3862 -13275 -3846 -13258
rect -4308 -13292 -4106 -13275
rect -5066 -13330 -4106 -13292
rect -4048 -13292 -3846 -13275
rect -3290 -13275 -3274 -13258
rect -1826 -13184 -1810 -13167
rect -1254 -13167 -1052 -13150
rect -994 -13150 -34 -13112
rect -994 -13167 -792 -13150
rect -1254 -13184 -1238 -13167
rect -1826 -13200 -1238 -13184
rect -2844 -13258 -2256 -13242
rect -2844 -13275 -2828 -13258
rect -3290 -13292 -3088 -13275
rect -4048 -13330 -3088 -13292
rect -3030 -13292 -2828 -13275
rect -2272 -13275 -2256 -13258
rect -808 -13184 -792 -13167
rect -236 -13167 -34 -13150
rect -236 -13184 -220 -13167
rect -808 -13200 -220 -13184
rect -1826 -13258 -1238 -13242
rect -1826 -13275 -1810 -13258
rect -2272 -13292 -2070 -13275
rect -3030 -13330 -2070 -13292
rect -2012 -13292 -1810 -13275
rect -1254 -13275 -1238 -13258
rect -808 -13258 -220 -13242
rect -808 -13275 -792 -13258
rect -1254 -13292 -1052 -13275
rect -2012 -13330 -1052 -13292
rect -994 -13292 -792 -13275
rect -236 -13275 -220 -13258
rect -236 -13292 -34 -13275
rect -994 -13330 -34 -13292
rect 2628 -13492 3588 -13454
rect 2628 -13509 2830 -13492
rect 2814 -13526 2830 -13509
rect 3386 -13509 3588 -13492
rect 3646 -13492 4606 -13454
rect 3646 -13509 3848 -13492
rect 3386 -13526 3402 -13509
rect 2814 -13542 3402 -13526
rect 3832 -13526 3848 -13509
rect 4404 -13509 4606 -13492
rect 4664 -13492 5624 -13454
rect 4664 -13509 4866 -13492
rect 4404 -13526 4420 -13509
rect 3832 -13542 4420 -13526
rect 4850 -13526 4866 -13509
rect 5422 -13509 5624 -13492
rect 5682 -13492 6642 -13454
rect 5682 -13509 5884 -13492
rect 5422 -13526 5438 -13509
rect 4850 -13542 5438 -13526
rect 5868 -13526 5884 -13509
rect 6440 -13509 6642 -13492
rect 6700 -13492 7660 -13454
rect 6700 -13509 6902 -13492
rect 6440 -13526 6456 -13509
rect 5868 -13542 6456 -13526
rect 6886 -13526 6902 -13509
rect 7458 -13509 7660 -13492
rect 7718 -13492 8678 -13454
rect 7718 -13509 7920 -13492
rect 7458 -13526 7474 -13509
rect 6886 -13542 7474 -13526
rect 7904 -13526 7920 -13509
rect 8476 -13509 8678 -13492
rect 8736 -13492 9696 -13454
rect 8736 -13509 8938 -13492
rect 8476 -13526 8492 -13509
rect 7904 -13542 8492 -13526
rect 8922 -13526 8938 -13509
rect 9494 -13509 9696 -13492
rect 9754 -13492 10714 -13454
rect 9754 -13509 9956 -13492
rect 9494 -13526 9510 -13509
rect 8922 -13542 9510 -13526
rect 9940 -13526 9956 -13509
rect 10512 -13509 10714 -13492
rect 10772 -13492 11732 -13454
rect 10772 -13509 10974 -13492
rect 10512 -13526 10528 -13509
rect 9940 -13542 10528 -13526
rect 10958 -13526 10974 -13509
rect 11530 -13509 11732 -13492
rect 11790 -13492 12750 -13454
rect 11790 -13509 11992 -13492
rect 11530 -13526 11546 -13509
rect 10958 -13542 11546 -13526
rect 11976 -13526 11992 -13509
rect 12548 -13509 12750 -13492
rect 12808 -13492 13768 -13454
rect 12808 -13509 13010 -13492
rect 12548 -13526 12564 -13509
rect 11976 -13542 12564 -13526
rect 12994 -13526 13010 -13509
rect 13566 -13509 13768 -13492
rect 13826 -13492 14786 -13454
rect 13826 -13509 14028 -13492
rect 13566 -13526 13582 -13509
rect 12994 -13542 13582 -13526
rect 14012 -13526 14028 -13509
rect 14584 -13509 14786 -13492
rect 14844 -13492 15804 -13454
rect 14844 -13509 15046 -13492
rect 14584 -13526 14600 -13509
rect 14012 -13542 14600 -13526
rect 15030 -13526 15046 -13509
rect 15602 -13509 15804 -13492
rect 15862 -13492 16822 -13454
rect 15862 -13509 16064 -13492
rect 15602 -13526 15618 -13509
rect 15030 -13542 15618 -13526
rect 16048 -13526 16064 -13509
rect 16620 -13509 16822 -13492
rect 16880 -13492 17840 -13454
rect 16880 -13509 17082 -13492
rect 16620 -13526 16636 -13509
rect 16048 -13542 16636 -13526
rect 17066 -13526 17082 -13509
rect 17638 -13509 17840 -13492
rect 17898 -13492 18858 -13454
rect 17898 -13509 18100 -13492
rect 17638 -13526 17654 -13509
rect 17066 -13542 17654 -13526
rect 18084 -13526 18100 -13509
rect 18656 -13509 18858 -13492
rect 18916 -13492 19876 -13454
rect 18916 -13509 19118 -13492
rect 18656 -13526 18672 -13509
rect 18084 -13542 18672 -13526
rect 19102 -13526 19118 -13509
rect 19674 -13509 19876 -13492
rect 19934 -13492 20894 -13454
rect 19934 -13509 20136 -13492
rect 19674 -13526 19690 -13509
rect 19102 -13542 19690 -13526
rect 20120 -13526 20136 -13509
rect 20692 -13509 20894 -13492
rect 20952 -13492 21912 -13454
rect 20952 -13509 21154 -13492
rect 20692 -13526 20708 -13509
rect 20120 -13542 20708 -13526
rect 21138 -13526 21154 -13509
rect 21710 -13509 21912 -13492
rect 21970 -13492 22930 -13454
rect 21970 -13509 22172 -13492
rect 21710 -13526 21726 -13509
rect 21138 -13542 21726 -13526
rect 22156 -13526 22172 -13509
rect 22728 -13509 22930 -13492
rect 22728 -13526 22744 -13509
rect 22156 -13542 22744 -13526
rect -9138 -13968 -8178 -13930
rect -9138 -13985 -8936 -13968
rect -8952 -14002 -8936 -13985
rect -8380 -13985 -8178 -13968
rect -8120 -13968 -7160 -13930
rect -8120 -13985 -7918 -13968
rect -8380 -14002 -8364 -13985
rect -8952 -14018 -8364 -14002
rect -7934 -14002 -7918 -13985
rect -7362 -13985 -7160 -13968
rect -7102 -13968 -6142 -13930
rect -7102 -13985 -6900 -13968
rect -7362 -14002 -7346 -13985
rect -7934 -14018 -7346 -14002
rect -8952 -14076 -8364 -14060
rect -8952 -14093 -8936 -14076
rect -9138 -14110 -8936 -14093
rect -8380 -14093 -8364 -14076
rect -6916 -14002 -6900 -13985
rect -6344 -13985 -6142 -13968
rect -6084 -13968 -5124 -13930
rect -6084 -13985 -5882 -13968
rect -6344 -14002 -6328 -13985
rect -6916 -14018 -6328 -14002
rect -7934 -14076 -7346 -14060
rect -7934 -14093 -7918 -14076
rect -8380 -14110 -8178 -14093
rect -9138 -14148 -8178 -14110
rect -8120 -14110 -7918 -14093
rect -7362 -14093 -7346 -14076
rect -5898 -14002 -5882 -13985
rect -5326 -13985 -5124 -13968
rect -5066 -13968 -4106 -13930
rect -5066 -13985 -4864 -13968
rect -5326 -14002 -5310 -13985
rect -5898 -14018 -5310 -14002
rect -6916 -14076 -6328 -14060
rect -6916 -14093 -6900 -14076
rect -7362 -14110 -7160 -14093
rect -8120 -14148 -7160 -14110
rect -7102 -14110 -6900 -14093
rect -6344 -14093 -6328 -14076
rect -4880 -14002 -4864 -13985
rect -4308 -13985 -4106 -13968
rect -4048 -13968 -3088 -13930
rect -4048 -13985 -3846 -13968
rect -4308 -14002 -4292 -13985
rect -4880 -14018 -4292 -14002
rect -5898 -14076 -5310 -14060
rect -5898 -14093 -5882 -14076
rect -6344 -14110 -6142 -14093
rect -7102 -14148 -6142 -14110
rect -6084 -14110 -5882 -14093
rect -5326 -14093 -5310 -14076
rect -3862 -14002 -3846 -13985
rect -3290 -13985 -3088 -13968
rect -3030 -13968 -2070 -13930
rect -3030 -13985 -2828 -13968
rect -3290 -14002 -3274 -13985
rect -3862 -14018 -3274 -14002
rect -4880 -14076 -4292 -14060
rect -4880 -14093 -4864 -14076
rect -5326 -14110 -5124 -14093
rect -6084 -14148 -5124 -14110
rect -5066 -14110 -4864 -14093
rect -4308 -14093 -4292 -14076
rect -2844 -14002 -2828 -13985
rect -2272 -13985 -2070 -13968
rect -2012 -13968 -1052 -13930
rect -2012 -13985 -1810 -13968
rect -2272 -14002 -2256 -13985
rect -2844 -14018 -2256 -14002
rect -3862 -14076 -3274 -14060
rect -3862 -14093 -3846 -14076
rect -4308 -14110 -4106 -14093
rect -5066 -14148 -4106 -14110
rect -4048 -14110 -3846 -14093
rect -3290 -14093 -3274 -14076
rect -1826 -14002 -1810 -13985
rect -1254 -13985 -1052 -13968
rect -994 -13968 -34 -13930
rect -994 -13985 -792 -13968
rect -1254 -14002 -1238 -13985
rect -1826 -14018 -1238 -14002
rect -2844 -14076 -2256 -14060
rect -2844 -14093 -2828 -14076
rect -3290 -14110 -3088 -14093
rect -4048 -14148 -3088 -14110
rect -3030 -14110 -2828 -14093
rect -2272 -14093 -2256 -14076
rect -808 -14002 -792 -13985
rect -236 -13985 -34 -13968
rect -236 -14002 -220 -13985
rect -808 -14018 -220 -14002
rect -1826 -14076 -1238 -14060
rect -1826 -14093 -1810 -14076
rect -2272 -14110 -2070 -14093
rect -3030 -14148 -2070 -14110
rect -2012 -14110 -1810 -14093
rect -1254 -14093 -1238 -14076
rect -808 -14076 -220 -14060
rect -808 -14093 -792 -14076
rect -1254 -14110 -1052 -14093
rect -2012 -14148 -1052 -14110
rect -994 -14110 -792 -14093
rect -236 -14093 -220 -14076
rect -236 -14110 -34 -14093
rect -994 -14148 -34 -14110
rect 2814 -14160 3402 -14144
rect 2814 -14177 2830 -14160
rect 2628 -14194 2830 -14177
rect 3386 -14177 3402 -14160
rect 3832 -14160 4420 -14144
rect 3832 -14177 3848 -14160
rect 3386 -14194 3588 -14177
rect 2628 -14232 3588 -14194
rect 3646 -14194 3848 -14177
rect 4404 -14177 4420 -14160
rect 4850 -14160 5438 -14144
rect 4850 -14177 4866 -14160
rect 4404 -14194 4606 -14177
rect 3646 -14232 4606 -14194
rect 4664 -14194 4866 -14177
rect 5422 -14177 5438 -14160
rect 5868 -14160 6456 -14144
rect 5868 -14177 5884 -14160
rect 5422 -14194 5624 -14177
rect 4664 -14232 5624 -14194
rect 5682 -14194 5884 -14177
rect 6440 -14177 6456 -14160
rect 6886 -14160 7474 -14144
rect 6886 -14177 6902 -14160
rect 6440 -14194 6642 -14177
rect 5682 -14232 6642 -14194
rect 6700 -14194 6902 -14177
rect 7458 -14177 7474 -14160
rect 7904 -14160 8492 -14144
rect 7904 -14177 7920 -14160
rect 7458 -14194 7660 -14177
rect 6700 -14232 7660 -14194
rect 7718 -14194 7920 -14177
rect 8476 -14177 8492 -14160
rect 8922 -14160 9510 -14144
rect 8922 -14177 8938 -14160
rect 8476 -14194 8678 -14177
rect 7718 -14232 8678 -14194
rect 8736 -14194 8938 -14177
rect 9494 -14177 9510 -14160
rect 9940 -14160 10528 -14144
rect 9940 -14177 9956 -14160
rect 9494 -14194 9696 -14177
rect 8736 -14232 9696 -14194
rect 9754 -14194 9956 -14177
rect 10512 -14177 10528 -14160
rect 10958 -14160 11546 -14144
rect 10958 -14177 10974 -14160
rect 10512 -14194 10714 -14177
rect 9754 -14232 10714 -14194
rect 10772 -14194 10974 -14177
rect 11530 -14177 11546 -14160
rect 11976 -14160 12564 -14144
rect 11976 -14177 11992 -14160
rect 11530 -14194 11732 -14177
rect 10772 -14232 11732 -14194
rect 11790 -14194 11992 -14177
rect 12548 -14177 12564 -14160
rect 12994 -14160 13582 -14144
rect 12994 -14177 13010 -14160
rect 12548 -14194 12750 -14177
rect 11790 -14232 12750 -14194
rect 12808 -14194 13010 -14177
rect 13566 -14177 13582 -14160
rect 14012 -14160 14600 -14144
rect 14012 -14177 14028 -14160
rect 13566 -14194 13768 -14177
rect 12808 -14232 13768 -14194
rect 13826 -14194 14028 -14177
rect 14584 -14177 14600 -14160
rect 15030 -14160 15618 -14144
rect 15030 -14177 15046 -14160
rect 14584 -14194 14786 -14177
rect 13826 -14232 14786 -14194
rect 14844 -14194 15046 -14177
rect 15602 -14177 15618 -14160
rect 16048 -14160 16636 -14144
rect 16048 -14177 16064 -14160
rect 15602 -14194 15804 -14177
rect 14844 -14232 15804 -14194
rect 15862 -14194 16064 -14177
rect 16620 -14177 16636 -14160
rect 17066 -14160 17654 -14144
rect 17066 -14177 17082 -14160
rect 16620 -14194 16822 -14177
rect 15862 -14232 16822 -14194
rect 16880 -14194 17082 -14177
rect 17638 -14177 17654 -14160
rect 18084 -14160 18672 -14144
rect 18084 -14177 18100 -14160
rect 17638 -14194 17840 -14177
rect 16880 -14232 17840 -14194
rect 17898 -14194 18100 -14177
rect 18656 -14177 18672 -14160
rect 19102 -14160 19690 -14144
rect 19102 -14177 19118 -14160
rect 18656 -14194 18858 -14177
rect 17898 -14232 18858 -14194
rect 18916 -14194 19118 -14177
rect 19674 -14177 19690 -14160
rect 20120 -14160 20708 -14144
rect 20120 -14177 20136 -14160
rect 19674 -14194 19876 -14177
rect 18916 -14232 19876 -14194
rect 19934 -14194 20136 -14177
rect 20692 -14177 20708 -14160
rect 21138 -14160 21726 -14144
rect 21138 -14177 21154 -14160
rect 20692 -14194 20894 -14177
rect 19934 -14232 20894 -14194
rect 20952 -14194 21154 -14177
rect 21710 -14177 21726 -14160
rect 22156 -14160 22744 -14144
rect 22156 -14177 22172 -14160
rect 21710 -14194 21912 -14177
rect 20952 -14232 21912 -14194
rect 21970 -14194 22172 -14177
rect 22728 -14177 22744 -14160
rect 22728 -14194 22930 -14177
rect 21970 -14232 22930 -14194
rect -9138 -14786 -8178 -14748
rect -9138 -14803 -8936 -14786
rect -8952 -14820 -8936 -14803
rect -8380 -14803 -8178 -14786
rect -8120 -14786 -7160 -14748
rect -8120 -14803 -7918 -14786
rect -8380 -14820 -8364 -14803
rect -8952 -14836 -8364 -14820
rect -7934 -14820 -7918 -14803
rect -7362 -14803 -7160 -14786
rect -7102 -14786 -6142 -14748
rect -7102 -14803 -6900 -14786
rect -7362 -14820 -7346 -14803
rect -7934 -14836 -7346 -14820
rect -8952 -14894 -8364 -14878
rect -8952 -14911 -8936 -14894
rect -9138 -14928 -8936 -14911
rect -8380 -14911 -8364 -14894
rect -6916 -14820 -6900 -14803
rect -6344 -14803 -6142 -14786
rect -6084 -14786 -5124 -14748
rect -6084 -14803 -5882 -14786
rect -6344 -14820 -6328 -14803
rect -6916 -14836 -6328 -14820
rect -7934 -14894 -7346 -14878
rect -7934 -14911 -7918 -14894
rect -8380 -14928 -8178 -14911
rect -9138 -14966 -8178 -14928
rect -8120 -14928 -7918 -14911
rect -7362 -14911 -7346 -14894
rect -5898 -14820 -5882 -14803
rect -5326 -14803 -5124 -14786
rect -5066 -14786 -4106 -14748
rect -5066 -14803 -4864 -14786
rect -5326 -14820 -5310 -14803
rect -5898 -14836 -5310 -14820
rect -6916 -14894 -6328 -14878
rect -6916 -14911 -6900 -14894
rect -7362 -14928 -7160 -14911
rect -8120 -14966 -7160 -14928
rect -7102 -14928 -6900 -14911
rect -6344 -14911 -6328 -14894
rect -4880 -14820 -4864 -14803
rect -4308 -14803 -4106 -14786
rect -4048 -14786 -3088 -14748
rect -4048 -14803 -3846 -14786
rect -4308 -14820 -4292 -14803
rect -4880 -14836 -4292 -14820
rect -5898 -14894 -5310 -14878
rect -5898 -14911 -5882 -14894
rect -6344 -14928 -6142 -14911
rect -7102 -14966 -6142 -14928
rect -6084 -14928 -5882 -14911
rect -5326 -14911 -5310 -14894
rect -3862 -14820 -3846 -14803
rect -3290 -14803 -3088 -14786
rect -3030 -14786 -2070 -14748
rect -3030 -14803 -2828 -14786
rect -3290 -14820 -3274 -14803
rect -3862 -14836 -3274 -14820
rect -4880 -14894 -4292 -14878
rect -4880 -14911 -4864 -14894
rect -5326 -14928 -5124 -14911
rect -6084 -14966 -5124 -14928
rect -5066 -14928 -4864 -14911
rect -4308 -14911 -4292 -14894
rect -2844 -14820 -2828 -14803
rect -2272 -14803 -2070 -14786
rect -2012 -14786 -1052 -14748
rect -2012 -14803 -1810 -14786
rect -2272 -14820 -2256 -14803
rect -2844 -14836 -2256 -14820
rect -3862 -14894 -3274 -14878
rect -3862 -14911 -3846 -14894
rect -4308 -14928 -4106 -14911
rect -5066 -14966 -4106 -14928
rect -4048 -14928 -3846 -14911
rect -3290 -14911 -3274 -14894
rect -1826 -14820 -1810 -14803
rect -1254 -14803 -1052 -14786
rect -994 -14786 -34 -14748
rect -994 -14803 -792 -14786
rect -1254 -14820 -1238 -14803
rect -1826 -14836 -1238 -14820
rect -2844 -14894 -2256 -14878
rect -2844 -14911 -2828 -14894
rect -3290 -14928 -3088 -14911
rect -4048 -14966 -3088 -14928
rect -3030 -14928 -2828 -14911
rect -2272 -14911 -2256 -14894
rect -808 -14820 -792 -14803
rect -236 -14803 -34 -14786
rect -236 -14820 -220 -14803
rect -808 -14836 -220 -14820
rect -1826 -14894 -1238 -14878
rect -1826 -14911 -1810 -14894
rect -2272 -14928 -2070 -14911
rect -3030 -14966 -2070 -14928
rect -2012 -14928 -1810 -14911
rect -1254 -14911 -1238 -14894
rect -808 -14894 -220 -14878
rect -808 -14911 -792 -14894
rect -1254 -14928 -1052 -14911
rect -2012 -14966 -1052 -14928
rect -994 -14928 -792 -14911
rect -236 -14911 -220 -14894
rect 2628 -14870 3588 -14832
rect 2628 -14887 2830 -14870
rect 2814 -14904 2830 -14887
rect 3386 -14887 3588 -14870
rect 3646 -14870 4606 -14832
rect 3646 -14887 3848 -14870
rect 3386 -14904 3402 -14887
rect -236 -14928 -34 -14911
rect 2814 -14920 3402 -14904
rect 3832 -14904 3848 -14887
rect 4404 -14887 4606 -14870
rect 4664 -14870 5624 -14832
rect 4664 -14887 4866 -14870
rect 4404 -14904 4420 -14887
rect 3832 -14920 4420 -14904
rect 4850 -14904 4866 -14887
rect 5422 -14887 5624 -14870
rect 5682 -14870 6642 -14832
rect 5682 -14887 5884 -14870
rect 5422 -14904 5438 -14887
rect 4850 -14920 5438 -14904
rect 5868 -14904 5884 -14887
rect 6440 -14887 6642 -14870
rect 6700 -14870 7660 -14832
rect 6700 -14887 6902 -14870
rect 6440 -14904 6456 -14887
rect 5868 -14920 6456 -14904
rect 6886 -14904 6902 -14887
rect 7458 -14887 7660 -14870
rect 7718 -14870 8678 -14832
rect 7718 -14887 7920 -14870
rect 7458 -14904 7474 -14887
rect 6886 -14920 7474 -14904
rect 7904 -14904 7920 -14887
rect 8476 -14887 8678 -14870
rect 8736 -14870 9696 -14832
rect 8736 -14887 8938 -14870
rect 8476 -14904 8492 -14887
rect 7904 -14920 8492 -14904
rect 8922 -14904 8938 -14887
rect 9494 -14887 9696 -14870
rect 9754 -14870 10714 -14832
rect 9754 -14887 9956 -14870
rect 9494 -14904 9510 -14887
rect 8922 -14920 9510 -14904
rect 9940 -14904 9956 -14887
rect 10512 -14887 10714 -14870
rect 10772 -14870 11732 -14832
rect 10772 -14887 10974 -14870
rect 10512 -14904 10528 -14887
rect 9940 -14920 10528 -14904
rect 10958 -14904 10974 -14887
rect 11530 -14887 11732 -14870
rect 11790 -14870 12750 -14832
rect 11790 -14887 11992 -14870
rect 11530 -14904 11546 -14887
rect 10958 -14920 11546 -14904
rect 11976 -14904 11992 -14887
rect 12548 -14887 12750 -14870
rect 12808 -14870 13768 -14832
rect 12808 -14887 13010 -14870
rect 12548 -14904 12564 -14887
rect 11976 -14920 12564 -14904
rect 12994 -14904 13010 -14887
rect 13566 -14887 13768 -14870
rect 13826 -14870 14786 -14832
rect 13826 -14887 14028 -14870
rect 13566 -14904 13582 -14887
rect 12994 -14920 13582 -14904
rect 14012 -14904 14028 -14887
rect 14584 -14887 14786 -14870
rect 14844 -14870 15804 -14832
rect 14844 -14887 15046 -14870
rect 14584 -14904 14600 -14887
rect 14012 -14920 14600 -14904
rect 15030 -14904 15046 -14887
rect 15602 -14887 15804 -14870
rect 15862 -14870 16822 -14832
rect 15862 -14887 16064 -14870
rect 15602 -14904 15618 -14887
rect 15030 -14920 15618 -14904
rect 16048 -14904 16064 -14887
rect 16620 -14887 16822 -14870
rect 16880 -14870 17840 -14832
rect 16880 -14887 17082 -14870
rect 16620 -14904 16636 -14887
rect 16048 -14920 16636 -14904
rect 17066 -14904 17082 -14887
rect 17638 -14887 17840 -14870
rect 17898 -14870 18858 -14832
rect 17898 -14887 18100 -14870
rect 17638 -14904 17654 -14887
rect 17066 -14920 17654 -14904
rect 18084 -14904 18100 -14887
rect 18656 -14887 18858 -14870
rect 18916 -14870 19876 -14832
rect 18916 -14887 19118 -14870
rect 18656 -14904 18672 -14887
rect 18084 -14920 18672 -14904
rect 19102 -14904 19118 -14887
rect 19674 -14887 19876 -14870
rect 19934 -14870 20894 -14832
rect 19934 -14887 20136 -14870
rect 19674 -14904 19690 -14887
rect 19102 -14920 19690 -14904
rect 20120 -14904 20136 -14887
rect 20692 -14887 20894 -14870
rect 20952 -14870 21912 -14832
rect 20952 -14887 21154 -14870
rect 20692 -14904 20708 -14887
rect 20120 -14920 20708 -14904
rect 21138 -14904 21154 -14887
rect 21710 -14887 21912 -14870
rect 21970 -14870 22930 -14832
rect 21970 -14887 22172 -14870
rect 21710 -14904 21726 -14887
rect 21138 -14920 21726 -14904
rect 22156 -14904 22172 -14887
rect 22728 -14887 22930 -14870
rect 22728 -14904 22744 -14887
rect 22156 -14920 22744 -14904
rect -994 -14966 -34 -14928
rect 2814 -15392 3402 -15376
rect 2814 -15409 2830 -15392
rect 2628 -15426 2830 -15409
rect 3386 -15409 3402 -15392
rect 3832 -15392 4420 -15376
rect 3832 -15409 3848 -15392
rect 3386 -15426 3588 -15409
rect 2628 -15464 3588 -15426
rect 3646 -15426 3848 -15409
rect 4404 -15409 4420 -15392
rect 4850 -15392 5438 -15376
rect 4850 -15409 4866 -15392
rect 4404 -15426 4606 -15409
rect 3646 -15464 4606 -15426
rect 4664 -15426 4866 -15409
rect 5422 -15409 5438 -15392
rect 5868 -15392 6456 -15376
rect 5868 -15409 5884 -15392
rect 5422 -15426 5624 -15409
rect 4664 -15464 5624 -15426
rect 5682 -15426 5884 -15409
rect 6440 -15409 6456 -15392
rect 6886 -15392 7474 -15376
rect 6886 -15409 6902 -15392
rect 6440 -15426 6642 -15409
rect 5682 -15464 6642 -15426
rect 6700 -15426 6902 -15409
rect 7458 -15409 7474 -15392
rect 7904 -15392 8492 -15376
rect 7904 -15409 7920 -15392
rect 7458 -15426 7660 -15409
rect 6700 -15464 7660 -15426
rect 7718 -15426 7920 -15409
rect 8476 -15409 8492 -15392
rect 8922 -15392 9510 -15376
rect 8922 -15409 8938 -15392
rect 8476 -15426 8678 -15409
rect 7718 -15464 8678 -15426
rect 8736 -15426 8938 -15409
rect 9494 -15409 9510 -15392
rect 9940 -15392 10528 -15376
rect 9940 -15409 9956 -15392
rect 9494 -15426 9696 -15409
rect 8736 -15464 9696 -15426
rect 9754 -15426 9956 -15409
rect 10512 -15409 10528 -15392
rect 10958 -15392 11546 -15376
rect 10958 -15409 10974 -15392
rect 10512 -15426 10714 -15409
rect 9754 -15464 10714 -15426
rect 10772 -15426 10974 -15409
rect 11530 -15409 11546 -15392
rect 11976 -15392 12564 -15376
rect 11976 -15409 11992 -15392
rect 11530 -15426 11732 -15409
rect 10772 -15464 11732 -15426
rect 11790 -15426 11992 -15409
rect 12548 -15409 12564 -15392
rect 12994 -15392 13582 -15376
rect 12994 -15409 13010 -15392
rect 12548 -15426 12750 -15409
rect 11790 -15464 12750 -15426
rect 12808 -15426 13010 -15409
rect 13566 -15409 13582 -15392
rect 14012 -15392 14600 -15376
rect 14012 -15409 14028 -15392
rect 13566 -15426 13768 -15409
rect 12808 -15464 13768 -15426
rect 13826 -15426 14028 -15409
rect 14584 -15409 14600 -15392
rect 15030 -15392 15618 -15376
rect 15030 -15409 15046 -15392
rect 14584 -15426 14786 -15409
rect 13826 -15464 14786 -15426
rect 14844 -15426 15046 -15409
rect 15602 -15409 15618 -15392
rect 16048 -15392 16636 -15376
rect 16048 -15409 16064 -15392
rect 15602 -15426 15804 -15409
rect 14844 -15464 15804 -15426
rect 15862 -15426 16064 -15409
rect 16620 -15409 16636 -15392
rect 17066 -15392 17654 -15376
rect 17066 -15409 17082 -15392
rect 16620 -15426 16822 -15409
rect 15862 -15464 16822 -15426
rect 16880 -15426 17082 -15409
rect 17638 -15409 17654 -15392
rect 18084 -15392 18672 -15376
rect 18084 -15409 18100 -15392
rect 17638 -15426 17840 -15409
rect 16880 -15464 17840 -15426
rect 17898 -15426 18100 -15409
rect 18656 -15409 18672 -15392
rect 19102 -15392 19690 -15376
rect 19102 -15409 19118 -15392
rect 18656 -15426 18858 -15409
rect 17898 -15464 18858 -15426
rect 18916 -15426 19118 -15409
rect 19674 -15409 19690 -15392
rect 20120 -15392 20708 -15376
rect 20120 -15409 20136 -15392
rect 19674 -15426 19876 -15409
rect 18916 -15464 19876 -15426
rect 19934 -15426 20136 -15409
rect 20692 -15409 20708 -15392
rect 21138 -15392 21726 -15376
rect 21138 -15409 21154 -15392
rect 20692 -15426 20894 -15409
rect 19934 -15464 20894 -15426
rect 20952 -15426 21154 -15409
rect 21710 -15409 21726 -15392
rect 22156 -15392 22744 -15376
rect 22156 -15409 22172 -15392
rect 21710 -15426 21912 -15409
rect 20952 -15464 21912 -15426
rect 21970 -15426 22172 -15409
rect 22728 -15409 22744 -15392
rect 22728 -15426 22930 -15409
rect 21970 -15464 22930 -15426
rect -9138 -15604 -8178 -15566
rect -9138 -15621 -8936 -15604
rect -8952 -15638 -8936 -15621
rect -8380 -15621 -8178 -15604
rect -8120 -15604 -7160 -15566
rect -8120 -15621 -7918 -15604
rect -8380 -15638 -8364 -15621
rect -8952 -15654 -8364 -15638
rect -7934 -15638 -7918 -15621
rect -7362 -15621 -7160 -15604
rect -7102 -15604 -6142 -15566
rect -7102 -15621 -6900 -15604
rect -7362 -15638 -7346 -15621
rect -7934 -15654 -7346 -15638
rect -8952 -15712 -8364 -15696
rect -8952 -15729 -8936 -15712
rect -9138 -15746 -8936 -15729
rect -8380 -15729 -8364 -15712
rect -6916 -15638 -6900 -15621
rect -6344 -15621 -6142 -15604
rect -6084 -15604 -5124 -15566
rect -6084 -15621 -5882 -15604
rect -6344 -15638 -6328 -15621
rect -6916 -15654 -6328 -15638
rect -7934 -15712 -7346 -15696
rect -7934 -15729 -7918 -15712
rect -8380 -15746 -8178 -15729
rect -9138 -15784 -8178 -15746
rect -8120 -15746 -7918 -15729
rect -7362 -15729 -7346 -15712
rect -5898 -15638 -5882 -15621
rect -5326 -15621 -5124 -15604
rect -5066 -15604 -4106 -15566
rect -5066 -15621 -4864 -15604
rect -5326 -15638 -5310 -15621
rect -5898 -15654 -5310 -15638
rect -6916 -15712 -6328 -15696
rect -6916 -15729 -6900 -15712
rect -7362 -15746 -7160 -15729
rect -8120 -15784 -7160 -15746
rect -7102 -15746 -6900 -15729
rect -6344 -15729 -6328 -15712
rect -4880 -15638 -4864 -15621
rect -4308 -15621 -4106 -15604
rect -4048 -15604 -3088 -15566
rect -4048 -15621 -3846 -15604
rect -4308 -15638 -4292 -15621
rect -4880 -15654 -4292 -15638
rect -5898 -15712 -5310 -15696
rect -5898 -15729 -5882 -15712
rect -6344 -15746 -6142 -15729
rect -7102 -15784 -6142 -15746
rect -6084 -15746 -5882 -15729
rect -5326 -15729 -5310 -15712
rect -3862 -15638 -3846 -15621
rect -3290 -15621 -3088 -15604
rect -3030 -15604 -2070 -15566
rect -3030 -15621 -2828 -15604
rect -3290 -15638 -3274 -15621
rect -3862 -15654 -3274 -15638
rect -4880 -15712 -4292 -15696
rect -4880 -15729 -4864 -15712
rect -5326 -15746 -5124 -15729
rect -6084 -15784 -5124 -15746
rect -5066 -15746 -4864 -15729
rect -4308 -15729 -4292 -15712
rect -2844 -15638 -2828 -15621
rect -2272 -15621 -2070 -15604
rect -2012 -15604 -1052 -15566
rect -2012 -15621 -1810 -15604
rect -2272 -15638 -2256 -15621
rect -2844 -15654 -2256 -15638
rect -3862 -15712 -3274 -15696
rect -3862 -15729 -3846 -15712
rect -4308 -15746 -4106 -15729
rect -5066 -15784 -4106 -15746
rect -4048 -15746 -3846 -15729
rect -3290 -15729 -3274 -15712
rect -1826 -15638 -1810 -15621
rect -1254 -15621 -1052 -15604
rect -994 -15604 -34 -15566
rect -994 -15621 -792 -15604
rect -1254 -15638 -1238 -15621
rect -1826 -15654 -1238 -15638
rect -2844 -15712 -2256 -15696
rect -2844 -15729 -2828 -15712
rect -3290 -15746 -3088 -15729
rect -4048 -15784 -3088 -15746
rect -3030 -15746 -2828 -15729
rect -2272 -15729 -2256 -15712
rect -808 -15638 -792 -15621
rect -236 -15621 -34 -15604
rect -236 -15638 -220 -15621
rect -808 -15654 -220 -15638
rect -1826 -15712 -1238 -15696
rect -1826 -15729 -1810 -15712
rect -2272 -15746 -2070 -15729
rect -3030 -15784 -2070 -15746
rect -2012 -15746 -1810 -15729
rect -1254 -15729 -1238 -15712
rect -808 -15712 -220 -15696
rect -808 -15729 -792 -15712
rect -1254 -15746 -1052 -15729
rect -2012 -15784 -1052 -15746
rect -994 -15746 -792 -15729
rect -236 -15729 -220 -15712
rect -236 -15746 -34 -15729
rect -994 -15784 -34 -15746
rect 2628 -16102 3588 -16064
rect 2628 -16119 2830 -16102
rect 2814 -16136 2830 -16119
rect 3386 -16119 3588 -16102
rect 3646 -16102 4606 -16064
rect 3646 -16119 3848 -16102
rect 3386 -16136 3402 -16119
rect 2814 -16152 3402 -16136
rect 3832 -16136 3848 -16119
rect 4404 -16119 4606 -16102
rect 4664 -16102 5624 -16064
rect 4664 -16119 4866 -16102
rect 4404 -16136 4420 -16119
rect 3832 -16152 4420 -16136
rect 4850 -16136 4866 -16119
rect 5422 -16119 5624 -16102
rect 5682 -16102 6642 -16064
rect 5682 -16119 5884 -16102
rect 5422 -16136 5438 -16119
rect 4850 -16152 5438 -16136
rect 5868 -16136 5884 -16119
rect 6440 -16119 6642 -16102
rect 6700 -16102 7660 -16064
rect 6700 -16119 6902 -16102
rect 6440 -16136 6456 -16119
rect 5868 -16152 6456 -16136
rect 6886 -16136 6902 -16119
rect 7458 -16119 7660 -16102
rect 7718 -16102 8678 -16064
rect 7718 -16119 7920 -16102
rect 7458 -16136 7474 -16119
rect 6886 -16152 7474 -16136
rect 7904 -16136 7920 -16119
rect 8476 -16119 8678 -16102
rect 8736 -16102 9696 -16064
rect 8736 -16119 8938 -16102
rect 8476 -16136 8492 -16119
rect 7904 -16152 8492 -16136
rect 8922 -16136 8938 -16119
rect 9494 -16119 9696 -16102
rect 9754 -16102 10714 -16064
rect 9754 -16119 9956 -16102
rect 9494 -16136 9510 -16119
rect 8922 -16152 9510 -16136
rect 9940 -16136 9956 -16119
rect 10512 -16119 10714 -16102
rect 10772 -16102 11732 -16064
rect 10772 -16119 10974 -16102
rect 10512 -16136 10528 -16119
rect 9940 -16152 10528 -16136
rect 10958 -16136 10974 -16119
rect 11530 -16119 11732 -16102
rect 11790 -16102 12750 -16064
rect 11790 -16119 11992 -16102
rect 11530 -16136 11546 -16119
rect 10958 -16152 11546 -16136
rect 11976 -16136 11992 -16119
rect 12548 -16119 12750 -16102
rect 12808 -16102 13768 -16064
rect 12808 -16119 13010 -16102
rect 12548 -16136 12564 -16119
rect 11976 -16152 12564 -16136
rect 12994 -16136 13010 -16119
rect 13566 -16119 13768 -16102
rect 13826 -16102 14786 -16064
rect 13826 -16119 14028 -16102
rect 13566 -16136 13582 -16119
rect 12994 -16152 13582 -16136
rect 14012 -16136 14028 -16119
rect 14584 -16119 14786 -16102
rect 14844 -16102 15804 -16064
rect 14844 -16119 15046 -16102
rect 14584 -16136 14600 -16119
rect 14012 -16152 14600 -16136
rect 15030 -16136 15046 -16119
rect 15602 -16119 15804 -16102
rect 15862 -16102 16822 -16064
rect 15862 -16119 16064 -16102
rect 15602 -16136 15618 -16119
rect 15030 -16152 15618 -16136
rect 16048 -16136 16064 -16119
rect 16620 -16119 16822 -16102
rect 16880 -16102 17840 -16064
rect 16880 -16119 17082 -16102
rect 16620 -16136 16636 -16119
rect 16048 -16152 16636 -16136
rect 17066 -16136 17082 -16119
rect 17638 -16119 17840 -16102
rect 17898 -16102 18858 -16064
rect 17898 -16119 18100 -16102
rect 17638 -16136 17654 -16119
rect 17066 -16152 17654 -16136
rect 18084 -16136 18100 -16119
rect 18656 -16119 18858 -16102
rect 18916 -16102 19876 -16064
rect 18916 -16119 19118 -16102
rect 18656 -16136 18672 -16119
rect 18084 -16152 18672 -16136
rect 19102 -16136 19118 -16119
rect 19674 -16119 19876 -16102
rect 19934 -16102 20894 -16064
rect 19934 -16119 20136 -16102
rect 19674 -16136 19690 -16119
rect 19102 -16152 19690 -16136
rect 20120 -16136 20136 -16119
rect 20692 -16119 20894 -16102
rect 20952 -16102 21912 -16064
rect 20952 -16119 21154 -16102
rect 20692 -16136 20708 -16119
rect 20120 -16152 20708 -16136
rect 21138 -16136 21154 -16119
rect 21710 -16119 21912 -16102
rect 21970 -16102 22930 -16064
rect 21970 -16119 22172 -16102
rect 21710 -16136 21726 -16119
rect 21138 -16152 21726 -16136
rect 22156 -16136 22172 -16119
rect 22728 -16119 22930 -16102
rect 22728 -16136 22744 -16119
rect 22156 -16152 22744 -16136
rect -9138 -16422 -8178 -16384
rect -9138 -16439 -8936 -16422
rect -8952 -16456 -8936 -16439
rect -8380 -16439 -8178 -16422
rect -8120 -16422 -7160 -16384
rect -8120 -16439 -7918 -16422
rect -8380 -16456 -8364 -16439
rect -8952 -16472 -8364 -16456
rect -7934 -16456 -7918 -16439
rect -7362 -16439 -7160 -16422
rect -7102 -16422 -6142 -16384
rect -7102 -16439 -6900 -16422
rect -7362 -16456 -7346 -16439
rect -7934 -16472 -7346 -16456
rect -8952 -16530 -8364 -16514
rect -8952 -16547 -8936 -16530
rect -9138 -16564 -8936 -16547
rect -8380 -16547 -8364 -16530
rect -6916 -16456 -6900 -16439
rect -6344 -16439 -6142 -16422
rect -6084 -16422 -5124 -16384
rect -6084 -16439 -5882 -16422
rect -6344 -16456 -6328 -16439
rect -6916 -16472 -6328 -16456
rect -7934 -16530 -7346 -16514
rect -7934 -16547 -7918 -16530
rect -8380 -16564 -8178 -16547
rect -9138 -16602 -8178 -16564
rect -8120 -16564 -7918 -16547
rect -7362 -16547 -7346 -16530
rect -5898 -16456 -5882 -16439
rect -5326 -16439 -5124 -16422
rect -5066 -16422 -4106 -16384
rect -5066 -16439 -4864 -16422
rect -5326 -16456 -5310 -16439
rect -5898 -16472 -5310 -16456
rect -6916 -16530 -6328 -16514
rect -6916 -16547 -6900 -16530
rect -7362 -16564 -7160 -16547
rect -8120 -16602 -7160 -16564
rect -7102 -16564 -6900 -16547
rect -6344 -16547 -6328 -16530
rect -4880 -16456 -4864 -16439
rect -4308 -16439 -4106 -16422
rect -4048 -16422 -3088 -16384
rect -4048 -16439 -3846 -16422
rect -4308 -16456 -4292 -16439
rect -4880 -16472 -4292 -16456
rect -5898 -16530 -5310 -16514
rect -5898 -16547 -5882 -16530
rect -6344 -16564 -6142 -16547
rect -7102 -16602 -6142 -16564
rect -6084 -16564 -5882 -16547
rect -5326 -16547 -5310 -16530
rect -3862 -16456 -3846 -16439
rect -3290 -16439 -3088 -16422
rect -3030 -16422 -2070 -16384
rect -3030 -16439 -2828 -16422
rect -3290 -16456 -3274 -16439
rect -3862 -16472 -3274 -16456
rect -4880 -16530 -4292 -16514
rect -4880 -16547 -4864 -16530
rect -5326 -16564 -5124 -16547
rect -6084 -16602 -5124 -16564
rect -5066 -16564 -4864 -16547
rect -4308 -16547 -4292 -16530
rect -2844 -16456 -2828 -16439
rect -2272 -16439 -2070 -16422
rect -2012 -16422 -1052 -16384
rect -2012 -16439 -1810 -16422
rect -2272 -16456 -2256 -16439
rect -2844 -16472 -2256 -16456
rect -3862 -16530 -3274 -16514
rect -3862 -16547 -3846 -16530
rect -4308 -16564 -4106 -16547
rect -5066 -16602 -4106 -16564
rect -4048 -16564 -3846 -16547
rect -3290 -16547 -3274 -16530
rect -1826 -16456 -1810 -16439
rect -1254 -16439 -1052 -16422
rect -994 -16422 -34 -16384
rect -994 -16439 -792 -16422
rect -1254 -16456 -1238 -16439
rect -1826 -16472 -1238 -16456
rect -2844 -16530 -2256 -16514
rect -2844 -16547 -2828 -16530
rect -3290 -16564 -3088 -16547
rect -4048 -16602 -3088 -16564
rect -3030 -16564 -2828 -16547
rect -2272 -16547 -2256 -16530
rect -808 -16456 -792 -16439
rect -236 -16439 -34 -16422
rect -236 -16456 -220 -16439
rect -808 -16472 -220 -16456
rect -1826 -16530 -1238 -16514
rect -1826 -16547 -1810 -16530
rect -2272 -16564 -2070 -16547
rect -3030 -16602 -2070 -16564
rect -2012 -16564 -1810 -16547
rect -1254 -16547 -1238 -16530
rect -808 -16530 -220 -16514
rect -808 -16547 -792 -16530
rect -1254 -16564 -1052 -16547
rect -2012 -16602 -1052 -16564
rect -994 -16564 -792 -16547
rect -236 -16547 -220 -16530
rect -236 -16564 -34 -16547
rect -994 -16602 -34 -16564
rect 2812 -16626 3400 -16610
rect 2812 -16643 2828 -16626
rect 2626 -16660 2828 -16643
rect 3384 -16643 3400 -16626
rect 3830 -16626 4418 -16610
rect 3830 -16643 3846 -16626
rect 3384 -16660 3586 -16643
rect 2626 -16698 3586 -16660
rect 3644 -16660 3846 -16643
rect 4402 -16643 4418 -16626
rect 4848 -16626 5436 -16610
rect 4848 -16643 4864 -16626
rect 4402 -16660 4604 -16643
rect 3644 -16698 4604 -16660
rect 4662 -16660 4864 -16643
rect 5420 -16643 5436 -16626
rect 5866 -16626 6454 -16610
rect 5866 -16643 5882 -16626
rect 5420 -16660 5622 -16643
rect 4662 -16698 5622 -16660
rect 5680 -16660 5882 -16643
rect 6438 -16643 6454 -16626
rect 6884 -16626 7472 -16610
rect 6884 -16643 6900 -16626
rect 6438 -16660 6640 -16643
rect 5680 -16698 6640 -16660
rect 6698 -16660 6900 -16643
rect 7456 -16643 7472 -16626
rect 7902 -16626 8490 -16610
rect 7902 -16643 7918 -16626
rect 7456 -16660 7658 -16643
rect 6698 -16698 7658 -16660
rect 7716 -16660 7918 -16643
rect 8474 -16643 8490 -16626
rect 8920 -16626 9508 -16610
rect 8920 -16643 8936 -16626
rect 8474 -16660 8676 -16643
rect 7716 -16698 8676 -16660
rect 8734 -16660 8936 -16643
rect 9492 -16643 9508 -16626
rect 9938 -16626 10526 -16610
rect 9938 -16643 9954 -16626
rect 9492 -16660 9694 -16643
rect 8734 -16698 9694 -16660
rect 9752 -16660 9954 -16643
rect 10510 -16643 10526 -16626
rect 10956 -16626 11544 -16610
rect 10956 -16643 10972 -16626
rect 10510 -16660 10712 -16643
rect 9752 -16698 10712 -16660
rect 10770 -16660 10972 -16643
rect 11528 -16643 11544 -16626
rect 11974 -16626 12562 -16610
rect 11974 -16643 11990 -16626
rect 11528 -16660 11730 -16643
rect 10770 -16698 11730 -16660
rect 11788 -16660 11990 -16643
rect 12546 -16643 12562 -16626
rect 12992 -16626 13580 -16610
rect 12992 -16643 13008 -16626
rect 12546 -16660 12748 -16643
rect 11788 -16698 12748 -16660
rect 12806 -16660 13008 -16643
rect 13564 -16643 13580 -16626
rect 14010 -16626 14598 -16610
rect 14010 -16643 14026 -16626
rect 13564 -16660 13766 -16643
rect 12806 -16698 13766 -16660
rect 13824 -16660 14026 -16643
rect 14582 -16643 14598 -16626
rect 15028 -16626 15616 -16610
rect 15028 -16643 15044 -16626
rect 14582 -16660 14784 -16643
rect 13824 -16698 14784 -16660
rect 14842 -16660 15044 -16643
rect 15600 -16643 15616 -16626
rect 16046 -16626 16634 -16610
rect 16046 -16643 16062 -16626
rect 15600 -16660 15802 -16643
rect 14842 -16698 15802 -16660
rect 15860 -16660 16062 -16643
rect 16618 -16643 16634 -16626
rect 17064 -16626 17652 -16610
rect 17064 -16643 17080 -16626
rect 16618 -16660 16820 -16643
rect 15860 -16698 16820 -16660
rect 16878 -16660 17080 -16643
rect 17636 -16643 17652 -16626
rect 18082 -16626 18670 -16610
rect 18082 -16643 18098 -16626
rect 17636 -16660 17838 -16643
rect 16878 -16698 17838 -16660
rect 17896 -16660 18098 -16643
rect 18654 -16643 18670 -16626
rect 19100 -16626 19688 -16610
rect 19100 -16643 19116 -16626
rect 18654 -16660 18856 -16643
rect 17896 -16698 18856 -16660
rect 18914 -16660 19116 -16643
rect 19672 -16643 19688 -16626
rect 20118 -16626 20706 -16610
rect 20118 -16643 20134 -16626
rect 19672 -16660 19874 -16643
rect 18914 -16698 19874 -16660
rect 19932 -16660 20134 -16643
rect 20690 -16643 20706 -16626
rect 21136 -16626 21724 -16610
rect 21136 -16643 21152 -16626
rect 20690 -16660 20892 -16643
rect 19932 -16698 20892 -16660
rect 20950 -16660 21152 -16643
rect 21708 -16643 21724 -16626
rect 22154 -16626 22742 -16610
rect 22154 -16643 22170 -16626
rect 21708 -16660 21910 -16643
rect 20950 -16698 21910 -16660
rect 21968 -16660 22170 -16643
rect 22726 -16643 22742 -16626
rect 22726 -16660 22928 -16643
rect 21968 -16698 22928 -16660
rect -9138 -17240 -8178 -17202
rect -9138 -17257 -8936 -17240
rect -8952 -17274 -8936 -17257
rect -8380 -17257 -8178 -17240
rect -8120 -17240 -7160 -17202
rect -8120 -17257 -7918 -17240
rect -8380 -17274 -8364 -17257
rect -8952 -17290 -8364 -17274
rect -7934 -17274 -7918 -17257
rect -7362 -17257 -7160 -17240
rect -7102 -17240 -6142 -17202
rect -7102 -17257 -6900 -17240
rect -7362 -17274 -7346 -17257
rect -7934 -17290 -7346 -17274
rect -8952 -17348 -8364 -17332
rect -8952 -17365 -8936 -17348
rect -9138 -17382 -8936 -17365
rect -8380 -17365 -8364 -17348
rect -6916 -17274 -6900 -17257
rect -6344 -17257 -6142 -17240
rect -6084 -17240 -5124 -17202
rect -6084 -17257 -5882 -17240
rect -6344 -17274 -6328 -17257
rect -6916 -17290 -6328 -17274
rect -7934 -17348 -7346 -17332
rect -7934 -17365 -7918 -17348
rect -8380 -17382 -8178 -17365
rect -9138 -17420 -8178 -17382
rect -8120 -17382 -7918 -17365
rect -7362 -17365 -7346 -17348
rect -5898 -17274 -5882 -17257
rect -5326 -17257 -5124 -17240
rect -5066 -17240 -4106 -17202
rect -5066 -17257 -4864 -17240
rect -5326 -17274 -5310 -17257
rect -5898 -17290 -5310 -17274
rect -6916 -17348 -6328 -17332
rect -6916 -17365 -6900 -17348
rect -7362 -17382 -7160 -17365
rect -8120 -17420 -7160 -17382
rect -7102 -17382 -6900 -17365
rect -6344 -17365 -6328 -17348
rect -4880 -17274 -4864 -17257
rect -4308 -17257 -4106 -17240
rect -4048 -17240 -3088 -17202
rect -4048 -17257 -3846 -17240
rect -4308 -17274 -4292 -17257
rect -4880 -17290 -4292 -17274
rect -5898 -17348 -5310 -17332
rect -5898 -17365 -5882 -17348
rect -6344 -17382 -6142 -17365
rect -7102 -17420 -6142 -17382
rect -6084 -17382 -5882 -17365
rect -5326 -17365 -5310 -17348
rect -3862 -17274 -3846 -17257
rect -3290 -17257 -3088 -17240
rect -3030 -17240 -2070 -17202
rect -3030 -17257 -2828 -17240
rect -3290 -17274 -3274 -17257
rect -3862 -17290 -3274 -17274
rect -4880 -17348 -4292 -17332
rect -4880 -17365 -4864 -17348
rect -5326 -17382 -5124 -17365
rect -6084 -17420 -5124 -17382
rect -5066 -17382 -4864 -17365
rect -4308 -17365 -4292 -17348
rect -2844 -17274 -2828 -17257
rect -2272 -17257 -2070 -17240
rect -2012 -17240 -1052 -17202
rect -2012 -17257 -1810 -17240
rect -2272 -17274 -2256 -17257
rect -2844 -17290 -2256 -17274
rect -3862 -17348 -3274 -17332
rect -3862 -17365 -3846 -17348
rect -4308 -17382 -4106 -17365
rect -5066 -17420 -4106 -17382
rect -4048 -17382 -3846 -17365
rect -3290 -17365 -3274 -17348
rect -1826 -17274 -1810 -17257
rect -1254 -17257 -1052 -17240
rect -994 -17240 -34 -17202
rect -994 -17257 -792 -17240
rect -1254 -17274 -1238 -17257
rect -1826 -17290 -1238 -17274
rect -2844 -17348 -2256 -17332
rect -2844 -17365 -2828 -17348
rect -3290 -17382 -3088 -17365
rect -4048 -17420 -3088 -17382
rect -3030 -17382 -2828 -17365
rect -2272 -17365 -2256 -17348
rect -808 -17274 -792 -17257
rect -236 -17257 -34 -17240
rect -236 -17274 -220 -17257
rect -808 -17290 -220 -17274
rect -1826 -17348 -1238 -17332
rect -1826 -17365 -1810 -17348
rect -2272 -17382 -2070 -17365
rect -3030 -17420 -2070 -17382
rect -2012 -17382 -1810 -17365
rect -1254 -17365 -1238 -17348
rect -808 -17348 -220 -17332
rect -808 -17365 -792 -17348
rect -1254 -17382 -1052 -17365
rect -2012 -17420 -1052 -17382
rect -994 -17382 -792 -17365
rect -236 -17365 -220 -17348
rect 2626 -17336 3586 -17298
rect 2626 -17353 2828 -17336
rect -236 -17382 -34 -17365
rect -994 -17420 -34 -17382
rect 2812 -17370 2828 -17353
rect 3384 -17353 3586 -17336
rect 3644 -17336 4604 -17298
rect 3644 -17353 3846 -17336
rect 3384 -17370 3400 -17353
rect 2812 -17386 3400 -17370
rect 3830 -17370 3846 -17353
rect 4402 -17353 4604 -17336
rect 4662 -17336 5622 -17298
rect 4662 -17353 4864 -17336
rect 4402 -17370 4418 -17353
rect 3830 -17386 4418 -17370
rect 4848 -17370 4864 -17353
rect 5420 -17353 5622 -17336
rect 5680 -17336 6640 -17298
rect 5680 -17353 5882 -17336
rect 5420 -17370 5436 -17353
rect 4848 -17386 5436 -17370
rect 5866 -17370 5882 -17353
rect 6438 -17353 6640 -17336
rect 6698 -17336 7658 -17298
rect 6698 -17353 6900 -17336
rect 6438 -17370 6454 -17353
rect 5866 -17386 6454 -17370
rect 6884 -17370 6900 -17353
rect 7456 -17353 7658 -17336
rect 7716 -17336 8676 -17298
rect 7716 -17353 7918 -17336
rect 7456 -17370 7472 -17353
rect 6884 -17386 7472 -17370
rect 7902 -17370 7918 -17353
rect 8474 -17353 8676 -17336
rect 8734 -17336 9694 -17298
rect 8734 -17353 8936 -17336
rect 8474 -17370 8490 -17353
rect 7902 -17386 8490 -17370
rect 8920 -17370 8936 -17353
rect 9492 -17353 9694 -17336
rect 9752 -17336 10712 -17298
rect 9752 -17353 9954 -17336
rect 9492 -17370 9508 -17353
rect 8920 -17386 9508 -17370
rect 9938 -17370 9954 -17353
rect 10510 -17353 10712 -17336
rect 10770 -17336 11730 -17298
rect 10770 -17353 10972 -17336
rect 10510 -17370 10526 -17353
rect 9938 -17386 10526 -17370
rect 10956 -17370 10972 -17353
rect 11528 -17353 11730 -17336
rect 11788 -17336 12748 -17298
rect 11788 -17353 11990 -17336
rect 11528 -17370 11544 -17353
rect 10956 -17386 11544 -17370
rect 11974 -17370 11990 -17353
rect 12546 -17353 12748 -17336
rect 12806 -17336 13766 -17298
rect 12806 -17353 13008 -17336
rect 12546 -17370 12562 -17353
rect 11974 -17386 12562 -17370
rect 12992 -17370 13008 -17353
rect 13564 -17353 13766 -17336
rect 13824 -17336 14784 -17298
rect 13824 -17353 14026 -17336
rect 13564 -17370 13580 -17353
rect 12992 -17386 13580 -17370
rect 14010 -17370 14026 -17353
rect 14582 -17353 14784 -17336
rect 14842 -17336 15802 -17298
rect 14842 -17353 15044 -17336
rect 14582 -17370 14598 -17353
rect 14010 -17386 14598 -17370
rect 15028 -17370 15044 -17353
rect 15600 -17353 15802 -17336
rect 15860 -17336 16820 -17298
rect 15860 -17353 16062 -17336
rect 15600 -17370 15616 -17353
rect 15028 -17386 15616 -17370
rect 16046 -17370 16062 -17353
rect 16618 -17353 16820 -17336
rect 16878 -17336 17838 -17298
rect 16878 -17353 17080 -17336
rect 16618 -17370 16634 -17353
rect 16046 -17386 16634 -17370
rect 17064 -17370 17080 -17353
rect 17636 -17353 17838 -17336
rect 17896 -17336 18856 -17298
rect 17896 -17353 18098 -17336
rect 17636 -17370 17652 -17353
rect 17064 -17386 17652 -17370
rect 18082 -17370 18098 -17353
rect 18654 -17353 18856 -17336
rect 18914 -17336 19874 -17298
rect 18914 -17353 19116 -17336
rect 18654 -17370 18670 -17353
rect 18082 -17386 18670 -17370
rect 19100 -17370 19116 -17353
rect 19672 -17353 19874 -17336
rect 19932 -17336 20892 -17298
rect 19932 -17353 20134 -17336
rect 19672 -17370 19688 -17353
rect 19100 -17386 19688 -17370
rect 20118 -17370 20134 -17353
rect 20690 -17353 20892 -17336
rect 20950 -17336 21910 -17298
rect 20950 -17353 21152 -17336
rect 20690 -17370 20706 -17353
rect 20118 -17386 20706 -17370
rect 21136 -17370 21152 -17353
rect 21708 -17353 21910 -17336
rect 21968 -17336 22928 -17298
rect 21968 -17353 22170 -17336
rect 21708 -17370 21724 -17353
rect 21136 -17386 21724 -17370
rect 22154 -17370 22170 -17353
rect 22726 -17353 22928 -17336
rect 22726 -17370 22742 -17353
rect 22154 -17386 22742 -17370
rect 2812 -17860 3400 -17844
rect 2812 -17877 2828 -17860
rect 2626 -17894 2828 -17877
rect 3384 -17877 3400 -17860
rect 3830 -17860 4418 -17844
rect 3830 -17877 3846 -17860
rect 3384 -17894 3586 -17877
rect 2626 -17932 3586 -17894
rect 3644 -17894 3846 -17877
rect 4402 -17877 4418 -17860
rect 4848 -17860 5436 -17844
rect 4848 -17877 4864 -17860
rect 4402 -17894 4604 -17877
rect 3644 -17932 4604 -17894
rect 4662 -17894 4864 -17877
rect 5420 -17877 5436 -17860
rect 5866 -17860 6454 -17844
rect 5866 -17877 5882 -17860
rect 5420 -17894 5622 -17877
rect 4662 -17932 5622 -17894
rect 5680 -17894 5882 -17877
rect 6438 -17877 6454 -17860
rect 6884 -17860 7472 -17844
rect 6884 -17877 6900 -17860
rect 6438 -17894 6640 -17877
rect 5680 -17932 6640 -17894
rect 6698 -17894 6900 -17877
rect 7456 -17877 7472 -17860
rect 7902 -17860 8490 -17844
rect 7902 -17877 7918 -17860
rect 7456 -17894 7658 -17877
rect 6698 -17932 7658 -17894
rect 7716 -17894 7918 -17877
rect 8474 -17877 8490 -17860
rect 8920 -17860 9508 -17844
rect 8920 -17877 8936 -17860
rect 8474 -17894 8676 -17877
rect 7716 -17932 8676 -17894
rect 8734 -17894 8936 -17877
rect 9492 -17877 9508 -17860
rect 9938 -17860 10526 -17844
rect 9938 -17877 9954 -17860
rect 9492 -17894 9694 -17877
rect 8734 -17932 9694 -17894
rect 9752 -17894 9954 -17877
rect 10510 -17877 10526 -17860
rect 10956 -17860 11544 -17844
rect 10956 -17877 10972 -17860
rect 10510 -17894 10712 -17877
rect 9752 -17932 10712 -17894
rect 10770 -17894 10972 -17877
rect 11528 -17877 11544 -17860
rect 11974 -17860 12562 -17844
rect 11974 -17877 11990 -17860
rect 11528 -17894 11730 -17877
rect 10770 -17932 11730 -17894
rect 11788 -17894 11990 -17877
rect 12546 -17877 12562 -17860
rect 12992 -17860 13580 -17844
rect 12992 -17877 13008 -17860
rect 12546 -17894 12748 -17877
rect 11788 -17932 12748 -17894
rect 12806 -17894 13008 -17877
rect 13564 -17877 13580 -17860
rect 14010 -17860 14598 -17844
rect 14010 -17877 14026 -17860
rect 13564 -17894 13766 -17877
rect 12806 -17932 13766 -17894
rect 13824 -17894 14026 -17877
rect 14582 -17877 14598 -17860
rect 15028 -17860 15616 -17844
rect 15028 -17877 15044 -17860
rect 14582 -17894 14784 -17877
rect 13824 -17932 14784 -17894
rect 14842 -17894 15044 -17877
rect 15600 -17877 15616 -17860
rect 16046 -17860 16634 -17844
rect 16046 -17877 16062 -17860
rect 15600 -17894 15802 -17877
rect 14842 -17932 15802 -17894
rect 15860 -17894 16062 -17877
rect 16618 -17877 16634 -17860
rect 17064 -17860 17652 -17844
rect 17064 -17877 17080 -17860
rect 16618 -17894 16820 -17877
rect 15860 -17932 16820 -17894
rect 16878 -17894 17080 -17877
rect 17636 -17877 17652 -17860
rect 18082 -17860 18670 -17844
rect 18082 -17877 18098 -17860
rect 17636 -17894 17838 -17877
rect 16878 -17932 17838 -17894
rect 17896 -17894 18098 -17877
rect 18654 -17877 18670 -17860
rect 19100 -17860 19688 -17844
rect 19100 -17877 19116 -17860
rect 18654 -17894 18856 -17877
rect 17896 -17932 18856 -17894
rect 18914 -17894 19116 -17877
rect 19672 -17877 19688 -17860
rect 20118 -17860 20706 -17844
rect 20118 -17877 20134 -17860
rect 19672 -17894 19874 -17877
rect 18914 -17932 19874 -17894
rect 19932 -17894 20134 -17877
rect 20690 -17877 20706 -17860
rect 21136 -17860 21724 -17844
rect 21136 -17877 21152 -17860
rect 20690 -17894 20892 -17877
rect 19932 -17932 20892 -17894
rect 20950 -17894 21152 -17877
rect 21708 -17877 21724 -17860
rect 22154 -17860 22742 -17844
rect 22154 -17877 22170 -17860
rect 21708 -17894 21910 -17877
rect 20950 -17932 21910 -17894
rect 21968 -17894 22170 -17877
rect 22726 -17877 22742 -17860
rect 22726 -17894 22928 -17877
rect 21968 -17932 22928 -17894
rect -9138 -18058 -8178 -18020
rect -9138 -18075 -8936 -18058
rect -8952 -18092 -8936 -18075
rect -8380 -18075 -8178 -18058
rect -8120 -18058 -7160 -18020
rect -8120 -18075 -7918 -18058
rect -8380 -18092 -8364 -18075
rect -8952 -18108 -8364 -18092
rect -7934 -18092 -7918 -18075
rect -7362 -18075 -7160 -18058
rect -7102 -18058 -6142 -18020
rect -7102 -18075 -6900 -18058
rect -7362 -18092 -7346 -18075
rect -7934 -18108 -7346 -18092
rect -8952 -18166 -8364 -18150
rect -8952 -18183 -8936 -18166
rect -9138 -18200 -8936 -18183
rect -8380 -18183 -8364 -18166
rect -6916 -18092 -6900 -18075
rect -6344 -18075 -6142 -18058
rect -6084 -18058 -5124 -18020
rect -6084 -18075 -5882 -18058
rect -6344 -18092 -6328 -18075
rect -6916 -18108 -6328 -18092
rect -7934 -18166 -7346 -18150
rect -7934 -18183 -7918 -18166
rect -8380 -18200 -8178 -18183
rect -9138 -18238 -8178 -18200
rect -8120 -18200 -7918 -18183
rect -7362 -18183 -7346 -18166
rect -5898 -18092 -5882 -18075
rect -5326 -18075 -5124 -18058
rect -5066 -18058 -4106 -18020
rect -5066 -18075 -4864 -18058
rect -5326 -18092 -5310 -18075
rect -5898 -18108 -5310 -18092
rect -6916 -18166 -6328 -18150
rect -6916 -18183 -6900 -18166
rect -7362 -18200 -7160 -18183
rect -8120 -18238 -7160 -18200
rect -7102 -18200 -6900 -18183
rect -6344 -18183 -6328 -18166
rect -4880 -18092 -4864 -18075
rect -4308 -18075 -4106 -18058
rect -4048 -18058 -3088 -18020
rect -4048 -18075 -3846 -18058
rect -4308 -18092 -4292 -18075
rect -4880 -18108 -4292 -18092
rect -5898 -18166 -5310 -18150
rect -5898 -18183 -5882 -18166
rect -6344 -18200 -6142 -18183
rect -7102 -18238 -6142 -18200
rect -6084 -18200 -5882 -18183
rect -5326 -18183 -5310 -18166
rect -3862 -18092 -3846 -18075
rect -3290 -18075 -3088 -18058
rect -3030 -18058 -2070 -18020
rect -3030 -18075 -2828 -18058
rect -3290 -18092 -3274 -18075
rect -3862 -18108 -3274 -18092
rect -4880 -18166 -4292 -18150
rect -4880 -18183 -4864 -18166
rect -5326 -18200 -5124 -18183
rect -6084 -18238 -5124 -18200
rect -5066 -18200 -4864 -18183
rect -4308 -18183 -4292 -18166
rect -2844 -18092 -2828 -18075
rect -2272 -18075 -2070 -18058
rect -2012 -18058 -1052 -18020
rect -2012 -18075 -1810 -18058
rect -2272 -18092 -2256 -18075
rect -2844 -18108 -2256 -18092
rect -3862 -18166 -3274 -18150
rect -3862 -18183 -3846 -18166
rect -4308 -18200 -4106 -18183
rect -5066 -18238 -4106 -18200
rect -4048 -18200 -3846 -18183
rect -3290 -18183 -3274 -18166
rect -1826 -18092 -1810 -18075
rect -1254 -18075 -1052 -18058
rect -994 -18058 -34 -18020
rect -994 -18075 -792 -18058
rect -1254 -18092 -1238 -18075
rect -1826 -18108 -1238 -18092
rect -2844 -18166 -2256 -18150
rect -2844 -18183 -2828 -18166
rect -3290 -18200 -3088 -18183
rect -4048 -18238 -3088 -18200
rect -3030 -18200 -2828 -18183
rect -2272 -18183 -2256 -18166
rect -808 -18092 -792 -18075
rect -236 -18075 -34 -18058
rect -236 -18092 -220 -18075
rect -808 -18108 -220 -18092
rect -1826 -18166 -1238 -18150
rect -1826 -18183 -1810 -18166
rect -2272 -18200 -2070 -18183
rect -3030 -18238 -2070 -18200
rect -2012 -18200 -1810 -18183
rect -1254 -18183 -1238 -18166
rect -808 -18166 -220 -18150
rect -808 -18183 -792 -18166
rect -1254 -18200 -1052 -18183
rect -2012 -18238 -1052 -18200
rect -994 -18200 -792 -18183
rect -236 -18183 -220 -18166
rect -236 -18200 -34 -18183
rect -994 -18238 -34 -18200
rect 2626 -18570 3586 -18532
rect 2626 -18587 2828 -18570
rect 2812 -18604 2828 -18587
rect 3384 -18587 3586 -18570
rect 3644 -18570 4604 -18532
rect 3644 -18587 3846 -18570
rect 3384 -18604 3400 -18587
rect 2812 -18620 3400 -18604
rect 3830 -18604 3846 -18587
rect 4402 -18587 4604 -18570
rect 4662 -18570 5622 -18532
rect 4662 -18587 4864 -18570
rect 4402 -18604 4418 -18587
rect 3830 -18620 4418 -18604
rect 4848 -18604 4864 -18587
rect 5420 -18587 5622 -18570
rect 5680 -18570 6640 -18532
rect 5680 -18587 5882 -18570
rect 5420 -18604 5436 -18587
rect 4848 -18620 5436 -18604
rect 5866 -18604 5882 -18587
rect 6438 -18587 6640 -18570
rect 6698 -18570 7658 -18532
rect 6698 -18587 6900 -18570
rect 6438 -18604 6454 -18587
rect 5866 -18620 6454 -18604
rect 6884 -18604 6900 -18587
rect 7456 -18587 7658 -18570
rect 7716 -18570 8676 -18532
rect 7716 -18587 7918 -18570
rect 7456 -18604 7472 -18587
rect 6884 -18620 7472 -18604
rect 7902 -18604 7918 -18587
rect 8474 -18587 8676 -18570
rect 8734 -18570 9694 -18532
rect 8734 -18587 8936 -18570
rect 8474 -18604 8490 -18587
rect 7902 -18620 8490 -18604
rect 8920 -18604 8936 -18587
rect 9492 -18587 9694 -18570
rect 9752 -18570 10712 -18532
rect 9752 -18587 9954 -18570
rect 9492 -18604 9508 -18587
rect 8920 -18620 9508 -18604
rect 9938 -18604 9954 -18587
rect 10510 -18587 10712 -18570
rect 10770 -18570 11730 -18532
rect 10770 -18587 10972 -18570
rect 10510 -18604 10526 -18587
rect 9938 -18620 10526 -18604
rect 10956 -18604 10972 -18587
rect 11528 -18587 11730 -18570
rect 11788 -18570 12748 -18532
rect 11788 -18587 11990 -18570
rect 11528 -18604 11544 -18587
rect 10956 -18620 11544 -18604
rect 11974 -18604 11990 -18587
rect 12546 -18587 12748 -18570
rect 12806 -18570 13766 -18532
rect 12806 -18587 13008 -18570
rect 12546 -18604 12562 -18587
rect 11974 -18620 12562 -18604
rect 12992 -18604 13008 -18587
rect 13564 -18587 13766 -18570
rect 13824 -18570 14784 -18532
rect 13824 -18587 14026 -18570
rect 13564 -18604 13580 -18587
rect 12992 -18620 13580 -18604
rect 14010 -18604 14026 -18587
rect 14582 -18587 14784 -18570
rect 14842 -18570 15802 -18532
rect 14842 -18587 15044 -18570
rect 14582 -18604 14598 -18587
rect 14010 -18620 14598 -18604
rect 15028 -18604 15044 -18587
rect 15600 -18587 15802 -18570
rect 15860 -18570 16820 -18532
rect 15860 -18587 16062 -18570
rect 15600 -18604 15616 -18587
rect 15028 -18620 15616 -18604
rect 16046 -18604 16062 -18587
rect 16618 -18587 16820 -18570
rect 16878 -18570 17838 -18532
rect 16878 -18587 17080 -18570
rect 16618 -18604 16634 -18587
rect 16046 -18620 16634 -18604
rect 17064 -18604 17080 -18587
rect 17636 -18587 17838 -18570
rect 17896 -18570 18856 -18532
rect 17896 -18587 18098 -18570
rect 17636 -18604 17652 -18587
rect 17064 -18620 17652 -18604
rect 18082 -18604 18098 -18587
rect 18654 -18587 18856 -18570
rect 18914 -18570 19874 -18532
rect 18914 -18587 19116 -18570
rect 18654 -18604 18670 -18587
rect 18082 -18620 18670 -18604
rect 19100 -18604 19116 -18587
rect 19672 -18587 19874 -18570
rect 19932 -18570 20892 -18532
rect 19932 -18587 20134 -18570
rect 19672 -18604 19688 -18587
rect 19100 -18620 19688 -18604
rect 20118 -18604 20134 -18587
rect 20690 -18587 20892 -18570
rect 20950 -18570 21910 -18532
rect 20950 -18587 21152 -18570
rect 20690 -18604 20706 -18587
rect 20118 -18620 20706 -18604
rect 21136 -18604 21152 -18587
rect 21708 -18587 21910 -18570
rect 21968 -18570 22928 -18532
rect 21968 -18587 22170 -18570
rect 21708 -18604 21724 -18587
rect 21136 -18620 21724 -18604
rect 22154 -18604 22170 -18587
rect 22726 -18587 22928 -18570
rect 22726 -18604 22742 -18587
rect 22154 -18620 22742 -18604
rect -9138 -18876 -8178 -18838
rect -9138 -18893 -8936 -18876
rect -8952 -18910 -8936 -18893
rect -8380 -18893 -8178 -18876
rect -8120 -18876 -7160 -18838
rect -8120 -18893 -7918 -18876
rect -8380 -18910 -8364 -18893
rect -8952 -18926 -8364 -18910
rect -7934 -18910 -7918 -18893
rect -7362 -18893 -7160 -18876
rect -7102 -18876 -6142 -18838
rect -7102 -18893 -6900 -18876
rect -7362 -18910 -7346 -18893
rect -7934 -18926 -7346 -18910
rect -6916 -18910 -6900 -18893
rect -6344 -18893 -6142 -18876
rect -6084 -18876 -5124 -18838
rect -6084 -18893 -5882 -18876
rect -6344 -18910 -6328 -18893
rect -6916 -18926 -6328 -18910
rect -5898 -18910 -5882 -18893
rect -5326 -18893 -5124 -18876
rect -5066 -18876 -4106 -18838
rect -5066 -18893 -4864 -18876
rect -5326 -18910 -5310 -18893
rect -5898 -18926 -5310 -18910
rect -4880 -18910 -4864 -18893
rect -4308 -18893 -4106 -18876
rect -4048 -18876 -3088 -18838
rect -4048 -18893 -3846 -18876
rect -4308 -18910 -4292 -18893
rect -4880 -18926 -4292 -18910
rect -3862 -18910 -3846 -18893
rect -3290 -18893 -3088 -18876
rect -3030 -18876 -2070 -18838
rect -3030 -18893 -2828 -18876
rect -3290 -18910 -3274 -18893
rect -3862 -18926 -3274 -18910
rect -2844 -18910 -2828 -18893
rect -2272 -18893 -2070 -18876
rect -2012 -18876 -1052 -18838
rect -2012 -18893 -1810 -18876
rect -2272 -18910 -2256 -18893
rect -2844 -18926 -2256 -18910
rect -1826 -18910 -1810 -18893
rect -1254 -18893 -1052 -18876
rect -994 -18876 -34 -18838
rect -994 -18893 -792 -18876
rect -1254 -18910 -1238 -18893
rect -1826 -18926 -1238 -18910
rect -808 -18910 -792 -18893
rect -236 -18893 -34 -18876
rect -236 -18910 -220 -18893
rect -808 -18926 -220 -18910
rect 2812 -19092 3400 -19076
rect 2812 -19109 2828 -19092
rect 2626 -19126 2828 -19109
rect 3384 -19109 3400 -19092
rect 3830 -19092 4418 -19076
rect 3830 -19109 3846 -19092
rect 3384 -19126 3586 -19109
rect 2626 -19164 3586 -19126
rect 3644 -19126 3846 -19109
rect 4402 -19109 4418 -19092
rect 4848 -19092 5436 -19076
rect 4848 -19109 4864 -19092
rect 4402 -19126 4604 -19109
rect 3644 -19164 4604 -19126
rect 4662 -19126 4864 -19109
rect 5420 -19109 5436 -19092
rect 5866 -19092 6454 -19076
rect 5866 -19109 5882 -19092
rect 5420 -19126 5622 -19109
rect 4662 -19164 5622 -19126
rect 5680 -19126 5882 -19109
rect 6438 -19109 6454 -19092
rect 6884 -19092 7472 -19076
rect 6884 -19109 6900 -19092
rect 6438 -19126 6640 -19109
rect 5680 -19164 6640 -19126
rect 6698 -19126 6900 -19109
rect 7456 -19109 7472 -19092
rect 7902 -19092 8490 -19076
rect 7902 -19109 7918 -19092
rect 7456 -19126 7658 -19109
rect 6698 -19164 7658 -19126
rect 7716 -19126 7918 -19109
rect 8474 -19109 8490 -19092
rect 8920 -19092 9508 -19076
rect 8920 -19109 8936 -19092
rect 8474 -19126 8676 -19109
rect 7716 -19164 8676 -19126
rect 8734 -19126 8936 -19109
rect 9492 -19109 9508 -19092
rect 9938 -19092 10526 -19076
rect 9938 -19109 9954 -19092
rect 9492 -19126 9694 -19109
rect 8734 -19164 9694 -19126
rect 9752 -19126 9954 -19109
rect 10510 -19109 10526 -19092
rect 10956 -19092 11544 -19076
rect 10956 -19109 10972 -19092
rect 10510 -19126 10712 -19109
rect 9752 -19164 10712 -19126
rect 10770 -19126 10972 -19109
rect 11528 -19109 11544 -19092
rect 11974 -19092 12562 -19076
rect 11974 -19109 11990 -19092
rect 11528 -19126 11730 -19109
rect 10770 -19164 11730 -19126
rect 11788 -19126 11990 -19109
rect 12546 -19109 12562 -19092
rect 12992 -19092 13580 -19076
rect 12992 -19109 13008 -19092
rect 12546 -19126 12748 -19109
rect 11788 -19164 12748 -19126
rect 12806 -19126 13008 -19109
rect 13564 -19109 13580 -19092
rect 14010 -19092 14598 -19076
rect 14010 -19109 14026 -19092
rect 13564 -19126 13766 -19109
rect 12806 -19164 13766 -19126
rect 13824 -19126 14026 -19109
rect 14582 -19109 14598 -19092
rect 15028 -19092 15616 -19076
rect 15028 -19109 15044 -19092
rect 14582 -19126 14784 -19109
rect 13824 -19164 14784 -19126
rect 14842 -19126 15044 -19109
rect 15600 -19109 15616 -19092
rect 16046 -19092 16634 -19076
rect 16046 -19109 16062 -19092
rect 15600 -19126 15802 -19109
rect 14842 -19164 15802 -19126
rect 15860 -19126 16062 -19109
rect 16618 -19109 16634 -19092
rect 17064 -19092 17652 -19076
rect 17064 -19109 17080 -19092
rect 16618 -19126 16820 -19109
rect 15860 -19164 16820 -19126
rect 16878 -19126 17080 -19109
rect 17636 -19109 17652 -19092
rect 18082 -19092 18670 -19076
rect 18082 -19109 18098 -19092
rect 17636 -19126 17838 -19109
rect 16878 -19164 17838 -19126
rect 17896 -19126 18098 -19109
rect 18654 -19109 18670 -19092
rect 19100 -19092 19688 -19076
rect 19100 -19109 19116 -19092
rect 18654 -19126 18856 -19109
rect 17896 -19164 18856 -19126
rect 18914 -19126 19116 -19109
rect 19672 -19109 19688 -19092
rect 20118 -19092 20706 -19076
rect 20118 -19109 20134 -19092
rect 19672 -19126 19874 -19109
rect 18914 -19164 19874 -19126
rect 19932 -19126 20134 -19109
rect 20690 -19109 20706 -19092
rect 21136 -19092 21724 -19076
rect 21136 -19109 21152 -19092
rect 20690 -19126 20892 -19109
rect 19932 -19164 20892 -19126
rect 20950 -19126 21152 -19109
rect 21708 -19109 21724 -19092
rect 22154 -19092 22742 -19076
rect 22154 -19109 22170 -19092
rect 21708 -19126 21910 -19109
rect 20950 -19164 21910 -19126
rect 21968 -19126 22170 -19109
rect 22726 -19109 22742 -19092
rect 22726 -19126 22928 -19109
rect 21968 -19164 22928 -19126
rect 2626 -19802 3586 -19764
rect 2626 -19819 2828 -19802
rect 2812 -19836 2828 -19819
rect 3384 -19819 3586 -19802
rect 3644 -19802 4604 -19764
rect 3644 -19819 3846 -19802
rect 3384 -19836 3400 -19819
rect 2812 -19852 3400 -19836
rect 3830 -19836 3846 -19819
rect 4402 -19819 4604 -19802
rect 4662 -19802 5622 -19764
rect 4662 -19819 4864 -19802
rect 4402 -19836 4418 -19819
rect 3830 -19852 4418 -19836
rect 4848 -19836 4864 -19819
rect 5420 -19819 5622 -19802
rect 5680 -19802 6640 -19764
rect 5680 -19819 5882 -19802
rect 5420 -19836 5436 -19819
rect 4848 -19852 5436 -19836
rect 5866 -19836 5882 -19819
rect 6438 -19819 6640 -19802
rect 6698 -19802 7658 -19764
rect 6698 -19819 6900 -19802
rect 6438 -19836 6454 -19819
rect 5866 -19852 6454 -19836
rect 6884 -19836 6900 -19819
rect 7456 -19819 7658 -19802
rect 7716 -19802 8676 -19764
rect 7716 -19819 7918 -19802
rect 7456 -19836 7472 -19819
rect 6884 -19852 7472 -19836
rect 7902 -19836 7918 -19819
rect 8474 -19819 8676 -19802
rect 8734 -19802 9694 -19764
rect 8734 -19819 8936 -19802
rect 8474 -19836 8490 -19819
rect 7902 -19852 8490 -19836
rect 8920 -19836 8936 -19819
rect 9492 -19819 9694 -19802
rect 9752 -19802 10712 -19764
rect 9752 -19819 9954 -19802
rect 9492 -19836 9508 -19819
rect 8920 -19852 9508 -19836
rect 9938 -19836 9954 -19819
rect 10510 -19819 10712 -19802
rect 10770 -19802 11730 -19764
rect 10770 -19819 10972 -19802
rect 10510 -19836 10526 -19819
rect 9938 -19852 10526 -19836
rect 10956 -19836 10972 -19819
rect 11528 -19819 11730 -19802
rect 11788 -19802 12748 -19764
rect 11788 -19819 11990 -19802
rect 11528 -19836 11544 -19819
rect 10956 -19852 11544 -19836
rect 11974 -19836 11990 -19819
rect 12546 -19819 12748 -19802
rect 12806 -19802 13766 -19764
rect 12806 -19819 13008 -19802
rect 12546 -19836 12562 -19819
rect 11974 -19852 12562 -19836
rect 12992 -19836 13008 -19819
rect 13564 -19819 13766 -19802
rect 13824 -19802 14784 -19764
rect 13824 -19819 14026 -19802
rect 13564 -19836 13580 -19819
rect 12992 -19852 13580 -19836
rect 14010 -19836 14026 -19819
rect 14582 -19819 14784 -19802
rect 14842 -19802 15802 -19764
rect 14842 -19819 15044 -19802
rect 14582 -19836 14598 -19819
rect 14010 -19852 14598 -19836
rect 15028 -19836 15044 -19819
rect 15600 -19819 15802 -19802
rect 15860 -19802 16820 -19764
rect 15860 -19819 16062 -19802
rect 15600 -19836 15616 -19819
rect 15028 -19852 15616 -19836
rect 16046 -19836 16062 -19819
rect 16618 -19819 16820 -19802
rect 16878 -19802 17838 -19764
rect 16878 -19819 17080 -19802
rect 16618 -19836 16634 -19819
rect 16046 -19852 16634 -19836
rect 17064 -19836 17080 -19819
rect 17636 -19819 17838 -19802
rect 17896 -19802 18856 -19764
rect 17896 -19819 18098 -19802
rect 17636 -19836 17652 -19819
rect 17064 -19852 17652 -19836
rect 18082 -19836 18098 -19819
rect 18654 -19819 18856 -19802
rect 18914 -19802 19874 -19764
rect 18914 -19819 19116 -19802
rect 18654 -19836 18670 -19819
rect 18082 -19852 18670 -19836
rect 19100 -19836 19116 -19819
rect 19672 -19819 19874 -19802
rect 19932 -19802 20892 -19764
rect 19932 -19819 20134 -19802
rect 19672 -19836 19688 -19819
rect 19100 -19852 19688 -19836
rect 20118 -19836 20134 -19819
rect 20690 -19819 20892 -19802
rect 20950 -19802 21910 -19764
rect 20950 -19819 21152 -19802
rect 20690 -19836 20706 -19819
rect 20118 -19852 20706 -19836
rect 21136 -19836 21152 -19819
rect 21708 -19819 21910 -19802
rect 21968 -19802 22928 -19764
rect 21968 -19819 22170 -19802
rect 21708 -19836 21724 -19819
rect 21136 -19852 21724 -19836
rect 22154 -19836 22170 -19819
rect 22726 -19819 22928 -19802
rect 22726 -19836 22742 -19819
rect 22154 -19852 22742 -19836
rect -10276 -20190 -9688 -20174
rect -10276 -20207 -10260 -20190
rect -10462 -20224 -10260 -20207
rect -9704 -20207 -9688 -20190
rect -9258 -20190 -8670 -20174
rect -9258 -20207 -9242 -20190
rect -9704 -20224 -9502 -20207
rect -10462 -20262 -9502 -20224
rect -9444 -20224 -9242 -20207
rect -8686 -20207 -8670 -20190
rect -8240 -20190 -7652 -20174
rect -8240 -20207 -8224 -20190
rect -8686 -20224 -8484 -20207
rect -9444 -20262 -8484 -20224
rect -8426 -20224 -8224 -20207
rect -7668 -20207 -7652 -20190
rect -7222 -20190 -6634 -20174
rect -7222 -20207 -7206 -20190
rect -7668 -20224 -7466 -20207
rect -8426 -20262 -7466 -20224
rect -7408 -20224 -7206 -20207
rect -6650 -20207 -6634 -20190
rect -6204 -20190 -5616 -20174
rect -6204 -20207 -6188 -20190
rect -6650 -20224 -6448 -20207
rect -7408 -20262 -6448 -20224
rect -6390 -20224 -6188 -20207
rect -5632 -20207 -5616 -20190
rect -5186 -20190 -4598 -20174
rect -5186 -20207 -5170 -20190
rect -5632 -20224 -5430 -20207
rect -6390 -20262 -5430 -20224
rect -5372 -20224 -5170 -20207
rect -4614 -20207 -4598 -20190
rect -4168 -20190 -3580 -20174
rect -4168 -20207 -4152 -20190
rect -4614 -20224 -4412 -20207
rect -5372 -20262 -4412 -20224
rect -4354 -20224 -4152 -20207
rect -3596 -20207 -3580 -20190
rect -3150 -20190 -2562 -20174
rect -3150 -20207 -3134 -20190
rect -3596 -20224 -3394 -20207
rect -4354 -20262 -3394 -20224
rect -3336 -20224 -3134 -20207
rect -2578 -20207 -2562 -20190
rect -2132 -20190 -1544 -20174
rect -2132 -20207 -2116 -20190
rect -2578 -20224 -2376 -20207
rect -3336 -20262 -2376 -20224
rect -2318 -20224 -2116 -20207
rect -1560 -20207 -1544 -20190
rect -1114 -20190 -526 -20174
rect -1114 -20207 -1098 -20190
rect -1560 -20224 -1358 -20207
rect -2318 -20262 -1358 -20224
rect -1300 -20224 -1098 -20207
rect -542 -20207 -526 -20190
rect -96 -20190 492 -20174
rect -96 -20207 -80 -20190
rect -542 -20224 -340 -20207
rect -1300 -20262 -340 -20224
rect -282 -20224 -80 -20207
rect 476 -20207 492 -20190
rect 476 -20224 678 -20207
rect -282 -20262 678 -20224
rect 2812 -20326 3400 -20310
rect 2812 -20343 2828 -20326
rect 2626 -20360 2828 -20343
rect 3384 -20343 3400 -20326
rect 3830 -20326 4418 -20310
rect 3830 -20343 3846 -20326
rect 3384 -20360 3586 -20343
rect 2626 -20398 3586 -20360
rect 3644 -20360 3846 -20343
rect 4402 -20343 4418 -20326
rect 4848 -20326 5436 -20310
rect 4848 -20343 4864 -20326
rect 4402 -20360 4604 -20343
rect 3644 -20398 4604 -20360
rect 4662 -20360 4864 -20343
rect 5420 -20343 5436 -20326
rect 5866 -20326 6454 -20310
rect 5866 -20343 5882 -20326
rect 5420 -20360 5622 -20343
rect 4662 -20398 5622 -20360
rect 5680 -20360 5882 -20343
rect 6438 -20343 6454 -20326
rect 6884 -20326 7472 -20310
rect 6884 -20343 6900 -20326
rect 6438 -20360 6640 -20343
rect 5680 -20398 6640 -20360
rect 6698 -20360 6900 -20343
rect 7456 -20343 7472 -20326
rect 7902 -20326 8490 -20310
rect 7902 -20343 7918 -20326
rect 7456 -20360 7658 -20343
rect 6698 -20398 7658 -20360
rect 7716 -20360 7918 -20343
rect 8474 -20343 8490 -20326
rect 8920 -20326 9508 -20310
rect 8920 -20343 8936 -20326
rect 8474 -20360 8676 -20343
rect 7716 -20398 8676 -20360
rect 8734 -20360 8936 -20343
rect 9492 -20343 9508 -20326
rect 9938 -20326 10526 -20310
rect 9938 -20343 9954 -20326
rect 9492 -20360 9694 -20343
rect 8734 -20398 9694 -20360
rect 9752 -20360 9954 -20343
rect 10510 -20343 10526 -20326
rect 10956 -20326 11544 -20310
rect 10956 -20343 10972 -20326
rect 10510 -20360 10712 -20343
rect 9752 -20398 10712 -20360
rect 10770 -20360 10972 -20343
rect 11528 -20343 11544 -20326
rect 11974 -20326 12562 -20310
rect 11974 -20343 11990 -20326
rect 11528 -20360 11730 -20343
rect 10770 -20398 11730 -20360
rect 11788 -20360 11990 -20343
rect 12546 -20343 12562 -20326
rect 12992 -20326 13580 -20310
rect 12992 -20343 13008 -20326
rect 12546 -20360 12748 -20343
rect 11788 -20398 12748 -20360
rect 12806 -20360 13008 -20343
rect 13564 -20343 13580 -20326
rect 14010 -20326 14598 -20310
rect 14010 -20343 14026 -20326
rect 13564 -20360 13766 -20343
rect 12806 -20398 13766 -20360
rect 13824 -20360 14026 -20343
rect 14582 -20343 14598 -20326
rect 15028 -20326 15616 -20310
rect 15028 -20343 15044 -20326
rect 14582 -20360 14784 -20343
rect 13824 -20398 14784 -20360
rect 14842 -20360 15044 -20343
rect 15600 -20343 15616 -20326
rect 16046 -20326 16634 -20310
rect 16046 -20343 16062 -20326
rect 15600 -20360 15802 -20343
rect 14842 -20398 15802 -20360
rect 15860 -20360 16062 -20343
rect 16618 -20343 16634 -20326
rect 17064 -20326 17652 -20310
rect 17064 -20343 17080 -20326
rect 16618 -20360 16820 -20343
rect 15860 -20398 16820 -20360
rect 16878 -20360 17080 -20343
rect 17636 -20343 17652 -20326
rect 18082 -20326 18670 -20310
rect 18082 -20343 18098 -20326
rect 17636 -20360 17838 -20343
rect 16878 -20398 17838 -20360
rect 17896 -20360 18098 -20343
rect 18654 -20343 18670 -20326
rect 19100 -20326 19688 -20310
rect 19100 -20343 19116 -20326
rect 18654 -20360 18856 -20343
rect 17896 -20398 18856 -20360
rect 18914 -20360 19116 -20343
rect 19672 -20343 19688 -20326
rect 20118 -20326 20706 -20310
rect 20118 -20343 20134 -20326
rect 19672 -20360 19874 -20343
rect 18914 -20398 19874 -20360
rect 19932 -20360 20134 -20343
rect 20690 -20343 20706 -20326
rect 21136 -20326 21724 -20310
rect 21136 -20343 21152 -20326
rect 20690 -20360 20892 -20343
rect 19932 -20398 20892 -20360
rect 20950 -20360 21152 -20343
rect 21708 -20343 21724 -20326
rect 22154 -20326 22742 -20310
rect 22154 -20343 22170 -20326
rect 21708 -20360 21910 -20343
rect 20950 -20398 21910 -20360
rect 21968 -20360 22170 -20343
rect 22726 -20343 22742 -20326
rect 22726 -20360 22928 -20343
rect 21968 -20398 22928 -20360
rect -10462 -20900 -9502 -20862
rect -10462 -20917 -10260 -20900
rect -10276 -20934 -10260 -20917
rect -9704 -20917 -9502 -20900
rect -9444 -20900 -8484 -20862
rect -9444 -20917 -9242 -20900
rect -9704 -20934 -9688 -20917
rect -10276 -20950 -9688 -20934
rect -9258 -20934 -9242 -20917
rect -8686 -20917 -8484 -20900
rect -8426 -20900 -7466 -20862
rect -8426 -20917 -8224 -20900
rect -8686 -20934 -8670 -20917
rect -9258 -20950 -8670 -20934
rect -8240 -20934 -8224 -20917
rect -7668 -20917 -7466 -20900
rect -7408 -20900 -6448 -20862
rect -7408 -20917 -7206 -20900
rect -7668 -20934 -7652 -20917
rect -8240 -20950 -7652 -20934
rect -7222 -20934 -7206 -20917
rect -6650 -20917 -6448 -20900
rect -6390 -20900 -5430 -20862
rect -6390 -20917 -6188 -20900
rect -6650 -20934 -6634 -20917
rect -7222 -20950 -6634 -20934
rect -6204 -20934 -6188 -20917
rect -5632 -20917 -5430 -20900
rect -5372 -20900 -4412 -20862
rect -5372 -20917 -5170 -20900
rect -5632 -20934 -5616 -20917
rect -6204 -20950 -5616 -20934
rect -5186 -20934 -5170 -20917
rect -4614 -20917 -4412 -20900
rect -4354 -20900 -3394 -20862
rect -4354 -20917 -4152 -20900
rect -4614 -20934 -4598 -20917
rect -5186 -20950 -4598 -20934
rect -4168 -20934 -4152 -20917
rect -3596 -20917 -3394 -20900
rect -3336 -20900 -2376 -20862
rect -3336 -20917 -3134 -20900
rect -3596 -20934 -3580 -20917
rect -4168 -20950 -3580 -20934
rect -3150 -20934 -3134 -20917
rect -2578 -20917 -2376 -20900
rect -2318 -20900 -1358 -20862
rect -2318 -20917 -2116 -20900
rect -2578 -20934 -2562 -20917
rect -3150 -20950 -2562 -20934
rect -2132 -20934 -2116 -20917
rect -1560 -20917 -1358 -20900
rect -1300 -20900 -340 -20862
rect -1300 -20917 -1098 -20900
rect -1560 -20934 -1544 -20917
rect -2132 -20950 -1544 -20934
rect -1114 -20934 -1098 -20917
rect -542 -20917 -340 -20900
rect -282 -20900 678 -20862
rect -282 -20917 -80 -20900
rect -542 -20934 -526 -20917
rect -1114 -20950 -526 -20934
rect -96 -20934 -80 -20917
rect 476 -20917 678 -20900
rect 476 -20934 492 -20917
rect -96 -20950 492 -20934
rect 2626 -21036 3586 -20998
rect 2626 -21053 2828 -21036
rect 2812 -21070 2828 -21053
rect 3384 -21053 3586 -21036
rect 3644 -21036 4604 -20998
rect 3644 -21053 3846 -21036
rect 3384 -21070 3400 -21053
rect 2812 -21086 3400 -21070
rect 3830 -21070 3846 -21053
rect 4402 -21053 4604 -21036
rect 4662 -21036 5622 -20998
rect 4662 -21053 4864 -21036
rect 4402 -21070 4418 -21053
rect 3830 -21086 4418 -21070
rect 4848 -21070 4864 -21053
rect 5420 -21053 5622 -21036
rect 5680 -21036 6640 -20998
rect 5680 -21053 5882 -21036
rect 5420 -21070 5436 -21053
rect 4848 -21086 5436 -21070
rect 5866 -21070 5882 -21053
rect 6438 -21053 6640 -21036
rect 6698 -21036 7658 -20998
rect 6698 -21053 6900 -21036
rect 6438 -21070 6454 -21053
rect 5866 -21086 6454 -21070
rect 6884 -21070 6900 -21053
rect 7456 -21053 7658 -21036
rect 7716 -21036 8676 -20998
rect 7716 -21053 7918 -21036
rect 7456 -21070 7472 -21053
rect 6884 -21086 7472 -21070
rect 7902 -21070 7918 -21053
rect 8474 -21053 8676 -21036
rect 8734 -21036 9694 -20998
rect 8734 -21053 8936 -21036
rect 8474 -21070 8490 -21053
rect 7902 -21086 8490 -21070
rect 8920 -21070 8936 -21053
rect 9492 -21053 9694 -21036
rect 9752 -21036 10712 -20998
rect 9752 -21053 9954 -21036
rect 9492 -21070 9508 -21053
rect 8920 -21086 9508 -21070
rect 9938 -21070 9954 -21053
rect 10510 -21053 10712 -21036
rect 10770 -21036 11730 -20998
rect 10770 -21053 10972 -21036
rect 10510 -21070 10526 -21053
rect 9938 -21086 10526 -21070
rect 10956 -21070 10972 -21053
rect 11528 -21053 11730 -21036
rect 11788 -21036 12748 -20998
rect 11788 -21053 11990 -21036
rect 11528 -21070 11544 -21053
rect 10956 -21086 11544 -21070
rect 11974 -21070 11990 -21053
rect 12546 -21053 12748 -21036
rect 12806 -21036 13766 -20998
rect 12806 -21053 13008 -21036
rect 12546 -21070 12562 -21053
rect 11974 -21086 12562 -21070
rect 12992 -21070 13008 -21053
rect 13564 -21053 13766 -21036
rect 13824 -21036 14784 -20998
rect 13824 -21053 14026 -21036
rect 13564 -21070 13580 -21053
rect 12992 -21086 13580 -21070
rect 14010 -21070 14026 -21053
rect 14582 -21053 14784 -21036
rect 14842 -21036 15802 -20998
rect 14842 -21053 15044 -21036
rect 14582 -21070 14598 -21053
rect 14010 -21086 14598 -21070
rect 15028 -21070 15044 -21053
rect 15600 -21053 15802 -21036
rect 15860 -21036 16820 -20998
rect 15860 -21053 16062 -21036
rect 15600 -21070 15616 -21053
rect 15028 -21086 15616 -21070
rect 16046 -21070 16062 -21053
rect 16618 -21053 16820 -21036
rect 16878 -21036 17838 -20998
rect 16878 -21053 17080 -21036
rect 16618 -21070 16634 -21053
rect 16046 -21086 16634 -21070
rect 17064 -21070 17080 -21053
rect 17636 -21053 17838 -21036
rect 17896 -21036 18856 -20998
rect 17896 -21053 18098 -21036
rect 17636 -21070 17652 -21053
rect 17064 -21086 17652 -21070
rect 18082 -21070 18098 -21053
rect 18654 -21053 18856 -21036
rect 18914 -21036 19874 -20998
rect 18914 -21053 19116 -21036
rect 18654 -21070 18670 -21053
rect 18082 -21086 18670 -21070
rect 19100 -21070 19116 -21053
rect 19672 -21053 19874 -21036
rect 19932 -21036 20892 -20998
rect 19932 -21053 20134 -21036
rect 19672 -21070 19688 -21053
rect 19100 -21086 19688 -21070
rect 20118 -21070 20134 -21053
rect 20690 -21053 20892 -21036
rect 20950 -21036 21910 -20998
rect 20950 -21053 21152 -21036
rect 20690 -21070 20706 -21053
rect 20118 -21086 20706 -21070
rect 21136 -21070 21152 -21053
rect 21708 -21053 21910 -21036
rect 21968 -21036 22928 -20998
rect 21968 -21053 22170 -21036
rect 21708 -21070 21724 -21053
rect 21136 -21086 21724 -21070
rect 22154 -21070 22170 -21053
rect 22726 -21053 22928 -21036
rect 22726 -21070 22742 -21053
rect 22154 -21086 22742 -21070
rect -10276 -21302 -9688 -21286
rect -10276 -21319 -10260 -21302
rect -10462 -21336 -10260 -21319
rect -9704 -21319 -9688 -21302
rect -9258 -21302 -8670 -21286
rect -9258 -21319 -9242 -21302
rect -9704 -21336 -9502 -21319
rect -10462 -21374 -9502 -21336
rect -9444 -21336 -9242 -21319
rect -8686 -21319 -8670 -21302
rect -8240 -21302 -7652 -21286
rect -8240 -21319 -8224 -21302
rect -8686 -21336 -8484 -21319
rect -9444 -21374 -8484 -21336
rect -8426 -21336 -8224 -21319
rect -7668 -21319 -7652 -21302
rect -7222 -21302 -6634 -21286
rect -7222 -21319 -7206 -21302
rect -7668 -21336 -7466 -21319
rect -8426 -21374 -7466 -21336
rect -7408 -21336 -7206 -21319
rect -6650 -21319 -6634 -21302
rect -6204 -21302 -5616 -21286
rect -6204 -21319 -6188 -21302
rect -6650 -21336 -6448 -21319
rect -7408 -21374 -6448 -21336
rect -6390 -21336 -6188 -21319
rect -5632 -21319 -5616 -21302
rect -5186 -21302 -4598 -21286
rect -5186 -21319 -5170 -21302
rect -5632 -21336 -5430 -21319
rect -6390 -21374 -5430 -21336
rect -5372 -21336 -5170 -21319
rect -4614 -21319 -4598 -21302
rect -4168 -21302 -3580 -21286
rect -4168 -21319 -4152 -21302
rect -4614 -21336 -4412 -21319
rect -5372 -21374 -4412 -21336
rect -4354 -21336 -4152 -21319
rect -3596 -21319 -3580 -21302
rect -3150 -21302 -2562 -21286
rect -3150 -21319 -3134 -21302
rect -3596 -21336 -3394 -21319
rect -4354 -21374 -3394 -21336
rect -3336 -21336 -3134 -21319
rect -2578 -21319 -2562 -21302
rect -2132 -21302 -1544 -21286
rect -2132 -21319 -2116 -21302
rect -2578 -21336 -2376 -21319
rect -3336 -21374 -2376 -21336
rect -2318 -21336 -2116 -21319
rect -1560 -21319 -1544 -21302
rect -1114 -21302 -526 -21286
rect -1114 -21319 -1098 -21302
rect -1560 -21336 -1358 -21319
rect -2318 -21374 -1358 -21336
rect -1300 -21336 -1098 -21319
rect -542 -21319 -526 -21302
rect -96 -21302 492 -21286
rect -96 -21319 -80 -21302
rect -542 -21336 -340 -21319
rect -1300 -21374 -340 -21336
rect -282 -21336 -80 -21319
rect 476 -21319 492 -21302
rect 476 -21336 678 -21319
rect -282 -21374 678 -21336
rect 2812 -21560 3400 -21544
rect 2812 -21577 2828 -21560
rect 2626 -21594 2828 -21577
rect 3384 -21577 3400 -21560
rect 3830 -21560 4418 -21544
rect 3830 -21577 3846 -21560
rect 3384 -21594 3586 -21577
rect 2626 -21632 3586 -21594
rect 3644 -21594 3846 -21577
rect 4402 -21577 4418 -21560
rect 4848 -21560 5436 -21544
rect 4848 -21577 4864 -21560
rect 4402 -21594 4604 -21577
rect 3644 -21632 4604 -21594
rect 4662 -21594 4864 -21577
rect 5420 -21577 5436 -21560
rect 5866 -21560 6454 -21544
rect 5866 -21577 5882 -21560
rect 5420 -21594 5622 -21577
rect 4662 -21632 5622 -21594
rect 5680 -21594 5882 -21577
rect 6438 -21577 6454 -21560
rect 6884 -21560 7472 -21544
rect 6884 -21577 6900 -21560
rect 6438 -21594 6640 -21577
rect 5680 -21632 6640 -21594
rect 6698 -21594 6900 -21577
rect 7456 -21577 7472 -21560
rect 7902 -21560 8490 -21544
rect 7902 -21577 7918 -21560
rect 7456 -21594 7658 -21577
rect 6698 -21632 7658 -21594
rect 7716 -21594 7918 -21577
rect 8474 -21577 8490 -21560
rect 8920 -21560 9508 -21544
rect 8920 -21577 8936 -21560
rect 8474 -21594 8676 -21577
rect 7716 -21632 8676 -21594
rect 8734 -21594 8936 -21577
rect 9492 -21577 9508 -21560
rect 9938 -21560 10526 -21544
rect 9938 -21577 9954 -21560
rect 9492 -21594 9694 -21577
rect 8734 -21632 9694 -21594
rect 9752 -21594 9954 -21577
rect 10510 -21577 10526 -21560
rect 10956 -21560 11544 -21544
rect 10956 -21577 10972 -21560
rect 10510 -21594 10712 -21577
rect 9752 -21632 10712 -21594
rect 10770 -21594 10972 -21577
rect 11528 -21577 11544 -21560
rect 11974 -21560 12562 -21544
rect 11974 -21577 11990 -21560
rect 11528 -21594 11730 -21577
rect 10770 -21632 11730 -21594
rect 11788 -21594 11990 -21577
rect 12546 -21577 12562 -21560
rect 12992 -21560 13580 -21544
rect 12992 -21577 13008 -21560
rect 12546 -21594 12748 -21577
rect 11788 -21632 12748 -21594
rect 12806 -21594 13008 -21577
rect 13564 -21577 13580 -21560
rect 14010 -21560 14598 -21544
rect 14010 -21577 14026 -21560
rect 13564 -21594 13766 -21577
rect 12806 -21632 13766 -21594
rect 13824 -21594 14026 -21577
rect 14582 -21577 14598 -21560
rect 15028 -21560 15616 -21544
rect 15028 -21577 15044 -21560
rect 14582 -21594 14784 -21577
rect 13824 -21632 14784 -21594
rect 14842 -21594 15044 -21577
rect 15600 -21577 15616 -21560
rect 16046 -21560 16634 -21544
rect 16046 -21577 16062 -21560
rect 15600 -21594 15802 -21577
rect 14842 -21632 15802 -21594
rect 15860 -21594 16062 -21577
rect 16618 -21577 16634 -21560
rect 17064 -21560 17652 -21544
rect 17064 -21577 17080 -21560
rect 16618 -21594 16820 -21577
rect 15860 -21632 16820 -21594
rect 16878 -21594 17080 -21577
rect 17636 -21577 17652 -21560
rect 18082 -21560 18670 -21544
rect 18082 -21577 18098 -21560
rect 17636 -21594 17838 -21577
rect 16878 -21632 17838 -21594
rect 17896 -21594 18098 -21577
rect 18654 -21577 18670 -21560
rect 19100 -21560 19688 -21544
rect 19100 -21577 19116 -21560
rect 18654 -21594 18856 -21577
rect 17896 -21632 18856 -21594
rect 18914 -21594 19116 -21577
rect 19672 -21577 19688 -21560
rect 20118 -21560 20706 -21544
rect 20118 -21577 20134 -21560
rect 19672 -21594 19874 -21577
rect 18914 -21632 19874 -21594
rect 19932 -21594 20134 -21577
rect 20690 -21577 20706 -21560
rect 21136 -21560 21724 -21544
rect 21136 -21577 21152 -21560
rect 20690 -21594 20892 -21577
rect 19932 -21632 20892 -21594
rect 20950 -21594 21152 -21577
rect 21708 -21577 21724 -21560
rect 22154 -21560 22742 -21544
rect 22154 -21577 22170 -21560
rect 21708 -21594 21910 -21577
rect 20950 -21632 21910 -21594
rect 21968 -21594 22170 -21577
rect 22726 -21577 22742 -21560
rect 22726 -21594 22928 -21577
rect 21968 -21632 22928 -21594
rect -10462 -22012 -9502 -21974
rect -10462 -22029 -10260 -22012
rect -10276 -22046 -10260 -22029
rect -9704 -22029 -9502 -22012
rect -9444 -22012 -8484 -21974
rect -9444 -22029 -9242 -22012
rect -9704 -22046 -9688 -22029
rect -10276 -22062 -9688 -22046
rect -9258 -22046 -9242 -22029
rect -8686 -22029 -8484 -22012
rect -8426 -22012 -7466 -21974
rect -8426 -22029 -8224 -22012
rect -8686 -22046 -8670 -22029
rect -9258 -22062 -8670 -22046
rect -8240 -22046 -8224 -22029
rect -7668 -22029 -7466 -22012
rect -7408 -22012 -6448 -21974
rect -7408 -22029 -7206 -22012
rect -7668 -22046 -7652 -22029
rect -8240 -22062 -7652 -22046
rect -7222 -22046 -7206 -22029
rect -6650 -22029 -6448 -22012
rect -6390 -22012 -5430 -21974
rect -6390 -22029 -6188 -22012
rect -6650 -22046 -6634 -22029
rect -7222 -22062 -6634 -22046
rect -6204 -22046 -6188 -22029
rect -5632 -22029 -5430 -22012
rect -5372 -22012 -4412 -21974
rect -5372 -22029 -5170 -22012
rect -5632 -22046 -5616 -22029
rect -6204 -22062 -5616 -22046
rect -5186 -22046 -5170 -22029
rect -4614 -22029 -4412 -22012
rect -4354 -22012 -3394 -21974
rect -4354 -22029 -4152 -22012
rect -4614 -22046 -4598 -22029
rect -5186 -22062 -4598 -22046
rect -4168 -22046 -4152 -22029
rect -3596 -22029 -3394 -22012
rect -3336 -22012 -2376 -21974
rect -3336 -22029 -3134 -22012
rect -3596 -22046 -3580 -22029
rect -4168 -22062 -3580 -22046
rect -3150 -22046 -3134 -22029
rect -2578 -22029 -2376 -22012
rect -2318 -22012 -1358 -21974
rect -2318 -22029 -2116 -22012
rect -2578 -22046 -2562 -22029
rect -3150 -22062 -2562 -22046
rect -2132 -22046 -2116 -22029
rect -1560 -22029 -1358 -22012
rect -1300 -22012 -340 -21974
rect -1300 -22029 -1098 -22012
rect -1560 -22046 -1544 -22029
rect -2132 -22062 -1544 -22046
rect -1114 -22046 -1098 -22029
rect -542 -22029 -340 -22012
rect -282 -22012 678 -21974
rect -282 -22029 -80 -22012
rect -542 -22046 -526 -22029
rect -1114 -22062 -526 -22046
rect -96 -22046 -80 -22029
rect 476 -22029 678 -22012
rect 476 -22046 492 -22029
rect -96 -22062 492 -22046
rect 2626 -22270 3586 -22232
rect 2626 -22287 2828 -22270
rect 2812 -22304 2828 -22287
rect 3384 -22287 3586 -22270
rect 3644 -22270 4604 -22232
rect 3644 -22287 3846 -22270
rect 3384 -22304 3400 -22287
rect 2812 -22320 3400 -22304
rect 3830 -22304 3846 -22287
rect 4402 -22287 4604 -22270
rect 4662 -22270 5622 -22232
rect 4662 -22287 4864 -22270
rect 4402 -22304 4418 -22287
rect 3830 -22320 4418 -22304
rect 4848 -22304 4864 -22287
rect 5420 -22287 5622 -22270
rect 5680 -22270 6640 -22232
rect 5680 -22287 5882 -22270
rect 5420 -22304 5436 -22287
rect 4848 -22320 5436 -22304
rect 5866 -22304 5882 -22287
rect 6438 -22287 6640 -22270
rect 6698 -22270 7658 -22232
rect 6698 -22287 6900 -22270
rect 6438 -22304 6454 -22287
rect 5866 -22320 6454 -22304
rect 6884 -22304 6900 -22287
rect 7456 -22287 7658 -22270
rect 7716 -22270 8676 -22232
rect 7716 -22287 7918 -22270
rect 7456 -22304 7472 -22287
rect 6884 -22320 7472 -22304
rect 7902 -22304 7918 -22287
rect 8474 -22287 8676 -22270
rect 8734 -22270 9694 -22232
rect 8734 -22287 8936 -22270
rect 8474 -22304 8490 -22287
rect 7902 -22320 8490 -22304
rect 8920 -22304 8936 -22287
rect 9492 -22287 9694 -22270
rect 9752 -22270 10712 -22232
rect 9752 -22287 9954 -22270
rect 9492 -22304 9508 -22287
rect 8920 -22320 9508 -22304
rect 9938 -22304 9954 -22287
rect 10510 -22287 10712 -22270
rect 10770 -22270 11730 -22232
rect 10770 -22287 10972 -22270
rect 10510 -22304 10526 -22287
rect 9938 -22320 10526 -22304
rect 10956 -22304 10972 -22287
rect 11528 -22287 11730 -22270
rect 11788 -22270 12748 -22232
rect 11788 -22287 11990 -22270
rect 11528 -22304 11544 -22287
rect 10956 -22320 11544 -22304
rect 11974 -22304 11990 -22287
rect 12546 -22287 12748 -22270
rect 12806 -22270 13766 -22232
rect 12806 -22287 13008 -22270
rect 12546 -22304 12562 -22287
rect 11974 -22320 12562 -22304
rect 12992 -22304 13008 -22287
rect 13564 -22287 13766 -22270
rect 13824 -22270 14784 -22232
rect 13824 -22287 14026 -22270
rect 13564 -22304 13580 -22287
rect 12992 -22320 13580 -22304
rect 14010 -22304 14026 -22287
rect 14582 -22287 14784 -22270
rect 14842 -22270 15802 -22232
rect 14842 -22287 15044 -22270
rect 14582 -22304 14598 -22287
rect 14010 -22320 14598 -22304
rect 15028 -22304 15044 -22287
rect 15600 -22287 15802 -22270
rect 15860 -22270 16820 -22232
rect 15860 -22287 16062 -22270
rect 15600 -22304 15616 -22287
rect 15028 -22320 15616 -22304
rect 16046 -22304 16062 -22287
rect 16618 -22287 16820 -22270
rect 16878 -22270 17838 -22232
rect 16878 -22287 17080 -22270
rect 16618 -22304 16634 -22287
rect 16046 -22320 16634 -22304
rect 17064 -22304 17080 -22287
rect 17636 -22287 17838 -22270
rect 17896 -22270 18856 -22232
rect 17896 -22287 18098 -22270
rect 17636 -22304 17652 -22287
rect 17064 -22320 17652 -22304
rect 18082 -22304 18098 -22287
rect 18654 -22287 18856 -22270
rect 18914 -22270 19874 -22232
rect 18914 -22287 19116 -22270
rect 18654 -22304 18670 -22287
rect 18082 -22320 18670 -22304
rect 19100 -22304 19116 -22287
rect 19672 -22287 19874 -22270
rect 19932 -22270 20892 -22232
rect 19932 -22287 20134 -22270
rect 19672 -22304 19688 -22287
rect 19100 -22320 19688 -22304
rect 20118 -22304 20134 -22287
rect 20690 -22287 20892 -22270
rect 20950 -22270 21910 -22232
rect 20950 -22287 21152 -22270
rect 20690 -22304 20706 -22287
rect 20118 -22320 20706 -22304
rect 21136 -22304 21152 -22287
rect 21708 -22287 21910 -22270
rect 21968 -22270 22928 -22232
rect 21968 -22287 22170 -22270
rect 21708 -22304 21724 -22287
rect 21136 -22320 21724 -22304
rect 22154 -22304 22170 -22287
rect 22726 -22287 22928 -22270
rect 22726 -22304 22742 -22287
rect 22154 -22320 22742 -22304
rect -10276 -22414 -9688 -22398
rect -10276 -22431 -10260 -22414
rect -10462 -22448 -10260 -22431
rect -9704 -22431 -9688 -22414
rect -9258 -22414 -8670 -22398
rect -9258 -22431 -9242 -22414
rect -9704 -22448 -9502 -22431
rect -10462 -22486 -9502 -22448
rect -9444 -22448 -9242 -22431
rect -8686 -22431 -8670 -22414
rect -8240 -22414 -7652 -22398
rect -8240 -22431 -8224 -22414
rect -8686 -22448 -8484 -22431
rect -9444 -22486 -8484 -22448
rect -8426 -22448 -8224 -22431
rect -7668 -22431 -7652 -22414
rect -7222 -22414 -6634 -22398
rect -7222 -22431 -7206 -22414
rect -7668 -22448 -7466 -22431
rect -8426 -22486 -7466 -22448
rect -7408 -22448 -7206 -22431
rect -6650 -22431 -6634 -22414
rect -6204 -22414 -5616 -22398
rect -6204 -22431 -6188 -22414
rect -6650 -22448 -6448 -22431
rect -7408 -22486 -6448 -22448
rect -6390 -22448 -6188 -22431
rect -5632 -22431 -5616 -22414
rect -5186 -22414 -4598 -22398
rect -5186 -22431 -5170 -22414
rect -5632 -22448 -5430 -22431
rect -6390 -22486 -5430 -22448
rect -5372 -22448 -5170 -22431
rect -4614 -22431 -4598 -22414
rect -4168 -22414 -3580 -22398
rect -4168 -22431 -4152 -22414
rect -4614 -22448 -4412 -22431
rect -5372 -22486 -4412 -22448
rect -4354 -22448 -4152 -22431
rect -3596 -22431 -3580 -22414
rect -3150 -22414 -2562 -22398
rect -3150 -22431 -3134 -22414
rect -3596 -22448 -3394 -22431
rect -4354 -22486 -3394 -22448
rect -3336 -22448 -3134 -22431
rect -2578 -22431 -2562 -22414
rect -2132 -22414 -1544 -22398
rect -2132 -22431 -2116 -22414
rect -2578 -22448 -2376 -22431
rect -3336 -22486 -2376 -22448
rect -2318 -22448 -2116 -22431
rect -1560 -22431 -1544 -22414
rect -1114 -22414 -526 -22398
rect -1114 -22431 -1098 -22414
rect -1560 -22448 -1358 -22431
rect -2318 -22486 -1358 -22448
rect -1300 -22448 -1098 -22431
rect -542 -22431 -526 -22414
rect -96 -22414 492 -22398
rect -96 -22431 -80 -22414
rect -542 -22448 -340 -22431
rect -1300 -22486 -340 -22448
rect -282 -22448 -80 -22431
rect 476 -22431 492 -22414
rect 476 -22448 678 -22431
rect -282 -22486 678 -22448
rect 2812 -22792 3400 -22776
rect 2812 -22809 2828 -22792
rect 2626 -22826 2828 -22809
rect 3384 -22809 3400 -22792
rect 3830 -22792 4418 -22776
rect 3830 -22809 3846 -22792
rect 3384 -22826 3586 -22809
rect 2626 -22864 3586 -22826
rect 3644 -22826 3846 -22809
rect 4402 -22809 4418 -22792
rect 4848 -22792 5436 -22776
rect 4848 -22809 4864 -22792
rect 4402 -22826 4604 -22809
rect 3644 -22864 4604 -22826
rect 4662 -22826 4864 -22809
rect 5420 -22809 5436 -22792
rect 5866 -22792 6454 -22776
rect 5866 -22809 5882 -22792
rect 5420 -22826 5622 -22809
rect 4662 -22864 5622 -22826
rect 5680 -22826 5882 -22809
rect 6438 -22809 6454 -22792
rect 6884 -22792 7472 -22776
rect 6884 -22809 6900 -22792
rect 6438 -22826 6640 -22809
rect 5680 -22864 6640 -22826
rect 6698 -22826 6900 -22809
rect 7456 -22809 7472 -22792
rect 7902 -22792 8490 -22776
rect 7902 -22809 7918 -22792
rect 7456 -22826 7658 -22809
rect 6698 -22864 7658 -22826
rect 7716 -22826 7918 -22809
rect 8474 -22809 8490 -22792
rect 8920 -22792 9508 -22776
rect 8920 -22809 8936 -22792
rect 8474 -22826 8676 -22809
rect 7716 -22864 8676 -22826
rect 8734 -22826 8936 -22809
rect 9492 -22809 9508 -22792
rect 9938 -22792 10526 -22776
rect 9938 -22809 9954 -22792
rect 9492 -22826 9694 -22809
rect 8734 -22864 9694 -22826
rect 9752 -22826 9954 -22809
rect 10510 -22809 10526 -22792
rect 10956 -22792 11544 -22776
rect 10956 -22809 10972 -22792
rect 10510 -22826 10712 -22809
rect 9752 -22864 10712 -22826
rect 10770 -22826 10972 -22809
rect 11528 -22809 11544 -22792
rect 11974 -22792 12562 -22776
rect 11974 -22809 11990 -22792
rect 11528 -22826 11730 -22809
rect 10770 -22864 11730 -22826
rect 11788 -22826 11990 -22809
rect 12546 -22809 12562 -22792
rect 12992 -22792 13580 -22776
rect 12992 -22809 13008 -22792
rect 12546 -22826 12748 -22809
rect 11788 -22864 12748 -22826
rect 12806 -22826 13008 -22809
rect 13564 -22809 13580 -22792
rect 14010 -22792 14598 -22776
rect 14010 -22809 14026 -22792
rect 13564 -22826 13766 -22809
rect 12806 -22864 13766 -22826
rect 13824 -22826 14026 -22809
rect 14582 -22809 14598 -22792
rect 15028 -22792 15616 -22776
rect 15028 -22809 15044 -22792
rect 14582 -22826 14784 -22809
rect 13824 -22864 14784 -22826
rect 14842 -22826 15044 -22809
rect 15600 -22809 15616 -22792
rect 16046 -22792 16634 -22776
rect 16046 -22809 16062 -22792
rect 15600 -22826 15802 -22809
rect 14842 -22864 15802 -22826
rect 15860 -22826 16062 -22809
rect 16618 -22809 16634 -22792
rect 17064 -22792 17652 -22776
rect 17064 -22809 17080 -22792
rect 16618 -22826 16820 -22809
rect 15860 -22864 16820 -22826
rect 16878 -22826 17080 -22809
rect 17636 -22809 17652 -22792
rect 18082 -22792 18670 -22776
rect 18082 -22809 18098 -22792
rect 17636 -22826 17838 -22809
rect 16878 -22864 17838 -22826
rect 17896 -22826 18098 -22809
rect 18654 -22809 18670 -22792
rect 19100 -22792 19688 -22776
rect 19100 -22809 19116 -22792
rect 18654 -22826 18856 -22809
rect 17896 -22864 18856 -22826
rect 18914 -22826 19116 -22809
rect 19672 -22809 19688 -22792
rect 20118 -22792 20706 -22776
rect 20118 -22809 20134 -22792
rect 19672 -22826 19874 -22809
rect 18914 -22864 19874 -22826
rect 19932 -22826 20134 -22809
rect 20690 -22809 20706 -22792
rect 21136 -22792 21724 -22776
rect 21136 -22809 21152 -22792
rect 20690 -22826 20892 -22809
rect 19932 -22864 20892 -22826
rect 20950 -22826 21152 -22809
rect 21708 -22809 21724 -22792
rect 22154 -22792 22742 -22776
rect 22154 -22809 22170 -22792
rect 21708 -22826 21910 -22809
rect 20950 -22864 21910 -22826
rect 21968 -22826 22170 -22809
rect 22726 -22809 22742 -22792
rect 22726 -22826 22928 -22809
rect 21968 -22864 22928 -22826
rect -10462 -23124 -9502 -23086
rect -10462 -23141 -10260 -23124
rect -10276 -23158 -10260 -23141
rect -9704 -23141 -9502 -23124
rect -9444 -23124 -8484 -23086
rect -9444 -23141 -9242 -23124
rect -9704 -23158 -9688 -23141
rect -10276 -23174 -9688 -23158
rect -9258 -23158 -9242 -23141
rect -8686 -23141 -8484 -23124
rect -8426 -23124 -7466 -23086
rect -8426 -23141 -8224 -23124
rect -8686 -23158 -8670 -23141
rect -9258 -23174 -8670 -23158
rect -8240 -23158 -8224 -23141
rect -7668 -23141 -7466 -23124
rect -7408 -23124 -6448 -23086
rect -7408 -23141 -7206 -23124
rect -7668 -23158 -7652 -23141
rect -8240 -23174 -7652 -23158
rect -7222 -23158 -7206 -23141
rect -6650 -23141 -6448 -23124
rect -6390 -23124 -5430 -23086
rect -6390 -23141 -6188 -23124
rect -6650 -23158 -6634 -23141
rect -7222 -23174 -6634 -23158
rect -6204 -23158 -6188 -23141
rect -5632 -23141 -5430 -23124
rect -5372 -23124 -4412 -23086
rect -5372 -23141 -5170 -23124
rect -5632 -23158 -5616 -23141
rect -6204 -23174 -5616 -23158
rect -5186 -23158 -5170 -23141
rect -4614 -23141 -4412 -23124
rect -4354 -23124 -3394 -23086
rect -4354 -23141 -4152 -23124
rect -4614 -23158 -4598 -23141
rect -5186 -23174 -4598 -23158
rect -4168 -23158 -4152 -23141
rect -3596 -23141 -3394 -23124
rect -3336 -23124 -2376 -23086
rect -3336 -23141 -3134 -23124
rect -3596 -23158 -3580 -23141
rect -4168 -23174 -3580 -23158
rect -3150 -23158 -3134 -23141
rect -2578 -23141 -2376 -23124
rect -2318 -23124 -1358 -23086
rect -2318 -23141 -2116 -23124
rect -2578 -23158 -2562 -23141
rect -3150 -23174 -2562 -23158
rect -2132 -23158 -2116 -23141
rect -1560 -23141 -1358 -23124
rect -1300 -23124 -340 -23086
rect -1300 -23141 -1098 -23124
rect -1560 -23158 -1544 -23141
rect -2132 -23174 -1544 -23158
rect -1114 -23158 -1098 -23141
rect -542 -23141 -340 -23124
rect -282 -23124 678 -23086
rect -282 -23141 -80 -23124
rect -542 -23158 -526 -23141
rect -1114 -23174 -526 -23158
rect -96 -23158 -80 -23141
rect 476 -23141 678 -23124
rect 476 -23158 492 -23141
rect -96 -23174 492 -23158
rect 2626 -23502 3586 -23464
rect -10276 -23526 -9688 -23510
rect -10276 -23543 -10260 -23526
rect -10462 -23560 -10260 -23543
rect -9704 -23543 -9688 -23526
rect -9258 -23526 -8670 -23510
rect -9258 -23543 -9242 -23526
rect -9704 -23560 -9502 -23543
rect -10462 -23598 -9502 -23560
rect -9444 -23560 -9242 -23543
rect -8686 -23543 -8670 -23526
rect -8240 -23526 -7652 -23510
rect -8240 -23543 -8224 -23526
rect -8686 -23560 -8484 -23543
rect -9444 -23598 -8484 -23560
rect -8426 -23560 -8224 -23543
rect -7668 -23543 -7652 -23526
rect -7222 -23526 -6634 -23510
rect -7222 -23543 -7206 -23526
rect -7668 -23560 -7466 -23543
rect -8426 -23598 -7466 -23560
rect -7408 -23560 -7206 -23543
rect -6650 -23543 -6634 -23526
rect -6204 -23526 -5616 -23510
rect -6204 -23543 -6188 -23526
rect -6650 -23560 -6448 -23543
rect -7408 -23598 -6448 -23560
rect -6390 -23560 -6188 -23543
rect -5632 -23543 -5616 -23526
rect -5186 -23526 -4598 -23510
rect -5186 -23543 -5170 -23526
rect -5632 -23560 -5430 -23543
rect -6390 -23598 -5430 -23560
rect -5372 -23560 -5170 -23543
rect -4614 -23543 -4598 -23526
rect -4168 -23526 -3580 -23510
rect -4168 -23543 -4152 -23526
rect -4614 -23560 -4412 -23543
rect -5372 -23598 -4412 -23560
rect -4354 -23560 -4152 -23543
rect -3596 -23543 -3580 -23526
rect -3150 -23526 -2562 -23510
rect -3150 -23543 -3134 -23526
rect -3596 -23560 -3394 -23543
rect -4354 -23598 -3394 -23560
rect -3336 -23560 -3134 -23543
rect -2578 -23543 -2562 -23526
rect -2132 -23526 -1544 -23510
rect -2132 -23543 -2116 -23526
rect -2578 -23560 -2376 -23543
rect -3336 -23598 -2376 -23560
rect -2318 -23560 -2116 -23543
rect -1560 -23543 -1544 -23526
rect -1114 -23526 -526 -23510
rect -1114 -23543 -1098 -23526
rect -1560 -23560 -1358 -23543
rect -2318 -23598 -1358 -23560
rect -1300 -23560 -1098 -23543
rect -542 -23543 -526 -23526
rect -96 -23526 492 -23510
rect 2626 -23519 2828 -23502
rect -96 -23543 -80 -23526
rect -542 -23560 -340 -23543
rect -1300 -23598 -340 -23560
rect -282 -23560 -80 -23543
rect 476 -23543 492 -23526
rect 2812 -23536 2828 -23519
rect 3384 -23519 3586 -23502
rect 3644 -23502 4604 -23464
rect 3644 -23519 3846 -23502
rect 3384 -23536 3400 -23519
rect 476 -23560 678 -23543
rect 2812 -23552 3400 -23536
rect 3830 -23536 3846 -23519
rect 4402 -23519 4604 -23502
rect 4662 -23502 5622 -23464
rect 4662 -23519 4864 -23502
rect 4402 -23536 4418 -23519
rect 3830 -23552 4418 -23536
rect 4848 -23536 4864 -23519
rect 5420 -23519 5622 -23502
rect 5680 -23502 6640 -23464
rect 5680 -23519 5882 -23502
rect 5420 -23536 5436 -23519
rect 4848 -23552 5436 -23536
rect 5866 -23536 5882 -23519
rect 6438 -23519 6640 -23502
rect 6698 -23502 7658 -23464
rect 6698 -23519 6900 -23502
rect 6438 -23536 6454 -23519
rect 5866 -23552 6454 -23536
rect 6884 -23536 6900 -23519
rect 7456 -23519 7658 -23502
rect 7716 -23502 8676 -23464
rect 7716 -23519 7918 -23502
rect 7456 -23536 7472 -23519
rect 6884 -23552 7472 -23536
rect 7902 -23536 7918 -23519
rect 8474 -23519 8676 -23502
rect 8734 -23502 9694 -23464
rect 8734 -23519 8936 -23502
rect 8474 -23536 8490 -23519
rect 7902 -23552 8490 -23536
rect 8920 -23536 8936 -23519
rect 9492 -23519 9694 -23502
rect 9752 -23502 10712 -23464
rect 9752 -23519 9954 -23502
rect 9492 -23536 9508 -23519
rect 8920 -23552 9508 -23536
rect 9938 -23536 9954 -23519
rect 10510 -23519 10712 -23502
rect 10770 -23502 11730 -23464
rect 10770 -23519 10972 -23502
rect 10510 -23536 10526 -23519
rect 9938 -23552 10526 -23536
rect 10956 -23536 10972 -23519
rect 11528 -23519 11730 -23502
rect 11788 -23502 12748 -23464
rect 11788 -23519 11990 -23502
rect 11528 -23536 11544 -23519
rect 10956 -23552 11544 -23536
rect 11974 -23536 11990 -23519
rect 12546 -23519 12748 -23502
rect 12806 -23502 13766 -23464
rect 12806 -23519 13008 -23502
rect 12546 -23536 12562 -23519
rect 11974 -23552 12562 -23536
rect 12992 -23536 13008 -23519
rect 13564 -23519 13766 -23502
rect 13824 -23502 14784 -23464
rect 13824 -23519 14026 -23502
rect 13564 -23536 13580 -23519
rect 12992 -23552 13580 -23536
rect 14010 -23536 14026 -23519
rect 14582 -23519 14784 -23502
rect 14842 -23502 15802 -23464
rect 14842 -23519 15044 -23502
rect 14582 -23536 14598 -23519
rect 14010 -23552 14598 -23536
rect 15028 -23536 15044 -23519
rect 15600 -23519 15802 -23502
rect 15860 -23502 16820 -23464
rect 15860 -23519 16062 -23502
rect 15600 -23536 15616 -23519
rect 15028 -23552 15616 -23536
rect 16046 -23536 16062 -23519
rect 16618 -23519 16820 -23502
rect 16878 -23502 17838 -23464
rect 16878 -23519 17080 -23502
rect 16618 -23536 16634 -23519
rect 16046 -23552 16634 -23536
rect 17064 -23536 17080 -23519
rect 17636 -23519 17838 -23502
rect 17896 -23502 18856 -23464
rect 17896 -23519 18098 -23502
rect 17636 -23536 17652 -23519
rect 17064 -23552 17652 -23536
rect 18082 -23536 18098 -23519
rect 18654 -23519 18856 -23502
rect 18914 -23502 19874 -23464
rect 18914 -23519 19116 -23502
rect 18654 -23536 18670 -23519
rect 18082 -23552 18670 -23536
rect 19100 -23536 19116 -23519
rect 19672 -23519 19874 -23502
rect 19932 -23502 20892 -23464
rect 19932 -23519 20134 -23502
rect 19672 -23536 19688 -23519
rect 19100 -23552 19688 -23536
rect 20118 -23536 20134 -23519
rect 20690 -23519 20892 -23502
rect 20950 -23502 21910 -23464
rect 20950 -23519 21152 -23502
rect 20690 -23536 20706 -23519
rect 20118 -23552 20706 -23536
rect 21136 -23536 21152 -23519
rect 21708 -23519 21910 -23502
rect 21968 -23502 22928 -23464
rect 21968 -23519 22170 -23502
rect 21708 -23536 21724 -23519
rect 21136 -23552 21724 -23536
rect 22154 -23536 22170 -23519
rect 22726 -23519 22928 -23502
rect 22726 -23536 22742 -23519
rect 22154 -23552 22742 -23536
rect -282 -23598 678 -23560
rect 2812 -24026 3400 -24010
rect 2812 -24043 2828 -24026
rect 2626 -24060 2828 -24043
rect 3384 -24043 3400 -24026
rect 3830 -24026 4418 -24010
rect 3830 -24043 3846 -24026
rect 3384 -24060 3586 -24043
rect 2626 -24098 3586 -24060
rect 3644 -24060 3846 -24043
rect 4402 -24043 4418 -24026
rect 4848 -24026 5436 -24010
rect 4848 -24043 4864 -24026
rect 4402 -24060 4604 -24043
rect 3644 -24098 4604 -24060
rect 4662 -24060 4864 -24043
rect 5420 -24043 5436 -24026
rect 5866 -24026 6454 -24010
rect 5866 -24043 5882 -24026
rect 5420 -24060 5622 -24043
rect 4662 -24098 5622 -24060
rect 5680 -24060 5882 -24043
rect 6438 -24043 6454 -24026
rect 6884 -24026 7472 -24010
rect 6884 -24043 6900 -24026
rect 6438 -24060 6640 -24043
rect 5680 -24098 6640 -24060
rect 6698 -24060 6900 -24043
rect 7456 -24043 7472 -24026
rect 7902 -24026 8490 -24010
rect 7902 -24043 7918 -24026
rect 7456 -24060 7658 -24043
rect 6698 -24098 7658 -24060
rect 7716 -24060 7918 -24043
rect 8474 -24043 8490 -24026
rect 8920 -24026 9508 -24010
rect 8920 -24043 8936 -24026
rect 8474 -24060 8676 -24043
rect 7716 -24098 8676 -24060
rect 8734 -24060 8936 -24043
rect 9492 -24043 9508 -24026
rect 9938 -24026 10526 -24010
rect 9938 -24043 9954 -24026
rect 9492 -24060 9694 -24043
rect 8734 -24098 9694 -24060
rect 9752 -24060 9954 -24043
rect 10510 -24043 10526 -24026
rect 10956 -24026 11544 -24010
rect 10956 -24043 10972 -24026
rect 10510 -24060 10712 -24043
rect 9752 -24098 10712 -24060
rect 10770 -24060 10972 -24043
rect 11528 -24043 11544 -24026
rect 11974 -24026 12562 -24010
rect 11974 -24043 11990 -24026
rect 11528 -24060 11730 -24043
rect 10770 -24098 11730 -24060
rect 11788 -24060 11990 -24043
rect 12546 -24043 12562 -24026
rect 12992 -24026 13580 -24010
rect 12992 -24043 13008 -24026
rect 12546 -24060 12748 -24043
rect 11788 -24098 12748 -24060
rect 12806 -24060 13008 -24043
rect 13564 -24043 13580 -24026
rect 14010 -24026 14598 -24010
rect 14010 -24043 14026 -24026
rect 13564 -24060 13766 -24043
rect 12806 -24098 13766 -24060
rect 13824 -24060 14026 -24043
rect 14582 -24043 14598 -24026
rect 15028 -24026 15616 -24010
rect 15028 -24043 15044 -24026
rect 14582 -24060 14784 -24043
rect 13824 -24098 14784 -24060
rect 14842 -24060 15044 -24043
rect 15600 -24043 15616 -24026
rect 16046 -24026 16634 -24010
rect 16046 -24043 16062 -24026
rect 15600 -24060 15802 -24043
rect 14842 -24098 15802 -24060
rect 15860 -24060 16062 -24043
rect 16618 -24043 16634 -24026
rect 17064 -24026 17652 -24010
rect 17064 -24043 17080 -24026
rect 16618 -24060 16820 -24043
rect 15860 -24098 16820 -24060
rect 16878 -24060 17080 -24043
rect 17636 -24043 17652 -24026
rect 18082 -24026 18670 -24010
rect 18082 -24043 18098 -24026
rect 17636 -24060 17838 -24043
rect 16878 -24098 17838 -24060
rect 17896 -24060 18098 -24043
rect 18654 -24043 18670 -24026
rect 19100 -24026 19688 -24010
rect 19100 -24043 19116 -24026
rect 18654 -24060 18856 -24043
rect 17896 -24098 18856 -24060
rect 18914 -24060 19116 -24043
rect 19672 -24043 19688 -24026
rect 20118 -24026 20706 -24010
rect 20118 -24043 20134 -24026
rect 19672 -24060 19874 -24043
rect 18914 -24098 19874 -24060
rect 19932 -24060 20134 -24043
rect 20690 -24043 20706 -24026
rect 21136 -24026 21724 -24010
rect 21136 -24043 21152 -24026
rect 20690 -24060 20892 -24043
rect 19932 -24098 20892 -24060
rect 20950 -24060 21152 -24043
rect 21708 -24043 21724 -24026
rect 22154 -24026 22742 -24010
rect 22154 -24043 22170 -24026
rect 21708 -24060 21910 -24043
rect 20950 -24098 21910 -24060
rect 21968 -24060 22170 -24043
rect 22726 -24043 22742 -24026
rect 22726 -24060 22928 -24043
rect 21968 -24098 22928 -24060
rect -10462 -24236 -9502 -24198
rect -10462 -24253 -10260 -24236
rect -10276 -24270 -10260 -24253
rect -9704 -24253 -9502 -24236
rect -9444 -24236 -8484 -24198
rect -9444 -24253 -9242 -24236
rect -9704 -24270 -9688 -24253
rect -10276 -24286 -9688 -24270
rect -9258 -24270 -9242 -24253
rect -8686 -24253 -8484 -24236
rect -8426 -24236 -7466 -24198
rect -8426 -24253 -8224 -24236
rect -8686 -24270 -8670 -24253
rect -9258 -24286 -8670 -24270
rect -8240 -24270 -8224 -24253
rect -7668 -24253 -7466 -24236
rect -7408 -24236 -6448 -24198
rect -7408 -24253 -7206 -24236
rect -7668 -24270 -7652 -24253
rect -8240 -24286 -7652 -24270
rect -7222 -24270 -7206 -24253
rect -6650 -24253 -6448 -24236
rect -6390 -24236 -5430 -24198
rect -6390 -24253 -6188 -24236
rect -6650 -24270 -6634 -24253
rect -7222 -24286 -6634 -24270
rect -6204 -24270 -6188 -24253
rect -5632 -24253 -5430 -24236
rect -5372 -24236 -4412 -24198
rect -5372 -24253 -5170 -24236
rect -5632 -24270 -5616 -24253
rect -6204 -24286 -5616 -24270
rect -5186 -24270 -5170 -24253
rect -4614 -24253 -4412 -24236
rect -4354 -24236 -3394 -24198
rect -4354 -24253 -4152 -24236
rect -4614 -24270 -4598 -24253
rect -5186 -24286 -4598 -24270
rect -4168 -24270 -4152 -24253
rect -3596 -24253 -3394 -24236
rect -3336 -24236 -2376 -24198
rect -3336 -24253 -3134 -24236
rect -3596 -24270 -3580 -24253
rect -4168 -24286 -3580 -24270
rect -3150 -24270 -3134 -24253
rect -2578 -24253 -2376 -24236
rect -2318 -24236 -1358 -24198
rect -2318 -24253 -2116 -24236
rect -2578 -24270 -2562 -24253
rect -3150 -24286 -2562 -24270
rect -2132 -24270 -2116 -24253
rect -1560 -24253 -1358 -24236
rect -1300 -24236 -340 -24198
rect -1300 -24253 -1098 -24236
rect -1560 -24270 -1544 -24253
rect -2132 -24286 -1544 -24270
rect -1114 -24270 -1098 -24253
rect -542 -24253 -340 -24236
rect -282 -24236 678 -24198
rect -282 -24253 -80 -24236
rect -542 -24270 -526 -24253
rect -1114 -24286 -526 -24270
rect -96 -24270 -80 -24253
rect 476 -24253 678 -24236
rect 476 -24270 492 -24253
rect -96 -24286 492 -24270
rect 2626 -24736 3586 -24698
rect 2626 -24753 2828 -24736
rect 2812 -24770 2828 -24753
rect 3384 -24753 3586 -24736
rect 3644 -24736 4604 -24698
rect 3644 -24753 3846 -24736
rect 3384 -24770 3400 -24753
rect 2812 -24786 3400 -24770
rect 3830 -24770 3846 -24753
rect 4402 -24753 4604 -24736
rect 4662 -24736 5622 -24698
rect 4662 -24753 4864 -24736
rect 4402 -24770 4418 -24753
rect 3830 -24786 4418 -24770
rect 4848 -24770 4864 -24753
rect 5420 -24753 5622 -24736
rect 5680 -24736 6640 -24698
rect 5680 -24753 5882 -24736
rect 5420 -24770 5436 -24753
rect 4848 -24786 5436 -24770
rect 5866 -24770 5882 -24753
rect 6438 -24753 6640 -24736
rect 6698 -24736 7658 -24698
rect 6698 -24753 6900 -24736
rect 6438 -24770 6454 -24753
rect 5866 -24786 6454 -24770
rect 6884 -24770 6900 -24753
rect 7456 -24753 7658 -24736
rect 7716 -24736 8676 -24698
rect 7716 -24753 7918 -24736
rect 7456 -24770 7472 -24753
rect 6884 -24786 7472 -24770
rect 7902 -24770 7918 -24753
rect 8474 -24753 8676 -24736
rect 8734 -24736 9694 -24698
rect 8734 -24753 8936 -24736
rect 8474 -24770 8490 -24753
rect 7902 -24786 8490 -24770
rect 8920 -24770 8936 -24753
rect 9492 -24753 9694 -24736
rect 9752 -24736 10712 -24698
rect 9752 -24753 9954 -24736
rect 9492 -24770 9508 -24753
rect 8920 -24786 9508 -24770
rect 9938 -24770 9954 -24753
rect 10510 -24753 10712 -24736
rect 10770 -24736 11730 -24698
rect 10770 -24753 10972 -24736
rect 10510 -24770 10526 -24753
rect 9938 -24786 10526 -24770
rect 10956 -24770 10972 -24753
rect 11528 -24753 11730 -24736
rect 11788 -24736 12748 -24698
rect 11788 -24753 11990 -24736
rect 11528 -24770 11544 -24753
rect 10956 -24786 11544 -24770
rect 11974 -24770 11990 -24753
rect 12546 -24753 12748 -24736
rect 12806 -24736 13766 -24698
rect 12806 -24753 13008 -24736
rect 12546 -24770 12562 -24753
rect 11974 -24786 12562 -24770
rect 12992 -24770 13008 -24753
rect 13564 -24753 13766 -24736
rect 13824 -24736 14784 -24698
rect 13824 -24753 14026 -24736
rect 13564 -24770 13580 -24753
rect 12992 -24786 13580 -24770
rect 14010 -24770 14026 -24753
rect 14582 -24753 14784 -24736
rect 14842 -24736 15802 -24698
rect 14842 -24753 15044 -24736
rect 14582 -24770 14598 -24753
rect 14010 -24786 14598 -24770
rect 15028 -24770 15044 -24753
rect 15600 -24753 15802 -24736
rect 15860 -24736 16820 -24698
rect 15860 -24753 16062 -24736
rect 15600 -24770 15616 -24753
rect 15028 -24786 15616 -24770
rect 16046 -24770 16062 -24753
rect 16618 -24753 16820 -24736
rect 16878 -24736 17838 -24698
rect 16878 -24753 17080 -24736
rect 16618 -24770 16634 -24753
rect 16046 -24786 16634 -24770
rect 17064 -24770 17080 -24753
rect 17636 -24753 17838 -24736
rect 17896 -24736 18856 -24698
rect 17896 -24753 18098 -24736
rect 17636 -24770 17652 -24753
rect 17064 -24786 17652 -24770
rect 18082 -24770 18098 -24753
rect 18654 -24753 18856 -24736
rect 18914 -24736 19874 -24698
rect 18914 -24753 19116 -24736
rect 18654 -24770 18670 -24753
rect 18082 -24786 18670 -24770
rect 19100 -24770 19116 -24753
rect 19672 -24753 19874 -24736
rect 19932 -24736 20892 -24698
rect 19932 -24753 20134 -24736
rect 19672 -24770 19688 -24753
rect 19100 -24786 19688 -24770
rect 20118 -24770 20134 -24753
rect 20690 -24753 20892 -24736
rect 20950 -24736 21910 -24698
rect 20950 -24753 21152 -24736
rect 20690 -24770 20706 -24753
rect 20118 -24786 20706 -24770
rect 21136 -24770 21152 -24753
rect 21708 -24753 21910 -24736
rect 21968 -24736 22928 -24698
rect 21968 -24753 22170 -24736
rect 21708 -24770 21724 -24753
rect 21136 -24786 21724 -24770
rect 22154 -24770 22170 -24753
rect 22726 -24753 22928 -24736
rect 22726 -24770 22742 -24753
rect 22154 -24786 22742 -24770
rect -9818 -25068 -9230 -25052
rect -9818 -25085 -9802 -25068
rect -10004 -25102 -9802 -25085
rect -9246 -25085 -9230 -25068
rect -8800 -25068 -8212 -25052
rect -8800 -25085 -8784 -25068
rect -9246 -25102 -9044 -25085
rect -10004 -25140 -9044 -25102
rect -8986 -25102 -8784 -25085
rect -8228 -25085 -8212 -25068
rect -7782 -25068 -7194 -25052
rect -7782 -25085 -7766 -25068
rect -8228 -25102 -8026 -25085
rect -8986 -25140 -8026 -25102
rect -7968 -25102 -7766 -25085
rect -7210 -25085 -7194 -25068
rect -6764 -25068 -6176 -25052
rect -6764 -25085 -6748 -25068
rect -7210 -25102 -7008 -25085
rect -7968 -25140 -7008 -25102
rect -6950 -25102 -6748 -25085
rect -6192 -25085 -6176 -25068
rect -5746 -25068 -5158 -25052
rect -5746 -25085 -5730 -25068
rect -6192 -25102 -5990 -25085
rect -6950 -25140 -5990 -25102
rect -5932 -25102 -5730 -25085
rect -5174 -25085 -5158 -25068
rect -4728 -25068 -4140 -25052
rect -4728 -25085 -4712 -25068
rect -5174 -25102 -4972 -25085
rect -5932 -25140 -4972 -25102
rect -4914 -25102 -4712 -25085
rect -4156 -25085 -4140 -25068
rect -3710 -25068 -3122 -25052
rect -3710 -25085 -3694 -25068
rect -4156 -25102 -3954 -25085
rect -4914 -25140 -3954 -25102
rect -3896 -25102 -3694 -25085
rect -3138 -25085 -3122 -25068
rect -2692 -25068 -2104 -25052
rect -2692 -25085 -2676 -25068
rect -3138 -25102 -2936 -25085
rect -3896 -25140 -2936 -25102
rect -2878 -25102 -2676 -25085
rect -2120 -25085 -2104 -25068
rect -1674 -25068 -1086 -25052
rect -1674 -25085 -1658 -25068
rect -2120 -25102 -1918 -25085
rect -2878 -25140 -1918 -25102
rect -1860 -25102 -1658 -25085
rect -1102 -25085 -1086 -25068
rect -656 -25068 -68 -25052
rect -656 -25085 -640 -25068
rect -1102 -25102 -900 -25085
rect -1860 -25140 -900 -25102
rect -842 -25102 -640 -25085
rect -84 -25085 -68 -25068
rect -84 -25102 118 -25085
rect -842 -25140 118 -25102
rect 2812 -25258 3400 -25242
rect 2812 -25275 2828 -25258
rect 2626 -25292 2828 -25275
rect 3384 -25275 3400 -25258
rect 3830 -25258 4418 -25242
rect 3830 -25275 3846 -25258
rect 3384 -25292 3586 -25275
rect 2626 -25330 3586 -25292
rect 3644 -25292 3846 -25275
rect 4402 -25275 4418 -25258
rect 4848 -25258 5436 -25242
rect 4848 -25275 4864 -25258
rect 4402 -25292 4604 -25275
rect 3644 -25330 4604 -25292
rect 4662 -25292 4864 -25275
rect 5420 -25275 5436 -25258
rect 5866 -25258 6454 -25242
rect 5866 -25275 5882 -25258
rect 5420 -25292 5622 -25275
rect 4662 -25330 5622 -25292
rect 5680 -25292 5882 -25275
rect 6438 -25275 6454 -25258
rect 6884 -25258 7472 -25242
rect 6884 -25275 6900 -25258
rect 6438 -25292 6640 -25275
rect 5680 -25330 6640 -25292
rect 6698 -25292 6900 -25275
rect 7456 -25275 7472 -25258
rect 7902 -25258 8490 -25242
rect 7902 -25275 7918 -25258
rect 7456 -25292 7658 -25275
rect 6698 -25330 7658 -25292
rect 7716 -25292 7918 -25275
rect 8474 -25275 8490 -25258
rect 8920 -25258 9508 -25242
rect 8920 -25275 8936 -25258
rect 8474 -25292 8676 -25275
rect 7716 -25330 8676 -25292
rect 8734 -25292 8936 -25275
rect 9492 -25275 9508 -25258
rect 9938 -25258 10526 -25242
rect 9938 -25275 9954 -25258
rect 9492 -25292 9694 -25275
rect 8734 -25330 9694 -25292
rect 9752 -25292 9954 -25275
rect 10510 -25275 10526 -25258
rect 10956 -25258 11544 -25242
rect 10956 -25275 10972 -25258
rect 10510 -25292 10712 -25275
rect 9752 -25330 10712 -25292
rect 10770 -25292 10972 -25275
rect 11528 -25275 11544 -25258
rect 11974 -25258 12562 -25242
rect 11974 -25275 11990 -25258
rect 11528 -25292 11730 -25275
rect 10770 -25330 11730 -25292
rect 11788 -25292 11990 -25275
rect 12546 -25275 12562 -25258
rect 12992 -25258 13580 -25242
rect 12992 -25275 13008 -25258
rect 12546 -25292 12748 -25275
rect 11788 -25330 12748 -25292
rect 12806 -25292 13008 -25275
rect 13564 -25275 13580 -25258
rect 14010 -25258 14598 -25242
rect 14010 -25275 14026 -25258
rect 13564 -25292 13766 -25275
rect 12806 -25330 13766 -25292
rect 13824 -25292 14026 -25275
rect 14582 -25275 14598 -25258
rect 15028 -25258 15616 -25242
rect 15028 -25275 15044 -25258
rect 14582 -25292 14784 -25275
rect 13824 -25330 14784 -25292
rect 14842 -25292 15044 -25275
rect 15600 -25275 15616 -25258
rect 16046 -25258 16634 -25242
rect 16046 -25275 16062 -25258
rect 15600 -25292 15802 -25275
rect 14842 -25330 15802 -25292
rect 15860 -25292 16062 -25275
rect 16618 -25275 16634 -25258
rect 17064 -25258 17652 -25242
rect 17064 -25275 17080 -25258
rect 16618 -25292 16820 -25275
rect 15860 -25330 16820 -25292
rect 16878 -25292 17080 -25275
rect 17636 -25275 17652 -25258
rect 18082 -25258 18670 -25242
rect 18082 -25275 18098 -25258
rect 17636 -25292 17838 -25275
rect 16878 -25330 17838 -25292
rect 17896 -25292 18098 -25275
rect 18654 -25275 18670 -25258
rect 19100 -25258 19688 -25242
rect 19100 -25275 19116 -25258
rect 18654 -25292 18856 -25275
rect 17896 -25330 18856 -25292
rect 18914 -25292 19116 -25275
rect 19672 -25275 19688 -25258
rect 20118 -25258 20706 -25242
rect 20118 -25275 20134 -25258
rect 19672 -25292 19874 -25275
rect 18914 -25330 19874 -25292
rect 19932 -25292 20134 -25275
rect 20690 -25275 20706 -25258
rect 21136 -25258 21724 -25242
rect 21136 -25275 21152 -25258
rect 20690 -25292 20892 -25275
rect 19932 -25330 20892 -25292
rect 20950 -25292 21152 -25275
rect 21708 -25275 21724 -25258
rect 22154 -25258 22742 -25242
rect 22154 -25275 22170 -25258
rect 21708 -25292 21910 -25275
rect 20950 -25330 21910 -25292
rect 21968 -25292 22170 -25275
rect 22726 -25275 22742 -25258
rect 22726 -25292 22928 -25275
rect 21968 -25330 22928 -25292
rect -10004 -25778 -9044 -25740
rect -10004 -25795 -9802 -25778
rect -9818 -25812 -9802 -25795
rect -9246 -25795 -9044 -25778
rect -8986 -25778 -8026 -25740
rect -8986 -25795 -8784 -25778
rect -9246 -25812 -9230 -25795
rect -9818 -25828 -9230 -25812
rect -8800 -25812 -8784 -25795
rect -8228 -25795 -8026 -25778
rect -7968 -25778 -7008 -25740
rect -7968 -25795 -7766 -25778
rect -8228 -25812 -8212 -25795
rect -8800 -25828 -8212 -25812
rect -7782 -25812 -7766 -25795
rect -7210 -25795 -7008 -25778
rect -6950 -25778 -5990 -25740
rect -6950 -25795 -6748 -25778
rect -7210 -25812 -7194 -25795
rect -7782 -25828 -7194 -25812
rect -6764 -25812 -6748 -25795
rect -6192 -25795 -5990 -25778
rect -5932 -25778 -4972 -25740
rect -5932 -25795 -5730 -25778
rect -6192 -25812 -6176 -25795
rect -6764 -25828 -6176 -25812
rect -5746 -25812 -5730 -25795
rect -5174 -25795 -4972 -25778
rect -4914 -25778 -3954 -25740
rect -4914 -25795 -4712 -25778
rect -5174 -25812 -5158 -25795
rect -5746 -25828 -5158 -25812
rect -4728 -25812 -4712 -25795
rect -4156 -25795 -3954 -25778
rect -3896 -25778 -2936 -25740
rect -3896 -25795 -3694 -25778
rect -4156 -25812 -4140 -25795
rect -4728 -25828 -4140 -25812
rect -3710 -25812 -3694 -25795
rect -3138 -25795 -2936 -25778
rect -2878 -25778 -1918 -25740
rect -2878 -25795 -2676 -25778
rect -3138 -25812 -3122 -25795
rect -3710 -25828 -3122 -25812
rect -2692 -25812 -2676 -25795
rect -2120 -25795 -1918 -25778
rect -1860 -25778 -900 -25740
rect -1860 -25795 -1658 -25778
rect -2120 -25812 -2104 -25795
rect -2692 -25828 -2104 -25812
rect -1674 -25812 -1658 -25795
rect -1102 -25795 -900 -25778
rect -842 -25778 118 -25740
rect -842 -25795 -640 -25778
rect -1102 -25812 -1086 -25795
rect -1674 -25828 -1086 -25812
rect -656 -25812 -640 -25795
rect -84 -25795 118 -25778
rect -84 -25812 -68 -25795
rect -656 -25828 -68 -25812
rect 2626 -25968 3586 -25930
rect 2626 -25985 2828 -25968
rect 2812 -26002 2828 -25985
rect 3384 -25985 3586 -25968
rect 3644 -25968 4604 -25930
rect 3644 -25985 3846 -25968
rect 3384 -26002 3400 -25985
rect 2812 -26018 3400 -26002
rect 3830 -26002 3846 -25985
rect 4402 -25985 4604 -25968
rect 4662 -25968 5622 -25930
rect 4662 -25985 4864 -25968
rect 4402 -26002 4418 -25985
rect 3830 -26018 4418 -26002
rect 4848 -26002 4864 -25985
rect 5420 -25985 5622 -25968
rect 5680 -25968 6640 -25930
rect 5680 -25985 5882 -25968
rect 5420 -26002 5436 -25985
rect 4848 -26018 5436 -26002
rect 5866 -26002 5882 -25985
rect 6438 -25985 6640 -25968
rect 6698 -25968 7658 -25930
rect 6698 -25985 6900 -25968
rect 6438 -26002 6454 -25985
rect 5866 -26018 6454 -26002
rect 6884 -26002 6900 -25985
rect 7456 -25985 7658 -25968
rect 7716 -25968 8676 -25930
rect 7716 -25985 7918 -25968
rect 7456 -26002 7472 -25985
rect 6884 -26018 7472 -26002
rect 7902 -26002 7918 -25985
rect 8474 -25985 8676 -25968
rect 8734 -25968 9694 -25930
rect 8734 -25985 8936 -25968
rect 8474 -26002 8490 -25985
rect 7902 -26018 8490 -26002
rect 8920 -26002 8936 -25985
rect 9492 -25985 9694 -25968
rect 9752 -25968 10712 -25930
rect 9752 -25985 9954 -25968
rect 9492 -26002 9508 -25985
rect 8920 -26018 9508 -26002
rect 9938 -26002 9954 -25985
rect 10510 -25985 10712 -25968
rect 10770 -25968 11730 -25930
rect 10770 -25985 10972 -25968
rect 10510 -26002 10526 -25985
rect 9938 -26018 10526 -26002
rect 10956 -26002 10972 -25985
rect 11528 -25985 11730 -25968
rect 11788 -25968 12748 -25930
rect 11788 -25985 11990 -25968
rect 11528 -26002 11544 -25985
rect 10956 -26018 11544 -26002
rect 11974 -26002 11990 -25985
rect 12546 -25985 12748 -25968
rect 12806 -25968 13766 -25930
rect 12806 -25985 13008 -25968
rect 12546 -26002 12562 -25985
rect 11974 -26018 12562 -26002
rect 12992 -26002 13008 -25985
rect 13564 -25985 13766 -25968
rect 13824 -25968 14784 -25930
rect 13824 -25985 14026 -25968
rect 13564 -26002 13580 -25985
rect 12992 -26018 13580 -26002
rect 14010 -26002 14026 -25985
rect 14582 -25985 14784 -25968
rect 14842 -25968 15802 -25930
rect 14842 -25985 15044 -25968
rect 14582 -26002 14598 -25985
rect 14010 -26018 14598 -26002
rect 15028 -26002 15044 -25985
rect 15600 -25985 15802 -25968
rect 15860 -25968 16820 -25930
rect 15860 -25985 16062 -25968
rect 15600 -26002 15616 -25985
rect 15028 -26018 15616 -26002
rect 16046 -26002 16062 -25985
rect 16618 -25985 16820 -25968
rect 16878 -25968 17838 -25930
rect 16878 -25985 17080 -25968
rect 16618 -26002 16634 -25985
rect 16046 -26018 16634 -26002
rect 17064 -26002 17080 -25985
rect 17636 -25985 17838 -25968
rect 17896 -25968 18856 -25930
rect 17896 -25985 18098 -25968
rect 17636 -26002 17652 -25985
rect 17064 -26018 17652 -26002
rect 18082 -26002 18098 -25985
rect 18654 -25985 18856 -25968
rect 18914 -25968 19874 -25930
rect 18914 -25985 19116 -25968
rect 18654 -26002 18670 -25985
rect 18082 -26018 18670 -26002
rect 19100 -26002 19116 -25985
rect 19672 -25985 19874 -25968
rect 19932 -25968 20892 -25930
rect 19932 -25985 20134 -25968
rect 19672 -26002 19688 -25985
rect 19100 -26018 19688 -26002
rect 20118 -26002 20134 -25985
rect 20690 -25985 20892 -25968
rect 20950 -25968 21910 -25930
rect 20950 -25985 21152 -25968
rect 20690 -26002 20706 -25985
rect 20118 -26018 20706 -26002
rect 21136 -26002 21152 -25985
rect 21708 -25985 21910 -25968
rect 21968 -25968 22928 -25930
rect 21968 -25985 22170 -25968
rect 21708 -26002 21724 -25985
rect 21136 -26018 21724 -26002
rect 22154 -26002 22170 -25985
rect 22726 -25985 22928 -25968
rect 22726 -26002 22742 -25985
rect 22154 -26018 22742 -26002
<< polycont >>
rect 6736 1521 7292 1555
rect 7754 1521 8310 1555
rect 8772 1521 9328 1555
rect 9790 1521 10346 1555
rect 10808 1521 11364 1555
rect 11826 1521 12382 1555
rect 12844 1521 13400 1555
rect 13862 1521 14418 1555
rect 14880 1521 15436 1555
rect 15898 1521 16454 1555
rect 16916 1521 17472 1555
rect 17934 1521 18490 1555
rect 18952 1521 19508 1555
rect 19970 1521 20526 1555
rect 20988 1521 21544 1555
rect 22006 1521 22562 1555
rect 6736 793 7292 827
rect 7754 793 8310 827
rect 8772 793 9328 827
rect 9790 793 10346 827
rect 10808 793 11364 827
rect 11826 793 12382 827
rect 12844 793 13400 827
rect 13862 793 14418 827
rect 14880 793 15436 827
rect 15898 793 16454 827
rect 16916 793 17472 827
rect 17934 793 18490 827
rect 18952 793 19508 827
rect 19970 793 20526 827
rect 20988 793 21544 827
rect 22006 793 22562 827
rect 6736 385 7292 419
rect 7754 385 8310 419
rect 8772 385 9328 419
rect 9790 385 10346 419
rect 10808 385 11364 419
rect 11826 385 12382 419
rect 12844 385 13400 419
rect 13862 385 14418 419
rect 14880 385 15436 419
rect 15898 385 16454 419
rect 16916 385 17472 419
rect 17934 385 18490 419
rect 18952 385 19508 419
rect 19970 385 20526 419
rect 20988 385 21544 419
rect 22006 385 22562 419
rect 6736 -343 7292 -309
rect 7754 -343 8310 -309
rect 8772 -343 9328 -309
rect 9790 -343 10346 -309
rect 10808 -343 11364 -309
rect 11826 -343 12382 -309
rect 12844 -343 13400 -309
rect 13862 -343 14418 -309
rect 14880 -343 15436 -309
rect 15898 -343 16454 -309
rect 16916 -343 17472 -309
rect 17934 -343 18490 -309
rect 18952 -343 19508 -309
rect 19970 -343 20526 -309
rect 20988 -343 21544 -309
rect 22006 -343 22562 -309
rect 6736 -751 7292 -717
rect 7754 -751 8310 -717
rect 8772 -751 9328 -717
rect 9790 -751 10346 -717
rect 10808 -751 11364 -717
rect 11826 -751 12382 -717
rect 12844 -751 13400 -717
rect 13862 -751 14418 -717
rect 14880 -751 15436 -717
rect 15898 -751 16454 -717
rect 16916 -751 17472 -717
rect 17934 -751 18490 -717
rect 18952 -751 19508 -717
rect 19970 -751 20526 -717
rect 20988 -751 21544 -717
rect 22006 -751 22562 -717
rect 6736 -1479 7292 -1445
rect 7754 -1479 8310 -1445
rect 8772 -1479 9328 -1445
rect 9790 -1479 10346 -1445
rect 10808 -1479 11364 -1445
rect 11826 -1479 12382 -1445
rect 12844 -1479 13400 -1445
rect 13862 -1479 14418 -1445
rect 14880 -1479 15436 -1445
rect 15898 -1479 16454 -1445
rect 16916 -1479 17472 -1445
rect 17934 -1479 18490 -1445
rect 18952 -1479 19508 -1445
rect 19970 -1479 20526 -1445
rect 20988 -1479 21544 -1445
rect 22006 -1479 22562 -1445
rect 7930 -2389 8486 -2355
rect 8948 -2389 9504 -2355
rect 9966 -2389 10522 -2355
rect 10984 -2389 11540 -2355
rect 12002 -2389 12558 -2355
rect 13020 -2389 13576 -2355
rect 14038 -2389 14594 -2355
rect 15056 -2389 15612 -2355
rect 16074 -2389 16630 -2355
rect 17092 -2389 17648 -2355
rect 18110 -2389 18666 -2355
rect 19128 -2389 19684 -2355
rect 20146 -2389 20702 -2355
rect 21164 -2389 21720 -2355
rect 7930 -3117 8486 -3083
rect 8948 -3117 9504 -3083
rect 9966 -3117 10522 -3083
rect 10984 -3117 11540 -3083
rect 12002 -3117 12558 -3083
rect 13020 -3117 13576 -3083
rect 14038 -3117 14594 -3083
rect 15056 -3117 15612 -3083
rect 16074 -3117 16630 -3083
rect 17092 -3117 17648 -3083
rect 18110 -3117 18666 -3083
rect 19128 -3117 19684 -3083
rect 20146 -3117 20702 -3083
rect 21164 -3117 21720 -3083
rect 7930 -3421 8486 -3387
rect 8948 -3421 9504 -3387
rect 9966 -3421 10522 -3387
rect 10984 -3421 11540 -3387
rect 12002 -3421 12558 -3387
rect 13020 -3421 13576 -3387
rect 14038 -3421 14594 -3387
rect 15056 -3421 15612 -3387
rect 16074 -3421 16630 -3387
rect 17092 -3421 17648 -3387
rect 18110 -3421 18666 -3387
rect 19128 -3421 19684 -3387
rect 20146 -3421 20702 -3387
rect 21164 -3421 21720 -3387
rect 7930 -4149 8486 -4115
rect 8948 -4149 9504 -4115
rect 9966 -4149 10522 -4115
rect 10984 -4149 11540 -4115
rect 12002 -4149 12558 -4115
rect 13020 -4149 13576 -4115
rect 14038 -4149 14594 -4115
rect 15056 -4149 15612 -4115
rect 16074 -4149 16630 -4115
rect 17092 -4149 17648 -4115
rect 18110 -4149 18666 -4115
rect 19128 -4149 19684 -4115
rect 20146 -4149 20702 -4115
rect 21164 -4149 21720 -4115
rect 7722 -5025 8278 -4991
rect 8740 -5025 9296 -4991
rect 9758 -5025 10314 -4991
rect 10776 -5025 11332 -4991
rect 11794 -5025 12350 -4991
rect 12812 -5025 13368 -4991
rect 13830 -5025 14386 -4991
rect 14848 -5025 15404 -4991
rect 15866 -5025 16422 -4991
rect 16884 -5025 17440 -4991
rect 17902 -5025 18458 -4991
rect 18920 -5025 19476 -4991
rect 19938 -5025 20494 -4991
rect 20956 -5025 21512 -4991
rect 21974 -5025 22530 -4991
rect 2418 -5129 2974 -5095
rect 3436 -5129 3992 -5095
rect 4454 -5129 5010 -5095
rect 5472 -5129 6028 -5095
rect 7722 -5753 8278 -5719
rect 8740 -5753 9296 -5719
rect 9758 -5753 10314 -5719
rect 10776 -5753 11332 -5719
rect 11794 -5753 12350 -5719
rect 12812 -5753 13368 -5719
rect 13830 -5753 14386 -5719
rect 14848 -5753 15404 -5719
rect 15866 -5753 16422 -5719
rect 16884 -5753 17440 -5719
rect 17902 -5753 18458 -5719
rect 18920 -5753 19476 -5719
rect 19938 -5753 20494 -5719
rect 20956 -5753 21512 -5719
rect 21974 -5753 22530 -5719
rect 2418 -5857 2974 -5823
rect 3436 -5857 3992 -5823
rect 4454 -5857 5010 -5823
rect 5472 -5857 6028 -5823
rect 2418 -6161 2974 -6127
rect 3436 -6161 3992 -6127
rect 4454 -6161 5010 -6127
rect 5472 -6161 6028 -6127
rect 7722 -6281 8278 -6247
rect 8740 -6281 9296 -6247
rect 9758 -6281 10314 -6247
rect 10776 -6281 11332 -6247
rect 11794 -6281 12350 -6247
rect 12812 -6281 13368 -6247
rect 13830 -6281 14386 -6247
rect 14848 -6281 15404 -6247
rect 15866 -6281 16422 -6247
rect 16884 -6281 17440 -6247
rect 17902 -6281 18458 -6247
rect 18920 -6281 19476 -6247
rect 19938 -6281 20494 -6247
rect 20956 -6281 21512 -6247
rect 21974 -6281 22530 -6247
rect 2418 -6889 2974 -6855
rect 3436 -6889 3992 -6855
rect 4454 -6889 5010 -6855
rect 5472 -6889 6028 -6855
rect 7722 -7009 8278 -6975
rect 8740 -7009 9296 -6975
rect 9758 -7009 10314 -6975
rect 10776 -7009 11332 -6975
rect 11794 -7009 12350 -6975
rect 12812 -7009 13368 -6975
rect 13830 -7009 14386 -6975
rect 14848 -7009 15404 -6975
rect 15866 -7009 16422 -6975
rect 16884 -7009 17440 -6975
rect 17902 -7009 18458 -6975
rect 18920 -7009 19476 -6975
rect 19938 -7009 20494 -6975
rect 20956 -7009 21512 -6975
rect 21974 -7009 22530 -6975
rect 2418 -7193 2974 -7159
rect 3436 -7193 3992 -7159
rect 4454 -7193 5010 -7159
rect 5472 -7193 6028 -7159
rect 7722 -7537 8278 -7503
rect 8740 -7537 9296 -7503
rect 9758 -7537 10314 -7503
rect 10776 -7537 11332 -7503
rect 11794 -7537 12350 -7503
rect 12812 -7537 13368 -7503
rect 13830 -7537 14386 -7503
rect 14848 -7537 15404 -7503
rect 15866 -7537 16422 -7503
rect 16884 -7537 17440 -7503
rect 17902 -7537 18458 -7503
rect 18920 -7537 19476 -7503
rect 19938 -7537 20494 -7503
rect 20956 -7537 21512 -7503
rect 21974 -7537 22530 -7503
rect 2418 -7921 2974 -7887
rect 3436 -7921 3992 -7887
rect 4454 -7921 5010 -7887
rect 5472 -7921 6028 -7887
rect 2418 -8225 2974 -8191
rect 3436 -8225 3992 -8191
rect 4454 -8225 5010 -8191
rect 5472 -8225 6028 -8191
rect 7722 -8265 8278 -8231
rect 8740 -8265 9296 -8231
rect 9758 -8265 10314 -8231
rect 10776 -8265 11332 -8231
rect 11794 -8265 12350 -8231
rect 12812 -8265 13368 -8231
rect 13830 -8265 14386 -8231
rect 14848 -8265 15404 -8231
rect 15866 -8265 16422 -8231
rect 16884 -8265 17440 -8231
rect 17902 -8265 18458 -8231
rect 18920 -8265 19476 -8231
rect 19938 -8265 20494 -8231
rect 20956 -8265 21512 -8231
rect 21974 -8265 22530 -8231
rect 7722 -8793 8278 -8759
rect 8740 -8793 9296 -8759
rect 9758 -8793 10314 -8759
rect 10776 -8793 11332 -8759
rect 11794 -8793 12350 -8759
rect 12812 -8793 13368 -8759
rect 13830 -8793 14386 -8759
rect 14848 -8793 15404 -8759
rect 15866 -8793 16422 -8759
rect 16884 -8793 17440 -8759
rect 17902 -8793 18458 -8759
rect 18920 -8793 19476 -8759
rect 19938 -8793 20494 -8759
rect 20956 -8793 21512 -8759
rect 21974 -8793 22530 -8759
rect 2418 -8953 2974 -8919
rect 3436 -8953 3992 -8919
rect 4454 -8953 5010 -8919
rect 5472 -8953 6028 -8919
rect 7722 -9521 8278 -9487
rect 8740 -9521 9296 -9487
rect 9758 -9521 10314 -9487
rect 10776 -9521 11332 -9487
rect 11794 -9521 12350 -9487
rect 12812 -9521 13368 -9487
rect 13830 -9521 14386 -9487
rect 14848 -9521 15404 -9487
rect 15866 -9521 16422 -9487
rect 16884 -9521 17440 -9487
rect 17902 -9521 18458 -9487
rect 18920 -9521 19476 -9487
rect 19938 -9521 20494 -9487
rect 20956 -9521 21512 -9487
rect 21974 -9521 22530 -9487
rect 2830 -11998 3386 -11964
rect 3848 -11998 4404 -11964
rect 4866 -11998 5422 -11964
rect 5884 -11998 6440 -11964
rect 6902 -11998 7458 -11964
rect 7920 -11998 8476 -11964
rect 8938 -11998 9494 -11964
rect 9956 -11998 10512 -11964
rect 10974 -11998 11530 -11964
rect 11992 -11998 12548 -11964
rect 13010 -11998 13566 -11964
rect 14028 -11998 14584 -11964
rect 15046 -11998 15602 -11964
rect 16064 -11998 16620 -11964
rect 17082 -11998 17638 -11964
rect 18100 -11998 18656 -11964
rect 19118 -11998 19674 -11964
rect 20136 -11998 20692 -11964
rect 21154 -11998 21710 -11964
rect 22172 -11998 22728 -11964
rect -8936 -12474 -8380 -12440
rect -7918 -12474 -7362 -12440
rect -6900 -12474 -6344 -12440
rect -5882 -12474 -5326 -12440
rect -4864 -12474 -4308 -12440
rect -3846 -12474 -3290 -12440
rect -2828 -12474 -2272 -12440
rect -1810 -12474 -1254 -12440
rect -792 -12474 -236 -12440
rect 2830 -12708 3386 -12674
rect 3848 -12708 4404 -12674
rect 4866 -12708 5422 -12674
rect 5884 -12708 6440 -12674
rect 6902 -12708 7458 -12674
rect 7920 -12708 8476 -12674
rect 8938 -12708 9494 -12674
rect 9956 -12708 10512 -12674
rect 10974 -12708 11530 -12674
rect 11992 -12708 12548 -12674
rect 13010 -12708 13566 -12674
rect 14028 -12708 14584 -12674
rect 15046 -12708 15602 -12674
rect 16064 -12708 16620 -12674
rect 17082 -12708 17638 -12674
rect 18100 -12708 18656 -12674
rect 19118 -12708 19674 -12674
rect 20136 -12708 20692 -12674
rect 21154 -12708 21710 -12674
rect 22172 -12708 22728 -12674
rect 2830 -12816 3386 -12782
rect 3848 -12816 4404 -12782
rect 4866 -12816 5422 -12782
rect 5884 -12816 6440 -12782
rect 6902 -12816 7458 -12782
rect 7920 -12816 8476 -12782
rect 8938 -12816 9494 -12782
rect 9956 -12816 10512 -12782
rect 10974 -12816 11530 -12782
rect 11992 -12816 12548 -12782
rect 13010 -12816 13566 -12782
rect 14028 -12816 14584 -12782
rect 15046 -12816 15602 -12782
rect 16064 -12816 16620 -12782
rect 17082 -12816 17638 -12782
rect 18100 -12816 18656 -12782
rect 19118 -12816 19674 -12782
rect 20136 -12816 20692 -12782
rect 21154 -12816 21710 -12782
rect 22172 -12816 22728 -12782
rect -8936 -13184 -8380 -13150
rect -7918 -13184 -7362 -13150
rect -8936 -13292 -8380 -13258
rect -6900 -13184 -6344 -13150
rect -7918 -13292 -7362 -13258
rect -5882 -13184 -5326 -13150
rect -6900 -13292 -6344 -13258
rect -4864 -13184 -4308 -13150
rect -5882 -13292 -5326 -13258
rect -3846 -13184 -3290 -13150
rect -4864 -13292 -4308 -13258
rect -2828 -13184 -2272 -13150
rect -3846 -13292 -3290 -13258
rect -1810 -13184 -1254 -13150
rect -2828 -13292 -2272 -13258
rect -792 -13184 -236 -13150
rect -1810 -13292 -1254 -13258
rect -792 -13292 -236 -13258
rect 2830 -13526 3386 -13492
rect 3848 -13526 4404 -13492
rect 4866 -13526 5422 -13492
rect 5884 -13526 6440 -13492
rect 6902 -13526 7458 -13492
rect 7920 -13526 8476 -13492
rect 8938 -13526 9494 -13492
rect 9956 -13526 10512 -13492
rect 10974 -13526 11530 -13492
rect 11992 -13526 12548 -13492
rect 13010 -13526 13566 -13492
rect 14028 -13526 14584 -13492
rect 15046 -13526 15602 -13492
rect 16064 -13526 16620 -13492
rect 17082 -13526 17638 -13492
rect 18100 -13526 18656 -13492
rect 19118 -13526 19674 -13492
rect 20136 -13526 20692 -13492
rect 21154 -13526 21710 -13492
rect 22172 -13526 22728 -13492
rect -8936 -14002 -8380 -13968
rect -7918 -14002 -7362 -13968
rect -8936 -14110 -8380 -14076
rect -6900 -14002 -6344 -13968
rect -7918 -14110 -7362 -14076
rect -5882 -14002 -5326 -13968
rect -6900 -14110 -6344 -14076
rect -4864 -14002 -4308 -13968
rect -5882 -14110 -5326 -14076
rect -3846 -14002 -3290 -13968
rect -4864 -14110 -4308 -14076
rect -2828 -14002 -2272 -13968
rect -3846 -14110 -3290 -14076
rect -1810 -14002 -1254 -13968
rect -2828 -14110 -2272 -14076
rect -792 -14002 -236 -13968
rect -1810 -14110 -1254 -14076
rect -792 -14110 -236 -14076
rect 2830 -14194 3386 -14160
rect 3848 -14194 4404 -14160
rect 4866 -14194 5422 -14160
rect 5884 -14194 6440 -14160
rect 6902 -14194 7458 -14160
rect 7920 -14194 8476 -14160
rect 8938 -14194 9494 -14160
rect 9956 -14194 10512 -14160
rect 10974 -14194 11530 -14160
rect 11992 -14194 12548 -14160
rect 13010 -14194 13566 -14160
rect 14028 -14194 14584 -14160
rect 15046 -14194 15602 -14160
rect 16064 -14194 16620 -14160
rect 17082 -14194 17638 -14160
rect 18100 -14194 18656 -14160
rect 19118 -14194 19674 -14160
rect 20136 -14194 20692 -14160
rect 21154 -14194 21710 -14160
rect 22172 -14194 22728 -14160
rect -8936 -14820 -8380 -14786
rect -7918 -14820 -7362 -14786
rect -8936 -14928 -8380 -14894
rect -6900 -14820 -6344 -14786
rect -7918 -14928 -7362 -14894
rect -5882 -14820 -5326 -14786
rect -6900 -14928 -6344 -14894
rect -4864 -14820 -4308 -14786
rect -5882 -14928 -5326 -14894
rect -3846 -14820 -3290 -14786
rect -4864 -14928 -4308 -14894
rect -2828 -14820 -2272 -14786
rect -3846 -14928 -3290 -14894
rect -1810 -14820 -1254 -14786
rect -2828 -14928 -2272 -14894
rect -792 -14820 -236 -14786
rect -1810 -14928 -1254 -14894
rect -792 -14928 -236 -14894
rect 2830 -14904 3386 -14870
rect 3848 -14904 4404 -14870
rect 4866 -14904 5422 -14870
rect 5884 -14904 6440 -14870
rect 6902 -14904 7458 -14870
rect 7920 -14904 8476 -14870
rect 8938 -14904 9494 -14870
rect 9956 -14904 10512 -14870
rect 10974 -14904 11530 -14870
rect 11992 -14904 12548 -14870
rect 13010 -14904 13566 -14870
rect 14028 -14904 14584 -14870
rect 15046 -14904 15602 -14870
rect 16064 -14904 16620 -14870
rect 17082 -14904 17638 -14870
rect 18100 -14904 18656 -14870
rect 19118 -14904 19674 -14870
rect 20136 -14904 20692 -14870
rect 21154 -14904 21710 -14870
rect 22172 -14904 22728 -14870
rect 2830 -15426 3386 -15392
rect 3848 -15426 4404 -15392
rect 4866 -15426 5422 -15392
rect 5884 -15426 6440 -15392
rect 6902 -15426 7458 -15392
rect 7920 -15426 8476 -15392
rect 8938 -15426 9494 -15392
rect 9956 -15426 10512 -15392
rect 10974 -15426 11530 -15392
rect 11992 -15426 12548 -15392
rect 13010 -15426 13566 -15392
rect 14028 -15426 14584 -15392
rect 15046 -15426 15602 -15392
rect 16064 -15426 16620 -15392
rect 17082 -15426 17638 -15392
rect 18100 -15426 18656 -15392
rect 19118 -15426 19674 -15392
rect 20136 -15426 20692 -15392
rect 21154 -15426 21710 -15392
rect 22172 -15426 22728 -15392
rect -8936 -15638 -8380 -15604
rect -7918 -15638 -7362 -15604
rect -8936 -15746 -8380 -15712
rect -6900 -15638 -6344 -15604
rect -7918 -15746 -7362 -15712
rect -5882 -15638 -5326 -15604
rect -6900 -15746 -6344 -15712
rect -4864 -15638 -4308 -15604
rect -5882 -15746 -5326 -15712
rect -3846 -15638 -3290 -15604
rect -4864 -15746 -4308 -15712
rect -2828 -15638 -2272 -15604
rect -3846 -15746 -3290 -15712
rect -1810 -15638 -1254 -15604
rect -2828 -15746 -2272 -15712
rect -792 -15638 -236 -15604
rect -1810 -15746 -1254 -15712
rect -792 -15746 -236 -15712
rect 2830 -16136 3386 -16102
rect 3848 -16136 4404 -16102
rect 4866 -16136 5422 -16102
rect 5884 -16136 6440 -16102
rect 6902 -16136 7458 -16102
rect 7920 -16136 8476 -16102
rect 8938 -16136 9494 -16102
rect 9956 -16136 10512 -16102
rect 10974 -16136 11530 -16102
rect 11992 -16136 12548 -16102
rect 13010 -16136 13566 -16102
rect 14028 -16136 14584 -16102
rect 15046 -16136 15602 -16102
rect 16064 -16136 16620 -16102
rect 17082 -16136 17638 -16102
rect 18100 -16136 18656 -16102
rect 19118 -16136 19674 -16102
rect 20136 -16136 20692 -16102
rect 21154 -16136 21710 -16102
rect 22172 -16136 22728 -16102
rect -8936 -16456 -8380 -16422
rect -7918 -16456 -7362 -16422
rect -8936 -16564 -8380 -16530
rect -6900 -16456 -6344 -16422
rect -7918 -16564 -7362 -16530
rect -5882 -16456 -5326 -16422
rect -6900 -16564 -6344 -16530
rect -4864 -16456 -4308 -16422
rect -5882 -16564 -5326 -16530
rect -3846 -16456 -3290 -16422
rect -4864 -16564 -4308 -16530
rect -2828 -16456 -2272 -16422
rect -3846 -16564 -3290 -16530
rect -1810 -16456 -1254 -16422
rect -2828 -16564 -2272 -16530
rect -792 -16456 -236 -16422
rect -1810 -16564 -1254 -16530
rect -792 -16564 -236 -16530
rect 2828 -16660 3384 -16626
rect 3846 -16660 4402 -16626
rect 4864 -16660 5420 -16626
rect 5882 -16660 6438 -16626
rect 6900 -16660 7456 -16626
rect 7918 -16660 8474 -16626
rect 8936 -16660 9492 -16626
rect 9954 -16660 10510 -16626
rect 10972 -16660 11528 -16626
rect 11990 -16660 12546 -16626
rect 13008 -16660 13564 -16626
rect 14026 -16660 14582 -16626
rect 15044 -16660 15600 -16626
rect 16062 -16660 16618 -16626
rect 17080 -16660 17636 -16626
rect 18098 -16660 18654 -16626
rect 19116 -16660 19672 -16626
rect 20134 -16660 20690 -16626
rect 21152 -16660 21708 -16626
rect 22170 -16660 22726 -16626
rect -8936 -17274 -8380 -17240
rect -7918 -17274 -7362 -17240
rect -8936 -17382 -8380 -17348
rect -6900 -17274 -6344 -17240
rect -7918 -17382 -7362 -17348
rect -5882 -17274 -5326 -17240
rect -6900 -17382 -6344 -17348
rect -4864 -17274 -4308 -17240
rect -5882 -17382 -5326 -17348
rect -3846 -17274 -3290 -17240
rect -4864 -17382 -4308 -17348
rect -2828 -17274 -2272 -17240
rect -3846 -17382 -3290 -17348
rect -1810 -17274 -1254 -17240
rect -2828 -17382 -2272 -17348
rect -792 -17274 -236 -17240
rect -1810 -17382 -1254 -17348
rect -792 -17382 -236 -17348
rect 2828 -17370 3384 -17336
rect 3846 -17370 4402 -17336
rect 4864 -17370 5420 -17336
rect 5882 -17370 6438 -17336
rect 6900 -17370 7456 -17336
rect 7918 -17370 8474 -17336
rect 8936 -17370 9492 -17336
rect 9954 -17370 10510 -17336
rect 10972 -17370 11528 -17336
rect 11990 -17370 12546 -17336
rect 13008 -17370 13564 -17336
rect 14026 -17370 14582 -17336
rect 15044 -17370 15600 -17336
rect 16062 -17370 16618 -17336
rect 17080 -17370 17636 -17336
rect 18098 -17370 18654 -17336
rect 19116 -17370 19672 -17336
rect 20134 -17370 20690 -17336
rect 21152 -17370 21708 -17336
rect 22170 -17370 22726 -17336
rect 2828 -17894 3384 -17860
rect 3846 -17894 4402 -17860
rect 4864 -17894 5420 -17860
rect 5882 -17894 6438 -17860
rect 6900 -17894 7456 -17860
rect 7918 -17894 8474 -17860
rect 8936 -17894 9492 -17860
rect 9954 -17894 10510 -17860
rect 10972 -17894 11528 -17860
rect 11990 -17894 12546 -17860
rect 13008 -17894 13564 -17860
rect 14026 -17894 14582 -17860
rect 15044 -17894 15600 -17860
rect 16062 -17894 16618 -17860
rect 17080 -17894 17636 -17860
rect 18098 -17894 18654 -17860
rect 19116 -17894 19672 -17860
rect 20134 -17894 20690 -17860
rect 21152 -17894 21708 -17860
rect 22170 -17894 22726 -17860
rect -8936 -18092 -8380 -18058
rect -7918 -18092 -7362 -18058
rect -8936 -18200 -8380 -18166
rect -6900 -18092 -6344 -18058
rect -7918 -18200 -7362 -18166
rect -5882 -18092 -5326 -18058
rect -6900 -18200 -6344 -18166
rect -4864 -18092 -4308 -18058
rect -5882 -18200 -5326 -18166
rect -3846 -18092 -3290 -18058
rect -4864 -18200 -4308 -18166
rect -2828 -18092 -2272 -18058
rect -3846 -18200 -3290 -18166
rect -1810 -18092 -1254 -18058
rect -2828 -18200 -2272 -18166
rect -792 -18092 -236 -18058
rect -1810 -18200 -1254 -18166
rect -792 -18200 -236 -18166
rect 2828 -18604 3384 -18570
rect 3846 -18604 4402 -18570
rect 4864 -18604 5420 -18570
rect 5882 -18604 6438 -18570
rect 6900 -18604 7456 -18570
rect 7918 -18604 8474 -18570
rect 8936 -18604 9492 -18570
rect 9954 -18604 10510 -18570
rect 10972 -18604 11528 -18570
rect 11990 -18604 12546 -18570
rect 13008 -18604 13564 -18570
rect 14026 -18604 14582 -18570
rect 15044 -18604 15600 -18570
rect 16062 -18604 16618 -18570
rect 17080 -18604 17636 -18570
rect 18098 -18604 18654 -18570
rect 19116 -18604 19672 -18570
rect 20134 -18604 20690 -18570
rect 21152 -18604 21708 -18570
rect 22170 -18604 22726 -18570
rect -8936 -18910 -8380 -18876
rect -7918 -18910 -7362 -18876
rect -6900 -18910 -6344 -18876
rect -5882 -18910 -5326 -18876
rect -4864 -18910 -4308 -18876
rect -3846 -18910 -3290 -18876
rect -2828 -18910 -2272 -18876
rect -1810 -18910 -1254 -18876
rect -792 -18910 -236 -18876
rect 2828 -19126 3384 -19092
rect 3846 -19126 4402 -19092
rect 4864 -19126 5420 -19092
rect 5882 -19126 6438 -19092
rect 6900 -19126 7456 -19092
rect 7918 -19126 8474 -19092
rect 8936 -19126 9492 -19092
rect 9954 -19126 10510 -19092
rect 10972 -19126 11528 -19092
rect 11990 -19126 12546 -19092
rect 13008 -19126 13564 -19092
rect 14026 -19126 14582 -19092
rect 15044 -19126 15600 -19092
rect 16062 -19126 16618 -19092
rect 17080 -19126 17636 -19092
rect 18098 -19126 18654 -19092
rect 19116 -19126 19672 -19092
rect 20134 -19126 20690 -19092
rect 21152 -19126 21708 -19092
rect 22170 -19126 22726 -19092
rect 2828 -19836 3384 -19802
rect 3846 -19836 4402 -19802
rect 4864 -19836 5420 -19802
rect 5882 -19836 6438 -19802
rect 6900 -19836 7456 -19802
rect 7918 -19836 8474 -19802
rect 8936 -19836 9492 -19802
rect 9954 -19836 10510 -19802
rect 10972 -19836 11528 -19802
rect 11990 -19836 12546 -19802
rect 13008 -19836 13564 -19802
rect 14026 -19836 14582 -19802
rect 15044 -19836 15600 -19802
rect 16062 -19836 16618 -19802
rect 17080 -19836 17636 -19802
rect 18098 -19836 18654 -19802
rect 19116 -19836 19672 -19802
rect 20134 -19836 20690 -19802
rect 21152 -19836 21708 -19802
rect 22170 -19836 22726 -19802
rect -10260 -20224 -9704 -20190
rect -9242 -20224 -8686 -20190
rect -8224 -20224 -7668 -20190
rect -7206 -20224 -6650 -20190
rect -6188 -20224 -5632 -20190
rect -5170 -20224 -4614 -20190
rect -4152 -20224 -3596 -20190
rect -3134 -20224 -2578 -20190
rect -2116 -20224 -1560 -20190
rect -1098 -20224 -542 -20190
rect -80 -20224 476 -20190
rect 2828 -20360 3384 -20326
rect 3846 -20360 4402 -20326
rect 4864 -20360 5420 -20326
rect 5882 -20360 6438 -20326
rect 6900 -20360 7456 -20326
rect 7918 -20360 8474 -20326
rect 8936 -20360 9492 -20326
rect 9954 -20360 10510 -20326
rect 10972 -20360 11528 -20326
rect 11990 -20360 12546 -20326
rect 13008 -20360 13564 -20326
rect 14026 -20360 14582 -20326
rect 15044 -20360 15600 -20326
rect 16062 -20360 16618 -20326
rect 17080 -20360 17636 -20326
rect 18098 -20360 18654 -20326
rect 19116 -20360 19672 -20326
rect 20134 -20360 20690 -20326
rect 21152 -20360 21708 -20326
rect 22170 -20360 22726 -20326
rect -10260 -20934 -9704 -20900
rect -9242 -20934 -8686 -20900
rect -8224 -20934 -7668 -20900
rect -7206 -20934 -6650 -20900
rect -6188 -20934 -5632 -20900
rect -5170 -20934 -4614 -20900
rect -4152 -20934 -3596 -20900
rect -3134 -20934 -2578 -20900
rect -2116 -20934 -1560 -20900
rect -1098 -20934 -542 -20900
rect -80 -20934 476 -20900
rect 2828 -21070 3384 -21036
rect 3846 -21070 4402 -21036
rect 4864 -21070 5420 -21036
rect 5882 -21070 6438 -21036
rect 6900 -21070 7456 -21036
rect 7918 -21070 8474 -21036
rect 8936 -21070 9492 -21036
rect 9954 -21070 10510 -21036
rect 10972 -21070 11528 -21036
rect 11990 -21070 12546 -21036
rect 13008 -21070 13564 -21036
rect 14026 -21070 14582 -21036
rect 15044 -21070 15600 -21036
rect 16062 -21070 16618 -21036
rect 17080 -21070 17636 -21036
rect 18098 -21070 18654 -21036
rect 19116 -21070 19672 -21036
rect 20134 -21070 20690 -21036
rect 21152 -21070 21708 -21036
rect 22170 -21070 22726 -21036
rect -10260 -21336 -9704 -21302
rect -9242 -21336 -8686 -21302
rect -8224 -21336 -7668 -21302
rect -7206 -21336 -6650 -21302
rect -6188 -21336 -5632 -21302
rect -5170 -21336 -4614 -21302
rect -4152 -21336 -3596 -21302
rect -3134 -21336 -2578 -21302
rect -2116 -21336 -1560 -21302
rect -1098 -21336 -542 -21302
rect -80 -21336 476 -21302
rect 2828 -21594 3384 -21560
rect 3846 -21594 4402 -21560
rect 4864 -21594 5420 -21560
rect 5882 -21594 6438 -21560
rect 6900 -21594 7456 -21560
rect 7918 -21594 8474 -21560
rect 8936 -21594 9492 -21560
rect 9954 -21594 10510 -21560
rect 10972 -21594 11528 -21560
rect 11990 -21594 12546 -21560
rect 13008 -21594 13564 -21560
rect 14026 -21594 14582 -21560
rect 15044 -21594 15600 -21560
rect 16062 -21594 16618 -21560
rect 17080 -21594 17636 -21560
rect 18098 -21594 18654 -21560
rect 19116 -21594 19672 -21560
rect 20134 -21594 20690 -21560
rect 21152 -21594 21708 -21560
rect 22170 -21594 22726 -21560
rect -10260 -22046 -9704 -22012
rect -9242 -22046 -8686 -22012
rect -8224 -22046 -7668 -22012
rect -7206 -22046 -6650 -22012
rect -6188 -22046 -5632 -22012
rect -5170 -22046 -4614 -22012
rect -4152 -22046 -3596 -22012
rect -3134 -22046 -2578 -22012
rect -2116 -22046 -1560 -22012
rect -1098 -22046 -542 -22012
rect -80 -22046 476 -22012
rect 2828 -22304 3384 -22270
rect 3846 -22304 4402 -22270
rect 4864 -22304 5420 -22270
rect 5882 -22304 6438 -22270
rect 6900 -22304 7456 -22270
rect 7918 -22304 8474 -22270
rect 8936 -22304 9492 -22270
rect 9954 -22304 10510 -22270
rect 10972 -22304 11528 -22270
rect 11990 -22304 12546 -22270
rect 13008 -22304 13564 -22270
rect 14026 -22304 14582 -22270
rect 15044 -22304 15600 -22270
rect 16062 -22304 16618 -22270
rect 17080 -22304 17636 -22270
rect 18098 -22304 18654 -22270
rect 19116 -22304 19672 -22270
rect 20134 -22304 20690 -22270
rect 21152 -22304 21708 -22270
rect 22170 -22304 22726 -22270
rect -10260 -22448 -9704 -22414
rect -9242 -22448 -8686 -22414
rect -8224 -22448 -7668 -22414
rect -7206 -22448 -6650 -22414
rect -6188 -22448 -5632 -22414
rect -5170 -22448 -4614 -22414
rect -4152 -22448 -3596 -22414
rect -3134 -22448 -2578 -22414
rect -2116 -22448 -1560 -22414
rect -1098 -22448 -542 -22414
rect -80 -22448 476 -22414
rect 2828 -22826 3384 -22792
rect 3846 -22826 4402 -22792
rect 4864 -22826 5420 -22792
rect 5882 -22826 6438 -22792
rect 6900 -22826 7456 -22792
rect 7918 -22826 8474 -22792
rect 8936 -22826 9492 -22792
rect 9954 -22826 10510 -22792
rect 10972 -22826 11528 -22792
rect 11990 -22826 12546 -22792
rect 13008 -22826 13564 -22792
rect 14026 -22826 14582 -22792
rect 15044 -22826 15600 -22792
rect 16062 -22826 16618 -22792
rect 17080 -22826 17636 -22792
rect 18098 -22826 18654 -22792
rect 19116 -22826 19672 -22792
rect 20134 -22826 20690 -22792
rect 21152 -22826 21708 -22792
rect 22170 -22826 22726 -22792
rect -10260 -23158 -9704 -23124
rect -9242 -23158 -8686 -23124
rect -8224 -23158 -7668 -23124
rect -7206 -23158 -6650 -23124
rect -6188 -23158 -5632 -23124
rect -5170 -23158 -4614 -23124
rect -4152 -23158 -3596 -23124
rect -3134 -23158 -2578 -23124
rect -2116 -23158 -1560 -23124
rect -1098 -23158 -542 -23124
rect -80 -23158 476 -23124
rect -10260 -23560 -9704 -23526
rect -9242 -23560 -8686 -23526
rect -8224 -23560 -7668 -23526
rect -7206 -23560 -6650 -23526
rect -6188 -23560 -5632 -23526
rect -5170 -23560 -4614 -23526
rect -4152 -23560 -3596 -23526
rect -3134 -23560 -2578 -23526
rect -2116 -23560 -1560 -23526
rect -1098 -23560 -542 -23526
rect -80 -23560 476 -23526
rect 2828 -23536 3384 -23502
rect 3846 -23536 4402 -23502
rect 4864 -23536 5420 -23502
rect 5882 -23536 6438 -23502
rect 6900 -23536 7456 -23502
rect 7918 -23536 8474 -23502
rect 8936 -23536 9492 -23502
rect 9954 -23536 10510 -23502
rect 10972 -23536 11528 -23502
rect 11990 -23536 12546 -23502
rect 13008 -23536 13564 -23502
rect 14026 -23536 14582 -23502
rect 15044 -23536 15600 -23502
rect 16062 -23536 16618 -23502
rect 17080 -23536 17636 -23502
rect 18098 -23536 18654 -23502
rect 19116 -23536 19672 -23502
rect 20134 -23536 20690 -23502
rect 21152 -23536 21708 -23502
rect 22170 -23536 22726 -23502
rect 2828 -24060 3384 -24026
rect 3846 -24060 4402 -24026
rect 4864 -24060 5420 -24026
rect 5882 -24060 6438 -24026
rect 6900 -24060 7456 -24026
rect 7918 -24060 8474 -24026
rect 8936 -24060 9492 -24026
rect 9954 -24060 10510 -24026
rect 10972 -24060 11528 -24026
rect 11990 -24060 12546 -24026
rect 13008 -24060 13564 -24026
rect 14026 -24060 14582 -24026
rect 15044 -24060 15600 -24026
rect 16062 -24060 16618 -24026
rect 17080 -24060 17636 -24026
rect 18098 -24060 18654 -24026
rect 19116 -24060 19672 -24026
rect 20134 -24060 20690 -24026
rect 21152 -24060 21708 -24026
rect 22170 -24060 22726 -24026
rect -10260 -24270 -9704 -24236
rect -9242 -24270 -8686 -24236
rect -8224 -24270 -7668 -24236
rect -7206 -24270 -6650 -24236
rect -6188 -24270 -5632 -24236
rect -5170 -24270 -4614 -24236
rect -4152 -24270 -3596 -24236
rect -3134 -24270 -2578 -24236
rect -2116 -24270 -1560 -24236
rect -1098 -24270 -542 -24236
rect -80 -24270 476 -24236
rect 2828 -24770 3384 -24736
rect 3846 -24770 4402 -24736
rect 4864 -24770 5420 -24736
rect 5882 -24770 6438 -24736
rect 6900 -24770 7456 -24736
rect 7918 -24770 8474 -24736
rect 8936 -24770 9492 -24736
rect 9954 -24770 10510 -24736
rect 10972 -24770 11528 -24736
rect 11990 -24770 12546 -24736
rect 13008 -24770 13564 -24736
rect 14026 -24770 14582 -24736
rect 15044 -24770 15600 -24736
rect 16062 -24770 16618 -24736
rect 17080 -24770 17636 -24736
rect 18098 -24770 18654 -24736
rect 19116 -24770 19672 -24736
rect 20134 -24770 20690 -24736
rect 21152 -24770 21708 -24736
rect 22170 -24770 22726 -24736
rect -9802 -25102 -9246 -25068
rect -8784 -25102 -8228 -25068
rect -7766 -25102 -7210 -25068
rect -6748 -25102 -6192 -25068
rect -5730 -25102 -5174 -25068
rect -4712 -25102 -4156 -25068
rect -3694 -25102 -3138 -25068
rect -2676 -25102 -2120 -25068
rect -1658 -25102 -1102 -25068
rect -640 -25102 -84 -25068
rect 2828 -25292 3384 -25258
rect 3846 -25292 4402 -25258
rect 4864 -25292 5420 -25258
rect 5882 -25292 6438 -25258
rect 6900 -25292 7456 -25258
rect 7918 -25292 8474 -25258
rect 8936 -25292 9492 -25258
rect 9954 -25292 10510 -25258
rect 10972 -25292 11528 -25258
rect 11990 -25292 12546 -25258
rect 13008 -25292 13564 -25258
rect 14026 -25292 14582 -25258
rect 15044 -25292 15600 -25258
rect 16062 -25292 16618 -25258
rect 17080 -25292 17636 -25258
rect 18098 -25292 18654 -25258
rect 19116 -25292 19672 -25258
rect 20134 -25292 20690 -25258
rect 21152 -25292 21708 -25258
rect 22170 -25292 22726 -25258
rect -9802 -25812 -9246 -25778
rect -8784 -25812 -8228 -25778
rect -7766 -25812 -7210 -25778
rect -6748 -25812 -6192 -25778
rect -5730 -25812 -5174 -25778
rect -4712 -25812 -4156 -25778
rect -3694 -25812 -3138 -25778
rect -2676 -25812 -2120 -25778
rect -1658 -25812 -1102 -25778
rect -640 -25812 -84 -25778
rect 2828 -26002 3384 -25968
rect 3846 -26002 4402 -25968
rect 4864 -26002 5420 -25968
rect 5882 -26002 6438 -25968
rect 6900 -26002 7456 -25968
rect 7918 -26002 8474 -25968
rect 8936 -26002 9492 -25968
rect 9954 -26002 10510 -25968
rect 10972 -26002 11528 -25968
rect 11990 -26002 12546 -25968
rect 13008 -26002 13564 -25968
rect 14026 -26002 14582 -25968
rect 15044 -26002 15600 -25968
rect 16062 -26002 16618 -25968
rect 17080 -26002 17636 -25968
rect 18098 -26002 18654 -25968
rect 19116 -26002 19672 -25968
rect 20134 -26002 20690 -25968
rect 21152 -26002 21708 -25968
rect 22170 -26002 22726 -25968
<< locali >>
rect 378 4160 478 4322
rect 24722 4160 24822 4322
rect 6968 1778 7058 1808
rect 6968 1744 6996 1778
rect 7030 1744 7058 1778
rect 6968 1716 7058 1744
rect 7986 1778 8076 1808
rect 7986 1744 8014 1778
rect 8048 1744 8076 1778
rect 7986 1716 8076 1744
rect 9004 1778 9094 1808
rect 9004 1744 9032 1778
rect 9066 1744 9094 1778
rect 9004 1716 9094 1744
rect 10022 1778 10112 1808
rect 10022 1744 10050 1778
rect 10084 1744 10112 1778
rect 10022 1716 10112 1744
rect 11040 1778 11130 1808
rect 11040 1744 11068 1778
rect 11102 1744 11130 1778
rect 11040 1716 11130 1744
rect 12058 1778 12148 1808
rect 12058 1744 12086 1778
rect 12120 1744 12148 1778
rect 12058 1716 12148 1744
rect 13076 1778 13166 1808
rect 13076 1744 13104 1778
rect 13138 1744 13166 1778
rect 13076 1716 13166 1744
rect 14094 1778 14184 1808
rect 14094 1744 14122 1778
rect 14156 1744 14184 1778
rect 14094 1716 14184 1744
rect 15112 1778 15202 1808
rect 15112 1744 15140 1778
rect 15174 1744 15202 1778
rect 15112 1716 15202 1744
rect 16130 1778 16220 1808
rect 16130 1744 16158 1778
rect 16192 1744 16220 1778
rect 16130 1716 16220 1744
rect 17148 1778 17238 1808
rect 17148 1744 17176 1778
rect 17210 1744 17238 1778
rect 17148 1716 17238 1744
rect 18166 1778 18256 1808
rect 18166 1744 18194 1778
rect 18228 1744 18256 1778
rect 18166 1716 18256 1744
rect 19184 1778 19274 1808
rect 19184 1744 19212 1778
rect 19246 1744 19274 1778
rect 19184 1716 19274 1744
rect 20202 1778 20292 1808
rect 20202 1744 20230 1778
rect 20264 1744 20292 1778
rect 20202 1716 20292 1744
rect 21220 1778 21310 1808
rect 21220 1744 21248 1778
rect 21282 1744 21310 1778
rect 21220 1716 21310 1744
rect 22238 1778 22328 1808
rect 22238 1744 22266 1778
rect 22300 1744 22328 1778
rect 22238 1716 22328 1744
rect 6720 1521 6736 1555
rect 7292 1521 7308 1555
rect 7738 1521 7754 1555
rect 8310 1521 8326 1555
rect 8756 1521 8772 1555
rect 9328 1521 9344 1555
rect 9774 1521 9790 1555
rect 10346 1521 10362 1555
rect 10792 1521 10808 1555
rect 11364 1521 11380 1555
rect 11810 1521 11826 1555
rect 12382 1521 12398 1555
rect 12828 1521 12844 1555
rect 13400 1521 13416 1555
rect 13846 1521 13862 1555
rect 14418 1521 14434 1555
rect 14864 1521 14880 1555
rect 15436 1521 15452 1555
rect 15882 1521 15898 1555
rect 16454 1521 16470 1555
rect 16900 1521 16916 1555
rect 17472 1521 17488 1555
rect 17918 1521 17934 1555
rect 18490 1521 18506 1555
rect 18936 1521 18952 1555
rect 19508 1521 19524 1555
rect 19954 1521 19970 1555
rect 20526 1521 20542 1555
rect 20972 1521 20988 1555
rect 21544 1521 21560 1555
rect 21990 1521 22006 1555
rect 22562 1521 22578 1555
rect 6488 1462 6522 1478
rect 6488 870 6522 886
rect 7506 1462 7540 1478
rect 7506 870 7540 886
rect 8524 1462 8558 1478
rect 8524 870 8558 886
rect 9542 1462 9576 1478
rect 9542 870 9576 886
rect 10560 1462 10594 1478
rect 10560 870 10594 886
rect 11578 1462 11612 1478
rect 11578 870 11612 886
rect 12596 1462 12630 1478
rect 12596 870 12630 886
rect 13614 1462 13648 1478
rect 13614 870 13648 886
rect 14632 1462 14666 1478
rect 14632 870 14666 886
rect 15650 1462 15684 1478
rect 15650 870 15684 886
rect 16668 1462 16702 1478
rect 16668 870 16702 886
rect 17686 1462 17720 1478
rect 17686 870 17720 886
rect 18704 1462 18738 1478
rect 18704 870 18738 886
rect 19722 1462 19756 1478
rect 19722 870 19756 886
rect 20740 1462 20774 1478
rect 20740 870 20774 886
rect 21758 1462 21792 1478
rect 21758 870 21792 886
rect 22776 1462 22810 1478
rect 22776 870 22810 886
rect 6720 793 6736 827
rect 7292 793 7308 827
rect 7738 793 7754 827
rect 8310 793 8326 827
rect 8756 793 8772 827
rect 9328 793 9344 827
rect 9774 793 9790 827
rect 10346 793 10362 827
rect 10792 793 10808 827
rect 11364 793 11380 827
rect 11810 793 11826 827
rect 12382 793 12398 827
rect 12828 793 12844 827
rect 13400 793 13416 827
rect 13846 793 13862 827
rect 14418 793 14434 827
rect 14864 793 14880 827
rect 15436 793 15452 827
rect 15882 793 15898 827
rect 16454 793 16470 827
rect 16900 793 16916 827
rect 17472 793 17488 827
rect 17918 793 17934 827
rect 18490 793 18506 827
rect 18936 793 18952 827
rect 19508 793 19524 827
rect 19954 793 19970 827
rect 20526 793 20542 827
rect 20972 793 20988 827
rect 21544 793 21560 827
rect 21990 793 22006 827
rect 22562 793 22578 827
rect 6990 624 7080 654
rect 6990 590 7018 624
rect 7052 590 7080 624
rect 6990 562 7080 590
rect 8008 624 8098 654
rect 8008 590 8036 624
rect 8070 590 8098 624
rect 8008 562 8098 590
rect 9026 624 9116 654
rect 9026 590 9054 624
rect 9088 590 9116 624
rect 9026 562 9116 590
rect 10044 624 10134 654
rect 10044 590 10072 624
rect 10106 590 10134 624
rect 10044 562 10134 590
rect 11062 624 11152 654
rect 11062 590 11090 624
rect 11124 590 11152 624
rect 11062 562 11152 590
rect 12080 624 12170 654
rect 12080 590 12108 624
rect 12142 590 12170 624
rect 12080 562 12170 590
rect 13098 624 13188 654
rect 13098 590 13126 624
rect 13160 590 13188 624
rect 13098 562 13188 590
rect 14116 624 14206 654
rect 14116 590 14144 624
rect 14178 590 14206 624
rect 14116 562 14206 590
rect 15134 624 15224 654
rect 15134 590 15162 624
rect 15196 590 15224 624
rect 15134 562 15224 590
rect 16152 624 16242 654
rect 16152 590 16180 624
rect 16214 590 16242 624
rect 16152 562 16242 590
rect 17170 624 17260 654
rect 17170 590 17198 624
rect 17232 590 17260 624
rect 17170 562 17260 590
rect 18188 624 18278 654
rect 18188 590 18216 624
rect 18250 590 18278 624
rect 18188 562 18278 590
rect 19206 624 19296 654
rect 19206 590 19234 624
rect 19268 590 19296 624
rect 19206 562 19296 590
rect 20224 624 20314 654
rect 20224 590 20252 624
rect 20286 590 20314 624
rect 20224 562 20314 590
rect 21242 624 21332 654
rect 21242 590 21270 624
rect 21304 590 21332 624
rect 21242 562 21332 590
rect 22260 624 22350 654
rect 22260 590 22288 624
rect 22322 590 22350 624
rect 22260 562 22350 590
rect 6720 385 6736 419
rect 7292 385 7308 419
rect 7738 385 7754 419
rect 8310 385 8326 419
rect 8756 385 8772 419
rect 9328 385 9344 419
rect 9774 385 9790 419
rect 10346 385 10362 419
rect 10792 385 10808 419
rect 11364 385 11380 419
rect 11810 385 11826 419
rect 12382 385 12398 419
rect 12828 385 12844 419
rect 13400 385 13416 419
rect 13846 385 13862 419
rect 14418 385 14434 419
rect 14864 385 14880 419
rect 15436 385 15452 419
rect 15882 385 15898 419
rect 16454 385 16470 419
rect 16900 385 16916 419
rect 17472 385 17488 419
rect 17918 385 17934 419
rect 18490 385 18506 419
rect 18936 385 18952 419
rect 19508 385 19524 419
rect 19954 385 19970 419
rect 20526 385 20542 419
rect 20972 385 20988 419
rect 21544 385 21560 419
rect 21990 385 22006 419
rect 22562 385 22578 419
rect 6488 326 6522 342
rect 6488 -266 6522 -250
rect 7506 326 7540 342
rect 7506 -266 7540 -250
rect 8524 326 8558 342
rect 8524 -266 8558 -250
rect 9542 326 9576 342
rect 9542 -266 9576 -250
rect 10560 326 10594 342
rect 10560 -266 10594 -250
rect 11578 326 11612 342
rect 11578 -266 11612 -250
rect 12596 326 12630 342
rect 12596 -266 12630 -250
rect 13614 326 13648 342
rect 13614 -266 13648 -250
rect 14632 326 14666 342
rect 14632 -266 14666 -250
rect 15650 326 15684 342
rect 15650 -266 15684 -250
rect 16668 326 16702 342
rect 16668 -266 16702 -250
rect 17686 326 17720 342
rect 17686 -266 17720 -250
rect 18704 326 18738 342
rect 18704 -266 18738 -250
rect 19722 326 19756 342
rect 19722 -266 19756 -250
rect 20740 326 20774 342
rect 20740 -266 20774 -250
rect 21758 326 21792 342
rect 21758 -266 21792 -250
rect 22776 326 22810 342
rect 22776 -266 22810 -250
rect 6720 -343 6736 -309
rect 7292 -343 7308 -309
rect 7738 -343 7754 -309
rect 8310 -343 8326 -309
rect 8756 -343 8772 -309
rect 9328 -343 9344 -309
rect 9774 -343 9790 -309
rect 10346 -343 10362 -309
rect 10792 -343 10808 -309
rect 11364 -343 11380 -309
rect 11810 -343 11826 -309
rect 12382 -343 12398 -309
rect 12828 -343 12844 -309
rect 13400 -343 13416 -309
rect 13846 -343 13862 -309
rect 14418 -343 14434 -309
rect 14864 -343 14880 -309
rect 15436 -343 15452 -309
rect 15882 -343 15898 -309
rect 16454 -343 16470 -309
rect 16900 -343 16916 -309
rect 17472 -343 17488 -309
rect 17918 -343 17934 -309
rect 18490 -343 18506 -309
rect 18936 -343 18952 -309
rect 19508 -343 19524 -309
rect 19954 -343 19970 -309
rect 20526 -343 20542 -309
rect 20972 -343 20988 -309
rect 21544 -343 21560 -309
rect 21990 -343 22006 -309
rect 22562 -343 22578 -309
rect 6968 -508 7058 -478
rect 6968 -542 6996 -508
rect 7030 -542 7058 -508
rect 6968 -570 7058 -542
rect 7986 -508 8076 -478
rect 7986 -542 8014 -508
rect 8048 -542 8076 -508
rect 7986 -570 8076 -542
rect 9004 -508 9094 -478
rect 9004 -542 9032 -508
rect 9066 -542 9094 -508
rect 9004 -570 9094 -542
rect 10022 -508 10112 -478
rect 10022 -542 10050 -508
rect 10084 -542 10112 -508
rect 10022 -570 10112 -542
rect 11040 -508 11130 -478
rect 11040 -542 11068 -508
rect 11102 -542 11130 -508
rect 11040 -570 11130 -542
rect 12058 -508 12148 -478
rect 12058 -542 12086 -508
rect 12120 -542 12148 -508
rect 12058 -570 12148 -542
rect 13076 -508 13166 -478
rect 13076 -542 13104 -508
rect 13138 -542 13166 -508
rect 13076 -570 13166 -542
rect 14094 -508 14184 -478
rect 14094 -542 14122 -508
rect 14156 -542 14184 -508
rect 14094 -570 14184 -542
rect 15112 -508 15202 -478
rect 15112 -542 15140 -508
rect 15174 -542 15202 -508
rect 15112 -570 15202 -542
rect 16130 -508 16220 -478
rect 16130 -542 16158 -508
rect 16192 -542 16220 -508
rect 16130 -570 16220 -542
rect 17148 -508 17238 -478
rect 17148 -542 17176 -508
rect 17210 -542 17238 -508
rect 17148 -570 17238 -542
rect 18166 -508 18256 -478
rect 18166 -542 18194 -508
rect 18228 -542 18256 -508
rect 18166 -570 18256 -542
rect 19184 -508 19274 -478
rect 19184 -542 19212 -508
rect 19246 -542 19274 -508
rect 19184 -570 19274 -542
rect 20202 -508 20292 -478
rect 20202 -542 20230 -508
rect 20264 -542 20292 -508
rect 20202 -570 20292 -542
rect 21220 -508 21310 -478
rect 21220 -542 21248 -508
rect 21282 -542 21310 -508
rect 21220 -570 21310 -542
rect 22238 -508 22328 -478
rect 22238 -542 22266 -508
rect 22300 -542 22328 -508
rect 22238 -570 22328 -542
rect 6720 -751 6736 -717
rect 7292 -751 7308 -717
rect 7738 -751 7754 -717
rect 8310 -751 8326 -717
rect 8756 -751 8772 -717
rect 9328 -751 9344 -717
rect 9774 -751 9790 -717
rect 10346 -751 10362 -717
rect 10792 -751 10808 -717
rect 11364 -751 11380 -717
rect 11810 -751 11826 -717
rect 12382 -751 12398 -717
rect 12828 -751 12844 -717
rect 13400 -751 13416 -717
rect 13846 -751 13862 -717
rect 14418 -751 14434 -717
rect 14864 -751 14880 -717
rect 15436 -751 15452 -717
rect 15882 -751 15898 -717
rect 16454 -751 16470 -717
rect 16900 -751 16916 -717
rect 17472 -751 17488 -717
rect 17918 -751 17934 -717
rect 18490 -751 18506 -717
rect 18936 -751 18952 -717
rect 19508 -751 19524 -717
rect 19954 -751 19970 -717
rect 20526 -751 20542 -717
rect 20972 -751 20988 -717
rect 21544 -751 21560 -717
rect 21990 -751 22006 -717
rect 22562 -751 22578 -717
rect 6488 -810 6522 -794
rect 6488 -1402 6522 -1386
rect 7506 -810 7540 -794
rect 7506 -1402 7540 -1386
rect 8524 -810 8558 -794
rect 8524 -1402 8558 -1386
rect 9542 -810 9576 -794
rect 9542 -1402 9576 -1386
rect 10560 -810 10594 -794
rect 10560 -1402 10594 -1386
rect 11578 -810 11612 -794
rect 11578 -1402 11612 -1386
rect 12596 -810 12630 -794
rect 12596 -1402 12630 -1386
rect 13614 -810 13648 -794
rect 13614 -1402 13648 -1386
rect 14632 -810 14666 -794
rect 14632 -1402 14666 -1386
rect 15650 -810 15684 -794
rect 15650 -1402 15684 -1386
rect 16668 -810 16702 -794
rect 16668 -1402 16702 -1386
rect 17686 -810 17720 -794
rect 17686 -1402 17720 -1386
rect 18704 -810 18738 -794
rect 18704 -1402 18738 -1386
rect 19722 -810 19756 -794
rect 19722 -1402 19756 -1386
rect 20740 -810 20774 -794
rect 20740 -1402 20774 -1386
rect 21758 -810 21792 -794
rect 21758 -1402 21792 -1386
rect 22776 -810 22810 -794
rect 22776 -1402 22810 -1386
rect 6720 -1479 6736 -1445
rect 7292 -1479 7308 -1445
rect 7738 -1479 7754 -1445
rect 8310 -1479 8326 -1445
rect 8756 -1479 8772 -1445
rect 9328 -1479 9344 -1445
rect 9774 -1479 9790 -1445
rect 10346 -1479 10362 -1445
rect 10792 -1479 10808 -1445
rect 11364 -1479 11380 -1445
rect 11810 -1479 11826 -1445
rect 12382 -1479 12398 -1445
rect 12828 -1479 12844 -1445
rect 13400 -1479 13416 -1445
rect 13846 -1479 13862 -1445
rect 14418 -1479 14434 -1445
rect 14864 -1479 14880 -1445
rect 15436 -1479 15452 -1445
rect 15882 -1479 15898 -1445
rect 16454 -1479 16470 -1445
rect 16900 -1479 16916 -1445
rect 17472 -1479 17488 -1445
rect 17918 -1479 17934 -1445
rect 18490 -1479 18506 -1445
rect 18936 -1479 18952 -1445
rect 19508 -1479 19524 -1445
rect 19954 -1479 19970 -1445
rect 20526 -1479 20542 -1445
rect 20972 -1479 20988 -1445
rect 21544 -1479 21560 -1445
rect 21990 -1479 22006 -1445
rect 22562 -1479 22578 -1445
rect 6968 -1890 7058 -1860
rect 6968 -1924 6996 -1890
rect 7030 -1924 7058 -1890
rect 6968 -1952 7058 -1924
rect 7986 -1890 8076 -1860
rect 7986 -1924 8014 -1890
rect 8048 -1924 8076 -1890
rect 7986 -1952 8076 -1924
rect 9004 -1890 9094 -1860
rect 9004 -1924 9032 -1890
rect 9066 -1924 9094 -1890
rect 9004 -1952 9094 -1924
rect 10022 -1890 10112 -1860
rect 10022 -1924 10050 -1890
rect 10084 -1924 10112 -1890
rect 10022 -1952 10112 -1924
rect 11040 -1890 11130 -1860
rect 11040 -1924 11068 -1890
rect 11102 -1924 11130 -1890
rect 11040 -1952 11130 -1924
rect 12058 -1890 12148 -1860
rect 12058 -1924 12086 -1890
rect 12120 -1924 12148 -1890
rect 12058 -1952 12148 -1924
rect 13076 -1890 13166 -1860
rect 13076 -1924 13104 -1890
rect 13138 -1924 13166 -1890
rect 13076 -1952 13166 -1924
rect 14094 -1890 14184 -1860
rect 14094 -1924 14122 -1890
rect 14156 -1924 14184 -1890
rect 14094 -1952 14184 -1924
rect 15112 -1890 15202 -1860
rect 15112 -1924 15140 -1890
rect 15174 -1924 15202 -1890
rect 15112 -1952 15202 -1924
rect 16130 -1890 16220 -1860
rect 16130 -1924 16158 -1890
rect 16192 -1924 16220 -1890
rect 16130 -1952 16220 -1924
rect 17148 -1890 17238 -1860
rect 17148 -1924 17176 -1890
rect 17210 -1924 17238 -1890
rect 17148 -1952 17238 -1924
rect 18166 -1890 18256 -1860
rect 18166 -1924 18194 -1890
rect 18228 -1924 18256 -1890
rect 18166 -1952 18256 -1924
rect 19184 -1890 19274 -1860
rect 19184 -1924 19212 -1890
rect 19246 -1924 19274 -1890
rect 19184 -1952 19274 -1924
rect 20202 -1890 20292 -1860
rect 20202 -1924 20230 -1890
rect 20264 -1924 20292 -1890
rect 20202 -1952 20292 -1924
rect 21220 -1890 21310 -1860
rect 21220 -1924 21248 -1890
rect 21282 -1924 21310 -1890
rect 21220 -1952 21310 -1924
rect 22238 -1890 22328 -1860
rect 22238 -1924 22266 -1890
rect 22300 -1924 22328 -1890
rect 22238 -1952 22328 -1924
rect 7914 -2389 7930 -2355
rect 8486 -2389 8502 -2355
rect 8932 -2389 8948 -2355
rect 9504 -2389 9520 -2355
rect 9950 -2389 9966 -2355
rect 10522 -2389 10538 -2355
rect 10968 -2389 10984 -2355
rect 11540 -2389 11556 -2355
rect 11986 -2389 12002 -2355
rect 12558 -2389 12574 -2355
rect 13004 -2389 13020 -2355
rect 13576 -2389 13592 -2355
rect 14022 -2389 14038 -2355
rect 14594 -2389 14610 -2355
rect 15040 -2389 15056 -2355
rect 15612 -2389 15628 -2355
rect 16058 -2389 16074 -2355
rect 16630 -2389 16646 -2355
rect 17076 -2389 17092 -2355
rect 17648 -2389 17664 -2355
rect 18094 -2389 18110 -2355
rect 18666 -2389 18682 -2355
rect 19112 -2389 19128 -2355
rect 19684 -2389 19700 -2355
rect 20130 -2389 20146 -2355
rect 20702 -2389 20718 -2355
rect 21148 -2389 21164 -2355
rect 21720 -2389 21736 -2355
rect 7682 -2448 7716 -2432
rect 7682 -3040 7716 -3024
rect 8700 -2448 8734 -2432
rect 8700 -3040 8734 -3024
rect 9718 -2448 9752 -2432
rect 9718 -3040 9752 -3024
rect 10736 -2448 10770 -2432
rect 10736 -3040 10770 -3024
rect 11754 -2448 11788 -2432
rect 11754 -3040 11788 -3024
rect 12772 -2448 12806 -2432
rect 12772 -3040 12806 -3024
rect 13790 -2448 13824 -2432
rect 13790 -3040 13824 -3024
rect 14808 -2448 14842 -2432
rect 14808 -3040 14842 -3024
rect 15826 -2448 15860 -2432
rect 15826 -3040 15860 -3024
rect 16844 -2448 16878 -2432
rect 16844 -3040 16878 -3024
rect 17862 -2448 17896 -2432
rect 17862 -3040 17896 -3024
rect 18880 -2448 18914 -2432
rect 18880 -3040 18914 -3024
rect 19898 -2448 19932 -2432
rect 19898 -3040 19932 -3024
rect 20916 -2448 20950 -2432
rect 20916 -3040 20950 -3024
rect 21934 -2448 21968 -2432
rect 21934 -3040 21968 -3024
rect 7914 -3117 7930 -3083
rect 8486 -3117 8502 -3083
rect 8932 -3117 8948 -3083
rect 9504 -3117 9520 -3083
rect 9950 -3117 9966 -3083
rect 10522 -3117 10538 -3083
rect 10968 -3117 10984 -3083
rect 11540 -3117 11556 -3083
rect 11986 -3117 12002 -3083
rect 12558 -3117 12574 -3083
rect 13004 -3117 13020 -3083
rect 13576 -3117 13592 -3083
rect 14022 -3117 14038 -3083
rect 14594 -3117 14610 -3083
rect 15040 -3117 15056 -3083
rect 15612 -3117 15628 -3083
rect 16058 -3117 16074 -3083
rect 16630 -3117 16646 -3083
rect 17076 -3117 17092 -3083
rect 17648 -3117 17664 -3083
rect 18094 -3117 18110 -3083
rect 18666 -3117 18682 -3083
rect 19112 -3117 19128 -3083
rect 19684 -3117 19700 -3083
rect 20130 -3117 20146 -3083
rect 20702 -3117 20718 -3083
rect 21148 -3117 21164 -3083
rect 21720 -3117 21736 -3083
rect 7656 -3238 7746 -3208
rect 7656 -3272 7684 -3238
rect 7718 -3272 7746 -3238
rect 7656 -3300 7746 -3272
rect 8674 -3238 8764 -3208
rect 8674 -3272 8702 -3238
rect 8736 -3272 8764 -3238
rect 8674 -3300 8764 -3272
rect 9692 -3238 9782 -3208
rect 9692 -3272 9720 -3238
rect 9754 -3272 9782 -3238
rect 9692 -3300 9782 -3272
rect 10710 -3238 10800 -3208
rect 10710 -3272 10738 -3238
rect 10772 -3272 10800 -3238
rect 10710 -3300 10800 -3272
rect 11728 -3238 11818 -3208
rect 11728 -3272 11756 -3238
rect 11790 -3272 11818 -3238
rect 11728 -3300 11818 -3272
rect 12746 -3238 12836 -3208
rect 12746 -3272 12774 -3238
rect 12808 -3272 12836 -3238
rect 12746 -3300 12836 -3272
rect 13764 -3238 13854 -3208
rect 13764 -3272 13792 -3238
rect 13826 -3272 13854 -3238
rect 13764 -3300 13854 -3272
rect 14782 -3238 14872 -3208
rect 14782 -3272 14810 -3238
rect 14844 -3272 14872 -3238
rect 14782 -3300 14872 -3272
rect 15800 -3238 15890 -3208
rect 15800 -3272 15828 -3238
rect 15862 -3272 15890 -3238
rect 15800 -3300 15890 -3272
rect 16818 -3238 16908 -3208
rect 16818 -3272 16846 -3238
rect 16880 -3272 16908 -3238
rect 16818 -3300 16908 -3272
rect 17836 -3238 17926 -3208
rect 17836 -3272 17864 -3238
rect 17898 -3272 17926 -3238
rect 17836 -3300 17926 -3272
rect 18854 -3238 18944 -3208
rect 18854 -3272 18882 -3238
rect 18916 -3272 18944 -3238
rect 18854 -3300 18944 -3272
rect 19872 -3238 19962 -3208
rect 19872 -3272 19900 -3238
rect 19934 -3272 19962 -3238
rect 19872 -3300 19962 -3272
rect 20890 -3238 20980 -3208
rect 20890 -3272 20918 -3238
rect 20952 -3272 20980 -3238
rect 20890 -3300 20980 -3272
rect 21908 -3238 21998 -3208
rect 21908 -3272 21936 -3238
rect 21970 -3272 21998 -3238
rect 21908 -3300 21998 -3272
rect 7914 -3421 7930 -3387
rect 8486 -3421 8502 -3387
rect 8932 -3421 8948 -3387
rect 9504 -3421 9520 -3387
rect 9950 -3421 9966 -3387
rect 10522 -3421 10538 -3387
rect 10968 -3421 10984 -3387
rect 11540 -3421 11556 -3387
rect 11986 -3421 12002 -3387
rect 12558 -3421 12574 -3387
rect 13004 -3421 13020 -3387
rect 13576 -3421 13592 -3387
rect 14022 -3421 14038 -3387
rect 14594 -3421 14610 -3387
rect 15040 -3421 15056 -3387
rect 15612 -3421 15628 -3387
rect 16058 -3421 16074 -3387
rect 16630 -3421 16646 -3387
rect 17076 -3421 17092 -3387
rect 17648 -3421 17664 -3387
rect 18094 -3421 18110 -3387
rect 18666 -3421 18682 -3387
rect 19112 -3421 19128 -3387
rect 19684 -3421 19700 -3387
rect 20130 -3421 20146 -3387
rect 20702 -3421 20718 -3387
rect 21148 -3421 21164 -3387
rect 21720 -3421 21736 -3387
rect 7682 -3480 7716 -3464
rect 7682 -4072 7716 -4056
rect 8700 -3480 8734 -3464
rect 8700 -4072 8734 -4056
rect 9718 -3480 9752 -3464
rect 9718 -4072 9752 -4056
rect 10736 -3480 10770 -3464
rect 10736 -4072 10770 -4056
rect 11754 -3480 11788 -3464
rect 11754 -4072 11788 -4056
rect 12772 -3480 12806 -3464
rect 12772 -4072 12806 -4056
rect 13790 -3480 13824 -3464
rect 13790 -4072 13824 -4056
rect 14808 -3480 14842 -3464
rect 14808 -4072 14842 -4056
rect 15826 -3480 15860 -3464
rect 15826 -4072 15860 -4056
rect 16844 -3480 16878 -3464
rect 16844 -4072 16878 -4056
rect 17862 -3480 17896 -3464
rect 17862 -4072 17896 -4056
rect 18880 -3480 18914 -3464
rect 18880 -4072 18914 -4056
rect 19898 -3480 19932 -3464
rect 19898 -4072 19932 -4056
rect 20916 -3480 20950 -3464
rect 20916 -4072 20950 -4056
rect 21934 -3480 21968 -3464
rect 21934 -4072 21968 -4056
rect 7914 -4149 7930 -4115
rect 8486 -4149 8502 -4115
rect 8932 -4149 8948 -4115
rect 9504 -4149 9520 -4115
rect 9950 -4149 9966 -4115
rect 10522 -4149 10538 -4115
rect 10968 -4149 10984 -4115
rect 11540 -4149 11556 -4115
rect 11986 -4149 12002 -4115
rect 12558 -4149 12574 -4115
rect 13004 -4149 13020 -4115
rect 13576 -4149 13592 -4115
rect 14022 -4149 14038 -4115
rect 14594 -4149 14610 -4115
rect 15040 -4149 15056 -4115
rect 15612 -4149 15628 -4115
rect 16058 -4149 16074 -4115
rect 16630 -4149 16646 -4115
rect 17076 -4149 17092 -4115
rect 17648 -4149 17664 -4115
rect 18094 -4149 18110 -4115
rect 18666 -4149 18682 -4115
rect 19112 -4149 19128 -4115
rect 19684 -4149 19700 -4115
rect 20130 -4149 20146 -4115
rect 20702 -4149 20718 -4115
rect 21148 -4149 21164 -4115
rect 21720 -4149 21736 -4115
rect 7262 -4516 7352 -4486
rect 7262 -4550 7290 -4516
rect 7324 -4550 7352 -4516
rect 7262 -4578 7352 -4550
rect 8280 -4516 8370 -4486
rect 8280 -4550 8308 -4516
rect 8342 -4550 8370 -4516
rect 8280 -4578 8370 -4550
rect 9298 -4516 9388 -4486
rect 9298 -4550 9326 -4516
rect 9360 -4550 9388 -4516
rect 9298 -4578 9388 -4550
rect 10316 -4516 10406 -4486
rect 10316 -4550 10344 -4516
rect 10378 -4550 10406 -4516
rect 10316 -4578 10406 -4550
rect 11334 -4516 11424 -4486
rect 11334 -4550 11362 -4516
rect 11396 -4550 11424 -4516
rect 11334 -4578 11424 -4550
rect 12352 -4516 12442 -4486
rect 12352 -4550 12380 -4516
rect 12414 -4550 12442 -4516
rect 12352 -4578 12442 -4550
rect 13370 -4516 13460 -4486
rect 13370 -4550 13398 -4516
rect 13432 -4550 13460 -4516
rect 13370 -4578 13460 -4550
rect 14388 -4516 14478 -4486
rect 14388 -4550 14416 -4516
rect 14450 -4550 14478 -4516
rect 14388 -4578 14478 -4550
rect 15406 -4516 15496 -4486
rect 15406 -4550 15434 -4516
rect 15468 -4550 15496 -4516
rect 15406 -4578 15496 -4550
rect 16424 -4516 16514 -4486
rect 16424 -4550 16452 -4516
rect 16486 -4550 16514 -4516
rect 16424 -4578 16514 -4550
rect 17442 -4516 17532 -4486
rect 17442 -4550 17470 -4516
rect 17504 -4550 17532 -4516
rect 17442 -4578 17532 -4550
rect 18460 -4516 18550 -4486
rect 18460 -4550 18488 -4516
rect 18522 -4550 18550 -4516
rect 18460 -4578 18550 -4550
rect 19478 -4516 19568 -4486
rect 19478 -4550 19506 -4516
rect 19540 -4550 19568 -4516
rect 19478 -4578 19568 -4550
rect 20496 -4516 20586 -4486
rect 20496 -4550 20524 -4516
rect 20558 -4550 20586 -4516
rect 20496 -4578 20586 -4550
rect 21514 -4516 21604 -4486
rect 21514 -4550 21542 -4516
rect 21576 -4550 21604 -4516
rect 21514 -4578 21604 -4550
rect 22532 -4516 22622 -4486
rect 22532 -4550 22560 -4516
rect 22594 -4550 22622 -4516
rect 22532 -4578 22622 -4550
rect 2664 -4826 2754 -4796
rect 2664 -4860 2692 -4826
rect 2726 -4860 2754 -4826
rect 2664 -4888 2754 -4860
rect 3682 -4826 3772 -4796
rect 3682 -4860 3710 -4826
rect 3744 -4860 3772 -4826
rect 3682 -4888 3772 -4860
rect 4700 -4826 4790 -4796
rect 4700 -4860 4728 -4826
rect 4762 -4860 4790 -4826
rect 4700 -4888 4790 -4860
rect 5718 -4826 5808 -4796
rect 5718 -4860 5746 -4826
rect 5780 -4860 5808 -4826
rect 5718 -4888 5808 -4860
rect 7706 -5025 7722 -4991
rect 8278 -5025 8294 -4991
rect 8724 -5025 8740 -4991
rect 9296 -5025 9312 -4991
rect 9742 -5025 9758 -4991
rect 10314 -5025 10330 -4991
rect 10760 -5025 10776 -4991
rect 11332 -5025 11348 -4991
rect 11778 -5025 11794 -4991
rect 12350 -5025 12366 -4991
rect 12796 -5025 12812 -4991
rect 13368 -5025 13384 -4991
rect 13814 -5025 13830 -4991
rect 14386 -5025 14402 -4991
rect 14832 -5025 14848 -4991
rect 15404 -5025 15420 -4991
rect 15850 -5025 15866 -4991
rect 16422 -5025 16438 -4991
rect 16868 -5025 16884 -4991
rect 17440 -5025 17456 -4991
rect 17886 -5025 17902 -4991
rect 18458 -5025 18474 -4991
rect 18904 -5025 18920 -4991
rect 19476 -5025 19492 -4991
rect 19922 -5025 19938 -4991
rect 20494 -5025 20510 -4991
rect 20940 -5025 20956 -4991
rect 21512 -5025 21528 -4991
rect 21958 -5025 21974 -4991
rect 22530 -5025 22546 -4991
rect 7474 -5084 7508 -5068
rect 2402 -5129 2418 -5095
rect 2974 -5129 2990 -5095
rect 3420 -5129 3436 -5095
rect 3992 -5129 4008 -5095
rect 4438 -5129 4454 -5095
rect 5010 -5129 5026 -5095
rect 5456 -5129 5472 -5095
rect 6028 -5129 6044 -5095
rect 2170 -5188 2204 -5172
rect 2170 -5780 2204 -5764
rect 3188 -5188 3222 -5172
rect 3188 -5780 3222 -5764
rect 4206 -5188 4240 -5172
rect 4206 -5780 4240 -5764
rect 5224 -5188 5258 -5172
rect 5224 -5780 5258 -5764
rect 6242 -5188 6276 -5172
rect 7474 -5676 7508 -5660
rect 8492 -5084 8526 -5068
rect 8492 -5676 8526 -5660
rect 9510 -5084 9544 -5068
rect 9510 -5676 9544 -5660
rect 10528 -5084 10562 -5068
rect 10528 -5676 10562 -5660
rect 11546 -5084 11580 -5068
rect 11546 -5676 11580 -5660
rect 12564 -5084 12598 -5068
rect 12564 -5676 12598 -5660
rect 13582 -5084 13616 -5068
rect 13582 -5676 13616 -5660
rect 14600 -5084 14634 -5068
rect 14600 -5676 14634 -5660
rect 15618 -5084 15652 -5068
rect 15618 -5676 15652 -5660
rect 16636 -5084 16670 -5068
rect 16636 -5676 16670 -5660
rect 17654 -5084 17688 -5068
rect 17654 -5676 17688 -5660
rect 18672 -5084 18706 -5068
rect 18672 -5676 18706 -5660
rect 19690 -5084 19724 -5068
rect 19690 -5676 19724 -5660
rect 20708 -5084 20742 -5068
rect 20708 -5676 20742 -5660
rect 21726 -5084 21760 -5068
rect 21726 -5676 21760 -5660
rect 22744 -5084 22778 -5068
rect 22744 -5676 22778 -5660
rect 7706 -5753 7722 -5719
rect 8278 -5753 8294 -5719
rect 8724 -5753 8740 -5719
rect 9296 -5753 9312 -5719
rect 9742 -5753 9758 -5719
rect 10314 -5753 10330 -5719
rect 10760 -5753 10776 -5719
rect 11332 -5753 11348 -5719
rect 11778 -5753 11794 -5719
rect 12350 -5753 12366 -5719
rect 12796 -5753 12812 -5719
rect 13368 -5753 13384 -5719
rect 13814 -5753 13830 -5719
rect 14386 -5753 14402 -5719
rect 14832 -5753 14848 -5719
rect 15404 -5753 15420 -5719
rect 15850 -5753 15866 -5719
rect 16422 -5753 16438 -5719
rect 16868 -5753 16884 -5719
rect 17440 -5753 17456 -5719
rect 17886 -5753 17902 -5719
rect 18458 -5753 18474 -5719
rect 18904 -5753 18920 -5719
rect 19476 -5753 19492 -5719
rect 19922 -5753 19938 -5719
rect 20494 -5753 20510 -5719
rect 20940 -5753 20956 -5719
rect 21512 -5753 21528 -5719
rect 21958 -5753 21974 -5719
rect 22530 -5753 22546 -5719
rect 6242 -5780 6276 -5764
rect 2402 -5857 2418 -5823
rect 2974 -5857 2990 -5823
rect 3420 -5857 3436 -5823
rect 3992 -5857 4008 -5823
rect 4438 -5857 4454 -5823
rect 5010 -5857 5026 -5823
rect 5456 -5857 5472 -5823
rect 6028 -5857 6044 -5823
rect 2140 -5980 2230 -5950
rect 2140 -6014 2168 -5980
rect 2202 -6014 2230 -5980
rect 2140 -6042 2230 -6014
rect 3158 -5980 3248 -5950
rect 3158 -6014 3186 -5980
rect 3220 -6014 3248 -5980
rect 3158 -6042 3248 -6014
rect 4176 -5980 4266 -5950
rect 4176 -6014 4204 -5980
rect 4238 -6014 4266 -5980
rect 4176 -6042 4266 -6014
rect 5194 -5980 5284 -5950
rect 5194 -6014 5222 -5980
rect 5256 -6014 5284 -5980
rect 5194 -6042 5284 -6014
rect 7352 -5964 7442 -5934
rect 7352 -5998 7380 -5964
rect 7414 -5998 7442 -5964
rect 7352 -6026 7442 -5998
rect 8370 -5964 8460 -5934
rect 8370 -5998 8398 -5964
rect 8432 -5998 8460 -5964
rect 8370 -6026 8460 -5998
rect 9388 -5964 9478 -5934
rect 9388 -5998 9416 -5964
rect 9450 -5998 9478 -5964
rect 9388 -6026 9478 -5998
rect 10406 -5964 10496 -5934
rect 10406 -5998 10434 -5964
rect 10468 -5998 10496 -5964
rect 10406 -6026 10496 -5998
rect 11424 -5964 11514 -5934
rect 11424 -5998 11452 -5964
rect 11486 -5998 11514 -5964
rect 11424 -6026 11514 -5998
rect 12442 -5964 12532 -5934
rect 12442 -5998 12470 -5964
rect 12504 -5998 12532 -5964
rect 12442 -6026 12532 -5998
rect 13460 -5964 13550 -5934
rect 13460 -5998 13488 -5964
rect 13522 -5998 13550 -5964
rect 13460 -6026 13550 -5998
rect 14478 -5964 14568 -5934
rect 14478 -5998 14506 -5964
rect 14540 -5998 14568 -5964
rect 14478 -6026 14568 -5998
rect 15496 -5964 15586 -5934
rect 15496 -5998 15524 -5964
rect 15558 -5998 15586 -5964
rect 15496 -6026 15586 -5998
rect 16514 -5964 16604 -5934
rect 16514 -5998 16542 -5964
rect 16576 -5998 16604 -5964
rect 16514 -6026 16604 -5998
rect 17532 -5964 17622 -5934
rect 17532 -5998 17560 -5964
rect 17594 -5998 17622 -5964
rect 17532 -6026 17622 -5998
rect 18550 -5964 18640 -5934
rect 18550 -5998 18578 -5964
rect 18612 -5998 18640 -5964
rect 18550 -6026 18640 -5998
rect 19568 -5964 19658 -5934
rect 19568 -5998 19596 -5964
rect 19630 -5998 19658 -5964
rect 19568 -6026 19658 -5998
rect 20586 -5964 20676 -5934
rect 20586 -5998 20614 -5964
rect 20648 -5998 20676 -5964
rect 20586 -6026 20676 -5998
rect 21604 -5964 21694 -5934
rect 21604 -5998 21632 -5964
rect 21666 -5998 21694 -5964
rect 21604 -6026 21694 -5998
rect 22622 -5964 22712 -5934
rect 22622 -5998 22650 -5964
rect 22684 -5998 22712 -5964
rect 22622 -6026 22712 -5998
rect 2402 -6161 2418 -6127
rect 2974 -6161 2990 -6127
rect 3420 -6161 3436 -6127
rect 3992 -6161 4008 -6127
rect 4438 -6161 4454 -6127
rect 5010 -6161 5026 -6127
rect 5456 -6161 5472 -6127
rect 6028 -6161 6044 -6127
rect 2170 -6220 2204 -6204
rect 2170 -6812 2204 -6796
rect 3188 -6220 3222 -6204
rect 3188 -6812 3222 -6796
rect 4206 -6220 4240 -6204
rect 4206 -6812 4240 -6796
rect 5224 -6220 5258 -6204
rect 5224 -6812 5258 -6796
rect 6242 -6220 6276 -6204
rect 7706 -6281 7722 -6247
rect 8278 -6281 8294 -6247
rect 8724 -6281 8740 -6247
rect 9296 -6281 9312 -6247
rect 9742 -6281 9758 -6247
rect 10314 -6281 10330 -6247
rect 10760 -6281 10776 -6247
rect 11332 -6281 11348 -6247
rect 11778 -6281 11794 -6247
rect 12350 -6281 12366 -6247
rect 12796 -6281 12812 -6247
rect 13368 -6281 13384 -6247
rect 13814 -6281 13830 -6247
rect 14386 -6281 14402 -6247
rect 14832 -6281 14848 -6247
rect 15404 -6281 15420 -6247
rect 15850 -6281 15866 -6247
rect 16422 -6281 16438 -6247
rect 16868 -6281 16884 -6247
rect 17440 -6281 17456 -6247
rect 17886 -6281 17902 -6247
rect 18458 -6281 18474 -6247
rect 18904 -6281 18920 -6247
rect 19476 -6281 19492 -6247
rect 19922 -6281 19938 -6247
rect 20494 -6281 20510 -6247
rect 20940 -6281 20956 -6247
rect 21512 -6281 21528 -6247
rect 21958 -6281 21974 -6247
rect 22530 -6281 22546 -6247
rect 6242 -6812 6276 -6796
rect 7474 -6340 7508 -6324
rect 2402 -6889 2418 -6855
rect 2974 -6889 2990 -6855
rect 3420 -6889 3436 -6855
rect 3992 -6889 4008 -6855
rect 4438 -6889 4454 -6855
rect 5010 -6889 5026 -6855
rect 5456 -6889 5472 -6855
rect 6028 -6889 6044 -6855
rect 7474 -6932 7508 -6916
rect 8492 -6340 8526 -6324
rect 8492 -6932 8526 -6916
rect 9510 -6340 9544 -6324
rect 9510 -6932 9544 -6916
rect 10528 -6340 10562 -6324
rect 10528 -6932 10562 -6916
rect 11546 -6340 11580 -6324
rect 11546 -6932 11580 -6916
rect 12564 -6340 12598 -6324
rect 12564 -6932 12598 -6916
rect 13582 -6340 13616 -6324
rect 13582 -6932 13616 -6916
rect 14600 -6340 14634 -6324
rect 14600 -6932 14634 -6916
rect 15618 -6340 15652 -6324
rect 15618 -6932 15652 -6916
rect 16636 -6340 16670 -6324
rect 16636 -6932 16670 -6916
rect 17654 -6340 17688 -6324
rect 17654 -6932 17688 -6916
rect 18672 -6340 18706 -6324
rect 18672 -6932 18706 -6916
rect 19690 -6340 19724 -6324
rect 19690 -6932 19724 -6916
rect 20708 -6340 20742 -6324
rect 20708 -6932 20742 -6916
rect 21726 -6340 21760 -6324
rect 21726 -6932 21760 -6916
rect 22744 -6340 22778 -6324
rect 22744 -6932 22778 -6916
rect 2150 -7008 2240 -6978
rect 2150 -7042 2178 -7008
rect 2212 -7042 2240 -7008
rect 2150 -7070 2240 -7042
rect 3168 -7008 3258 -6978
rect 3168 -7042 3196 -7008
rect 3230 -7042 3258 -7008
rect 3168 -7070 3258 -7042
rect 4186 -7008 4276 -6978
rect 4186 -7042 4214 -7008
rect 4248 -7042 4276 -7008
rect 4186 -7070 4276 -7042
rect 5204 -7008 5294 -6978
rect 5204 -7042 5232 -7008
rect 5266 -7042 5294 -7008
rect 7706 -7009 7722 -6975
rect 8278 -7009 8294 -6975
rect 8724 -7009 8740 -6975
rect 9296 -7009 9312 -6975
rect 9742 -7009 9758 -6975
rect 10314 -7009 10330 -6975
rect 10760 -7009 10776 -6975
rect 11332 -7009 11348 -6975
rect 11778 -7009 11794 -6975
rect 12350 -7009 12366 -6975
rect 12796 -7009 12812 -6975
rect 13368 -7009 13384 -6975
rect 13814 -7009 13830 -6975
rect 14386 -7009 14402 -6975
rect 14832 -7009 14848 -6975
rect 15404 -7009 15420 -6975
rect 15850 -7009 15866 -6975
rect 16422 -7009 16438 -6975
rect 16868 -7009 16884 -6975
rect 17440 -7009 17456 -6975
rect 17886 -7009 17902 -6975
rect 18458 -7009 18474 -6975
rect 18904 -7009 18920 -6975
rect 19476 -7009 19492 -6975
rect 19922 -7009 19938 -6975
rect 20494 -7009 20510 -6975
rect 20940 -7009 20956 -6975
rect 21512 -7009 21528 -6975
rect 21958 -7009 21974 -6975
rect 22530 -7009 22546 -6975
rect 5204 -7070 5294 -7042
rect 2402 -7193 2418 -7159
rect 2974 -7193 2990 -7159
rect 3420 -7193 3436 -7159
rect 3992 -7193 4008 -7159
rect 4438 -7193 4454 -7159
rect 5010 -7193 5026 -7159
rect 5456 -7193 5472 -7159
rect 6028 -7193 6044 -7159
rect 7376 -7232 7466 -7202
rect 2170 -7252 2204 -7236
rect 2170 -7844 2204 -7828
rect 3188 -7252 3222 -7236
rect 3188 -7844 3222 -7828
rect 4206 -7252 4240 -7236
rect 4206 -7844 4240 -7828
rect 5224 -7252 5258 -7236
rect 5224 -7844 5258 -7828
rect 6242 -7252 6276 -7236
rect 7376 -7266 7404 -7232
rect 7438 -7266 7466 -7232
rect 7376 -7294 7466 -7266
rect 8394 -7232 8484 -7202
rect 8394 -7266 8422 -7232
rect 8456 -7266 8484 -7232
rect 8394 -7294 8484 -7266
rect 9412 -7232 9502 -7202
rect 9412 -7266 9440 -7232
rect 9474 -7266 9502 -7232
rect 9412 -7294 9502 -7266
rect 10430 -7232 10520 -7202
rect 10430 -7266 10458 -7232
rect 10492 -7266 10520 -7232
rect 10430 -7294 10520 -7266
rect 11448 -7232 11538 -7202
rect 11448 -7266 11476 -7232
rect 11510 -7266 11538 -7232
rect 11448 -7294 11538 -7266
rect 12466 -7232 12556 -7202
rect 12466 -7266 12494 -7232
rect 12528 -7266 12556 -7232
rect 12466 -7294 12556 -7266
rect 13484 -7232 13574 -7202
rect 13484 -7266 13512 -7232
rect 13546 -7266 13574 -7232
rect 13484 -7294 13574 -7266
rect 14502 -7232 14592 -7202
rect 14502 -7266 14530 -7232
rect 14564 -7266 14592 -7232
rect 14502 -7294 14592 -7266
rect 15520 -7232 15610 -7202
rect 15520 -7266 15548 -7232
rect 15582 -7266 15610 -7232
rect 15520 -7294 15610 -7266
rect 16538 -7232 16628 -7202
rect 16538 -7266 16566 -7232
rect 16600 -7266 16628 -7232
rect 16538 -7294 16628 -7266
rect 17556 -7232 17646 -7202
rect 17556 -7266 17584 -7232
rect 17618 -7266 17646 -7232
rect 17556 -7294 17646 -7266
rect 18574 -7232 18664 -7202
rect 18574 -7266 18602 -7232
rect 18636 -7266 18664 -7232
rect 18574 -7294 18664 -7266
rect 19592 -7232 19682 -7202
rect 19592 -7266 19620 -7232
rect 19654 -7266 19682 -7232
rect 19592 -7294 19682 -7266
rect 20610 -7232 20700 -7202
rect 20610 -7266 20638 -7232
rect 20672 -7266 20700 -7232
rect 20610 -7294 20700 -7266
rect 21628 -7232 21718 -7202
rect 21628 -7266 21656 -7232
rect 21690 -7266 21718 -7232
rect 21628 -7294 21718 -7266
rect 22646 -7232 22736 -7202
rect 22646 -7266 22674 -7232
rect 22708 -7266 22736 -7232
rect 22646 -7294 22736 -7266
rect 7706 -7537 7722 -7503
rect 8278 -7537 8294 -7503
rect 8724 -7537 8740 -7503
rect 9296 -7537 9312 -7503
rect 9742 -7537 9758 -7503
rect 10314 -7537 10330 -7503
rect 10760 -7537 10776 -7503
rect 11332 -7537 11348 -7503
rect 11778 -7537 11794 -7503
rect 12350 -7537 12366 -7503
rect 12796 -7537 12812 -7503
rect 13368 -7537 13384 -7503
rect 13814 -7537 13830 -7503
rect 14386 -7537 14402 -7503
rect 14832 -7537 14848 -7503
rect 15404 -7537 15420 -7503
rect 15850 -7537 15866 -7503
rect 16422 -7537 16438 -7503
rect 16868 -7537 16884 -7503
rect 17440 -7537 17456 -7503
rect 17886 -7537 17902 -7503
rect 18458 -7537 18474 -7503
rect 18904 -7537 18920 -7503
rect 19476 -7537 19492 -7503
rect 19922 -7537 19938 -7503
rect 20494 -7537 20510 -7503
rect 20940 -7537 20956 -7503
rect 21512 -7537 21528 -7503
rect 21958 -7537 21974 -7503
rect 22530 -7537 22546 -7503
rect 6242 -7844 6276 -7828
rect 7474 -7596 7508 -7580
rect 2402 -7921 2418 -7887
rect 2974 -7921 2990 -7887
rect 3420 -7921 3436 -7887
rect 3992 -7921 4008 -7887
rect 4438 -7921 4454 -7887
rect 5010 -7921 5026 -7887
rect 5456 -7921 5472 -7887
rect 6028 -7921 6044 -7887
rect 2140 -8036 2230 -8006
rect 2140 -8070 2168 -8036
rect 2202 -8070 2230 -8036
rect 2140 -8098 2230 -8070
rect 3158 -8036 3248 -8006
rect 3158 -8070 3186 -8036
rect 3220 -8070 3248 -8036
rect 3158 -8098 3248 -8070
rect 4176 -8036 4266 -8006
rect 4176 -8070 4204 -8036
rect 4238 -8070 4266 -8036
rect 4176 -8098 4266 -8070
rect 5194 -8036 5284 -8006
rect 5194 -8070 5222 -8036
rect 5256 -8070 5284 -8036
rect 5194 -8098 5284 -8070
rect 7474 -8188 7508 -8172
rect 8492 -7596 8526 -7580
rect 8492 -8188 8526 -8172
rect 9510 -7596 9544 -7580
rect 9510 -8188 9544 -8172
rect 10528 -7596 10562 -7580
rect 10528 -8188 10562 -8172
rect 11546 -7596 11580 -7580
rect 11546 -8188 11580 -8172
rect 12564 -7596 12598 -7580
rect 12564 -8188 12598 -8172
rect 13582 -7596 13616 -7580
rect 13582 -8188 13616 -8172
rect 14600 -7596 14634 -7580
rect 14600 -8188 14634 -8172
rect 15618 -7596 15652 -7580
rect 15618 -8188 15652 -8172
rect 16636 -7596 16670 -7580
rect 16636 -8188 16670 -8172
rect 17654 -7596 17688 -7580
rect 17654 -8188 17688 -8172
rect 18672 -7596 18706 -7580
rect 18672 -8188 18706 -8172
rect 19690 -7596 19724 -7580
rect 19690 -8188 19724 -8172
rect 20708 -7596 20742 -7580
rect 20708 -8188 20742 -8172
rect 21726 -7596 21760 -7580
rect 21726 -8188 21760 -8172
rect 22744 -7596 22778 -7580
rect 22744 -8188 22778 -8172
rect 2402 -8225 2418 -8191
rect 2974 -8225 2990 -8191
rect 3420 -8225 3436 -8191
rect 3992 -8225 4008 -8191
rect 4438 -8225 4454 -8191
rect 5010 -8225 5026 -8191
rect 5456 -8225 5472 -8191
rect 6028 -8225 6044 -8191
rect 7706 -8265 7722 -8231
rect 8278 -8265 8294 -8231
rect 8724 -8265 8740 -8231
rect 9296 -8265 9312 -8231
rect 9742 -8265 9758 -8231
rect 10314 -8265 10330 -8231
rect 10760 -8265 10776 -8231
rect 11332 -8265 11348 -8231
rect 11778 -8265 11794 -8231
rect 12350 -8265 12366 -8231
rect 12796 -8265 12812 -8231
rect 13368 -8265 13384 -8231
rect 13814 -8265 13830 -8231
rect 14386 -8265 14402 -8231
rect 14832 -8265 14848 -8231
rect 15404 -8265 15420 -8231
rect 15850 -8265 15866 -8231
rect 16422 -8265 16438 -8231
rect 16868 -8265 16884 -8231
rect 17440 -8265 17456 -8231
rect 17886 -8265 17902 -8231
rect 18458 -8265 18474 -8231
rect 18904 -8265 18920 -8231
rect 19476 -8265 19492 -8231
rect 19922 -8265 19938 -8231
rect 20494 -8265 20510 -8231
rect 20940 -8265 20956 -8231
rect 21512 -8265 21528 -8231
rect 21958 -8265 21974 -8231
rect 22530 -8265 22546 -8231
rect 2170 -8284 2204 -8268
rect 2170 -8876 2204 -8860
rect 3188 -8284 3222 -8268
rect 3188 -8876 3222 -8860
rect 4206 -8284 4240 -8268
rect 4206 -8876 4240 -8860
rect 5224 -8284 5258 -8268
rect 5224 -8876 5258 -8860
rect 6242 -8284 6276 -8268
rect 7240 -8476 7330 -8446
rect 7240 -8510 7268 -8476
rect 7302 -8510 7330 -8476
rect 7240 -8538 7330 -8510
rect 8258 -8476 8348 -8446
rect 8258 -8510 8286 -8476
rect 8320 -8510 8348 -8476
rect 8258 -8538 8348 -8510
rect 9276 -8476 9366 -8446
rect 9276 -8510 9304 -8476
rect 9338 -8510 9366 -8476
rect 9276 -8538 9366 -8510
rect 10294 -8476 10384 -8446
rect 10294 -8510 10322 -8476
rect 10356 -8510 10384 -8476
rect 10294 -8538 10384 -8510
rect 11312 -8476 11402 -8446
rect 11312 -8510 11340 -8476
rect 11374 -8510 11402 -8476
rect 11312 -8538 11402 -8510
rect 12330 -8476 12420 -8446
rect 12330 -8510 12358 -8476
rect 12392 -8510 12420 -8476
rect 12330 -8538 12420 -8510
rect 13348 -8476 13438 -8446
rect 13348 -8510 13376 -8476
rect 13410 -8510 13438 -8476
rect 13348 -8538 13438 -8510
rect 14366 -8476 14456 -8446
rect 14366 -8510 14394 -8476
rect 14428 -8510 14456 -8476
rect 14366 -8538 14456 -8510
rect 15384 -8476 15474 -8446
rect 15384 -8510 15412 -8476
rect 15446 -8510 15474 -8476
rect 15384 -8538 15474 -8510
rect 16402 -8476 16492 -8446
rect 16402 -8510 16430 -8476
rect 16464 -8510 16492 -8476
rect 16402 -8538 16492 -8510
rect 17420 -8476 17510 -8446
rect 17420 -8510 17448 -8476
rect 17482 -8510 17510 -8476
rect 17420 -8538 17510 -8510
rect 18438 -8476 18528 -8446
rect 18438 -8510 18466 -8476
rect 18500 -8510 18528 -8476
rect 18438 -8538 18528 -8510
rect 19456 -8476 19546 -8446
rect 19456 -8510 19484 -8476
rect 19518 -8510 19546 -8476
rect 19456 -8538 19546 -8510
rect 20474 -8476 20564 -8446
rect 20474 -8510 20502 -8476
rect 20536 -8510 20564 -8476
rect 20474 -8538 20564 -8510
rect 21492 -8476 21582 -8446
rect 21492 -8510 21520 -8476
rect 21554 -8510 21582 -8476
rect 21492 -8538 21582 -8510
rect 22510 -8476 22600 -8446
rect 22510 -8510 22538 -8476
rect 22572 -8510 22600 -8476
rect 22510 -8538 22600 -8510
rect 7706 -8793 7722 -8759
rect 8278 -8793 8294 -8759
rect 8724 -8793 8740 -8759
rect 9296 -8793 9312 -8759
rect 9742 -8793 9758 -8759
rect 10314 -8793 10330 -8759
rect 10760 -8793 10776 -8759
rect 11332 -8793 11348 -8759
rect 11778 -8793 11794 -8759
rect 12350 -8793 12366 -8759
rect 12796 -8793 12812 -8759
rect 13368 -8793 13384 -8759
rect 13814 -8793 13830 -8759
rect 14386 -8793 14402 -8759
rect 14832 -8793 14848 -8759
rect 15404 -8793 15420 -8759
rect 15850 -8793 15866 -8759
rect 16422 -8793 16438 -8759
rect 16868 -8793 16884 -8759
rect 17440 -8793 17456 -8759
rect 17886 -8793 17902 -8759
rect 18458 -8793 18474 -8759
rect 18904 -8793 18920 -8759
rect 19476 -8793 19492 -8759
rect 19922 -8793 19938 -8759
rect 20494 -8793 20510 -8759
rect 20940 -8793 20956 -8759
rect 21512 -8793 21528 -8759
rect 21958 -8793 21974 -8759
rect 22530 -8793 22546 -8759
rect 6242 -8876 6276 -8860
rect 7474 -8852 7508 -8836
rect 2402 -8953 2418 -8919
rect 2974 -8953 2990 -8919
rect 3420 -8953 3436 -8919
rect 3992 -8953 4008 -8919
rect 4438 -8953 4454 -8919
rect 5010 -8953 5026 -8919
rect 5456 -8953 5472 -8919
rect 6028 -8953 6044 -8919
rect 2664 -9188 2754 -9158
rect 2664 -9222 2692 -9188
rect 2726 -9222 2754 -9188
rect 2664 -9250 2754 -9222
rect 3682 -9188 3772 -9158
rect 3682 -9222 3710 -9188
rect 3744 -9222 3772 -9188
rect 3682 -9250 3772 -9222
rect 4700 -9188 4790 -9158
rect 4700 -9222 4728 -9188
rect 4762 -9222 4790 -9188
rect 4700 -9250 4790 -9222
rect 5718 -9188 5808 -9158
rect 5718 -9222 5746 -9188
rect 5780 -9222 5808 -9188
rect 5718 -9250 5808 -9222
rect 7474 -9444 7508 -9428
rect 8492 -8852 8526 -8836
rect 8492 -9444 8526 -9428
rect 9510 -8852 9544 -8836
rect 9510 -9444 9544 -9428
rect 10528 -8852 10562 -8836
rect 10528 -9444 10562 -9428
rect 11546 -8852 11580 -8836
rect 11546 -9444 11580 -9428
rect 12564 -8852 12598 -8836
rect 12564 -9444 12598 -9428
rect 13582 -8852 13616 -8836
rect 13582 -9444 13616 -9428
rect 14600 -8852 14634 -8836
rect 14600 -9444 14634 -9428
rect 15618 -8852 15652 -8836
rect 15618 -9444 15652 -9428
rect 16636 -8852 16670 -8836
rect 16636 -9444 16670 -9428
rect 17654 -8852 17688 -8836
rect 17654 -9444 17688 -9428
rect 18672 -8852 18706 -8836
rect 18672 -9444 18706 -9428
rect 19690 -8852 19724 -8836
rect 19690 -9444 19724 -9428
rect 20708 -8852 20742 -8836
rect 20708 -9444 20742 -9428
rect 21726 -8852 21760 -8836
rect 21726 -9444 21760 -9428
rect 22744 -8852 22778 -8836
rect 22744 -9444 22778 -9428
rect 7706 -9521 7722 -9487
rect 8278 -9521 8294 -9487
rect 8724 -9521 8740 -9487
rect 9296 -9521 9312 -9487
rect 9742 -9521 9758 -9487
rect 10314 -9521 10330 -9487
rect 10760 -9521 10776 -9487
rect 11332 -9521 11348 -9487
rect 11778 -9521 11794 -9487
rect 12350 -9521 12366 -9487
rect 12796 -9521 12812 -9487
rect 13368 -9521 13384 -9487
rect 13814 -9521 13830 -9487
rect 14386 -9521 14402 -9487
rect 14832 -9521 14848 -9487
rect 15404 -9521 15420 -9487
rect 15850 -9521 15866 -9487
rect 16422 -9521 16438 -9487
rect 16868 -9521 16884 -9487
rect 17440 -9521 17456 -9487
rect 17886 -9521 17902 -9487
rect 18458 -9521 18474 -9487
rect 18904 -9521 18920 -9487
rect 19476 -9521 19492 -9487
rect 19922 -9521 19938 -9487
rect 20494 -9521 20510 -9487
rect 20940 -9521 20956 -9487
rect 21512 -9521 21528 -9487
rect 21958 -9521 21974 -9487
rect 22530 -9521 22546 -9487
rect 378 -10348 478 -10186
rect 24722 -10348 24822 -10186
rect -12322 -11340 -12222 -11178
rect 24822 -11340 24922 -11178
rect 3086 -11784 3168 -11760
rect 3086 -11818 3110 -11784
rect 3144 -11818 3168 -11784
rect 3086 -11842 3168 -11818
rect 4104 -11784 4186 -11760
rect 4104 -11818 4128 -11784
rect 4162 -11818 4186 -11784
rect 4104 -11842 4186 -11818
rect 5122 -11784 5204 -11760
rect 5122 -11818 5146 -11784
rect 5180 -11818 5204 -11784
rect 5122 -11842 5204 -11818
rect 6140 -11784 6222 -11760
rect 6140 -11818 6164 -11784
rect 6198 -11818 6222 -11784
rect 6140 -11842 6222 -11818
rect 7158 -11784 7240 -11760
rect 7158 -11818 7182 -11784
rect 7216 -11818 7240 -11784
rect 7158 -11842 7240 -11818
rect 8176 -11784 8258 -11760
rect 8176 -11818 8200 -11784
rect 8234 -11818 8258 -11784
rect 8176 -11842 8258 -11818
rect 9194 -11784 9276 -11760
rect 9194 -11818 9218 -11784
rect 9252 -11818 9276 -11784
rect 9194 -11842 9276 -11818
rect 10212 -11784 10294 -11760
rect 10212 -11818 10236 -11784
rect 10270 -11818 10294 -11784
rect 10212 -11842 10294 -11818
rect 11230 -11784 11312 -11760
rect 11230 -11818 11254 -11784
rect 11288 -11818 11312 -11784
rect 11230 -11842 11312 -11818
rect 12248 -11784 12330 -11760
rect 12248 -11818 12272 -11784
rect 12306 -11818 12330 -11784
rect 12248 -11842 12330 -11818
rect 13266 -11784 13348 -11760
rect 13266 -11818 13290 -11784
rect 13324 -11818 13348 -11784
rect 13266 -11842 13348 -11818
rect 14284 -11784 14366 -11760
rect 14284 -11818 14308 -11784
rect 14342 -11818 14366 -11784
rect 14284 -11842 14366 -11818
rect 15302 -11784 15384 -11760
rect 15302 -11818 15326 -11784
rect 15360 -11818 15384 -11784
rect 15302 -11842 15384 -11818
rect 16320 -11784 16402 -11760
rect 16320 -11818 16344 -11784
rect 16378 -11818 16402 -11784
rect 16320 -11842 16402 -11818
rect 17338 -11784 17420 -11760
rect 17338 -11818 17362 -11784
rect 17396 -11818 17420 -11784
rect 17338 -11842 17420 -11818
rect 18356 -11784 18438 -11760
rect 18356 -11818 18380 -11784
rect 18414 -11818 18438 -11784
rect 18356 -11842 18438 -11818
rect 19374 -11784 19456 -11760
rect 19374 -11818 19398 -11784
rect 19432 -11818 19456 -11784
rect 19374 -11842 19456 -11818
rect 20392 -11784 20474 -11760
rect 20392 -11818 20416 -11784
rect 20450 -11818 20474 -11784
rect 20392 -11842 20474 -11818
rect 21410 -11784 21492 -11760
rect 21410 -11818 21434 -11784
rect 21468 -11818 21492 -11784
rect 21410 -11842 21492 -11818
rect 22428 -11784 22510 -11760
rect 22428 -11818 22452 -11784
rect 22486 -11818 22510 -11784
rect 22428 -11842 22510 -11818
rect 2814 -11998 2830 -11964
rect 3386 -11998 3402 -11964
rect 3832 -11998 3848 -11964
rect 4404 -11998 4420 -11964
rect 4850 -11998 4866 -11964
rect 5422 -11998 5438 -11964
rect 5868 -11998 5884 -11964
rect 6440 -11998 6456 -11964
rect 6886 -11998 6902 -11964
rect 7458 -11998 7474 -11964
rect 7904 -11998 7920 -11964
rect 8476 -11998 8492 -11964
rect 8922 -11998 8938 -11964
rect 9494 -11998 9510 -11964
rect 9940 -11998 9956 -11964
rect 10512 -11998 10528 -11964
rect 10958 -11998 10974 -11964
rect 11530 -11998 11546 -11964
rect 11976 -11998 11992 -11964
rect 12548 -11998 12564 -11964
rect 12994 -11998 13010 -11964
rect 13566 -11998 13582 -11964
rect 14012 -11998 14028 -11964
rect 14584 -11998 14600 -11964
rect 15030 -11998 15046 -11964
rect 15602 -11998 15618 -11964
rect 16048 -11998 16064 -11964
rect 16620 -11998 16636 -11964
rect 17066 -11998 17082 -11964
rect 17638 -11998 17654 -11964
rect 18084 -11998 18100 -11964
rect 18656 -11998 18672 -11964
rect 19102 -11998 19118 -11964
rect 19674 -11998 19690 -11964
rect 20120 -11998 20136 -11964
rect 20692 -11998 20708 -11964
rect 21138 -11998 21154 -11964
rect 21710 -11998 21726 -11964
rect 22156 -11998 22172 -11964
rect 22728 -11998 22744 -11964
rect 2582 -12048 2616 -12032
rect -9208 -12386 -9126 -12362
rect -9208 -12420 -9184 -12386
rect -9150 -12420 -9126 -12386
rect -9208 -12444 -9126 -12420
rect -8190 -12386 -8108 -12362
rect -8190 -12420 -8166 -12386
rect -8132 -12420 -8108 -12386
rect -8952 -12474 -8936 -12440
rect -8380 -12474 -8364 -12440
rect -8190 -12444 -8108 -12420
rect -7172 -12386 -7090 -12362
rect -7172 -12420 -7148 -12386
rect -7114 -12420 -7090 -12386
rect -7934 -12474 -7918 -12440
rect -7362 -12474 -7346 -12440
rect -7172 -12444 -7090 -12420
rect -6154 -12386 -6072 -12362
rect -6154 -12420 -6130 -12386
rect -6096 -12420 -6072 -12386
rect -6916 -12474 -6900 -12440
rect -6344 -12474 -6328 -12440
rect -6154 -12444 -6072 -12420
rect -5136 -12386 -5054 -12362
rect -5136 -12420 -5112 -12386
rect -5078 -12420 -5054 -12386
rect -5898 -12474 -5882 -12440
rect -5326 -12474 -5310 -12440
rect -5136 -12444 -5054 -12420
rect -4118 -12386 -4036 -12362
rect -4118 -12420 -4094 -12386
rect -4060 -12420 -4036 -12386
rect -4880 -12474 -4864 -12440
rect -4308 -12474 -4292 -12440
rect -4118 -12444 -4036 -12420
rect -3100 -12386 -3018 -12362
rect -3100 -12420 -3076 -12386
rect -3042 -12420 -3018 -12386
rect -3862 -12474 -3846 -12440
rect -3290 -12474 -3274 -12440
rect -3100 -12444 -3018 -12420
rect -2082 -12386 -2000 -12362
rect -2082 -12420 -2058 -12386
rect -2024 -12420 -2000 -12386
rect -2844 -12474 -2828 -12440
rect -2272 -12474 -2256 -12440
rect -2082 -12444 -2000 -12420
rect -1064 -12386 -982 -12362
rect -1064 -12420 -1040 -12386
rect -1006 -12420 -982 -12386
rect -1826 -12474 -1810 -12440
rect -1254 -12474 -1238 -12440
rect -1064 -12444 -982 -12420
rect -36 -12386 46 -12362
rect -36 -12420 -12 -12386
rect 22 -12420 46 -12386
rect -808 -12474 -792 -12440
rect -236 -12474 -220 -12440
rect -36 -12444 46 -12420
rect -9184 -12524 -9150 -12508
rect -9184 -13116 -9150 -13100
rect -8166 -12524 -8132 -12508
rect -8166 -13116 -8132 -13100
rect -7148 -12524 -7114 -12508
rect -7148 -13116 -7114 -13100
rect -6130 -12524 -6096 -12508
rect -6130 -13116 -6096 -13100
rect -5112 -12524 -5078 -12508
rect -5112 -13116 -5078 -13100
rect -4094 -12524 -4060 -12508
rect -4094 -13116 -4060 -13100
rect -3076 -12524 -3042 -12508
rect -3076 -13116 -3042 -13100
rect -2058 -12524 -2024 -12508
rect -2058 -13116 -2024 -13100
rect -1040 -12524 -1006 -12508
rect -1040 -13116 -1006 -13100
rect -22 -12524 12 -12508
rect 2582 -12640 2616 -12624
rect 3600 -12048 3634 -12032
rect 3600 -12640 3634 -12624
rect 4618 -12048 4652 -12032
rect 4618 -12640 4652 -12624
rect 5636 -12048 5670 -12032
rect 5636 -12640 5670 -12624
rect 6654 -12048 6688 -12032
rect 6654 -12640 6688 -12624
rect 7672 -12048 7706 -12032
rect 7672 -12640 7706 -12624
rect 8690 -12048 8724 -12032
rect 8690 -12640 8724 -12624
rect 9708 -12048 9742 -12032
rect 9708 -12640 9742 -12624
rect 10726 -12048 10760 -12032
rect 10726 -12640 10760 -12624
rect 11744 -12048 11778 -12032
rect 11744 -12640 11778 -12624
rect 12762 -12048 12796 -12032
rect 12762 -12640 12796 -12624
rect 13780 -12048 13814 -12032
rect 13780 -12640 13814 -12624
rect 14798 -12048 14832 -12032
rect 14798 -12640 14832 -12624
rect 15816 -12048 15850 -12032
rect 15816 -12640 15850 -12624
rect 16834 -12048 16868 -12032
rect 16834 -12640 16868 -12624
rect 17852 -12048 17886 -12032
rect 17852 -12640 17886 -12624
rect 18870 -12048 18904 -12032
rect 18870 -12640 18904 -12624
rect 19888 -12048 19922 -12032
rect 19888 -12640 19922 -12624
rect 20906 -12048 20940 -12032
rect 20906 -12640 20940 -12624
rect 21924 -12048 21958 -12032
rect 21924 -12640 21958 -12624
rect 22942 -12048 22976 -12032
rect 22942 -12640 22976 -12624
rect 2814 -12708 2830 -12674
rect 3386 -12708 3402 -12674
rect 3832 -12708 3848 -12674
rect 4404 -12708 4420 -12674
rect 4850 -12708 4866 -12674
rect 5422 -12708 5438 -12674
rect 5868 -12708 5884 -12674
rect 6440 -12708 6456 -12674
rect 6886 -12708 6902 -12674
rect 7458 -12708 7474 -12674
rect 7904 -12708 7920 -12674
rect 8476 -12708 8492 -12674
rect 8922 -12708 8938 -12674
rect 9494 -12708 9510 -12674
rect 9940 -12708 9956 -12674
rect 10512 -12708 10528 -12674
rect 10958 -12708 10974 -12674
rect 11530 -12708 11546 -12674
rect 11976 -12708 11992 -12674
rect 12548 -12708 12564 -12674
rect 12994 -12708 13010 -12674
rect 13566 -12708 13582 -12674
rect 14012 -12708 14028 -12674
rect 14584 -12708 14600 -12674
rect 15030 -12708 15046 -12674
rect 15602 -12708 15618 -12674
rect 16048 -12708 16064 -12674
rect 16620 -12708 16636 -12674
rect 17066 -12708 17082 -12674
rect 17638 -12708 17654 -12674
rect 18084 -12708 18100 -12674
rect 18656 -12708 18672 -12674
rect 19102 -12708 19118 -12674
rect 19674 -12708 19690 -12674
rect 20120 -12708 20136 -12674
rect 20692 -12708 20708 -12674
rect 21138 -12708 21154 -12674
rect 21710 -12708 21726 -12674
rect 22156 -12708 22172 -12674
rect 22728 -12708 22744 -12674
rect 2814 -12816 2830 -12782
rect 3386 -12816 3402 -12782
rect 3832 -12816 3848 -12782
rect 4404 -12816 4420 -12782
rect 4850 -12816 4866 -12782
rect 5422 -12816 5438 -12782
rect 5868 -12816 5884 -12782
rect 6440 -12816 6456 -12782
rect 6886 -12816 6902 -12782
rect 7458 -12816 7474 -12782
rect 7904 -12816 7920 -12782
rect 8476 -12816 8492 -12782
rect 8922 -12816 8938 -12782
rect 9494 -12816 9510 -12782
rect 9940 -12816 9956 -12782
rect 10512 -12816 10528 -12782
rect 10958 -12816 10974 -12782
rect 11530 -12816 11546 -12782
rect 11976 -12816 11992 -12782
rect 12548 -12816 12564 -12782
rect 12994 -12816 13010 -12782
rect 13566 -12816 13582 -12782
rect 14012 -12816 14028 -12782
rect 14584 -12816 14600 -12782
rect 15030 -12816 15046 -12782
rect 15602 -12816 15618 -12782
rect 16048 -12816 16064 -12782
rect 16620 -12816 16636 -12782
rect 17066 -12816 17082 -12782
rect 17638 -12816 17654 -12782
rect 18084 -12816 18100 -12782
rect 18656 -12816 18672 -12782
rect 19102 -12816 19118 -12782
rect 19674 -12816 19690 -12782
rect 20120 -12816 20136 -12782
rect 20692 -12816 20708 -12782
rect 21138 -12816 21154 -12782
rect 21710 -12816 21726 -12782
rect 22156 -12816 22172 -12782
rect 22728 -12816 22744 -12782
rect -22 -13116 12 -13100
rect 2582 -12866 2616 -12850
rect -9208 -13204 -9126 -13180
rect -8952 -13184 -8936 -13150
rect -8380 -13184 -8364 -13150
rect -9208 -13238 -9184 -13204
rect -9150 -13238 -9126 -13204
rect -9208 -13262 -9126 -13238
rect -8190 -13204 -8108 -13180
rect -7934 -13184 -7918 -13150
rect -7362 -13184 -7346 -13150
rect -8190 -13238 -8166 -13204
rect -8132 -13238 -8108 -13204
rect -8952 -13292 -8936 -13258
rect -8380 -13292 -8364 -13258
rect -8190 -13262 -8108 -13238
rect -7172 -13204 -7090 -13180
rect -6916 -13184 -6900 -13150
rect -6344 -13184 -6328 -13150
rect -7172 -13238 -7148 -13204
rect -7114 -13238 -7090 -13204
rect -7934 -13292 -7918 -13258
rect -7362 -13292 -7346 -13258
rect -7172 -13262 -7090 -13238
rect -6154 -13204 -6072 -13180
rect -5898 -13184 -5882 -13150
rect -5326 -13184 -5310 -13150
rect -6154 -13238 -6130 -13204
rect -6096 -13238 -6072 -13204
rect -6916 -13292 -6900 -13258
rect -6344 -13292 -6328 -13258
rect -6154 -13262 -6072 -13238
rect -5136 -13204 -5054 -13180
rect -4880 -13184 -4864 -13150
rect -4308 -13184 -4292 -13150
rect -5136 -13238 -5112 -13204
rect -5078 -13238 -5054 -13204
rect -5898 -13292 -5882 -13258
rect -5326 -13292 -5310 -13258
rect -5136 -13262 -5054 -13238
rect -4118 -13204 -4036 -13180
rect -3862 -13184 -3846 -13150
rect -3290 -13184 -3274 -13150
rect -4118 -13238 -4094 -13204
rect -4060 -13238 -4036 -13204
rect -4880 -13292 -4864 -13258
rect -4308 -13292 -4292 -13258
rect -4118 -13262 -4036 -13238
rect -3100 -13204 -3018 -13180
rect -2844 -13184 -2828 -13150
rect -2272 -13184 -2256 -13150
rect -3100 -13238 -3076 -13204
rect -3042 -13238 -3018 -13204
rect -3862 -13292 -3846 -13258
rect -3290 -13292 -3274 -13258
rect -3100 -13262 -3018 -13238
rect -2082 -13204 -2000 -13180
rect -1826 -13184 -1810 -13150
rect -1254 -13184 -1238 -13150
rect -2082 -13238 -2058 -13204
rect -2024 -13238 -2000 -13204
rect -2844 -13292 -2828 -13258
rect -2272 -13292 -2256 -13258
rect -2082 -13262 -2000 -13238
rect -1064 -13204 -982 -13180
rect -808 -13184 -792 -13150
rect -236 -13184 -220 -13150
rect -1064 -13238 -1040 -13204
rect -1006 -13238 -982 -13204
rect -1826 -13292 -1810 -13258
rect -1254 -13292 -1238 -13258
rect -1064 -13262 -982 -13238
rect -36 -13204 46 -13180
rect -36 -13238 -12 -13204
rect 22 -13238 46 -13204
rect -808 -13292 -792 -13258
rect -236 -13292 -220 -13258
rect -36 -13262 46 -13238
rect -3592 -13294 -3532 -13292
rect -9184 -13342 -9150 -13326
rect -9184 -13934 -9150 -13918
rect -8166 -13342 -8132 -13326
rect -8166 -13934 -8132 -13918
rect -7148 -13342 -7114 -13326
rect -7148 -13934 -7114 -13918
rect -6130 -13342 -6096 -13326
rect -6130 -13934 -6096 -13918
rect -5112 -13342 -5078 -13326
rect -5112 -13934 -5078 -13918
rect -4094 -13342 -4060 -13326
rect -4094 -13934 -4060 -13918
rect -3076 -13342 -3042 -13326
rect -3076 -13934 -3042 -13918
rect -2058 -13342 -2024 -13326
rect -2058 -13934 -2024 -13918
rect -1040 -13342 -1006 -13326
rect -1040 -13934 -1006 -13918
rect -22 -13342 12 -13326
rect 2582 -13458 2616 -13442
rect 3600 -12866 3634 -12850
rect 3600 -13458 3634 -13442
rect 4618 -12866 4652 -12850
rect 4618 -13458 4652 -13442
rect 5636 -12866 5670 -12850
rect 5636 -13458 5670 -13442
rect 6654 -12866 6688 -12850
rect 6654 -13458 6688 -13442
rect 7672 -12866 7706 -12850
rect 7672 -13458 7706 -13442
rect 8690 -12866 8724 -12850
rect 8690 -13458 8724 -13442
rect 9708 -12866 9742 -12850
rect 9708 -13458 9742 -13442
rect 10726 -12866 10760 -12850
rect 10726 -13458 10760 -13442
rect 11744 -12866 11778 -12850
rect 11744 -13458 11778 -13442
rect 12762 -12866 12796 -12850
rect 12762 -13458 12796 -13442
rect 13780 -12866 13814 -12850
rect 13780 -13458 13814 -13442
rect 14798 -12866 14832 -12850
rect 14798 -13458 14832 -13442
rect 15816 -12866 15850 -12850
rect 15816 -13458 15850 -13442
rect 16834 -12866 16868 -12850
rect 16834 -13458 16868 -13442
rect 17852 -12866 17886 -12850
rect 17852 -13458 17886 -13442
rect 18870 -12866 18904 -12850
rect 18870 -13458 18904 -13442
rect 19888 -12866 19922 -12850
rect 19888 -13458 19922 -13442
rect 20906 -12866 20940 -12850
rect 20906 -13458 20940 -13442
rect 21924 -12866 21958 -12850
rect 21924 -13458 21958 -13442
rect 22942 -12866 22976 -12850
rect 22942 -13458 22976 -13442
rect 2814 -13526 2830 -13492
rect 3386 -13526 3402 -13492
rect 3832 -13526 3848 -13492
rect 4404 -13526 4420 -13492
rect 4850 -13526 4866 -13492
rect 5422 -13526 5438 -13492
rect 5868 -13526 5884 -13492
rect 6440 -13526 6456 -13492
rect 6886 -13526 6902 -13492
rect 7458 -13526 7474 -13492
rect 7904 -13526 7920 -13492
rect 8476 -13526 8492 -13492
rect 8922 -13526 8938 -13492
rect 9494 -13526 9510 -13492
rect 9940 -13526 9956 -13492
rect 10512 -13526 10528 -13492
rect 10958 -13526 10974 -13492
rect 11530 -13526 11546 -13492
rect 11976 -13526 11992 -13492
rect 12548 -13526 12564 -13492
rect 12994 -13526 13010 -13492
rect 13566 -13526 13582 -13492
rect 14012 -13526 14028 -13492
rect 14584 -13526 14600 -13492
rect 15030 -13526 15046 -13492
rect 15602 -13526 15618 -13492
rect 16048 -13526 16064 -13492
rect 16620 -13526 16636 -13492
rect 17066 -13526 17082 -13492
rect 17638 -13526 17654 -13492
rect 18084 -13526 18100 -13492
rect 18656 -13526 18672 -13492
rect 19102 -13526 19118 -13492
rect 19674 -13526 19690 -13492
rect 20120 -13526 20136 -13492
rect 20692 -13526 20708 -13492
rect 21138 -13526 21154 -13492
rect 21710 -13526 21726 -13492
rect 22156 -13526 22172 -13492
rect 22728 -13526 22744 -13492
rect 3098 -13810 3180 -13786
rect 3098 -13844 3122 -13810
rect 3156 -13844 3180 -13810
rect 3098 -13868 3180 -13844
rect 4116 -13810 4198 -13786
rect 4116 -13844 4140 -13810
rect 4174 -13844 4198 -13810
rect 4116 -13868 4198 -13844
rect 5134 -13810 5216 -13786
rect 5134 -13844 5158 -13810
rect 5192 -13844 5216 -13810
rect 5134 -13868 5216 -13844
rect 6152 -13810 6234 -13786
rect 6152 -13844 6176 -13810
rect 6210 -13844 6234 -13810
rect 6152 -13868 6234 -13844
rect 7170 -13810 7252 -13786
rect 7170 -13844 7194 -13810
rect 7228 -13844 7252 -13810
rect 7170 -13868 7252 -13844
rect 8188 -13810 8270 -13786
rect 8188 -13844 8212 -13810
rect 8246 -13844 8270 -13810
rect 8188 -13868 8270 -13844
rect 9206 -13810 9288 -13786
rect 9206 -13844 9230 -13810
rect 9264 -13844 9288 -13810
rect 9206 -13868 9288 -13844
rect 10224 -13810 10306 -13786
rect 10224 -13844 10248 -13810
rect 10282 -13844 10306 -13810
rect 10224 -13868 10306 -13844
rect 11242 -13810 11324 -13786
rect 11242 -13844 11266 -13810
rect 11300 -13844 11324 -13810
rect 11242 -13868 11324 -13844
rect 12260 -13810 12342 -13786
rect 12260 -13844 12284 -13810
rect 12318 -13844 12342 -13810
rect 12260 -13868 12342 -13844
rect 13278 -13810 13360 -13786
rect 13278 -13844 13302 -13810
rect 13336 -13844 13360 -13810
rect 13278 -13868 13360 -13844
rect 14296 -13810 14378 -13786
rect 14296 -13844 14320 -13810
rect 14354 -13844 14378 -13810
rect 14296 -13868 14378 -13844
rect 15314 -13810 15396 -13786
rect 15314 -13844 15338 -13810
rect 15372 -13844 15396 -13810
rect 15314 -13868 15396 -13844
rect 16332 -13810 16414 -13786
rect 16332 -13844 16356 -13810
rect 16390 -13844 16414 -13810
rect 16332 -13868 16414 -13844
rect 17350 -13810 17432 -13786
rect 17350 -13844 17374 -13810
rect 17408 -13844 17432 -13810
rect 17350 -13868 17432 -13844
rect 18368 -13810 18450 -13786
rect 18368 -13844 18392 -13810
rect 18426 -13844 18450 -13810
rect 18368 -13868 18450 -13844
rect 19386 -13810 19468 -13786
rect 19386 -13844 19410 -13810
rect 19444 -13844 19468 -13810
rect 19386 -13868 19468 -13844
rect 20404 -13810 20486 -13786
rect 20404 -13844 20428 -13810
rect 20462 -13844 20486 -13810
rect 20404 -13868 20486 -13844
rect 21422 -13810 21504 -13786
rect 21422 -13844 21446 -13810
rect 21480 -13844 21504 -13810
rect 21422 -13868 21504 -13844
rect 22440 -13810 22522 -13786
rect 22440 -13844 22464 -13810
rect 22498 -13844 22522 -13810
rect 22440 -13868 22522 -13844
rect -22 -13934 12 -13918
rect -7660 -13968 -7600 -13966
rect -6646 -13968 -6586 -13966
rect -2572 -13968 -2512 -13966
rect -1556 -13968 -1496 -13966
rect -9208 -14022 -9126 -13998
rect -8952 -14002 -8936 -13968
rect -8380 -14002 -8364 -13968
rect -9208 -14056 -9184 -14022
rect -9150 -14056 -9126 -14022
rect -9208 -14080 -9126 -14056
rect -8190 -14022 -8108 -13998
rect -7934 -14002 -7918 -13968
rect -7362 -14002 -7346 -13968
rect -8190 -14056 -8166 -14022
rect -8132 -14056 -8108 -14022
rect -8952 -14110 -8936 -14076
rect -8380 -14110 -8364 -14076
rect -8190 -14080 -8108 -14056
rect -7172 -14022 -7090 -13998
rect -6916 -14002 -6900 -13968
rect -6344 -14002 -6328 -13968
rect -7172 -14056 -7148 -14022
rect -7114 -14056 -7090 -14022
rect -7934 -14110 -7918 -14076
rect -7362 -14110 -7346 -14076
rect -7172 -14080 -7090 -14056
rect -6154 -14022 -6072 -13998
rect -5898 -14002 -5882 -13968
rect -5326 -14002 -5310 -13968
rect -6154 -14056 -6130 -14022
rect -6096 -14056 -6072 -14022
rect -6916 -14110 -6900 -14076
rect -6344 -14110 -6328 -14076
rect -6154 -14080 -6072 -14056
rect -5136 -14022 -5054 -13998
rect -4880 -14002 -4864 -13968
rect -4308 -14002 -4292 -13968
rect -5136 -14056 -5112 -14022
rect -5078 -14056 -5054 -14022
rect -5898 -14110 -5882 -14076
rect -5326 -14110 -5310 -14076
rect -5136 -14080 -5054 -14056
rect -4118 -14022 -4036 -13998
rect -3862 -14002 -3846 -13968
rect -3290 -14002 -3274 -13968
rect -4118 -14056 -4094 -14022
rect -4060 -14056 -4036 -14022
rect -4880 -14110 -4864 -14076
rect -4308 -14110 -4292 -14076
rect -4118 -14080 -4036 -14056
rect -3100 -14022 -3018 -13998
rect -2844 -14002 -2828 -13968
rect -2272 -14002 -2256 -13968
rect -3100 -14056 -3076 -14022
rect -3042 -14056 -3018 -14022
rect -3862 -14110 -3846 -14076
rect -3290 -14110 -3274 -14076
rect -3100 -14080 -3018 -14056
rect -2082 -14022 -2000 -13998
rect -1826 -14002 -1810 -13968
rect -1254 -14002 -1238 -13968
rect -2082 -14056 -2058 -14022
rect -2024 -14056 -2000 -14022
rect -2844 -14110 -2828 -14076
rect -2272 -14110 -2256 -14076
rect -2082 -14080 -2000 -14056
rect -1064 -14022 -982 -13998
rect -808 -14002 -792 -13968
rect -236 -14002 -220 -13968
rect -1064 -14056 -1040 -14022
rect -1006 -14056 -982 -14022
rect -1826 -14110 -1810 -14076
rect -1254 -14110 -1238 -14076
rect -1064 -14080 -982 -14056
rect -36 -14022 46 -13998
rect -36 -14056 -12 -14022
rect 22 -14056 46 -14022
rect -808 -14110 -792 -14076
rect -236 -14110 -220 -14076
rect -36 -14080 46 -14056
rect -9184 -14160 -9150 -14144
rect -9184 -14752 -9150 -14736
rect -8166 -14160 -8132 -14144
rect -8166 -14752 -8132 -14736
rect -7148 -14160 -7114 -14144
rect -7148 -14752 -7114 -14736
rect -6130 -14160 -6096 -14144
rect -6130 -14752 -6096 -14736
rect -5112 -14160 -5078 -14144
rect -5112 -14752 -5078 -14736
rect -4094 -14160 -4060 -14144
rect -4094 -14752 -4060 -14736
rect -3076 -14160 -3042 -14144
rect -3076 -14752 -3042 -14736
rect -2058 -14160 -2024 -14144
rect -2058 -14752 -2024 -14736
rect -1040 -14160 -1006 -14144
rect -1040 -14752 -1006 -14736
rect -22 -14160 12 -14144
rect 2814 -14194 2830 -14160
rect 3386 -14194 3402 -14160
rect 3832 -14194 3848 -14160
rect 4404 -14194 4420 -14160
rect 4850 -14194 4866 -14160
rect 5422 -14194 5438 -14160
rect 5868 -14194 5884 -14160
rect 6440 -14194 6456 -14160
rect 6886 -14194 6902 -14160
rect 7458 -14194 7474 -14160
rect 7904 -14194 7920 -14160
rect 8476 -14194 8492 -14160
rect 8922 -14194 8938 -14160
rect 9494 -14194 9510 -14160
rect 9940 -14194 9956 -14160
rect 10512 -14194 10528 -14160
rect 10958 -14194 10974 -14160
rect 11530 -14194 11546 -14160
rect 11976 -14194 11992 -14160
rect 12548 -14194 12564 -14160
rect 12994 -14194 13010 -14160
rect 13566 -14194 13582 -14160
rect 14012 -14194 14028 -14160
rect 14584 -14194 14600 -14160
rect 15030 -14194 15046 -14160
rect 15602 -14194 15618 -14160
rect 16048 -14194 16064 -14160
rect 16620 -14194 16636 -14160
rect 17066 -14194 17082 -14160
rect 17638 -14194 17654 -14160
rect 18084 -14194 18100 -14160
rect 18656 -14194 18672 -14160
rect 19102 -14194 19118 -14160
rect 19674 -14194 19690 -14160
rect 20120 -14194 20136 -14160
rect 20692 -14194 20708 -14160
rect 21138 -14194 21154 -14160
rect 21710 -14194 21726 -14160
rect 22156 -14194 22172 -14160
rect 22728 -14194 22744 -14160
rect 12238 -14200 12298 -14194
rect -22 -14752 12 -14736
rect 2582 -14244 2616 -14228
rect -7656 -14786 -7596 -14784
rect -6642 -14786 -6582 -14784
rect -2568 -14786 -2508 -14784
rect -1552 -14786 -1492 -14784
rect -9208 -14840 -9126 -14816
rect -8952 -14820 -8936 -14786
rect -8380 -14820 -8364 -14786
rect -9208 -14874 -9184 -14840
rect -9150 -14874 -9126 -14840
rect -9208 -14898 -9126 -14874
rect -8190 -14840 -8108 -14816
rect -7934 -14820 -7918 -14786
rect -7362 -14820 -7346 -14786
rect -8190 -14874 -8166 -14840
rect -8132 -14874 -8108 -14840
rect -8952 -14928 -8936 -14894
rect -8380 -14928 -8364 -14894
rect -8190 -14898 -8108 -14874
rect -7172 -14840 -7090 -14816
rect -6916 -14820 -6900 -14786
rect -6344 -14820 -6328 -14786
rect -7172 -14874 -7148 -14840
rect -7114 -14874 -7090 -14840
rect -7934 -14928 -7918 -14894
rect -7362 -14928 -7346 -14894
rect -7172 -14898 -7090 -14874
rect -6154 -14840 -6072 -14816
rect -5898 -14820 -5882 -14786
rect -5326 -14820 -5310 -14786
rect -6154 -14874 -6130 -14840
rect -6096 -14874 -6072 -14840
rect -6916 -14928 -6900 -14894
rect -6344 -14928 -6328 -14894
rect -6154 -14898 -6072 -14874
rect -5136 -14840 -5054 -14816
rect -4880 -14820 -4864 -14786
rect -4308 -14820 -4292 -14786
rect -5136 -14874 -5112 -14840
rect -5078 -14874 -5054 -14840
rect -5898 -14928 -5882 -14894
rect -5326 -14928 -5310 -14894
rect -5136 -14898 -5054 -14874
rect -4118 -14840 -4036 -14816
rect -3862 -14820 -3846 -14786
rect -3290 -14820 -3274 -14786
rect -4118 -14874 -4094 -14840
rect -4060 -14874 -4036 -14840
rect -4880 -14928 -4864 -14894
rect -4308 -14928 -4292 -14894
rect -4118 -14898 -4036 -14874
rect -3100 -14840 -3018 -14816
rect -2844 -14820 -2828 -14786
rect -2272 -14820 -2256 -14786
rect -3100 -14874 -3076 -14840
rect -3042 -14874 -3018 -14840
rect -3862 -14928 -3846 -14894
rect -3290 -14928 -3274 -14894
rect -3100 -14898 -3018 -14874
rect -2082 -14840 -2000 -14816
rect -1826 -14820 -1810 -14786
rect -1254 -14820 -1238 -14786
rect -2082 -14874 -2058 -14840
rect -2024 -14874 -2000 -14840
rect -2844 -14928 -2828 -14894
rect -2272 -14928 -2256 -14894
rect -2082 -14898 -2000 -14874
rect -1064 -14840 -982 -14816
rect -808 -14820 -792 -14786
rect -236 -14820 -220 -14786
rect -1064 -14874 -1040 -14840
rect -1006 -14874 -982 -14840
rect -1826 -14928 -1810 -14894
rect -1254 -14928 -1238 -14894
rect -1064 -14898 -982 -14874
rect -36 -14840 46 -14816
rect 2582 -14836 2616 -14820
rect 3600 -14244 3634 -14228
rect 3600 -14836 3634 -14820
rect 4618 -14244 4652 -14228
rect 4618 -14836 4652 -14820
rect 5636 -14244 5670 -14228
rect 5636 -14836 5670 -14820
rect 6654 -14244 6688 -14228
rect 6654 -14836 6688 -14820
rect 7672 -14244 7706 -14228
rect 7672 -14836 7706 -14820
rect 8690 -14244 8724 -14228
rect 8690 -14836 8724 -14820
rect 9708 -14244 9742 -14228
rect 9708 -14836 9742 -14820
rect 10726 -14244 10760 -14228
rect 10726 -14836 10760 -14820
rect 11744 -14244 11778 -14228
rect 11744 -14836 11778 -14820
rect 12762 -14244 12796 -14228
rect 12762 -14836 12796 -14820
rect 13780 -14244 13814 -14228
rect 13780 -14836 13814 -14820
rect 14798 -14244 14832 -14228
rect 14798 -14836 14832 -14820
rect 15816 -14244 15850 -14228
rect 15816 -14836 15850 -14820
rect 16834 -14244 16868 -14228
rect 16834 -14836 16868 -14820
rect 17852 -14244 17886 -14228
rect 17852 -14836 17886 -14820
rect 18870 -14244 18904 -14228
rect 18870 -14836 18904 -14820
rect 19888 -14244 19922 -14228
rect 19888 -14836 19922 -14820
rect 20906 -14244 20940 -14228
rect 20906 -14836 20940 -14820
rect 21924 -14244 21958 -14228
rect 21924 -14836 21958 -14820
rect 22942 -14244 22976 -14228
rect 22942 -14836 22976 -14820
rect -36 -14874 -12 -14840
rect 22 -14874 46 -14840
rect 8166 -14870 8226 -14864
rect 10202 -14870 10262 -14864
rect 11222 -14870 11282 -14864
rect 16294 -14870 16354 -14864
rect -808 -14928 -792 -14894
rect -236 -14928 -220 -14894
rect -36 -14898 46 -14874
rect 2814 -14904 2830 -14870
rect 3386 -14904 3402 -14870
rect 3832 -14904 3848 -14870
rect 4404 -14904 4420 -14870
rect 4850 -14904 4866 -14870
rect 5422 -14904 5438 -14870
rect 5868 -14904 5884 -14870
rect 6440 -14904 6456 -14870
rect 6886 -14904 6902 -14870
rect 7458 -14904 7474 -14870
rect 7904 -14904 7920 -14870
rect 8476 -14904 8492 -14870
rect 8922 -14904 8938 -14870
rect 9494 -14904 9510 -14870
rect 9940 -14904 9956 -14870
rect 10512 -14904 10528 -14870
rect 10958 -14904 10974 -14870
rect 11530 -14904 11546 -14870
rect 11976 -14904 11992 -14870
rect 12548 -14904 12564 -14870
rect 12994 -14904 13010 -14870
rect 13566 -14904 13582 -14870
rect 14012 -14904 14028 -14870
rect 14584 -14904 14600 -14870
rect 15030 -14904 15046 -14870
rect 15602 -14904 15618 -14870
rect 16048 -14904 16064 -14870
rect 16620 -14904 16636 -14870
rect 17066 -14904 17082 -14870
rect 17638 -14904 17654 -14870
rect 18084 -14904 18100 -14870
rect 18656 -14904 18672 -14870
rect 19102 -14904 19118 -14870
rect 19674 -14904 19690 -14870
rect 20120 -14904 20136 -14870
rect 20692 -14904 20708 -14870
rect 21138 -14904 21154 -14870
rect 21710 -14904 21726 -14870
rect 22156 -14904 22172 -14870
rect 22728 -14904 22744 -14870
rect -9184 -14978 -9150 -14962
rect -9184 -15570 -9150 -15554
rect -8166 -14978 -8132 -14962
rect -8166 -15570 -8132 -15554
rect -7148 -14978 -7114 -14962
rect -7148 -15570 -7114 -15554
rect -6130 -14978 -6096 -14962
rect -6130 -15570 -6096 -15554
rect -5112 -14978 -5078 -14962
rect -5112 -15570 -5078 -15554
rect -4094 -14978 -4060 -14962
rect -4094 -15570 -4060 -15554
rect -3076 -14978 -3042 -14962
rect -3076 -15570 -3042 -15554
rect -2058 -14978 -2024 -14962
rect -2058 -15570 -2024 -15554
rect -1040 -14978 -1006 -14962
rect -1040 -15570 -1006 -15554
rect -22 -14978 12 -14962
rect 3086 -15116 3168 -15092
rect 3086 -15150 3110 -15116
rect 3144 -15150 3168 -15116
rect 3086 -15174 3168 -15150
rect 4104 -15116 4186 -15092
rect 4104 -15150 4128 -15116
rect 4162 -15150 4186 -15116
rect 4104 -15174 4186 -15150
rect 5122 -15116 5204 -15092
rect 5122 -15150 5146 -15116
rect 5180 -15150 5204 -15116
rect 5122 -15174 5204 -15150
rect 6140 -15116 6222 -15092
rect 6140 -15150 6164 -15116
rect 6198 -15150 6222 -15116
rect 6140 -15174 6222 -15150
rect 7158 -15116 7240 -15092
rect 7158 -15150 7182 -15116
rect 7216 -15150 7240 -15116
rect 7158 -15174 7240 -15150
rect 8176 -15116 8258 -15092
rect 8176 -15150 8200 -15116
rect 8234 -15150 8258 -15116
rect 8176 -15174 8258 -15150
rect 9194 -15116 9276 -15092
rect 9194 -15150 9218 -15116
rect 9252 -15150 9276 -15116
rect 9194 -15174 9276 -15150
rect 10212 -15116 10294 -15092
rect 10212 -15150 10236 -15116
rect 10270 -15150 10294 -15116
rect 10212 -15174 10294 -15150
rect 11230 -15116 11312 -15092
rect 11230 -15150 11254 -15116
rect 11288 -15150 11312 -15116
rect 11230 -15174 11312 -15150
rect 12248 -15116 12330 -15092
rect 12248 -15150 12272 -15116
rect 12306 -15150 12330 -15116
rect 12248 -15174 12330 -15150
rect 13266 -15116 13348 -15092
rect 13266 -15150 13290 -15116
rect 13324 -15150 13348 -15116
rect 13266 -15174 13348 -15150
rect 14284 -15116 14366 -15092
rect 14284 -15150 14308 -15116
rect 14342 -15150 14366 -15116
rect 14284 -15174 14366 -15150
rect 15302 -15116 15384 -15092
rect 15302 -15150 15326 -15116
rect 15360 -15150 15384 -15116
rect 15302 -15174 15384 -15150
rect 16320 -15116 16402 -15092
rect 16320 -15150 16344 -15116
rect 16378 -15150 16402 -15116
rect 16320 -15174 16402 -15150
rect 17338 -15116 17420 -15092
rect 17338 -15150 17362 -15116
rect 17396 -15150 17420 -15116
rect 17338 -15174 17420 -15150
rect 18356 -15116 18438 -15092
rect 18356 -15150 18380 -15116
rect 18414 -15150 18438 -15116
rect 18356 -15174 18438 -15150
rect 19374 -15116 19456 -15092
rect 19374 -15150 19398 -15116
rect 19432 -15150 19456 -15116
rect 19374 -15174 19456 -15150
rect 20392 -15116 20474 -15092
rect 20392 -15150 20416 -15116
rect 20450 -15150 20474 -15116
rect 20392 -15174 20474 -15150
rect 21410 -15116 21492 -15092
rect 21410 -15150 21434 -15116
rect 21468 -15150 21492 -15116
rect 21410 -15174 21492 -15150
rect 22428 -15116 22510 -15092
rect 22428 -15150 22452 -15116
rect 22486 -15150 22510 -15116
rect 22428 -15174 22510 -15150
rect 2814 -15426 2830 -15392
rect 3386 -15426 3402 -15392
rect 3832 -15426 3848 -15392
rect 4404 -15426 4420 -15392
rect 4850 -15426 4866 -15392
rect 5422 -15426 5438 -15392
rect 5868 -15426 5884 -15392
rect 6440 -15426 6456 -15392
rect 6886 -15426 6902 -15392
rect 7458 -15426 7474 -15392
rect 7904 -15426 7920 -15392
rect 8476 -15426 8492 -15392
rect 8922 -15426 8938 -15392
rect 9494 -15426 9510 -15392
rect 9940 -15426 9956 -15392
rect 10512 -15426 10528 -15392
rect 10958 -15426 10974 -15392
rect 11530 -15426 11546 -15392
rect 11976 -15426 11992 -15392
rect 12548 -15426 12564 -15392
rect 12994 -15426 13010 -15392
rect 13566 -15426 13582 -15392
rect 14012 -15426 14028 -15392
rect 14584 -15426 14600 -15392
rect 15030 -15426 15046 -15392
rect 15602 -15426 15618 -15392
rect 16048 -15426 16064 -15392
rect 16620 -15426 16636 -15392
rect 17066 -15426 17082 -15392
rect 17638 -15426 17654 -15392
rect 18084 -15426 18100 -15392
rect 18656 -15426 18672 -15392
rect 19102 -15426 19118 -15392
rect 19674 -15426 19690 -15392
rect 20120 -15426 20136 -15392
rect 20692 -15426 20708 -15392
rect 21138 -15426 21154 -15392
rect 21710 -15426 21726 -15392
rect 22156 -15426 22172 -15392
rect 22728 -15426 22744 -15392
rect 4100 -15430 4160 -15426
rect 5116 -15430 5176 -15426
rect 9192 -15434 9252 -15426
rect 13258 -15430 13318 -15426
rect 15292 -15430 15352 -15426
rect 21404 -15430 21464 -15426
rect -22 -15570 12 -15554
rect 2582 -15476 2616 -15460
rect -9208 -15658 -9126 -15634
rect -8952 -15638 -8936 -15604
rect -8380 -15638 -8364 -15604
rect -9208 -15692 -9184 -15658
rect -9150 -15692 -9126 -15658
rect -9208 -15716 -9126 -15692
rect -8190 -15658 -8108 -15634
rect -7934 -15638 -7918 -15604
rect -7362 -15638 -7346 -15604
rect -8190 -15692 -8166 -15658
rect -8132 -15692 -8108 -15658
rect -8952 -15746 -8936 -15712
rect -8380 -15746 -8364 -15712
rect -8190 -15716 -8108 -15692
rect -7172 -15658 -7090 -15634
rect -6916 -15638 -6900 -15604
rect -6344 -15638 -6328 -15604
rect -7172 -15692 -7148 -15658
rect -7114 -15692 -7090 -15658
rect -7934 -15746 -7918 -15712
rect -7362 -15746 -7346 -15712
rect -7172 -15716 -7090 -15692
rect -6154 -15658 -6072 -15634
rect -5898 -15638 -5882 -15604
rect -5326 -15638 -5310 -15604
rect -6154 -15692 -6130 -15658
rect -6096 -15692 -6072 -15658
rect -6916 -15746 -6900 -15712
rect -6344 -15746 -6328 -15712
rect -6154 -15716 -6072 -15692
rect -5136 -15658 -5054 -15634
rect -4880 -15638 -4864 -15604
rect -4308 -15638 -4292 -15604
rect -5136 -15692 -5112 -15658
rect -5078 -15692 -5054 -15658
rect -5898 -15746 -5882 -15712
rect -5326 -15746 -5310 -15712
rect -5136 -15716 -5054 -15692
rect -4118 -15658 -4036 -15634
rect -3862 -15638 -3846 -15604
rect -3290 -15638 -3274 -15604
rect -4118 -15692 -4094 -15658
rect -4060 -15692 -4036 -15658
rect -4880 -15746 -4864 -15712
rect -4308 -15746 -4292 -15712
rect -4118 -15716 -4036 -15692
rect -3100 -15658 -3018 -15634
rect -2844 -15638 -2828 -15604
rect -2272 -15638 -2256 -15604
rect -3100 -15692 -3076 -15658
rect -3042 -15692 -3018 -15658
rect -3862 -15746 -3846 -15712
rect -3290 -15746 -3274 -15712
rect -3100 -15716 -3018 -15692
rect -2082 -15658 -2000 -15634
rect -1826 -15638 -1810 -15604
rect -1254 -15638 -1238 -15604
rect -2082 -15692 -2058 -15658
rect -2024 -15692 -2000 -15658
rect -2844 -15746 -2828 -15712
rect -2272 -15746 -2256 -15712
rect -2082 -15716 -2000 -15692
rect -1064 -15658 -982 -15634
rect -808 -15638 -792 -15604
rect -236 -15638 -220 -15604
rect -1064 -15692 -1040 -15658
rect -1006 -15692 -982 -15658
rect -1826 -15746 -1810 -15712
rect -1254 -15746 -1238 -15712
rect -1064 -15716 -982 -15692
rect -36 -15658 46 -15634
rect -36 -15692 -12 -15658
rect 22 -15692 46 -15658
rect -808 -15746 -792 -15712
rect -236 -15746 -220 -15712
rect -36 -15716 46 -15692
rect -3596 -15748 -3536 -15746
rect -9184 -15796 -9150 -15780
rect -9184 -16388 -9150 -16372
rect -8166 -15796 -8132 -15780
rect -8166 -16388 -8132 -16372
rect -7148 -15796 -7114 -15780
rect -7148 -16388 -7114 -16372
rect -6130 -15796 -6096 -15780
rect -6130 -16388 -6096 -16372
rect -5112 -15796 -5078 -15780
rect -5112 -16388 -5078 -16372
rect -4094 -15796 -4060 -15780
rect -4094 -16388 -4060 -16372
rect -3076 -15796 -3042 -15780
rect -3076 -16388 -3042 -16372
rect -2058 -15796 -2024 -15780
rect -2058 -16388 -2024 -16372
rect -1040 -15796 -1006 -15780
rect -1040 -16388 -1006 -16372
rect -22 -15796 12 -15780
rect 2582 -16068 2616 -16052
rect 3600 -15476 3634 -15460
rect 3600 -16068 3634 -16052
rect 4618 -15476 4652 -15460
rect 4618 -16068 4652 -16052
rect 5636 -15476 5670 -15460
rect 5636 -16068 5670 -16052
rect 6654 -15476 6688 -15460
rect 6654 -16068 6688 -16052
rect 7672 -15476 7706 -15460
rect 7672 -16068 7706 -16052
rect 8690 -15476 8724 -15460
rect 8690 -16068 8724 -16052
rect 9708 -15476 9742 -15460
rect 9708 -16068 9742 -16052
rect 10726 -15476 10760 -15460
rect 10726 -16068 10760 -16052
rect 11744 -15476 11778 -15460
rect 11744 -16068 11778 -16052
rect 12762 -15476 12796 -15460
rect 12762 -16068 12796 -16052
rect 13780 -15476 13814 -15460
rect 13780 -16068 13814 -16052
rect 14798 -15476 14832 -15460
rect 14798 -16068 14832 -16052
rect 15816 -15476 15850 -15460
rect 15816 -16068 15850 -16052
rect 16834 -15476 16868 -15460
rect 16834 -16068 16868 -16052
rect 17852 -15476 17886 -15460
rect 17852 -16068 17886 -16052
rect 18870 -15476 18904 -15460
rect 18870 -16068 18904 -16052
rect 19888 -15476 19922 -15460
rect 19888 -16068 19922 -16052
rect 20906 -15476 20940 -15460
rect 20906 -16068 20940 -16052
rect 21924 -15476 21958 -15460
rect 21924 -16068 21958 -16052
rect 22942 -15476 22976 -15460
rect 22976 -16052 22982 -16004
rect 22942 -16068 22976 -16052
rect 6126 -16102 6186 -16100
rect 2814 -16136 2830 -16102
rect 3386 -16136 3402 -16102
rect 3832 -16136 3848 -16102
rect 4404 -16136 4420 -16102
rect 4850 -16136 4866 -16102
rect 5422 -16136 5438 -16102
rect 5868 -16136 5884 -16102
rect 6440 -16136 6456 -16102
rect 6886 -16136 6902 -16102
rect 7458 -16136 7474 -16102
rect 7904 -16136 7920 -16102
rect 8476 -16136 8492 -16102
rect 8922 -16136 8938 -16102
rect 9494 -16136 9510 -16102
rect 9940 -16136 9956 -16102
rect 10512 -16136 10528 -16102
rect 10958 -16136 10974 -16102
rect 11530 -16136 11546 -16102
rect 11976 -16136 11992 -16102
rect 12548 -16136 12564 -16102
rect 12994 -16136 13010 -16102
rect 13566 -16136 13582 -16102
rect 14012 -16136 14028 -16102
rect 14584 -16136 14600 -16102
rect 15030 -16136 15046 -16102
rect 15602 -16136 15618 -16102
rect 16048 -16136 16064 -16102
rect 16620 -16136 16636 -16102
rect 17066 -16136 17082 -16102
rect 17638 -16136 17654 -16102
rect 18084 -16136 18100 -16102
rect 18656 -16136 18672 -16102
rect 19102 -16136 19118 -16102
rect 19674 -16136 19690 -16102
rect 20120 -16136 20136 -16102
rect 20692 -16136 20708 -16102
rect 21138 -16136 21154 -16102
rect 21710 -16136 21726 -16102
rect 22156 -16136 22172 -16102
rect 22728 -16136 22744 -16102
rect 8160 -16140 8220 -16136
rect 17318 -16150 17378 -16136
rect 18352 -16150 18412 -16136
rect -22 -16388 12 -16372
rect 3074 -16352 3156 -16328
rect 3074 -16386 3098 -16352
rect 3132 -16386 3156 -16352
rect 3074 -16410 3156 -16386
rect 4092 -16352 4174 -16328
rect 4092 -16386 4116 -16352
rect 4150 -16386 4174 -16352
rect 4092 -16410 4174 -16386
rect 5110 -16352 5192 -16328
rect 5110 -16386 5134 -16352
rect 5168 -16386 5192 -16352
rect 5110 -16410 5192 -16386
rect 6128 -16352 6210 -16328
rect 6128 -16386 6152 -16352
rect 6186 -16386 6210 -16352
rect 6128 -16410 6210 -16386
rect 7146 -16352 7228 -16328
rect 7146 -16386 7170 -16352
rect 7204 -16386 7228 -16352
rect 7146 -16410 7228 -16386
rect 8164 -16352 8246 -16328
rect 8164 -16386 8188 -16352
rect 8222 -16386 8246 -16352
rect 8164 -16410 8246 -16386
rect 9182 -16352 9264 -16328
rect 9182 -16386 9206 -16352
rect 9240 -16386 9264 -16352
rect 9182 -16410 9264 -16386
rect 10200 -16352 10282 -16328
rect 10200 -16386 10224 -16352
rect 10258 -16386 10282 -16352
rect 10200 -16410 10282 -16386
rect 11218 -16352 11300 -16328
rect 11218 -16386 11242 -16352
rect 11276 -16386 11300 -16352
rect 11218 -16410 11300 -16386
rect 12236 -16352 12318 -16328
rect 12236 -16386 12260 -16352
rect 12294 -16386 12318 -16352
rect 12236 -16410 12318 -16386
rect 13254 -16352 13336 -16328
rect 13254 -16386 13278 -16352
rect 13312 -16386 13336 -16352
rect 13254 -16410 13336 -16386
rect 14272 -16352 14354 -16328
rect 14272 -16386 14296 -16352
rect 14330 -16386 14354 -16352
rect 14272 -16410 14354 -16386
rect 15290 -16352 15372 -16328
rect 15290 -16386 15314 -16352
rect 15348 -16386 15372 -16352
rect 15290 -16410 15372 -16386
rect 16308 -16352 16390 -16328
rect 16308 -16386 16332 -16352
rect 16366 -16386 16390 -16352
rect 16308 -16410 16390 -16386
rect 17326 -16352 17408 -16328
rect 17326 -16386 17350 -16352
rect 17384 -16386 17408 -16352
rect 17326 -16410 17408 -16386
rect 18344 -16352 18426 -16328
rect 18344 -16386 18368 -16352
rect 18402 -16386 18426 -16352
rect 18344 -16410 18426 -16386
rect 19362 -16352 19444 -16328
rect 19362 -16386 19386 -16352
rect 19420 -16386 19444 -16352
rect 19362 -16410 19444 -16386
rect 20380 -16352 20462 -16328
rect 20380 -16386 20404 -16352
rect 20438 -16386 20462 -16352
rect 20380 -16410 20462 -16386
rect 21398 -16352 21480 -16328
rect 21398 -16386 21422 -16352
rect 21456 -16386 21480 -16352
rect 21398 -16410 21480 -16386
rect 22416 -16352 22498 -16328
rect 22416 -16386 22440 -16352
rect 22474 -16386 22498 -16352
rect 22416 -16410 22498 -16386
rect -7670 -16422 -7610 -16420
rect -6656 -16422 -6596 -16420
rect -2582 -16422 -2522 -16420
rect -1566 -16422 -1506 -16420
rect -9208 -16476 -9126 -16452
rect -8952 -16456 -8936 -16422
rect -8380 -16456 -8364 -16422
rect -9208 -16510 -9184 -16476
rect -9150 -16510 -9126 -16476
rect -9208 -16534 -9126 -16510
rect -8190 -16476 -8108 -16452
rect -7934 -16456 -7918 -16422
rect -7362 -16456 -7346 -16422
rect -8190 -16510 -8166 -16476
rect -8132 -16510 -8108 -16476
rect -8952 -16564 -8936 -16530
rect -8380 -16564 -8364 -16530
rect -8190 -16534 -8108 -16510
rect -7172 -16476 -7090 -16452
rect -6916 -16456 -6900 -16422
rect -6344 -16456 -6328 -16422
rect -7172 -16510 -7148 -16476
rect -7114 -16510 -7090 -16476
rect -7934 -16564 -7918 -16530
rect -7362 -16564 -7346 -16530
rect -7172 -16534 -7090 -16510
rect -6154 -16476 -6072 -16452
rect -5898 -16456 -5882 -16422
rect -5326 -16456 -5310 -16422
rect -6154 -16510 -6130 -16476
rect -6096 -16510 -6072 -16476
rect -6916 -16564 -6900 -16530
rect -6344 -16564 -6328 -16530
rect -6154 -16534 -6072 -16510
rect -5136 -16476 -5054 -16452
rect -4880 -16456 -4864 -16422
rect -4308 -16456 -4292 -16422
rect -5136 -16510 -5112 -16476
rect -5078 -16510 -5054 -16476
rect -5898 -16564 -5882 -16530
rect -5326 -16564 -5310 -16530
rect -5136 -16534 -5054 -16510
rect -4118 -16476 -4036 -16452
rect -3862 -16456 -3846 -16422
rect -3290 -16456 -3274 -16422
rect -4118 -16510 -4094 -16476
rect -4060 -16510 -4036 -16476
rect -4880 -16564 -4864 -16530
rect -4308 -16564 -4292 -16530
rect -4118 -16534 -4036 -16510
rect -3100 -16476 -3018 -16452
rect -2844 -16456 -2828 -16422
rect -2272 -16456 -2256 -16422
rect -3100 -16510 -3076 -16476
rect -3042 -16510 -3018 -16476
rect -3862 -16564 -3846 -16530
rect -3290 -16564 -3274 -16530
rect -3100 -16534 -3018 -16510
rect -2082 -16476 -2000 -16452
rect -1826 -16456 -1810 -16422
rect -1254 -16456 -1238 -16422
rect -2082 -16510 -2058 -16476
rect -2024 -16510 -2000 -16476
rect -2844 -16564 -2828 -16530
rect -2272 -16564 -2256 -16530
rect -2082 -16534 -2000 -16510
rect -1064 -16476 -982 -16452
rect -808 -16456 -792 -16422
rect -236 -16456 -220 -16422
rect -1064 -16510 -1040 -16476
rect -1006 -16510 -982 -16476
rect -1826 -16564 -1810 -16530
rect -1254 -16564 -1238 -16530
rect -1064 -16534 -982 -16510
rect -36 -16476 46 -16452
rect -36 -16510 -12 -16476
rect 22 -16510 46 -16476
rect -808 -16564 -792 -16530
rect -236 -16564 -220 -16530
rect -36 -16534 46 -16510
rect -9184 -16614 -9150 -16598
rect -9184 -17206 -9150 -17190
rect -8166 -16614 -8132 -16598
rect -8166 -17206 -8132 -17190
rect -7148 -16614 -7114 -16598
rect -7148 -17206 -7114 -17190
rect -6130 -16614 -6096 -16598
rect -6130 -17206 -6096 -17190
rect -5112 -16614 -5078 -16598
rect -5112 -17206 -5078 -17190
rect -4094 -16614 -4060 -16598
rect -4094 -17206 -4060 -17190
rect -3076 -16614 -3042 -16598
rect -3076 -17206 -3042 -17190
rect -2058 -16614 -2024 -16598
rect -2058 -17206 -2024 -17190
rect -1040 -16614 -1006 -16598
rect -1040 -17206 -1006 -17190
rect -22 -16614 12 -16598
rect 2812 -16660 2828 -16626
rect 3384 -16660 3400 -16626
rect 3830 -16660 3846 -16626
rect 4402 -16660 4418 -16626
rect 4848 -16660 4864 -16626
rect 5420 -16660 5436 -16626
rect 5866 -16660 5882 -16626
rect 6438 -16660 6454 -16626
rect 6884 -16660 6900 -16626
rect 7456 -16660 7472 -16626
rect 7902 -16660 7918 -16626
rect 8474 -16660 8490 -16626
rect 8920 -16660 8936 -16626
rect 9492 -16660 9508 -16626
rect 9938 -16660 9954 -16626
rect 10510 -16660 10526 -16626
rect 10956 -16660 10972 -16626
rect 11528 -16660 11544 -16626
rect 11974 -16660 11990 -16626
rect 12546 -16660 12562 -16626
rect 12992 -16660 13008 -16626
rect 13564 -16660 13580 -16626
rect 14010 -16660 14026 -16626
rect 14582 -16660 14598 -16626
rect 15028 -16660 15044 -16626
rect 15600 -16660 15616 -16626
rect 16046 -16660 16062 -16626
rect 16618 -16660 16634 -16626
rect 17064 -16660 17080 -16626
rect 17636 -16660 17652 -16626
rect 18082 -16660 18098 -16626
rect 18654 -16660 18670 -16626
rect 19100 -16660 19116 -16626
rect 19672 -16660 19688 -16626
rect 20118 -16660 20134 -16626
rect 20690 -16660 20706 -16626
rect 21136 -16660 21152 -16626
rect 21708 -16660 21724 -16626
rect 22154 -16660 22170 -16626
rect 22726 -16660 22742 -16626
rect 5122 -16664 5182 -16660
rect -22 -17206 12 -17190
rect 2580 -16710 2614 -16694
rect -7666 -17240 -7606 -17238
rect -6652 -17240 -6592 -17238
rect -2578 -17240 -2518 -17238
rect -1562 -17240 -1502 -17238
rect -9208 -17294 -9126 -17270
rect -8952 -17274 -8936 -17240
rect -8380 -17274 -8364 -17240
rect -9208 -17328 -9184 -17294
rect -9150 -17328 -9126 -17294
rect -9208 -17352 -9126 -17328
rect -8190 -17294 -8108 -17270
rect -7934 -17274 -7918 -17240
rect -7362 -17274 -7346 -17240
rect -8190 -17328 -8166 -17294
rect -8132 -17328 -8108 -17294
rect -8952 -17382 -8936 -17348
rect -8380 -17382 -8364 -17348
rect -8190 -17352 -8108 -17328
rect -7172 -17294 -7090 -17270
rect -6916 -17274 -6900 -17240
rect -6344 -17274 -6328 -17240
rect -7172 -17328 -7148 -17294
rect -7114 -17328 -7090 -17294
rect -7934 -17382 -7918 -17348
rect -7362 -17382 -7346 -17348
rect -7172 -17352 -7090 -17328
rect -6154 -17294 -6072 -17270
rect -5898 -17274 -5882 -17240
rect -5326 -17274 -5310 -17240
rect -6154 -17328 -6130 -17294
rect -6096 -17328 -6072 -17294
rect -6916 -17382 -6900 -17348
rect -6344 -17382 -6328 -17348
rect -6154 -17352 -6072 -17328
rect -5136 -17294 -5054 -17270
rect -4880 -17274 -4864 -17240
rect -4308 -17274 -4292 -17240
rect -5136 -17328 -5112 -17294
rect -5078 -17328 -5054 -17294
rect -5898 -17382 -5882 -17348
rect -5326 -17382 -5310 -17348
rect -5136 -17352 -5054 -17328
rect -4118 -17294 -4036 -17270
rect -3862 -17274 -3846 -17240
rect -3290 -17274 -3274 -17240
rect -4118 -17328 -4094 -17294
rect -4060 -17328 -4036 -17294
rect -4880 -17382 -4864 -17348
rect -4308 -17382 -4292 -17348
rect -4118 -17352 -4036 -17328
rect -3100 -17294 -3018 -17270
rect -2844 -17274 -2828 -17240
rect -2272 -17274 -2256 -17240
rect -3100 -17328 -3076 -17294
rect -3042 -17328 -3018 -17294
rect -3862 -17382 -3846 -17348
rect -3290 -17382 -3274 -17348
rect -3100 -17352 -3018 -17328
rect -2082 -17294 -2000 -17270
rect -1826 -17274 -1810 -17240
rect -1254 -17274 -1238 -17240
rect -2082 -17328 -2058 -17294
rect -2024 -17328 -2000 -17294
rect -2844 -17382 -2828 -17348
rect -2272 -17382 -2256 -17348
rect -2082 -17352 -2000 -17328
rect -1064 -17294 -982 -17270
rect -808 -17274 -792 -17240
rect -236 -17274 -220 -17240
rect -1064 -17328 -1040 -17294
rect -1006 -17328 -982 -17294
rect -1826 -17382 -1810 -17348
rect -1254 -17382 -1238 -17348
rect -1064 -17352 -982 -17328
rect -36 -17294 46 -17270
rect -36 -17328 -12 -17294
rect 22 -17328 46 -17294
rect 2580 -17302 2614 -17286
rect 3598 -16710 3632 -16694
rect 3598 -17302 3632 -17286
rect 4616 -16710 4650 -16694
rect 4616 -17302 4650 -17286
rect 5634 -16710 5668 -16694
rect 5634 -17302 5668 -17286
rect 6652 -16710 6686 -16694
rect 6652 -17302 6686 -17286
rect 7670 -16710 7704 -16694
rect 7670 -17302 7704 -17286
rect 8688 -16710 8722 -16694
rect 8688 -17302 8722 -17286
rect 9706 -16710 9740 -16694
rect 9706 -17302 9740 -17286
rect 10724 -16710 10758 -16694
rect 10724 -17302 10758 -17286
rect 11742 -16710 11776 -16694
rect 11742 -17302 11776 -17286
rect 12760 -16710 12794 -16694
rect 12760 -17302 12794 -17286
rect 13778 -16710 13812 -16694
rect 13778 -17302 13812 -17286
rect 14796 -16710 14830 -16694
rect 14796 -17302 14830 -17286
rect 15814 -16710 15848 -16694
rect 15814 -17302 15848 -17286
rect 16832 -16710 16866 -16694
rect 16832 -17302 16866 -17286
rect 17850 -16710 17884 -16694
rect 17850 -17302 17884 -17286
rect 18868 -16710 18902 -16694
rect 18868 -17302 18902 -17286
rect 19886 -16710 19920 -16694
rect 19886 -17302 19920 -17286
rect 20904 -16710 20938 -16694
rect 20904 -17302 20938 -17286
rect 21922 -16710 21956 -16694
rect 21922 -17302 21956 -17286
rect 22940 -16710 22974 -16694
rect 22940 -17302 22974 -17286
rect -808 -17382 -792 -17348
rect -236 -17382 -220 -17348
rect -36 -17352 46 -17328
rect 10190 -17336 10250 -17332
rect 11218 -17336 11278 -17334
rect 13262 -17336 13322 -17332
rect 2812 -17370 2828 -17336
rect 3384 -17370 3400 -17336
rect 3830 -17370 3846 -17336
rect 4402 -17370 4418 -17336
rect 4848 -17370 4864 -17336
rect 5420 -17370 5436 -17336
rect 5866 -17370 5882 -17336
rect 6438 -17370 6454 -17336
rect 6884 -17370 6900 -17336
rect 7456 -17370 7472 -17336
rect 7902 -17370 7918 -17336
rect 8474 -17370 8490 -17336
rect 8920 -17370 8936 -17336
rect 9492 -17370 9508 -17336
rect 9938 -17370 9954 -17336
rect 10510 -17370 10526 -17336
rect 10956 -17370 10972 -17336
rect 11528 -17370 11544 -17336
rect 11974 -17370 11990 -17336
rect 12546 -17370 12562 -17336
rect 12992 -17370 13008 -17336
rect 13564 -17370 13580 -17336
rect 14010 -17370 14026 -17336
rect 14582 -17370 14598 -17336
rect 15028 -17370 15044 -17336
rect 15600 -17370 15616 -17336
rect 16046 -17370 16062 -17336
rect 16618 -17370 16634 -17336
rect 17064 -17370 17080 -17336
rect 17636 -17370 17652 -17336
rect 18082 -17370 18098 -17336
rect 18654 -17370 18670 -17336
rect 19100 -17370 19116 -17336
rect 19672 -17370 19688 -17336
rect 20118 -17370 20134 -17336
rect 20690 -17370 20706 -17336
rect 21136 -17370 21152 -17336
rect 21708 -17370 21724 -17336
rect 22154 -17370 22170 -17336
rect 22726 -17370 22742 -17336
rect -9184 -17432 -9150 -17416
rect -9184 -18024 -9150 -18008
rect -8166 -17432 -8132 -17416
rect -8166 -18024 -8132 -18008
rect -7148 -17432 -7114 -17416
rect -7148 -18024 -7114 -18008
rect -6130 -17432 -6096 -17416
rect -6130 -18024 -6096 -18008
rect -5112 -17432 -5078 -17416
rect -5112 -18024 -5078 -18008
rect -4094 -17432 -4060 -17416
rect -4094 -18024 -4060 -18008
rect -3076 -17432 -3042 -17416
rect -3076 -18024 -3042 -18008
rect -2058 -17432 -2024 -17416
rect -2058 -18024 -2024 -18008
rect -1040 -17432 -1006 -17416
rect -1040 -18024 -1006 -18008
rect -22 -17432 12 -17416
rect 3074 -17576 3156 -17552
rect 3074 -17610 3098 -17576
rect 3132 -17610 3156 -17576
rect 3074 -17634 3156 -17610
rect 4092 -17576 4174 -17552
rect 4092 -17610 4116 -17576
rect 4150 -17610 4174 -17576
rect 4092 -17634 4174 -17610
rect 5110 -17576 5192 -17552
rect 5110 -17610 5134 -17576
rect 5168 -17610 5192 -17576
rect 5110 -17634 5192 -17610
rect 6128 -17576 6210 -17552
rect 6128 -17610 6152 -17576
rect 6186 -17610 6210 -17576
rect 6128 -17634 6210 -17610
rect 7146 -17576 7228 -17552
rect 7146 -17610 7170 -17576
rect 7204 -17610 7228 -17576
rect 7146 -17634 7228 -17610
rect 8164 -17576 8246 -17552
rect 8164 -17610 8188 -17576
rect 8222 -17610 8246 -17576
rect 8164 -17634 8246 -17610
rect 9182 -17576 9264 -17552
rect 9182 -17610 9206 -17576
rect 9240 -17610 9264 -17576
rect 9182 -17634 9264 -17610
rect 10200 -17576 10282 -17552
rect 10200 -17610 10224 -17576
rect 10258 -17610 10282 -17576
rect 10200 -17634 10282 -17610
rect 11218 -17576 11300 -17552
rect 11218 -17610 11242 -17576
rect 11276 -17610 11300 -17576
rect 11218 -17634 11300 -17610
rect 12236 -17576 12318 -17552
rect 12236 -17610 12260 -17576
rect 12294 -17610 12318 -17576
rect 12236 -17634 12318 -17610
rect 13254 -17576 13336 -17552
rect 13254 -17610 13278 -17576
rect 13312 -17610 13336 -17576
rect 13254 -17634 13336 -17610
rect 14272 -17576 14354 -17552
rect 14272 -17610 14296 -17576
rect 14330 -17610 14354 -17576
rect 14272 -17634 14354 -17610
rect 15290 -17576 15372 -17552
rect 15290 -17610 15314 -17576
rect 15348 -17610 15372 -17576
rect 15290 -17634 15372 -17610
rect 16308 -17576 16390 -17552
rect 16308 -17610 16332 -17576
rect 16366 -17610 16390 -17576
rect 16308 -17634 16390 -17610
rect 17326 -17576 17408 -17552
rect 17326 -17610 17350 -17576
rect 17384 -17610 17408 -17576
rect 17326 -17634 17408 -17610
rect 18344 -17576 18426 -17552
rect 18344 -17610 18368 -17576
rect 18402 -17610 18426 -17576
rect 18344 -17634 18426 -17610
rect 19362 -17576 19444 -17552
rect 19362 -17610 19386 -17576
rect 19420 -17610 19444 -17576
rect 19362 -17634 19444 -17610
rect 20380 -17576 20462 -17552
rect 20380 -17610 20404 -17576
rect 20438 -17610 20462 -17576
rect 20380 -17634 20462 -17610
rect 21398 -17576 21480 -17552
rect 21398 -17610 21422 -17576
rect 21456 -17610 21480 -17576
rect 21398 -17634 21480 -17610
rect 22416 -17576 22498 -17552
rect 22416 -17610 22440 -17576
rect 22474 -17610 22498 -17576
rect 22416 -17634 22498 -17610
rect 2812 -17894 2828 -17860
rect 3384 -17894 3400 -17860
rect 3830 -17894 3846 -17860
rect 4402 -17894 4418 -17860
rect 4848 -17894 4864 -17860
rect 5420 -17894 5436 -17860
rect 5866 -17894 5882 -17860
rect 6438 -17894 6454 -17860
rect 6884 -17894 6900 -17860
rect 7456 -17894 7472 -17860
rect 7902 -17894 7918 -17860
rect 8474 -17894 8490 -17860
rect 8920 -17894 8936 -17860
rect 9492 -17894 9508 -17860
rect 9938 -17894 9954 -17860
rect 10510 -17894 10526 -17860
rect 10956 -17894 10972 -17860
rect 11528 -17894 11544 -17860
rect 11974 -17894 11990 -17860
rect 12546 -17894 12562 -17860
rect 12992 -17894 13008 -17860
rect 13564 -17894 13580 -17860
rect 14010 -17894 14026 -17860
rect 14582 -17894 14598 -17860
rect 15028 -17894 15044 -17860
rect 15600 -17894 15616 -17860
rect 16046 -17894 16062 -17860
rect 16618 -17894 16634 -17860
rect 17064 -17894 17080 -17860
rect 17636 -17894 17652 -17860
rect 18082 -17894 18098 -17860
rect 18654 -17894 18670 -17860
rect 19100 -17894 19116 -17860
rect 19672 -17894 19688 -17860
rect 20118 -17894 20134 -17860
rect 20690 -17894 20706 -17860
rect 21136 -17894 21152 -17860
rect 21708 -17894 21724 -17860
rect 22154 -17894 22170 -17860
rect 22726 -17894 22742 -17860
rect -22 -18024 12 -18008
rect 2580 -17944 2614 -17928
rect -8692 -18058 -8632 -18056
rect -7666 -18058 -7606 -18054
rect -6652 -18058 -6592 -18054
rect -5632 -18058 -5572 -18056
rect -4610 -18058 -4550 -18056
rect -2578 -18058 -2518 -18054
rect -1562 -18058 -1502 -18054
rect -542 -18058 -482 -18056
rect -9208 -18112 -9126 -18088
rect -8952 -18092 -8936 -18058
rect -8380 -18092 -8364 -18058
rect -9208 -18146 -9184 -18112
rect -9150 -18146 -9126 -18112
rect -9208 -18170 -9126 -18146
rect -8190 -18112 -8108 -18088
rect -7934 -18092 -7918 -18058
rect -7362 -18092 -7346 -18058
rect -8190 -18146 -8166 -18112
rect -8132 -18146 -8108 -18112
rect -8952 -18200 -8936 -18166
rect -8380 -18200 -8364 -18166
rect -8190 -18170 -8108 -18146
rect -7172 -18112 -7090 -18088
rect -6916 -18092 -6900 -18058
rect -6344 -18092 -6328 -18058
rect -7172 -18146 -7148 -18112
rect -7114 -18146 -7090 -18112
rect -7934 -18200 -7918 -18166
rect -7362 -18200 -7346 -18166
rect -7172 -18170 -7090 -18146
rect -6154 -18112 -6072 -18088
rect -5898 -18092 -5882 -18058
rect -5326 -18092 -5310 -18058
rect -6154 -18146 -6130 -18112
rect -6096 -18146 -6072 -18112
rect -6916 -18200 -6900 -18166
rect -6344 -18200 -6328 -18166
rect -6154 -18170 -6072 -18146
rect -5136 -18112 -5054 -18088
rect -4880 -18092 -4864 -18058
rect -4308 -18092 -4292 -18058
rect -5136 -18146 -5112 -18112
rect -5078 -18146 -5054 -18112
rect -5898 -18200 -5882 -18166
rect -5326 -18200 -5310 -18166
rect -5136 -18170 -5054 -18146
rect -4118 -18112 -4036 -18088
rect -3862 -18092 -3846 -18058
rect -3290 -18092 -3274 -18058
rect -4118 -18146 -4094 -18112
rect -4060 -18146 -4036 -18112
rect -4880 -18200 -4864 -18166
rect -4308 -18200 -4292 -18166
rect -4118 -18170 -4036 -18146
rect -3100 -18112 -3018 -18088
rect -2844 -18092 -2828 -18058
rect -2272 -18092 -2256 -18058
rect -3100 -18146 -3076 -18112
rect -3042 -18146 -3018 -18112
rect -3862 -18200 -3846 -18166
rect -3290 -18200 -3274 -18166
rect -3100 -18170 -3018 -18146
rect -2082 -18112 -2000 -18088
rect -1826 -18092 -1810 -18058
rect -1254 -18092 -1238 -18058
rect -2082 -18146 -2058 -18112
rect -2024 -18146 -2000 -18112
rect -2844 -18200 -2828 -18166
rect -2272 -18200 -2256 -18166
rect -2082 -18170 -2000 -18146
rect -1064 -18112 -982 -18088
rect -808 -18092 -792 -18058
rect -236 -18092 -220 -18058
rect -1064 -18146 -1040 -18112
rect -1006 -18146 -982 -18112
rect -1826 -18200 -1810 -18166
rect -1254 -18200 -1238 -18166
rect -1064 -18170 -982 -18146
rect -36 -18112 46 -18088
rect -36 -18146 -12 -18112
rect 22 -18146 46 -18112
rect -808 -18200 -792 -18166
rect -236 -18200 -220 -18166
rect -36 -18170 46 -18146
rect -9184 -18250 -9150 -18234
rect -9184 -18842 -9150 -18826
rect -8166 -18250 -8132 -18234
rect -8166 -18842 -8132 -18826
rect -7148 -18250 -7114 -18234
rect -7148 -18842 -7114 -18826
rect -6130 -18250 -6096 -18234
rect -6130 -18842 -6096 -18826
rect -5112 -18250 -5078 -18234
rect -5112 -18842 -5078 -18826
rect -4094 -18250 -4060 -18234
rect -4094 -18842 -4060 -18826
rect -3076 -18250 -3042 -18234
rect -3076 -18842 -3042 -18826
rect -2058 -18250 -2024 -18234
rect -2058 -18842 -2024 -18826
rect -1040 -18250 -1006 -18234
rect -1040 -18842 -1006 -18826
rect -22 -18250 12 -18234
rect 2580 -18536 2614 -18520
rect 3598 -17944 3632 -17928
rect 3598 -18536 3632 -18520
rect 4616 -17944 4650 -17928
rect 4616 -18536 4650 -18520
rect 5634 -17944 5668 -17928
rect 5634 -18536 5668 -18520
rect 6652 -17944 6686 -17928
rect 6652 -18536 6686 -18520
rect 7670 -17944 7704 -17928
rect 7670 -18536 7704 -18520
rect 8688 -17944 8722 -17928
rect 8688 -18536 8722 -18520
rect 9706 -17944 9740 -17928
rect 9706 -18536 9740 -18520
rect 10724 -17944 10758 -17928
rect 10724 -18536 10758 -18520
rect 11742 -17944 11776 -17928
rect 11742 -18536 11776 -18520
rect 12760 -17944 12794 -17928
rect 12760 -18536 12794 -18520
rect 13778 -17944 13812 -17928
rect 13778 -18536 13812 -18520
rect 14796 -17944 14830 -17928
rect 14796 -18536 14830 -18520
rect 15814 -17944 15848 -17928
rect 15814 -18536 15848 -18520
rect 16832 -17944 16866 -17928
rect 16832 -18536 16866 -18520
rect 17850 -17944 17884 -17928
rect 17850 -18536 17884 -18520
rect 18868 -17944 18902 -17928
rect 18868 -18536 18902 -18520
rect 19886 -17944 19920 -17928
rect 19886 -18536 19920 -18520
rect 20904 -17944 20938 -17928
rect 20904 -18536 20938 -18520
rect 21922 -17944 21956 -17928
rect 21922 -18536 21956 -18520
rect 22940 -17944 22974 -17928
rect 22940 -18536 22974 -18520
rect 2812 -18604 2828 -18570
rect 3384 -18604 3400 -18570
rect 3830 -18604 3846 -18570
rect 4402 -18604 4418 -18570
rect 4848 -18604 4864 -18570
rect 5420 -18604 5436 -18570
rect 5866 -18604 5882 -18570
rect 6438 -18604 6454 -18570
rect 6884 -18604 6900 -18570
rect 7456 -18604 7472 -18570
rect 7902 -18604 7918 -18570
rect 8474 -18604 8490 -18570
rect 8920 -18604 8936 -18570
rect 9492 -18604 9508 -18570
rect 9938 -18604 9954 -18570
rect 10510 -18604 10526 -18570
rect 10956 -18604 10972 -18570
rect 11528 -18604 11544 -18570
rect 11974 -18604 11990 -18570
rect 12546 -18604 12562 -18570
rect 12992 -18604 13008 -18570
rect 13564 -18604 13580 -18570
rect 14010 -18604 14026 -18570
rect 14582 -18604 14598 -18570
rect 15028 -18604 15044 -18570
rect 15600 -18604 15616 -18570
rect 16046 -18604 16062 -18570
rect 16618 -18604 16634 -18570
rect 17064 -18604 17080 -18570
rect 17636 -18604 17652 -18570
rect 18082 -18604 18098 -18570
rect 18654 -18604 18670 -18570
rect 19100 -18604 19116 -18570
rect 19672 -18604 19688 -18570
rect 20118 -18604 20134 -18570
rect 20690 -18604 20706 -18570
rect 21136 -18604 21152 -18570
rect 21708 -18604 21724 -18570
rect 22154 -18604 22170 -18570
rect 22726 -18604 22742 -18570
rect -22 -18842 12 -18826
rect 3086 -18812 3168 -18788
rect 3086 -18846 3110 -18812
rect 3144 -18846 3168 -18812
rect 3086 -18870 3168 -18846
rect 4104 -18812 4186 -18788
rect 4104 -18846 4128 -18812
rect 4162 -18846 4186 -18812
rect 4104 -18870 4186 -18846
rect 5122 -18812 5204 -18788
rect 5122 -18846 5146 -18812
rect 5180 -18846 5204 -18812
rect 5122 -18870 5204 -18846
rect 6140 -18812 6222 -18788
rect 6140 -18846 6164 -18812
rect 6198 -18846 6222 -18812
rect 6140 -18870 6222 -18846
rect 7158 -18812 7240 -18788
rect 7158 -18846 7182 -18812
rect 7216 -18846 7240 -18812
rect 7158 -18870 7240 -18846
rect 8176 -18812 8258 -18788
rect 8176 -18846 8200 -18812
rect 8234 -18846 8258 -18812
rect 8176 -18870 8258 -18846
rect 9194 -18812 9276 -18788
rect 9194 -18846 9218 -18812
rect 9252 -18846 9276 -18812
rect 9194 -18870 9276 -18846
rect 10212 -18812 10294 -18788
rect 10212 -18846 10236 -18812
rect 10270 -18846 10294 -18812
rect 10212 -18870 10294 -18846
rect 11230 -18812 11312 -18788
rect 11230 -18846 11254 -18812
rect 11288 -18846 11312 -18812
rect 11230 -18870 11312 -18846
rect 12248 -18812 12330 -18788
rect 12248 -18846 12272 -18812
rect 12306 -18846 12330 -18812
rect 12248 -18870 12330 -18846
rect 13266 -18812 13348 -18788
rect 13266 -18846 13290 -18812
rect 13324 -18846 13348 -18812
rect 13266 -18870 13348 -18846
rect 14284 -18812 14366 -18788
rect 14284 -18846 14308 -18812
rect 14342 -18846 14366 -18812
rect 14284 -18870 14366 -18846
rect 15302 -18812 15384 -18788
rect 15302 -18846 15326 -18812
rect 15360 -18846 15384 -18812
rect 15302 -18870 15384 -18846
rect 16320 -18812 16402 -18788
rect 16320 -18846 16344 -18812
rect 16378 -18846 16402 -18812
rect 16320 -18870 16402 -18846
rect 17338 -18812 17420 -18788
rect 17338 -18846 17362 -18812
rect 17396 -18846 17420 -18812
rect 17338 -18870 17420 -18846
rect 18356 -18812 18438 -18788
rect 18356 -18846 18380 -18812
rect 18414 -18846 18438 -18812
rect 18356 -18870 18438 -18846
rect 19374 -18812 19456 -18788
rect 19374 -18846 19398 -18812
rect 19432 -18846 19456 -18812
rect 19374 -18870 19456 -18846
rect 20392 -18812 20474 -18788
rect 20392 -18846 20416 -18812
rect 20450 -18846 20474 -18812
rect 20392 -18870 20474 -18846
rect 21410 -18812 21492 -18788
rect 21410 -18846 21434 -18812
rect 21468 -18846 21492 -18812
rect 21410 -18870 21492 -18846
rect 22428 -18812 22510 -18788
rect 22428 -18846 22452 -18812
rect 22486 -18846 22510 -18812
rect 22428 -18870 22510 -18846
rect -8952 -18910 -8936 -18876
rect -8380 -18910 -8364 -18876
rect -7934 -18910 -7918 -18876
rect -7362 -18910 -7346 -18876
rect -6916 -18910 -6900 -18876
rect -6344 -18910 -6328 -18876
rect -5898 -18910 -5882 -18876
rect -5326 -18910 -5310 -18876
rect -4880 -18910 -4864 -18876
rect -4308 -18910 -4292 -18876
rect -3862 -18910 -3846 -18876
rect -3290 -18910 -3274 -18876
rect -2844 -18910 -2828 -18876
rect -2272 -18910 -2256 -18876
rect -1826 -18910 -1810 -18876
rect -1254 -18910 -1238 -18876
rect -808 -18910 -792 -18876
rect -236 -18910 -220 -18876
rect -9220 -19006 -9138 -18982
rect -9220 -19040 -9196 -19006
rect -9162 -19040 -9138 -19006
rect -9220 -19064 -9138 -19040
rect -8202 -19006 -8120 -18982
rect -8202 -19040 -8178 -19006
rect -8144 -19040 -8120 -19006
rect -8202 -19064 -8120 -19040
rect -7184 -19006 -7102 -18982
rect -7184 -19040 -7160 -19006
rect -7126 -19040 -7102 -19006
rect -7184 -19064 -7102 -19040
rect -6166 -19006 -6084 -18982
rect -6166 -19040 -6142 -19006
rect -6108 -19040 -6084 -19006
rect -6166 -19064 -6084 -19040
rect -5148 -19006 -5066 -18982
rect -5148 -19040 -5124 -19006
rect -5090 -19040 -5066 -19006
rect -5148 -19064 -5066 -19040
rect -4130 -19006 -4048 -18982
rect -4130 -19040 -4106 -19006
rect -4072 -19040 -4048 -19006
rect -4130 -19064 -4048 -19040
rect -3112 -19006 -3030 -18982
rect -3112 -19040 -3088 -19006
rect -3054 -19040 -3030 -19006
rect -3112 -19064 -3030 -19040
rect -2094 -19006 -2012 -18982
rect -2094 -19040 -2070 -19006
rect -2036 -19040 -2012 -19006
rect -2094 -19064 -2012 -19040
rect -1076 -19006 -994 -18982
rect -1076 -19040 -1052 -19006
rect -1018 -19040 -994 -19006
rect -1076 -19064 -994 -19040
rect -48 -19006 34 -18982
rect -48 -19040 -24 -19006
rect 10 -19040 34 -19006
rect -48 -19064 34 -19040
rect 2812 -19126 2828 -19092
rect 3384 -19126 3400 -19092
rect 3830 -19126 3846 -19092
rect 4402 -19126 4418 -19092
rect 4848 -19126 4864 -19092
rect 5420 -19126 5436 -19092
rect 5866 -19126 5882 -19092
rect 6438 -19126 6454 -19092
rect 6884 -19126 6900 -19092
rect 7456 -19126 7472 -19092
rect 7902 -19126 7918 -19092
rect 8474 -19126 8490 -19092
rect 8920 -19126 8936 -19092
rect 9492 -19126 9508 -19092
rect 9938 -19126 9954 -19092
rect 10510 -19126 10526 -19092
rect 10956 -19126 10972 -19092
rect 11528 -19126 11544 -19092
rect 11974 -19126 11990 -19092
rect 12546 -19126 12562 -19092
rect 12992 -19126 13008 -19092
rect 13564 -19126 13580 -19092
rect 14010 -19126 14026 -19092
rect 14582 -19126 14598 -19092
rect 15028 -19126 15044 -19092
rect 15600 -19126 15616 -19092
rect 16046 -19126 16062 -19092
rect 16618 -19126 16634 -19092
rect 17064 -19126 17080 -19092
rect 17636 -19126 17652 -19092
rect 18082 -19126 18098 -19092
rect 18654 -19126 18670 -19092
rect 19100 -19126 19116 -19092
rect 19672 -19126 19688 -19092
rect 20118 -19126 20134 -19092
rect 20690 -19126 20706 -19092
rect 21136 -19126 21152 -19092
rect 21708 -19126 21724 -19092
rect 22154 -19126 22170 -19092
rect 22726 -19126 22742 -19092
rect 2580 -19176 2614 -19160
rect 2580 -19768 2614 -19752
rect 3598 -19176 3632 -19160
rect 3598 -19768 3632 -19752
rect 4616 -19176 4650 -19160
rect 4616 -19768 4650 -19752
rect 5634 -19176 5668 -19160
rect 5634 -19768 5668 -19752
rect 6652 -19176 6686 -19160
rect 6652 -19768 6686 -19752
rect 7670 -19176 7704 -19160
rect 7670 -19768 7704 -19752
rect 8688 -19176 8722 -19160
rect 8688 -19768 8722 -19752
rect 9706 -19176 9740 -19160
rect 9706 -19768 9740 -19752
rect 10724 -19176 10758 -19160
rect 10724 -19768 10758 -19752
rect 11742 -19176 11776 -19160
rect 11742 -19768 11776 -19752
rect 12760 -19176 12794 -19160
rect 12760 -19768 12794 -19752
rect 13778 -19176 13812 -19160
rect 13778 -19768 13812 -19752
rect 14796 -19176 14830 -19160
rect 14796 -19768 14830 -19752
rect 15814 -19176 15848 -19160
rect 15814 -19768 15848 -19752
rect 16832 -19176 16866 -19160
rect 16832 -19768 16866 -19752
rect 17850 -19176 17884 -19160
rect 17850 -19768 17884 -19752
rect 18868 -19176 18902 -19160
rect 18868 -19768 18902 -19752
rect 19886 -19176 19920 -19160
rect 19886 -19768 19920 -19752
rect 20904 -19176 20938 -19160
rect 20904 -19768 20938 -19752
rect 21922 -19176 21956 -19160
rect 21922 -19768 21956 -19752
rect 22940 -19176 22974 -19160
rect 22940 -19768 22974 -19752
rect 11230 -19802 11290 -19800
rect 13274 -19802 13334 -19798
rect 21408 -19802 21468 -19800
rect 2812 -19836 2828 -19802
rect 3384 -19836 3400 -19802
rect 3830 -19836 3846 -19802
rect 4402 -19836 4418 -19802
rect 4848 -19836 4864 -19802
rect 5420 -19836 5436 -19802
rect 5866 -19836 5882 -19802
rect 6438 -19836 6454 -19802
rect 6884 -19836 6900 -19802
rect 7456 -19836 7472 -19802
rect 7902 -19836 7918 -19802
rect 8474 -19836 8490 -19802
rect 8920 -19836 8936 -19802
rect 9492 -19836 9508 -19802
rect 9938 -19836 9954 -19802
rect 10510 -19836 10526 -19802
rect 10956 -19836 10972 -19802
rect 11528 -19836 11544 -19802
rect 11974 -19836 11990 -19802
rect 12546 -19836 12562 -19802
rect 12992 -19836 13008 -19802
rect 13564 -19836 13580 -19802
rect 14010 -19836 14026 -19802
rect 14582 -19836 14598 -19802
rect 15028 -19836 15044 -19802
rect 15600 -19836 15616 -19802
rect 16046 -19836 16062 -19802
rect 16618 -19836 16634 -19802
rect 17064 -19836 17080 -19802
rect 17636 -19836 17652 -19802
rect 18082 -19836 18098 -19802
rect 18654 -19836 18670 -19802
rect 19100 -19836 19116 -19802
rect 19672 -19836 19688 -19802
rect 20118 -19836 20134 -19802
rect 20690 -19836 20706 -19802
rect 21136 -19836 21152 -19802
rect 21708 -19836 21724 -19802
rect 22154 -19836 22170 -19802
rect 22726 -19836 22742 -19802
rect -10016 -19954 -9934 -19930
rect -10016 -19988 -9992 -19954
rect -9958 -19988 -9934 -19954
rect -10016 -20012 -9934 -19988
rect -8998 -19954 -8916 -19930
rect -8998 -19988 -8974 -19954
rect -8940 -19988 -8916 -19954
rect -8998 -20012 -8916 -19988
rect -7980 -19954 -7898 -19930
rect -7980 -19988 -7956 -19954
rect -7922 -19988 -7898 -19954
rect -7980 -20012 -7898 -19988
rect -6962 -19954 -6880 -19930
rect -6962 -19988 -6938 -19954
rect -6904 -19988 -6880 -19954
rect -6962 -20012 -6880 -19988
rect -5944 -19954 -5862 -19930
rect -5944 -19988 -5920 -19954
rect -5886 -19988 -5862 -19954
rect -5944 -20012 -5862 -19988
rect -4926 -19954 -4844 -19930
rect -4926 -19988 -4902 -19954
rect -4868 -19988 -4844 -19954
rect -4926 -20012 -4844 -19988
rect -3908 -19954 -3826 -19930
rect -3908 -19988 -3884 -19954
rect -3850 -19988 -3826 -19954
rect -3908 -20012 -3826 -19988
rect -2890 -19954 -2808 -19930
rect -2890 -19988 -2866 -19954
rect -2832 -19988 -2808 -19954
rect -2890 -20012 -2808 -19988
rect -1872 -19954 -1790 -19930
rect -1872 -19988 -1848 -19954
rect -1814 -19988 -1790 -19954
rect -1872 -20012 -1790 -19988
rect -854 -19954 -772 -19930
rect -854 -19988 -830 -19954
rect -796 -19988 -772 -19954
rect -854 -20012 -772 -19988
rect 164 -19954 246 -19930
rect 164 -19988 188 -19954
rect 222 -19988 246 -19954
rect 164 -20012 246 -19988
rect 3086 -20060 3168 -20036
rect 3086 -20094 3110 -20060
rect 3144 -20094 3168 -20060
rect 3086 -20118 3168 -20094
rect 4104 -20060 4186 -20036
rect 4104 -20094 4128 -20060
rect 4162 -20094 4186 -20060
rect 4104 -20118 4186 -20094
rect 5122 -20060 5204 -20036
rect 5122 -20094 5146 -20060
rect 5180 -20094 5204 -20060
rect 5122 -20118 5204 -20094
rect 6140 -20060 6222 -20036
rect 6140 -20094 6164 -20060
rect 6198 -20094 6222 -20060
rect 6140 -20118 6222 -20094
rect 7158 -20060 7240 -20036
rect 7158 -20094 7182 -20060
rect 7216 -20094 7240 -20060
rect 7158 -20118 7240 -20094
rect 8176 -20060 8258 -20036
rect 8176 -20094 8200 -20060
rect 8234 -20094 8258 -20060
rect 8176 -20118 8258 -20094
rect 9194 -20060 9276 -20036
rect 9194 -20094 9218 -20060
rect 9252 -20094 9276 -20060
rect 9194 -20118 9276 -20094
rect 10212 -20060 10294 -20036
rect 10212 -20094 10236 -20060
rect 10270 -20094 10294 -20060
rect 10212 -20118 10294 -20094
rect 11230 -20060 11312 -20036
rect 11230 -20094 11254 -20060
rect 11288 -20094 11312 -20060
rect 11230 -20118 11312 -20094
rect 12248 -20060 12330 -20036
rect 12248 -20094 12272 -20060
rect 12306 -20094 12330 -20060
rect 12248 -20118 12330 -20094
rect 13266 -20060 13348 -20036
rect 13266 -20094 13290 -20060
rect 13324 -20094 13348 -20060
rect 13266 -20118 13348 -20094
rect 14284 -20060 14366 -20036
rect 14284 -20094 14308 -20060
rect 14342 -20094 14366 -20060
rect 14284 -20118 14366 -20094
rect 15302 -20060 15384 -20036
rect 15302 -20094 15326 -20060
rect 15360 -20094 15384 -20060
rect 15302 -20118 15384 -20094
rect 16320 -20060 16402 -20036
rect 16320 -20094 16344 -20060
rect 16378 -20094 16402 -20060
rect 16320 -20118 16402 -20094
rect 17338 -20060 17420 -20036
rect 17338 -20094 17362 -20060
rect 17396 -20094 17420 -20060
rect 17338 -20118 17420 -20094
rect 18356 -20060 18438 -20036
rect 18356 -20094 18380 -20060
rect 18414 -20094 18438 -20060
rect 18356 -20118 18438 -20094
rect 19374 -20060 19456 -20036
rect 19374 -20094 19398 -20060
rect 19432 -20094 19456 -20060
rect 19374 -20118 19456 -20094
rect 20392 -20060 20474 -20036
rect 20392 -20094 20416 -20060
rect 20450 -20094 20474 -20060
rect 20392 -20118 20474 -20094
rect 21410 -20060 21492 -20036
rect 21410 -20094 21434 -20060
rect 21468 -20094 21492 -20060
rect 21410 -20118 21492 -20094
rect 22428 -20060 22510 -20036
rect 22428 -20094 22452 -20060
rect 22486 -20094 22510 -20060
rect 22428 -20118 22510 -20094
rect -10276 -20224 -10260 -20190
rect -9704 -20224 -9688 -20190
rect -9258 -20224 -9242 -20190
rect -8686 -20224 -8670 -20190
rect -8240 -20224 -8224 -20190
rect -7668 -20224 -7652 -20190
rect -7222 -20224 -7206 -20190
rect -6650 -20224 -6634 -20190
rect -6204 -20224 -6188 -20190
rect -5632 -20224 -5616 -20190
rect -5186 -20224 -5170 -20190
rect -4614 -20224 -4598 -20190
rect -4168 -20224 -4152 -20190
rect -3596 -20224 -3580 -20190
rect -3150 -20224 -3134 -20190
rect -2578 -20224 -2562 -20190
rect -2132 -20224 -2116 -20190
rect -1560 -20224 -1544 -20190
rect -1114 -20224 -1098 -20190
rect -542 -20224 -526 -20190
rect -96 -20224 -80 -20190
rect 476 -20224 492 -20190
rect -10508 -20274 -10474 -20258
rect -10508 -20866 -10474 -20850
rect -9490 -20274 -9456 -20258
rect -9490 -20866 -9456 -20850
rect -8472 -20274 -8438 -20258
rect -8472 -20866 -8438 -20850
rect -7454 -20274 -7420 -20258
rect -7454 -20866 -7420 -20850
rect -6436 -20274 -6402 -20258
rect -6436 -20866 -6402 -20850
rect -5418 -20274 -5384 -20258
rect -5418 -20866 -5384 -20850
rect -4400 -20274 -4366 -20258
rect -4400 -20866 -4366 -20850
rect -3382 -20274 -3348 -20258
rect -3382 -20866 -3348 -20850
rect -2364 -20274 -2330 -20258
rect -2364 -20866 -2330 -20850
rect -1346 -20274 -1312 -20258
rect -1346 -20866 -1312 -20850
rect -328 -20274 -294 -20258
rect -328 -20866 -294 -20850
rect 690 -20274 724 -20258
rect 2812 -20360 2828 -20326
rect 3384 -20360 3400 -20326
rect 3830 -20360 3846 -20326
rect 4402 -20360 4418 -20326
rect 4848 -20360 4864 -20326
rect 5420 -20360 5436 -20326
rect 5866 -20360 5882 -20326
rect 6438 -20360 6454 -20326
rect 6884 -20360 6900 -20326
rect 7456 -20360 7472 -20326
rect 7902 -20360 7918 -20326
rect 8474 -20360 8490 -20326
rect 8920 -20360 8936 -20326
rect 9492 -20360 9508 -20326
rect 9938 -20360 9954 -20326
rect 10510 -20360 10526 -20326
rect 10956 -20360 10972 -20326
rect 11528 -20360 11544 -20326
rect 11974 -20360 11990 -20326
rect 12546 -20360 12562 -20326
rect 12992 -20360 13008 -20326
rect 13564 -20360 13580 -20326
rect 14010 -20360 14026 -20326
rect 14582 -20360 14598 -20326
rect 15028 -20360 15044 -20326
rect 15600 -20360 15616 -20326
rect 16046 -20360 16062 -20326
rect 16618 -20360 16634 -20326
rect 17064 -20360 17080 -20326
rect 17636 -20360 17652 -20326
rect 18082 -20360 18098 -20326
rect 18654 -20360 18670 -20326
rect 19100 -20360 19116 -20326
rect 19672 -20360 19688 -20326
rect 20118 -20360 20134 -20326
rect 20690 -20360 20706 -20326
rect 21136 -20360 21152 -20326
rect 21708 -20360 21724 -20326
rect 22154 -20360 22170 -20326
rect 22726 -20360 22742 -20326
rect 690 -20866 724 -20850
rect 2580 -20410 2614 -20394
rect -10276 -20934 -10260 -20900
rect -9704 -20934 -9688 -20900
rect -9258 -20934 -9242 -20900
rect -8686 -20934 -8670 -20900
rect -8240 -20934 -8224 -20900
rect -7668 -20934 -7652 -20900
rect -7222 -20934 -7206 -20900
rect -6650 -20934 -6634 -20900
rect -6204 -20934 -6188 -20900
rect -5632 -20934 -5616 -20900
rect -5186 -20934 -5170 -20900
rect -4614 -20934 -4598 -20900
rect -4168 -20934 -4152 -20900
rect -3596 -20934 -3580 -20900
rect -3150 -20934 -3134 -20900
rect -2578 -20934 -2562 -20900
rect -2132 -20934 -2116 -20900
rect -1560 -20934 -1544 -20900
rect -1114 -20934 -1098 -20900
rect -542 -20934 -526 -20900
rect -96 -20934 -80 -20900
rect 476 -20934 492 -20900
rect 2580 -21002 2614 -20986
rect 3598 -20410 3632 -20394
rect 3598 -21002 3632 -20986
rect 4616 -20410 4650 -20394
rect 4616 -21002 4650 -20986
rect 5634 -20410 5668 -20394
rect 5634 -21002 5668 -20986
rect 6652 -20410 6686 -20394
rect 6652 -21002 6686 -20986
rect 7670 -20410 7704 -20394
rect 7670 -21002 7704 -20986
rect 8688 -20410 8722 -20394
rect 8688 -21002 8722 -20986
rect 9706 -20410 9740 -20394
rect 9706 -21002 9740 -20986
rect 10724 -20410 10758 -20394
rect 10724 -21002 10758 -20986
rect 11742 -20410 11776 -20394
rect 11742 -21002 11776 -20986
rect 12760 -20410 12794 -20394
rect 12760 -21002 12794 -20986
rect 13778 -20410 13812 -20394
rect 13778 -21002 13812 -20986
rect 14796 -20410 14830 -20394
rect 14796 -21002 14830 -20986
rect 15814 -20410 15848 -20394
rect 15814 -21002 15848 -20986
rect 16832 -20410 16866 -20394
rect 16832 -21002 16866 -20986
rect 17850 -20410 17884 -20394
rect 17850 -21002 17884 -20986
rect 18868 -20410 18902 -20394
rect 18868 -21002 18902 -20986
rect 19886 -20410 19920 -20394
rect 19886 -21002 19920 -20986
rect 20904 -20410 20938 -20394
rect 20904 -21002 20938 -20986
rect 21922 -20410 21956 -20394
rect 21922 -21002 21956 -20986
rect 22940 -20410 22974 -20394
rect 22940 -21002 22974 -20986
rect 5106 -21036 5166 -21032
rect 2812 -21070 2828 -21036
rect 3384 -21070 3400 -21036
rect 3830 -21070 3846 -21036
rect 4402 -21070 4418 -21036
rect 4848 -21070 4864 -21036
rect 5420 -21070 5436 -21036
rect 5866 -21070 5882 -21036
rect 6438 -21070 6454 -21036
rect 6884 -21070 6900 -21036
rect 7456 -21070 7472 -21036
rect 7902 -21070 7918 -21036
rect 8474 -21070 8490 -21036
rect 8920 -21070 8936 -21036
rect 9492 -21070 9508 -21036
rect 9938 -21070 9954 -21036
rect 10510 -21070 10526 -21036
rect 10956 -21070 10972 -21036
rect 11528 -21070 11544 -21036
rect 11974 -21070 11990 -21036
rect 12546 -21070 12562 -21036
rect 12992 -21070 13008 -21036
rect 13564 -21070 13580 -21036
rect 14010 -21070 14026 -21036
rect 14582 -21070 14598 -21036
rect 15028 -21070 15044 -21036
rect 15600 -21070 15616 -21036
rect 16046 -21070 16062 -21036
rect 16618 -21070 16634 -21036
rect 17064 -21070 17080 -21036
rect 17636 -21070 17652 -21036
rect 18082 -21070 18098 -21036
rect 18654 -21070 18670 -21036
rect 19100 -21070 19116 -21036
rect 19672 -21070 19688 -21036
rect 20118 -21070 20134 -21036
rect 20690 -21070 20706 -21036
rect 21136 -21070 21152 -21036
rect 21708 -21070 21724 -21036
rect 22154 -21070 22170 -21036
rect 22726 -21070 22742 -21036
rect -10004 -21096 -9922 -21072
rect -10004 -21130 -9980 -21096
rect -9946 -21130 -9922 -21096
rect -10004 -21154 -9922 -21130
rect -8986 -21096 -8904 -21072
rect -8986 -21130 -8962 -21096
rect -8928 -21130 -8904 -21096
rect -8986 -21154 -8904 -21130
rect -7968 -21096 -7886 -21072
rect -7968 -21130 -7944 -21096
rect -7910 -21130 -7886 -21096
rect -7968 -21154 -7886 -21130
rect -6950 -21096 -6868 -21072
rect -6950 -21130 -6926 -21096
rect -6892 -21130 -6868 -21096
rect -6950 -21154 -6868 -21130
rect -5932 -21096 -5850 -21072
rect -5932 -21130 -5908 -21096
rect -5874 -21130 -5850 -21096
rect -5932 -21154 -5850 -21130
rect -4914 -21096 -4832 -21072
rect -4914 -21130 -4890 -21096
rect -4856 -21130 -4832 -21096
rect -4914 -21154 -4832 -21130
rect -3896 -21096 -3814 -21072
rect -3896 -21130 -3872 -21096
rect -3838 -21130 -3814 -21096
rect -3896 -21154 -3814 -21130
rect -2878 -21096 -2796 -21072
rect -2878 -21130 -2854 -21096
rect -2820 -21130 -2796 -21096
rect -2878 -21154 -2796 -21130
rect -1860 -21096 -1778 -21072
rect -1860 -21130 -1836 -21096
rect -1802 -21130 -1778 -21096
rect -1860 -21154 -1778 -21130
rect -842 -21096 -760 -21072
rect -842 -21130 -818 -21096
rect -784 -21130 -760 -21096
rect -842 -21154 -760 -21130
rect 176 -21096 258 -21072
rect 176 -21130 200 -21096
rect 234 -21130 258 -21096
rect 176 -21154 258 -21130
rect 3062 -21296 3144 -21272
rect -10276 -21336 -10260 -21302
rect -9704 -21336 -9688 -21302
rect -9258 -21336 -9242 -21302
rect -8686 -21336 -8670 -21302
rect -8240 -21336 -8224 -21302
rect -7668 -21336 -7652 -21302
rect -7222 -21336 -7206 -21302
rect -6650 -21336 -6634 -21302
rect -6204 -21336 -6188 -21302
rect -5632 -21336 -5616 -21302
rect -5186 -21336 -5170 -21302
rect -4614 -21336 -4598 -21302
rect -4168 -21336 -4152 -21302
rect -3596 -21336 -3580 -21302
rect -3150 -21336 -3134 -21302
rect -2578 -21336 -2562 -21302
rect -2132 -21336 -2116 -21302
rect -1560 -21336 -1544 -21302
rect -1114 -21336 -1098 -21302
rect -542 -21336 -526 -21302
rect -96 -21336 -80 -21302
rect 476 -21336 492 -21302
rect 3062 -21330 3086 -21296
rect 3120 -21330 3144 -21296
rect 3062 -21354 3144 -21330
rect 4080 -21296 4162 -21272
rect 4080 -21330 4104 -21296
rect 4138 -21330 4162 -21296
rect 4080 -21354 4162 -21330
rect 5098 -21296 5180 -21272
rect 5098 -21330 5122 -21296
rect 5156 -21330 5180 -21296
rect 5098 -21354 5180 -21330
rect 6116 -21296 6198 -21272
rect 6116 -21330 6140 -21296
rect 6174 -21330 6198 -21296
rect 6116 -21354 6198 -21330
rect 7134 -21296 7216 -21272
rect 7134 -21330 7158 -21296
rect 7192 -21330 7216 -21296
rect 7134 -21354 7216 -21330
rect 8152 -21296 8234 -21272
rect 8152 -21330 8176 -21296
rect 8210 -21330 8234 -21296
rect 8152 -21354 8234 -21330
rect 9170 -21296 9252 -21272
rect 9170 -21330 9194 -21296
rect 9228 -21330 9252 -21296
rect 9170 -21354 9252 -21330
rect 10188 -21296 10270 -21272
rect 10188 -21330 10212 -21296
rect 10246 -21330 10270 -21296
rect 10188 -21354 10270 -21330
rect 11206 -21296 11288 -21272
rect 11206 -21330 11230 -21296
rect 11264 -21330 11288 -21296
rect 11206 -21354 11288 -21330
rect 12224 -21296 12306 -21272
rect 12224 -21330 12248 -21296
rect 12282 -21330 12306 -21296
rect 12224 -21354 12306 -21330
rect 13242 -21296 13324 -21272
rect 13242 -21330 13266 -21296
rect 13300 -21330 13324 -21296
rect 13242 -21354 13324 -21330
rect 14260 -21296 14342 -21272
rect 14260 -21330 14284 -21296
rect 14318 -21330 14342 -21296
rect 14260 -21354 14342 -21330
rect 15278 -21296 15360 -21272
rect 15278 -21330 15302 -21296
rect 15336 -21330 15360 -21296
rect 15278 -21354 15360 -21330
rect 16296 -21296 16378 -21272
rect 16296 -21330 16320 -21296
rect 16354 -21330 16378 -21296
rect 16296 -21354 16378 -21330
rect 17314 -21296 17396 -21272
rect 17314 -21330 17338 -21296
rect 17372 -21330 17396 -21296
rect 17314 -21354 17396 -21330
rect 18332 -21296 18414 -21272
rect 18332 -21330 18356 -21296
rect 18390 -21330 18414 -21296
rect 18332 -21354 18414 -21330
rect 19350 -21296 19432 -21272
rect 19350 -21330 19374 -21296
rect 19408 -21330 19432 -21296
rect 19350 -21354 19432 -21330
rect 20368 -21296 20450 -21272
rect 20368 -21330 20392 -21296
rect 20426 -21330 20450 -21296
rect 20368 -21354 20450 -21330
rect 21386 -21296 21468 -21272
rect 21386 -21330 21410 -21296
rect 21444 -21330 21468 -21296
rect 21386 -21354 21468 -21330
rect 22404 -21296 22486 -21272
rect 22404 -21330 22428 -21296
rect 22462 -21330 22486 -21296
rect 22404 -21354 22486 -21330
rect -10508 -21386 -10474 -21370
rect -10508 -21978 -10474 -21962
rect -9490 -21386 -9456 -21370
rect -9490 -21978 -9456 -21962
rect -8472 -21386 -8438 -21370
rect -8472 -21978 -8438 -21962
rect -7454 -21386 -7420 -21370
rect -7454 -21978 -7420 -21962
rect -6436 -21386 -6402 -21370
rect -6436 -21978 -6402 -21962
rect -5418 -21386 -5384 -21370
rect -5418 -21978 -5384 -21962
rect -4400 -21386 -4366 -21370
rect -4400 -21978 -4366 -21962
rect -3382 -21386 -3348 -21370
rect -3382 -21978 -3348 -21962
rect -2364 -21386 -2330 -21370
rect -2364 -21978 -2330 -21962
rect -1346 -21386 -1312 -21370
rect -1346 -21978 -1312 -21962
rect -328 -21386 -294 -21370
rect -328 -21978 -294 -21962
rect 690 -21386 724 -21370
rect 2812 -21594 2828 -21560
rect 3384 -21594 3400 -21560
rect 3830 -21594 3846 -21560
rect 4402 -21594 4418 -21560
rect 4848 -21594 4864 -21560
rect 5420 -21594 5436 -21560
rect 5866 -21594 5882 -21560
rect 6438 -21594 6454 -21560
rect 6884 -21594 6900 -21560
rect 7456 -21594 7472 -21560
rect 7902 -21594 7918 -21560
rect 8474 -21594 8490 -21560
rect 8920 -21594 8936 -21560
rect 9492 -21594 9508 -21560
rect 9938 -21594 9954 -21560
rect 10510 -21594 10526 -21560
rect 10956 -21594 10972 -21560
rect 11528 -21594 11544 -21560
rect 11974 -21594 11990 -21560
rect 12546 -21594 12562 -21560
rect 12992 -21594 13008 -21560
rect 13564 -21594 13580 -21560
rect 14010 -21594 14026 -21560
rect 14582 -21594 14598 -21560
rect 15028 -21594 15044 -21560
rect 15600 -21594 15616 -21560
rect 16046 -21594 16062 -21560
rect 16618 -21594 16634 -21560
rect 17064 -21594 17080 -21560
rect 17636 -21594 17652 -21560
rect 18082 -21594 18098 -21560
rect 18654 -21594 18670 -21560
rect 19100 -21594 19116 -21560
rect 19672 -21594 19688 -21560
rect 20118 -21594 20134 -21560
rect 20690 -21594 20706 -21560
rect 21136 -21594 21152 -21560
rect 21708 -21594 21724 -21560
rect 22154 -21594 22170 -21560
rect 22726 -21594 22742 -21560
rect 690 -21978 724 -21962
rect 2580 -21644 2614 -21628
rect -10276 -22046 -10260 -22012
rect -9704 -22046 -9688 -22012
rect -9258 -22046 -9242 -22012
rect -8686 -22046 -8670 -22012
rect -8240 -22046 -8224 -22012
rect -7668 -22046 -7652 -22012
rect -7222 -22046 -7206 -22012
rect -6650 -22046 -6634 -22012
rect -6204 -22046 -6188 -22012
rect -5632 -22046 -5616 -22012
rect -5186 -22046 -5170 -22012
rect -4614 -22046 -4598 -22012
rect -4168 -22046 -4152 -22012
rect -3596 -22046 -3580 -22012
rect -3150 -22046 -3134 -22012
rect -2578 -22046 -2562 -22012
rect -2132 -22046 -2116 -22012
rect -1560 -22046 -1544 -22012
rect -1114 -22046 -1098 -22012
rect -542 -22046 -526 -22012
rect -96 -22046 -80 -22012
rect 476 -22046 492 -22012
rect -10026 -22204 -9944 -22180
rect -10026 -22238 -10002 -22204
rect -9968 -22238 -9944 -22204
rect -10026 -22262 -9944 -22238
rect -9008 -22204 -8926 -22180
rect -9008 -22238 -8984 -22204
rect -8950 -22238 -8926 -22204
rect -9008 -22262 -8926 -22238
rect -7990 -22204 -7908 -22180
rect -7990 -22238 -7966 -22204
rect -7932 -22238 -7908 -22204
rect -7990 -22262 -7908 -22238
rect -6972 -22204 -6890 -22180
rect -6972 -22238 -6948 -22204
rect -6914 -22238 -6890 -22204
rect -6972 -22262 -6890 -22238
rect -5954 -22204 -5872 -22180
rect -5954 -22238 -5930 -22204
rect -5896 -22238 -5872 -22204
rect -5954 -22262 -5872 -22238
rect -4936 -22204 -4854 -22180
rect -4936 -22238 -4912 -22204
rect -4878 -22238 -4854 -22204
rect -4936 -22262 -4854 -22238
rect -3918 -22204 -3836 -22180
rect -3918 -22238 -3894 -22204
rect -3860 -22238 -3836 -22204
rect -3918 -22262 -3836 -22238
rect -2900 -22204 -2818 -22180
rect -2900 -22238 -2876 -22204
rect -2842 -22238 -2818 -22204
rect -2900 -22262 -2818 -22238
rect -1882 -22204 -1800 -22180
rect -1882 -22238 -1858 -22204
rect -1824 -22238 -1800 -22204
rect -1882 -22262 -1800 -22238
rect -864 -22204 -782 -22180
rect -864 -22238 -840 -22204
rect -806 -22238 -782 -22204
rect -864 -22262 -782 -22238
rect 154 -22204 236 -22180
rect 154 -22238 178 -22204
rect 212 -22238 236 -22204
rect 2580 -22236 2614 -22220
rect 3598 -21644 3632 -21628
rect 3598 -22236 3632 -22220
rect 4616 -21644 4650 -21628
rect 4616 -22236 4650 -22220
rect 5634 -21644 5668 -21628
rect 5634 -22236 5668 -22220
rect 6652 -21644 6686 -21628
rect 6652 -22236 6686 -22220
rect 7670 -21644 7704 -21628
rect 7670 -22236 7704 -22220
rect 8688 -21644 8722 -21628
rect 8688 -22236 8722 -22220
rect 9706 -21644 9740 -21628
rect 9706 -22236 9740 -22220
rect 10724 -21644 10758 -21628
rect 10724 -22236 10758 -22220
rect 11742 -21644 11776 -21628
rect 11742 -22236 11776 -22220
rect 12760 -21644 12794 -21628
rect 12760 -22236 12794 -22220
rect 13778 -21644 13812 -21628
rect 13778 -22236 13812 -22220
rect 14796 -21644 14830 -21628
rect 14796 -22236 14830 -22220
rect 15814 -21644 15848 -21628
rect 15814 -22236 15848 -22220
rect 16832 -21644 16866 -21628
rect 16832 -22236 16866 -22220
rect 17850 -21644 17884 -21628
rect 17850 -22236 17884 -22220
rect 18868 -21644 18902 -21628
rect 18868 -22236 18902 -22220
rect 19886 -21644 19920 -21628
rect 19886 -22236 19920 -22220
rect 20904 -21644 20938 -21628
rect 20904 -22236 20938 -22220
rect 21922 -21644 21956 -21628
rect 21922 -22236 21956 -22220
rect 22940 -21644 22974 -21628
rect 22940 -22236 22974 -22220
rect 154 -22262 236 -22238
rect 11230 -22270 11290 -22268
rect 13274 -22270 13334 -22266
rect 16312 -22270 16372 -22266
rect 2812 -22304 2828 -22270
rect 3384 -22304 3400 -22270
rect 3830 -22304 3846 -22270
rect 4402 -22304 4418 -22270
rect 4848 -22304 4864 -22270
rect 5420 -22304 5436 -22270
rect 5866 -22304 5882 -22270
rect 6438 -22304 6454 -22270
rect 6884 -22304 6900 -22270
rect 7456 -22304 7472 -22270
rect 7902 -22304 7918 -22270
rect 8474 -22304 8490 -22270
rect 8920 -22304 8936 -22270
rect 9492 -22304 9508 -22270
rect 9938 -22304 9954 -22270
rect 10510 -22304 10526 -22270
rect 10956 -22304 10972 -22270
rect 11528 -22304 11544 -22270
rect 11974 -22304 11990 -22270
rect 12546 -22304 12562 -22270
rect 12992 -22304 13008 -22270
rect 13564 -22304 13580 -22270
rect 14010 -22304 14026 -22270
rect 14582 -22304 14598 -22270
rect 15028 -22304 15044 -22270
rect 15600 -22304 15616 -22270
rect 16046 -22304 16062 -22270
rect 16618 -22304 16634 -22270
rect 17064 -22304 17080 -22270
rect 17636 -22304 17652 -22270
rect 18082 -22304 18098 -22270
rect 18654 -22304 18670 -22270
rect 19100 -22304 19116 -22270
rect 19672 -22304 19688 -22270
rect 20118 -22304 20134 -22270
rect 20690 -22304 20706 -22270
rect 21136 -22304 21152 -22270
rect 21708 -22304 21724 -22270
rect 22154 -22304 22170 -22270
rect 22726 -22304 22742 -22270
rect -10276 -22448 -10260 -22414
rect -9704 -22448 -9688 -22414
rect -9258 -22448 -9242 -22414
rect -8686 -22448 -8670 -22414
rect -8240 -22448 -8224 -22414
rect -7668 -22448 -7652 -22414
rect -7222 -22448 -7206 -22414
rect -6650 -22448 -6634 -22414
rect -6204 -22448 -6188 -22414
rect -5632 -22448 -5616 -22414
rect -5186 -22448 -5170 -22414
rect -4614 -22448 -4598 -22414
rect -4168 -22448 -4152 -22414
rect -3596 -22448 -3580 -22414
rect -3150 -22448 -3134 -22414
rect -2578 -22448 -2562 -22414
rect -2132 -22448 -2116 -22414
rect -1560 -22448 -1544 -22414
rect -1114 -22448 -1098 -22414
rect -542 -22448 -526 -22414
rect -96 -22448 -80 -22414
rect 476 -22448 492 -22414
rect -10508 -22498 -10474 -22482
rect -10508 -23090 -10474 -23074
rect -9490 -22498 -9456 -22482
rect -9490 -23090 -9456 -23074
rect -8472 -22498 -8438 -22482
rect -8472 -23090 -8438 -23074
rect -7454 -22498 -7420 -22482
rect -7454 -23090 -7420 -23074
rect -6436 -22498 -6402 -22482
rect -6436 -23090 -6402 -23074
rect -5418 -22498 -5384 -22482
rect -5418 -23090 -5384 -23074
rect -4400 -22498 -4366 -22482
rect -4400 -23090 -4366 -23074
rect -3382 -22498 -3348 -22482
rect -3382 -23090 -3348 -23074
rect -2364 -22498 -2330 -22482
rect -2364 -23090 -2330 -23074
rect -1346 -22498 -1312 -22482
rect -1346 -23090 -1312 -23074
rect -328 -22498 -294 -22482
rect -328 -23090 -294 -23074
rect 690 -22498 724 -22482
rect 3074 -22520 3156 -22496
rect 3074 -22554 3098 -22520
rect 3132 -22554 3156 -22520
rect 3074 -22578 3156 -22554
rect 4092 -22520 4174 -22496
rect 4092 -22554 4116 -22520
rect 4150 -22554 4174 -22520
rect 4092 -22578 4174 -22554
rect 5110 -22520 5192 -22496
rect 5110 -22554 5134 -22520
rect 5168 -22554 5192 -22520
rect 5110 -22578 5192 -22554
rect 6128 -22520 6210 -22496
rect 6128 -22554 6152 -22520
rect 6186 -22554 6210 -22520
rect 6128 -22578 6210 -22554
rect 7146 -22520 7228 -22496
rect 7146 -22554 7170 -22520
rect 7204 -22554 7228 -22520
rect 7146 -22578 7228 -22554
rect 8164 -22520 8246 -22496
rect 8164 -22554 8188 -22520
rect 8222 -22554 8246 -22520
rect 8164 -22578 8246 -22554
rect 9182 -22520 9264 -22496
rect 9182 -22554 9206 -22520
rect 9240 -22554 9264 -22520
rect 9182 -22578 9264 -22554
rect 10200 -22520 10282 -22496
rect 10200 -22554 10224 -22520
rect 10258 -22554 10282 -22520
rect 10200 -22578 10282 -22554
rect 11218 -22520 11300 -22496
rect 11218 -22554 11242 -22520
rect 11276 -22554 11300 -22520
rect 11218 -22578 11300 -22554
rect 12236 -22520 12318 -22496
rect 12236 -22554 12260 -22520
rect 12294 -22554 12318 -22520
rect 12236 -22578 12318 -22554
rect 13254 -22520 13336 -22496
rect 13254 -22554 13278 -22520
rect 13312 -22554 13336 -22520
rect 13254 -22578 13336 -22554
rect 14272 -22520 14354 -22496
rect 14272 -22554 14296 -22520
rect 14330 -22554 14354 -22520
rect 14272 -22578 14354 -22554
rect 15290 -22520 15372 -22496
rect 15290 -22554 15314 -22520
rect 15348 -22554 15372 -22520
rect 15290 -22578 15372 -22554
rect 16308 -22520 16390 -22496
rect 16308 -22554 16332 -22520
rect 16366 -22554 16390 -22520
rect 16308 -22578 16390 -22554
rect 17326 -22520 17408 -22496
rect 17326 -22554 17350 -22520
rect 17384 -22554 17408 -22520
rect 17326 -22578 17408 -22554
rect 18344 -22520 18426 -22496
rect 18344 -22554 18368 -22520
rect 18402 -22554 18426 -22520
rect 18344 -22578 18426 -22554
rect 19362 -22520 19444 -22496
rect 19362 -22554 19386 -22520
rect 19420 -22554 19444 -22520
rect 19362 -22578 19444 -22554
rect 20380 -22520 20462 -22496
rect 20380 -22554 20404 -22520
rect 20438 -22554 20462 -22520
rect 20380 -22578 20462 -22554
rect 21398 -22520 21480 -22496
rect 21398 -22554 21422 -22520
rect 21456 -22554 21480 -22520
rect 21398 -22578 21480 -22554
rect 22416 -22520 22498 -22496
rect 22416 -22554 22440 -22520
rect 22474 -22554 22498 -22520
rect 22416 -22578 22498 -22554
rect 2812 -22826 2828 -22792
rect 3384 -22826 3400 -22792
rect 3830 -22826 3846 -22792
rect 4402 -22826 4418 -22792
rect 4848 -22826 4864 -22792
rect 5420 -22826 5436 -22792
rect 5866 -22826 5882 -22792
rect 6438 -22826 6454 -22792
rect 6884 -22826 6900 -22792
rect 7456 -22826 7472 -22792
rect 7902 -22826 7918 -22792
rect 8474 -22826 8490 -22792
rect 8920 -22826 8936 -22792
rect 9492 -22826 9508 -22792
rect 9938 -22826 9954 -22792
rect 10510 -22826 10526 -22792
rect 10956 -22826 10972 -22792
rect 11528 -22826 11544 -22792
rect 11974 -22826 11990 -22792
rect 12546 -22826 12562 -22792
rect 12992 -22826 13008 -22792
rect 13564 -22826 13580 -22792
rect 14010 -22826 14026 -22792
rect 14582 -22826 14598 -22792
rect 15028 -22826 15044 -22792
rect 15600 -22826 15616 -22792
rect 16046 -22826 16062 -22792
rect 16618 -22826 16634 -22792
rect 17064 -22826 17080 -22792
rect 17636 -22826 17652 -22792
rect 18082 -22826 18098 -22792
rect 18654 -22826 18670 -22792
rect 19100 -22826 19116 -22792
rect 19672 -22826 19688 -22792
rect 20118 -22826 20134 -22792
rect 20690 -22826 20706 -22792
rect 21136 -22826 21152 -22792
rect 21708 -22826 21724 -22792
rect 22154 -22826 22170 -22792
rect 22726 -22826 22742 -22792
rect 6134 -22828 6194 -22826
rect 690 -23090 724 -23074
rect 2580 -22876 2614 -22860
rect -10276 -23158 -10260 -23124
rect -9704 -23158 -9688 -23124
rect -9258 -23158 -9242 -23124
rect -8686 -23158 -8670 -23124
rect -8240 -23158 -8224 -23124
rect -7668 -23158 -7652 -23124
rect -7222 -23158 -7206 -23124
rect -6650 -23158 -6634 -23124
rect -6204 -23158 -6188 -23124
rect -5632 -23158 -5616 -23124
rect -5186 -23158 -5170 -23124
rect -4614 -23158 -4598 -23124
rect -4168 -23158 -4152 -23124
rect -3596 -23158 -3580 -23124
rect -3150 -23158 -3134 -23124
rect -2578 -23158 -2562 -23124
rect -2132 -23158 -2116 -23124
rect -1560 -23158 -1544 -23124
rect -1114 -23158 -1098 -23124
rect -542 -23158 -526 -23124
rect -96 -23158 -80 -23124
rect 476 -23158 492 -23124
rect -10026 -23310 -9944 -23286
rect -10026 -23344 -10002 -23310
rect -9968 -23344 -9944 -23310
rect -10026 -23368 -9944 -23344
rect -9008 -23310 -8926 -23286
rect -9008 -23344 -8984 -23310
rect -8950 -23344 -8926 -23310
rect -9008 -23368 -8926 -23344
rect -7990 -23310 -7908 -23286
rect -7990 -23344 -7966 -23310
rect -7932 -23344 -7908 -23310
rect -7990 -23368 -7908 -23344
rect -6972 -23310 -6890 -23286
rect -6972 -23344 -6948 -23310
rect -6914 -23344 -6890 -23310
rect -6972 -23368 -6890 -23344
rect -5954 -23310 -5872 -23286
rect -5954 -23344 -5930 -23310
rect -5896 -23344 -5872 -23310
rect -5954 -23368 -5872 -23344
rect -4936 -23310 -4854 -23286
rect -4936 -23344 -4912 -23310
rect -4878 -23344 -4854 -23310
rect -4936 -23368 -4854 -23344
rect -3918 -23310 -3836 -23286
rect -3918 -23344 -3894 -23310
rect -3860 -23344 -3836 -23310
rect -3918 -23368 -3836 -23344
rect -2900 -23310 -2818 -23286
rect -2900 -23344 -2876 -23310
rect -2842 -23344 -2818 -23310
rect -2900 -23368 -2818 -23344
rect -1882 -23310 -1800 -23286
rect -1882 -23344 -1858 -23310
rect -1824 -23344 -1800 -23310
rect -1882 -23368 -1800 -23344
rect -864 -23310 -782 -23286
rect -864 -23344 -840 -23310
rect -806 -23344 -782 -23310
rect -864 -23368 -782 -23344
rect 154 -23310 236 -23286
rect 154 -23344 178 -23310
rect 212 -23344 236 -23310
rect 154 -23368 236 -23344
rect 2580 -23468 2614 -23452
rect 3598 -22876 3632 -22860
rect 3598 -23468 3632 -23452
rect 4616 -22876 4650 -22860
rect 4616 -23468 4650 -23452
rect 5634 -22876 5668 -22860
rect 5634 -23468 5668 -23452
rect 6652 -22876 6686 -22860
rect 6652 -23468 6686 -23452
rect 7670 -22876 7704 -22860
rect 7670 -23468 7704 -23452
rect 8688 -22876 8722 -22860
rect 8688 -23468 8722 -23452
rect 9706 -22876 9740 -22860
rect 9706 -23468 9740 -23452
rect 10724 -22876 10758 -22860
rect 10724 -23468 10758 -23452
rect 11742 -22876 11776 -22860
rect 11742 -23468 11776 -23452
rect 12760 -22876 12794 -22860
rect 12760 -23468 12794 -23452
rect 13778 -22876 13812 -22860
rect 13778 -23468 13812 -23452
rect 14796 -22876 14830 -22860
rect 14796 -23468 14830 -23452
rect 15814 -22876 15848 -22860
rect 15814 -23468 15848 -23452
rect 16832 -22876 16866 -22860
rect 16832 -23468 16866 -23452
rect 17850 -22876 17884 -22860
rect 17850 -23468 17884 -23452
rect 18868 -22876 18902 -22860
rect 18868 -23468 18902 -23452
rect 19886 -22876 19920 -22860
rect 19886 -23468 19920 -23452
rect 20904 -22876 20938 -22860
rect 20904 -23468 20938 -23452
rect 21922 -22876 21956 -22860
rect 21922 -23468 21956 -23452
rect 22940 -22876 22974 -22860
rect 22940 -23468 22974 -23452
rect 10206 -23502 10266 -23492
rect -10276 -23560 -10260 -23526
rect -9704 -23560 -9688 -23526
rect -9258 -23560 -9242 -23526
rect -8686 -23560 -8670 -23526
rect -8240 -23560 -8224 -23526
rect -7668 -23560 -7652 -23526
rect -7222 -23560 -7206 -23526
rect -6650 -23560 -6634 -23526
rect -6204 -23560 -6188 -23526
rect -5632 -23560 -5616 -23526
rect -5186 -23560 -5170 -23526
rect -4614 -23560 -4598 -23526
rect -4168 -23560 -4152 -23526
rect -3596 -23560 -3580 -23526
rect -3150 -23560 -3134 -23526
rect -2578 -23560 -2562 -23526
rect -2132 -23560 -2116 -23526
rect -1560 -23560 -1544 -23526
rect -1114 -23560 -1098 -23526
rect -542 -23560 -526 -23526
rect -96 -23560 -80 -23526
rect 476 -23560 492 -23526
rect 2812 -23536 2828 -23502
rect 3384 -23536 3400 -23502
rect 3830 -23536 3846 -23502
rect 4402 -23536 4418 -23502
rect 4848 -23536 4864 -23502
rect 5420 -23536 5436 -23502
rect 5866 -23536 5882 -23502
rect 6438 -23536 6454 -23502
rect 6884 -23536 6900 -23502
rect 7456 -23536 7472 -23502
rect 7902 -23536 7918 -23502
rect 8474 -23536 8490 -23502
rect 8920 -23536 8936 -23502
rect 9492 -23536 9508 -23502
rect 9938 -23536 9954 -23502
rect 10510 -23536 10526 -23502
rect 10956 -23536 10972 -23502
rect 11528 -23536 11544 -23502
rect 11974 -23536 11990 -23502
rect 12546 -23536 12562 -23502
rect 12992 -23536 13008 -23502
rect 13564 -23536 13580 -23502
rect 14010 -23536 14026 -23502
rect 14582 -23536 14598 -23502
rect 15028 -23536 15044 -23502
rect 15600 -23536 15616 -23502
rect 16046 -23536 16062 -23502
rect 16618 -23536 16634 -23502
rect 17064 -23536 17080 -23502
rect 17636 -23536 17652 -23502
rect 18082 -23536 18098 -23502
rect 18654 -23536 18670 -23502
rect 19100 -23536 19116 -23502
rect 19672 -23536 19688 -23502
rect 20118 -23536 20134 -23502
rect 20690 -23536 20706 -23502
rect 21136 -23536 21152 -23502
rect 21708 -23536 21724 -23502
rect 22154 -23536 22170 -23502
rect 22726 -23536 22742 -23502
rect -10508 -23610 -10474 -23594
rect -10508 -24202 -10474 -24186
rect -9490 -23610 -9456 -23594
rect -9490 -24202 -9456 -24186
rect -8472 -23610 -8438 -23594
rect -8472 -24202 -8438 -24186
rect -7454 -23610 -7420 -23594
rect -7454 -24202 -7420 -24186
rect -6436 -23610 -6402 -23594
rect -6436 -24202 -6402 -24186
rect -5418 -23610 -5384 -23594
rect -5418 -24202 -5384 -24186
rect -4400 -23610 -4366 -23594
rect -4400 -24202 -4366 -24186
rect -3382 -23610 -3348 -23594
rect -3382 -24202 -3348 -24186
rect -2364 -23610 -2330 -23594
rect -2364 -24202 -2330 -24186
rect -1346 -23610 -1312 -23594
rect -1346 -24202 -1312 -24186
rect -328 -23610 -294 -23594
rect -328 -24202 -294 -24186
rect 690 -23610 724 -23594
rect 3074 -23756 3156 -23732
rect 3074 -23790 3098 -23756
rect 3132 -23790 3156 -23756
rect 3074 -23814 3156 -23790
rect 4092 -23756 4174 -23732
rect 4092 -23790 4116 -23756
rect 4150 -23790 4174 -23756
rect 4092 -23814 4174 -23790
rect 5110 -23756 5192 -23732
rect 5110 -23790 5134 -23756
rect 5168 -23790 5192 -23756
rect 5110 -23814 5192 -23790
rect 6128 -23756 6210 -23732
rect 6128 -23790 6152 -23756
rect 6186 -23790 6210 -23756
rect 6128 -23814 6210 -23790
rect 7146 -23756 7228 -23732
rect 7146 -23790 7170 -23756
rect 7204 -23790 7228 -23756
rect 7146 -23814 7228 -23790
rect 8164 -23756 8246 -23732
rect 8164 -23790 8188 -23756
rect 8222 -23790 8246 -23756
rect 8164 -23814 8246 -23790
rect 9182 -23756 9264 -23732
rect 9182 -23790 9206 -23756
rect 9240 -23790 9264 -23756
rect 9182 -23814 9264 -23790
rect 10200 -23756 10282 -23732
rect 10200 -23790 10224 -23756
rect 10258 -23790 10282 -23756
rect 10200 -23814 10282 -23790
rect 11218 -23756 11300 -23732
rect 11218 -23790 11242 -23756
rect 11276 -23790 11300 -23756
rect 11218 -23814 11300 -23790
rect 12236 -23756 12318 -23732
rect 12236 -23790 12260 -23756
rect 12294 -23790 12318 -23756
rect 12236 -23814 12318 -23790
rect 13254 -23756 13336 -23732
rect 13254 -23790 13278 -23756
rect 13312 -23790 13336 -23756
rect 13254 -23814 13336 -23790
rect 14272 -23756 14354 -23732
rect 14272 -23790 14296 -23756
rect 14330 -23790 14354 -23756
rect 14272 -23814 14354 -23790
rect 15290 -23756 15372 -23732
rect 15290 -23790 15314 -23756
rect 15348 -23790 15372 -23756
rect 15290 -23814 15372 -23790
rect 16308 -23756 16390 -23732
rect 16308 -23790 16332 -23756
rect 16366 -23790 16390 -23756
rect 16308 -23814 16390 -23790
rect 17326 -23756 17408 -23732
rect 17326 -23790 17350 -23756
rect 17384 -23790 17408 -23756
rect 17326 -23814 17408 -23790
rect 18344 -23756 18426 -23732
rect 18344 -23790 18368 -23756
rect 18402 -23790 18426 -23756
rect 18344 -23814 18426 -23790
rect 19362 -23756 19444 -23732
rect 19362 -23790 19386 -23756
rect 19420 -23790 19444 -23756
rect 19362 -23814 19444 -23790
rect 20380 -23756 20462 -23732
rect 20380 -23790 20404 -23756
rect 20438 -23790 20462 -23756
rect 20380 -23814 20462 -23790
rect 21398 -23756 21480 -23732
rect 21398 -23790 21422 -23756
rect 21456 -23790 21480 -23756
rect 21398 -23814 21480 -23790
rect 22416 -23756 22498 -23732
rect 22416 -23790 22440 -23756
rect 22474 -23790 22498 -23756
rect 22416 -23814 22498 -23790
rect 2812 -24060 2828 -24026
rect 3384 -24060 3400 -24026
rect 3830 -24060 3846 -24026
rect 4402 -24060 4418 -24026
rect 4848 -24060 4864 -24026
rect 5420 -24060 5436 -24026
rect 5866 -24060 5882 -24026
rect 6438 -24060 6454 -24026
rect 6884 -24060 6900 -24026
rect 7456 -24060 7472 -24026
rect 7902 -24060 7918 -24026
rect 8474 -24060 8490 -24026
rect 8920 -24060 8936 -24026
rect 9492 -24060 9508 -24026
rect 9938 -24060 9954 -24026
rect 10510 -24060 10526 -24026
rect 10956 -24060 10972 -24026
rect 11528 -24060 11544 -24026
rect 11974 -24060 11990 -24026
rect 12546 -24060 12562 -24026
rect 12992 -24060 13008 -24026
rect 13564 -24060 13580 -24026
rect 14010 -24060 14026 -24026
rect 14582 -24060 14598 -24026
rect 15028 -24060 15044 -24026
rect 15600 -24060 15616 -24026
rect 16046 -24060 16062 -24026
rect 16618 -24060 16634 -24026
rect 17064 -24060 17080 -24026
rect 17636 -24060 17652 -24026
rect 18082 -24060 18098 -24026
rect 18654 -24060 18670 -24026
rect 19100 -24060 19116 -24026
rect 19672 -24060 19688 -24026
rect 20118 -24060 20134 -24026
rect 20690 -24060 20706 -24026
rect 21136 -24060 21152 -24026
rect 21708 -24060 21724 -24026
rect 22154 -24060 22170 -24026
rect 22726 -24060 22742 -24026
rect 6120 -24062 6180 -24060
rect 690 -24202 724 -24186
rect 2580 -24110 2614 -24094
rect -10276 -24270 -10260 -24236
rect -9704 -24270 -9688 -24236
rect -9258 -24270 -9242 -24236
rect -8686 -24270 -8670 -24236
rect -8240 -24270 -8224 -24236
rect -7668 -24270 -7652 -24236
rect -7222 -24270 -7206 -24236
rect -6650 -24270 -6634 -24236
rect -6204 -24270 -6188 -24236
rect -5632 -24270 -5616 -24236
rect -5186 -24270 -5170 -24236
rect -4614 -24270 -4598 -24236
rect -4168 -24270 -4152 -24236
rect -3596 -24270 -3580 -24236
rect -3150 -24270 -3134 -24236
rect -2578 -24270 -2562 -24236
rect -2132 -24270 -2116 -24236
rect -1560 -24270 -1544 -24236
rect -1114 -24270 -1098 -24236
rect -542 -24270 -526 -24236
rect -96 -24270 -80 -24236
rect 476 -24270 492 -24236
rect -10026 -24652 -9944 -24628
rect -10026 -24686 -10002 -24652
rect -9968 -24686 -9944 -24652
rect -10026 -24710 -9944 -24686
rect -9008 -24652 -8926 -24628
rect -9008 -24686 -8984 -24652
rect -8950 -24686 -8926 -24652
rect -9008 -24710 -8926 -24686
rect -7990 -24652 -7908 -24628
rect -7990 -24686 -7966 -24652
rect -7932 -24686 -7908 -24652
rect -7990 -24710 -7908 -24686
rect -6972 -24652 -6890 -24628
rect -6972 -24686 -6948 -24652
rect -6914 -24686 -6890 -24652
rect -6972 -24710 -6890 -24686
rect -5954 -24652 -5872 -24628
rect -5954 -24686 -5930 -24652
rect -5896 -24686 -5872 -24652
rect -5954 -24710 -5872 -24686
rect -4936 -24652 -4854 -24628
rect -4936 -24686 -4912 -24652
rect -4878 -24686 -4854 -24652
rect -4936 -24710 -4854 -24686
rect -3918 -24652 -3836 -24628
rect -3918 -24686 -3894 -24652
rect -3860 -24686 -3836 -24652
rect -3918 -24710 -3836 -24686
rect -2900 -24652 -2818 -24628
rect -2900 -24686 -2876 -24652
rect -2842 -24686 -2818 -24652
rect -2900 -24710 -2818 -24686
rect -1882 -24652 -1800 -24628
rect -1882 -24686 -1858 -24652
rect -1824 -24686 -1800 -24652
rect -1882 -24710 -1800 -24686
rect -864 -24652 -782 -24628
rect -864 -24686 -840 -24652
rect -806 -24686 -782 -24652
rect -864 -24710 -782 -24686
rect 154 -24652 236 -24628
rect 154 -24686 178 -24652
rect 212 -24686 236 -24652
rect 154 -24710 236 -24686
rect 2580 -24702 2614 -24686
rect 3598 -24110 3632 -24094
rect 3598 -24702 3632 -24686
rect 4616 -24110 4650 -24094
rect 4616 -24702 4650 -24686
rect 5634 -24110 5668 -24094
rect 5634 -24702 5668 -24686
rect 6652 -24110 6686 -24094
rect 6652 -24702 6686 -24686
rect 7670 -24110 7704 -24094
rect 7670 -24702 7704 -24686
rect 8688 -24110 8722 -24094
rect 8688 -24702 8722 -24686
rect 9706 -24110 9740 -24094
rect 9706 -24702 9740 -24686
rect 10724 -24110 10758 -24094
rect 10724 -24702 10758 -24686
rect 11742 -24110 11776 -24094
rect 11742 -24702 11776 -24686
rect 12760 -24110 12794 -24094
rect 12760 -24702 12794 -24686
rect 13778 -24110 13812 -24094
rect 13778 -24702 13812 -24686
rect 14796 -24110 14830 -24094
rect 14796 -24702 14830 -24686
rect 15814 -24110 15848 -24094
rect 15814 -24702 15848 -24686
rect 16832 -24110 16866 -24094
rect 16832 -24702 16866 -24686
rect 17850 -24110 17884 -24094
rect 17850 -24702 17884 -24686
rect 18868 -24110 18902 -24094
rect 18868 -24702 18902 -24686
rect 19886 -24110 19920 -24094
rect 19886 -24702 19920 -24686
rect 20904 -24110 20938 -24094
rect 20904 -24702 20938 -24686
rect 21922 -24110 21956 -24094
rect 21922 -24702 21956 -24686
rect 22940 -24110 22974 -24094
rect 22940 -24702 22974 -24686
rect 4088 -24736 4148 -24734
rect 10200 -24736 10260 -24734
rect 12234 -24736 12294 -24734
rect 16300 -24736 16360 -24730
rect 20376 -24736 20436 -24734
rect 21392 -24736 21452 -24734
rect 2812 -24770 2828 -24736
rect 3384 -24770 3400 -24736
rect 3830 -24770 3846 -24736
rect 4402 -24770 4418 -24736
rect 4848 -24770 4864 -24736
rect 5420 -24770 5436 -24736
rect 5866 -24770 5882 -24736
rect 6438 -24770 6454 -24736
rect 6884 -24770 6900 -24736
rect 7456 -24770 7472 -24736
rect 7902 -24770 7918 -24736
rect 8474 -24770 8490 -24736
rect 8920 -24770 8936 -24736
rect 9492 -24770 9508 -24736
rect 9938 -24770 9954 -24736
rect 10510 -24770 10526 -24736
rect 10956 -24770 10972 -24736
rect 11528 -24770 11544 -24736
rect 11974 -24770 11990 -24736
rect 12546 -24770 12562 -24736
rect 12992 -24770 13008 -24736
rect 13564 -24770 13580 -24736
rect 14010 -24770 14026 -24736
rect 14582 -24770 14598 -24736
rect 15028 -24770 15044 -24736
rect 15600 -24770 15616 -24736
rect 16046 -24770 16062 -24736
rect 16618 -24770 16634 -24736
rect 17064 -24770 17080 -24736
rect 17636 -24770 17652 -24736
rect 18082 -24770 18098 -24736
rect 18654 -24770 18670 -24736
rect 19100 -24770 19116 -24736
rect 19672 -24770 19688 -24736
rect 20118 -24770 20134 -24736
rect 20690 -24770 20706 -24736
rect 21136 -24770 21152 -24736
rect 21708 -24770 21724 -24736
rect 22154 -24770 22170 -24736
rect 22726 -24770 22742 -24736
rect 3086 -25002 3168 -24978
rect 3086 -25036 3110 -25002
rect 3144 -25036 3168 -25002
rect 3086 -25060 3168 -25036
rect 4104 -25002 4186 -24978
rect 4104 -25036 4128 -25002
rect 4162 -25036 4186 -25002
rect 4104 -25060 4186 -25036
rect 5122 -25002 5204 -24978
rect 5122 -25036 5146 -25002
rect 5180 -25036 5204 -25002
rect 5122 -25060 5204 -25036
rect 6140 -25002 6222 -24978
rect 6140 -25036 6164 -25002
rect 6198 -25036 6222 -25002
rect 6140 -25060 6222 -25036
rect 7158 -25002 7240 -24978
rect 7158 -25036 7182 -25002
rect 7216 -25036 7240 -25002
rect 7158 -25060 7240 -25036
rect 8176 -25002 8258 -24978
rect 8176 -25036 8200 -25002
rect 8234 -25036 8258 -25002
rect 8176 -25060 8258 -25036
rect 9194 -25002 9276 -24978
rect 9194 -25036 9218 -25002
rect 9252 -25036 9276 -25002
rect 9194 -25060 9276 -25036
rect 10212 -25002 10294 -24978
rect 10212 -25036 10236 -25002
rect 10270 -25036 10294 -25002
rect 10212 -25060 10294 -25036
rect 11230 -25002 11312 -24978
rect 11230 -25036 11254 -25002
rect 11288 -25036 11312 -25002
rect 11230 -25060 11312 -25036
rect 12248 -25002 12330 -24978
rect 12248 -25036 12272 -25002
rect 12306 -25036 12330 -25002
rect 12248 -25060 12330 -25036
rect 13266 -25002 13348 -24978
rect 13266 -25036 13290 -25002
rect 13324 -25036 13348 -25002
rect 13266 -25060 13348 -25036
rect 14284 -25002 14366 -24978
rect 14284 -25036 14308 -25002
rect 14342 -25036 14366 -25002
rect 14284 -25060 14366 -25036
rect 15302 -25002 15384 -24978
rect 15302 -25036 15326 -25002
rect 15360 -25036 15384 -25002
rect 15302 -25060 15384 -25036
rect 16320 -25002 16402 -24978
rect 16320 -25036 16344 -25002
rect 16378 -25036 16402 -25002
rect 16320 -25060 16402 -25036
rect 17338 -25002 17420 -24978
rect 17338 -25036 17362 -25002
rect 17396 -25036 17420 -25002
rect 17338 -25060 17420 -25036
rect 18356 -25002 18438 -24978
rect 18356 -25036 18380 -25002
rect 18414 -25036 18438 -25002
rect 18356 -25060 18438 -25036
rect 19374 -25002 19456 -24978
rect 19374 -25036 19398 -25002
rect 19432 -25036 19456 -25002
rect 19374 -25060 19456 -25036
rect 20392 -25002 20474 -24978
rect 20392 -25036 20416 -25002
rect 20450 -25036 20474 -25002
rect 20392 -25060 20474 -25036
rect 21410 -25002 21492 -24978
rect 21410 -25036 21434 -25002
rect 21468 -25036 21492 -25002
rect 21410 -25060 21492 -25036
rect 22428 -25002 22510 -24978
rect 22428 -25036 22452 -25002
rect 22486 -25036 22510 -25002
rect 22428 -25060 22510 -25036
rect -9818 -25102 -9802 -25068
rect -9246 -25102 -9230 -25068
rect -8800 -25102 -8784 -25068
rect -8228 -25102 -8212 -25068
rect -7782 -25102 -7766 -25068
rect -7210 -25102 -7194 -25068
rect -6764 -25102 -6748 -25068
rect -6192 -25102 -6176 -25068
rect -5746 -25102 -5730 -25068
rect -5174 -25102 -5158 -25068
rect -4728 -25102 -4712 -25068
rect -4156 -25102 -4140 -25068
rect -3710 -25102 -3694 -25068
rect -3138 -25102 -3122 -25068
rect -2692 -25102 -2676 -25068
rect -2120 -25102 -2104 -25068
rect -1674 -25102 -1658 -25068
rect -1102 -25102 -1086 -25068
rect -656 -25102 -640 -25068
rect -84 -25102 -68 -25068
rect -10050 -25152 -10016 -25136
rect -10050 -25744 -10016 -25728
rect -9032 -25152 -8998 -25136
rect -9032 -25744 -8998 -25728
rect -8014 -25152 -7980 -25136
rect -8014 -25744 -7980 -25728
rect -6996 -25152 -6962 -25136
rect -6996 -25744 -6962 -25728
rect -5978 -25152 -5944 -25136
rect -5978 -25744 -5944 -25728
rect -4960 -25152 -4926 -25136
rect -4960 -25744 -4926 -25728
rect -3942 -25152 -3908 -25136
rect -3942 -25744 -3908 -25728
rect -2924 -25152 -2890 -25136
rect -2924 -25744 -2890 -25728
rect -1906 -25152 -1872 -25136
rect -1906 -25744 -1872 -25728
rect -888 -25152 -854 -25136
rect -888 -25744 -854 -25728
rect 130 -25152 164 -25136
rect 2812 -25292 2828 -25258
rect 3384 -25292 3400 -25258
rect 3830 -25292 3846 -25258
rect 4402 -25292 4418 -25258
rect 4848 -25292 4864 -25258
rect 5420 -25292 5436 -25258
rect 5866 -25292 5882 -25258
rect 6438 -25292 6454 -25258
rect 6884 -25292 6900 -25258
rect 7456 -25292 7472 -25258
rect 7902 -25292 7918 -25258
rect 8474 -25292 8490 -25258
rect 8920 -25292 8936 -25258
rect 9492 -25292 9508 -25258
rect 9938 -25292 9954 -25258
rect 10510 -25292 10526 -25258
rect 10956 -25292 10972 -25258
rect 11528 -25292 11544 -25258
rect 11974 -25292 11990 -25258
rect 12546 -25292 12562 -25258
rect 12992 -25292 13008 -25258
rect 13564 -25292 13580 -25258
rect 14010 -25292 14026 -25258
rect 14582 -25292 14598 -25258
rect 15028 -25292 15044 -25258
rect 15600 -25292 15616 -25258
rect 16046 -25292 16062 -25258
rect 16618 -25292 16634 -25258
rect 17064 -25292 17080 -25258
rect 17636 -25292 17652 -25258
rect 18082 -25292 18098 -25258
rect 18654 -25292 18670 -25258
rect 19100 -25292 19116 -25258
rect 19672 -25292 19688 -25258
rect 20118 -25292 20134 -25258
rect 20690 -25292 20706 -25258
rect 21136 -25292 21152 -25258
rect 21708 -25292 21724 -25258
rect 22154 -25292 22170 -25258
rect 22726 -25292 22742 -25258
rect 130 -25744 164 -25728
rect 2580 -25342 2614 -25326
rect -9818 -25812 -9802 -25778
rect -9246 -25812 -9230 -25778
rect -8800 -25812 -8784 -25778
rect -8228 -25812 -8212 -25778
rect -7782 -25812 -7766 -25778
rect -7210 -25812 -7194 -25778
rect -6764 -25812 -6748 -25778
rect -6192 -25812 -6176 -25778
rect -5746 -25812 -5730 -25778
rect -5174 -25812 -5158 -25778
rect -4728 -25812 -4712 -25778
rect -4156 -25812 -4140 -25778
rect -3710 -25812 -3694 -25778
rect -3138 -25812 -3122 -25778
rect -2692 -25812 -2676 -25778
rect -2120 -25812 -2104 -25778
rect -1674 -25812 -1658 -25778
rect -1102 -25812 -1086 -25778
rect -656 -25812 -640 -25778
rect -84 -25812 -68 -25778
rect 2580 -25934 2614 -25918
rect 3598 -25342 3632 -25326
rect 3598 -25934 3632 -25918
rect 4616 -25342 4650 -25326
rect 4616 -25934 4650 -25918
rect 5634 -25342 5668 -25326
rect 5634 -25934 5668 -25918
rect 6652 -25342 6686 -25326
rect 6652 -25934 6686 -25918
rect 7670 -25342 7704 -25326
rect 7670 -25934 7704 -25918
rect 8688 -25342 8722 -25326
rect 8688 -25934 8722 -25918
rect 9706 -25342 9740 -25326
rect 9706 -25934 9740 -25918
rect 10724 -25342 10758 -25326
rect 10724 -25934 10758 -25918
rect 11742 -25342 11776 -25326
rect 11742 -25934 11776 -25918
rect 12760 -25342 12794 -25326
rect 12760 -25934 12794 -25918
rect 13778 -25342 13812 -25326
rect 13778 -25934 13812 -25918
rect 14796 -25342 14830 -25326
rect 14796 -25934 14830 -25918
rect 15814 -25342 15848 -25326
rect 15814 -25934 15848 -25918
rect 16832 -25342 16866 -25326
rect 16832 -25934 16866 -25918
rect 17850 -25342 17884 -25326
rect 17850 -25934 17884 -25918
rect 18868 -25342 18902 -25326
rect 18868 -25934 18902 -25918
rect 19886 -25342 19920 -25326
rect 19886 -25934 19920 -25918
rect 20904 -25342 20938 -25326
rect 20904 -25934 20938 -25918
rect 21922 -25342 21956 -25326
rect 21922 -25934 21956 -25918
rect 22940 -25342 22974 -25326
rect 22940 -25934 22974 -25918
rect 2812 -26002 2828 -25968
rect 3384 -26002 3400 -25968
rect 3830 -26002 3846 -25968
rect 4402 -26002 4418 -25968
rect 4848 -26002 4864 -25968
rect 5420 -26002 5436 -25968
rect 5866 -26002 5882 -25968
rect 6438 -26002 6454 -25968
rect 6884 -26002 6900 -25968
rect 7456 -26002 7472 -25968
rect 7902 -26002 7918 -25968
rect 8474 -26002 8490 -25968
rect 8920 -26002 8936 -25968
rect 9492 -26002 9508 -25968
rect 9938 -26002 9954 -25968
rect 10510 -26002 10526 -25968
rect 10956 -26002 10972 -25968
rect 11528 -26002 11544 -25968
rect 11974 -26002 11990 -25968
rect 12546 -26002 12562 -25968
rect 12992 -26002 13008 -25968
rect 13564 -26002 13580 -25968
rect 14010 -26002 14026 -25968
rect 14582 -26002 14598 -25968
rect 15028 -26002 15044 -25968
rect 15600 -26002 15616 -25968
rect 16046 -26002 16062 -25968
rect 16618 -26002 16634 -25968
rect 17064 -26002 17080 -25968
rect 17636 -26002 17652 -25968
rect 18082 -26002 18098 -25968
rect 18654 -26002 18670 -25968
rect 19100 -26002 19116 -25968
rect 19672 -26002 19688 -25968
rect 20118 -26002 20134 -25968
rect 20690 -26002 20706 -25968
rect 21136 -26002 21152 -25968
rect 21708 -26002 21724 -25968
rect 22154 -26002 22170 -25968
rect 22726 -26002 22742 -25968
rect -10216 -26098 -10134 -26074
rect -10216 -26132 -10192 -26098
rect -10158 -26132 -10134 -26098
rect -10216 -26156 -10134 -26132
rect -9198 -26098 -9116 -26074
rect -9198 -26132 -9174 -26098
rect -9140 -26132 -9116 -26098
rect -9198 -26156 -9116 -26132
rect -8180 -26098 -8098 -26074
rect -8180 -26132 -8156 -26098
rect -8122 -26132 -8098 -26098
rect -8180 -26156 -8098 -26132
rect -7162 -26098 -7080 -26074
rect -7162 -26132 -7138 -26098
rect -7104 -26132 -7080 -26098
rect -7162 -26156 -7080 -26132
rect -6144 -26098 -6062 -26074
rect -6144 -26132 -6120 -26098
rect -6086 -26132 -6062 -26098
rect -6144 -26156 -6062 -26132
rect -5126 -26098 -5044 -26074
rect -5126 -26132 -5102 -26098
rect -5068 -26132 -5044 -26098
rect -5126 -26156 -5044 -26132
rect -4108 -26098 -4026 -26074
rect -4108 -26132 -4084 -26098
rect -4050 -26132 -4026 -26098
rect -4108 -26156 -4026 -26132
rect -3090 -26098 -3008 -26074
rect -3090 -26132 -3066 -26098
rect -3032 -26132 -3008 -26098
rect -3090 -26156 -3008 -26132
rect -2072 -26098 -1990 -26074
rect -2072 -26132 -2048 -26098
rect -2014 -26132 -1990 -26098
rect -2072 -26156 -1990 -26132
rect -1054 -26098 -972 -26074
rect -1054 -26132 -1030 -26098
rect -996 -26132 -972 -26098
rect -1054 -26156 -972 -26132
rect -36 -26098 46 -26074
rect -36 -26132 -12 -26098
rect 22 -26132 46 -26098
rect -36 -26156 46 -26132
rect 3074 -26180 3156 -26156
rect 3074 -26214 3098 -26180
rect 3132 -26214 3156 -26180
rect 3074 -26238 3156 -26214
rect 4092 -26180 4174 -26156
rect 4092 -26214 4116 -26180
rect 4150 -26214 4174 -26180
rect 4092 -26238 4174 -26214
rect 5110 -26180 5192 -26156
rect 5110 -26214 5134 -26180
rect 5168 -26214 5192 -26180
rect 5110 -26238 5192 -26214
rect 6128 -26180 6210 -26156
rect 6128 -26214 6152 -26180
rect 6186 -26214 6210 -26180
rect 6128 -26238 6210 -26214
rect 7146 -26180 7228 -26156
rect 7146 -26214 7170 -26180
rect 7204 -26214 7228 -26180
rect 7146 -26238 7228 -26214
rect 8164 -26180 8246 -26156
rect 8164 -26214 8188 -26180
rect 8222 -26214 8246 -26180
rect 8164 -26238 8246 -26214
rect 9182 -26180 9264 -26156
rect 9182 -26214 9206 -26180
rect 9240 -26214 9264 -26180
rect 9182 -26238 9264 -26214
rect 10200 -26180 10282 -26156
rect 10200 -26214 10224 -26180
rect 10258 -26214 10282 -26180
rect 10200 -26238 10282 -26214
rect 11218 -26180 11300 -26156
rect 11218 -26214 11242 -26180
rect 11276 -26214 11300 -26180
rect 11218 -26238 11300 -26214
rect 12236 -26180 12318 -26156
rect 12236 -26214 12260 -26180
rect 12294 -26214 12318 -26180
rect 12236 -26238 12318 -26214
rect 13254 -26180 13336 -26156
rect 13254 -26214 13278 -26180
rect 13312 -26214 13336 -26180
rect 13254 -26238 13336 -26214
rect 14272 -26180 14354 -26156
rect 14272 -26214 14296 -26180
rect 14330 -26214 14354 -26180
rect 14272 -26238 14354 -26214
rect 15290 -26180 15372 -26156
rect 15290 -26214 15314 -26180
rect 15348 -26214 15372 -26180
rect 15290 -26238 15372 -26214
rect 16308 -26180 16390 -26156
rect 16308 -26214 16332 -26180
rect 16366 -26214 16390 -26180
rect 16308 -26238 16390 -26214
rect 17326 -26180 17408 -26156
rect 17326 -26214 17350 -26180
rect 17384 -26214 17408 -26180
rect 17326 -26238 17408 -26214
rect 18344 -26180 18426 -26156
rect 18344 -26214 18368 -26180
rect 18402 -26214 18426 -26180
rect 18344 -26238 18426 -26214
rect 19362 -26180 19444 -26156
rect 19362 -26214 19386 -26180
rect 19420 -26214 19444 -26180
rect 19362 -26238 19444 -26214
rect 20380 -26180 20462 -26156
rect 20380 -26214 20404 -26180
rect 20438 -26214 20462 -26180
rect 20380 -26238 20462 -26214
rect 21398 -26180 21480 -26156
rect 21398 -26214 21422 -26180
rect 21456 -26214 21480 -26180
rect 21398 -26238 21480 -26214
rect 22416 -26180 22498 -26156
rect 22416 -26214 22440 -26180
rect 22474 -26214 22498 -26180
rect 22416 -26238 22498 -26214
rect -12322 -27222 -12222 -27060
rect 24822 -27222 24922 -27060
<< viali >>
rect 478 4222 540 4322
rect 540 4222 24660 4322
rect 24660 4222 24722 4322
rect 378 -9728 478 3702
rect 6782 1521 7246 1555
rect 7800 1521 8264 1555
rect 8818 1521 9282 1555
rect 9836 1521 10300 1555
rect 10854 1521 11318 1555
rect 11872 1521 12336 1555
rect 12890 1521 13354 1555
rect 13908 1521 14372 1555
rect 14926 1521 15390 1555
rect 15944 1521 16408 1555
rect 16962 1521 17426 1555
rect 17980 1521 18444 1555
rect 18998 1521 19462 1555
rect 20016 1521 20480 1555
rect 21034 1521 21498 1555
rect 22052 1521 22516 1555
rect 6488 886 6522 1462
rect 7506 886 7540 1462
rect 8524 886 8558 1462
rect 9542 886 9576 1462
rect 10560 886 10594 1462
rect 11578 886 11612 1462
rect 12596 886 12630 1462
rect 13614 886 13648 1462
rect 14632 886 14666 1462
rect 15650 886 15684 1462
rect 16668 886 16702 1462
rect 17686 886 17720 1462
rect 18704 886 18738 1462
rect 19722 886 19756 1462
rect 20740 886 20774 1462
rect 21758 886 21792 1462
rect 22776 886 22810 1462
rect 6782 793 7246 827
rect 7800 793 8264 827
rect 8818 793 9282 827
rect 9836 793 10300 827
rect 10854 793 11318 827
rect 11872 793 12336 827
rect 12890 793 13354 827
rect 13908 793 14372 827
rect 14926 793 15390 827
rect 15944 793 16408 827
rect 16962 793 17426 827
rect 17980 793 18444 827
rect 18998 793 19462 827
rect 20016 793 20480 827
rect 21034 793 21498 827
rect 22052 793 22516 827
rect 6782 385 7246 419
rect 7800 385 8264 419
rect 8818 385 9282 419
rect 9836 385 10300 419
rect 10854 385 11318 419
rect 11872 385 12336 419
rect 12890 385 13354 419
rect 13908 385 14372 419
rect 14926 385 15390 419
rect 15944 385 16408 419
rect 16962 385 17426 419
rect 17980 385 18444 419
rect 18998 385 19462 419
rect 20016 385 20480 419
rect 21034 385 21498 419
rect 22052 385 22516 419
rect 6488 -250 6522 326
rect 7506 -250 7540 326
rect 8524 -250 8558 326
rect 9542 -250 9576 326
rect 10560 -250 10594 326
rect 11578 -250 11612 326
rect 12596 -250 12630 326
rect 13614 -250 13648 326
rect 14632 -250 14666 326
rect 15650 -250 15684 326
rect 16668 -250 16702 326
rect 17686 -250 17720 326
rect 18704 -250 18738 326
rect 19722 -250 19756 326
rect 20740 -250 20774 326
rect 21758 -250 21792 326
rect 22776 -250 22810 326
rect 6782 -343 7246 -309
rect 7800 -343 8264 -309
rect 8818 -343 9282 -309
rect 9836 -343 10300 -309
rect 10854 -343 11318 -309
rect 11872 -343 12336 -309
rect 12890 -343 13354 -309
rect 13908 -343 14372 -309
rect 14926 -343 15390 -309
rect 15944 -343 16408 -309
rect 16962 -343 17426 -309
rect 17980 -343 18444 -309
rect 18998 -343 19462 -309
rect 20016 -343 20480 -309
rect 21034 -343 21498 -309
rect 22052 -343 22516 -309
rect 6782 -751 7246 -717
rect 7800 -751 8264 -717
rect 8818 -751 9282 -717
rect 9836 -751 10300 -717
rect 10854 -751 11318 -717
rect 11872 -751 12336 -717
rect 12890 -751 13354 -717
rect 13908 -751 14372 -717
rect 14926 -751 15390 -717
rect 15944 -751 16408 -717
rect 16962 -751 17426 -717
rect 17980 -751 18444 -717
rect 18998 -751 19462 -717
rect 20016 -751 20480 -717
rect 21034 -751 21498 -717
rect 22052 -751 22516 -717
rect 6488 -1386 6522 -810
rect 7506 -1386 7540 -810
rect 8524 -1386 8558 -810
rect 9542 -1386 9576 -810
rect 10560 -1386 10594 -810
rect 11578 -1386 11612 -810
rect 12596 -1386 12630 -810
rect 13614 -1386 13648 -810
rect 14632 -1386 14666 -810
rect 15650 -1386 15684 -810
rect 16668 -1386 16702 -810
rect 17686 -1386 17720 -810
rect 18704 -1386 18738 -810
rect 19722 -1386 19756 -810
rect 20740 -1386 20774 -810
rect 21758 -1386 21792 -810
rect 22776 -1386 22810 -810
rect 6782 -1479 7246 -1445
rect 7800 -1479 8264 -1445
rect 8818 -1479 9282 -1445
rect 9836 -1479 10300 -1445
rect 10854 -1479 11318 -1445
rect 11872 -1479 12336 -1445
rect 12890 -1479 13354 -1445
rect 13908 -1479 14372 -1445
rect 14926 -1479 15390 -1445
rect 15944 -1479 16408 -1445
rect 16962 -1479 17426 -1445
rect 17980 -1479 18444 -1445
rect 18998 -1479 19462 -1445
rect 20016 -1479 20480 -1445
rect 21034 -1479 21498 -1445
rect 22052 -1479 22516 -1445
rect 7976 -2389 8440 -2355
rect 8994 -2389 9458 -2355
rect 10012 -2389 10476 -2355
rect 11030 -2389 11494 -2355
rect 12048 -2389 12512 -2355
rect 13066 -2389 13530 -2355
rect 14084 -2389 14548 -2355
rect 15102 -2389 15566 -2355
rect 16120 -2389 16584 -2355
rect 17138 -2389 17602 -2355
rect 18156 -2389 18620 -2355
rect 19174 -2389 19638 -2355
rect 20192 -2389 20656 -2355
rect 21210 -2389 21674 -2355
rect 7682 -3024 7716 -2448
rect 8700 -3024 8734 -2448
rect 9718 -3024 9752 -2448
rect 10736 -3024 10770 -2448
rect 11754 -3024 11788 -2448
rect 12772 -3024 12806 -2448
rect 13790 -3024 13824 -2448
rect 14808 -3024 14842 -2448
rect 15826 -3024 15860 -2448
rect 16844 -3024 16878 -2448
rect 17862 -3024 17896 -2448
rect 18880 -3024 18914 -2448
rect 19898 -3024 19932 -2448
rect 20916 -3024 20950 -2448
rect 21934 -3024 21968 -2448
rect 7976 -3117 8440 -3083
rect 8994 -3117 9458 -3083
rect 10012 -3117 10476 -3083
rect 11030 -3117 11494 -3083
rect 12048 -3117 12512 -3083
rect 13066 -3117 13530 -3083
rect 14084 -3117 14548 -3083
rect 15102 -3117 15566 -3083
rect 16120 -3117 16584 -3083
rect 17138 -3117 17602 -3083
rect 18156 -3117 18620 -3083
rect 19174 -3117 19638 -3083
rect 20192 -3117 20656 -3083
rect 21210 -3117 21674 -3083
rect 7976 -3421 8440 -3387
rect 8994 -3421 9458 -3387
rect 10012 -3421 10476 -3387
rect 11030 -3421 11494 -3387
rect 12048 -3421 12512 -3387
rect 13066 -3421 13530 -3387
rect 14084 -3421 14548 -3387
rect 15102 -3421 15566 -3387
rect 16120 -3421 16584 -3387
rect 17138 -3421 17602 -3387
rect 18156 -3421 18620 -3387
rect 19174 -3421 19638 -3387
rect 20192 -3421 20656 -3387
rect 21210 -3421 21674 -3387
rect 7682 -4056 7716 -3480
rect 8700 -4056 8734 -3480
rect 9718 -4056 9752 -3480
rect 10736 -4056 10770 -3480
rect 11754 -4056 11788 -3480
rect 12772 -4056 12806 -3480
rect 13790 -4056 13824 -3480
rect 14808 -4056 14842 -3480
rect 15826 -4056 15860 -3480
rect 16844 -4056 16878 -3480
rect 17862 -4056 17896 -3480
rect 18880 -4056 18914 -3480
rect 19898 -4056 19932 -3480
rect 20916 -4056 20950 -3480
rect 21934 -4056 21968 -3480
rect 7976 -4149 8440 -4115
rect 8994 -4149 9458 -4115
rect 10012 -4149 10476 -4115
rect 11030 -4149 11494 -4115
rect 12048 -4149 12512 -4115
rect 13066 -4149 13530 -4115
rect 14084 -4149 14548 -4115
rect 15102 -4149 15566 -4115
rect 16120 -4149 16584 -4115
rect 17138 -4149 17602 -4115
rect 18156 -4149 18620 -4115
rect 19174 -4149 19638 -4115
rect 20192 -4149 20656 -4115
rect 21210 -4149 21674 -4115
rect 7768 -5025 8232 -4991
rect 8786 -5025 9250 -4991
rect 9804 -5025 10268 -4991
rect 10822 -5025 11286 -4991
rect 11840 -5025 12304 -4991
rect 12858 -5025 13322 -4991
rect 13876 -5025 14340 -4991
rect 14894 -5025 15358 -4991
rect 15912 -5025 16376 -4991
rect 16930 -5025 17394 -4991
rect 17948 -5025 18412 -4991
rect 18966 -5025 19430 -4991
rect 19984 -5025 20448 -4991
rect 21002 -5025 21466 -4991
rect 22020 -5025 22484 -4991
rect 2464 -5129 2928 -5095
rect 3482 -5129 3946 -5095
rect 4500 -5129 4964 -5095
rect 5518 -5129 5982 -5095
rect 2170 -5764 2204 -5188
rect 3188 -5764 3222 -5188
rect 4206 -5764 4240 -5188
rect 5224 -5764 5258 -5188
rect 6242 -5764 6276 -5188
rect 7474 -5660 7508 -5084
rect 8492 -5660 8526 -5084
rect 9510 -5660 9544 -5084
rect 10528 -5660 10562 -5084
rect 11546 -5660 11580 -5084
rect 12564 -5660 12598 -5084
rect 13582 -5660 13616 -5084
rect 14600 -5660 14634 -5084
rect 15618 -5660 15652 -5084
rect 16636 -5660 16670 -5084
rect 17654 -5660 17688 -5084
rect 18672 -5660 18706 -5084
rect 19690 -5660 19724 -5084
rect 20708 -5660 20742 -5084
rect 21726 -5660 21760 -5084
rect 22744 -5660 22778 -5084
rect 7768 -5753 8232 -5719
rect 8786 -5753 9250 -5719
rect 9804 -5753 10268 -5719
rect 10822 -5753 11286 -5719
rect 11840 -5753 12304 -5719
rect 12858 -5753 13322 -5719
rect 13876 -5753 14340 -5719
rect 14894 -5753 15358 -5719
rect 15912 -5753 16376 -5719
rect 16930 -5753 17394 -5719
rect 17948 -5753 18412 -5719
rect 18966 -5753 19430 -5719
rect 19984 -5753 20448 -5719
rect 21002 -5753 21466 -5719
rect 22020 -5753 22484 -5719
rect 2464 -5857 2928 -5823
rect 3482 -5857 3946 -5823
rect 4500 -5857 4964 -5823
rect 5518 -5857 5982 -5823
rect 2464 -6161 2928 -6127
rect 3482 -6161 3946 -6127
rect 4500 -6161 4964 -6127
rect 5518 -6161 5982 -6127
rect 2170 -6796 2204 -6220
rect 3188 -6796 3222 -6220
rect 4206 -6796 4240 -6220
rect 5224 -6796 5258 -6220
rect 6242 -6796 6276 -6220
rect 7768 -6281 8232 -6247
rect 8786 -6281 9250 -6247
rect 9804 -6281 10268 -6247
rect 10822 -6281 11286 -6247
rect 11840 -6281 12304 -6247
rect 12858 -6281 13322 -6247
rect 13876 -6281 14340 -6247
rect 14894 -6281 15358 -6247
rect 15912 -6281 16376 -6247
rect 16930 -6281 17394 -6247
rect 17948 -6281 18412 -6247
rect 18966 -6281 19430 -6247
rect 19984 -6281 20448 -6247
rect 21002 -6281 21466 -6247
rect 22020 -6281 22484 -6247
rect 2464 -6889 2928 -6855
rect 3482 -6889 3946 -6855
rect 4500 -6889 4964 -6855
rect 5518 -6889 5982 -6855
rect 7474 -6916 7508 -6340
rect 8492 -6916 8526 -6340
rect 9510 -6916 9544 -6340
rect 10528 -6916 10562 -6340
rect 11546 -6916 11580 -6340
rect 12564 -6916 12598 -6340
rect 13582 -6916 13616 -6340
rect 14600 -6916 14634 -6340
rect 15618 -6916 15652 -6340
rect 16636 -6916 16670 -6340
rect 17654 -6916 17688 -6340
rect 18672 -6916 18706 -6340
rect 19690 -6916 19724 -6340
rect 20708 -6916 20742 -6340
rect 21726 -6916 21760 -6340
rect 22744 -6916 22778 -6340
rect 7768 -7009 8232 -6975
rect 8786 -7009 9250 -6975
rect 9804 -7009 10268 -6975
rect 10822 -7009 11286 -6975
rect 11840 -7009 12304 -6975
rect 12858 -7009 13322 -6975
rect 13876 -7009 14340 -6975
rect 14894 -7009 15358 -6975
rect 15912 -7009 16376 -6975
rect 16930 -7009 17394 -6975
rect 17948 -7009 18412 -6975
rect 18966 -7009 19430 -6975
rect 19984 -7009 20448 -6975
rect 21002 -7009 21466 -6975
rect 22020 -7009 22484 -6975
rect 2464 -7193 2928 -7159
rect 3482 -7193 3946 -7159
rect 4500 -7193 4964 -7159
rect 5518 -7193 5982 -7159
rect 2170 -7828 2204 -7252
rect 3188 -7828 3222 -7252
rect 4206 -7828 4240 -7252
rect 5224 -7828 5258 -7252
rect 6242 -7828 6276 -7252
rect 7768 -7537 8232 -7503
rect 8786 -7537 9250 -7503
rect 9804 -7537 10268 -7503
rect 10822 -7537 11286 -7503
rect 11840 -7537 12304 -7503
rect 12858 -7537 13322 -7503
rect 13876 -7537 14340 -7503
rect 14894 -7537 15358 -7503
rect 15912 -7537 16376 -7503
rect 16930 -7537 17394 -7503
rect 17948 -7537 18412 -7503
rect 18966 -7537 19430 -7503
rect 19984 -7537 20448 -7503
rect 21002 -7537 21466 -7503
rect 22020 -7537 22484 -7503
rect 2464 -7921 2928 -7887
rect 3482 -7921 3946 -7887
rect 4500 -7921 4964 -7887
rect 5518 -7921 5982 -7887
rect 7474 -8172 7508 -7596
rect 8492 -8172 8526 -7596
rect 9510 -8172 9544 -7596
rect 10528 -8172 10562 -7596
rect 11546 -8172 11580 -7596
rect 12564 -8172 12598 -7596
rect 13582 -8172 13616 -7596
rect 14600 -8172 14634 -7596
rect 15618 -8172 15652 -7596
rect 16636 -8172 16670 -7596
rect 17654 -8172 17688 -7596
rect 18672 -8172 18706 -7596
rect 19690 -8172 19724 -7596
rect 20708 -8172 20742 -7596
rect 21726 -8172 21760 -7596
rect 22744 -8172 22778 -7596
rect 2464 -8225 2928 -8191
rect 3482 -8225 3946 -8191
rect 4500 -8225 4964 -8191
rect 5518 -8225 5982 -8191
rect 7768 -8265 8232 -8231
rect 8786 -8265 9250 -8231
rect 9804 -8265 10268 -8231
rect 10822 -8265 11286 -8231
rect 11840 -8265 12304 -8231
rect 12858 -8265 13322 -8231
rect 13876 -8265 14340 -8231
rect 14894 -8265 15358 -8231
rect 15912 -8265 16376 -8231
rect 16930 -8265 17394 -8231
rect 17948 -8265 18412 -8231
rect 18966 -8265 19430 -8231
rect 19984 -8265 20448 -8231
rect 21002 -8265 21466 -8231
rect 22020 -8265 22484 -8231
rect 2170 -8860 2204 -8284
rect 3188 -8860 3222 -8284
rect 4206 -8860 4240 -8284
rect 5224 -8860 5258 -8284
rect 6242 -8860 6276 -8284
rect 7768 -8793 8232 -8759
rect 8786 -8793 9250 -8759
rect 9804 -8793 10268 -8759
rect 10822 -8793 11286 -8759
rect 11840 -8793 12304 -8759
rect 12858 -8793 13322 -8759
rect 13876 -8793 14340 -8759
rect 14894 -8793 15358 -8759
rect 15912 -8793 16376 -8759
rect 16930 -8793 17394 -8759
rect 17948 -8793 18412 -8759
rect 18966 -8793 19430 -8759
rect 19984 -8793 20448 -8759
rect 21002 -8793 21466 -8759
rect 22020 -8793 22484 -8759
rect 2464 -8953 2928 -8919
rect 3482 -8953 3946 -8919
rect 4500 -8953 4964 -8919
rect 5518 -8953 5982 -8919
rect 7474 -9428 7508 -8852
rect 8492 -9428 8526 -8852
rect 9510 -9428 9544 -8852
rect 10528 -9428 10562 -8852
rect 11546 -9428 11580 -8852
rect 12564 -9428 12598 -8852
rect 13582 -9428 13616 -8852
rect 14600 -9428 14634 -8852
rect 15618 -9428 15652 -8852
rect 16636 -9428 16670 -8852
rect 17654 -9428 17688 -8852
rect 18672 -9428 18706 -8852
rect 19690 -9428 19724 -8852
rect 20708 -9428 20742 -8852
rect 21726 -9428 21760 -8852
rect 22744 -9428 22778 -8852
rect 7768 -9521 8232 -9487
rect 8786 -9521 9250 -9487
rect 9804 -9521 10268 -9487
rect 10822 -9521 11286 -9487
rect 11840 -9521 12304 -9487
rect 12858 -9521 13322 -9487
rect 13876 -9521 14340 -9487
rect 14894 -9521 15358 -9487
rect 15912 -9521 16376 -9487
rect 16930 -9521 17394 -9487
rect 17948 -9521 18412 -9487
rect 18966 -9521 19430 -9487
rect 19984 -9521 20448 -9487
rect 21002 -9521 21466 -9487
rect 22020 -9521 22484 -9487
rect 24722 -9728 24822 3702
rect 478 -10348 540 -10248
rect 540 -10348 24660 -10248
rect 24660 -10348 24722 -10248
rect -12222 -11278 -12160 -11178
rect -12160 -11278 24760 -11178
rect 24760 -11278 24822 -11178
rect 2876 -11998 3340 -11964
rect 3894 -11998 4358 -11964
rect 4912 -11998 5376 -11964
rect 5930 -11998 6394 -11964
rect 6948 -11998 7412 -11964
rect 7966 -11998 8430 -11964
rect 8984 -11998 9448 -11964
rect 10002 -11998 10466 -11964
rect 11020 -11998 11484 -11964
rect 12038 -11998 12502 -11964
rect 13056 -11998 13520 -11964
rect 14074 -11998 14538 -11964
rect 15092 -11998 15556 -11964
rect 16110 -11998 16574 -11964
rect 17128 -11998 17592 -11964
rect 18146 -11998 18610 -11964
rect 19164 -11998 19628 -11964
rect 20182 -11998 20646 -11964
rect 21200 -11998 21664 -11964
rect 22218 -11998 22682 -11964
rect -12322 -26330 -12222 -12070
rect -8890 -12474 -8426 -12440
rect -7872 -12474 -7408 -12440
rect -6854 -12474 -6390 -12440
rect -5836 -12474 -5372 -12440
rect -4818 -12474 -4354 -12440
rect -3800 -12474 -3336 -12440
rect -2782 -12474 -2318 -12440
rect -1764 -12474 -1300 -12440
rect -746 -12474 -282 -12440
rect -9184 -13100 -9150 -12524
rect -8166 -13100 -8132 -12524
rect -7148 -13100 -7114 -12524
rect -6130 -13100 -6096 -12524
rect -5112 -13100 -5078 -12524
rect -4094 -13100 -4060 -12524
rect -3076 -13100 -3042 -12524
rect -2058 -13100 -2024 -12524
rect -1040 -13100 -1006 -12524
rect -22 -13100 12 -12524
rect 2582 -12624 2616 -12048
rect 3600 -12624 3634 -12048
rect 4618 -12624 4652 -12048
rect 5636 -12624 5670 -12048
rect 6654 -12624 6688 -12048
rect 7672 -12624 7706 -12048
rect 8690 -12624 8724 -12048
rect 9708 -12624 9742 -12048
rect 10726 -12624 10760 -12048
rect 11744 -12624 11778 -12048
rect 12762 -12624 12796 -12048
rect 13780 -12624 13814 -12048
rect 14798 -12624 14832 -12048
rect 15816 -12624 15850 -12048
rect 16834 -12624 16868 -12048
rect 17852 -12624 17886 -12048
rect 18870 -12624 18904 -12048
rect 19888 -12624 19922 -12048
rect 20906 -12624 20940 -12048
rect 21924 -12624 21958 -12048
rect 22942 -12624 22976 -12048
rect 2876 -12708 3340 -12674
rect 3894 -12708 4358 -12674
rect 4912 -12708 5376 -12674
rect 5930 -12708 6394 -12674
rect 6948 -12708 7412 -12674
rect 7966 -12708 8430 -12674
rect 8984 -12708 9448 -12674
rect 10002 -12708 10466 -12674
rect 11020 -12708 11484 -12674
rect 12038 -12708 12502 -12674
rect 13056 -12708 13520 -12674
rect 14074 -12708 14538 -12674
rect 15092 -12708 15556 -12674
rect 16110 -12708 16574 -12674
rect 17128 -12708 17592 -12674
rect 18146 -12708 18610 -12674
rect 19164 -12708 19628 -12674
rect 20182 -12708 20646 -12674
rect 21200 -12708 21664 -12674
rect 22218 -12708 22682 -12674
rect 2876 -12816 3340 -12782
rect 3894 -12816 4358 -12782
rect 4912 -12816 5376 -12782
rect 5930 -12816 6394 -12782
rect 6948 -12816 7412 -12782
rect 7966 -12816 8430 -12782
rect 8984 -12816 9448 -12782
rect 10002 -12816 10466 -12782
rect 11020 -12816 11484 -12782
rect 12038 -12816 12502 -12782
rect 13056 -12816 13520 -12782
rect 14074 -12816 14538 -12782
rect 15092 -12816 15556 -12782
rect 16110 -12816 16574 -12782
rect 17128 -12816 17592 -12782
rect 18146 -12816 18610 -12782
rect 19164 -12816 19628 -12782
rect 20182 -12816 20646 -12782
rect 21200 -12816 21664 -12782
rect 22218 -12816 22682 -12782
rect -8890 -13184 -8426 -13150
rect -7872 -13184 -7408 -13150
rect -8890 -13292 -8426 -13258
rect -6854 -13184 -6390 -13150
rect -7872 -13292 -7408 -13258
rect -5836 -13184 -5372 -13150
rect -6854 -13292 -6390 -13258
rect -4818 -13184 -4354 -13150
rect -5836 -13292 -5372 -13258
rect -3800 -13184 -3336 -13150
rect -4818 -13292 -4354 -13258
rect -2782 -13184 -2318 -13150
rect -3800 -13292 -3336 -13258
rect -1764 -13184 -1300 -13150
rect -2782 -13292 -2318 -13258
rect -746 -13184 -282 -13150
rect -1764 -13292 -1300 -13258
rect -746 -13292 -282 -13258
rect -9184 -13918 -9150 -13342
rect -8166 -13918 -8132 -13342
rect -7148 -13918 -7114 -13342
rect -6130 -13918 -6096 -13342
rect -5112 -13918 -5078 -13342
rect -4094 -13918 -4060 -13342
rect -3076 -13918 -3042 -13342
rect -2058 -13918 -2024 -13342
rect -1040 -13918 -1006 -13342
rect -22 -13918 12 -13342
rect 2582 -13442 2616 -12866
rect 3600 -13442 3634 -12866
rect 4618 -13442 4652 -12866
rect 5636 -13442 5670 -12866
rect 6654 -13442 6688 -12866
rect 7672 -13442 7706 -12866
rect 8690 -13442 8724 -12866
rect 9708 -13442 9742 -12866
rect 10726 -13442 10760 -12866
rect 11744 -13442 11778 -12866
rect 12762 -13442 12796 -12866
rect 13780 -13442 13814 -12866
rect 14798 -13442 14832 -12866
rect 15816 -13442 15850 -12866
rect 16834 -13442 16868 -12866
rect 17852 -13442 17886 -12866
rect 18870 -13442 18904 -12866
rect 19888 -13442 19922 -12866
rect 20906 -13442 20940 -12866
rect 21924 -13442 21958 -12866
rect 22942 -13442 22976 -12866
rect 2876 -13526 3340 -13492
rect 3894 -13526 4358 -13492
rect 4912 -13526 5376 -13492
rect 5930 -13526 6394 -13492
rect 6948 -13526 7412 -13492
rect 7966 -13526 8430 -13492
rect 8984 -13526 9448 -13492
rect 10002 -13526 10466 -13492
rect 11020 -13526 11484 -13492
rect 12038 -13526 12502 -13492
rect 13056 -13526 13520 -13492
rect 14074 -13526 14538 -13492
rect 15092 -13526 15556 -13492
rect 16110 -13526 16574 -13492
rect 17128 -13526 17592 -13492
rect 18146 -13526 18610 -13492
rect 19164 -13526 19628 -13492
rect 20182 -13526 20646 -13492
rect 21200 -13526 21664 -13492
rect 22218 -13526 22682 -13492
rect -8890 -14002 -8426 -13968
rect -7872 -14002 -7408 -13968
rect -8890 -14110 -8426 -14076
rect -6854 -14002 -6390 -13968
rect -7872 -14110 -7408 -14076
rect -5836 -14002 -5372 -13968
rect -6854 -14110 -6390 -14076
rect -4818 -14002 -4354 -13968
rect -5836 -14110 -5372 -14076
rect -3800 -14002 -3336 -13968
rect -4818 -14110 -4354 -14076
rect -2782 -14002 -2318 -13968
rect -3800 -14110 -3336 -14076
rect -1764 -14002 -1300 -13968
rect -2782 -14110 -2318 -14076
rect -746 -14002 -282 -13968
rect -1764 -14110 -1300 -14076
rect -746 -14110 -282 -14076
rect -9184 -14736 -9150 -14160
rect -8166 -14736 -8132 -14160
rect -7148 -14736 -7114 -14160
rect -6130 -14736 -6096 -14160
rect -5112 -14736 -5078 -14160
rect -4094 -14736 -4060 -14160
rect -3076 -14736 -3042 -14160
rect -2058 -14736 -2024 -14160
rect -1040 -14736 -1006 -14160
rect -22 -14736 12 -14160
rect 2876 -14194 3340 -14160
rect 3894 -14194 4358 -14160
rect 4912 -14194 5376 -14160
rect 5930 -14194 6394 -14160
rect 6948 -14194 7412 -14160
rect 7966 -14194 8430 -14160
rect 8984 -14194 9448 -14160
rect 10002 -14194 10466 -14160
rect 11020 -14194 11484 -14160
rect 12038 -14194 12502 -14160
rect 13056 -14194 13520 -14160
rect 14074 -14194 14538 -14160
rect 15092 -14194 15556 -14160
rect 16110 -14194 16574 -14160
rect 17128 -14194 17592 -14160
rect 18146 -14194 18610 -14160
rect 19164 -14194 19628 -14160
rect 20182 -14194 20646 -14160
rect 21200 -14194 21664 -14160
rect 22218 -14194 22682 -14160
rect -8890 -14820 -8426 -14786
rect -7872 -14820 -7408 -14786
rect -8890 -14928 -8426 -14894
rect -6854 -14820 -6390 -14786
rect -7872 -14928 -7408 -14894
rect -5836 -14820 -5372 -14786
rect -6854 -14928 -6390 -14894
rect -4818 -14820 -4354 -14786
rect -5836 -14928 -5372 -14894
rect -3800 -14820 -3336 -14786
rect -4818 -14928 -4354 -14894
rect -2782 -14820 -2318 -14786
rect -3800 -14928 -3336 -14894
rect -1764 -14820 -1300 -14786
rect -2782 -14928 -2318 -14894
rect -746 -14820 -282 -14786
rect -1764 -14928 -1300 -14894
rect 2582 -14820 2616 -14244
rect 3600 -14820 3634 -14244
rect 4618 -14820 4652 -14244
rect 5636 -14820 5670 -14244
rect 6654 -14820 6688 -14244
rect 7672 -14820 7706 -14244
rect 8690 -14820 8724 -14244
rect 9708 -14820 9742 -14244
rect 10726 -14820 10760 -14244
rect 11744 -14820 11778 -14244
rect 12762 -14820 12796 -14244
rect 13780 -14820 13814 -14244
rect 14798 -14820 14832 -14244
rect 15816 -14820 15850 -14244
rect 16834 -14820 16868 -14244
rect 17852 -14820 17886 -14244
rect 18870 -14820 18904 -14244
rect 19888 -14820 19922 -14244
rect 20906 -14820 20940 -14244
rect 21924 -14820 21958 -14244
rect 22942 -14820 22976 -14244
rect -746 -14928 -282 -14894
rect 2876 -14904 3340 -14870
rect 3894 -14904 4358 -14870
rect 4912 -14904 5376 -14870
rect 5930 -14904 6394 -14870
rect 6948 -14904 7412 -14870
rect 7966 -14904 8430 -14870
rect 8984 -14904 9448 -14870
rect 10002 -14904 10466 -14870
rect 11020 -14904 11484 -14870
rect 12038 -14904 12502 -14870
rect 13056 -14904 13520 -14870
rect 14074 -14904 14538 -14870
rect 15092 -14904 15556 -14870
rect 16110 -14904 16574 -14870
rect 17128 -14904 17592 -14870
rect 18146 -14904 18610 -14870
rect 19164 -14904 19628 -14870
rect 20182 -14904 20646 -14870
rect 21200 -14904 21664 -14870
rect 22218 -14904 22682 -14870
rect -9184 -15554 -9150 -14978
rect -8166 -15554 -8132 -14978
rect -7148 -15554 -7114 -14978
rect -6130 -15554 -6096 -14978
rect -5112 -15554 -5078 -14978
rect -4094 -15554 -4060 -14978
rect -3076 -15554 -3042 -14978
rect -2058 -15554 -2024 -14978
rect -1040 -15554 -1006 -14978
rect -22 -15554 12 -14978
rect 2876 -15426 3340 -15392
rect 3894 -15426 4358 -15392
rect 4912 -15426 5376 -15392
rect 5930 -15426 6394 -15392
rect 6948 -15426 7412 -15392
rect 7966 -15426 8430 -15392
rect 8984 -15426 9448 -15392
rect 10002 -15426 10466 -15392
rect 11020 -15426 11484 -15392
rect 12038 -15426 12502 -15392
rect 13056 -15426 13520 -15392
rect 14074 -15426 14538 -15392
rect 15092 -15426 15556 -15392
rect 16110 -15426 16574 -15392
rect 17128 -15426 17592 -15392
rect 18146 -15426 18610 -15392
rect 19164 -15426 19628 -15392
rect 20182 -15426 20646 -15392
rect 21200 -15426 21664 -15392
rect 22218 -15426 22682 -15392
rect -8890 -15638 -8426 -15604
rect -7872 -15638 -7408 -15604
rect -8890 -15746 -8426 -15712
rect -6854 -15638 -6390 -15604
rect -7872 -15746 -7408 -15712
rect -5836 -15638 -5372 -15604
rect -6854 -15746 -6390 -15712
rect -4818 -15638 -4354 -15604
rect -5836 -15746 -5372 -15712
rect -3800 -15638 -3336 -15604
rect -4818 -15746 -4354 -15712
rect -2782 -15638 -2318 -15604
rect -3800 -15746 -3336 -15712
rect -1764 -15638 -1300 -15604
rect -2782 -15746 -2318 -15712
rect -746 -15638 -282 -15604
rect -1764 -15746 -1300 -15712
rect -746 -15746 -282 -15712
rect -9184 -16372 -9150 -15796
rect -8166 -16372 -8132 -15796
rect -7148 -16372 -7114 -15796
rect -6130 -16372 -6096 -15796
rect -5112 -16372 -5078 -15796
rect -4094 -16372 -4060 -15796
rect -3076 -16372 -3042 -15796
rect -2058 -16372 -2024 -15796
rect -1040 -16372 -1006 -15796
rect -22 -16372 12 -15796
rect 2582 -16052 2616 -15476
rect 3600 -16052 3634 -15476
rect 4618 -16052 4652 -15476
rect 5636 -16052 5670 -15476
rect 6654 -16052 6688 -15476
rect 7672 -16052 7706 -15476
rect 8690 -16052 8724 -15476
rect 9708 -16052 9742 -15476
rect 10726 -16052 10760 -15476
rect 11744 -16052 11778 -15476
rect 12762 -16052 12796 -15476
rect 13780 -16052 13814 -15476
rect 14798 -16052 14832 -15476
rect 15816 -16052 15850 -15476
rect 16834 -16052 16868 -15476
rect 17852 -16052 17886 -15476
rect 18870 -16052 18904 -15476
rect 19888 -16052 19922 -15476
rect 20906 -16052 20940 -15476
rect 21924 -16052 21958 -15476
rect 22942 -16052 22976 -15476
rect 2876 -16136 3340 -16102
rect 3894 -16136 4358 -16102
rect 4912 -16136 5376 -16102
rect 5930 -16136 6394 -16102
rect 6948 -16136 7412 -16102
rect 7966 -16136 8430 -16102
rect 8984 -16136 9448 -16102
rect 10002 -16136 10466 -16102
rect 11020 -16136 11484 -16102
rect 12038 -16136 12502 -16102
rect 13056 -16136 13520 -16102
rect 14074 -16136 14538 -16102
rect 15092 -16136 15556 -16102
rect 16110 -16136 16574 -16102
rect 17128 -16136 17592 -16102
rect 18146 -16136 18610 -16102
rect 19164 -16136 19628 -16102
rect 20182 -16136 20646 -16102
rect 21200 -16136 21664 -16102
rect 22218 -16136 22682 -16102
rect -8890 -16456 -8426 -16422
rect -7872 -16456 -7408 -16422
rect -8890 -16564 -8426 -16530
rect -6854 -16456 -6390 -16422
rect -7872 -16564 -7408 -16530
rect -5836 -16456 -5372 -16422
rect -6854 -16564 -6390 -16530
rect -4818 -16456 -4354 -16422
rect -5836 -16564 -5372 -16530
rect -3800 -16456 -3336 -16422
rect -4818 -16564 -4354 -16530
rect -2782 -16456 -2318 -16422
rect -3800 -16564 -3336 -16530
rect -1764 -16456 -1300 -16422
rect -2782 -16564 -2318 -16530
rect -746 -16456 -282 -16422
rect -1764 -16564 -1300 -16530
rect -746 -16564 -282 -16530
rect -9184 -17190 -9150 -16614
rect -8166 -17190 -8132 -16614
rect -7148 -17190 -7114 -16614
rect -6130 -17190 -6096 -16614
rect -5112 -17190 -5078 -16614
rect -4094 -17190 -4060 -16614
rect -3076 -17190 -3042 -16614
rect -2058 -17190 -2024 -16614
rect -1040 -17190 -1006 -16614
rect -22 -17190 12 -16614
rect 2874 -16660 3338 -16626
rect 3892 -16660 4356 -16626
rect 4910 -16660 5374 -16626
rect 5928 -16660 6392 -16626
rect 6946 -16660 7410 -16626
rect 7964 -16660 8428 -16626
rect 8982 -16660 9446 -16626
rect 10000 -16660 10464 -16626
rect 11018 -16660 11482 -16626
rect 12036 -16660 12500 -16626
rect 13054 -16660 13518 -16626
rect 14072 -16660 14536 -16626
rect 15090 -16660 15554 -16626
rect 16108 -16660 16572 -16626
rect 17126 -16660 17590 -16626
rect 18144 -16660 18608 -16626
rect 19162 -16660 19626 -16626
rect 20180 -16660 20644 -16626
rect 21198 -16660 21662 -16626
rect 22216 -16660 22680 -16626
rect -8890 -17274 -8426 -17240
rect -7872 -17274 -7408 -17240
rect -8890 -17382 -8426 -17348
rect -6854 -17274 -6390 -17240
rect -7872 -17382 -7408 -17348
rect -5836 -17274 -5372 -17240
rect -6854 -17382 -6390 -17348
rect -4818 -17274 -4354 -17240
rect -5836 -17382 -5372 -17348
rect -3800 -17274 -3336 -17240
rect -4818 -17382 -4354 -17348
rect -2782 -17274 -2318 -17240
rect -3800 -17382 -3336 -17348
rect -1764 -17274 -1300 -17240
rect -2782 -17382 -2318 -17348
rect -746 -17274 -282 -17240
rect -1764 -17382 -1300 -17348
rect 2580 -17286 2614 -16710
rect 3598 -17286 3632 -16710
rect 4616 -17286 4650 -16710
rect 5634 -17286 5668 -16710
rect 6652 -17286 6686 -16710
rect 7670 -17286 7704 -16710
rect 8688 -17286 8722 -16710
rect 9706 -17286 9740 -16710
rect 10724 -17286 10758 -16710
rect 11742 -17286 11776 -16710
rect 12760 -17286 12794 -16710
rect 13778 -17286 13812 -16710
rect 14796 -17286 14830 -16710
rect 15814 -17286 15848 -16710
rect 16832 -17286 16866 -16710
rect 17850 -17286 17884 -16710
rect 18868 -17286 18902 -16710
rect 19886 -17286 19920 -16710
rect 20904 -17286 20938 -16710
rect 21922 -17286 21956 -16710
rect 22940 -17286 22974 -16710
rect -746 -17382 -282 -17348
rect 2874 -17370 3338 -17336
rect 3892 -17370 4356 -17336
rect 4910 -17370 5374 -17336
rect 5928 -17370 6392 -17336
rect 6946 -17370 7410 -17336
rect 7964 -17370 8428 -17336
rect 8982 -17370 9446 -17336
rect 10000 -17370 10464 -17336
rect 11018 -17370 11482 -17336
rect 12036 -17370 12500 -17336
rect 13054 -17370 13518 -17336
rect 14072 -17370 14536 -17336
rect 15090 -17370 15554 -17336
rect 16108 -17370 16572 -17336
rect 17126 -17370 17590 -17336
rect 18144 -17370 18608 -17336
rect 19162 -17370 19626 -17336
rect 20180 -17370 20644 -17336
rect 21198 -17370 21662 -17336
rect 22216 -17370 22680 -17336
rect -9184 -18008 -9150 -17432
rect -8166 -18008 -8132 -17432
rect -7148 -18008 -7114 -17432
rect -6130 -18008 -6096 -17432
rect -5112 -18008 -5078 -17432
rect -4094 -18008 -4060 -17432
rect -3076 -18008 -3042 -17432
rect -2058 -18008 -2024 -17432
rect -1040 -18008 -1006 -17432
rect -22 -18008 12 -17432
rect 2874 -17894 3338 -17860
rect 3892 -17894 4356 -17860
rect 4910 -17894 5374 -17860
rect 5928 -17894 6392 -17860
rect 6946 -17894 7410 -17860
rect 7964 -17894 8428 -17860
rect 8982 -17894 9446 -17860
rect 10000 -17894 10464 -17860
rect 11018 -17894 11482 -17860
rect 12036 -17894 12500 -17860
rect 13054 -17894 13518 -17860
rect 14072 -17894 14536 -17860
rect 15090 -17894 15554 -17860
rect 16108 -17894 16572 -17860
rect 17126 -17894 17590 -17860
rect 18144 -17894 18608 -17860
rect 19162 -17894 19626 -17860
rect 20180 -17894 20644 -17860
rect 21198 -17894 21662 -17860
rect 22216 -17894 22680 -17860
rect -8890 -18092 -8426 -18058
rect -7872 -18092 -7408 -18058
rect -8890 -18200 -8426 -18166
rect -6854 -18092 -6390 -18058
rect -7872 -18200 -7408 -18166
rect -5836 -18092 -5372 -18058
rect -6854 -18200 -6390 -18166
rect -4818 -18092 -4354 -18058
rect -5836 -18200 -5372 -18166
rect -3800 -18092 -3336 -18058
rect -4818 -18200 -4354 -18166
rect -2782 -18092 -2318 -18058
rect -3800 -18200 -3336 -18166
rect -1764 -18092 -1300 -18058
rect -2782 -18200 -2318 -18166
rect -746 -18092 -282 -18058
rect -1764 -18200 -1300 -18166
rect -746 -18200 -282 -18166
rect -9184 -18826 -9150 -18250
rect -8166 -18826 -8132 -18250
rect -7148 -18826 -7114 -18250
rect -6130 -18826 -6096 -18250
rect -5112 -18826 -5078 -18250
rect -4094 -18826 -4060 -18250
rect -3076 -18826 -3042 -18250
rect -2058 -18826 -2024 -18250
rect -1040 -18826 -1006 -18250
rect -22 -18826 12 -18250
rect 2580 -18520 2614 -17944
rect 3598 -18520 3632 -17944
rect 4616 -18520 4650 -17944
rect 5634 -18520 5668 -17944
rect 6652 -18520 6686 -17944
rect 7670 -18520 7704 -17944
rect 8688 -18520 8722 -17944
rect 9706 -18520 9740 -17944
rect 10724 -18520 10758 -17944
rect 11742 -18520 11776 -17944
rect 12760 -18520 12794 -17944
rect 13778 -18520 13812 -17944
rect 14796 -18520 14830 -17944
rect 15814 -18520 15848 -17944
rect 16832 -18520 16866 -17944
rect 17850 -18520 17884 -17944
rect 18868 -18520 18902 -17944
rect 19886 -18520 19920 -17944
rect 20904 -18520 20938 -17944
rect 21922 -18520 21956 -17944
rect 22940 -18520 22974 -17944
rect 2874 -18604 3338 -18570
rect 3892 -18604 4356 -18570
rect 4910 -18604 5374 -18570
rect 5928 -18604 6392 -18570
rect 6946 -18604 7410 -18570
rect 7964 -18604 8428 -18570
rect 8982 -18604 9446 -18570
rect 10000 -18604 10464 -18570
rect 11018 -18604 11482 -18570
rect 12036 -18604 12500 -18570
rect 13054 -18604 13518 -18570
rect 14072 -18604 14536 -18570
rect 15090 -18604 15554 -18570
rect 16108 -18604 16572 -18570
rect 17126 -18604 17590 -18570
rect 18144 -18604 18608 -18570
rect 19162 -18604 19626 -18570
rect 20180 -18604 20644 -18570
rect 21198 -18604 21662 -18570
rect 22216 -18604 22680 -18570
rect -8890 -18910 -8426 -18876
rect -7872 -18910 -7408 -18876
rect -6854 -18910 -6390 -18876
rect -5836 -18910 -5372 -18876
rect -4818 -18910 -4354 -18876
rect -3800 -18910 -3336 -18876
rect -2782 -18910 -2318 -18876
rect -1764 -18910 -1300 -18876
rect -746 -18910 -282 -18876
rect 2874 -19126 3338 -19092
rect 3892 -19126 4356 -19092
rect 4910 -19126 5374 -19092
rect 5928 -19126 6392 -19092
rect 6946 -19126 7410 -19092
rect 7964 -19126 8428 -19092
rect 8982 -19126 9446 -19092
rect 10000 -19126 10464 -19092
rect 11018 -19126 11482 -19092
rect 12036 -19126 12500 -19092
rect 13054 -19126 13518 -19092
rect 14072 -19126 14536 -19092
rect 15090 -19126 15554 -19092
rect 16108 -19126 16572 -19092
rect 17126 -19126 17590 -19092
rect 18144 -19126 18608 -19092
rect 19162 -19126 19626 -19092
rect 20180 -19126 20644 -19092
rect 21198 -19126 21662 -19092
rect 22216 -19126 22680 -19092
rect 2580 -19752 2614 -19176
rect 3598 -19752 3632 -19176
rect 4616 -19752 4650 -19176
rect 5634 -19752 5668 -19176
rect 6652 -19752 6686 -19176
rect 7670 -19752 7704 -19176
rect 8688 -19752 8722 -19176
rect 9706 -19752 9740 -19176
rect 10724 -19752 10758 -19176
rect 11742 -19752 11776 -19176
rect 12760 -19752 12794 -19176
rect 13778 -19752 13812 -19176
rect 14796 -19752 14830 -19176
rect 15814 -19752 15848 -19176
rect 16832 -19752 16866 -19176
rect 17850 -19752 17884 -19176
rect 18868 -19752 18902 -19176
rect 19886 -19752 19920 -19176
rect 20904 -19752 20938 -19176
rect 21922 -19752 21956 -19176
rect 22940 -19752 22974 -19176
rect 2874 -19836 3338 -19802
rect 3892 -19836 4356 -19802
rect 4910 -19836 5374 -19802
rect 5928 -19836 6392 -19802
rect 6946 -19836 7410 -19802
rect 7964 -19836 8428 -19802
rect 8982 -19836 9446 -19802
rect 10000 -19836 10464 -19802
rect 11018 -19836 11482 -19802
rect 12036 -19836 12500 -19802
rect 13054 -19836 13518 -19802
rect 14072 -19836 14536 -19802
rect 15090 -19836 15554 -19802
rect 16108 -19836 16572 -19802
rect 17126 -19836 17590 -19802
rect 18144 -19836 18608 -19802
rect 19162 -19836 19626 -19802
rect 20180 -19836 20644 -19802
rect 21198 -19836 21662 -19802
rect 22216 -19836 22680 -19802
rect -10214 -20224 -9750 -20190
rect -9196 -20224 -8732 -20190
rect -8178 -20224 -7714 -20190
rect -7160 -20224 -6696 -20190
rect -6142 -20224 -5678 -20190
rect -5124 -20224 -4660 -20190
rect -4106 -20224 -3642 -20190
rect -3088 -20224 -2624 -20190
rect -2070 -20224 -1606 -20190
rect -1052 -20224 -588 -20190
rect -34 -20224 430 -20190
rect -10508 -20850 -10474 -20274
rect -9490 -20850 -9456 -20274
rect -8472 -20850 -8438 -20274
rect -7454 -20850 -7420 -20274
rect -6436 -20850 -6402 -20274
rect -5418 -20850 -5384 -20274
rect -4400 -20850 -4366 -20274
rect -3382 -20850 -3348 -20274
rect -2364 -20850 -2330 -20274
rect -1346 -20850 -1312 -20274
rect -328 -20850 -294 -20274
rect 690 -20850 724 -20274
rect 2874 -20360 3338 -20326
rect 3892 -20360 4356 -20326
rect 4910 -20360 5374 -20326
rect 5928 -20360 6392 -20326
rect 6946 -20360 7410 -20326
rect 7964 -20360 8428 -20326
rect 8982 -20360 9446 -20326
rect 10000 -20360 10464 -20326
rect 11018 -20360 11482 -20326
rect 12036 -20360 12500 -20326
rect 13054 -20360 13518 -20326
rect 14072 -20360 14536 -20326
rect 15090 -20360 15554 -20326
rect 16108 -20360 16572 -20326
rect 17126 -20360 17590 -20326
rect 18144 -20360 18608 -20326
rect 19162 -20360 19626 -20326
rect 20180 -20360 20644 -20326
rect 21198 -20360 21662 -20326
rect 22216 -20360 22680 -20326
rect -10214 -20934 -9750 -20900
rect -9196 -20934 -8732 -20900
rect -8178 -20934 -7714 -20900
rect -7160 -20934 -6696 -20900
rect -6142 -20934 -5678 -20900
rect -5124 -20934 -4660 -20900
rect -4106 -20934 -3642 -20900
rect -3088 -20934 -2624 -20900
rect -2070 -20934 -1606 -20900
rect -1052 -20934 -588 -20900
rect -34 -20934 430 -20900
rect 2580 -20986 2614 -20410
rect 3598 -20986 3632 -20410
rect 4616 -20986 4650 -20410
rect 5634 -20986 5668 -20410
rect 6652 -20986 6686 -20410
rect 7670 -20986 7704 -20410
rect 8688 -20986 8722 -20410
rect 9706 -20986 9740 -20410
rect 10724 -20986 10758 -20410
rect 11742 -20986 11776 -20410
rect 12760 -20986 12794 -20410
rect 13778 -20986 13812 -20410
rect 14796 -20986 14830 -20410
rect 15814 -20986 15848 -20410
rect 16832 -20986 16866 -20410
rect 17850 -20986 17884 -20410
rect 18868 -20986 18902 -20410
rect 19886 -20986 19920 -20410
rect 20904 -20986 20938 -20410
rect 21922 -20986 21956 -20410
rect 22940 -20986 22974 -20410
rect 2874 -21070 3338 -21036
rect 3892 -21070 4356 -21036
rect 4910 -21070 5374 -21036
rect 5928 -21070 6392 -21036
rect 6946 -21070 7410 -21036
rect 7964 -21070 8428 -21036
rect 8982 -21070 9446 -21036
rect 10000 -21070 10464 -21036
rect 11018 -21070 11482 -21036
rect 12036 -21070 12500 -21036
rect 13054 -21070 13518 -21036
rect 14072 -21070 14536 -21036
rect 15090 -21070 15554 -21036
rect 16108 -21070 16572 -21036
rect 17126 -21070 17590 -21036
rect 18144 -21070 18608 -21036
rect 19162 -21070 19626 -21036
rect 20180 -21070 20644 -21036
rect 21198 -21070 21662 -21036
rect 22216 -21070 22680 -21036
rect -10214 -21336 -9750 -21302
rect -9196 -21336 -8732 -21302
rect -8178 -21336 -7714 -21302
rect -7160 -21336 -6696 -21302
rect -6142 -21336 -5678 -21302
rect -5124 -21336 -4660 -21302
rect -4106 -21336 -3642 -21302
rect -3088 -21336 -2624 -21302
rect -2070 -21336 -1606 -21302
rect -1052 -21336 -588 -21302
rect -34 -21336 430 -21302
rect -10508 -21962 -10474 -21386
rect -9490 -21962 -9456 -21386
rect -8472 -21962 -8438 -21386
rect -7454 -21962 -7420 -21386
rect -6436 -21962 -6402 -21386
rect -5418 -21962 -5384 -21386
rect -4400 -21962 -4366 -21386
rect -3382 -21962 -3348 -21386
rect -2364 -21962 -2330 -21386
rect -1346 -21962 -1312 -21386
rect -328 -21962 -294 -21386
rect 690 -21962 724 -21386
rect 2874 -21594 3338 -21560
rect 3892 -21594 4356 -21560
rect 4910 -21594 5374 -21560
rect 5928 -21594 6392 -21560
rect 6946 -21594 7410 -21560
rect 7964 -21594 8428 -21560
rect 8982 -21594 9446 -21560
rect 10000 -21594 10464 -21560
rect 11018 -21594 11482 -21560
rect 12036 -21594 12500 -21560
rect 13054 -21594 13518 -21560
rect 14072 -21594 14536 -21560
rect 15090 -21594 15554 -21560
rect 16108 -21594 16572 -21560
rect 17126 -21594 17590 -21560
rect 18144 -21594 18608 -21560
rect 19162 -21594 19626 -21560
rect 20180 -21594 20644 -21560
rect 21198 -21594 21662 -21560
rect 22216 -21594 22680 -21560
rect -10214 -22046 -9750 -22012
rect -9196 -22046 -8732 -22012
rect -8178 -22046 -7714 -22012
rect -7160 -22046 -6696 -22012
rect -6142 -22046 -5678 -22012
rect -5124 -22046 -4660 -22012
rect -4106 -22046 -3642 -22012
rect -3088 -22046 -2624 -22012
rect -2070 -22046 -1606 -22012
rect -1052 -22046 -588 -22012
rect -34 -22046 430 -22012
rect 2580 -22220 2614 -21644
rect 3598 -22220 3632 -21644
rect 4616 -22220 4650 -21644
rect 5634 -22220 5668 -21644
rect 6652 -22220 6686 -21644
rect 7670 -22220 7704 -21644
rect 8688 -22220 8722 -21644
rect 9706 -22220 9740 -21644
rect 10724 -22220 10758 -21644
rect 11742 -22220 11776 -21644
rect 12760 -22220 12794 -21644
rect 13778 -22220 13812 -21644
rect 14796 -22220 14830 -21644
rect 15814 -22220 15848 -21644
rect 16832 -22220 16866 -21644
rect 17850 -22220 17884 -21644
rect 18868 -22220 18902 -21644
rect 19886 -22220 19920 -21644
rect 20904 -22220 20938 -21644
rect 21922 -22220 21956 -21644
rect 22940 -22220 22974 -21644
rect 2874 -22304 3338 -22270
rect 3892 -22304 4356 -22270
rect 4910 -22304 5374 -22270
rect 5928 -22304 6392 -22270
rect 6946 -22304 7410 -22270
rect 7964 -22304 8428 -22270
rect 8982 -22304 9446 -22270
rect 10000 -22304 10464 -22270
rect 11018 -22304 11482 -22270
rect 12036 -22304 12500 -22270
rect 13054 -22304 13518 -22270
rect 14072 -22304 14536 -22270
rect 15090 -22304 15554 -22270
rect 16108 -22304 16572 -22270
rect 17126 -22304 17590 -22270
rect 18144 -22304 18608 -22270
rect 19162 -22304 19626 -22270
rect 20180 -22304 20644 -22270
rect 21198 -22304 21662 -22270
rect 22216 -22304 22680 -22270
rect -10214 -22448 -9750 -22414
rect -9196 -22448 -8732 -22414
rect -8178 -22448 -7714 -22414
rect -7160 -22448 -6696 -22414
rect -6142 -22448 -5678 -22414
rect -5124 -22448 -4660 -22414
rect -4106 -22448 -3642 -22414
rect -3088 -22448 -2624 -22414
rect -2070 -22448 -1606 -22414
rect -1052 -22448 -588 -22414
rect -34 -22448 430 -22414
rect -10508 -23074 -10474 -22498
rect -9490 -23074 -9456 -22498
rect -8472 -23074 -8438 -22498
rect -7454 -23074 -7420 -22498
rect -6436 -23074 -6402 -22498
rect -5418 -23074 -5384 -22498
rect -4400 -23074 -4366 -22498
rect -3382 -23074 -3348 -22498
rect -2364 -23074 -2330 -22498
rect -1346 -23074 -1312 -22498
rect -328 -23074 -294 -22498
rect 690 -23074 724 -22498
rect 2874 -22826 3338 -22792
rect 3892 -22826 4356 -22792
rect 4910 -22826 5374 -22792
rect 5928 -22826 6392 -22792
rect 6946 -22826 7410 -22792
rect 7964 -22826 8428 -22792
rect 8982 -22826 9446 -22792
rect 10000 -22826 10464 -22792
rect 11018 -22826 11482 -22792
rect 12036 -22826 12500 -22792
rect 13054 -22826 13518 -22792
rect 14072 -22826 14536 -22792
rect 15090 -22826 15554 -22792
rect 16108 -22826 16572 -22792
rect 17126 -22826 17590 -22792
rect 18144 -22826 18608 -22792
rect 19162 -22826 19626 -22792
rect 20180 -22826 20644 -22792
rect 21198 -22826 21662 -22792
rect 22216 -22826 22680 -22792
rect -10214 -23158 -9750 -23124
rect -9196 -23158 -8732 -23124
rect -8178 -23158 -7714 -23124
rect -7160 -23158 -6696 -23124
rect -6142 -23158 -5678 -23124
rect -5124 -23158 -4660 -23124
rect -4106 -23158 -3642 -23124
rect -3088 -23158 -2624 -23124
rect -2070 -23158 -1606 -23124
rect -1052 -23158 -588 -23124
rect -34 -23158 430 -23124
rect 2580 -23452 2614 -22876
rect 3598 -23452 3632 -22876
rect 4616 -23452 4650 -22876
rect 5634 -23452 5668 -22876
rect 6652 -23452 6686 -22876
rect 7670 -23452 7704 -22876
rect 8688 -23452 8722 -22876
rect 9706 -23452 9740 -22876
rect 10724 -23452 10758 -22876
rect 11742 -23452 11776 -22876
rect 12760 -23452 12794 -22876
rect 13778 -23452 13812 -22876
rect 14796 -23452 14830 -22876
rect 15814 -23452 15848 -22876
rect 16832 -23452 16866 -22876
rect 17850 -23452 17884 -22876
rect 18868 -23452 18902 -22876
rect 19886 -23452 19920 -22876
rect 20904 -23452 20938 -22876
rect 21922 -23452 21956 -22876
rect 22940 -23452 22974 -22876
rect -10214 -23560 -9750 -23526
rect -9196 -23560 -8732 -23526
rect -8178 -23560 -7714 -23526
rect -7160 -23560 -6696 -23526
rect -6142 -23560 -5678 -23526
rect -5124 -23560 -4660 -23526
rect -4106 -23560 -3642 -23526
rect -3088 -23560 -2624 -23526
rect -2070 -23560 -1606 -23526
rect -1052 -23560 -588 -23526
rect -34 -23560 430 -23526
rect 2874 -23536 3338 -23502
rect 3892 -23536 4356 -23502
rect 4910 -23536 5374 -23502
rect 5928 -23536 6392 -23502
rect 6946 -23536 7410 -23502
rect 7964 -23536 8428 -23502
rect 8982 -23536 9446 -23502
rect 10000 -23536 10464 -23502
rect 11018 -23536 11482 -23502
rect 12036 -23536 12500 -23502
rect 13054 -23536 13518 -23502
rect 14072 -23536 14536 -23502
rect 15090 -23536 15554 -23502
rect 16108 -23536 16572 -23502
rect 17126 -23536 17590 -23502
rect 18144 -23536 18608 -23502
rect 19162 -23536 19626 -23502
rect 20180 -23536 20644 -23502
rect 21198 -23536 21662 -23502
rect 22216 -23536 22680 -23502
rect -10508 -24186 -10474 -23610
rect -9490 -24186 -9456 -23610
rect -8472 -24186 -8438 -23610
rect -7454 -24186 -7420 -23610
rect -6436 -24186 -6402 -23610
rect -5418 -24186 -5384 -23610
rect -4400 -24186 -4366 -23610
rect -3382 -24186 -3348 -23610
rect -2364 -24186 -2330 -23610
rect -1346 -24186 -1312 -23610
rect -328 -24186 -294 -23610
rect 690 -24186 724 -23610
rect 2874 -24060 3338 -24026
rect 3892 -24060 4356 -24026
rect 4910 -24060 5374 -24026
rect 5928 -24060 6392 -24026
rect 6946 -24060 7410 -24026
rect 7964 -24060 8428 -24026
rect 8982 -24060 9446 -24026
rect 10000 -24060 10464 -24026
rect 11018 -24060 11482 -24026
rect 12036 -24060 12500 -24026
rect 13054 -24060 13518 -24026
rect 14072 -24060 14536 -24026
rect 15090 -24060 15554 -24026
rect 16108 -24060 16572 -24026
rect 17126 -24060 17590 -24026
rect 18144 -24060 18608 -24026
rect 19162 -24060 19626 -24026
rect 20180 -24060 20644 -24026
rect 21198 -24060 21662 -24026
rect 22216 -24060 22680 -24026
rect -10214 -24270 -9750 -24236
rect -9196 -24270 -8732 -24236
rect -8178 -24270 -7714 -24236
rect -7160 -24270 -6696 -24236
rect -6142 -24270 -5678 -24236
rect -5124 -24270 -4660 -24236
rect -4106 -24270 -3642 -24236
rect -3088 -24270 -2624 -24236
rect -2070 -24270 -1606 -24236
rect -1052 -24270 -588 -24236
rect -34 -24270 430 -24236
rect 2580 -24686 2614 -24110
rect 3598 -24686 3632 -24110
rect 4616 -24686 4650 -24110
rect 5634 -24686 5668 -24110
rect 6652 -24686 6686 -24110
rect 7670 -24686 7704 -24110
rect 8688 -24686 8722 -24110
rect 9706 -24686 9740 -24110
rect 10724 -24686 10758 -24110
rect 11742 -24686 11776 -24110
rect 12760 -24686 12794 -24110
rect 13778 -24686 13812 -24110
rect 14796 -24686 14830 -24110
rect 15814 -24686 15848 -24110
rect 16832 -24686 16866 -24110
rect 17850 -24686 17884 -24110
rect 18868 -24686 18902 -24110
rect 19886 -24686 19920 -24110
rect 20904 -24686 20938 -24110
rect 21922 -24686 21956 -24110
rect 22940 -24686 22974 -24110
rect 2874 -24770 3338 -24736
rect 3892 -24770 4356 -24736
rect 4910 -24770 5374 -24736
rect 5928 -24770 6392 -24736
rect 6946 -24770 7410 -24736
rect 7964 -24770 8428 -24736
rect 8982 -24770 9446 -24736
rect 10000 -24770 10464 -24736
rect 11018 -24770 11482 -24736
rect 12036 -24770 12500 -24736
rect 13054 -24770 13518 -24736
rect 14072 -24770 14536 -24736
rect 15090 -24770 15554 -24736
rect 16108 -24770 16572 -24736
rect 17126 -24770 17590 -24736
rect 18144 -24770 18608 -24736
rect 19162 -24770 19626 -24736
rect 20180 -24770 20644 -24736
rect 21198 -24770 21662 -24736
rect 22216 -24770 22680 -24736
rect -9756 -25102 -9292 -25068
rect -8738 -25102 -8274 -25068
rect -7720 -25102 -7256 -25068
rect -6702 -25102 -6238 -25068
rect -5684 -25102 -5220 -25068
rect -4666 -25102 -4202 -25068
rect -3648 -25102 -3184 -25068
rect -2630 -25102 -2166 -25068
rect -1612 -25102 -1148 -25068
rect -594 -25102 -130 -25068
rect -10050 -25728 -10016 -25152
rect -9032 -25728 -8998 -25152
rect -8014 -25728 -7980 -25152
rect -6996 -25728 -6962 -25152
rect -5978 -25728 -5944 -25152
rect -4960 -25728 -4926 -25152
rect -3942 -25728 -3908 -25152
rect -2924 -25728 -2890 -25152
rect -1906 -25728 -1872 -25152
rect -888 -25728 -854 -25152
rect 130 -25728 164 -25152
rect 2874 -25292 3338 -25258
rect 3892 -25292 4356 -25258
rect 4910 -25292 5374 -25258
rect 5928 -25292 6392 -25258
rect 6946 -25292 7410 -25258
rect 7964 -25292 8428 -25258
rect 8982 -25292 9446 -25258
rect 10000 -25292 10464 -25258
rect 11018 -25292 11482 -25258
rect 12036 -25292 12500 -25258
rect 13054 -25292 13518 -25258
rect 14072 -25292 14536 -25258
rect 15090 -25292 15554 -25258
rect 16108 -25292 16572 -25258
rect 17126 -25292 17590 -25258
rect 18144 -25292 18608 -25258
rect 19162 -25292 19626 -25258
rect 20180 -25292 20644 -25258
rect 21198 -25292 21662 -25258
rect 22216 -25292 22680 -25258
rect -9756 -25812 -9292 -25778
rect -8738 -25812 -8274 -25778
rect -7720 -25812 -7256 -25778
rect -6702 -25812 -6238 -25778
rect -5684 -25812 -5220 -25778
rect -4666 -25812 -4202 -25778
rect -3648 -25812 -3184 -25778
rect -2630 -25812 -2166 -25778
rect -1612 -25812 -1148 -25778
rect -594 -25812 -130 -25778
rect 2580 -25918 2614 -25342
rect 3598 -25918 3632 -25342
rect 4616 -25918 4650 -25342
rect 5634 -25918 5668 -25342
rect 6652 -25918 6686 -25342
rect 7670 -25918 7704 -25342
rect 8688 -25918 8722 -25342
rect 9706 -25918 9740 -25342
rect 10724 -25918 10758 -25342
rect 11742 -25918 11776 -25342
rect 12760 -25918 12794 -25342
rect 13778 -25918 13812 -25342
rect 14796 -25918 14830 -25342
rect 15814 -25918 15848 -25342
rect 16832 -25918 16866 -25342
rect 17850 -25918 17884 -25342
rect 18868 -25918 18902 -25342
rect 19886 -25918 19920 -25342
rect 20904 -25918 20938 -25342
rect 21922 -25918 21956 -25342
rect 22940 -25918 22974 -25342
rect 2874 -26002 3338 -25968
rect 3892 -26002 4356 -25968
rect 4910 -26002 5374 -25968
rect 5928 -26002 6392 -25968
rect 6946 -26002 7410 -25968
rect 7964 -26002 8428 -25968
rect 8982 -26002 9446 -25968
rect 10000 -26002 10464 -25968
rect 11018 -26002 11482 -25968
rect 12036 -26002 12500 -25968
rect 13054 -26002 13518 -25968
rect 14072 -26002 14536 -25968
rect 15090 -26002 15554 -25968
rect 16108 -26002 16572 -25968
rect 17126 -26002 17590 -25968
rect 18144 -26002 18608 -25968
rect 19162 -26002 19626 -25968
rect 20180 -26002 20644 -25968
rect 21198 -26002 21662 -25968
rect 22216 -26002 22680 -25968
rect 24822 -26330 24922 -12070
rect -12222 -27222 -12160 -27122
rect -12160 -27222 24760 -27122
rect 24760 -27222 24822 -27122
<< metal1 >>
rect 372 4322 24828 4328
rect 372 4222 478 4322
rect 24722 4222 24828 4322
rect 372 4216 24828 4222
rect 372 3702 484 4216
rect 1084 3916 1094 4216
rect 24106 3916 24116 4216
rect 372 -9728 378 3702
rect 478 -9728 484 3702
rect 3998 3834 20878 3866
rect 3998 3620 4061 3834
rect 20846 3620 20878 3834
rect 3998 3598 4048 3620
rect 4108 3598 4484 3620
rect 4544 3598 4922 3620
rect 4982 3598 5356 3620
rect 5416 3600 20878 3620
rect 24716 3702 24828 4216
rect 5416 3598 8352 3600
rect 8512 2124 8572 3600
rect 10548 2124 10608 3600
rect 11052 2124 11112 3600
rect 11560 2124 11620 3600
rect 12072 2124 12132 3600
rect 12586 2124 12646 3600
rect 14618 2124 14678 3600
rect 16658 2124 16718 3600
rect 17148 2124 17208 3600
rect 17668 2124 17728 3600
rect 18176 2124 18236 3600
rect 18690 2124 18750 3600
rect 20726 2124 20786 3600
rect 8512 2064 20786 2124
rect 7980 1858 7986 1918
rect 8046 1858 8052 1918
rect 6474 1642 7552 1702
rect 6474 1462 6534 1642
rect 6978 1561 7038 1642
rect 6770 1555 7258 1561
rect 6770 1521 6782 1555
rect 7246 1521 7258 1555
rect 6770 1515 7258 1521
rect 6474 1422 6488 1462
rect 6482 886 6488 1422
rect 6522 1422 6534 1462
rect 7492 1462 7552 1642
rect 7986 1561 8046 1858
rect 8512 1672 8572 2064
rect 9062 1858 9068 1918
rect 9128 1858 9134 1918
rect 10020 1858 10026 1918
rect 10086 1858 10092 1918
rect 8506 1612 8512 1672
rect 8572 1612 8578 1672
rect 7788 1555 8276 1561
rect 7788 1521 7800 1555
rect 8264 1521 8276 1555
rect 7788 1515 8276 1521
rect 7492 1436 7506 1462
rect 6522 886 6528 1422
rect 7500 922 7506 1436
rect 6482 874 6528 886
rect 7494 886 7506 922
rect 7540 1436 7552 1462
rect 8512 1462 8572 1612
rect 9068 1561 9128 1858
rect 10026 1561 10086 1858
rect 10548 1672 10608 2064
rect 10542 1612 10548 1672
rect 10608 1612 10614 1672
rect 8806 1555 9294 1561
rect 8806 1521 8818 1555
rect 9282 1521 9294 1555
rect 8806 1515 9294 1521
rect 9824 1555 10312 1561
rect 9824 1521 9836 1555
rect 10300 1521 10312 1555
rect 9824 1515 10312 1521
rect 10026 1512 10086 1515
rect 8512 1438 8524 1462
rect 7540 922 7546 1436
rect 8518 926 8524 1438
rect 7540 886 7554 922
rect 6770 827 7258 833
rect 6770 793 6782 827
rect 7246 793 7258 827
rect 6770 787 7258 793
rect 7494 740 7554 886
rect 8514 886 8524 926
rect 8558 1438 8572 1462
rect 9536 1462 9582 1474
rect 8558 926 8564 1438
rect 8558 886 8574 926
rect 9536 914 9542 1462
rect 7998 833 8058 834
rect 7788 827 8276 833
rect 7788 793 7800 827
rect 8264 793 8276 827
rect 7788 787 8276 793
rect 6324 680 6330 740
rect 6390 680 6396 740
rect 7488 680 7494 740
rect 7554 680 7560 740
rect 6194 476 6200 536
rect 6260 476 6266 536
rect 4186 -1708 4192 -1648
rect 4252 -1708 4258 -1648
rect 2014 -5024 3236 -4964
rect 2014 -6940 2074 -5024
rect 2156 -5188 2216 -5024
rect 2668 -5089 2728 -5024
rect 2452 -5095 2940 -5089
rect 2452 -5129 2464 -5095
rect 2928 -5129 2940 -5095
rect 2452 -5135 2940 -5129
rect 2156 -5238 2170 -5188
rect 2164 -5764 2170 -5238
rect 2204 -5238 2216 -5188
rect 3176 -5188 3236 -5024
rect 3470 -5095 3958 -5089
rect 3470 -5129 3482 -5095
rect 3946 -5129 3958 -5095
rect 3470 -5135 3958 -5129
rect 2204 -5764 2210 -5238
rect 3176 -5240 3188 -5188
rect 2164 -5776 2210 -5764
rect 3182 -5764 3188 -5240
rect 3222 -5240 3236 -5188
rect 4192 -5188 4252 -1708
rect 6200 -2080 6260 476
rect 6330 -1934 6390 680
rect 7488 476 7494 536
rect 7554 476 7560 536
rect 6770 419 7258 425
rect 6770 385 6782 419
rect 7246 385 7258 419
rect 6770 379 7258 385
rect 6482 326 6528 338
rect 6482 -214 6488 326
rect 6476 -250 6488 -214
rect 6522 -214 6528 326
rect 7494 326 7554 476
rect 7998 425 8058 787
rect 7788 419 8276 425
rect 7788 385 7800 419
rect 8264 385 8276 419
rect 7788 379 8276 385
rect 7998 376 8058 379
rect 7494 288 7506 326
rect 6522 -250 6536 -214
rect 7500 -220 7506 288
rect 6476 -400 6536 -250
rect 7494 -250 7506 -220
rect 7540 288 7554 326
rect 8514 326 8574 886
rect 9530 886 9542 914
rect 9576 914 9582 1462
rect 10548 1462 10608 1612
rect 11052 1561 11112 2064
rect 10842 1555 11330 1561
rect 10842 1521 10854 1555
rect 11318 1521 11330 1555
rect 10842 1515 11330 1521
rect 10548 1438 10560 1462
rect 10554 944 10560 1438
rect 9576 886 9590 914
rect 8806 827 9294 833
rect 8806 793 8818 827
rect 9282 793 9294 827
rect 8806 787 9294 793
rect 9530 636 9590 886
rect 10538 886 10560 944
rect 10594 1438 10608 1462
rect 11560 1462 11620 2064
rect 12072 1561 12132 2064
rect 12586 1674 12646 2064
rect 13084 1858 13090 1918
rect 13150 1858 13156 1918
rect 14102 1858 14108 1918
rect 14168 1858 14174 1918
rect 12580 1614 12586 1674
rect 12646 1614 12652 1674
rect 11860 1555 12348 1561
rect 11860 1521 11872 1555
rect 12336 1521 12348 1555
rect 11860 1515 12348 1521
rect 10594 944 10600 1438
rect 11560 1392 11578 1462
rect 10594 886 10602 944
rect 9824 827 10312 833
rect 9824 793 9836 827
rect 10300 793 10312 827
rect 9824 787 10312 793
rect 9524 576 9530 636
rect 9590 576 9596 636
rect 8806 419 9294 425
rect 8806 385 8818 419
rect 9282 385 9294 419
rect 8806 379 9294 385
rect 9824 419 10312 425
rect 9824 385 9836 419
rect 10300 385 10312 419
rect 9824 379 10312 385
rect 7540 -220 7546 288
rect 8514 286 8524 326
rect 7540 -250 7554 -220
rect 8518 -224 8524 286
rect 6770 -309 7258 -303
rect 6770 -343 6782 -309
rect 7246 -343 7258 -309
rect 6770 -349 7258 -343
rect 6988 -400 7048 -349
rect 7494 -400 7554 -250
rect 8510 -250 8524 -224
rect 8558 286 8574 326
rect 9536 326 9582 338
rect 8558 -224 8564 286
rect 8558 -250 8570 -224
rect 9536 -230 9542 326
rect 7980 -303 8040 -296
rect 7788 -309 8276 -303
rect 7788 -343 7800 -309
rect 8264 -343 8276 -309
rect 7788 -349 8276 -343
rect 6476 -460 7554 -400
rect 7488 -604 7548 -602
rect 6478 -664 7548 -604
rect 6478 -810 6538 -664
rect 6988 -711 7048 -664
rect 6770 -717 7258 -711
rect 6770 -751 6782 -717
rect 7246 -751 7258 -717
rect 6770 -757 7258 -751
rect 6478 -842 6488 -810
rect 6482 -1386 6488 -842
rect 6522 -842 6538 -810
rect 7488 -810 7548 -664
rect 7980 -614 8040 -349
rect 7980 -711 8040 -674
rect 8510 -396 8570 -250
rect 9528 -250 9542 -230
rect 9576 -230 9582 326
rect 10538 326 10602 886
rect 11572 886 11578 1392
rect 11612 1392 11620 1462
rect 12586 1462 12646 1614
rect 13090 1561 13150 1858
rect 14108 1561 14168 1858
rect 14618 1674 14678 2064
rect 15126 1858 15132 1918
rect 15192 1858 15198 1918
rect 16138 1858 16144 1918
rect 16204 1858 16210 1918
rect 14610 1614 14616 1674
rect 14676 1614 14682 1674
rect 12878 1555 13366 1561
rect 12878 1521 12890 1555
rect 13354 1521 13366 1555
rect 12878 1515 13366 1521
rect 13896 1555 14384 1561
rect 13896 1521 13908 1555
rect 14372 1521 14384 1555
rect 13896 1515 14384 1521
rect 12586 1422 12596 1462
rect 11612 886 11618 1392
rect 12590 940 12596 1422
rect 11572 874 11618 886
rect 12574 886 12596 940
rect 12630 1422 12646 1462
rect 13608 1462 13654 1474
rect 12630 940 12636 1422
rect 12630 886 12638 940
rect 13608 926 13614 1462
rect 10842 827 11330 833
rect 10842 793 10854 827
rect 11318 793 11330 827
rect 10842 787 11330 793
rect 11860 827 12348 833
rect 11860 793 11872 827
rect 12336 793 12348 827
rect 11860 787 12348 793
rect 11560 576 11566 636
rect 11626 576 11632 636
rect 10842 419 11330 425
rect 10842 385 10854 419
rect 11318 385 11330 419
rect 10842 379 11330 385
rect 10538 296 10560 326
rect 10554 -222 10560 296
rect 9576 -250 9588 -230
rect 9008 -303 9068 -302
rect 8806 -309 9294 -303
rect 8806 -343 8818 -309
rect 9282 -343 9294 -309
rect 8806 -349 9294 -343
rect 9008 -396 9068 -349
rect 9528 -396 9588 -250
rect 10546 -250 10560 -222
rect 10594 296 10602 326
rect 11566 326 11626 576
rect 11860 419 12348 425
rect 11860 385 11872 419
rect 12336 385 12348 419
rect 11860 379 12348 385
rect 10594 -222 10600 296
rect 11566 288 11578 326
rect 11572 -214 11578 288
rect 10594 -224 10606 -222
rect 10594 -250 10610 -224
rect 10036 -303 10096 -298
rect 9824 -309 10312 -303
rect 9824 -343 9836 -309
rect 10300 -343 10312 -309
rect 9824 -349 10312 -343
rect 10036 -396 10096 -349
rect 8510 -398 10096 -396
rect 10546 -398 10610 -250
rect 11564 -250 11578 -214
rect 11612 288 11626 326
rect 12574 326 12638 886
rect 13604 886 13614 926
rect 13648 926 13654 1462
rect 14618 1462 14678 1614
rect 15132 1561 15192 1858
rect 16144 1561 16204 1858
rect 16658 1676 16718 2064
rect 16652 1616 16658 1676
rect 16718 1616 16724 1676
rect 14914 1555 15402 1561
rect 14914 1521 14926 1555
rect 15390 1521 15402 1555
rect 14914 1515 15402 1521
rect 15932 1555 16420 1561
rect 15932 1521 15944 1555
rect 16408 1521 16420 1555
rect 15932 1515 16420 1521
rect 14618 1422 14632 1462
rect 14626 942 14632 1422
rect 13648 886 13664 926
rect 13092 833 13152 836
rect 12878 827 13366 833
rect 12878 793 12890 827
rect 13354 793 13366 827
rect 12878 787 13366 793
rect 13092 425 13152 787
rect 13604 740 13664 886
rect 14616 886 14632 942
rect 14666 1422 14678 1462
rect 15644 1462 15690 1474
rect 14666 942 14672 1422
rect 14666 886 14680 942
rect 15644 924 15650 1462
rect 14110 833 14170 842
rect 13896 827 14384 833
rect 13896 793 13908 827
rect 14372 793 14384 827
rect 13896 787 14384 793
rect 13598 680 13604 740
rect 13664 680 13670 740
rect 13594 476 13600 536
rect 13660 476 13666 536
rect 12878 419 13366 425
rect 12878 385 12890 419
rect 13354 385 13366 419
rect 12878 379 13366 385
rect 13092 378 13152 379
rect 12574 292 12596 326
rect 11612 -214 11618 288
rect 12590 -214 12596 292
rect 11612 -250 11628 -214
rect 10842 -309 11330 -303
rect 10842 -343 10854 -309
rect 11318 -343 11330 -309
rect 10842 -349 11330 -343
rect 8510 -456 10036 -398
rect 7788 -717 8276 -711
rect 7788 -751 7800 -717
rect 8264 -751 8276 -717
rect 7788 -757 8276 -751
rect 7488 -842 7506 -810
rect 6522 -1386 6528 -842
rect 7500 -1344 7506 -842
rect 6482 -1398 6528 -1386
rect 7488 -1386 7506 -1344
rect 7540 -842 7548 -810
rect 8510 -810 8570 -456
rect 10540 -458 10546 -398
rect 10606 -458 10612 -398
rect 10036 -464 10096 -458
rect 9522 -560 9528 -496
rect 9592 -560 9598 -496
rect 9012 -674 9018 -614
rect 9078 -674 9084 -614
rect 9528 -654 9592 -560
rect 9018 -711 9078 -674
rect 8806 -717 9294 -711
rect 8806 -751 8818 -717
rect 9282 -751 9294 -717
rect 8806 -757 9294 -751
rect 7540 -1344 7546 -842
rect 8510 -862 8524 -810
rect 7540 -1386 7552 -1344
rect 8518 -1350 8524 -862
rect 6770 -1445 7258 -1439
rect 6770 -1479 6782 -1445
rect 7246 -1479 7258 -1445
rect 6770 -1485 7258 -1479
rect 7488 -1594 7552 -1386
rect 8510 -1386 8524 -1350
rect 8558 -862 8570 -810
rect 9528 -810 9594 -654
rect 10024 -674 10030 -614
rect 10090 -674 10096 -614
rect 10030 -711 10090 -674
rect 9824 -717 10312 -711
rect 9824 -751 9836 -717
rect 10300 -751 10312 -717
rect 9824 -757 10312 -751
rect 10030 -758 10090 -757
rect 9528 -860 9542 -810
rect 8558 -1350 8564 -862
rect 8558 -1386 8570 -1350
rect 9536 -1362 9542 -860
rect 7788 -1445 8276 -1439
rect 7788 -1479 7800 -1445
rect 8264 -1479 8276 -1445
rect 7788 -1485 8276 -1479
rect 7044 -1654 7552 -1594
rect 6324 -1994 6330 -1934
rect 6390 -1994 6396 -1934
rect 6200 -2140 6620 -2080
rect 6560 -4952 6620 -2140
rect 6680 -4402 6686 -4342
rect 6746 -4402 6752 -4342
rect 5210 -5020 6420 -4960
rect 6554 -5012 6560 -4952
rect 6620 -5012 6626 -4952
rect 4488 -5095 4976 -5089
rect 4488 -5129 4500 -5095
rect 4964 -5129 4976 -5095
rect 4488 -5135 4976 -5129
rect 3222 -5764 3228 -5240
rect 3182 -5776 3228 -5764
rect 4192 -5764 4206 -5188
rect 4240 -5764 4252 -5188
rect 5210 -5188 5270 -5020
rect 5722 -5089 5782 -5020
rect 5506 -5095 5994 -5089
rect 5506 -5129 5518 -5095
rect 5982 -5129 5994 -5095
rect 5506 -5135 5994 -5129
rect 5210 -5236 5224 -5188
rect 2452 -5823 2940 -5817
rect 2452 -5857 2464 -5823
rect 2928 -5857 2940 -5823
rect 2452 -5863 2940 -5857
rect 3470 -5823 3958 -5817
rect 3470 -5857 3482 -5823
rect 3946 -5857 3958 -5823
rect 3470 -5863 3958 -5857
rect 3676 -5906 3736 -5863
rect 3670 -5966 3676 -5906
rect 3736 -5966 3742 -5906
rect 3778 -6078 3784 -6018
rect 3844 -6078 3850 -6018
rect 3784 -6121 3844 -6078
rect 2452 -6127 2940 -6121
rect 2452 -6161 2464 -6127
rect 2928 -6161 2940 -6127
rect 2452 -6167 2940 -6161
rect 3470 -6127 3958 -6121
rect 3470 -6161 3482 -6127
rect 3946 -6161 3958 -6127
rect 3470 -6167 3958 -6161
rect 2164 -6220 2210 -6208
rect 2164 -6738 2170 -6220
rect 2154 -6796 2170 -6738
rect 2204 -6738 2210 -6220
rect 3182 -6220 3228 -6208
rect 2204 -6796 2214 -6738
rect 3182 -6746 3188 -6220
rect 2008 -7000 2014 -6940
rect 2074 -7000 2080 -6940
rect 1888 -8028 1948 -8022
rect 2014 -8028 2074 -7000
rect 2154 -7050 2214 -6796
rect 3174 -6796 3188 -6746
rect 3222 -6746 3228 -6220
rect 4192 -6220 4252 -5764
rect 5218 -5764 5224 -5236
rect 5258 -5236 5270 -5188
rect 6228 -5188 6288 -5020
rect 6228 -5234 6242 -5188
rect 5258 -5764 5264 -5236
rect 5218 -5776 5264 -5764
rect 6236 -5764 6242 -5234
rect 6276 -5234 6288 -5188
rect 6276 -5764 6282 -5234
rect 6236 -5776 6282 -5764
rect 4488 -5823 4976 -5817
rect 4488 -5857 4500 -5823
rect 4964 -5857 4976 -5823
rect 4488 -5863 4976 -5857
rect 5506 -5823 5994 -5817
rect 5506 -5857 5518 -5823
rect 5982 -5857 5994 -5823
rect 5506 -5863 5994 -5857
rect 4568 -6018 4628 -5863
rect 4692 -5966 4698 -5906
rect 4758 -5966 4764 -5906
rect 4562 -6078 4568 -6018
rect 4628 -6078 4634 -6018
rect 4698 -6121 4758 -5966
rect 4488 -6127 4976 -6121
rect 4488 -6161 4500 -6127
rect 4964 -6161 4976 -6127
rect 4488 -6167 4976 -6161
rect 5506 -6127 5994 -6121
rect 5506 -6161 5518 -6127
rect 5982 -6161 5994 -6127
rect 5506 -6167 5994 -6161
rect 3222 -6796 3234 -6746
rect 2452 -6855 2940 -6849
rect 2452 -6889 2464 -6855
rect 2928 -6889 2940 -6855
rect 2452 -6895 2940 -6889
rect 2656 -7050 2716 -6895
rect 3174 -7050 3234 -6796
rect 4192 -6796 4206 -6220
rect 4240 -6796 4252 -6220
rect 5218 -6220 5264 -6208
rect 5218 -6710 5224 -6220
rect 3470 -6855 3958 -6849
rect 3470 -6889 3482 -6855
rect 3946 -6889 3958 -6855
rect 3470 -6895 3958 -6889
rect 2154 -7110 3174 -7050
rect 3234 -7110 3240 -7050
rect 2154 -7252 2214 -7110
rect 2656 -7153 2716 -7110
rect 2452 -7159 2940 -7153
rect 2452 -7193 2464 -7159
rect 2928 -7193 2940 -7159
rect 2452 -7199 2940 -7193
rect 2154 -7312 2170 -7252
rect 2164 -7828 2170 -7312
rect 2204 -7312 2214 -7252
rect 3174 -7252 3234 -7110
rect 3684 -7153 3744 -6895
rect 3470 -7159 3958 -7153
rect 3470 -7193 3482 -7159
rect 3946 -7193 3958 -7159
rect 3470 -7199 3958 -7193
rect 2204 -7828 2210 -7312
rect 3174 -7316 3188 -7252
rect 2164 -7840 2210 -7828
rect 3182 -7828 3188 -7316
rect 3222 -7316 3234 -7252
rect 4192 -7252 4252 -6796
rect 5208 -6796 5224 -6710
rect 5258 -6710 5264 -6220
rect 6236 -6220 6282 -6208
rect 5258 -6796 5268 -6710
rect 6236 -6750 6242 -6220
rect 4488 -6855 4976 -6849
rect 4488 -6889 4500 -6855
rect 4964 -6889 4976 -6855
rect 4488 -6895 4976 -6889
rect 4702 -7153 4762 -6895
rect 5208 -6940 5268 -6796
rect 6228 -6796 6242 -6750
rect 6276 -6750 6282 -6220
rect 6276 -6796 6288 -6750
rect 5506 -6855 5994 -6849
rect 5506 -6889 5518 -6855
rect 5982 -6889 5994 -6855
rect 5506 -6895 5994 -6889
rect 5722 -6940 5782 -6895
rect 6228 -6940 6288 -6796
rect 5202 -7000 5208 -6940
rect 5268 -7000 6288 -6940
rect 4488 -7159 4976 -7153
rect 4488 -7193 4500 -7159
rect 4964 -7193 4976 -7159
rect 4488 -7199 4976 -7193
rect 3222 -7828 3228 -7316
rect 3182 -7840 3228 -7828
rect 4192 -7828 4206 -7252
rect 4240 -7828 4252 -7252
rect 5208 -7252 5268 -7000
rect 5722 -7153 5782 -7000
rect 5506 -7159 5994 -7153
rect 5506 -7193 5518 -7159
rect 5982 -7193 5994 -7159
rect 5506 -7199 5994 -7193
rect 5208 -7308 5224 -7252
rect 2452 -7887 2940 -7881
rect 2452 -7921 2464 -7887
rect 2928 -7921 2940 -7887
rect 2452 -7927 2940 -7921
rect 3470 -7887 3958 -7881
rect 3470 -7921 3482 -7887
rect 3946 -7921 3958 -7887
rect 3470 -7927 3958 -7921
rect 3690 -7974 3750 -7927
rect 1948 -8088 3238 -8028
rect 3684 -8034 3690 -7974
rect 3750 -8034 3756 -7974
rect 1888 -8094 1948 -8088
rect 2152 -8284 2212 -8088
rect 2660 -8185 2720 -8088
rect 2452 -8191 2940 -8185
rect 2452 -8225 2464 -8191
rect 2928 -8225 2940 -8191
rect 2452 -8231 2940 -8225
rect 2152 -8336 2170 -8284
rect 2164 -8860 2170 -8336
rect 2204 -8336 2212 -8284
rect 3178 -8284 3238 -8088
rect 3790 -8134 3796 -8074
rect 3856 -8134 3862 -8074
rect 3796 -8185 3856 -8134
rect 3470 -8191 3958 -8185
rect 3470 -8225 3482 -8191
rect 3946 -8225 3958 -8191
rect 3470 -8231 3958 -8225
rect 3178 -8332 3188 -8284
rect 2204 -8860 2210 -8336
rect 2164 -8872 2210 -8860
rect 3182 -8860 3188 -8332
rect 3222 -8332 3238 -8284
rect 4192 -8284 4252 -7828
rect 5218 -7828 5224 -7308
rect 5258 -7308 5268 -7252
rect 6228 -7252 6288 -7000
rect 6360 -7050 6420 -5020
rect 6354 -7110 6360 -7050
rect 6420 -7110 6426 -7050
rect 6228 -7288 6242 -7252
rect 5258 -7828 5264 -7308
rect 5218 -7840 5264 -7828
rect 6236 -7828 6242 -7288
rect 6276 -7288 6288 -7252
rect 6276 -7828 6282 -7288
rect 6236 -7840 6282 -7828
rect 4488 -7887 4976 -7881
rect 4488 -7921 4500 -7887
rect 4964 -7921 4976 -7887
rect 4488 -7927 4976 -7921
rect 5506 -7887 5994 -7881
rect 5506 -7921 5518 -7887
rect 5982 -7921 5994 -7887
rect 5506 -7927 5994 -7921
rect 4582 -8074 4642 -7927
rect 4694 -8034 4700 -7974
rect 4760 -8034 4766 -7974
rect 6360 -8028 6420 -7110
rect 6546 -7238 6552 -7178
rect 6612 -7238 6618 -7178
rect 4576 -8134 4582 -8074
rect 4642 -8134 4648 -8074
rect 4700 -8185 4760 -8034
rect 5208 -8088 6420 -8028
rect 4488 -8191 4976 -8185
rect 4488 -8225 4500 -8191
rect 4964 -8225 4976 -8191
rect 4488 -8231 4976 -8225
rect 3222 -8860 3228 -8332
rect 4192 -8358 4206 -8284
rect 3182 -8872 3228 -8860
rect 4200 -8860 4206 -8358
rect 4240 -8358 4252 -8284
rect 5208 -8284 5268 -8088
rect 5710 -8185 5770 -8088
rect 5506 -8191 5994 -8185
rect 5506 -8225 5518 -8191
rect 5982 -8225 5994 -8191
rect 5506 -8231 5994 -8225
rect 5208 -8314 5224 -8284
rect 4240 -8860 4246 -8358
rect 5218 -8778 5224 -8314
rect 4200 -8872 4246 -8860
rect 5210 -8860 5224 -8778
rect 5258 -8314 5268 -8284
rect 6228 -8284 6288 -8088
rect 5258 -8778 5264 -8314
rect 6228 -8352 6242 -8284
rect 5258 -8860 5270 -8778
rect 4688 -8913 4748 -8909
rect 2452 -8919 2940 -8913
rect 2452 -8953 2464 -8919
rect 2928 -8953 2940 -8919
rect 2452 -8959 2940 -8953
rect 3470 -8919 3958 -8913
rect 3470 -8953 3482 -8919
rect 3946 -8953 3958 -8919
rect 3470 -8959 3958 -8953
rect 4488 -8919 4976 -8913
rect 4488 -8953 4500 -8919
rect 4964 -8953 4976 -8919
rect 4488 -8959 4976 -8953
rect 1402 -9084 1462 -9078
rect 3682 -9084 3742 -8959
rect 1462 -9144 3742 -9084
rect 1402 -9150 1462 -9144
rect 1542 -9260 1602 -9254
rect 4688 -9260 4748 -8959
rect 1602 -9320 4748 -9260
rect 1542 -9326 1602 -9320
rect 2442 -9434 2502 -9428
rect 5210 -9434 5270 -8860
rect 6236 -8860 6242 -8352
rect 6276 -8352 6288 -8284
rect 6276 -8860 6282 -8352
rect 6236 -8872 6282 -8860
rect 5506 -8919 5994 -8913
rect 5506 -8953 5518 -8919
rect 5982 -8953 5994 -8919
rect 5506 -8959 5994 -8953
rect 2502 -9494 5270 -9434
rect 2442 -9500 2502 -9494
rect 1282 -9584 1342 -9578
rect 6552 -9584 6612 -7238
rect 6686 -8330 6746 -4402
rect 6796 -5012 6802 -4952
rect 6862 -5012 6868 -4952
rect 6802 -7074 6862 -5012
rect 7044 -5916 7104 -1654
rect 7488 -1784 7552 -1654
rect 7482 -1848 7488 -1784
rect 7552 -1848 7558 -1784
rect 7312 -1934 7372 -1928
rect 7312 -4870 7372 -1994
rect 7990 -2040 8050 -1485
rect 8510 -1536 8570 -1386
rect 9526 -1386 9542 -1362
rect 9576 -856 9594 -810
rect 10546 -810 10610 -458
rect 11040 -606 11100 -349
rect 11564 -496 11628 -250
rect 12580 -250 12596 -214
rect 12630 292 12638 326
rect 13600 326 13660 476
rect 14110 425 14170 787
rect 13896 419 14384 425
rect 13896 385 13908 419
rect 14372 385 14384 419
rect 13896 379 14384 385
rect 13600 300 13614 326
rect 12630 -214 12636 292
rect 12630 -216 12640 -214
rect 12630 -250 12644 -216
rect 11860 -309 12348 -303
rect 11860 -343 11872 -309
rect 12336 -343 12348 -309
rect 11860 -349 12348 -343
rect 11398 -560 11404 -496
rect 11468 -560 11628 -496
rect 12064 -606 12124 -349
rect 12580 -398 12644 -250
rect 13608 -250 13614 300
rect 13648 300 13660 326
rect 14616 326 14680 886
rect 15638 886 15650 924
rect 15684 924 15690 1462
rect 16658 1462 16718 1616
rect 17148 1561 17208 2064
rect 17668 1676 17728 2064
rect 17662 1616 17668 1676
rect 17728 1616 17734 1676
rect 16950 1555 17438 1561
rect 16950 1521 16962 1555
rect 17426 1521 17438 1555
rect 16950 1515 17438 1521
rect 16658 1424 16668 1462
rect 16662 926 16668 1424
rect 15684 886 15698 924
rect 15126 833 15186 839
rect 14914 827 15402 833
rect 14914 793 14926 827
rect 15390 793 15402 827
rect 14914 787 15402 793
rect 15126 425 15186 787
rect 15638 740 15698 886
rect 16654 886 16668 926
rect 16702 1424 16718 1462
rect 17668 1462 17728 1616
rect 18176 1561 18236 2064
rect 18690 1676 18750 2064
rect 19196 1858 19202 1918
rect 19262 1858 19268 1918
rect 20208 1858 20214 1918
rect 20274 1858 20280 1918
rect 18684 1616 18690 1676
rect 18750 1616 18756 1676
rect 17968 1555 18456 1561
rect 17968 1521 17980 1555
rect 18444 1521 18456 1555
rect 17968 1515 18456 1521
rect 18176 1512 18236 1515
rect 16702 926 16708 1424
rect 17668 1392 17686 1462
rect 16702 886 16718 926
rect 16138 833 16198 839
rect 15932 827 16420 833
rect 15932 793 15944 827
rect 16408 793 16420 827
rect 15932 787 16420 793
rect 15632 680 15638 740
rect 15698 680 15704 740
rect 16138 536 16198 787
rect 15630 476 15636 536
rect 15696 476 15702 536
rect 16132 476 16138 536
rect 16198 476 16204 536
rect 14914 419 15402 425
rect 14914 385 14926 419
rect 15390 385 15402 419
rect 14914 379 15402 385
rect 15126 376 15186 379
rect 13648 -250 13654 300
rect 14616 294 14632 326
rect 14626 -202 14632 294
rect 13608 -262 13654 -250
rect 14618 -250 14632 -202
rect 14666 294 14680 326
rect 15636 326 15696 476
rect 16138 425 16198 476
rect 15932 419 16420 425
rect 15932 385 15944 419
rect 16408 385 16420 419
rect 15932 379 16420 385
rect 16138 376 16198 379
rect 15636 294 15650 326
rect 14666 -202 14672 294
rect 14666 -204 14678 -202
rect 14666 -250 14682 -204
rect 15644 -220 15650 294
rect 13092 -303 13152 -296
rect 12878 -309 13366 -303
rect 12878 -343 12890 -309
rect 13354 -343 13366 -309
rect 12878 -349 13366 -343
rect 13896 -309 14384 -303
rect 13896 -343 13908 -309
rect 14372 -343 14384 -309
rect 13896 -349 14384 -343
rect 12574 -458 12580 -398
rect 12640 -458 12646 -398
rect 11034 -666 11040 -606
rect 11100 -666 11106 -606
rect 12058 -666 12064 -606
rect 12124 -666 12130 -606
rect 10842 -717 11330 -711
rect 10842 -751 10854 -717
rect 11318 -751 11330 -717
rect 10842 -757 11330 -751
rect 11860 -717 12348 -711
rect 11860 -751 11872 -717
rect 12336 -751 12348 -717
rect 11860 -757 12348 -751
rect 9576 -860 9592 -856
rect 10546 -858 10560 -810
rect 9576 -1362 9582 -860
rect 10554 -1360 10560 -858
rect 9576 -1386 9590 -1362
rect 8806 -1445 9294 -1439
rect 8806 -1479 8818 -1445
rect 9282 -1479 9294 -1445
rect 8806 -1485 9294 -1479
rect 8504 -1596 8510 -1536
rect 8570 -1596 8576 -1536
rect 9032 -2040 9092 -1485
rect 9526 -1646 9590 -1386
rect 10546 -1386 10560 -1360
rect 10594 -858 10610 -810
rect 11572 -810 11618 -798
rect 10594 -1360 10600 -858
rect 11572 -1330 11578 -810
rect 10594 -1362 10606 -1360
rect 10594 -1386 10610 -1362
rect 9824 -1445 10312 -1439
rect 9824 -1479 9836 -1445
rect 10300 -1479 10312 -1445
rect 9824 -1485 10312 -1479
rect 9520 -1710 9526 -1646
rect 9590 -1710 9596 -1646
rect 10032 -2040 10092 -1485
rect 10546 -1536 10610 -1386
rect 11566 -1386 11578 -1330
rect 11612 -1330 11618 -810
rect 12580 -810 12644 -458
rect 13092 -606 13152 -349
rect 13086 -666 13092 -606
rect 13152 -666 13158 -606
rect 13092 -711 13152 -666
rect 14120 -711 14180 -349
rect 14618 -400 14682 -250
rect 15638 -250 15650 -220
rect 15684 294 15696 326
rect 16654 326 16718 886
rect 17680 886 17686 1392
rect 17720 1392 17728 1462
rect 18690 1462 18750 1616
rect 19202 1561 19262 1858
rect 20214 1561 20274 1858
rect 20726 1676 20786 2064
rect 21226 1858 21232 1918
rect 21292 1858 21298 1918
rect 20720 1616 20726 1676
rect 20786 1616 20792 1676
rect 18986 1555 19474 1561
rect 18986 1521 18998 1555
rect 19462 1521 19474 1555
rect 18986 1515 19474 1521
rect 20004 1555 20492 1561
rect 20004 1521 20016 1555
rect 20480 1521 20492 1555
rect 20004 1515 20492 1521
rect 18690 1434 18704 1462
rect 17720 886 17726 1392
rect 18698 934 18704 1434
rect 17680 874 17726 886
rect 18690 886 18704 934
rect 18738 1434 18750 1462
rect 19716 1462 19762 1474
rect 18738 934 18744 1434
rect 18738 886 18750 934
rect 19716 918 19722 1462
rect 16950 827 17438 833
rect 16950 793 16962 827
rect 17426 793 17438 827
rect 16950 787 17438 793
rect 17968 827 18456 833
rect 17968 793 17980 827
rect 18444 793 18456 827
rect 17968 787 18456 793
rect 17666 576 17672 636
rect 17732 576 17738 636
rect 17152 476 17158 536
rect 17218 476 17224 536
rect 17158 425 17218 476
rect 16950 419 17438 425
rect 16950 385 16962 419
rect 17426 385 17438 419
rect 16950 379 17438 385
rect 15684 -220 15690 294
rect 16654 278 16668 326
rect 16662 -206 16668 278
rect 15684 -250 15698 -220
rect 15138 -303 15198 -291
rect 14914 -309 15402 -303
rect 14914 -343 14926 -309
rect 15390 -343 15402 -309
rect 14914 -349 15402 -343
rect 14612 -460 14618 -400
rect 14678 -460 14684 -400
rect 12878 -717 13366 -711
rect 12878 -751 12890 -717
rect 13354 -751 13366 -717
rect 12878 -757 13366 -751
rect 13896 -717 14384 -711
rect 13896 -751 13908 -717
rect 14372 -751 14384 -717
rect 13896 -757 14384 -751
rect 14120 -764 14180 -757
rect 12580 -870 12596 -810
rect 11612 -1386 11626 -1330
rect 12590 -1352 12596 -870
rect 11068 -1439 11128 -1436
rect 10842 -1445 11330 -1439
rect 10842 -1479 10854 -1445
rect 11318 -1479 11330 -1445
rect 10842 -1485 11330 -1479
rect 11068 -1536 11128 -1485
rect 11566 -1536 11626 -1386
rect 12580 -1386 12596 -1352
rect 12630 -870 12644 -810
rect 13608 -810 13654 -798
rect 12630 -1352 12636 -870
rect 12630 -1354 12640 -1352
rect 13608 -1354 13614 -810
rect 12630 -1386 12644 -1354
rect 11860 -1445 12348 -1439
rect 11860 -1479 11872 -1445
rect 12336 -1479 12348 -1445
rect 11860 -1485 12348 -1479
rect 10540 -1596 10546 -1536
rect 10606 -1596 10612 -1536
rect 11062 -1596 11068 -1536
rect 11128 -1596 11134 -1536
rect 11560 -1596 11566 -1536
rect 11626 -1596 11632 -1536
rect 12040 -1540 12100 -1485
rect 12580 -1532 12644 -1386
rect 13598 -1386 13614 -1354
rect 13648 -1354 13654 -810
rect 14618 -810 14682 -460
rect 15138 -711 15198 -349
rect 15638 -498 15698 -250
rect 16654 -250 16668 -206
rect 16702 278 16718 326
rect 17672 326 17732 576
rect 18178 476 18184 536
rect 18244 476 18250 536
rect 18690 532 18750 886
rect 19706 886 19722 918
rect 19756 918 19762 1462
rect 20726 1462 20786 1616
rect 21232 1561 21292 1858
rect 21746 1624 22826 1684
rect 21022 1555 21510 1561
rect 21022 1521 21034 1555
rect 21498 1521 21510 1555
rect 21022 1515 21510 1521
rect 20726 1430 20740 1462
rect 20734 924 20740 1430
rect 19756 886 19766 918
rect 18986 827 19474 833
rect 18986 793 18998 827
rect 19462 793 19474 827
rect 18986 787 19474 793
rect 19706 636 19766 886
rect 20730 886 20740 924
rect 20774 1430 20786 1462
rect 21746 1462 21806 1624
rect 22248 1561 22308 1624
rect 22040 1555 22528 1561
rect 22040 1521 22052 1555
rect 22516 1521 22528 1555
rect 22040 1515 22528 1521
rect 21746 1432 21758 1462
rect 20774 924 20780 1430
rect 21752 926 21758 1432
rect 20774 886 20790 924
rect 20004 827 20492 833
rect 20004 793 20016 827
rect 20480 793 20492 827
rect 20004 787 20492 793
rect 19700 576 19706 636
rect 19766 576 19772 636
rect 20730 538 20790 886
rect 21746 886 21758 926
rect 21792 1432 21806 1462
rect 22766 1462 22826 1624
rect 21792 926 21798 1432
rect 22766 1416 22776 1462
rect 21792 886 21806 926
rect 21210 833 21270 845
rect 21022 827 21510 833
rect 21022 793 21034 827
rect 21498 793 21510 827
rect 21022 787 21510 793
rect 20730 532 20794 538
rect 18184 425 18244 476
rect 18684 472 18690 532
rect 18750 472 18756 532
rect 19198 472 19204 532
rect 19264 472 19270 532
rect 19702 472 19708 532
rect 19768 472 19774 532
rect 20208 472 20214 532
rect 20274 472 20280 532
rect 20730 472 20734 532
rect 17968 419 18456 425
rect 17968 385 17980 419
rect 18444 385 18456 419
rect 17968 379 18456 385
rect 17672 302 17686 326
rect 16702 -206 16708 278
rect 16702 -208 16714 -206
rect 16702 -250 16718 -208
rect 16138 -303 16198 -295
rect 15932 -309 16420 -303
rect 15932 -343 15944 -309
rect 16408 -343 16420 -309
rect 15932 -349 16420 -343
rect 15632 -558 15638 -498
rect 15698 -558 15704 -498
rect 16138 -711 16198 -349
rect 16654 -400 16718 -250
rect 17680 -250 17686 302
rect 17720 302 17732 326
rect 18690 326 18750 472
rect 19204 425 19264 472
rect 18986 419 19474 425
rect 18986 385 18998 419
rect 19462 385 19474 419
rect 18986 379 19474 385
rect 17720 -250 17726 302
rect 18690 282 18704 326
rect 18698 -214 18704 282
rect 17680 -262 17726 -250
rect 18690 -250 18704 -214
rect 18738 282 18750 326
rect 19708 326 19768 472
rect 20214 425 20274 472
rect 20730 466 20794 472
rect 20004 419 20492 425
rect 20004 385 20016 419
rect 20480 385 20492 419
rect 20004 379 20492 385
rect 19708 298 19722 326
rect 18738 -214 18744 282
rect 19716 -180 19722 298
rect 18738 -250 18750 -214
rect 16950 -309 17438 -303
rect 16950 -343 16962 -309
rect 17426 -343 17438 -309
rect 16950 -349 17438 -343
rect 17968 -309 18456 -303
rect 17968 -343 17980 -309
rect 18444 -343 18456 -309
rect 17968 -349 18456 -343
rect 18690 -400 18750 -250
rect 19706 -250 19722 -180
rect 19756 298 19768 326
rect 20730 326 20790 466
rect 21210 425 21270 787
rect 21746 740 21806 886
rect 22770 886 22776 1416
rect 22810 1416 22826 1462
rect 22810 886 22816 1416
rect 22770 874 22816 886
rect 22040 827 22528 833
rect 22040 793 22052 827
rect 22516 793 22528 827
rect 22040 787 22528 793
rect 21740 680 21746 740
rect 21806 680 21812 740
rect 22990 680 22996 740
rect 23056 680 23062 740
rect 21750 464 22820 524
rect 21022 419 21510 425
rect 21022 385 21034 419
rect 21498 385 21510 419
rect 21022 379 21510 385
rect 19756 -180 19762 298
rect 20730 290 20740 326
rect 19756 -250 19766 -180
rect 20734 -218 20740 290
rect 18986 -309 19474 -303
rect 18986 -343 18998 -309
rect 19462 -343 19474 -309
rect 18986 -349 19474 -343
rect 19192 -400 19252 -349
rect 16648 -460 16654 -400
rect 16714 -460 16720 -400
rect 17148 -460 17154 -400
rect 17214 -460 17220 -400
rect 17662 -460 17668 -400
rect 17728 -460 17734 -400
rect 18186 -460 18192 -400
rect 18252 -460 18258 -400
rect 18684 -460 18690 -400
rect 18750 -460 18756 -400
rect 19186 -460 19192 -400
rect 19252 -460 19258 -400
rect 19706 -402 19766 -250
rect 20724 -250 20740 -218
rect 20774 290 20790 326
rect 21750 326 21810 464
rect 22256 425 22316 464
rect 22040 419 22528 425
rect 22040 385 22052 419
rect 22516 385 22528 419
rect 22040 379 22528 385
rect 21750 298 21758 326
rect 20774 -218 20780 290
rect 20774 -220 20784 -218
rect 21752 -220 21758 298
rect 20774 -250 20788 -220
rect 20214 -303 20274 -296
rect 20004 -309 20492 -303
rect 20004 -343 20016 -309
rect 20480 -343 20492 -309
rect 20004 -349 20492 -343
rect 20214 -402 20274 -349
rect 20724 -402 20788 -250
rect 21746 -250 21758 -220
rect 21792 298 21810 326
rect 22760 326 22820 464
rect 21792 -220 21798 298
rect 22760 292 22776 326
rect 21792 -250 21806 -220
rect 21210 -303 21270 -297
rect 21022 -309 21510 -303
rect 21022 -343 21034 -309
rect 21498 -343 21510 -309
rect 21022 -349 21510 -343
rect 14914 -717 15402 -711
rect 14914 -751 14926 -717
rect 15390 -751 15402 -717
rect 14914 -757 15402 -751
rect 15932 -717 16420 -711
rect 15932 -751 15944 -717
rect 16408 -751 16420 -717
rect 15932 -757 16420 -751
rect 16138 -758 16198 -757
rect 14618 -850 14632 -810
rect 14626 -1326 14632 -850
rect 13648 -1386 13662 -1354
rect 12878 -1445 13366 -1439
rect 12878 -1479 12890 -1445
rect 13354 -1479 13366 -1445
rect 12878 -1485 13366 -1479
rect 7422 -2100 7428 -2040
rect 7488 -2100 7494 -2040
rect 7984 -2100 7990 -2040
rect 8050 -2100 8056 -2040
rect 9026 -2100 9032 -2040
rect 9092 -2100 9098 -2040
rect 10026 -2100 10032 -2040
rect 10092 -2100 10098 -2040
rect 7428 -4682 7488 -2100
rect 12040 -2138 12100 -1600
rect 12548 -1536 12644 -1532
rect 12548 -1538 12580 -1536
rect 12640 -1596 12646 -1536
rect 13034 -1596 13040 -1536
rect 13100 -1596 13106 -1536
rect 12548 -2138 12608 -1598
rect 13040 -2138 13100 -1596
rect 13194 -2040 13254 -1485
rect 13598 -1788 13662 -1386
rect 14616 -1386 14632 -1326
rect 14666 -850 14682 -810
rect 15644 -810 15690 -798
rect 14666 -1326 14672 -850
rect 14666 -1386 14676 -1326
rect 15644 -1350 15650 -810
rect 13896 -1445 14384 -1439
rect 13896 -1479 13908 -1445
rect 14372 -1479 14384 -1445
rect 13896 -1485 14384 -1479
rect 13598 -1858 13662 -1852
rect 14084 -1534 14144 -1528
rect 13188 -2100 13194 -2040
rect 13254 -2100 13260 -2040
rect 14084 -2138 14144 -1594
rect 14204 -2040 14264 -1485
rect 14616 -1536 14676 -1386
rect 15634 -1386 15650 -1350
rect 15684 -1350 15690 -810
rect 16654 -810 16718 -460
rect 17154 -711 17214 -460
rect 16950 -717 17438 -711
rect 16950 -751 16962 -717
rect 17426 -751 17438 -717
rect 16950 -757 17438 -751
rect 16654 -862 16668 -810
rect 16662 -1344 16668 -862
rect 15684 -1386 15698 -1350
rect 14914 -1445 15402 -1439
rect 14914 -1479 14926 -1445
rect 15390 -1479 15402 -1445
rect 14914 -1485 15402 -1479
rect 14610 -1596 14616 -1536
rect 14676 -1596 14682 -1536
rect 15146 -2040 15206 -1485
rect 15634 -1930 15698 -1386
rect 16654 -1386 16668 -1344
rect 16702 -862 16718 -810
rect 17668 -810 17728 -460
rect 18192 -711 18252 -460
rect 17968 -717 18456 -711
rect 17968 -751 17980 -717
rect 18444 -751 18456 -717
rect 17968 -757 18456 -751
rect 16702 -1344 16708 -862
rect 17668 -864 17686 -810
rect 17680 -940 17686 -864
rect 16702 -1346 16714 -1344
rect 16702 -1386 16718 -1346
rect 15932 -1445 16420 -1439
rect 15932 -1479 15944 -1445
rect 16408 -1479 16420 -1445
rect 15932 -1485 16420 -1479
rect 16128 -1534 16188 -1528
rect 16654 -1534 16718 -1386
rect 17672 -1386 17686 -940
rect 17720 -864 17728 -810
rect 18690 -810 18750 -460
rect 19700 -462 19706 -402
rect 19766 -462 19772 -402
rect 20208 -462 20214 -402
rect 20274 -462 20280 -402
rect 20718 -462 20724 -402
rect 20784 -462 20790 -402
rect 19190 -674 19196 -614
rect 19256 -674 19262 -614
rect 20202 -674 20208 -614
rect 20268 -674 20274 -614
rect 19196 -711 19256 -674
rect 20208 -711 20268 -674
rect 18986 -717 19474 -711
rect 18986 -751 18998 -717
rect 19462 -751 19474 -717
rect 18986 -757 19474 -751
rect 20004 -717 20492 -711
rect 20004 -751 20016 -717
rect 20480 -751 20492 -717
rect 20004 -757 20492 -751
rect 18690 -864 18704 -810
rect 17720 -940 17726 -864
rect 17720 -1386 17732 -940
rect 18698 -1356 18704 -864
rect 17150 -1439 17210 -1430
rect 16950 -1445 17438 -1439
rect 16950 -1479 16962 -1445
rect 17426 -1479 17438 -1445
rect 16950 -1485 17438 -1479
rect 15628 -1994 15634 -1930
rect 15698 -1994 15704 -1930
rect 14198 -2100 14204 -2040
rect 14264 -2100 14270 -2040
rect 15140 -2100 15146 -2040
rect 15206 -2100 15212 -2040
rect 16128 -2138 16188 -1594
rect 16622 -1538 16718 -1534
rect 16622 -1540 16654 -1538
rect 16714 -1598 16720 -1538
rect 17150 -1544 17210 -1485
rect 17672 -1534 17732 -1386
rect 18690 -1386 18704 -1356
rect 18738 -864 18750 -810
rect 19716 -810 19762 -798
rect 18738 -1356 18744 -864
rect 19716 -1352 19722 -810
rect 18738 -1358 18750 -1356
rect 18738 -1386 18754 -1358
rect 18150 -1439 18210 -1436
rect 17968 -1445 18456 -1439
rect 17968 -1479 17980 -1445
rect 18444 -1479 18456 -1445
rect 17968 -1485 18456 -1479
rect 16622 -2138 16682 -1600
rect 17150 -2138 17210 -1604
rect 17638 -1540 17732 -1534
rect 17698 -1542 17732 -1540
rect 17638 -1602 17672 -1600
rect 17638 -1608 17732 -1602
rect 18150 -1544 18210 -1485
rect 18690 -1540 18754 -1386
rect 19706 -1386 19722 -1352
rect 19756 -1352 19762 -810
rect 20724 -810 20788 -462
rect 21210 -614 21270 -349
rect 21746 -498 21806 -250
rect 22770 -250 22776 292
rect 22810 292 22820 326
rect 22810 -250 22816 292
rect 22770 -262 22816 -250
rect 22040 -309 22528 -303
rect 22040 -343 22052 -309
rect 22516 -343 22528 -309
rect 22040 -349 22528 -343
rect 21740 -558 21746 -498
rect 21806 -558 21812 -498
rect 21748 -612 21808 -610
rect 21204 -674 21210 -614
rect 21270 -674 21276 -614
rect 21748 -672 22820 -612
rect 21210 -711 21270 -674
rect 21022 -717 21510 -711
rect 21022 -751 21034 -717
rect 21498 -751 21510 -717
rect 21022 -757 21510 -751
rect 21210 -760 21270 -757
rect 20724 -856 20740 -810
rect 19756 -1386 19770 -1352
rect 20734 -1356 20740 -856
rect 18986 -1445 19474 -1439
rect 18986 -1479 18998 -1445
rect 19462 -1479 19474 -1445
rect 18986 -1485 19474 -1479
rect 18684 -1600 18690 -1540
rect 18750 -1600 18756 -1540
rect 17638 -2138 17698 -1608
rect 18150 -2138 18210 -1604
rect 19706 -1646 19770 -1386
rect 20724 -1386 20740 -1356
rect 20774 -856 20788 -810
rect 21748 -810 21808 -672
rect 22252 -711 22312 -672
rect 22040 -717 22528 -711
rect 22040 -751 22052 -717
rect 22516 -751 22528 -717
rect 22040 -757 22528 -751
rect 21748 -836 21758 -810
rect 20774 -1356 20780 -856
rect 21752 -1298 21758 -836
rect 20774 -1358 20784 -1356
rect 20774 -1386 20788 -1358
rect 20004 -1445 20492 -1439
rect 20004 -1479 20016 -1445
rect 20480 -1479 20492 -1445
rect 20004 -1485 20492 -1479
rect 20724 -1540 20788 -1386
rect 21740 -1386 21758 -1298
rect 21792 -836 21808 -810
rect 22760 -810 22820 -672
rect 21792 -1298 21798 -836
rect 22760 -860 22776 -810
rect 21792 -1386 21800 -1298
rect 21022 -1445 21510 -1439
rect 21022 -1479 21034 -1445
rect 21498 -1479 21510 -1445
rect 21022 -1485 21510 -1479
rect 20718 -1600 20724 -1540
rect 20784 -1600 20790 -1540
rect 19700 -1710 19706 -1646
rect 19770 -1710 19776 -1646
rect 21740 -1934 21800 -1386
rect 22770 -1386 22776 -860
rect 22810 -860 22820 -810
rect 22810 -1386 22816 -860
rect 22770 -1398 22816 -1386
rect 22040 -1445 22528 -1439
rect 22040 -1479 22052 -1445
rect 22516 -1479 22528 -1445
rect 22040 -1485 22528 -1479
rect 22996 -1778 23056 680
rect 22992 -1784 23056 -1778
rect 22992 -1854 23056 -1848
rect 21734 -1994 21740 -1934
rect 21800 -1994 21806 -1934
rect 9704 -2198 19944 -2138
rect 7536 -2302 7542 -2242
rect 7602 -2302 7608 -2242
rect 7542 -4216 7602 -2302
rect 7964 -2355 8452 -2349
rect 7964 -2389 7976 -2355
rect 8440 -2389 8452 -2355
rect 7964 -2395 8452 -2389
rect 8982 -2355 9470 -2349
rect 8982 -2389 8994 -2355
rect 9458 -2389 9470 -2355
rect 8982 -2395 9470 -2389
rect 7676 -2448 7722 -2436
rect 7676 -2994 7682 -2448
rect 7668 -3024 7682 -2994
rect 7716 -2994 7722 -2448
rect 8694 -2448 8740 -2436
rect 7716 -3024 7728 -2994
rect 8694 -3000 8700 -2448
rect 7668 -3176 7728 -3024
rect 8686 -3024 8700 -3000
rect 8734 -3000 8740 -2448
rect 9704 -2448 9764 -2198
rect 10714 -2302 10720 -2242
rect 10780 -2302 10786 -2242
rect 10000 -2355 10488 -2349
rect 10000 -2389 10012 -2355
rect 10476 -2389 10488 -2355
rect 10000 -2395 10488 -2389
rect 8734 -3024 8746 -3000
rect 7964 -3083 8452 -3077
rect 7964 -3117 7976 -3083
rect 8440 -3117 8452 -3083
rect 7964 -3123 8452 -3117
rect 8180 -3176 8240 -3123
rect 8686 -3176 8746 -3024
rect 9704 -3024 9718 -2448
rect 9752 -3024 9764 -2448
rect 10720 -2448 10780 -2302
rect 11018 -2355 11506 -2349
rect 11018 -2389 11030 -2355
rect 11494 -2389 11506 -2355
rect 11018 -2395 11506 -2389
rect 10720 -2512 10736 -2448
rect 8982 -3083 9470 -3077
rect 8982 -3117 8994 -3083
rect 9458 -3117 9470 -3083
rect 8982 -3123 9470 -3117
rect 7668 -3178 8746 -3176
rect 7668 -3236 8686 -3178
rect 8680 -3238 8686 -3236
rect 8746 -3238 8752 -3178
rect 9190 -3286 9250 -3123
rect 9184 -3346 9190 -3286
rect 9250 -3346 9256 -3286
rect 9190 -3381 9250 -3346
rect 7964 -3387 8452 -3381
rect 7964 -3421 7976 -3387
rect 8440 -3421 8452 -3387
rect 7964 -3427 8452 -3421
rect 8982 -3387 9470 -3381
rect 8982 -3421 8994 -3387
rect 9458 -3421 9470 -3387
rect 8982 -3427 9470 -3421
rect 7676 -3480 7722 -3468
rect 7676 -4000 7682 -3480
rect 7668 -4056 7682 -4000
rect 7716 -4000 7722 -3480
rect 8694 -3480 8740 -3468
rect 7716 -4056 7728 -4000
rect 8694 -4026 8700 -3480
rect 7668 -4216 7728 -4056
rect 8682 -4056 8700 -4026
rect 8734 -4026 8740 -3480
rect 9704 -3480 9764 -3024
rect 10730 -3024 10736 -2512
rect 10770 -2512 10780 -2448
rect 11742 -2448 11802 -2198
rect 12036 -2355 12524 -2349
rect 12036 -2389 12048 -2355
rect 12512 -2389 12524 -2355
rect 12036 -2395 12524 -2389
rect 13054 -2355 13542 -2349
rect 13054 -2389 13066 -2355
rect 13530 -2389 13542 -2355
rect 13054 -2395 13542 -2389
rect 10770 -3024 10776 -2512
rect 10730 -3036 10776 -3024
rect 11742 -3024 11754 -2448
rect 11788 -3024 11802 -2448
rect 12766 -2448 12812 -2436
rect 12766 -2960 12772 -2448
rect 10210 -3077 10270 -3071
rect 10000 -3083 10488 -3077
rect 10000 -3117 10012 -3083
rect 10476 -3117 10488 -3083
rect 10000 -3123 10488 -3117
rect 11018 -3083 11506 -3077
rect 11018 -3117 11030 -3083
rect 11494 -3117 11506 -3083
rect 11018 -3123 11506 -3117
rect 10210 -3280 10270 -3123
rect 10714 -3238 10720 -3178
rect 10780 -3238 10786 -3178
rect 10210 -3286 10272 -3280
rect 10210 -3346 10212 -3286
rect 10210 -3352 10272 -3346
rect 10210 -3381 10270 -3352
rect 10000 -3387 10488 -3381
rect 10000 -3421 10012 -3387
rect 10476 -3421 10488 -3387
rect 10000 -3427 10488 -3421
rect 8734 -4056 8742 -4026
rect 7964 -4115 8452 -4109
rect 7964 -4149 7976 -4115
rect 8440 -4149 8452 -4115
rect 7964 -4155 8452 -4149
rect 8170 -4216 8230 -4155
rect 8682 -4210 8742 -4056
rect 9704 -4056 9718 -3480
rect 9752 -4056 9764 -3480
rect 10720 -3480 10780 -3238
rect 11232 -3280 11292 -3123
rect 11230 -3286 11292 -3280
rect 11290 -3346 11292 -3286
rect 11230 -3352 11292 -3346
rect 11232 -3381 11292 -3352
rect 11018 -3387 11506 -3381
rect 11018 -3421 11030 -3387
rect 11494 -3421 11506 -3387
rect 11018 -3427 11506 -3421
rect 11232 -3434 11292 -3427
rect 10720 -3526 10736 -3480
rect 8982 -4115 9470 -4109
rect 8982 -4149 8994 -4115
rect 9458 -4149 9470 -4115
rect 8982 -4155 9470 -4149
rect 8676 -4216 8682 -4210
rect 7542 -4270 8682 -4216
rect 8742 -4270 8748 -4210
rect 7542 -4276 8748 -4270
rect 9188 -4344 9248 -4155
rect 9188 -4410 9248 -4404
rect 9704 -4552 9764 -4056
rect 10730 -4056 10736 -3526
rect 10770 -3526 10780 -3480
rect 11742 -3480 11802 -3024
rect 12762 -3024 12772 -2960
rect 12806 -2960 12812 -2448
rect 13780 -2448 13840 -2198
rect 14782 -2302 14788 -2242
rect 14848 -2302 14854 -2242
rect 14072 -2355 14560 -2349
rect 14072 -2389 14084 -2355
rect 14548 -2389 14560 -2355
rect 14072 -2395 14560 -2389
rect 12806 -3024 12822 -2960
rect 12036 -3083 12524 -3077
rect 12036 -3117 12048 -3083
rect 12512 -3117 12524 -3083
rect 12036 -3123 12524 -3117
rect 12252 -3280 12312 -3123
rect 12762 -3178 12822 -3024
rect 13780 -3024 13790 -2448
rect 13824 -3024 13840 -2448
rect 14788 -2448 14848 -2302
rect 15090 -2355 15578 -2349
rect 15090 -2389 15102 -2355
rect 15566 -2389 15578 -2355
rect 15090 -2395 15578 -2389
rect 14788 -2522 14808 -2448
rect 13268 -3077 13328 -3075
rect 13054 -3083 13542 -3077
rect 13054 -3117 13066 -3083
rect 13530 -3117 13542 -3083
rect 13054 -3123 13542 -3117
rect 12756 -3238 12762 -3178
rect 12822 -3238 12828 -3178
rect 12252 -3286 12314 -3280
rect 12252 -3346 12254 -3286
rect 12252 -3352 12314 -3346
rect 13268 -3286 13328 -3123
rect 12252 -3381 12312 -3352
rect 13268 -3381 13328 -3346
rect 12036 -3387 12524 -3381
rect 12036 -3421 12048 -3387
rect 12512 -3421 12524 -3387
rect 12036 -3427 12524 -3421
rect 13054 -3387 13542 -3381
rect 13054 -3421 13066 -3387
rect 13530 -3421 13542 -3387
rect 13054 -3427 13542 -3421
rect 10770 -4056 10776 -3526
rect 10730 -4068 10776 -4056
rect 11742 -4056 11754 -3480
rect 11788 -4056 11802 -3480
rect 12766 -3480 12812 -3468
rect 12766 -3990 12772 -3480
rect 10202 -4109 10262 -4106
rect 10000 -4115 10488 -4109
rect 10000 -4149 10012 -4115
rect 10476 -4149 10488 -4115
rect 10000 -4155 10488 -4149
rect 11018 -4115 11506 -4109
rect 11018 -4149 11030 -4115
rect 11494 -4149 11506 -4115
rect 11018 -4155 11506 -4149
rect 10202 -4348 10262 -4155
rect 11234 -4340 11294 -4155
rect 11234 -4406 11294 -4400
rect 10202 -4414 10262 -4408
rect 11742 -4552 11802 -4056
rect 12762 -4056 12772 -3990
rect 12806 -3990 12812 -3480
rect 13780 -3480 13840 -3024
rect 14802 -3024 14808 -2522
rect 14842 -3024 14848 -2448
rect 14802 -3036 14848 -3024
rect 15816 -2448 15876 -2198
rect 16108 -2355 16596 -2349
rect 16108 -2389 16120 -2355
rect 16584 -2389 16596 -2355
rect 16108 -2395 16596 -2389
rect 17126 -2355 17614 -2349
rect 17126 -2389 17138 -2355
rect 17602 -2389 17614 -2355
rect 17126 -2395 17614 -2389
rect 15816 -3024 15826 -2448
rect 15860 -3024 15876 -2448
rect 16838 -2448 16884 -2436
rect 16838 -2960 16844 -2448
rect 14072 -3083 14560 -3077
rect 14072 -3117 14084 -3083
rect 14548 -3117 14560 -3083
rect 14072 -3123 14560 -3117
rect 15090 -3083 15578 -3077
rect 15090 -3117 15102 -3083
rect 15566 -3117 15578 -3083
rect 15090 -3123 15578 -3117
rect 14284 -3280 14344 -3123
rect 14782 -3238 14788 -3178
rect 14848 -3238 14854 -3178
rect 14284 -3286 14346 -3280
rect 14284 -3346 14286 -3286
rect 14284 -3352 14346 -3346
rect 14284 -3381 14344 -3352
rect 14072 -3387 14560 -3381
rect 14072 -3421 14084 -3387
rect 14548 -3421 14560 -3387
rect 14072 -3427 14560 -3421
rect 12806 -4056 12822 -3990
rect 12036 -4115 12524 -4109
rect 12036 -4149 12048 -4115
rect 12512 -4149 12524 -4115
rect 12036 -4155 12524 -4149
rect 12232 -4340 12292 -4155
rect 12762 -4210 12822 -4056
rect 13780 -4056 13790 -3480
rect 13824 -4056 13840 -3480
rect 14788 -3480 14848 -3238
rect 15294 -3280 15354 -3123
rect 15294 -3286 15356 -3280
rect 15294 -3346 15296 -3286
rect 15294 -3352 15356 -3346
rect 15294 -3381 15354 -3352
rect 15090 -3387 15578 -3381
rect 15090 -3421 15102 -3387
rect 15566 -3421 15578 -3387
rect 15090 -3427 15578 -3421
rect 14788 -3542 14808 -3480
rect 14802 -3964 14808 -3542
rect 13276 -4109 13336 -4096
rect 13054 -4115 13542 -4109
rect 13054 -4149 13066 -4115
rect 13530 -4149 13542 -4115
rect 13054 -4155 13542 -4149
rect 12756 -4270 12762 -4210
rect 12822 -4270 12828 -4210
rect 12232 -4406 12292 -4400
rect 13276 -4340 13336 -4155
rect 13276 -4406 13336 -4400
rect 13780 -4552 13840 -4056
rect 14798 -4056 14808 -3964
rect 14842 -3964 14848 -3480
rect 15816 -3480 15876 -3024
rect 16830 -3024 16844 -2960
rect 16878 -2960 16884 -2448
rect 17846 -2448 17906 -2198
rect 18858 -2302 18864 -2242
rect 18924 -2302 18930 -2242
rect 18144 -2355 18632 -2349
rect 18144 -2389 18156 -2355
rect 18620 -2389 18632 -2355
rect 18144 -2395 18632 -2389
rect 17846 -2858 17862 -2448
rect 17856 -2952 17862 -2858
rect 16878 -3024 16890 -2960
rect 16316 -3077 16376 -3075
rect 16108 -3083 16596 -3077
rect 16108 -3117 16120 -3083
rect 16584 -3117 16596 -3083
rect 16108 -3123 16596 -3117
rect 16316 -3280 16376 -3123
rect 16830 -3178 16890 -3024
rect 17846 -3024 17862 -2952
rect 17896 -2858 17906 -2448
rect 18864 -2448 18924 -2302
rect 19162 -2355 19650 -2349
rect 19162 -2389 19174 -2355
rect 19638 -2389 19650 -2355
rect 19162 -2395 19650 -2389
rect 18864 -2512 18880 -2448
rect 17896 -2952 17902 -2858
rect 17896 -3024 17906 -2952
rect 17330 -3077 17390 -3075
rect 17126 -3083 17614 -3077
rect 17126 -3117 17138 -3083
rect 17602 -3117 17614 -3083
rect 17126 -3123 17614 -3117
rect 16824 -3238 16830 -3178
rect 16890 -3238 16896 -3178
rect 17330 -3280 17390 -3123
rect 16316 -3286 16378 -3280
rect 16316 -3346 16318 -3286
rect 16316 -3352 16378 -3346
rect 17330 -3286 17392 -3280
rect 17330 -3346 17332 -3286
rect 17330 -3352 17392 -3346
rect 16316 -3381 16376 -3352
rect 17330 -3381 17390 -3352
rect 16108 -3387 16596 -3381
rect 16108 -3421 16120 -3387
rect 16584 -3421 16596 -3387
rect 16108 -3427 16596 -3421
rect 17126 -3387 17614 -3381
rect 17126 -3421 17138 -3387
rect 17602 -3421 17614 -3387
rect 17126 -3427 17614 -3421
rect 14842 -4056 14858 -3964
rect 14280 -4109 14340 -4106
rect 14072 -4115 14560 -4109
rect 14072 -4149 14084 -4115
rect 14548 -4149 14560 -4115
rect 14072 -4155 14560 -4149
rect 14280 -4344 14340 -4155
rect 14280 -4410 14340 -4404
rect 14798 -4460 14858 -4056
rect 15816 -4056 15826 -3480
rect 15860 -4056 15876 -3480
rect 16838 -3480 16884 -3468
rect 16838 -3974 16844 -3480
rect 15296 -4109 15356 -4102
rect 15090 -4115 15578 -4109
rect 15090 -4149 15102 -4115
rect 15566 -4149 15578 -4115
rect 15090 -4155 15578 -4149
rect 15296 -4344 15356 -4155
rect 15296 -4410 15356 -4404
rect 14588 -4520 14858 -4460
rect 9704 -4612 14080 -4552
rect 14140 -4612 14146 -4552
rect 7428 -4742 11596 -4682
rect 7306 -4930 7312 -4870
rect 7372 -4930 7378 -4870
rect 8472 -4930 8478 -4870
rect 8538 -4930 8544 -4870
rect 7038 -5976 7044 -5916
rect 7104 -5976 7110 -5916
rect 6796 -7134 6802 -7074
rect 6862 -7134 6868 -7074
rect 6792 -7348 6798 -7288
rect 6858 -7348 6864 -7288
rect 6680 -8390 6686 -8330
rect 6746 -8390 6752 -8330
rect 1342 -9644 6612 -9584
rect 1282 -9650 1342 -9644
rect -13992 -10182 -2722 -10122
rect -13992 -10670 -13926 -10182
rect -13698 -10378 -2722 -10182
rect 372 -10242 484 -9728
rect 2336 -9846 2396 -9840
rect 6798 -9846 6858 -7348
rect 7044 -9588 7104 -5976
rect 7174 -6074 7180 -6014
rect 7240 -6074 7246 -6014
rect 7038 -9648 7044 -9588
rect 7104 -9648 7110 -9588
rect 7180 -9718 7240 -6074
rect 7312 -8538 7372 -4930
rect 7756 -4991 8244 -4985
rect 7756 -5025 7768 -4991
rect 8232 -5025 8244 -4991
rect 7756 -5031 8244 -5025
rect 7468 -5084 7514 -5072
rect 7468 -5624 7474 -5084
rect 7460 -5660 7474 -5624
rect 7508 -5624 7514 -5084
rect 8478 -5084 8538 -4930
rect 8774 -4991 9262 -4985
rect 8774 -5025 8786 -4991
rect 9250 -5025 9262 -4991
rect 8774 -5031 9262 -5025
rect 8478 -5110 8492 -5084
rect 7508 -5660 7520 -5624
rect 8486 -5636 8492 -5110
rect 7460 -5818 7520 -5660
rect 8476 -5660 8492 -5636
rect 8526 -5110 8538 -5084
rect 9494 -5084 9554 -4742
rect 10508 -4930 10514 -4870
rect 10574 -4930 10580 -4870
rect 9792 -4991 10280 -4985
rect 9792 -5025 9804 -4991
rect 10268 -5025 10280 -4991
rect 9792 -5031 10280 -5025
rect 8526 -5636 8532 -5110
rect 9494 -5130 9510 -5084
rect 9504 -5636 9510 -5130
rect 8526 -5660 8536 -5636
rect 7756 -5719 8244 -5713
rect 7756 -5753 7768 -5719
rect 8232 -5753 8244 -5719
rect 7756 -5759 8244 -5753
rect 7974 -5818 8034 -5759
rect 8476 -5818 8536 -5660
rect 9496 -5660 9510 -5636
rect 9544 -5130 9554 -5084
rect 10514 -5084 10574 -4930
rect 11016 -4934 11022 -4870
rect 11086 -4934 11092 -4870
rect 11022 -4985 11086 -4934
rect 10810 -4991 11298 -4985
rect 10810 -5025 10822 -4991
rect 11286 -5025 11298 -4991
rect 10810 -5031 11298 -5025
rect 10514 -5108 10528 -5084
rect 9544 -5636 9550 -5130
rect 9544 -5660 9556 -5636
rect 8774 -5719 9262 -5713
rect 8774 -5753 8786 -5719
rect 9250 -5753 9262 -5719
rect 8774 -5759 9262 -5753
rect 7460 -5878 8536 -5818
rect 8966 -6120 9026 -5759
rect 9496 -5818 9556 -5660
rect 10522 -5660 10528 -5108
rect 10562 -5108 10574 -5084
rect 11536 -5084 11596 -4742
rect 12040 -4985 12100 -4612
rect 11828 -4991 12316 -4985
rect 11828 -5025 11840 -4991
rect 12304 -5025 12316 -4991
rect 11828 -5031 12316 -5025
rect 10562 -5660 10568 -5108
rect 11536 -5138 11546 -5084
rect 11540 -5632 11546 -5138
rect 10522 -5672 10568 -5660
rect 11532 -5660 11546 -5632
rect 11580 -5138 11596 -5084
rect 12548 -5084 12608 -4612
rect 13040 -4985 13100 -4612
rect 14078 -4985 14138 -4612
rect 12846 -4991 13334 -4985
rect 12846 -5025 12858 -4991
rect 13322 -5025 13334 -4991
rect 12846 -5031 13334 -5025
rect 13864 -4991 14352 -4985
rect 13864 -5025 13876 -4991
rect 14340 -5025 14352 -4991
rect 13864 -5031 14352 -5025
rect 11580 -5632 11586 -5138
rect 11580 -5660 11592 -5632
rect 9792 -5719 10280 -5713
rect 9792 -5753 9804 -5719
rect 10268 -5753 10280 -5719
rect 9792 -5759 10280 -5753
rect 10810 -5719 11298 -5713
rect 10810 -5753 10822 -5719
rect 11286 -5753 11298 -5719
rect 10810 -5759 11298 -5753
rect 9490 -5878 9496 -5818
rect 9556 -5878 9562 -5818
rect 10004 -5872 10064 -5759
rect 11010 -5872 11070 -5759
rect 11532 -5818 11592 -5660
rect 12548 -5660 12564 -5084
rect 12598 -5660 12608 -5084
rect 13576 -5084 13622 -5072
rect 13576 -5636 13582 -5084
rect 11828 -5719 12316 -5713
rect 11828 -5753 11840 -5719
rect 12304 -5753 12316 -5719
rect 11828 -5759 12316 -5753
rect 12042 -5814 12102 -5759
rect 12548 -5814 12608 -5660
rect 13568 -5660 13582 -5636
rect 13616 -5636 13622 -5084
rect 14588 -5084 14648 -4520
rect 15816 -4552 15876 -4056
rect 16830 -4056 16844 -3974
rect 16878 -3974 16884 -3480
rect 17846 -3480 17906 -3024
rect 18874 -3024 18880 -2512
rect 18914 -2512 18924 -2448
rect 19884 -2448 19944 -2198
rect 22054 -2302 22060 -2242
rect 22120 -2302 22126 -2242
rect 20180 -2355 20668 -2349
rect 20180 -2389 20192 -2355
rect 20656 -2389 20668 -2355
rect 20180 -2395 20668 -2389
rect 21198 -2355 21686 -2349
rect 21198 -2389 21210 -2355
rect 21674 -2389 21686 -2355
rect 21198 -2395 21686 -2389
rect 18914 -3024 18920 -2512
rect 18874 -3036 18920 -3024
rect 19884 -3024 19898 -2448
rect 19932 -3024 19944 -2448
rect 20910 -2448 20956 -2436
rect 20910 -2948 20916 -2448
rect 18362 -3077 18422 -3075
rect 19372 -3077 19432 -3075
rect 18144 -3083 18632 -3077
rect 18144 -3117 18156 -3083
rect 18620 -3117 18632 -3083
rect 18144 -3123 18632 -3117
rect 19162 -3083 19650 -3077
rect 19162 -3117 19174 -3083
rect 19638 -3117 19650 -3083
rect 19162 -3123 19650 -3117
rect 18362 -3280 18422 -3123
rect 18860 -3238 18866 -3178
rect 18926 -3238 18932 -3178
rect 18362 -3286 18424 -3280
rect 18362 -3346 18364 -3286
rect 18362 -3352 18424 -3346
rect 18362 -3381 18422 -3352
rect 18144 -3387 18632 -3381
rect 18144 -3421 18156 -3387
rect 18620 -3421 18632 -3387
rect 18144 -3427 18632 -3421
rect 16878 -4056 16890 -3974
rect 16108 -4115 16596 -4109
rect 16108 -4149 16120 -4115
rect 16584 -4149 16596 -4115
rect 16108 -4155 16596 -4149
rect 16300 -4344 16360 -4155
rect 16830 -4210 16890 -4056
rect 17846 -4056 17862 -3480
rect 17896 -4056 17906 -3480
rect 18866 -3480 18926 -3238
rect 19372 -3280 19432 -3123
rect 19372 -3286 19434 -3280
rect 19372 -3346 19374 -3286
rect 19372 -3352 19434 -3346
rect 19372 -3381 19432 -3352
rect 19162 -3387 19650 -3381
rect 19162 -3421 19174 -3387
rect 19638 -3421 19650 -3387
rect 19162 -3427 19650 -3421
rect 18866 -3548 18880 -3480
rect 17126 -4115 17614 -4109
rect 17126 -4149 17138 -4115
rect 17602 -4149 17614 -4115
rect 17126 -4155 17614 -4149
rect 16824 -4270 16830 -4210
rect 16890 -4270 16896 -4210
rect 16300 -4410 16360 -4404
rect 17332 -4340 17392 -4155
rect 17332 -4406 17392 -4400
rect 15090 -4812 15096 -4748
rect 15160 -4812 15166 -4748
rect 15096 -4870 15160 -4812
rect 15816 -4842 15876 -4612
rect 17846 -4452 17906 -4056
rect 18874 -4056 18880 -3548
rect 18914 -3548 18926 -3480
rect 19884 -3480 19944 -3024
rect 20902 -3024 20916 -2948
rect 20950 -2948 20956 -2448
rect 21928 -2448 21974 -2436
rect 20950 -3024 20962 -2948
rect 21928 -2998 21934 -2448
rect 20180 -3083 20668 -3077
rect 20180 -3117 20192 -3083
rect 20656 -3117 20668 -3083
rect 20180 -3123 20668 -3117
rect 20394 -3280 20454 -3123
rect 20902 -3176 20962 -3024
rect 21918 -3024 21934 -2998
rect 21968 -2998 21974 -2448
rect 21968 -3024 21978 -2998
rect 21198 -3083 21686 -3077
rect 21198 -3117 21210 -3083
rect 21674 -3117 21686 -3083
rect 21198 -3123 21686 -3117
rect 21424 -3176 21484 -3123
rect 21918 -3176 21978 -3024
rect 20902 -3178 21978 -3176
rect 20896 -3238 20902 -3178
rect 20962 -3236 21978 -3178
rect 20962 -3238 20968 -3236
rect 20394 -3286 20456 -3280
rect 20394 -3346 20396 -3286
rect 20394 -3352 20456 -3346
rect 20394 -3381 20454 -3352
rect 20180 -3387 20668 -3381
rect 20180 -3421 20192 -3387
rect 20656 -3421 20668 -3387
rect 20180 -3427 20668 -3421
rect 21198 -3387 21686 -3381
rect 21198 -3421 21210 -3387
rect 21674 -3421 21686 -3387
rect 21198 -3427 21686 -3421
rect 18914 -4056 18920 -3548
rect 18874 -4068 18920 -4056
rect 19884 -4056 19898 -3480
rect 19932 -4056 19944 -3480
rect 20910 -3480 20956 -3468
rect 20910 -3980 20916 -3480
rect 18348 -4109 18408 -4106
rect 18144 -4115 18632 -4109
rect 18144 -4149 18156 -4115
rect 18620 -4149 18632 -4115
rect 18144 -4155 18632 -4149
rect 19162 -4115 19650 -4109
rect 19162 -4149 19174 -4115
rect 19638 -4149 19650 -4115
rect 19162 -4155 19650 -4149
rect 18348 -4344 18408 -4155
rect 18348 -4410 18408 -4404
rect 19376 -4344 19436 -4155
rect 19376 -4410 19436 -4404
rect 19884 -4452 19944 -4056
rect 20898 -4056 20916 -3980
rect 20950 -3980 20956 -3480
rect 21928 -3480 21974 -3468
rect 20950 -4056 20958 -3980
rect 21928 -3984 21934 -3480
rect 20396 -4109 20456 -4106
rect 20180 -4115 20668 -4109
rect 20180 -4149 20192 -4115
rect 20656 -4149 20668 -4115
rect 20180 -4155 20668 -4149
rect 20396 -4344 20456 -4155
rect 20898 -4206 20958 -4056
rect 21918 -4056 21934 -3984
rect 21968 -3984 21974 -3480
rect 21968 -4056 21978 -3984
rect 21198 -4115 21686 -4109
rect 21198 -4149 21210 -4115
rect 21674 -4149 21686 -4115
rect 21198 -4155 21686 -4149
rect 21386 -4206 21446 -4155
rect 21918 -4206 21978 -4056
rect 22060 -4206 22120 -2302
rect 20896 -4210 22120 -4206
rect 20892 -4270 20898 -4210
rect 20958 -4266 22120 -4210
rect 20958 -4270 20964 -4266
rect 22848 -4402 22854 -4342
rect 22914 -4402 22920 -4342
rect 20396 -4410 20456 -4404
rect 17846 -4512 19944 -4452
rect 17846 -4842 17906 -4512
rect 21708 -4628 21714 -4568
rect 21774 -4628 21780 -4568
rect 19154 -4812 19160 -4748
rect 19224 -4812 19230 -4748
rect 20178 -4812 20184 -4748
rect 20248 -4812 20254 -4748
rect 21190 -4812 21196 -4748
rect 21260 -4812 21266 -4748
rect 15092 -4934 15098 -4870
rect 15162 -4934 15168 -4870
rect 15816 -4902 18210 -4842
rect 19160 -4866 19224 -4812
rect 15096 -4985 15160 -4934
rect 16128 -4985 16188 -4902
rect 14882 -4991 15370 -4985
rect 14882 -5025 14894 -4991
rect 15358 -5025 15370 -4991
rect 14882 -5031 15370 -5025
rect 15900 -4991 16388 -4985
rect 15900 -5025 15912 -4991
rect 16376 -5025 16388 -4991
rect 15900 -5031 16388 -5025
rect 13616 -5660 13628 -5636
rect 12846 -5719 13334 -5713
rect 12846 -5753 12858 -5719
rect 13322 -5753 13334 -5719
rect 12846 -5759 13334 -5753
rect 13062 -5814 13122 -5759
rect 13568 -5814 13628 -5660
rect 14588 -5660 14600 -5084
rect 14634 -5660 14648 -5084
rect 15612 -5084 15658 -5072
rect 15612 -5582 15618 -5084
rect 13864 -5719 14352 -5713
rect 13864 -5753 13876 -5719
rect 14340 -5753 14352 -5719
rect 13864 -5759 14352 -5753
rect 14072 -5814 14132 -5759
rect 9496 -6014 9556 -5878
rect 10004 -5932 11070 -5872
rect 11526 -5878 11532 -5818
rect 11592 -5878 11598 -5818
rect 11868 -5876 11874 -5816
rect 11934 -5876 11940 -5816
rect 12042 -5874 14132 -5814
rect 14588 -5816 14648 -5660
rect 15606 -5660 15618 -5582
rect 15652 -5582 15658 -5084
rect 16622 -5084 16682 -4902
rect 17150 -4985 17210 -4902
rect 16918 -4991 17406 -4985
rect 16918 -5025 16930 -4991
rect 17394 -5025 17406 -4991
rect 16918 -5031 17406 -5025
rect 17150 -5032 17210 -5031
rect 15652 -5660 15666 -5582
rect 14882 -5719 15370 -5713
rect 14882 -5753 14894 -5719
rect 15358 -5753 15370 -5719
rect 14882 -5759 15370 -5753
rect 9490 -6074 9496 -6014
rect 9556 -6074 9562 -6014
rect 10004 -6120 10064 -5932
rect 10510 -6072 10516 -6012
rect 10576 -6072 10582 -6012
rect 8476 -6184 8482 -6124
rect 8542 -6184 8548 -6124
rect 8966 -6180 10064 -6120
rect 10516 -6124 10576 -6072
rect 7756 -6247 8244 -6241
rect 7756 -6281 7768 -6247
rect 8232 -6281 8244 -6247
rect 7756 -6287 8244 -6281
rect 7468 -6340 7514 -6328
rect 7468 -6880 7474 -6340
rect 7464 -6916 7474 -6880
rect 7508 -6880 7514 -6340
rect 8482 -6340 8542 -6184
rect 8966 -6241 9026 -6180
rect 10004 -6241 10064 -6180
rect 10510 -6184 10516 -6124
rect 10576 -6184 10582 -6124
rect 8774 -6247 9262 -6241
rect 8774 -6281 8786 -6247
rect 9250 -6281 9262 -6247
rect 8774 -6287 9262 -6281
rect 9792 -6247 10280 -6241
rect 9792 -6281 9804 -6247
rect 10268 -6281 10280 -6247
rect 9792 -6287 10280 -6281
rect 8482 -6366 8492 -6340
rect 7508 -6916 7524 -6880
rect 8486 -6892 8492 -6366
rect 7464 -7074 7524 -6916
rect 8480 -6916 8492 -6892
rect 8526 -6366 8542 -6340
rect 9504 -6340 9550 -6328
rect 8526 -6892 8532 -6366
rect 9504 -6890 9510 -6340
rect 8526 -6916 8540 -6892
rect 7756 -6975 8244 -6969
rect 7756 -7009 7768 -6975
rect 8232 -7009 8244 -6975
rect 7756 -7015 8244 -7009
rect 7978 -7074 8038 -7015
rect 8480 -7074 8540 -6916
rect 9498 -6916 9510 -6890
rect 9544 -6890 9550 -6340
rect 10516 -6340 10576 -6184
rect 11010 -6241 11070 -5932
rect 11874 -6130 11934 -5876
rect 11532 -6190 11934 -6130
rect 10810 -6247 11298 -6241
rect 10810 -6281 10822 -6247
rect 11286 -6281 11298 -6247
rect 10810 -6287 11298 -6281
rect 10516 -6362 10528 -6340
rect 9544 -6916 9558 -6890
rect 8960 -6969 9020 -6968
rect 8774 -6975 9262 -6969
rect 8774 -7009 8786 -6975
rect 9250 -7009 9262 -6975
rect 8774 -7015 9262 -7009
rect 7464 -7134 8540 -7074
rect 7464 -7288 7524 -7134
rect 7458 -7348 7464 -7288
rect 7524 -7348 7530 -7288
rect 7462 -7458 8538 -7398
rect 7462 -7596 7522 -7458
rect 7976 -7497 8036 -7458
rect 7756 -7503 8244 -7497
rect 7756 -7537 7768 -7503
rect 8232 -7537 8244 -7503
rect 7756 -7543 8244 -7537
rect 7462 -7630 7474 -7596
rect 7468 -8172 7474 -7630
rect 7508 -7630 7522 -7596
rect 8478 -7596 8538 -7458
rect 8960 -7497 9020 -7015
rect 9498 -7178 9558 -6916
rect 10522 -6916 10528 -6362
rect 10562 -6362 10576 -6340
rect 11532 -6340 11592 -6190
rect 11828 -6247 12316 -6241
rect 11828 -6281 11840 -6247
rect 12304 -6281 12316 -6247
rect 11828 -6287 12316 -6281
rect 10562 -6916 10568 -6362
rect 11532 -6398 11546 -6340
rect 11540 -6886 11546 -6398
rect 10522 -6928 10568 -6916
rect 11534 -6916 11546 -6886
rect 11580 -6398 11592 -6340
rect 12548 -6340 12608 -5874
rect 14582 -5876 14588 -5816
rect 14648 -5876 14654 -5816
rect 15606 -6012 15666 -5660
rect 16622 -5660 16636 -5084
rect 16670 -5660 16682 -5084
rect 15900 -5719 16388 -5713
rect 15900 -5753 15912 -5719
rect 16376 -5753 16388 -5719
rect 15900 -5759 16388 -5753
rect 16116 -5814 16176 -5759
rect 16622 -5814 16682 -5660
rect 17638 -5084 17698 -4902
rect 18150 -4985 18210 -4902
rect 18654 -4930 18660 -4870
rect 18720 -4930 18726 -4870
rect 17936 -4991 18424 -4985
rect 17936 -5025 17948 -4991
rect 18412 -5025 18424 -4991
rect 17936 -5031 18424 -5025
rect 18150 -5038 18210 -5031
rect 17638 -5660 17654 -5084
rect 17688 -5660 17698 -5084
rect 18660 -5084 18720 -4930
rect 19160 -4985 19224 -4930
rect 20184 -4985 20248 -4812
rect 20688 -4930 20694 -4870
rect 20754 -4930 20760 -4870
rect 18954 -4991 19442 -4985
rect 18954 -5025 18966 -4991
rect 19430 -5025 19442 -4991
rect 18954 -5031 19442 -5025
rect 19972 -4991 20460 -4985
rect 19972 -5025 19984 -4991
rect 20448 -5025 20460 -4991
rect 19972 -5031 20460 -5025
rect 18660 -5112 18672 -5084
rect 16918 -5719 17406 -5713
rect 16918 -5753 16930 -5719
rect 17394 -5753 17406 -5719
rect 16918 -5759 17406 -5753
rect 17142 -5814 17202 -5759
rect 17638 -5814 17698 -5660
rect 18666 -5660 18672 -5112
rect 18706 -5112 18720 -5084
rect 19684 -5084 19730 -5072
rect 18706 -5660 18712 -5112
rect 19684 -5636 19690 -5084
rect 18666 -5672 18712 -5660
rect 19676 -5660 19690 -5636
rect 19724 -5636 19730 -5084
rect 20694 -5084 20754 -4930
rect 21196 -4985 21260 -4812
rect 21714 -4866 21774 -4628
rect 21714 -4926 22790 -4866
rect 20990 -4991 21478 -4985
rect 20990 -5025 21002 -4991
rect 21466 -5025 21478 -4991
rect 20990 -5031 21478 -5025
rect 20694 -5108 20708 -5084
rect 19724 -5660 19736 -5636
rect 17936 -5719 18424 -5713
rect 17936 -5753 17948 -5719
rect 18412 -5753 18424 -5719
rect 17936 -5759 18424 -5753
rect 18954 -5719 19442 -5713
rect 18954 -5753 18966 -5719
rect 19430 -5753 19442 -5719
rect 18954 -5759 19442 -5753
rect 18154 -5814 18214 -5759
rect 16116 -5874 18214 -5814
rect 15600 -6072 15606 -6012
rect 15666 -6072 15672 -6012
rect 13566 -6186 13572 -6126
rect 13632 -6186 13638 -6126
rect 15600 -6186 15606 -6126
rect 15666 -6186 15672 -6126
rect 12846 -6247 13334 -6241
rect 12846 -6281 12858 -6247
rect 13322 -6281 13334 -6247
rect 12846 -6287 13334 -6281
rect 12548 -6384 12564 -6340
rect 11580 -6886 11586 -6398
rect 12558 -6886 12564 -6384
rect 11580 -6916 11594 -6886
rect 9998 -6969 10058 -6968
rect 11004 -6969 11064 -6968
rect 9792 -6975 10280 -6969
rect 9792 -7009 9804 -6975
rect 10268 -7009 10280 -6975
rect 9792 -7015 10280 -7009
rect 10810 -6975 11298 -6969
rect 10810 -7009 10822 -6975
rect 11286 -7009 11298 -6975
rect 10810 -7015 11298 -7009
rect 9498 -7244 9558 -7238
rect 9492 -7442 9498 -7382
rect 9558 -7442 9564 -7382
rect 8774 -7503 9262 -7497
rect 8774 -7537 8786 -7503
rect 9250 -7537 9262 -7503
rect 8774 -7543 9262 -7537
rect 8478 -7618 8492 -7596
rect 7508 -8172 7514 -7630
rect 8486 -8144 8492 -7618
rect 7468 -8184 7514 -8172
rect 8480 -8172 8492 -8144
rect 8526 -7618 8538 -7596
rect 9498 -7596 9558 -7442
rect 9998 -7497 10058 -7015
rect 11004 -7497 11064 -7015
rect 11534 -7178 11594 -6916
rect 12550 -6916 12564 -6886
rect 12598 -6384 12608 -6340
rect 13572 -6340 13632 -6186
rect 13864 -6247 14352 -6241
rect 13864 -6281 13876 -6247
rect 14340 -6281 14352 -6247
rect 13864 -6287 14352 -6281
rect 14882 -6247 15370 -6241
rect 14882 -6281 14894 -6247
rect 15358 -6281 15370 -6247
rect 14882 -6287 15370 -6281
rect 13572 -6368 13582 -6340
rect 12598 -6886 12604 -6384
rect 12598 -6916 12610 -6886
rect 11828 -6975 12316 -6969
rect 11828 -7009 11840 -6975
rect 12304 -7009 12316 -6975
rect 11828 -7015 12316 -7009
rect 12054 -7070 12114 -7015
rect 12550 -7070 12610 -6916
rect 13576 -6916 13582 -6368
rect 13616 -6368 13632 -6340
rect 14594 -6340 14640 -6328
rect 13616 -6916 13622 -6368
rect 14594 -6892 14600 -6340
rect 13576 -6928 13622 -6916
rect 14588 -6916 14600 -6892
rect 14634 -6892 14640 -6340
rect 15606 -6340 15666 -6186
rect 15900 -6247 16388 -6241
rect 15900 -6281 15912 -6247
rect 16376 -6281 16388 -6247
rect 15900 -6287 16388 -6281
rect 16918 -6247 17406 -6241
rect 16918 -6281 16930 -6247
rect 17394 -6281 17406 -6247
rect 16918 -6287 17406 -6281
rect 15606 -6370 15618 -6340
rect 15612 -6888 15618 -6370
rect 14634 -6916 14648 -6892
rect 12846 -6975 13334 -6969
rect 12846 -7009 12858 -6975
rect 13322 -7009 13334 -6975
rect 12846 -7015 13334 -7009
rect 13864 -6975 14352 -6969
rect 13864 -7009 13876 -6975
rect 14340 -7009 14352 -6975
rect 13864 -7015 14352 -7009
rect 13066 -7070 13126 -7015
rect 12054 -7130 13126 -7070
rect 11528 -7238 11534 -7178
rect 11594 -7238 11600 -7178
rect 11526 -7340 11532 -7280
rect 11592 -7340 11598 -7280
rect 11532 -7382 11592 -7340
rect 11526 -7442 11532 -7382
rect 11592 -7442 11598 -7382
rect 9792 -7503 10280 -7497
rect 9792 -7537 9804 -7503
rect 10268 -7537 10280 -7503
rect 9792 -7543 10280 -7537
rect 10810 -7503 11298 -7497
rect 10810 -7537 10822 -7503
rect 11286 -7537 11298 -7503
rect 10810 -7543 11298 -7537
rect 8526 -8144 8532 -7618
rect 9498 -7620 9510 -7596
rect 8526 -8172 8540 -8144
rect 7756 -8231 8244 -8225
rect 7756 -8265 7768 -8231
rect 8232 -8265 8244 -8231
rect 7756 -8271 8244 -8265
rect 8480 -8330 8540 -8172
rect 9504 -8172 9510 -7620
rect 9544 -7620 9558 -7596
rect 10522 -7596 10568 -7584
rect 9544 -8172 9550 -7620
rect 10522 -8148 10528 -7596
rect 9504 -8184 9550 -8172
rect 10516 -8172 10528 -8148
rect 10562 -8148 10568 -7596
rect 11532 -7596 11592 -7442
rect 11828 -7503 12316 -7497
rect 11828 -7537 11840 -7503
rect 12304 -7537 12316 -7503
rect 11828 -7543 12316 -7537
rect 11532 -7624 11546 -7596
rect 10562 -8172 10576 -8148
rect 11540 -8153 11546 -7624
rect 8972 -8225 9032 -8218
rect 10010 -8225 10070 -8218
rect 8774 -8231 9262 -8225
rect 8774 -8265 8786 -8231
rect 9250 -8265 9262 -8231
rect 8774 -8271 9262 -8265
rect 9792 -8231 10280 -8225
rect 9792 -8265 9804 -8231
rect 10268 -8265 10280 -8231
rect 9792 -8271 10280 -8265
rect 8474 -8390 8480 -8330
rect 8540 -8390 8546 -8330
rect 7306 -8598 7312 -8538
rect 7372 -8598 7378 -8538
rect 7462 -8696 8538 -8636
rect 7462 -8852 7522 -8696
rect 7976 -8753 8036 -8696
rect 7756 -8759 8244 -8753
rect 7756 -8793 7768 -8759
rect 8232 -8793 8244 -8759
rect 7756 -8799 8244 -8793
rect 7462 -8890 7474 -8852
rect 7468 -9428 7474 -8890
rect 7508 -8890 7522 -8852
rect 8478 -8852 8538 -8696
rect 8972 -8753 9032 -8271
rect 9488 -8700 9494 -8640
rect 9554 -8700 9560 -8640
rect 8774 -8759 9262 -8753
rect 8774 -8793 8786 -8759
rect 9250 -8793 9262 -8759
rect 8774 -8799 9262 -8793
rect 8478 -8878 8492 -8852
rect 7508 -9428 7514 -8890
rect 8486 -9402 8492 -8878
rect 7468 -9440 7514 -9428
rect 8476 -9428 8492 -9402
rect 8526 -8878 8538 -8852
rect 9494 -8852 9554 -8700
rect 10010 -8753 10070 -8271
rect 10516 -8330 10576 -8172
rect 11534 -8172 11546 -8153
rect 11580 -7624 11592 -7596
rect 12550 -7596 12610 -7130
rect 13562 -7134 13568 -7074
rect 13628 -7134 13634 -7074
rect 12846 -7503 13334 -7497
rect 12846 -7537 12858 -7503
rect 13322 -7537 13334 -7503
rect 12846 -7543 13334 -7537
rect 11580 -8153 11586 -7624
rect 12550 -7634 12564 -7596
rect 12558 -8138 12564 -7634
rect 11580 -8172 11594 -8153
rect 11016 -8225 11076 -8218
rect 10810 -8231 11298 -8225
rect 10810 -8265 10822 -8231
rect 11286 -8265 11298 -8231
rect 10810 -8271 11298 -8265
rect 10510 -8390 10516 -8330
rect 10576 -8390 10582 -8330
rect 10516 -8438 10576 -8390
rect 10510 -8498 10516 -8438
rect 10576 -8498 10582 -8438
rect 11016 -8488 11076 -8271
rect 11534 -8322 11594 -8172
rect 12548 -8172 12564 -8138
rect 12598 -7634 12610 -7596
rect 13568 -7596 13628 -7134
rect 14070 -7236 14130 -7015
rect 14588 -7074 14648 -6916
rect 15606 -6916 15618 -6888
rect 15652 -6370 15666 -6340
rect 16630 -6340 16676 -6328
rect 15652 -6888 15658 -6370
rect 16630 -6888 16636 -6340
rect 15652 -6916 15666 -6888
rect 15100 -6969 15160 -6962
rect 14882 -6975 15370 -6969
rect 14882 -7009 14894 -6975
rect 15358 -7009 15370 -6975
rect 14882 -7015 15370 -7009
rect 14582 -7134 14588 -7074
rect 14648 -7134 14654 -7074
rect 15100 -7236 15160 -7015
rect 14070 -7296 15160 -7236
rect 14070 -7497 14130 -7296
rect 14582 -7440 14588 -7380
rect 14648 -7440 14654 -7380
rect 13864 -7503 14352 -7497
rect 13864 -7537 13876 -7503
rect 14340 -7537 14352 -7503
rect 13864 -7543 14352 -7537
rect 14070 -7548 14130 -7543
rect 13568 -7620 13582 -7596
rect 12598 -8138 12604 -7634
rect 12598 -8172 12608 -8138
rect 13576 -8142 13582 -7620
rect 11828 -8231 12316 -8225
rect 11828 -8265 11840 -8231
rect 12304 -8265 12316 -8231
rect 11828 -8271 12316 -8265
rect 12052 -8322 12112 -8271
rect 12548 -8322 12608 -8172
rect 13570 -8172 13582 -8142
rect 13616 -7620 13628 -7596
rect 14588 -7596 14648 -7440
rect 15100 -7497 15160 -7296
rect 15606 -7380 15666 -6916
rect 16624 -6916 16636 -6888
rect 16670 -6888 16676 -6340
rect 17638 -6340 17698 -5874
rect 18656 -6186 18662 -6126
rect 18722 -6186 18728 -6126
rect 17936 -6247 18424 -6241
rect 17936 -6281 17948 -6247
rect 18412 -6281 18424 -6247
rect 17936 -6287 18424 -6281
rect 17638 -6360 17654 -6340
rect 17648 -6888 17654 -6360
rect 16670 -6916 16684 -6888
rect 16112 -6969 16172 -6962
rect 15900 -6975 16388 -6969
rect 15900 -7009 15912 -6975
rect 16376 -7009 16388 -6975
rect 15900 -7015 16388 -7009
rect 15600 -7440 15606 -7380
rect 15666 -7440 15672 -7380
rect 16112 -7497 16172 -7015
rect 16624 -7074 16684 -6916
rect 17638 -6916 17654 -6888
rect 17688 -6360 17698 -6340
rect 18662 -6340 18722 -6186
rect 19162 -6241 19222 -5759
rect 19676 -5818 19736 -5660
rect 20702 -5660 20708 -5108
rect 20742 -5108 20754 -5084
rect 21714 -5084 21774 -4926
rect 22228 -4985 22288 -4926
rect 22008 -4991 22496 -4985
rect 22008 -5025 22020 -4991
rect 22484 -5025 22496 -4991
rect 22008 -5031 22496 -5025
rect 20742 -5660 20748 -5108
rect 21714 -5120 21726 -5084
rect 21720 -5632 21726 -5120
rect 20702 -5672 20748 -5660
rect 21712 -5660 21726 -5632
rect 21760 -5120 21774 -5084
rect 22730 -5084 22790 -4926
rect 22730 -5108 22744 -5084
rect 21760 -5632 21766 -5120
rect 21760 -5660 21772 -5632
rect 21192 -5713 21252 -5707
rect 19972 -5719 20460 -5713
rect 19972 -5753 19984 -5719
rect 20448 -5753 20460 -5719
rect 19972 -5759 20460 -5753
rect 20990 -5719 21478 -5713
rect 20990 -5753 21002 -5719
rect 21466 -5753 21478 -5719
rect 20990 -5759 21478 -5753
rect 19670 -5878 19676 -5818
rect 19736 -5878 19742 -5818
rect 20186 -6241 20246 -5759
rect 20690 -6186 20696 -6126
rect 20756 -6186 20762 -6126
rect 18954 -6247 19442 -6241
rect 18954 -6281 18966 -6247
rect 19430 -6281 19442 -6247
rect 18954 -6287 19442 -6281
rect 19972 -6247 20460 -6241
rect 19972 -6281 19984 -6247
rect 20448 -6281 20460 -6247
rect 19972 -6287 20460 -6281
rect 17688 -6888 17694 -6360
rect 18662 -6368 18672 -6340
rect 17688 -6916 17698 -6888
rect 16918 -6975 17406 -6969
rect 16918 -7009 16930 -6975
rect 17394 -7009 17406 -6975
rect 16918 -7015 17406 -7009
rect 17142 -7072 17202 -7015
rect 17638 -7072 17698 -6916
rect 18666 -6916 18672 -6368
rect 18706 -6368 18722 -6340
rect 19684 -6340 19730 -6328
rect 18706 -6916 18712 -6368
rect 19684 -6880 19690 -6340
rect 18666 -6928 18712 -6916
rect 19674 -6916 19690 -6880
rect 19724 -6880 19730 -6340
rect 20696 -6340 20756 -6186
rect 21192 -6241 21252 -5759
rect 21712 -5818 21772 -5660
rect 22738 -5660 22744 -5108
rect 22778 -5108 22790 -5084
rect 22778 -5660 22784 -5108
rect 22738 -5672 22784 -5660
rect 22008 -5719 22496 -5713
rect 22008 -5753 22020 -5719
rect 22484 -5753 22496 -5719
rect 22008 -5759 22496 -5753
rect 21706 -5878 21712 -5818
rect 21772 -5878 21778 -5818
rect 21714 -6180 22790 -6120
rect 20990 -6247 21478 -6241
rect 20990 -6281 21002 -6247
rect 21466 -6281 21478 -6247
rect 20990 -6287 21478 -6281
rect 20696 -6364 20708 -6340
rect 19724 -6916 19734 -6880
rect 20702 -6888 20708 -6364
rect 19156 -6969 19216 -6968
rect 17936 -6975 18424 -6969
rect 17936 -7009 17948 -6975
rect 18412 -7009 18424 -6975
rect 17936 -7015 18424 -7009
rect 18954 -6975 19442 -6969
rect 18954 -7009 18966 -6975
rect 19430 -7009 19442 -6975
rect 18954 -7015 19442 -7009
rect 18154 -7072 18214 -7015
rect 16618 -7134 16624 -7074
rect 16684 -7134 16690 -7074
rect 17142 -7132 18214 -7072
rect 16616 -7440 16622 -7380
rect 16682 -7440 16688 -7380
rect 14882 -7503 15370 -7497
rect 14882 -7537 14894 -7503
rect 15358 -7537 15370 -7503
rect 14882 -7543 15370 -7537
rect 15900 -7503 16388 -7497
rect 15900 -7537 15912 -7503
rect 16376 -7537 16388 -7503
rect 15900 -7543 16388 -7537
rect 14588 -7618 14600 -7596
rect 13616 -8142 13622 -7620
rect 13616 -8172 13630 -8142
rect 12846 -8231 13334 -8225
rect 12846 -8265 12858 -8231
rect 13322 -8265 13334 -8231
rect 12846 -8271 13334 -8265
rect 13064 -8322 13124 -8271
rect 11528 -8382 11534 -8322
rect 11594 -8382 11600 -8322
rect 12052 -8382 13124 -8322
rect 13330 -8382 13336 -8322
rect 13396 -8382 13402 -8322
rect 13570 -8328 13630 -8172
rect 14594 -8172 14600 -7618
rect 14634 -7618 14648 -7596
rect 15612 -7596 15658 -7584
rect 14634 -8172 14640 -7618
rect 15612 -8146 15618 -7596
rect 14594 -8184 14640 -8172
rect 15606 -8172 15618 -8146
rect 15652 -8146 15658 -7596
rect 16622 -7596 16682 -7440
rect 16918 -7503 17406 -7497
rect 16918 -7537 16930 -7503
rect 17394 -7537 17406 -7503
rect 16918 -7543 17406 -7537
rect 16622 -7622 16636 -7596
rect 15652 -8172 15666 -8146
rect 13864 -8231 14352 -8225
rect 13864 -8265 13876 -8231
rect 14340 -8265 14352 -8231
rect 13864 -8271 14352 -8265
rect 14882 -8231 15370 -8225
rect 14882 -8265 14894 -8231
rect 15358 -8265 15370 -8231
rect 14882 -8271 15370 -8265
rect 11016 -8548 11792 -8488
rect 11016 -8753 11076 -8548
rect 11522 -8700 11528 -8640
rect 11588 -8700 11594 -8640
rect 11732 -8652 11792 -8548
rect 9792 -8759 10280 -8753
rect 9792 -8793 9804 -8759
rect 10268 -8793 10280 -8759
rect 9792 -8799 10280 -8793
rect 10810 -8759 11298 -8753
rect 10810 -8793 10822 -8759
rect 11286 -8793 11298 -8759
rect 10810 -8799 11298 -8793
rect 9494 -8878 9510 -8852
rect 8526 -9402 8532 -8878
rect 8526 -9428 8536 -9402
rect 7756 -9487 8244 -9481
rect 7756 -9521 7768 -9487
rect 8232 -9521 8244 -9487
rect 7756 -9527 8244 -9521
rect 8476 -9588 8536 -9428
rect 9504 -9428 9510 -8878
rect 9544 -8878 9554 -8852
rect 10522 -8852 10568 -8840
rect 9544 -9428 9550 -8878
rect 10522 -9406 10528 -8852
rect 9504 -9440 9550 -9428
rect 10512 -9428 10528 -9406
rect 10562 -9406 10568 -8852
rect 11528 -8852 11588 -8700
rect 11726 -8712 11732 -8652
rect 11792 -8712 11798 -8652
rect 11828 -8759 12316 -8753
rect 11828 -8793 11840 -8759
rect 12304 -8793 12316 -8759
rect 11828 -8799 12316 -8793
rect 11528 -8882 11546 -8852
rect 11540 -9392 11546 -8882
rect 10562 -9428 10572 -9406
rect 8774 -9487 9262 -9481
rect 8774 -9521 8786 -9487
rect 9250 -9521 9262 -9487
rect 8774 -9527 9262 -9521
rect 9792 -9487 10280 -9481
rect 9792 -9521 9804 -9487
rect 10268 -9521 10280 -9487
rect 9792 -9527 10280 -9521
rect 8470 -9648 8476 -9588
rect 8536 -9648 8542 -9588
rect 8984 -9702 9044 -9527
rect 10008 -9702 10068 -9527
rect 10512 -9588 10572 -9428
rect 11534 -9428 11546 -9392
rect 11580 -8882 11588 -8852
rect 12548 -8852 12608 -8382
rect 13336 -8592 13396 -8382
rect 13564 -8388 13570 -8328
rect 13630 -8388 13636 -8328
rect 14066 -8450 14126 -8271
rect 15094 -8450 15154 -8271
rect 15606 -8328 15666 -8172
rect 16630 -8172 16636 -7622
rect 16670 -7622 16682 -7596
rect 17638 -7596 17698 -7132
rect 18652 -7238 18658 -7178
rect 18718 -7238 18724 -7178
rect 17936 -7503 18424 -7497
rect 17936 -7537 17948 -7503
rect 18412 -7537 18424 -7503
rect 17936 -7543 18424 -7537
rect 16670 -8172 16676 -7622
rect 17638 -7626 17654 -7596
rect 17648 -8140 17654 -7626
rect 16630 -8184 16676 -8172
rect 17636 -8172 17654 -8140
rect 17688 -7626 17698 -7596
rect 18658 -7596 18718 -7238
rect 19156 -7497 19216 -7015
rect 19520 -7120 19526 -7060
rect 19586 -7120 19592 -7060
rect 19526 -7380 19586 -7120
rect 19674 -7170 19734 -6916
rect 20694 -6916 20708 -6888
rect 20742 -6364 20756 -6340
rect 21714 -6340 21774 -6180
rect 22228 -6241 22288 -6180
rect 22008 -6247 22496 -6241
rect 22008 -6281 22020 -6247
rect 22484 -6281 22496 -6247
rect 22008 -6287 22496 -6281
rect 20742 -6888 20748 -6364
rect 21714 -6374 21726 -6340
rect 21720 -6876 21726 -6374
rect 20742 -6916 20754 -6888
rect 20180 -6969 20240 -6968
rect 19972 -6975 20460 -6969
rect 19972 -7009 19984 -6975
rect 20448 -7009 20460 -6975
rect 19972 -7015 20460 -7009
rect 19668 -7230 19674 -7170
rect 19734 -7230 19740 -7170
rect 19520 -7440 19526 -7380
rect 19586 -7440 19592 -7380
rect 19672 -7438 19678 -7378
rect 19738 -7438 19744 -7378
rect 18954 -7503 19442 -7497
rect 18954 -7537 18966 -7503
rect 19430 -7537 19442 -7503
rect 18954 -7543 19442 -7537
rect 17688 -8140 17694 -7626
rect 18658 -7628 18672 -7596
rect 18666 -8140 18672 -7628
rect 17688 -8172 17696 -8140
rect 15900 -8231 16388 -8225
rect 15900 -8265 15912 -8231
rect 16376 -8265 16388 -8231
rect 15900 -8271 16388 -8265
rect 16918 -8231 17406 -8225
rect 16918 -8265 16930 -8231
rect 17394 -8265 17406 -8231
rect 16918 -8271 17406 -8265
rect 15600 -8388 15606 -8328
rect 15666 -8388 15672 -8328
rect 14066 -8510 15154 -8450
rect 15598 -8498 15604 -8438
rect 15664 -8498 15670 -8438
rect 13336 -8652 14644 -8592
rect 12846 -8759 13334 -8753
rect 12846 -8793 12858 -8759
rect 13322 -8793 13334 -8759
rect 12846 -8799 13334 -8793
rect 13864 -8759 14352 -8753
rect 13864 -8793 13876 -8759
rect 14340 -8793 14352 -8759
rect 13864 -8799 14352 -8793
rect 11580 -9392 11586 -8882
rect 12548 -8910 12564 -8852
rect 11580 -9428 11594 -9392
rect 12558 -9396 12564 -8910
rect 10810 -9487 11298 -9481
rect 10810 -9521 10822 -9487
rect 11286 -9521 11298 -9487
rect 10810 -9527 11298 -9521
rect 10506 -9648 10512 -9588
rect 10572 -9648 10578 -9588
rect 11014 -9702 11074 -9527
rect 7174 -9778 7180 -9718
rect 7240 -9778 7246 -9718
rect 8984 -9762 11074 -9702
rect 2332 -9906 2336 -9846
rect 2396 -9906 6858 -9846
rect 2336 -9912 2396 -9906
rect 2216 -9964 2276 -9958
rect 7180 -9964 7240 -9778
rect 2276 -10024 7240 -9964
rect 2216 -10030 2276 -10024
rect 1770 -10082 1830 -10076
rect 8984 -10082 9044 -9762
rect 11014 -9972 11074 -9762
rect 11534 -9858 11594 -9428
rect 12548 -9428 12564 -9396
rect 12598 -8910 12608 -8852
rect 13576 -8852 13622 -8840
rect 12598 -9396 12604 -8910
rect 13576 -9384 13582 -8852
rect 12598 -9428 12608 -9396
rect 11828 -9487 12316 -9481
rect 11828 -9521 11840 -9487
rect 12304 -9521 12316 -9487
rect 11828 -9527 12316 -9521
rect 12052 -9582 12112 -9527
rect 12548 -9582 12608 -9428
rect 13570 -9428 13582 -9384
rect 13616 -9384 13622 -8852
rect 14584 -8852 14644 -8652
rect 15094 -8652 15154 -8510
rect 15094 -8753 15154 -8712
rect 14882 -8759 15370 -8753
rect 14882 -8793 14894 -8759
rect 15358 -8793 15370 -8759
rect 14882 -8799 15370 -8793
rect 14584 -8904 14600 -8852
rect 13616 -9428 13630 -9384
rect 12846 -9487 13334 -9481
rect 12846 -9521 12858 -9487
rect 13322 -9521 13334 -9487
rect 12846 -9527 13334 -9521
rect 13064 -9582 13124 -9527
rect 13570 -9582 13630 -9428
rect 14594 -9428 14600 -8904
rect 14634 -8904 14644 -8852
rect 15604 -8852 15664 -8498
rect 16110 -8652 16170 -8271
rect 17140 -8324 17200 -8271
rect 17636 -8324 17696 -8172
rect 18660 -8172 18672 -8140
rect 18706 -7628 18718 -7596
rect 19678 -7596 19738 -7438
rect 20180 -7497 20240 -7015
rect 20694 -7280 20754 -6916
rect 21714 -6916 21726 -6876
rect 21760 -6374 21774 -6340
rect 22730 -6340 22790 -6180
rect 22730 -6362 22744 -6340
rect 21760 -6876 21766 -6374
rect 21760 -6916 21774 -6876
rect 21186 -6969 21246 -6962
rect 20990 -6975 21478 -6969
rect 20990 -7009 21002 -6975
rect 21466 -7009 21478 -6975
rect 20990 -7015 21478 -7009
rect 20688 -7340 20694 -7280
rect 20754 -7340 20760 -7280
rect 21186 -7497 21246 -7015
rect 21714 -7170 21774 -6916
rect 22738 -6916 22744 -6362
rect 22778 -6362 22790 -6340
rect 22778 -6916 22784 -6362
rect 22738 -6928 22784 -6916
rect 22008 -6975 22496 -6969
rect 22008 -7009 22020 -6975
rect 22484 -7009 22496 -6975
rect 22008 -7015 22496 -7009
rect 22854 -7170 22914 -4402
rect 22996 -4570 23056 -1854
rect 23284 -4270 23290 -4210
rect 23350 -4270 23356 -4210
rect 22996 -4636 23056 -4630
rect 23132 -4930 23138 -4870
rect 23198 -4930 23204 -4870
rect 22972 -6072 22978 -6012
rect 23038 -6072 23044 -6012
rect 21708 -7230 21714 -7170
rect 21774 -7230 21780 -7170
rect 22848 -7230 22854 -7170
rect 22914 -7230 22920 -7170
rect 21706 -7438 21712 -7378
rect 21772 -7438 21778 -7378
rect 19972 -7503 20460 -7497
rect 19972 -7537 19984 -7503
rect 20448 -7537 20460 -7503
rect 19972 -7543 20460 -7537
rect 20990 -7503 21478 -7497
rect 20990 -7537 21002 -7503
rect 21466 -7537 21478 -7503
rect 20990 -7543 21478 -7537
rect 19678 -7616 19690 -7596
rect 18706 -8140 18712 -7628
rect 18706 -8172 18720 -8140
rect 17936 -8231 18424 -8225
rect 17936 -8265 17948 -8231
rect 18412 -8265 18424 -8231
rect 17936 -8271 18424 -8265
rect 18152 -8324 18212 -8271
rect 17140 -8384 18212 -8324
rect 18660 -8326 18720 -8172
rect 19684 -8172 19690 -7616
rect 19724 -7616 19738 -7596
rect 20702 -7596 20748 -7584
rect 19724 -8172 19730 -7616
rect 20702 -8144 20708 -7596
rect 19684 -8184 19730 -8172
rect 20696 -8172 20708 -8144
rect 20742 -8144 20748 -7596
rect 21712 -7596 21772 -7438
rect 22008 -7503 22496 -7497
rect 22008 -7537 22020 -7503
rect 22484 -7537 22496 -7503
rect 22008 -7543 22496 -7537
rect 21712 -7620 21726 -7596
rect 21720 -8136 21726 -7620
rect 20742 -8172 20756 -8144
rect 19168 -8225 19228 -8218
rect 20192 -8225 20252 -8218
rect 18954 -8231 19442 -8225
rect 18954 -8265 18966 -8231
rect 19430 -8265 19442 -8231
rect 18954 -8271 19442 -8265
rect 19972 -8231 20460 -8225
rect 19972 -8265 19984 -8231
rect 20448 -8265 20460 -8231
rect 19972 -8271 20460 -8265
rect 16110 -8718 16170 -8712
rect 15900 -8759 16388 -8753
rect 15900 -8793 15912 -8759
rect 16376 -8793 16388 -8759
rect 15900 -8799 16388 -8793
rect 16918 -8759 17406 -8753
rect 16918 -8793 16930 -8759
rect 17394 -8793 17406 -8759
rect 16918 -8799 17406 -8793
rect 14634 -9428 14640 -8904
rect 15604 -8916 15618 -8852
rect 14594 -9440 14640 -9428
rect 15612 -9428 15618 -8916
rect 15652 -8916 15664 -8852
rect 16630 -8852 16676 -8840
rect 15652 -9428 15658 -8916
rect 16630 -9400 16636 -8852
rect 15612 -9440 15658 -9428
rect 16622 -9428 16636 -9400
rect 16670 -9400 16676 -8852
rect 17636 -8852 17696 -8384
rect 18654 -8386 18660 -8326
rect 18720 -8386 18726 -8326
rect 19168 -8646 19228 -8271
rect 19168 -8652 19230 -8646
rect 19168 -8712 19170 -8652
rect 19676 -8700 19682 -8640
rect 19742 -8700 19748 -8640
rect 19168 -8718 19230 -8712
rect 19168 -8753 19228 -8718
rect 17936 -8759 18424 -8753
rect 17936 -8793 17948 -8759
rect 18412 -8793 18424 -8759
rect 17936 -8799 18424 -8793
rect 18954 -8759 19442 -8753
rect 18954 -8793 18966 -8759
rect 19430 -8793 19442 -8759
rect 18954 -8799 19442 -8793
rect 17636 -8890 17654 -8852
rect 17648 -9398 17654 -8890
rect 16670 -9428 16682 -9400
rect 13864 -9487 14352 -9481
rect 13864 -9521 13876 -9487
rect 14340 -9521 14352 -9487
rect 13864 -9527 14352 -9521
rect 14882 -9487 15370 -9481
rect 14882 -9521 14894 -9487
rect 15358 -9521 15370 -9487
rect 14882 -9527 15370 -9521
rect 15900 -9487 16388 -9481
rect 15900 -9521 15912 -9487
rect 16376 -9521 16388 -9487
rect 15900 -9527 16388 -9521
rect 14080 -9582 14140 -9527
rect 16106 -9582 16166 -9527
rect 16622 -9582 16682 -9428
rect 17636 -9428 17654 -9398
rect 17688 -8890 17696 -8852
rect 18666 -8852 18712 -8840
rect 17688 -9398 17694 -8890
rect 17688 -9428 17696 -9398
rect 18666 -9402 18672 -8852
rect 16918 -9487 17406 -9481
rect 16918 -9521 16930 -9487
rect 17394 -9521 17406 -9487
rect 16918 -9527 17406 -9521
rect 17140 -9582 17200 -9527
rect 17636 -9582 17696 -9428
rect 18664 -9428 18672 -9402
rect 18706 -9402 18712 -8852
rect 19682 -8852 19742 -8700
rect 20192 -8753 20252 -8271
rect 20696 -8326 20756 -8172
rect 21712 -8172 21726 -8136
rect 21760 -7620 21772 -7596
rect 22738 -7596 22784 -7584
rect 21760 -8136 21766 -7620
rect 21760 -8172 21772 -8136
rect 22738 -8148 22744 -7596
rect 21198 -8225 21258 -8212
rect 20990 -8231 21478 -8225
rect 20990 -8265 21002 -8231
rect 21466 -8265 21478 -8231
rect 20990 -8271 21478 -8265
rect 20690 -8386 20696 -8326
rect 20756 -8386 20762 -8326
rect 21198 -8753 21258 -8271
rect 21712 -8330 21772 -8172
rect 22728 -8172 22744 -8148
rect 22778 -8148 22784 -7596
rect 22778 -8172 22788 -8148
rect 22008 -8231 22496 -8225
rect 22008 -8265 22020 -8231
rect 22484 -8265 22496 -8231
rect 22008 -8271 22496 -8265
rect 22226 -8330 22286 -8271
rect 22728 -8330 22788 -8172
rect 21712 -8390 22788 -8330
rect 22854 -8438 22914 -7230
rect 22978 -7378 23038 -6072
rect 22972 -7438 22978 -7378
rect 23038 -7438 23044 -7378
rect 22848 -8498 22854 -8438
rect 22914 -8498 22920 -8438
rect 21710 -8700 21716 -8640
rect 21776 -8700 21782 -8640
rect 19972 -8759 20460 -8753
rect 19972 -8793 19984 -8759
rect 20448 -8793 20460 -8759
rect 19972 -8799 20460 -8793
rect 20990 -8759 21478 -8753
rect 20990 -8793 21002 -8759
rect 21466 -8793 21478 -8759
rect 20990 -8799 21478 -8793
rect 19682 -8878 19690 -8852
rect 18706 -9428 18724 -9402
rect 17936 -9487 18424 -9481
rect 17936 -9521 17948 -9487
rect 18412 -9521 18424 -9487
rect 17936 -9527 18424 -9521
rect 18152 -9582 18212 -9527
rect 12052 -9642 18212 -9582
rect 18664 -9588 18724 -9428
rect 19684 -9428 19690 -8878
rect 19724 -8878 19742 -8852
rect 20702 -8852 20748 -8840
rect 19724 -9428 19730 -8878
rect 20702 -9406 20708 -8852
rect 19684 -9440 19730 -9428
rect 20700 -9428 20708 -9406
rect 20742 -9406 20748 -8852
rect 21716 -8852 21776 -8700
rect 22008 -8759 22496 -8753
rect 22008 -8793 22020 -8759
rect 22484 -8793 22496 -8759
rect 22008 -8799 22496 -8793
rect 21716 -8882 21726 -8852
rect 21720 -9390 21726 -8882
rect 20742 -9428 20760 -9406
rect 19172 -9481 19232 -9474
rect 18954 -9487 19442 -9481
rect 18954 -9521 18966 -9487
rect 19430 -9521 19442 -9487
rect 18954 -9527 19442 -9521
rect 19972 -9487 20460 -9481
rect 19972 -9521 19984 -9487
rect 20448 -9521 20460 -9487
rect 19972 -9527 20460 -9521
rect 18658 -9648 18664 -9588
rect 18724 -9648 18730 -9588
rect 19172 -9700 19232 -9527
rect 20192 -9700 20252 -9527
rect 20700 -9588 20760 -9428
rect 21714 -9428 21726 -9390
rect 21760 -8882 21776 -8852
rect 22738 -8852 22784 -8840
rect 21760 -9390 21766 -8882
rect 21760 -9428 21774 -9390
rect 22738 -9402 22744 -8852
rect 20990 -9487 21478 -9481
rect 20990 -9521 21002 -9487
rect 21466 -9521 21478 -9487
rect 20990 -9527 21478 -9521
rect 20694 -9648 20700 -9588
rect 20760 -9648 20766 -9588
rect 21194 -9700 21254 -9527
rect 21714 -9584 21774 -9428
rect 22730 -9428 22744 -9402
rect 22778 -9402 22784 -8852
rect 22778 -9428 22790 -9402
rect 22008 -9487 22496 -9481
rect 22008 -9521 22020 -9487
rect 22484 -9521 22496 -9487
rect 22008 -9527 22496 -9521
rect 22228 -9584 22288 -9527
rect 22730 -9584 22790 -9428
rect 21714 -9644 22790 -9584
rect 19172 -9760 21254 -9700
rect 11528 -9918 11534 -9858
rect 11594 -9918 11600 -9858
rect 19172 -9972 19232 -9760
rect 23138 -9858 23198 -4930
rect 23290 -6126 23350 -4270
rect 23284 -6186 23290 -6126
rect 23350 -6186 23356 -6126
rect 24716 -9728 24722 3702
rect 24822 -9728 24828 3702
rect 23132 -9918 23138 -9858
rect 23198 -9918 23204 -9858
rect 11014 -10032 19232 -9972
rect 1830 -10142 9044 -10082
rect 1770 -10148 1830 -10142
rect 24716 -10242 24828 -9728
rect 372 -10248 24828 -10242
rect 372 -10348 478 -10248
rect 24722 -10348 24828 -10248
rect 372 -10354 24828 -10348
rect -2866 -10670 -2722 -10378
rect -13992 -10978 -2722 -10670
rect -13992 -11172 -1640 -10978
rect -13992 -11178 24928 -11172
rect -13992 -11278 -12222 -11178
rect 24822 -11278 24928 -11178
rect -13992 -11284 24928 -11278
rect -13992 -11300 -1642 -11284
rect -12328 -12070 -12216 -11300
rect 1888 -11358 1948 -11352
rect 2210 -11408 2216 -11348
rect 2276 -11408 2282 -11348
rect 2336 -11356 2396 -11350
rect 1276 -11554 1282 -11494
rect 1342 -11554 1348 -11494
rect 1396 -11552 1402 -11492
rect 1462 -11552 1468 -11492
rect 1536 -11534 1542 -11474
rect 1602 -11534 1608 -11474
rect 1764 -11518 1770 -11458
rect 1830 -11518 1836 -11458
rect 1144 -11682 1150 -11622
rect 1210 -11682 1216 -11622
rect -12328 -26330 -12322 -12070
rect -12222 -26330 -12216 -12070
rect -1568 -12280 -1562 -12220
rect -1502 -12280 -1496 -12220
rect -1562 -12324 -1502 -12280
rect -9196 -12384 -1502 -12324
rect -9196 -12524 -9136 -12384
rect -8686 -12434 -8626 -12384
rect -8902 -12440 -8414 -12434
rect -8902 -12474 -8890 -12440
rect -8426 -12474 -8414 -12440
rect -8902 -12480 -8414 -12474
rect -9196 -12554 -9184 -12524
rect -9190 -13082 -9184 -12554
rect -9200 -13100 -9184 -13082
rect -9150 -12554 -9136 -12524
rect -8180 -12524 -8120 -12384
rect -7678 -12434 -7618 -12384
rect -6650 -12434 -6590 -12384
rect -7884 -12440 -7396 -12434
rect -7884 -12474 -7872 -12440
rect -7408 -12474 -7396 -12440
rect -7884 -12480 -7396 -12474
rect -6866 -12440 -6378 -12434
rect -6866 -12474 -6854 -12440
rect -6390 -12474 -6378 -12440
rect -6866 -12480 -6378 -12474
rect -8180 -12548 -8166 -12524
rect -9150 -13082 -9144 -12554
rect -8172 -13078 -8166 -12548
rect -9150 -13100 -9140 -13082
rect -9200 -13342 -9140 -13100
rect -8180 -13100 -8166 -13078
rect -8132 -12548 -8120 -12524
rect -7154 -12524 -7108 -12512
rect -8132 -13078 -8126 -12548
rect -7154 -13076 -7148 -12524
rect -8132 -13100 -8120 -13078
rect -8902 -13150 -8414 -13144
rect -8902 -13184 -8890 -13150
rect -8426 -13184 -8414 -13150
rect -8902 -13190 -8414 -13184
rect -8686 -13252 -8626 -13190
rect -8902 -13258 -8414 -13252
rect -8902 -13292 -8890 -13258
rect -8426 -13292 -8414 -13258
rect -8902 -13298 -8414 -13292
rect -9200 -13372 -9184 -13342
rect -9190 -13896 -9184 -13372
rect -9198 -13918 -9184 -13896
rect -9150 -13372 -9140 -13342
rect -8180 -13342 -8120 -13100
rect -7160 -13100 -7148 -13076
rect -7114 -13076 -7108 -12524
rect -6142 -12524 -6082 -12384
rect -5636 -12434 -5576 -12384
rect -4622 -12434 -4562 -12384
rect -5848 -12440 -5360 -12434
rect -5848 -12474 -5836 -12440
rect -5372 -12474 -5360 -12440
rect -5848 -12480 -5360 -12474
rect -4830 -12440 -4342 -12434
rect -4830 -12474 -4818 -12440
rect -4354 -12474 -4342 -12440
rect -4830 -12480 -4342 -12474
rect -6142 -12562 -6130 -12524
rect -7114 -13100 -7100 -13076
rect -6136 -13080 -6130 -12562
rect -7884 -13150 -7396 -13144
rect -7884 -13184 -7872 -13150
rect -7408 -13184 -7396 -13150
rect -7884 -13190 -7396 -13184
rect -7682 -13252 -7622 -13190
rect -7884 -13258 -7396 -13252
rect -7884 -13292 -7872 -13258
rect -7408 -13292 -7396 -13258
rect -7884 -13298 -7396 -13292
rect -8180 -13368 -8166 -13342
rect -9150 -13896 -9144 -13372
rect -8172 -13892 -8166 -13368
rect -9150 -13918 -9138 -13896
rect -9198 -14160 -9138 -13918
rect -8178 -13918 -8166 -13892
rect -8132 -13368 -8120 -13342
rect -7160 -13342 -7100 -13100
rect -6142 -13100 -6130 -13080
rect -6096 -12562 -6082 -12524
rect -5118 -12524 -5072 -12512
rect -4106 -12524 -4046 -12384
rect -3590 -12434 -3530 -12384
rect -2584 -12434 -2524 -12384
rect -3812 -12440 -3324 -12434
rect -3812 -12474 -3800 -12440
rect -3336 -12474 -3324 -12440
rect -3812 -12480 -3324 -12474
rect -2794 -12440 -2306 -12434
rect -2794 -12474 -2782 -12440
rect -2318 -12474 -2306 -12440
rect -2794 -12480 -2306 -12474
rect -6096 -13080 -6090 -12562
rect -5118 -13072 -5112 -12524
rect -6096 -13100 -6082 -13080
rect -6866 -13150 -6378 -13144
rect -6866 -13184 -6854 -13150
rect -6390 -13184 -6378 -13150
rect -6866 -13190 -6378 -13184
rect -6652 -13252 -6592 -13190
rect -6866 -13258 -6378 -13252
rect -6866 -13292 -6854 -13258
rect -6390 -13292 -6378 -13258
rect -6866 -13298 -6378 -13292
rect -7160 -13366 -7148 -13342
rect -8132 -13892 -8126 -13368
rect -7154 -13890 -7148 -13366
rect -8132 -13918 -8118 -13892
rect -8902 -13968 -8414 -13962
rect -8902 -14002 -8890 -13968
rect -8426 -14002 -8414 -13968
rect -8902 -14008 -8414 -14002
rect -8686 -14070 -8626 -14008
rect -8902 -14076 -8414 -14070
rect -8902 -14110 -8890 -14076
rect -8426 -14110 -8414 -14076
rect -8902 -14116 -8414 -14110
rect -9198 -14186 -9184 -14160
rect -9190 -14724 -9184 -14186
rect -9198 -14736 -9184 -14724
rect -9150 -14186 -9138 -14160
rect -8178 -14160 -8118 -13918
rect -7158 -13918 -7148 -13890
rect -7114 -13366 -7100 -13342
rect -6142 -13342 -6082 -13100
rect -5122 -13100 -5112 -13072
rect -5078 -13072 -5072 -12524
rect -4108 -12558 -4094 -12524
rect -4106 -12570 -4094 -12558
rect -5078 -13100 -5062 -13072
rect -4100 -13080 -4094 -12570
rect -5848 -13150 -5360 -13144
rect -5848 -13184 -5836 -13150
rect -5372 -13184 -5360 -13150
rect -5848 -13190 -5360 -13184
rect -5650 -13252 -5590 -13190
rect -5848 -13258 -5360 -13252
rect -5848 -13292 -5836 -13258
rect -5372 -13292 -5360 -13258
rect -5848 -13298 -5360 -13292
rect -7114 -13890 -7108 -13366
rect -6142 -13370 -6130 -13342
rect -7114 -13918 -7098 -13890
rect -6136 -13894 -6130 -13370
rect -7884 -13968 -7396 -13962
rect -7884 -14002 -7872 -13968
rect -7408 -14002 -7396 -13968
rect -7884 -14008 -7396 -14002
rect -7670 -14070 -7610 -14008
rect -7884 -14076 -7396 -14070
rect -7884 -14110 -7872 -14076
rect -7408 -14110 -7396 -14076
rect -7884 -14116 -7396 -14110
rect -8178 -14182 -8166 -14160
rect -9150 -14724 -9144 -14186
rect -8172 -14720 -8166 -14182
rect -9150 -14736 -9138 -14724
rect -9198 -14978 -9138 -14736
rect -8178 -14736 -8166 -14720
rect -8132 -14182 -8118 -14160
rect -7158 -14160 -7098 -13918
rect -6140 -13918 -6130 -13894
rect -6096 -13370 -6082 -13342
rect -5122 -13342 -5062 -13100
rect -4110 -13100 -4094 -13080
rect -4060 -12570 -4046 -12524
rect -3082 -12524 -3036 -12512
rect -4060 -13080 -4054 -12570
rect -3082 -13080 -3076 -12524
rect -4060 -13100 -4050 -13080
rect -4830 -13150 -4342 -13144
rect -4830 -13184 -4818 -13150
rect -4354 -13184 -4342 -13150
rect -4830 -13190 -4342 -13184
rect -4620 -13252 -4560 -13190
rect -4830 -13258 -4342 -13252
rect -4830 -13292 -4818 -13258
rect -4354 -13292 -4342 -13258
rect -4830 -13298 -4342 -13292
rect -5122 -13362 -5112 -13342
rect -6096 -13894 -6090 -13370
rect -5118 -13886 -5112 -13362
rect -6096 -13918 -6080 -13894
rect -6866 -13968 -6378 -13962
rect -6866 -14002 -6854 -13968
rect -6390 -14002 -6378 -13968
rect -6866 -14008 -6378 -14002
rect -6652 -14070 -6592 -14008
rect -6866 -14076 -6378 -14070
rect -6866 -14110 -6854 -14076
rect -6390 -14110 -6378 -14076
rect -6866 -14116 -6378 -14110
rect -7158 -14180 -7148 -14160
rect -8132 -14720 -8126 -14182
rect -7154 -14718 -7148 -14180
rect -8132 -14736 -8118 -14720
rect -8902 -14786 -8414 -14780
rect -8902 -14820 -8890 -14786
rect -8426 -14820 -8414 -14786
rect -8902 -14826 -8414 -14820
rect -8692 -14888 -8632 -14826
rect -8902 -14894 -8414 -14888
rect -8902 -14928 -8890 -14894
rect -8426 -14928 -8414 -14894
rect -8902 -14934 -8414 -14928
rect -9198 -15014 -9184 -14978
rect -9190 -15536 -9184 -15014
rect -9198 -15554 -9184 -15536
rect -9150 -15014 -9138 -14978
rect -8178 -14978 -8118 -14736
rect -7158 -14736 -7148 -14718
rect -7114 -14180 -7098 -14160
rect -6140 -14160 -6080 -13918
rect -5120 -13918 -5112 -13886
rect -5078 -13362 -5062 -13342
rect -4110 -13342 -4050 -13100
rect -3088 -13100 -3076 -13080
rect -3042 -13080 -3036 -12524
rect -2072 -12524 -2012 -12384
rect -1562 -12434 -1502 -12384
rect -42 -12414 -36 -12354
rect 24 -12414 30 -12354
rect -1776 -12440 -1288 -12434
rect -1776 -12474 -1764 -12440
rect -1300 -12474 -1288 -12440
rect -1776 -12480 -1288 -12474
rect -758 -12440 -270 -12434
rect -758 -12474 -746 -12440
rect -282 -12474 -270 -12440
rect -758 -12480 -270 -12474
rect -2072 -12560 -2058 -12524
rect -2064 -13080 -2058 -12560
rect -3042 -13100 -3028 -13080
rect -3812 -13150 -3324 -13144
rect -3812 -13184 -3800 -13150
rect -3336 -13184 -3324 -13150
rect -3812 -13190 -3324 -13184
rect -3604 -13252 -3544 -13190
rect -3812 -13258 -3324 -13252
rect -3812 -13292 -3800 -13258
rect -3336 -13292 -3324 -13258
rect -3812 -13298 -3324 -13292
rect -5078 -13886 -5072 -13362
rect -4110 -13370 -4094 -13342
rect -5078 -13918 -5060 -13886
rect -4100 -13894 -4094 -13370
rect -5848 -13968 -5360 -13962
rect -5848 -14002 -5836 -13968
rect -5372 -14002 -5360 -13968
rect -5848 -14008 -5360 -14002
rect -5650 -14070 -5590 -14008
rect -5848 -14076 -5360 -14070
rect -5848 -14110 -5836 -14076
rect -5372 -14110 -5360 -14076
rect -5848 -14116 -5360 -14110
rect -7114 -14718 -7108 -14180
rect -6140 -14184 -6130 -14160
rect -7114 -14736 -7098 -14718
rect -6136 -14722 -6130 -14184
rect -7884 -14786 -7396 -14780
rect -7884 -14820 -7872 -14786
rect -7408 -14820 -7396 -14786
rect -7884 -14826 -7396 -14820
rect -7670 -14888 -7610 -14826
rect -7884 -14894 -7396 -14888
rect -7884 -14928 -7872 -14894
rect -7408 -14928 -7396 -14894
rect -7884 -14934 -7396 -14928
rect -8178 -15010 -8166 -14978
rect -9150 -15536 -9144 -15014
rect -8172 -15532 -8166 -15010
rect -9150 -15554 -9138 -15536
rect -9198 -15796 -9138 -15554
rect -8178 -15554 -8166 -15532
rect -8132 -15010 -8118 -14978
rect -7158 -14978 -7098 -14736
rect -6140 -14736 -6130 -14722
rect -6096 -14184 -6080 -14160
rect -5120 -14160 -5060 -13918
rect -4108 -13918 -4094 -13894
rect -4060 -13370 -4050 -13342
rect -3088 -13342 -3028 -13100
rect -2068 -13100 -2058 -13080
rect -2024 -12560 -2012 -12524
rect -1046 -12524 -1000 -12512
rect -2024 -13080 -2018 -12560
rect -1046 -13076 -1040 -12524
rect -2024 -13100 -2008 -13080
rect -2794 -13150 -2306 -13144
rect -2794 -13184 -2782 -13150
rect -2318 -13184 -2306 -13150
rect -2794 -13190 -2306 -13184
rect -2582 -13252 -2522 -13190
rect -2794 -13258 -2306 -13252
rect -2794 -13292 -2782 -13258
rect -2318 -13292 -2306 -13258
rect -2794 -13298 -2306 -13292
rect -3088 -13370 -3076 -13342
rect -4060 -13894 -4054 -13370
rect -3082 -13894 -3076 -13370
rect -4060 -13918 -4048 -13894
rect -4830 -13968 -4342 -13962
rect -4830 -14002 -4818 -13968
rect -4354 -14002 -4342 -13968
rect -4830 -14008 -4342 -14002
rect -4620 -14070 -4560 -14008
rect -4830 -14076 -4342 -14070
rect -4830 -14110 -4818 -14076
rect -4354 -14110 -4342 -14076
rect -4830 -14116 -4342 -14110
rect -5120 -14176 -5112 -14160
rect -6096 -14722 -6090 -14184
rect -5118 -14714 -5112 -14176
rect -6096 -14736 -6080 -14722
rect -6866 -14786 -6378 -14780
rect -6866 -14820 -6854 -14786
rect -6390 -14820 -6378 -14786
rect -6866 -14826 -6378 -14820
rect -6658 -14888 -6598 -14826
rect -6866 -14894 -6378 -14888
rect -6866 -14928 -6854 -14894
rect -6390 -14928 -6378 -14894
rect -6866 -14934 -6378 -14928
rect -7158 -15008 -7148 -14978
rect -8132 -15532 -8126 -15010
rect -7154 -15530 -7148 -15008
rect -8132 -15554 -8118 -15532
rect -8902 -15604 -8414 -15598
rect -8902 -15638 -8890 -15604
rect -8426 -15638 -8414 -15604
rect -8902 -15644 -8414 -15638
rect -8694 -15706 -8634 -15644
rect -8902 -15712 -8414 -15706
rect -8902 -15746 -8890 -15712
rect -8426 -15746 -8414 -15712
rect -8902 -15752 -8414 -15746
rect -9198 -15826 -9184 -15796
rect -9190 -16356 -9184 -15826
rect -9198 -16372 -9184 -16356
rect -9150 -15826 -9138 -15796
rect -8178 -15796 -8118 -15554
rect -7158 -15554 -7148 -15530
rect -7114 -15008 -7098 -14978
rect -6140 -14978 -6080 -14736
rect -5120 -14736 -5112 -14714
rect -5078 -14176 -5060 -14160
rect -4108 -14160 -4048 -13918
rect -3086 -13918 -3076 -13894
rect -3042 -13370 -3028 -13342
rect -2068 -13342 -2008 -13100
rect -1052 -13100 -1040 -13076
rect -1006 -13076 -1000 -12524
rect -36 -12524 24 -12414
rect -36 -12560 -22 -12524
rect -1006 -13100 -992 -13076
rect -28 -13080 -22 -12560
rect -1776 -13150 -1288 -13144
rect -1776 -13184 -1764 -13150
rect -1300 -13184 -1288 -13150
rect -1776 -13190 -1288 -13184
rect -1570 -13252 -1510 -13190
rect -1776 -13258 -1288 -13252
rect -1776 -13292 -1764 -13258
rect -1300 -13292 -1288 -13258
rect -1776 -13298 -1288 -13292
rect -2068 -13370 -2058 -13342
rect -3042 -13894 -3036 -13370
rect -2064 -13894 -2058 -13370
rect -3042 -13918 -3026 -13894
rect -3812 -13968 -3324 -13962
rect -3812 -14002 -3800 -13968
rect -3336 -14002 -3324 -13968
rect -3812 -14008 -3324 -14002
rect -3604 -14070 -3544 -14008
rect -3812 -14076 -3324 -14070
rect -3812 -14110 -3800 -14076
rect -3336 -14110 -3324 -14076
rect -3812 -14116 -3324 -14110
rect -5078 -14714 -5072 -14176
rect -4108 -14184 -4094 -14160
rect -5078 -14736 -5060 -14714
rect -4100 -14722 -4094 -14184
rect -5848 -14786 -5360 -14780
rect -5848 -14820 -5836 -14786
rect -5372 -14820 -5360 -14786
rect -5848 -14826 -5360 -14820
rect -5656 -14888 -5596 -14826
rect -5848 -14894 -5360 -14888
rect -5848 -14928 -5836 -14894
rect -5372 -14928 -5360 -14894
rect -5848 -14934 -5360 -14928
rect -7114 -15530 -7108 -15008
rect -6140 -15012 -6130 -14978
rect -7114 -15554 -7098 -15530
rect -6136 -15534 -6130 -15012
rect -7884 -15604 -7396 -15598
rect -7884 -15638 -7872 -15604
rect -7408 -15638 -7396 -15604
rect -7884 -15644 -7396 -15638
rect -7676 -15706 -7616 -15644
rect -7884 -15712 -7396 -15706
rect -7884 -15746 -7872 -15712
rect -7408 -15746 -7396 -15712
rect -7884 -15752 -7396 -15746
rect -8178 -15822 -8166 -15796
rect -9150 -16356 -9144 -15826
rect -8172 -16352 -8166 -15822
rect -9150 -16372 -9138 -16356
rect -9198 -16614 -9138 -16372
rect -8178 -16372 -8166 -16352
rect -8132 -15822 -8118 -15796
rect -7158 -15796 -7098 -15554
rect -6140 -15554 -6130 -15534
rect -6096 -15012 -6080 -14978
rect -5120 -14978 -5060 -14736
rect -4108 -14736 -4094 -14722
rect -4060 -14184 -4048 -14160
rect -3086 -14160 -3026 -13918
rect -2066 -13918 -2058 -13894
rect -2024 -13370 -2008 -13342
rect -1052 -13342 -992 -13100
rect -30 -13100 -22 -13080
rect 12 -12560 24 -12524
rect 12 -13080 18 -12560
rect 12 -13100 30 -13080
rect -758 -13150 -270 -13144
rect -758 -13184 -746 -13150
rect -282 -13184 -270 -13150
rect -758 -13190 -270 -13184
rect -550 -13252 -490 -13190
rect -758 -13258 -270 -13252
rect -758 -13292 -746 -13258
rect -282 -13292 -270 -13258
rect -758 -13298 -270 -13292
rect -1052 -13366 -1040 -13342
rect -2024 -13894 -2018 -13370
rect -1046 -13890 -1040 -13366
rect -2024 -13918 -2006 -13894
rect -2794 -13968 -2306 -13962
rect -2794 -14002 -2782 -13968
rect -2318 -14002 -2306 -13968
rect -2794 -14008 -2306 -14002
rect -2582 -14070 -2522 -14008
rect -2794 -14076 -2306 -14070
rect -2794 -14110 -2782 -14076
rect -2318 -14110 -2306 -14076
rect -2794 -14116 -2306 -14110
rect -3086 -14184 -3076 -14160
rect -4060 -14722 -4054 -14184
rect -3082 -14722 -3076 -14184
rect -4060 -14736 -4048 -14722
rect -4830 -14786 -4342 -14780
rect -4830 -14820 -4818 -14786
rect -4354 -14820 -4342 -14786
rect -4830 -14826 -4342 -14820
rect -4626 -14888 -4566 -14826
rect -4830 -14894 -4342 -14888
rect -4830 -14928 -4818 -14894
rect -4354 -14928 -4342 -14894
rect -4830 -14934 -4342 -14928
rect -5120 -15004 -5112 -14978
rect -6096 -15534 -6090 -15012
rect -5118 -15526 -5112 -15004
rect -6096 -15554 -6080 -15534
rect -6866 -15604 -6378 -15598
rect -6866 -15638 -6854 -15604
rect -6390 -15638 -6378 -15604
rect -6866 -15644 -6378 -15638
rect -6660 -15706 -6600 -15644
rect -6866 -15712 -6378 -15706
rect -6866 -15746 -6854 -15712
rect -6390 -15746 -6378 -15712
rect -6866 -15752 -6378 -15746
rect -7158 -15820 -7148 -15796
rect -8132 -16352 -8126 -15822
rect -7154 -16350 -7148 -15820
rect -8132 -16372 -8118 -16352
rect -8902 -16422 -8414 -16416
rect -8902 -16456 -8890 -16422
rect -8426 -16456 -8414 -16422
rect -8902 -16462 -8414 -16456
rect -8692 -16524 -8632 -16462
rect -8902 -16530 -8414 -16524
rect -8902 -16564 -8890 -16530
rect -8426 -16564 -8414 -16530
rect -8902 -16570 -8414 -16564
rect -9198 -16646 -9184 -16614
rect -9190 -17168 -9184 -16646
rect -9198 -17190 -9184 -17168
rect -9150 -16646 -9138 -16614
rect -8178 -16614 -8118 -16372
rect -7158 -16372 -7148 -16350
rect -7114 -15820 -7098 -15796
rect -6140 -15796 -6080 -15554
rect -5120 -15554 -5112 -15526
rect -5078 -15004 -5060 -14978
rect -4108 -14978 -4048 -14736
rect -3086 -14736 -3076 -14722
rect -3042 -14184 -3026 -14160
rect -2066 -14160 -2006 -13918
rect -1050 -13918 -1040 -13890
rect -1006 -13366 -992 -13342
rect -30 -13342 30 -13100
rect -1006 -13890 -1000 -13366
rect -30 -13370 -22 -13342
rect -1006 -13918 -990 -13890
rect -1776 -13968 -1288 -13962
rect -1776 -14002 -1764 -13968
rect -1300 -14002 -1288 -13968
rect -1776 -14008 -1288 -14002
rect -1570 -14070 -1510 -14008
rect -1776 -14076 -1288 -14070
rect -1776 -14110 -1764 -14076
rect -1300 -14110 -1288 -14076
rect -1776 -14116 -1288 -14110
rect -2066 -14184 -2058 -14160
rect -3042 -14722 -3036 -14184
rect -2064 -14722 -2058 -14184
rect -3042 -14736 -3026 -14722
rect -3812 -14786 -3324 -14780
rect -3812 -14820 -3800 -14786
rect -3336 -14820 -3324 -14786
rect -3812 -14826 -3324 -14820
rect -3610 -14888 -3550 -14826
rect -3812 -14894 -3324 -14888
rect -3812 -14928 -3800 -14894
rect -3336 -14928 -3324 -14894
rect -3812 -14934 -3324 -14928
rect -5078 -15526 -5072 -15004
rect -4108 -15012 -4094 -14978
rect -5078 -15554 -5060 -15526
rect -4100 -15534 -4094 -15012
rect -5848 -15604 -5360 -15598
rect -5848 -15638 -5836 -15604
rect -5372 -15638 -5360 -15604
rect -5848 -15644 -5360 -15638
rect -5658 -15706 -5598 -15644
rect -5848 -15712 -5360 -15706
rect -5848 -15746 -5836 -15712
rect -5372 -15746 -5360 -15712
rect -5848 -15752 -5360 -15746
rect -7114 -16350 -7108 -15820
rect -6140 -15824 -6130 -15796
rect -7114 -16372 -7098 -16350
rect -6136 -16354 -6130 -15824
rect -7884 -16422 -7396 -16416
rect -7884 -16456 -7872 -16422
rect -7408 -16456 -7396 -16422
rect -7884 -16462 -7396 -16456
rect -7678 -16524 -7618 -16462
rect -7884 -16530 -7396 -16524
rect -7884 -16564 -7872 -16530
rect -7408 -16564 -7396 -16530
rect -7884 -16570 -7396 -16564
rect -8178 -16642 -8166 -16614
rect -9150 -17168 -9144 -16646
rect -8172 -17164 -8166 -16642
rect -9150 -17190 -9138 -17168
rect -9198 -17432 -9138 -17190
rect -8178 -17190 -8166 -17164
rect -8132 -16642 -8118 -16614
rect -7158 -16614 -7098 -16372
rect -6140 -16372 -6130 -16354
rect -6096 -15824 -6080 -15796
rect -5120 -15796 -5060 -15554
rect -4108 -15554 -4094 -15534
rect -4060 -15012 -4048 -14978
rect -3086 -14978 -3026 -14736
rect -2066 -14736 -2058 -14722
rect -2024 -14184 -2006 -14160
rect -1050 -14160 -990 -13918
rect -28 -13918 -22 -13370
rect 12 -13370 30 -13342
rect 12 -13894 18 -13370
rect 12 -13918 32 -13894
rect -758 -13968 -270 -13962
rect -758 -14002 -746 -13968
rect -282 -14002 -270 -13968
rect -758 -14008 -270 -14002
rect -550 -14070 -490 -14008
rect -758 -14076 -270 -14070
rect -758 -14110 -746 -14076
rect -282 -14110 -270 -14076
rect -758 -14116 -270 -14110
rect -1050 -14180 -1040 -14160
rect -2024 -14722 -2018 -14184
rect -1046 -14718 -1040 -14180
rect -2024 -14736 -2006 -14722
rect -2794 -14786 -2306 -14780
rect -2794 -14820 -2782 -14786
rect -2318 -14820 -2306 -14786
rect -2794 -14826 -2306 -14820
rect -2588 -14888 -2528 -14826
rect -2794 -14894 -2306 -14888
rect -2794 -14928 -2782 -14894
rect -2318 -14928 -2306 -14894
rect -2794 -14934 -2306 -14928
rect -3086 -15012 -3076 -14978
rect -4060 -15534 -4054 -15012
rect -3082 -15534 -3076 -15012
rect -4060 -15554 -4048 -15534
rect -4830 -15604 -4342 -15598
rect -4830 -15638 -4818 -15604
rect -4354 -15638 -4342 -15604
rect -4830 -15644 -4342 -15638
rect -4628 -15706 -4568 -15644
rect -4830 -15712 -4342 -15706
rect -4830 -15746 -4818 -15712
rect -4354 -15746 -4342 -15712
rect -4830 -15752 -4342 -15746
rect -5120 -15816 -5112 -15796
rect -6096 -16354 -6090 -15824
rect -5118 -16346 -5112 -15816
rect -6096 -16372 -6080 -16354
rect -6866 -16422 -6378 -16416
rect -6866 -16456 -6854 -16422
rect -6390 -16456 -6378 -16422
rect -6866 -16462 -6378 -16456
rect -6658 -16524 -6598 -16462
rect -6866 -16530 -6378 -16524
rect -6866 -16564 -6854 -16530
rect -6390 -16564 -6378 -16530
rect -6866 -16570 -6378 -16564
rect -7158 -16640 -7148 -16614
rect -8132 -17164 -8126 -16642
rect -7154 -17162 -7148 -16640
rect -8132 -17190 -8118 -17164
rect -8902 -17240 -8414 -17234
rect -8902 -17274 -8890 -17240
rect -8426 -17274 -8414 -17240
rect -8902 -17280 -8414 -17274
rect -8690 -17342 -8630 -17280
rect -8902 -17348 -8414 -17342
rect -8902 -17382 -8890 -17348
rect -8426 -17382 -8414 -17348
rect -8902 -17388 -8414 -17382
rect -9198 -17458 -9184 -17432
rect -9190 -17986 -9184 -17458
rect -9198 -18008 -9184 -17986
rect -9150 -17458 -9138 -17432
rect -8178 -17432 -8118 -17190
rect -7158 -17190 -7148 -17162
rect -7114 -16640 -7098 -16614
rect -6140 -16614 -6080 -16372
rect -5120 -16372 -5112 -16346
rect -5078 -15816 -5060 -15796
rect -4108 -15796 -4048 -15554
rect -3086 -15554 -3076 -15534
rect -3042 -15012 -3026 -14978
rect -2066 -14978 -2006 -14736
rect -1050 -14736 -1040 -14718
rect -1006 -14180 -990 -14160
rect -28 -14160 32 -13918
rect -1006 -14718 -1000 -14180
rect -1006 -14736 -990 -14718
rect -1776 -14786 -1288 -14780
rect -1776 -14820 -1764 -14786
rect -1300 -14820 -1288 -14786
rect -1776 -14826 -1288 -14820
rect -1576 -14888 -1516 -14826
rect -1776 -14894 -1288 -14888
rect -1776 -14928 -1764 -14894
rect -1300 -14928 -1288 -14894
rect -1776 -14934 -1288 -14928
rect -2066 -15012 -2058 -14978
rect -3042 -15534 -3036 -15012
rect -2064 -15534 -2058 -15012
rect -3042 -15554 -3026 -15534
rect -3812 -15604 -3324 -15598
rect -3812 -15638 -3800 -15604
rect -3336 -15638 -3324 -15604
rect -3812 -15644 -3324 -15638
rect -3612 -15706 -3552 -15644
rect -3812 -15712 -3324 -15706
rect -3812 -15746 -3800 -15712
rect -3336 -15746 -3324 -15712
rect -3812 -15752 -3324 -15746
rect -5078 -16346 -5072 -15816
rect -4108 -15824 -4094 -15796
rect -5078 -16372 -5060 -16346
rect -4100 -16354 -4094 -15824
rect -5848 -16422 -5360 -16416
rect -5848 -16456 -5836 -16422
rect -5372 -16456 -5360 -16422
rect -5848 -16462 -5360 -16456
rect -5656 -16524 -5596 -16462
rect -5848 -16530 -5360 -16524
rect -5848 -16564 -5836 -16530
rect -5372 -16564 -5360 -16530
rect -5848 -16570 -5360 -16564
rect -7114 -17162 -7108 -16640
rect -6140 -16644 -6130 -16614
rect -7114 -17190 -7098 -17162
rect -6136 -17166 -6130 -16644
rect -7884 -17240 -7396 -17234
rect -7884 -17274 -7872 -17240
rect -7408 -17274 -7396 -17240
rect -7884 -17280 -7396 -17274
rect -7676 -17342 -7616 -17280
rect -7884 -17348 -7396 -17342
rect -7884 -17382 -7872 -17348
rect -7408 -17382 -7396 -17348
rect -7884 -17388 -7396 -17382
rect -8178 -17454 -8166 -17432
rect -9150 -17986 -9144 -17458
rect -8172 -17982 -8166 -17454
rect -9150 -18008 -9138 -17986
rect -9198 -18250 -9138 -18008
rect -8178 -18008 -8166 -17982
rect -8132 -17454 -8118 -17432
rect -7158 -17432 -7098 -17190
rect -6140 -17190 -6130 -17166
rect -6096 -16644 -6080 -16614
rect -5120 -16614 -5060 -16372
rect -4108 -16372 -4094 -16354
rect -4060 -15824 -4048 -15796
rect -3086 -15796 -3026 -15554
rect -2066 -15554 -2058 -15534
rect -2024 -15012 -2006 -14978
rect -1050 -14978 -990 -14736
rect -28 -14736 -22 -14160
rect 12 -14184 32 -14160
rect 12 -14722 18 -14184
rect 12 -14736 32 -14722
rect -758 -14786 -270 -14780
rect -758 -14820 -746 -14786
rect -282 -14820 -270 -14786
rect -758 -14826 -270 -14820
rect -556 -14888 -496 -14826
rect -758 -14894 -270 -14888
rect -758 -14928 -746 -14894
rect -282 -14928 -270 -14894
rect -758 -14934 -270 -14928
rect -1050 -15008 -1040 -14978
rect -2024 -15534 -2018 -15012
rect -1046 -15530 -1040 -15008
rect -2024 -15554 -2006 -15534
rect -2794 -15604 -2306 -15598
rect -2794 -15638 -2782 -15604
rect -2318 -15638 -2306 -15604
rect -2794 -15644 -2306 -15638
rect -2590 -15706 -2530 -15644
rect -2794 -15712 -2306 -15706
rect -2794 -15746 -2782 -15712
rect -2318 -15746 -2306 -15712
rect -2794 -15752 -2306 -15746
rect -3086 -15824 -3076 -15796
rect -4060 -16354 -4054 -15824
rect -3082 -16354 -3076 -15824
rect -4060 -16372 -4048 -16354
rect -4830 -16422 -4342 -16416
rect -4830 -16456 -4818 -16422
rect -4354 -16456 -4342 -16422
rect -4830 -16462 -4342 -16456
rect -4626 -16524 -4566 -16462
rect -4830 -16530 -4342 -16524
rect -4830 -16564 -4818 -16530
rect -4354 -16564 -4342 -16530
rect -4830 -16570 -4342 -16564
rect -5120 -16636 -5112 -16614
rect -6096 -17166 -6090 -16644
rect -5118 -17158 -5112 -16636
rect -6096 -17190 -6080 -17166
rect -6866 -17240 -6378 -17234
rect -6866 -17274 -6854 -17240
rect -6390 -17274 -6378 -17240
rect -6866 -17280 -6378 -17274
rect -6656 -17342 -6596 -17280
rect -6866 -17348 -6378 -17342
rect -6866 -17382 -6854 -17348
rect -6390 -17382 -6378 -17348
rect -6866 -17388 -6378 -17382
rect -7158 -17452 -7148 -17432
rect -8132 -17982 -8126 -17454
rect -7154 -17980 -7148 -17452
rect -8132 -18008 -8118 -17982
rect -8902 -18058 -8414 -18052
rect -8902 -18092 -8890 -18058
rect -8426 -18092 -8414 -18058
rect -8902 -18098 -8414 -18092
rect -8688 -18160 -8628 -18098
rect -8902 -18166 -8414 -18160
rect -8902 -18200 -8890 -18166
rect -8426 -18200 -8414 -18166
rect -8902 -18206 -8414 -18200
rect -9198 -18276 -9184 -18250
rect -9190 -18826 -9184 -18276
rect -9150 -18276 -9138 -18250
rect -8178 -18250 -8118 -18008
rect -7158 -18008 -7148 -17980
rect -7114 -17452 -7098 -17432
rect -6140 -17432 -6080 -17190
rect -5120 -17190 -5112 -17158
rect -5078 -16636 -5060 -16614
rect -4108 -16614 -4048 -16372
rect -3086 -16372 -3076 -16354
rect -3042 -15824 -3026 -15796
rect -2066 -15796 -2006 -15554
rect -1050 -15554 -1040 -15530
rect -1006 -15008 -990 -14978
rect -28 -14978 32 -14736
rect -1006 -15530 -1000 -15008
rect -1006 -15554 -990 -15530
rect -1776 -15604 -1288 -15598
rect -1776 -15638 -1764 -15604
rect -1300 -15638 -1288 -15604
rect -1776 -15644 -1288 -15638
rect -1578 -15706 -1518 -15644
rect -1776 -15712 -1288 -15706
rect -1776 -15746 -1764 -15712
rect -1300 -15746 -1288 -15712
rect -1776 -15752 -1288 -15746
rect -2066 -15824 -2058 -15796
rect -3042 -16354 -3036 -15824
rect -2064 -16354 -2058 -15824
rect -3042 -16372 -3026 -16354
rect -3812 -16422 -3324 -16416
rect -3812 -16456 -3800 -16422
rect -3336 -16456 -3324 -16422
rect -3812 -16462 -3324 -16456
rect -3610 -16524 -3550 -16462
rect -3812 -16530 -3324 -16524
rect -3812 -16564 -3800 -16530
rect -3336 -16564 -3324 -16530
rect -3812 -16570 -3324 -16564
rect -5078 -17158 -5072 -16636
rect -4108 -16644 -4094 -16614
rect -5078 -17190 -5060 -17158
rect -4100 -17166 -4094 -16644
rect -5848 -17240 -5360 -17234
rect -5848 -17274 -5836 -17240
rect -5372 -17274 -5360 -17240
rect -5848 -17280 -5360 -17274
rect -5654 -17342 -5594 -17280
rect -5848 -17348 -5360 -17342
rect -5848 -17382 -5836 -17348
rect -5372 -17382 -5360 -17348
rect -5848 -17388 -5360 -17382
rect -7114 -17980 -7108 -17452
rect -6140 -17456 -6130 -17432
rect -7114 -18008 -7098 -17980
rect -6136 -17984 -6130 -17456
rect -7884 -18058 -7396 -18052
rect -7884 -18092 -7872 -18058
rect -7408 -18092 -7396 -18058
rect -7884 -18098 -7396 -18092
rect -7674 -18160 -7614 -18098
rect -7884 -18166 -7396 -18160
rect -7884 -18200 -7872 -18166
rect -7408 -18200 -7396 -18166
rect -7884 -18206 -7396 -18200
rect -8178 -18272 -8166 -18250
rect -9150 -18826 -9144 -18276
rect -9190 -18838 -9144 -18826
rect -8172 -18826 -8166 -18272
rect -8132 -18272 -8118 -18250
rect -7158 -18250 -7098 -18008
rect -6140 -18008 -6130 -17984
rect -6096 -17456 -6080 -17432
rect -5120 -17432 -5060 -17190
rect -4108 -17190 -4094 -17166
rect -4060 -16644 -4048 -16614
rect -3086 -16614 -3026 -16372
rect -2066 -16372 -2058 -16354
rect -2024 -15824 -2006 -15796
rect -1050 -15796 -990 -15554
rect -28 -15554 -22 -14978
rect 12 -15012 32 -14978
rect 12 -15534 18 -15012
rect 12 -15554 32 -15534
rect -758 -15604 -270 -15598
rect -758 -15638 -746 -15604
rect -282 -15638 -270 -15604
rect -758 -15644 -270 -15638
rect -558 -15706 -498 -15644
rect -758 -15712 -270 -15706
rect -758 -15746 -746 -15712
rect -282 -15746 -270 -15712
rect -758 -15752 -270 -15746
rect -1050 -15820 -1040 -15796
rect -2024 -16354 -2018 -15824
rect -1046 -16350 -1040 -15820
rect -2024 -16372 -2006 -16354
rect -2794 -16422 -2306 -16416
rect -2794 -16456 -2782 -16422
rect -2318 -16456 -2306 -16422
rect -2794 -16462 -2306 -16456
rect -2588 -16524 -2528 -16462
rect -2794 -16530 -2306 -16524
rect -2794 -16564 -2782 -16530
rect -2318 -16564 -2306 -16530
rect -2794 -16570 -2306 -16564
rect -3086 -16644 -3076 -16614
rect -4060 -17166 -4054 -16644
rect -3082 -17166 -3076 -16644
rect -4060 -17190 -4048 -17166
rect -4830 -17240 -4342 -17234
rect -4830 -17274 -4818 -17240
rect -4354 -17274 -4342 -17240
rect -4830 -17280 -4342 -17274
rect -4624 -17342 -4564 -17280
rect -4830 -17348 -4342 -17342
rect -4830 -17382 -4818 -17348
rect -4354 -17382 -4342 -17348
rect -4830 -17388 -4342 -17382
rect -5120 -17448 -5112 -17432
rect -6096 -17984 -6090 -17456
rect -5118 -17976 -5112 -17448
rect -6096 -18008 -6080 -17984
rect -6866 -18058 -6378 -18052
rect -6866 -18092 -6854 -18058
rect -6390 -18092 -6378 -18058
rect -6866 -18098 -6378 -18092
rect -6654 -18160 -6594 -18098
rect -6866 -18166 -6378 -18160
rect -6866 -18200 -6854 -18166
rect -6390 -18200 -6378 -18166
rect -6866 -18206 -6378 -18200
rect -7158 -18270 -7148 -18250
rect -8132 -18826 -8126 -18272
rect -7154 -18780 -7148 -18270
rect -8172 -18838 -8126 -18826
rect -7164 -18826 -7148 -18780
rect -7114 -18270 -7098 -18250
rect -6140 -18250 -6080 -18008
rect -5120 -18008 -5112 -17976
rect -5078 -17448 -5060 -17432
rect -4108 -17432 -4048 -17190
rect -3086 -17190 -3076 -17166
rect -3042 -16644 -3026 -16614
rect -2066 -16614 -2006 -16372
rect -1050 -16372 -1040 -16350
rect -1006 -15820 -990 -15796
rect -28 -15796 32 -15554
rect -1006 -16350 -1000 -15820
rect -1006 -16372 -990 -16350
rect -1776 -16422 -1288 -16416
rect -1776 -16456 -1764 -16422
rect -1300 -16456 -1288 -16422
rect -1776 -16462 -1288 -16456
rect -1576 -16524 -1516 -16462
rect -1776 -16530 -1288 -16524
rect -1776 -16564 -1764 -16530
rect -1300 -16564 -1288 -16530
rect -1776 -16570 -1288 -16564
rect -2066 -16644 -2058 -16614
rect -3042 -17166 -3036 -16644
rect -2064 -17166 -2058 -16644
rect -3042 -17190 -3026 -17166
rect -3812 -17240 -3324 -17234
rect -3812 -17274 -3800 -17240
rect -3336 -17274 -3324 -17240
rect -3812 -17280 -3324 -17274
rect -3608 -17342 -3548 -17280
rect -3812 -17348 -3324 -17342
rect -3812 -17382 -3800 -17348
rect -3336 -17382 -3324 -17348
rect -3812 -17388 -3324 -17382
rect -5078 -17976 -5072 -17448
rect -4108 -17456 -4094 -17432
rect -5078 -18008 -5060 -17976
rect -4100 -17984 -4094 -17456
rect -5848 -18058 -5360 -18052
rect -5848 -18092 -5836 -18058
rect -5372 -18092 -5360 -18058
rect -5848 -18098 -5360 -18092
rect -5652 -18160 -5592 -18098
rect -5848 -18166 -5360 -18160
rect -5848 -18200 -5836 -18166
rect -5372 -18200 -5360 -18166
rect -5848 -18206 -5360 -18200
rect -7114 -18780 -7108 -18270
rect -6140 -18274 -6130 -18250
rect -7114 -18826 -7104 -18780
rect -8902 -18876 -8414 -18870
rect -8902 -18910 -8890 -18876
rect -8426 -18910 -8414 -18876
rect -8902 -18916 -8414 -18910
rect -7884 -18876 -7396 -18870
rect -7884 -18910 -7872 -18876
rect -7408 -18910 -7396 -18876
rect -7884 -18916 -7396 -18910
rect -7164 -19000 -7104 -18826
rect -6136 -18826 -6130 -18274
rect -6096 -18274 -6080 -18250
rect -5120 -18250 -5060 -18008
rect -4108 -18008 -4094 -17984
rect -4060 -17456 -4048 -17432
rect -3086 -17432 -3026 -17190
rect -2066 -17190 -2058 -17166
rect -2024 -16644 -2006 -16614
rect -1050 -16614 -990 -16372
rect -28 -16372 -22 -15796
rect 12 -15824 32 -15796
rect 12 -16354 18 -15824
rect 12 -16372 32 -16354
rect -758 -16422 -270 -16416
rect -758 -16456 -746 -16422
rect -282 -16456 -270 -16422
rect -758 -16462 -270 -16456
rect -556 -16524 -496 -16462
rect -758 -16530 -270 -16524
rect -758 -16564 -746 -16530
rect -282 -16564 -270 -16530
rect -758 -16570 -270 -16564
rect -1050 -16640 -1040 -16614
rect -2024 -17166 -2018 -16644
rect -1046 -17162 -1040 -16640
rect -2024 -17190 -2006 -17166
rect -2794 -17240 -2306 -17234
rect -2794 -17274 -2782 -17240
rect -2318 -17274 -2306 -17240
rect -2794 -17280 -2306 -17274
rect -2586 -17342 -2526 -17280
rect -2794 -17348 -2306 -17342
rect -2794 -17382 -2782 -17348
rect -2318 -17382 -2306 -17348
rect -2794 -17388 -2306 -17382
rect -3086 -17456 -3076 -17432
rect -4060 -17984 -4054 -17456
rect -3082 -17984 -3076 -17456
rect -4060 -18008 -4048 -17984
rect -4830 -18058 -4342 -18052
rect -4830 -18092 -4818 -18058
rect -4354 -18092 -4342 -18058
rect -4830 -18098 -4342 -18092
rect -4622 -18160 -4562 -18098
rect -4830 -18166 -4342 -18160
rect -4830 -18200 -4818 -18166
rect -4354 -18200 -4342 -18166
rect -4830 -18206 -4342 -18200
rect -5120 -18266 -5112 -18250
rect -6096 -18826 -6090 -18274
rect -5118 -18778 -5112 -18266
rect -6136 -18838 -6090 -18826
rect -5126 -18826 -5112 -18778
rect -5078 -18266 -5060 -18250
rect -4108 -18250 -4048 -18008
rect -3086 -18008 -3076 -17984
rect -3042 -17456 -3026 -17432
rect -2066 -17432 -2006 -17190
rect -1050 -17190 -1040 -17162
rect -1006 -16640 -990 -16614
rect -28 -16614 32 -16372
rect -1006 -17162 -1000 -16640
rect -1006 -17190 -990 -17162
rect -1776 -17240 -1288 -17234
rect -1776 -17274 -1764 -17240
rect -1300 -17274 -1288 -17240
rect -1776 -17280 -1288 -17274
rect -1574 -17342 -1514 -17280
rect -1776 -17348 -1288 -17342
rect -1776 -17382 -1764 -17348
rect -1300 -17382 -1288 -17348
rect -1776 -17388 -1288 -17382
rect -2066 -17456 -2058 -17432
rect -3042 -17984 -3036 -17456
rect -2064 -17984 -2058 -17456
rect -3042 -18008 -3026 -17984
rect -3812 -18058 -3324 -18052
rect -3812 -18092 -3800 -18058
rect -3336 -18092 -3324 -18058
rect -3812 -18098 -3324 -18092
rect -3606 -18160 -3546 -18098
rect -3812 -18166 -3324 -18160
rect -3812 -18200 -3800 -18166
rect -3336 -18200 -3324 -18166
rect -3812 -18206 -3324 -18200
rect -5078 -18778 -5072 -18266
rect -4108 -18274 -4094 -18250
rect -5078 -18826 -5066 -18778
rect -6866 -18876 -6378 -18870
rect -6866 -18910 -6854 -18876
rect -6390 -18910 -6378 -18876
rect -6866 -18916 -6378 -18910
rect -5848 -18876 -5360 -18870
rect -5848 -18910 -5836 -18876
rect -5372 -18910 -5360 -18876
rect -5848 -18916 -5360 -18910
rect -5126 -19000 -5066 -18826
rect -4100 -18826 -4094 -18274
rect -4060 -18274 -4048 -18250
rect -3086 -18250 -3026 -18008
rect -2066 -18008 -2058 -17984
rect -2024 -17456 -2006 -17432
rect -1050 -17432 -990 -17190
rect -28 -17190 -22 -16614
rect 12 -16644 32 -16614
rect 12 -17166 18 -16644
rect 12 -17190 32 -17166
rect -758 -17240 -270 -17234
rect -758 -17274 -746 -17240
rect -282 -17274 -270 -17240
rect -758 -17280 -270 -17274
rect -554 -17342 -494 -17280
rect -758 -17348 -270 -17342
rect -758 -17382 -746 -17348
rect -282 -17382 -270 -17348
rect -758 -17388 -270 -17382
rect -1050 -17452 -1040 -17432
rect -2024 -17984 -2018 -17456
rect -1046 -17980 -1040 -17452
rect -2024 -18008 -2006 -17984
rect -2794 -18058 -2306 -18052
rect -2794 -18092 -2782 -18058
rect -2318 -18092 -2306 -18058
rect -2794 -18098 -2306 -18092
rect -2584 -18160 -2524 -18098
rect -2794 -18166 -2306 -18160
rect -2794 -18200 -2782 -18166
rect -2318 -18200 -2306 -18166
rect -2794 -18206 -2306 -18200
rect -3086 -18274 -3076 -18250
rect -4060 -18826 -4054 -18274
rect -3082 -18782 -3076 -18274
rect -4100 -18838 -4054 -18826
rect -3090 -18826 -3076 -18782
rect -3042 -18274 -3026 -18250
rect -2066 -18250 -2006 -18008
rect -1050 -18008 -1040 -17980
rect -1006 -17452 -990 -17432
rect -28 -17432 32 -17190
rect -1006 -17980 -1000 -17452
rect -1006 -18008 -990 -17980
rect -1776 -18058 -1288 -18052
rect -1776 -18092 -1764 -18058
rect -1300 -18092 -1288 -18058
rect -1776 -18098 -1288 -18092
rect -1572 -18160 -1512 -18098
rect -1776 -18166 -1288 -18160
rect -1776 -18200 -1764 -18166
rect -1300 -18200 -1288 -18166
rect -1776 -18206 -1288 -18200
rect -2066 -18274 -2058 -18250
rect -3042 -18782 -3036 -18274
rect -3042 -18826 -3030 -18782
rect -4830 -18876 -4342 -18870
rect -4830 -18910 -4818 -18876
rect -4354 -18910 -4342 -18876
rect -4830 -18916 -4342 -18910
rect -3812 -18876 -3324 -18870
rect -3812 -18910 -3800 -18876
rect -3336 -18910 -3324 -18876
rect -3812 -18916 -3324 -18910
rect -3090 -19000 -3030 -18826
rect -2064 -18826 -2058 -18274
rect -2024 -18274 -2006 -18250
rect -1050 -18250 -990 -18008
rect -28 -18008 -22 -17432
rect 12 -17456 32 -17432
rect 12 -17984 18 -17456
rect 12 -18008 32 -17984
rect -758 -18058 -270 -18052
rect -758 -18092 -746 -18058
rect -282 -18092 -270 -18058
rect -758 -18098 -270 -18092
rect -552 -18160 -492 -18098
rect -758 -18166 -270 -18160
rect -758 -18200 -746 -18166
rect -282 -18200 -270 -18166
rect -758 -18206 -270 -18200
rect -1050 -18270 -1040 -18250
rect -2024 -18826 -2018 -18274
rect -1046 -18784 -1040 -18270
rect -2064 -18838 -2018 -18826
rect -1054 -18826 -1040 -18784
rect -1006 -18270 -990 -18250
rect -28 -18250 32 -18008
rect -1006 -18784 -1000 -18270
rect -28 -18772 -22 -18250
rect -1006 -18826 -994 -18784
rect -2794 -18876 -2306 -18870
rect -2794 -18910 -2782 -18876
rect -2318 -18910 -2306 -18876
rect -2794 -18916 -2306 -18910
rect -1776 -18876 -1288 -18870
rect -1776 -18910 -1764 -18876
rect -1300 -18910 -1288 -18876
rect -1776 -18916 -1288 -18910
rect -1054 -19000 -994 -18826
rect -34 -18826 -22 -18772
rect 12 -18274 32 -18250
rect 12 -18772 18 -18274
rect 12 -18826 26 -18772
rect 1150 -18822 1210 -11682
rect -758 -18876 -270 -18870
rect -758 -18910 -746 -18876
rect -282 -18910 -270 -18876
rect -758 -18916 -270 -18910
rect -540 -19000 -480 -18916
rect -34 -19000 26 -18826
rect 1144 -18882 1150 -18822
rect 1210 -18882 1216 -18822
rect -7164 -19060 1130 -19000
rect -3404 -19808 -3398 -19748
rect -3338 -19808 -3332 -19748
rect -9508 -19894 -9448 -19888
rect -5434 -19954 -5428 -19894
rect -5368 -19954 -5362 -19894
rect -10668 -20082 -10662 -20022
rect -10602 -20082 -10596 -20022
rect -10662 -22254 -10602 -20082
rect -9508 -20086 -9448 -19954
rect -7990 -20082 -7984 -20022
rect -7924 -20082 -7918 -20022
rect -6958 -20082 -6952 -20022
rect -6892 -20082 -6886 -20022
rect -10524 -20146 -9448 -20086
rect -10524 -20274 -10464 -20146
rect -10016 -20184 -9956 -20146
rect -10226 -20190 -9738 -20184
rect -10226 -20224 -10214 -20190
rect -9750 -20224 -9738 -20190
rect -10226 -20230 -9738 -20224
rect -10524 -20320 -10508 -20274
rect -10514 -20850 -10508 -20320
rect -10474 -20320 -10464 -20274
rect -9508 -20274 -9448 -20146
rect -7984 -20184 -7924 -20082
rect -6952 -20184 -6892 -20082
rect -9208 -20190 -8720 -20184
rect -9208 -20224 -9196 -20190
rect -8732 -20224 -8720 -20190
rect -9208 -20230 -8720 -20224
rect -8190 -20190 -7702 -20184
rect -8190 -20224 -8178 -20190
rect -7714 -20224 -7702 -20190
rect -8190 -20230 -7702 -20224
rect -7172 -20190 -6684 -20184
rect -7172 -20224 -7160 -20190
rect -6696 -20224 -6684 -20190
rect -7172 -20230 -6684 -20224
rect -6154 -20190 -5666 -20184
rect -6154 -20224 -6142 -20190
rect -5678 -20224 -5666 -20190
rect -6154 -20230 -5666 -20224
rect -9508 -20314 -9490 -20274
rect -10474 -20850 -10468 -20320
rect -10514 -20862 -10468 -20850
rect -9496 -20850 -9490 -20314
rect -9456 -20314 -9448 -20274
rect -8478 -20274 -8432 -20262
rect -9456 -20850 -9450 -20314
rect -8478 -20786 -8472 -20274
rect -9496 -20862 -9450 -20850
rect -8486 -20850 -8472 -20786
rect -8438 -20786 -8432 -20274
rect -7460 -20274 -7414 -20262
rect -8438 -20850 -8426 -20786
rect -7460 -20804 -7454 -20274
rect -10226 -20900 -9738 -20894
rect -10226 -20934 -10214 -20900
rect -9750 -20934 -9738 -20900
rect -10226 -20940 -9738 -20934
rect -9208 -20900 -8720 -20894
rect -9208 -20934 -9196 -20900
rect -8732 -20934 -8720 -20900
rect -9208 -20940 -8720 -20934
rect -9004 -20984 -8944 -20940
rect -9010 -21044 -9004 -20984
rect -8944 -21044 -8938 -20984
rect -9510 -21148 -9504 -21088
rect -9444 -21148 -9438 -21088
rect -9504 -21190 -9444 -21148
rect -10524 -21250 -9444 -21190
rect -10524 -21386 -10464 -21250
rect -10020 -21296 -9960 -21250
rect -10226 -21302 -9738 -21296
rect -10226 -21336 -10214 -21302
rect -9750 -21336 -9738 -21302
rect -10226 -21342 -9738 -21336
rect -10524 -21432 -10508 -21386
rect -10514 -21962 -10508 -21432
rect -10474 -21432 -10464 -21386
rect -9504 -21386 -9444 -21250
rect -8486 -21192 -8426 -20850
rect -7468 -20850 -7454 -20804
rect -7420 -20804 -7414 -20274
rect -6442 -20274 -6396 -20262
rect -6442 -20788 -6436 -20274
rect -7420 -20850 -7408 -20804
rect -8190 -20900 -7702 -20894
rect -8190 -20934 -8178 -20900
rect -7714 -20934 -7702 -20900
rect -8190 -20940 -7702 -20934
rect -7986 -21044 -7980 -20984
rect -7920 -21044 -7914 -20984
rect -9208 -21302 -8720 -21296
rect -9208 -21336 -9196 -21302
rect -8732 -21336 -8720 -21302
rect -9208 -21342 -8720 -21336
rect -10474 -21962 -10468 -21432
rect -10514 -21974 -10468 -21962
rect -9504 -21962 -9490 -21386
rect -9456 -21962 -9444 -21386
rect -10226 -22012 -9738 -22006
rect -10226 -22046 -10214 -22012
rect -9750 -22046 -9738 -22012
rect -10226 -22052 -9738 -22046
rect -10668 -22314 -10662 -22254
rect -10602 -22314 -10596 -22254
rect -10662 -24380 -10602 -22314
rect -10226 -22414 -9738 -22408
rect -10226 -22448 -10214 -22414
rect -9750 -22448 -9738 -22414
rect -10226 -22454 -9738 -22448
rect -10514 -22498 -10468 -22486
rect -10514 -23040 -10508 -22498
rect -10520 -23074 -10508 -23040
rect -10474 -23040 -10468 -22498
rect -9504 -22498 -9444 -21962
rect -8486 -21386 -8426 -21252
rect -7980 -21296 -7920 -21044
rect -7468 -21088 -7408 -20850
rect -6450 -20850 -6436 -20788
rect -6402 -20788 -6396 -20274
rect -5428 -20274 -5368 -19954
rect -3898 -20082 -3892 -20022
rect -3832 -20082 -3826 -20022
rect -3892 -20184 -3832 -20082
rect -5136 -20190 -4648 -20184
rect -5136 -20224 -5124 -20190
rect -4660 -20224 -4648 -20190
rect -5136 -20230 -4648 -20224
rect -4118 -20190 -3630 -20184
rect -4118 -20224 -4106 -20190
rect -3642 -20224 -3630 -20190
rect -4118 -20230 -3630 -20224
rect -5428 -20338 -5418 -20274
rect -6402 -20850 -6390 -20788
rect -7172 -20900 -6684 -20894
rect -7172 -20934 -7160 -20900
rect -6696 -20934 -6684 -20900
rect -7172 -20940 -6684 -20934
rect -6954 -21044 -6948 -20984
rect -6888 -21044 -6882 -20984
rect -7474 -21148 -7468 -21088
rect -7408 -21148 -7402 -21088
rect -6948 -21296 -6888 -21044
rect -6450 -21192 -6390 -20850
rect -5424 -20850 -5418 -20338
rect -5384 -20338 -5368 -20274
rect -4406 -20274 -4360 -20262
rect -5384 -20850 -5378 -20338
rect -4406 -20778 -4400 -20274
rect -5424 -20862 -5378 -20850
rect -4418 -20850 -4400 -20778
rect -4366 -20778 -4360 -20274
rect -3398 -20274 -3338 -19808
rect -1374 -19954 -1368 -19894
rect -1308 -19954 -1302 -19894
rect 810 -19954 816 -19894
rect 876 -19954 882 -19894
rect -2902 -20082 -2896 -20022
rect -2836 -20082 -2830 -20022
rect -2896 -20184 -2836 -20082
rect -3100 -20190 -2612 -20184
rect -3100 -20224 -3088 -20190
rect -2624 -20224 -2612 -20190
rect -3100 -20230 -2612 -20224
rect -2082 -20190 -1594 -20184
rect -2082 -20224 -2070 -20190
rect -1606 -20224 -1594 -20190
rect -2082 -20230 -1594 -20224
rect -2896 -20232 -2836 -20230
rect -1368 -20262 -1308 -19954
rect -1064 -20190 -576 -20184
rect -1064 -20224 -1052 -20190
rect -588 -20224 -576 -20190
rect -1064 -20230 -576 -20224
rect -46 -20190 442 -20184
rect -46 -20224 -34 -20190
rect 430 -20224 442 -20190
rect -46 -20230 442 -20224
rect -4366 -20850 -4358 -20778
rect -6154 -20900 -5666 -20894
rect -6154 -20934 -6142 -20900
rect -5678 -20934 -5666 -20900
rect -6154 -20940 -5666 -20934
rect -5136 -20900 -4648 -20894
rect -5136 -20934 -5124 -20900
rect -4660 -20934 -4648 -20900
rect -5136 -20940 -4648 -20934
rect -5948 -20984 -5888 -20940
rect -4928 -20984 -4868 -20940
rect -5954 -21044 -5948 -20984
rect -5888 -21044 -5882 -20984
rect -4934 -21044 -4928 -20984
rect -4868 -21044 -4862 -20984
rect -5438 -21148 -5432 -21088
rect -5372 -21148 -5366 -21088
rect -8190 -21302 -7702 -21296
rect -8190 -21336 -8178 -21302
rect -7714 -21336 -7702 -21302
rect -8190 -21342 -7702 -21336
rect -7172 -21302 -6684 -21296
rect -7172 -21336 -7160 -21302
rect -6696 -21336 -6684 -21302
rect -7172 -21342 -6684 -21336
rect -8486 -21962 -8472 -21386
rect -8438 -21962 -8426 -21386
rect -7460 -21386 -7414 -21374
rect -7460 -21924 -7454 -21386
rect -9208 -22012 -8720 -22006
rect -9208 -22046 -9196 -22012
rect -8732 -22046 -8720 -22012
rect -9208 -22052 -8720 -22046
rect -9012 -22254 -8952 -22052
rect -9018 -22314 -9012 -22254
rect -8952 -22314 -8946 -22254
rect -9012 -22408 -8952 -22314
rect -9208 -22414 -8720 -22408
rect -9208 -22448 -9196 -22414
rect -8732 -22448 -8720 -22414
rect -9208 -22454 -8720 -22448
rect -9504 -22570 -9490 -22498
rect -10474 -23074 -10460 -23040
rect -9496 -23044 -9490 -22570
rect -10520 -23206 -10460 -23074
rect -9500 -23074 -9490 -23044
rect -9456 -22570 -9444 -22498
rect -8486 -22498 -8426 -21962
rect -7474 -21962 -7454 -21924
rect -7420 -21962 -7414 -21386
rect -8190 -22012 -7702 -22006
rect -8190 -22046 -8178 -22012
rect -7714 -22046 -7702 -22012
rect -8190 -22052 -7702 -22046
rect -7474 -22134 -7414 -21962
rect -6450 -21386 -6390 -21252
rect -6154 -21302 -5666 -21296
rect -6154 -21336 -6142 -21302
rect -5678 -21336 -5666 -21302
rect -6154 -21342 -5666 -21336
rect -6450 -21962 -6436 -21386
rect -6402 -21962 -6390 -21386
rect -7172 -22012 -6684 -22006
rect -7172 -22046 -7160 -22012
rect -6696 -22046 -6684 -22012
rect -7172 -22052 -6684 -22046
rect -7480 -22194 -7474 -22134
rect -7414 -22194 -7408 -22134
rect -8190 -22414 -7702 -22408
rect -8190 -22448 -8178 -22414
rect -7714 -22448 -7702 -22414
rect -8190 -22454 -7702 -22448
rect -9456 -23044 -9450 -22570
rect -9456 -23074 -9440 -23044
rect -10226 -23124 -9738 -23118
rect -10226 -23158 -10214 -23124
rect -9750 -23158 -9738 -23124
rect -10226 -23164 -9738 -23158
rect -10028 -23206 -9968 -23164
rect -9500 -23206 -9440 -23074
rect -8486 -23074 -8472 -22498
rect -8438 -23074 -8426 -22498
rect -7474 -22498 -7414 -22194
rect -7172 -22414 -6684 -22408
rect -7172 -22448 -7160 -22414
rect -6696 -22448 -6684 -22414
rect -7172 -22454 -6684 -22448
rect -7474 -22568 -7454 -22498
rect -9208 -23124 -8720 -23118
rect -9208 -23158 -9196 -23124
rect -8732 -23158 -8720 -23124
rect -9208 -23164 -8720 -23158
rect -10520 -23266 -9440 -23206
rect -9500 -23306 -9440 -23266
rect -8486 -23198 -8426 -23074
rect -7460 -23074 -7454 -22568
rect -7420 -23074 -7414 -22498
rect -7460 -23086 -7414 -23074
rect -6450 -22498 -6390 -21962
rect -5432 -21386 -5372 -21148
rect -4418 -21192 -4358 -20850
rect -3398 -20850 -3382 -20274
rect -3348 -20850 -3338 -20274
rect -2370 -20274 -2324 -20262
rect -2370 -20788 -2364 -20274
rect -4118 -20900 -3630 -20894
rect -4118 -20934 -4106 -20900
rect -3642 -20934 -3630 -20900
rect -4118 -20940 -3630 -20934
rect -3914 -21044 -3908 -20984
rect -3848 -21044 -3842 -20984
rect -4424 -21252 -4418 -21192
rect -4358 -21252 -4352 -21192
rect -5136 -21302 -4648 -21296
rect -5136 -21336 -5124 -21302
rect -4660 -21336 -4648 -21302
rect -5136 -21342 -4648 -21336
rect -5432 -21962 -5418 -21386
rect -5384 -21962 -5372 -21386
rect -6154 -22012 -5666 -22006
rect -6154 -22046 -6142 -22012
rect -5678 -22046 -5666 -22012
rect -6154 -22052 -5666 -22046
rect -5942 -22254 -5882 -22052
rect -5948 -22314 -5942 -22254
rect -5882 -22314 -5876 -22254
rect -5942 -22408 -5882 -22314
rect -6154 -22414 -5666 -22408
rect -6154 -22448 -6142 -22414
rect -5678 -22448 -5666 -22414
rect -6154 -22454 -5666 -22448
rect -6450 -23074 -6436 -22498
rect -6402 -23074 -6390 -22498
rect -5432 -22498 -5372 -21962
rect -4418 -21386 -4358 -21252
rect -3908 -21296 -3848 -21044
rect -3398 -21088 -3338 -20850
rect -2384 -20850 -2364 -20788
rect -2330 -20850 -2324 -20274
rect -1368 -20274 -1306 -20262
rect -1368 -20306 -1346 -20274
rect -3100 -20900 -2612 -20894
rect -3100 -20934 -3088 -20900
rect -2624 -20934 -2612 -20900
rect -3100 -20940 -2612 -20934
rect -2898 -20984 -2838 -20978
rect -3404 -21148 -3398 -21088
rect -3338 -21148 -3332 -21088
rect -2898 -21296 -2838 -21044
rect -2384 -21192 -2324 -20850
rect -1352 -20850 -1346 -20306
rect -1312 -20850 -1306 -20274
rect -334 -20274 -288 -20262
rect -334 -20816 -328 -20274
rect -1352 -20862 -1306 -20850
rect -340 -20850 -328 -20816
rect -294 -20816 -288 -20274
rect 684 -20274 730 -20262
rect 684 -20796 690 -20274
rect -294 -20850 -280 -20816
rect -2082 -20900 -1594 -20894
rect -2082 -20934 -2070 -20900
rect -1606 -20934 -1594 -20900
rect -2082 -20940 -1594 -20934
rect -1064 -20900 -576 -20894
rect -1064 -20934 -1052 -20900
rect -588 -20934 -576 -20900
rect -1064 -20940 -576 -20934
rect -1884 -20984 -1824 -20940
rect -866 -20984 -806 -20940
rect -1890 -21044 -1884 -20984
rect -1824 -21044 -1818 -20984
rect -866 -21050 -806 -21044
rect -340 -21078 -280 -20850
rect 676 -20850 690 -20796
rect 724 -20796 730 -20274
rect 724 -20850 736 -20796
rect -46 -20900 442 -20894
rect -46 -20934 -34 -20900
rect 430 -20934 442 -20900
rect -46 -20940 442 -20934
rect 164 -21078 224 -20940
rect 676 -21078 736 -20850
rect -1368 -21148 -1362 -21088
rect -1302 -21148 -1296 -21088
rect -340 -21138 736 -21078
rect -4118 -21302 -3630 -21296
rect -4118 -21336 -4106 -21302
rect -3642 -21336 -3630 -21302
rect -4118 -21342 -3630 -21336
rect -3100 -21302 -2612 -21296
rect -3100 -21336 -3088 -21302
rect -2624 -21336 -2612 -21302
rect -3100 -21342 -2612 -21336
rect -4418 -21962 -4400 -21386
rect -4366 -21962 -4358 -21386
rect -3388 -21386 -3342 -21374
rect -3388 -21906 -3382 -21386
rect -5136 -22012 -4648 -22006
rect -5136 -22046 -5124 -22012
rect -4660 -22046 -4648 -22012
rect -5136 -22052 -4648 -22046
rect -4934 -22254 -4874 -22052
rect -4940 -22314 -4934 -22254
rect -4874 -22314 -4868 -22254
rect -4934 -22408 -4874 -22314
rect -5136 -22414 -4648 -22408
rect -5136 -22448 -5124 -22414
rect -4660 -22448 -4648 -22414
rect -5136 -22454 -4648 -22448
rect -5432 -22604 -5418 -22498
rect -5424 -23012 -5418 -22604
rect -8190 -23124 -7702 -23118
rect -8190 -23158 -8178 -23124
rect -7714 -23158 -7702 -23124
rect -8190 -23164 -7702 -23158
rect -7172 -23124 -6684 -23118
rect -7172 -23158 -7160 -23124
rect -6696 -23158 -6684 -23124
rect -7172 -23164 -6684 -23158
rect -9506 -23366 -9500 -23306
rect -9440 -23366 -9434 -23306
rect -9012 -23478 -9006 -23418
rect -8946 -23478 -8940 -23418
rect -9006 -23520 -8946 -23478
rect -10226 -23526 -9738 -23520
rect -10226 -23560 -10214 -23526
rect -9750 -23560 -9738 -23526
rect -10226 -23566 -9738 -23560
rect -9208 -23526 -8720 -23520
rect -9208 -23560 -9196 -23526
rect -8732 -23560 -8720 -23526
rect -9208 -23566 -8720 -23560
rect -10514 -23610 -10468 -23598
rect -10514 -24144 -10508 -23610
rect -10524 -24186 -10508 -24144
rect -10474 -24144 -10468 -23610
rect -9496 -23610 -9450 -23598
rect -10474 -24186 -10464 -24144
rect -9496 -24150 -9490 -23610
rect -10524 -24330 -10464 -24186
rect -9506 -24186 -9490 -24150
rect -9456 -24150 -9450 -23610
rect -8486 -23610 -8426 -23258
rect -7982 -23418 -7922 -23164
rect -7470 -23366 -7464 -23306
rect -7404 -23366 -7398 -23306
rect -7988 -23478 -7982 -23418
rect -7922 -23478 -7916 -23418
rect -8190 -23526 -7702 -23520
rect -8190 -23560 -8178 -23526
rect -7714 -23560 -7702 -23526
rect -8190 -23566 -7702 -23560
rect -8486 -23712 -8472 -23610
rect -9456 -24186 -9446 -24150
rect -10226 -24236 -9738 -24230
rect -10226 -24270 -10214 -24236
rect -9750 -24270 -9738 -24236
rect -10226 -24276 -9738 -24270
rect -10020 -24330 -9960 -24276
rect -9506 -24330 -9446 -24186
rect -8478 -24186 -8472 -23712
rect -8438 -23712 -8426 -23610
rect -7464 -23610 -7404 -23366
rect -6950 -23418 -6890 -23164
rect -6450 -23198 -6390 -23074
rect -5428 -23074 -5418 -23012
rect -5384 -22604 -5372 -22498
rect -4418 -22498 -4358 -21962
rect -3398 -21962 -3382 -21906
rect -3348 -21906 -3342 -21386
rect -2384 -21386 -2324 -21252
rect -2082 -21302 -1594 -21296
rect -2082 -21336 -2070 -21302
rect -1606 -21336 -1594 -21302
rect -2082 -21342 -1594 -21336
rect -3348 -21962 -3338 -21906
rect -4118 -22012 -3630 -22006
rect -4118 -22046 -4106 -22012
rect -3642 -22046 -3630 -22012
rect -4118 -22052 -3630 -22046
rect -3398 -22134 -3338 -21962
rect -2384 -21962 -2364 -21386
rect -2330 -21962 -2324 -21386
rect -3100 -22012 -2612 -22006
rect -3100 -22046 -3088 -22012
rect -2624 -22046 -2612 -22012
rect -3100 -22052 -2612 -22046
rect -3404 -22194 -3398 -22134
rect -3338 -22194 -3332 -22134
rect -4118 -22414 -3630 -22408
rect -4118 -22448 -4106 -22414
rect -3642 -22448 -3630 -22414
rect -4118 -22454 -3630 -22448
rect -5384 -23012 -5378 -22604
rect -5384 -23074 -5368 -23012
rect -6154 -23124 -5666 -23118
rect -6154 -23158 -6142 -23124
rect -5678 -23158 -5666 -23124
rect -6154 -23164 -5666 -23158
rect -6956 -23478 -6950 -23418
rect -6890 -23478 -6884 -23418
rect -7172 -23526 -6684 -23520
rect -7172 -23560 -7160 -23526
rect -6696 -23560 -6684 -23526
rect -7172 -23566 -6684 -23560
rect -7464 -23650 -7454 -23610
rect -8438 -24186 -8432 -23712
rect -8478 -24198 -8432 -24186
rect -7460 -24186 -7454 -23650
rect -7420 -23650 -7404 -23610
rect -6450 -23610 -6390 -23258
rect -5428 -23306 -5368 -23074
rect -4418 -23074 -4400 -22498
rect -4366 -23074 -4358 -22498
rect -3398 -22498 -3338 -22194
rect -3100 -22414 -2612 -22408
rect -3100 -22448 -3088 -22414
rect -2624 -22448 -2612 -22414
rect -3100 -22454 -2612 -22448
rect -3398 -22540 -3382 -22498
rect -5136 -23124 -4648 -23118
rect -5136 -23158 -5124 -23124
rect -4660 -23158 -4648 -23124
rect -5136 -23164 -4648 -23158
rect -4418 -23198 -4358 -23074
rect -3388 -23074 -3382 -22540
rect -3348 -22540 -3338 -22498
rect -2384 -22498 -2324 -21962
rect -1362 -21386 -1302 -21148
rect -340 -21192 -280 -21138
rect -1064 -21302 -576 -21296
rect -1064 -21336 -1052 -21302
rect -588 -21336 -576 -21302
rect -1064 -21342 -576 -21336
rect -1362 -21962 -1346 -21386
rect -1312 -21962 -1302 -21386
rect -2082 -22012 -1594 -22006
rect -2082 -22046 -2070 -22012
rect -1606 -22046 -1594 -22012
rect -2082 -22052 -1594 -22046
rect -1872 -22254 -1812 -22052
rect -1878 -22314 -1872 -22254
rect -1812 -22314 -1806 -22254
rect -1872 -22408 -1812 -22314
rect -2082 -22414 -1594 -22408
rect -2082 -22448 -2070 -22414
rect -1606 -22448 -1594 -22414
rect -2082 -22454 -1594 -22448
rect -3348 -23074 -3342 -22540
rect -3388 -23086 -3342 -23074
rect -2384 -23074 -2364 -22498
rect -2330 -23074 -2324 -22498
rect -1362 -22498 -1302 -21962
rect -340 -21386 -280 -21252
rect 164 -21296 224 -21138
rect -46 -21302 442 -21296
rect -46 -21336 -34 -21302
rect 430 -21336 442 -21302
rect -46 -21342 442 -21336
rect -340 -21962 -328 -21386
rect -294 -21962 -280 -21386
rect -1064 -22012 -576 -22006
rect -1064 -22046 -1052 -22012
rect -588 -22046 -576 -22012
rect -1064 -22052 -576 -22046
rect -846 -22254 -786 -22052
rect -340 -22198 -280 -21962
rect 676 -21386 736 -21138
rect 676 -21962 690 -21386
rect 724 -21962 736 -21386
rect -46 -22012 442 -22006
rect -46 -22046 -34 -22012
rect 430 -22046 442 -22012
rect -46 -22052 442 -22046
rect 160 -22198 220 -22052
rect 676 -22198 736 -21962
rect 816 -22134 876 -19954
rect 930 -21044 936 -20984
rect 996 -21044 1002 -20984
rect 810 -22194 816 -22134
rect 876 -22194 882 -22134
rect -852 -22314 -846 -22254
rect -786 -22314 -780 -22254
rect -340 -22258 736 -22198
rect -846 -22408 -786 -22314
rect -1064 -22414 -576 -22408
rect -1064 -22448 -1052 -22414
rect -588 -22448 -576 -22414
rect -1064 -22454 -576 -22448
rect -1362 -22554 -1346 -22498
rect -1352 -23028 -1346 -22554
rect -4118 -23124 -3630 -23118
rect -4118 -23158 -4106 -23124
rect -3642 -23158 -3630 -23124
rect -4118 -23164 -3630 -23158
rect -3100 -23124 -2612 -23118
rect -3100 -23158 -3088 -23124
rect -2624 -23158 -2612 -23124
rect -3100 -23164 -2612 -23158
rect -5434 -23366 -5428 -23306
rect -5368 -23366 -5362 -23306
rect -5956 -23478 -5950 -23418
rect -5890 -23478 -5884 -23418
rect -4936 -23478 -4930 -23418
rect -4870 -23478 -4864 -23418
rect -5950 -23520 -5890 -23478
rect -4930 -23520 -4870 -23478
rect -6154 -23526 -5666 -23520
rect -6154 -23560 -6142 -23526
rect -5678 -23560 -5666 -23526
rect -6154 -23566 -5666 -23560
rect -5136 -23526 -4648 -23520
rect -5136 -23560 -5124 -23526
rect -4660 -23560 -4648 -23526
rect -5136 -23566 -4648 -23560
rect -6450 -23648 -6436 -23610
rect -7420 -24186 -7414 -23650
rect -7460 -24198 -7414 -24186
rect -6442 -24186 -6436 -23648
rect -6402 -23648 -6390 -23610
rect -5424 -23610 -5378 -23598
rect -6402 -24186 -6396 -23648
rect -5424 -24126 -5418 -23610
rect -6442 -24198 -6396 -24186
rect -5426 -24186 -5418 -24126
rect -5384 -24126 -5378 -23610
rect -4418 -23610 -4358 -23258
rect -3910 -23418 -3850 -23164
rect -3400 -23366 -3394 -23306
rect -3334 -23366 -3328 -23306
rect -3916 -23478 -3910 -23418
rect -3850 -23478 -3844 -23418
rect -4118 -23526 -3630 -23520
rect -4118 -23560 -4106 -23526
rect -3642 -23560 -3630 -23526
rect -4118 -23566 -3630 -23560
rect -4418 -23670 -4400 -23610
rect -5384 -24186 -5366 -24126
rect -9208 -24236 -8720 -24230
rect -9208 -24270 -9196 -24236
rect -8732 -24270 -8720 -24236
rect -9208 -24276 -8720 -24270
rect -8190 -24236 -7702 -24230
rect -8190 -24270 -8178 -24236
rect -7714 -24270 -7702 -24236
rect -8190 -24276 -7702 -24270
rect -7172 -24236 -6684 -24230
rect -7172 -24270 -7160 -24236
rect -6696 -24270 -6684 -24236
rect -7172 -24276 -6684 -24270
rect -6154 -24236 -5666 -24230
rect -6154 -24270 -6142 -24236
rect -5678 -24270 -5666 -24236
rect -6154 -24276 -5666 -24270
rect -10668 -24440 -10662 -24380
rect -10602 -24440 -10596 -24380
rect -10524 -24390 -9446 -24330
rect -7992 -24380 -7932 -24276
rect -6960 -24380 -6900 -24276
rect -9506 -24510 -9446 -24390
rect -7998 -24440 -7992 -24380
rect -7932 -24440 -7926 -24380
rect -6966 -24440 -6960 -24380
rect -6900 -24440 -6894 -24380
rect -5426 -24510 -5366 -24186
rect -4406 -24186 -4400 -23670
rect -4366 -23670 -4358 -23610
rect -3394 -23610 -3334 -23366
rect -2900 -23418 -2840 -23164
rect -2900 -23484 -2840 -23478
rect -2384 -23198 -2324 -23074
rect -1358 -23074 -1346 -23028
rect -1312 -22554 -1302 -22498
rect -340 -22498 -280 -22258
rect 160 -22408 220 -22258
rect -46 -22414 442 -22408
rect -46 -22448 -34 -22414
rect 430 -22448 442 -22414
rect -46 -22454 442 -22448
rect -1312 -23028 -1306 -22554
rect -1312 -23074 -1298 -23028
rect -2082 -23124 -1594 -23118
rect -2082 -23158 -2070 -23124
rect -1606 -23158 -1594 -23124
rect -2082 -23164 -1594 -23158
rect -3100 -23526 -2612 -23520
rect -3100 -23560 -3088 -23526
rect -2624 -23560 -2612 -23526
rect -3100 -23566 -2612 -23560
rect -3394 -23656 -3382 -23610
rect -4366 -24186 -4360 -23670
rect -4406 -24198 -4360 -24186
rect -3388 -24186 -3382 -23656
rect -3348 -23656 -3334 -23610
rect -2384 -23610 -2324 -23258
rect -1358 -23306 -1298 -23074
rect -340 -23074 -328 -22498
rect -294 -23074 -280 -22498
rect -1064 -23124 -576 -23118
rect -1064 -23158 -1052 -23124
rect -588 -23158 -576 -23124
rect -1064 -23164 -576 -23158
rect -340 -23198 -280 -23074
rect 676 -22498 736 -22258
rect 676 -23074 690 -22498
rect 724 -23074 736 -22498
rect -46 -23124 442 -23118
rect -46 -23158 -34 -23124
rect 430 -23158 442 -23124
rect -46 -23164 442 -23158
rect -346 -23258 -340 -23198
rect -280 -23258 -274 -23198
rect -1364 -23366 -1358 -23306
rect -1298 -23366 -1292 -23306
rect -340 -23310 -280 -23258
rect 168 -23310 228 -23164
rect 676 -23310 736 -23074
rect -340 -23370 736 -23310
rect -868 -23418 -808 -23412
rect -1892 -23478 -1886 -23418
rect -1826 -23478 -1820 -23418
rect -1886 -23520 -1826 -23478
rect -868 -23520 -808 -23478
rect -2082 -23526 -1594 -23520
rect -2082 -23560 -2070 -23526
rect -1606 -23560 -1594 -23526
rect -2082 -23566 -1594 -23560
rect -1064 -23526 -576 -23520
rect -1064 -23560 -1052 -23526
rect -588 -23560 -576 -23526
rect -1064 -23566 -576 -23560
rect -2384 -23652 -2364 -23610
rect -3348 -24186 -3342 -23656
rect -3388 -24198 -3342 -24186
rect -2370 -24186 -2364 -23652
rect -2330 -24186 -2324 -23610
rect -1352 -23610 -1306 -23598
rect -1352 -24158 -1346 -23610
rect -2370 -24198 -2324 -24186
rect -1366 -24186 -1346 -24158
rect -1312 -24186 -1306 -23610
rect -340 -23610 -280 -23370
rect 168 -23520 228 -23370
rect -46 -23526 442 -23520
rect -46 -23560 -34 -23526
rect 430 -23560 442 -23526
rect -46 -23566 442 -23560
rect -340 -23674 -328 -23610
rect -5136 -24236 -4648 -24230
rect -5136 -24270 -5124 -24236
rect -4660 -24270 -4648 -24236
rect -5136 -24276 -4648 -24270
rect -4118 -24236 -3630 -24230
rect -4118 -24270 -4106 -24236
rect -3642 -24270 -3630 -24236
rect -4118 -24276 -3630 -24270
rect -3100 -24236 -2612 -24230
rect -3100 -24270 -3088 -24236
rect -2624 -24270 -2612 -24236
rect -3100 -24276 -2612 -24270
rect -2082 -24236 -1594 -24230
rect -2082 -24270 -2070 -24236
rect -1606 -24270 -1594 -24236
rect -2082 -24276 -1594 -24270
rect -3900 -24380 -3840 -24276
rect -2904 -24380 -2844 -24276
rect -3906 -24440 -3900 -24380
rect -3840 -24440 -3834 -24380
rect -2910 -24440 -2904 -24380
rect -2844 -24440 -2838 -24380
rect -1366 -24510 -1306 -24186
rect -334 -24186 -328 -23674
rect -294 -23674 -280 -23610
rect 676 -23610 736 -23370
rect 676 -23652 690 -23610
rect -294 -24186 -288 -23674
rect -334 -24198 -288 -24186
rect 684 -24186 690 -23652
rect 724 -23652 736 -23610
rect 724 -24186 730 -23652
rect 684 -24198 730 -24186
rect -1064 -24236 -576 -24230
rect -1064 -24270 -1052 -24236
rect -588 -24270 -576 -24236
rect -1064 -24276 -576 -24270
rect -46 -24236 442 -24230
rect -46 -24270 -34 -24236
rect 430 -24270 442 -24236
rect -46 -24276 442 -24270
rect 816 -24510 876 -22194
rect 936 -23418 996 -21044
rect 930 -23478 936 -23418
rect 996 -23478 1002 -23418
rect -5432 -24570 -5426 -24510
rect -5366 -24570 -5360 -24510
rect -1372 -24570 -1366 -24510
rect -1306 -24570 -1300 -24510
rect 810 -24570 816 -24510
rect 876 -24570 882 -24510
rect -9506 -24576 -9446 -24570
rect -10064 -24976 172 -24916
rect -10064 -25152 -10004 -24976
rect -9564 -25062 -9504 -24976
rect -9768 -25068 -9280 -25062
rect -9768 -25102 -9756 -25068
rect -9292 -25102 -9280 -25068
rect -9768 -25108 -9280 -25102
rect -10064 -25186 -10050 -25152
rect -10056 -25728 -10050 -25186
rect -10016 -25186 -10004 -25152
rect -9042 -25152 -8982 -24976
rect -8544 -25062 -8484 -24976
rect -7510 -25062 -7450 -24976
rect -6488 -25062 -6428 -24976
rect -5498 -25062 -5438 -24976
rect -8750 -25068 -8262 -25062
rect -8750 -25102 -8738 -25068
rect -8274 -25102 -8262 -25068
rect -8750 -25108 -8262 -25102
rect -7732 -25068 -7244 -25062
rect -7732 -25102 -7720 -25068
rect -7256 -25102 -7244 -25068
rect -7732 -25108 -7244 -25102
rect -6714 -25068 -6226 -25062
rect -6714 -25102 -6702 -25068
rect -6238 -25102 -6226 -25068
rect -6714 -25108 -6226 -25102
rect -5696 -25068 -5208 -25062
rect -5696 -25102 -5684 -25068
rect -5220 -25102 -5208 -25068
rect -5696 -25108 -5208 -25102
rect -10016 -25728 -10010 -25186
rect -9042 -25196 -9032 -25152
rect -10056 -25740 -10010 -25728
rect -9038 -25728 -9032 -25196
rect -8998 -25196 -8982 -25152
rect -8020 -25152 -7974 -25140
rect -8998 -25728 -8992 -25196
rect -8020 -25670 -8014 -25152
rect -9038 -25740 -8992 -25728
rect -8028 -25728 -8014 -25670
rect -7980 -25670 -7974 -25152
rect -7002 -25152 -6956 -25140
rect -7980 -25728 -7968 -25670
rect -7002 -25694 -6996 -25152
rect -9768 -25778 -9280 -25772
rect -9768 -25812 -9756 -25778
rect -9292 -25812 -9280 -25778
rect -9768 -25818 -9280 -25812
rect -8750 -25778 -8262 -25772
rect -8750 -25812 -8738 -25778
rect -8274 -25812 -8262 -25778
rect -8750 -25818 -8262 -25812
rect -8028 -25876 -7968 -25728
rect -7010 -25728 -6996 -25694
rect -6962 -25694 -6956 -25152
rect -5984 -25152 -5938 -25140
rect -5984 -25682 -5978 -25152
rect -6962 -25728 -6950 -25694
rect -7732 -25778 -7244 -25772
rect -7732 -25812 -7720 -25778
rect -7256 -25812 -7244 -25778
rect -7732 -25818 -7244 -25812
rect -8034 -25936 -8028 -25876
rect -7968 -25936 -7962 -25876
rect -12328 -27116 -12216 -26330
rect -8028 -26430 -7968 -25936
rect -7010 -25988 -6950 -25728
rect -5990 -25728 -5978 -25682
rect -5944 -25682 -5938 -25152
rect -4974 -25152 -4914 -24976
rect -4464 -25062 -4404 -24976
rect -3474 -25062 -3414 -24976
rect -2442 -25062 -2382 -24976
rect -1438 -25062 -1378 -24976
rect -4678 -25068 -4190 -25062
rect -4678 -25102 -4666 -25068
rect -4202 -25102 -4190 -25068
rect -4678 -25108 -4190 -25102
rect -3660 -25068 -3172 -25062
rect -3660 -25102 -3648 -25068
rect -3184 -25102 -3172 -25068
rect -3660 -25108 -3172 -25102
rect -2642 -25068 -2154 -25062
rect -2642 -25102 -2630 -25068
rect -2166 -25102 -2154 -25068
rect -2642 -25108 -2154 -25102
rect -1624 -25068 -1136 -25062
rect -1624 -25102 -1612 -25068
rect -1148 -25102 -1136 -25068
rect -1624 -25108 -1136 -25102
rect -4464 -25110 -4404 -25108
rect -2442 -25110 -2382 -25108
rect -4974 -25194 -4960 -25152
rect -5944 -25728 -5930 -25682
rect -6714 -25778 -6226 -25772
rect -6714 -25812 -6702 -25778
rect -6238 -25812 -6226 -25778
rect -6714 -25818 -6226 -25812
rect -5990 -25876 -5930 -25728
rect -4966 -25728 -4960 -25194
rect -4926 -25194 -4914 -25152
rect -3948 -25152 -3902 -25140
rect -4926 -25728 -4920 -25194
rect -3948 -25682 -3942 -25152
rect -4966 -25740 -4920 -25728
rect -3954 -25728 -3942 -25682
rect -3908 -25682 -3902 -25152
rect -2930 -25152 -2884 -25140
rect -3908 -25728 -3894 -25682
rect -2930 -25690 -2924 -25152
rect -5696 -25778 -5208 -25772
rect -5696 -25812 -5684 -25778
rect -5220 -25812 -5208 -25778
rect -5696 -25818 -5208 -25812
rect -4678 -25778 -4190 -25772
rect -4678 -25812 -4666 -25778
rect -4202 -25812 -4190 -25778
rect -4678 -25818 -4190 -25812
rect -3954 -25876 -3894 -25728
rect -2936 -25728 -2924 -25690
rect -2890 -25690 -2884 -25152
rect -1912 -25152 -1866 -25140
rect -2890 -25728 -2876 -25690
rect -1912 -25696 -1906 -25152
rect -3660 -25778 -3172 -25772
rect -3660 -25812 -3648 -25778
rect -3184 -25812 -3172 -25778
rect -3660 -25818 -3172 -25812
rect -5996 -25936 -5990 -25876
rect -5930 -25936 -5924 -25876
rect -3960 -25936 -3954 -25876
rect -3894 -25936 -3888 -25876
rect -7016 -26048 -7010 -25988
rect -6950 -26048 -6944 -25988
rect -5990 -26430 -5930 -25936
rect -3954 -26430 -3894 -25936
rect -2936 -25988 -2876 -25728
rect -1918 -25728 -1906 -25696
rect -1872 -25696 -1866 -25152
rect -898 -25152 -838 -24976
rect -418 -25062 -358 -24976
rect -606 -25068 -118 -25062
rect -606 -25102 -594 -25068
rect -130 -25102 -118 -25068
rect -606 -25108 -118 -25102
rect -898 -25220 -888 -25152
rect -1872 -25728 -1858 -25696
rect -2642 -25778 -2154 -25772
rect -2642 -25812 -2630 -25778
rect -2166 -25812 -2154 -25778
rect -2642 -25818 -2154 -25812
rect -1918 -25876 -1858 -25728
rect -894 -25728 -888 -25220
rect -854 -25220 -838 -25152
rect 112 -25152 172 -24976
rect 112 -25192 130 -25152
rect -854 -25728 -848 -25220
rect -894 -25740 -848 -25728
rect 124 -25728 130 -25192
rect 164 -25192 172 -25152
rect 164 -25728 170 -25192
rect 124 -25740 170 -25728
rect -1624 -25778 -1136 -25772
rect -1624 -25812 -1612 -25778
rect -1148 -25812 -1136 -25778
rect -1624 -25818 -1136 -25812
rect -606 -25778 -118 -25772
rect -606 -25812 -594 -25778
rect -130 -25812 -118 -25778
rect -606 -25818 -118 -25812
rect -1924 -25936 -1918 -25876
rect -1858 -25936 -1852 -25876
rect -2942 -26048 -2936 -25988
rect -2876 -26048 -2870 -25988
rect -1918 -26430 -1858 -25936
rect 1070 -25988 1130 -19060
rect 1282 -19894 1342 -11554
rect 1276 -19954 1282 -19894
rect 1342 -19954 1348 -19894
rect 1402 -20022 1462 -11552
rect 1396 -20082 1402 -20022
rect 1462 -20082 1468 -20022
rect 1542 -20984 1602 -11534
rect 1654 -11672 1660 -11612
rect 1720 -11672 1726 -11612
rect 1660 -17740 1720 -11672
rect 1770 -12354 1830 -11518
rect 1764 -12414 1770 -12354
rect 1830 -12414 1836 -12354
rect 1888 -15274 1948 -11418
rect 2216 -12220 2276 -11408
rect 2210 -12280 2216 -12220
rect 2276 -12280 2282 -12220
rect 2006 -13638 2012 -13578
rect 2072 -13638 2078 -13578
rect 1886 -15280 1948 -15274
rect 1946 -15340 1948 -15280
rect 1886 -15346 1948 -15340
rect 1654 -17800 1660 -17740
rect 1720 -17800 1726 -17740
rect 1536 -21044 1542 -20984
rect 1602 -21044 1608 -20984
rect 1888 -21342 1948 -15346
rect 2012 -16274 2072 -13638
rect 2218 -13974 2224 -13914
rect 2284 -13974 2290 -13914
rect 2114 -15234 2120 -15174
rect 2180 -15234 2186 -15174
rect 2006 -16334 2012 -16274
rect 2072 -16334 2078 -16274
rect 2120 -21192 2180 -15234
rect 2224 -16510 2284 -13974
rect 2336 -16396 2396 -11416
rect 2442 -11492 2502 -11486
rect 2442 -14036 2502 -11552
rect 13248 -11848 13254 -11842
rect 2568 -11902 13254 -11848
rect 13314 -11848 13320 -11842
rect 18352 -11848 18358 -11842
rect 13314 -11902 18358 -11848
rect 18418 -11848 18424 -11842
rect 22418 -11848 22478 -11842
rect 18418 -11902 22418 -11848
rect 2568 -11908 22418 -11902
rect 22478 -11908 22990 -11848
rect 2568 -12048 2628 -11908
rect 3090 -11958 3150 -11908
rect 4100 -11958 4160 -11908
rect 2864 -11964 3352 -11958
rect 2864 -11998 2876 -11964
rect 3340 -11998 3352 -11964
rect 2864 -12004 3352 -11998
rect 3882 -11964 4370 -11958
rect 3882 -11998 3894 -11964
rect 4358 -11998 4370 -11964
rect 3882 -12004 4370 -11998
rect 4100 -12010 4160 -12004
rect 2568 -12624 2582 -12048
rect 2616 -12624 2628 -12048
rect 3594 -12048 3640 -12036
rect 3594 -12590 3600 -12048
rect 2568 -12866 2628 -12624
rect 3586 -12624 3600 -12590
rect 3634 -12590 3640 -12048
rect 4606 -12048 4666 -11908
rect 5130 -11958 5190 -11908
rect 6142 -11958 6202 -11908
rect 4900 -11964 5388 -11958
rect 4900 -11998 4912 -11964
rect 5376 -11998 5388 -11964
rect 4900 -12004 5388 -11998
rect 5918 -11964 6406 -11958
rect 5918 -11998 5930 -11964
rect 6394 -11998 6406 -11964
rect 5918 -12004 6406 -11998
rect 6142 -12010 6202 -12004
rect 3634 -12624 3646 -12590
rect 2864 -12674 3352 -12668
rect 2864 -12708 2876 -12674
rect 3340 -12708 3352 -12674
rect 2864 -12714 3352 -12708
rect 3080 -12776 3140 -12714
rect 2864 -12782 3352 -12776
rect 2864 -12816 2876 -12782
rect 3340 -12816 3352 -12782
rect 2864 -12822 3352 -12816
rect 3080 -12828 3140 -12822
rect 2568 -13442 2582 -12866
rect 2616 -13442 2628 -12866
rect 2568 -13914 2628 -13442
rect 3586 -12866 3646 -12624
rect 4606 -12624 4618 -12048
rect 4652 -12624 4666 -12048
rect 5630 -12048 5676 -12036
rect 5630 -12578 5636 -12048
rect 4086 -12668 4146 -12666
rect 3882 -12674 4370 -12668
rect 3882 -12708 3894 -12674
rect 4358 -12708 4370 -12674
rect 3882 -12714 4370 -12708
rect 4086 -12776 4146 -12714
rect 3882 -12782 4370 -12776
rect 3882 -12816 3894 -12782
rect 4358 -12816 4370 -12782
rect 3882 -12822 4370 -12816
rect 3586 -13442 3600 -12866
rect 3634 -13442 3646 -12866
rect 4606 -12866 4666 -12624
rect 5620 -12624 5636 -12578
rect 5670 -12578 5676 -12048
rect 6638 -12048 6698 -11908
rect 7154 -11958 7214 -11908
rect 8154 -11958 8214 -11908
rect 6936 -11964 7424 -11958
rect 6936 -11998 6948 -11964
rect 7412 -11998 7424 -11964
rect 6936 -12004 7424 -11998
rect 7954 -11964 8442 -11958
rect 7954 -11998 7966 -11964
rect 8430 -11998 8442 -11964
rect 7954 -12004 8442 -11998
rect 5670 -12624 5680 -12578
rect 5098 -12668 5158 -12660
rect 4900 -12674 5388 -12668
rect 4900 -12708 4912 -12674
rect 5376 -12708 5388 -12674
rect 4900 -12714 5388 -12708
rect 5098 -12776 5158 -12714
rect 4900 -12782 5388 -12776
rect 4900 -12816 4912 -12782
rect 5376 -12816 5388 -12782
rect 4900 -12822 5388 -12816
rect 4606 -12924 4618 -12866
rect 2864 -13492 3352 -13486
rect 2864 -13526 2876 -13492
rect 3340 -13526 3352 -13492
rect 2864 -13532 3352 -13526
rect 3586 -13578 3646 -13442
rect 4612 -13442 4618 -12924
rect 4652 -12924 4666 -12866
rect 5620 -12866 5680 -12624
rect 6638 -12624 6654 -12048
rect 6688 -12624 6698 -12048
rect 7666 -12048 7712 -12036
rect 7666 -12584 7672 -12048
rect 5918 -12674 6406 -12668
rect 5918 -12708 5930 -12674
rect 6394 -12708 6406 -12674
rect 5918 -12714 6406 -12708
rect 6120 -12776 6180 -12714
rect 5918 -12782 6406 -12776
rect 5918 -12816 5930 -12782
rect 6394 -12816 6406 -12782
rect 5918 -12822 6406 -12816
rect 6120 -12828 6180 -12822
rect 4652 -13442 4658 -12924
rect 4612 -13454 4658 -13442
rect 5620 -13442 5636 -12866
rect 5670 -13442 5680 -12866
rect 6638 -12866 6698 -12624
rect 7656 -12624 7672 -12584
rect 7706 -12584 7712 -12048
rect 8676 -12048 8736 -11908
rect 9188 -11958 9248 -11908
rect 10200 -11958 10260 -11908
rect 8972 -11964 9460 -11958
rect 8972 -11998 8984 -11964
rect 9448 -11998 9460 -11964
rect 8972 -12004 9460 -11998
rect 9990 -11964 10478 -11958
rect 9990 -11998 10002 -11964
rect 10466 -11998 10478 -11964
rect 9990 -12004 10478 -11998
rect 7706 -12624 7716 -12584
rect 6936 -12674 7424 -12668
rect 6936 -12708 6948 -12674
rect 7412 -12708 7424 -12674
rect 6936 -12714 7424 -12708
rect 7132 -12776 7192 -12714
rect 6936 -12782 7424 -12776
rect 6936 -12816 6948 -12782
rect 7412 -12816 7424 -12782
rect 6936 -12822 7424 -12816
rect 7132 -12828 7192 -12822
rect 6638 -12928 6654 -12866
rect 3882 -13492 4370 -13486
rect 3882 -13526 3894 -13492
rect 4358 -13526 4370 -13492
rect 3882 -13532 4370 -13526
rect 4900 -13492 5388 -13486
rect 4900 -13526 4912 -13492
rect 5376 -13526 5388 -13492
rect 4900 -13532 5388 -13526
rect 5620 -13580 5680 -13442
rect 6648 -13442 6654 -12928
rect 6688 -12928 6698 -12866
rect 7656 -12866 7716 -12624
rect 8676 -12624 8690 -12048
rect 8724 -12624 8736 -12048
rect 9702 -12048 9748 -12036
rect 9702 -12584 9708 -12048
rect 7954 -12674 8442 -12668
rect 7954 -12708 7966 -12674
rect 8430 -12708 8442 -12674
rect 7954 -12714 8442 -12708
rect 8162 -12776 8222 -12714
rect 7954 -12782 8442 -12776
rect 7954 -12816 7966 -12782
rect 8430 -12816 8442 -12782
rect 7954 -12822 8442 -12816
rect 8162 -12828 8222 -12822
rect 6688 -13442 6694 -12928
rect 6648 -13454 6694 -13442
rect 7656 -13442 7672 -12866
rect 7706 -13442 7716 -12866
rect 8676 -12866 8736 -12624
rect 9694 -12624 9708 -12584
rect 9742 -12584 9748 -12048
rect 10712 -12048 10772 -11908
rect 11224 -11958 11284 -11908
rect 12236 -11958 12296 -11908
rect 11008 -11964 11496 -11958
rect 11008 -11998 11020 -11964
rect 11484 -11998 11496 -11964
rect 11008 -12004 11496 -11998
rect 12026 -11964 12514 -11958
rect 12026 -11998 12038 -11964
rect 12502 -11998 12514 -11964
rect 12026 -12004 12514 -11998
rect 9742 -12624 9754 -12584
rect 9168 -12668 9228 -12666
rect 8972 -12674 9460 -12668
rect 8972 -12708 8984 -12674
rect 9448 -12708 9460 -12674
rect 8972 -12714 9460 -12708
rect 9168 -12776 9228 -12714
rect 8972 -12782 9460 -12776
rect 8972 -12816 8984 -12782
rect 9448 -12816 9460 -12782
rect 8972 -12822 9460 -12816
rect 8676 -12908 8690 -12866
rect 5918 -13492 6406 -13486
rect 5918 -13526 5930 -13492
rect 6394 -13526 6406 -13492
rect 5918 -13532 6406 -13526
rect 6936 -13492 7424 -13486
rect 6936 -13526 6948 -13492
rect 7412 -13526 7424 -13492
rect 6936 -13532 7424 -13526
rect 7656 -13580 7716 -13442
rect 8684 -13442 8690 -12908
rect 8724 -12908 8736 -12866
rect 9694 -12866 9754 -12624
rect 10712 -12624 10726 -12048
rect 10760 -12624 10772 -12048
rect 11738 -12048 11784 -12036
rect 11738 -12578 11744 -12048
rect 10190 -12668 10250 -12666
rect 9990 -12674 10478 -12668
rect 9990 -12708 10002 -12674
rect 10466 -12708 10478 -12674
rect 9990 -12714 10478 -12708
rect 10190 -12776 10250 -12714
rect 9990 -12782 10478 -12776
rect 9990 -12816 10002 -12782
rect 10466 -12816 10478 -12782
rect 9990 -12822 10478 -12816
rect 8724 -13442 8730 -12908
rect 8684 -13454 8730 -13442
rect 9694 -13442 9708 -12866
rect 9742 -13442 9754 -12866
rect 10712 -12866 10772 -12624
rect 11732 -12624 11744 -12578
rect 11778 -12578 11784 -12048
rect 12744 -12048 12804 -11908
rect 13258 -11958 13318 -11908
rect 14270 -11958 14330 -11908
rect 13044 -11964 13532 -11958
rect 13044 -11998 13056 -11964
rect 13520 -11998 13532 -11964
rect 13044 -12004 13532 -11998
rect 14062 -11964 14550 -11958
rect 14062 -11998 14074 -11964
rect 14538 -11998 14550 -11964
rect 14062 -12004 14550 -11998
rect 14270 -12010 14330 -12004
rect 11778 -12624 11792 -12578
rect 11008 -12674 11496 -12668
rect 11008 -12708 11020 -12674
rect 11484 -12708 11496 -12674
rect 11008 -12714 11496 -12708
rect 11214 -12776 11274 -12714
rect 11008 -12782 11496 -12776
rect 11008 -12816 11020 -12782
rect 11484 -12816 11496 -12782
rect 11008 -12822 11496 -12816
rect 11214 -12828 11274 -12822
rect 10712 -12916 10726 -12866
rect 7954 -13492 8442 -13486
rect 7954 -13526 7966 -13492
rect 8430 -13526 8442 -13492
rect 7954 -13532 8442 -13526
rect 8972 -13492 9460 -13486
rect 8972 -13526 8984 -13492
rect 9448 -13526 9460 -13492
rect 8972 -13532 9460 -13526
rect 9694 -13580 9754 -13442
rect 10720 -13442 10726 -12916
rect 10760 -12916 10772 -12866
rect 11732 -12866 11792 -12624
rect 12744 -12624 12762 -12048
rect 12796 -12624 12804 -12048
rect 13774 -12048 13820 -12036
rect 13774 -12578 13780 -12048
rect 12220 -12668 12280 -12666
rect 12026 -12674 12514 -12668
rect 12026 -12708 12038 -12674
rect 12502 -12708 12514 -12674
rect 12026 -12714 12514 -12708
rect 12220 -12776 12280 -12714
rect 12026 -12782 12514 -12776
rect 12026 -12816 12038 -12782
rect 12502 -12816 12514 -12782
rect 12026 -12822 12514 -12816
rect 10760 -13442 10766 -12916
rect 10720 -13454 10766 -13442
rect 11732 -13442 11744 -12866
rect 11778 -13442 11792 -12866
rect 12744 -12866 12804 -12624
rect 13766 -12624 13780 -12578
rect 13814 -12578 13820 -12048
rect 14782 -12048 14842 -11908
rect 15294 -11958 15354 -11908
rect 16312 -11958 16372 -11908
rect 15080 -11964 15568 -11958
rect 15080 -11998 15092 -11964
rect 15556 -11998 15568 -11964
rect 15080 -12004 15568 -11998
rect 16098 -11964 16586 -11958
rect 16098 -11998 16110 -11964
rect 16574 -11998 16586 -11964
rect 16098 -12004 16586 -11998
rect 15294 -12010 15354 -12004
rect 13814 -12624 13826 -12578
rect 13244 -12668 13304 -12660
rect 13044 -12674 13532 -12668
rect 13044 -12708 13056 -12674
rect 13520 -12708 13532 -12674
rect 13044 -12714 13532 -12708
rect 13244 -12776 13304 -12714
rect 13044 -12782 13532 -12776
rect 13044 -12816 13056 -12782
rect 13520 -12816 13532 -12782
rect 13044 -12822 13532 -12816
rect 12744 -12914 12762 -12866
rect 9990 -13492 10478 -13486
rect 9990 -13526 10002 -13492
rect 10466 -13526 10478 -13492
rect 9990 -13532 10478 -13526
rect 11008 -13492 11496 -13486
rect 11008 -13526 11020 -13492
rect 11484 -13526 11496 -13492
rect 11008 -13532 11496 -13526
rect 11732 -13580 11792 -13442
rect 12756 -13442 12762 -12914
rect 12796 -12914 12804 -12866
rect 13766 -12866 13826 -12624
rect 14782 -12624 14798 -12048
rect 14832 -12624 14842 -12048
rect 15810 -12048 15856 -12036
rect 15810 -12578 15816 -12048
rect 14266 -12668 14326 -12666
rect 14062 -12674 14550 -12668
rect 14062 -12708 14074 -12674
rect 14538 -12708 14550 -12674
rect 14062 -12714 14550 -12708
rect 14266 -12776 14326 -12714
rect 14062 -12782 14550 -12776
rect 14062 -12816 14074 -12782
rect 14538 -12816 14550 -12782
rect 14062 -12822 14550 -12816
rect 12796 -13442 12802 -12914
rect 12756 -13454 12802 -13442
rect 13766 -13442 13780 -12866
rect 13814 -13442 13826 -12866
rect 14782 -12866 14842 -12624
rect 15802 -12624 15816 -12578
rect 15850 -12578 15856 -12048
rect 16818 -12048 16878 -11908
rect 17334 -11958 17394 -11908
rect 18358 -11958 18418 -11908
rect 17116 -11964 17604 -11958
rect 17116 -11998 17128 -11964
rect 17592 -11998 17604 -11964
rect 17116 -12004 17604 -11998
rect 18134 -11964 18622 -11958
rect 18134 -11998 18146 -11964
rect 18610 -11998 18622 -11964
rect 18134 -12004 18622 -11998
rect 15850 -12624 15862 -12578
rect 15278 -12668 15338 -12666
rect 15080 -12674 15568 -12668
rect 15080 -12708 15092 -12674
rect 15556 -12708 15568 -12674
rect 15080 -12714 15568 -12708
rect 15278 -12776 15338 -12714
rect 15080 -12782 15568 -12776
rect 15080 -12816 15092 -12782
rect 15556 -12816 15568 -12782
rect 15080 -12822 15568 -12816
rect 14782 -12916 14798 -12866
rect 12026 -13492 12514 -13486
rect 12026 -13526 12038 -13492
rect 12502 -13526 12514 -13492
rect 12026 -13532 12514 -13526
rect 13044 -13492 13532 -13486
rect 13044 -13526 13056 -13492
rect 13520 -13526 13532 -13492
rect 13044 -13532 13532 -13526
rect 13766 -13580 13826 -13442
rect 14792 -13442 14798 -12916
rect 14832 -12916 14842 -12866
rect 15802 -12866 15862 -12624
rect 16818 -12624 16834 -12048
rect 16868 -12624 16878 -12048
rect 17846 -12048 17892 -12036
rect 17846 -12554 17852 -12048
rect 16098 -12674 16586 -12668
rect 16098 -12708 16110 -12674
rect 16574 -12708 16586 -12674
rect 16098 -12714 16586 -12708
rect 16290 -12776 16350 -12714
rect 16098 -12782 16586 -12776
rect 16098 -12816 16110 -12782
rect 16574 -12816 16586 -12782
rect 16098 -12822 16586 -12816
rect 16290 -12828 16350 -12822
rect 14832 -13442 14838 -12916
rect 14792 -13454 14838 -13442
rect 15802 -13442 15816 -12866
rect 15850 -13442 15862 -12866
rect 16818 -12866 16878 -12624
rect 17840 -12624 17852 -12554
rect 17886 -12554 17892 -12048
rect 18854 -12048 18914 -11908
rect 19376 -11958 19436 -11908
rect 20388 -11958 20448 -11908
rect 19152 -11964 19640 -11958
rect 19152 -11998 19164 -11964
rect 19628 -11998 19640 -11964
rect 19152 -12004 19640 -11998
rect 20170 -11964 20658 -11958
rect 20170 -11998 20182 -11964
rect 20646 -11998 20658 -11964
rect 20170 -12004 20658 -11998
rect 17886 -12624 17900 -12554
rect 17314 -12668 17374 -12660
rect 17116 -12674 17604 -12668
rect 17116 -12708 17128 -12674
rect 17592 -12708 17604 -12674
rect 17116 -12714 17604 -12708
rect 17314 -12776 17374 -12714
rect 17116 -12782 17604 -12776
rect 17116 -12816 17128 -12782
rect 17592 -12816 17604 -12782
rect 17116 -12822 17604 -12816
rect 16818 -12890 16834 -12866
rect 14062 -13492 14550 -13486
rect 14062 -13526 14074 -13492
rect 14538 -13526 14550 -13492
rect 14062 -13532 14550 -13526
rect 15080 -13492 15568 -13486
rect 15080 -13526 15092 -13492
rect 15556 -13526 15568 -13492
rect 15080 -13532 15568 -13526
rect 15802 -13580 15862 -13442
rect 16828 -13442 16834 -12890
rect 16868 -12890 16878 -12866
rect 17840 -12866 17900 -12624
rect 18854 -12624 18870 -12048
rect 18904 -12624 18914 -12048
rect 19882 -12048 19928 -12036
rect 19882 -12514 19888 -12048
rect 18134 -12674 18622 -12668
rect 18134 -12708 18146 -12674
rect 18610 -12708 18622 -12674
rect 18134 -12714 18622 -12708
rect 18336 -12776 18396 -12714
rect 18134 -12782 18622 -12776
rect 18134 -12816 18146 -12782
rect 18610 -12816 18622 -12782
rect 18134 -12822 18622 -12816
rect 18336 -12834 18396 -12822
rect 16868 -13442 16874 -12890
rect 16828 -13454 16874 -13442
rect 17840 -13442 17852 -12866
rect 17886 -13442 17900 -12866
rect 18854 -12866 18914 -12624
rect 19874 -12624 19888 -12514
rect 19922 -12514 19928 -12048
rect 20892 -12048 20952 -11908
rect 21398 -11958 21458 -11908
rect 22416 -11914 22478 -11908
rect 22416 -11958 22476 -11914
rect 21188 -11964 21676 -11958
rect 21188 -11998 21200 -11964
rect 21664 -11998 21676 -11964
rect 21188 -12004 21676 -11998
rect 22206 -11964 22694 -11958
rect 22206 -11998 22218 -11964
rect 22682 -11998 22694 -11964
rect 22206 -12004 22694 -11998
rect 19922 -12624 19934 -12514
rect 19354 -12668 19414 -12666
rect 19152 -12674 19640 -12668
rect 19152 -12708 19164 -12674
rect 19628 -12708 19640 -12674
rect 19152 -12714 19640 -12708
rect 19354 -12776 19414 -12714
rect 19152 -12782 19640 -12776
rect 19152 -12816 19164 -12782
rect 19628 -12816 19640 -12782
rect 19152 -12822 19640 -12816
rect 18854 -12908 18870 -12866
rect 16098 -13492 16586 -13486
rect 16098 -13526 16110 -13492
rect 16574 -13526 16586 -13492
rect 16098 -13532 16586 -13526
rect 17116 -13492 17604 -13486
rect 17116 -13526 17128 -13492
rect 17592 -13526 17604 -13492
rect 17116 -13532 17604 -13526
rect 17840 -13580 17900 -13442
rect 18864 -13442 18870 -12908
rect 18904 -12908 18914 -12866
rect 19874 -12866 19934 -12624
rect 20892 -12624 20906 -12048
rect 20940 -12624 20952 -12048
rect 21918 -12048 21964 -12036
rect 21918 -12564 21924 -12048
rect 20384 -12668 20444 -12654
rect 20170 -12674 20658 -12668
rect 20170 -12708 20182 -12674
rect 20646 -12708 20658 -12674
rect 20170 -12714 20658 -12708
rect 20384 -12776 20444 -12714
rect 20170 -12782 20658 -12776
rect 20170 -12816 20182 -12782
rect 20646 -12816 20658 -12782
rect 20170 -12822 20658 -12816
rect 18904 -13442 18910 -12908
rect 18864 -13454 18910 -13442
rect 19874 -13442 19888 -12866
rect 19922 -13442 19934 -12866
rect 20892 -12866 20952 -12624
rect 21910 -12624 21924 -12564
rect 21958 -12564 21964 -12048
rect 22930 -12048 22990 -11908
rect 21958 -12624 21970 -12564
rect 21396 -12668 21456 -12654
rect 21188 -12674 21676 -12668
rect 21188 -12708 21200 -12674
rect 21664 -12708 21676 -12674
rect 21188 -12714 21676 -12708
rect 21396 -12776 21456 -12714
rect 21188 -12782 21676 -12776
rect 21188 -12816 21200 -12782
rect 21664 -12816 21676 -12782
rect 21188 -12822 21676 -12816
rect 20892 -12908 20906 -12866
rect 18134 -13492 18622 -13486
rect 18134 -13526 18146 -13492
rect 18610 -13526 18622 -13492
rect 18134 -13532 18622 -13526
rect 19152 -13492 19640 -13486
rect 19152 -13526 19164 -13492
rect 19628 -13526 19640 -13492
rect 19152 -13532 19640 -13526
rect 19874 -13580 19934 -13442
rect 20900 -13442 20906 -12908
rect 20940 -12908 20952 -12866
rect 21910 -12866 21970 -12624
rect 22930 -12624 22942 -12048
rect 22976 -12624 22990 -12048
rect 22206 -12674 22694 -12668
rect 22206 -12708 22218 -12674
rect 22682 -12708 22694 -12674
rect 22206 -12714 22694 -12708
rect 22396 -12776 22456 -12714
rect 22930 -12716 22990 -12624
rect 24816 -12070 24928 -11284
rect 22930 -12776 23710 -12716
rect 22206 -12782 22694 -12776
rect 22206 -12816 22218 -12782
rect 22682 -12816 22694 -12782
rect 22206 -12822 22694 -12816
rect 22396 -12828 22456 -12822
rect 20940 -13442 20946 -12908
rect 20900 -13454 20946 -13442
rect 21910 -13442 21924 -12866
rect 21958 -13442 21970 -12866
rect 22930 -12866 22990 -12776
rect 22930 -12916 22942 -12866
rect 20170 -13492 20658 -13486
rect 20170 -13526 20182 -13492
rect 20646 -13526 20658 -13492
rect 20170 -13532 20658 -13526
rect 21188 -13492 21676 -13486
rect 21188 -13526 21200 -13492
rect 21664 -13526 21676 -13492
rect 21188 -13532 21676 -13526
rect 21910 -13580 21970 -13442
rect 22936 -13442 22942 -12916
rect 22976 -12916 22990 -12866
rect 22976 -13442 22982 -12916
rect 22936 -13454 22982 -13442
rect 22206 -13492 22694 -13486
rect 22206 -13526 22218 -13492
rect 22682 -13526 22694 -13492
rect 22206 -13532 22694 -13526
rect 3646 -13638 23588 -13580
rect 3586 -13640 23588 -13638
rect 3586 -13644 3646 -13640
rect 4594 -13854 4600 -13794
rect 4660 -13854 4666 -13794
rect 6634 -13854 6640 -13794
rect 6700 -13854 6706 -13794
rect 8674 -13854 8680 -13794
rect 8740 -13854 8746 -13794
rect 10704 -13854 10710 -13794
rect 10770 -13854 10776 -13794
rect 12744 -13854 12750 -13794
rect 12810 -13854 12816 -13794
rect 14776 -13854 14782 -13794
rect 14842 -13854 14848 -13794
rect 16816 -13854 16822 -13794
rect 16882 -13854 16888 -13794
rect 18852 -13854 18858 -13794
rect 18918 -13854 18924 -13794
rect 20886 -13854 20892 -13794
rect 20952 -13854 20958 -13794
rect 2562 -13974 2568 -13914
rect 2628 -13974 2634 -13914
rect 4086 -13980 4092 -13920
rect 4152 -13980 4158 -13920
rect 2436 -14096 2442 -14036
rect 2502 -14096 2508 -14036
rect 2442 -16170 2502 -14096
rect 4092 -14154 4152 -13980
rect 2864 -14160 3352 -14154
rect 2864 -14194 2876 -14160
rect 3340 -14194 3352 -14160
rect 2864 -14200 3352 -14194
rect 3882 -14160 4370 -14154
rect 3882 -14194 3894 -14160
rect 4358 -14194 4370 -14160
rect 3882 -14200 4370 -14194
rect 2576 -14244 2622 -14232
rect 3594 -14244 3640 -14232
rect 4600 -14244 4660 -13854
rect 5106 -13920 5166 -13914
rect 5106 -14154 5166 -13980
rect 6128 -13920 6188 -13914
rect 6128 -14154 6188 -13980
rect 4900 -14160 5388 -14154
rect 4900 -14194 4912 -14160
rect 5376 -14194 5388 -14160
rect 4900 -14200 5388 -14194
rect 5918 -14160 6406 -14154
rect 5918 -14194 5930 -14160
rect 6394 -14194 6406 -14160
rect 5918 -14200 6406 -14194
rect 5630 -14244 5676 -14232
rect 2568 -14278 2582 -14244
rect 2576 -14770 2582 -14278
rect 2568 -14820 2582 -14770
rect 2616 -14278 2628 -14244
rect 2616 -14770 2622 -14278
rect 3586 -14292 3600 -14244
rect 2616 -14820 2628 -14770
rect 3594 -14784 3600 -14292
rect 2568 -14958 2628 -14820
rect 3586 -14820 3600 -14784
rect 3634 -14292 3646 -14244
rect 3634 -14784 3640 -14292
rect 4600 -14312 4618 -14244
rect 4612 -14756 4618 -14312
rect 3634 -14820 3646 -14784
rect 2864 -14870 3352 -14864
rect 2864 -14904 2876 -14870
rect 3340 -14904 3352 -14870
rect 2864 -14910 3352 -14904
rect 3070 -14958 3130 -14910
rect 3586 -14958 3646 -14820
rect 4604 -14820 4618 -14756
rect 4652 -14276 4664 -14244
rect 4652 -14312 4660 -14276
rect 4652 -14756 4658 -14312
rect 4652 -14820 4664 -14756
rect 5630 -14774 5636 -14244
rect 5626 -14792 5636 -14774
rect 5624 -14820 5636 -14792
rect 5670 -14774 5676 -14244
rect 6640 -14244 6700 -13854
rect 7142 -13920 7202 -13914
rect 7140 -13980 7142 -13974
rect 8168 -13920 8228 -13914
rect 7140 -13986 7202 -13980
rect 8166 -13980 8168 -13974
rect 8166 -13986 8228 -13980
rect 7140 -14154 7200 -13986
rect 7650 -14096 7656 -14036
rect 7716 -14096 7722 -14036
rect 6936 -14160 7424 -14154
rect 6936 -14194 6948 -14160
rect 7412 -14194 7424 -14160
rect 6936 -14200 7424 -14194
rect 6640 -14298 6654 -14244
rect 6648 -14748 6654 -14298
rect 6644 -14772 6654 -14748
rect 5670 -14820 5686 -14774
rect 6642 -14820 6654 -14772
rect 6688 -14298 6700 -14244
rect 7656 -14244 7716 -14096
rect 8166 -14154 8226 -13986
rect 7954 -14160 8442 -14154
rect 7954 -14194 7966 -14160
rect 8430 -14194 8442 -14160
rect 7954 -14200 8442 -14194
rect 7656 -14286 7672 -14244
rect 6688 -14748 6694 -14298
rect 7666 -14744 7672 -14286
rect 6688 -14820 6704 -14748
rect 7656 -14820 7672 -14744
rect 7706 -14286 7716 -14244
rect 8680 -14244 8740 -13854
rect 9180 -13920 9240 -13914
rect 9180 -14154 9240 -13980
rect 10216 -13920 10276 -13914
rect 10216 -14154 10276 -13980
rect 8972 -14160 9460 -14154
rect 8972 -14194 8984 -14160
rect 9448 -14194 9460 -14160
rect 8972 -14200 9460 -14194
rect 9990 -14160 10478 -14154
rect 9990 -14194 10002 -14160
rect 10466 -14194 10478 -14160
rect 9990 -14200 10478 -14194
rect 9702 -14244 9748 -14232
rect 10710 -14244 10770 -13854
rect 11222 -13920 11282 -13914
rect 12230 -13980 12236 -13920
rect 12296 -13980 12302 -13920
rect 11222 -14154 11282 -13980
rect 12236 -14154 12296 -13980
rect 11008 -14160 11496 -14154
rect 11008 -14194 11020 -14160
rect 11484 -14194 11496 -14160
rect 11008 -14200 11496 -14194
rect 12026 -14160 12514 -14154
rect 12026 -14194 12038 -14160
rect 12502 -14194 12514 -14160
rect 12026 -14200 12514 -14194
rect 7706 -14744 7712 -14286
rect 8680 -14318 8690 -14244
rect 7706 -14760 7716 -14744
rect 7706 -14820 7720 -14760
rect 8684 -14764 8690 -14318
rect 8676 -14820 8690 -14764
rect 8724 -14318 8740 -14244
rect 9696 -14294 9708 -14244
rect 8724 -14764 8730 -14318
rect 9702 -14756 9708 -14294
rect 8724 -14820 8736 -14764
rect 9696 -14784 9708 -14756
rect 9694 -14820 9708 -14784
rect 9742 -14294 9756 -14244
rect 9742 -14756 9748 -14294
rect 10710 -14312 10726 -14244
rect 10720 -14744 10726 -14312
rect 9742 -14820 9756 -14756
rect 3882 -14870 4370 -14864
rect 3882 -14904 3894 -14870
rect 4358 -14904 4370 -14870
rect 3882 -14910 4370 -14904
rect 2568 -15018 3646 -14958
rect 3586 -15174 3646 -15018
rect 4096 -15068 4156 -14910
rect 4604 -14958 4664 -14820
rect 4900 -14870 5388 -14864
rect 4900 -14904 4912 -14870
rect 5376 -14904 5388 -14870
rect 4900 -14910 5388 -14904
rect 4598 -15018 4604 -14958
rect 4664 -15018 4670 -14958
rect 4090 -15128 4096 -15068
rect 4156 -15128 4162 -15068
rect 3580 -15234 3586 -15174
rect 3646 -15234 3652 -15174
rect 2566 -15340 2572 -15280
rect 2632 -15340 2638 -15280
rect 3064 -15340 3070 -15280
rect 3130 -15340 3136 -15280
rect 3576 -15340 3582 -15280
rect 3642 -15340 3648 -15280
rect 2572 -15476 2632 -15340
rect 3070 -15386 3130 -15340
rect 2864 -15392 3352 -15386
rect 2864 -15426 2876 -15392
rect 3340 -15426 3352 -15392
rect 2864 -15432 3352 -15426
rect 2572 -15516 2582 -15476
rect 2576 -16052 2582 -15516
rect 2616 -15516 2632 -15476
rect 3582 -15476 3642 -15340
rect 4096 -15386 4156 -15128
rect 3882 -15392 4370 -15386
rect 3882 -15426 3894 -15392
rect 4358 -15426 4370 -15392
rect 3882 -15432 4370 -15426
rect 2616 -16052 2622 -15516
rect 3582 -15522 3600 -15476
rect 2576 -16064 2622 -16052
rect 3594 -16052 3600 -15522
rect 3634 -15522 3642 -15476
rect 4604 -15476 4664 -15018
rect 5118 -15068 5178 -14910
rect 5112 -15128 5118 -15068
rect 5178 -15128 5184 -15068
rect 5118 -15386 5178 -15128
rect 5626 -15174 5686 -14820
rect 5918 -14870 6406 -14864
rect 5918 -14904 5930 -14870
rect 6394 -14904 6406 -14870
rect 5918 -14910 6406 -14904
rect 6132 -15068 6192 -14910
rect 6644 -14958 6704 -14820
rect 7666 -14832 7712 -14820
rect 6936 -14870 7424 -14864
rect 6936 -14904 6948 -14870
rect 7412 -14904 7424 -14870
rect 6936 -14910 7424 -14904
rect 7954 -14870 8442 -14864
rect 7954 -14904 7966 -14870
rect 8430 -14904 8442 -14870
rect 7954 -14910 8442 -14904
rect 6638 -15018 6644 -14958
rect 6704 -15018 6710 -14958
rect 6126 -15128 6132 -15068
rect 6192 -15128 6198 -15068
rect 5620 -15234 5626 -15174
rect 5686 -15234 5692 -15174
rect 6132 -15386 6192 -15128
rect 4900 -15392 5388 -15386
rect 4900 -15426 4912 -15392
rect 5376 -15426 5388 -15392
rect 4900 -15432 5388 -15426
rect 5918 -15392 6406 -15386
rect 5918 -15426 5930 -15392
rect 6394 -15426 6406 -15392
rect 5918 -15432 6406 -15426
rect 5630 -15476 5676 -15464
rect 6644 -15476 6704 -15018
rect 7146 -15068 7206 -14910
rect 8164 -15068 8224 -14910
rect 8676 -14958 8736 -14820
rect 8972 -14870 9460 -14864
rect 8972 -14904 8984 -14870
rect 9448 -14904 9460 -14870
rect 8972 -14910 9460 -14904
rect 8670 -15018 8676 -14958
rect 8736 -15018 8742 -14958
rect 7140 -15128 7146 -15068
rect 7206 -15128 7212 -15068
rect 8158 -15128 8164 -15068
rect 8224 -15128 8230 -15068
rect 7146 -15386 7206 -15128
rect 7650 -15234 7656 -15174
rect 7716 -15234 7722 -15174
rect 6936 -15392 7424 -15386
rect 6936 -15426 6948 -15392
rect 7412 -15426 7424 -15392
rect 6936 -15432 7424 -15426
rect 4604 -15514 4618 -15476
rect 3634 -16052 3640 -15522
rect 4612 -15994 4618 -15514
rect 3594 -16064 3640 -16052
rect 4598 -16052 4618 -15994
rect 4652 -15514 4664 -15476
rect 4652 -16052 4658 -15514
rect 5624 -15528 5636 -15476
rect 5630 -16032 5636 -15528
rect 2864 -16102 3352 -16096
rect 2864 -16136 2876 -16102
rect 3340 -16136 3352 -16102
rect 2864 -16142 3352 -16136
rect 3882 -16102 4370 -16096
rect 3882 -16136 3894 -16102
rect 4358 -16136 4370 -16102
rect 3882 -16142 4370 -16136
rect 2436 -16230 2442 -16170
rect 2502 -16230 2508 -16170
rect 4598 -16274 4658 -16052
rect 5620 -16052 5636 -16032
rect 5670 -15528 5684 -15476
rect 5670 -16032 5676 -15528
rect 6642 -15540 6654 -15476
rect 6648 -15988 6654 -15540
rect 5670 -16052 5680 -16032
rect 4900 -16102 5388 -16096
rect 4900 -16136 4912 -16102
rect 5376 -16136 5388 -16102
rect 4900 -16142 5388 -16136
rect 2560 -16334 2566 -16274
rect 2626 -16334 2632 -16274
rect 4080 -16334 4086 -16274
rect 4146 -16334 4152 -16274
rect 4592 -16334 4598 -16274
rect 4658 -16334 4664 -16274
rect 2330 -16456 2336 -16396
rect 2396 -16456 2402 -16396
rect 2218 -16570 2224 -16510
rect 2284 -16570 2290 -16510
rect 2336 -17638 2396 -16456
rect 2566 -16710 2626 -16334
rect 3066 -16570 3072 -16510
rect 3132 -16570 3138 -16510
rect 3072 -16620 3132 -16570
rect 4086 -16620 4146 -16334
rect 4598 -16568 4604 -16508
rect 4664 -16568 4670 -16508
rect 2862 -16626 3350 -16620
rect 2862 -16660 2874 -16626
rect 3338 -16660 3350 -16626
rect 2862 -16666 3350 -16660
rect 3880 -16626 4368 -16620
rect 3880 -16660 3892 -16626
rect 4356 -16660 4368 -16626
rect 3880 -16666 4368 -16660
rect 3592 -16710 3638 -16698
rect 4604 -16710 4664 -16568
rect 5102 -16620 5162 -16142
rect 5620 -16170 5680 -16052
rect 6634 -16052 6654 -15988
rect 6688 -15510 6704 -15476
rect 7656 -15476 7716 -15234
rect 8164 -15386 8224 -15128
rect 7954 -15392 8442 -15386
rect 7954 -15426 7966 -15392
rect 8430 -15426 8442 -15392
rect 7954 -15432 8442 -15426
rect 8676 -15476 8736 -15018
rect 9190 -15068 9250 -14910
rect 9696 -15028 9756 -14820
rect 10708 -14820 10726 -14744
rect 10760 -14312 10770 -14244
rect 11738 -14244 11784 -14232
rect 10760 -14744 10766 -14312
rect 10760 -14820 10768 -14744
rect 11738 -14758 11744 -14244
rect 11732 -14760 11744 -14758
rect 9990 -14870 10478 -14864
rect 9990 -14904 10002 -14870
rect 10466 -14904 10478 -14870
rect 9990 -14910 10478 -14904
rect 9184 -15128 9190 -15068
rect 9250 -15128 9256 -15068
rect 9696 -15088 9922 -15028
rect 10210 -15068 10270 -14910
rect 10708 -14958 10768 -14820
rect 11730 -14820 11744 -14760
rect 11778 -14758 11784 -14244
rect 12750 -14244 12810 -13854
rect 13252 -13920 13312 -13914
rect 13252 -14154 13312 -13980
rect 14260 -13920 14320 -13914
rect 14320 -13980 14322 -13974
rect 14260 -13986 14322 -13980
rect 14262 -14154 14322 -13986
rect 13044 -14160 13532 -14154
rect 13044 -14194 13056 -14160
rect 13520 -14194 13532 -14160
rect 13044 -14200 13532 -14194
rect 14062 -14160 14550 -14154
rect 14062 -14194 14074 -14160
rect 14538 -14194 14550 -14160
rect 14062 -14200 14550 -14194
rect 13774 -14244 13820 -14232
rect 14782 -14244 14842 -13854
rect 15276 -13920 15336 -13914
rect 16300 -13920 16360 -13914
rect 15336 -13980 15338 -13974
rect 15276 -13986 15338 -13980
rect 15278 -14154 15338 -13986
rect 16300 -14154 16360 -13980
rect 15080 -14160 15568 -14154
rect 15080 -14194 15092 -14160
rect 15556 -14194 15568 -14160
rect 15080 -14200 15568 -14194
rect 16098 -14160 16586 -14154
rect 16098 -14194 16110 -14160
rect 16574 -14194 16586 -14160
rect 16098 -14200 16586 -14194
rect 15810 -14244 15856 -14232
rect 16822 -14244 16882 -13854
rect 17322 -13920 17382 -13914
rect 18344 -13920 18404 -13914
rect 17322 -14154 17382 -13980
rect 18342 -13980 18344 -13974
rect 18342 -13986 18404 -13980
rect 17838 -14096 17844 -14036
rect 17904 -14096 17910 -14036
rect 17116 -14160 17604 -14154
rect 17116 -14194 17128 -14160
rect 17592 -14194 17604 -14160
rect 17116 -14200 17604 -14194
rect 12750 -14312 12762 -14244
rect 12756 -14754 12762 -14312
rect 11778 -14820 11792 -14758
rect 12744 -14820 12762 -14754
rect 12796 -14312 12810 -14244
rect 13764 -14278 13780 -14244
rect 12796 -14754 12802 -14312
rect 12796 -14820 12804 -14754
rect 13774 -14772 13780 -14278
rect 11008 -14870 11496 -14864
rect 11008 -14904 11020 -14870
rect 11484 -14904 11496 -14870
rect 11008 -14910 11496 -14904
rect 10702 -15018 10708 -14958
rect 10768 -15018 10774 -14958
rect 9190 -15386 9250 -15128
rect 9690 -15234 9696 -15174
rect 9756 -15234 9762 -15174
rect 8972 -15392 9460 -15386
rect 8972 -15426 8984 -15392
rect 9448 -15426 9460 -15392
rect 8972 -15432 9460 -15426
rect 9696 -15476 9756 -15234
rect 9862 -15280 9922 -15088
rect 10204 -15128 10210 -15068
rect 10270 -15128 10276 -15068
rect 9856 -15340 9862 -15280
rect 9922 -15340 9928 -15280
rect 10210 -15386 10270 -15128
rect 9990 -15392 10478 -15386
rect 9990 -15426 10002 -15392
rect 10466 -15426 10478 -15392
rect 9990 -15432 10478 -15426
rect 6688 -15540 6702 -15510
rect 7656 -15520 7672 -15476
rect 6688 -16052 6694 -15540
rect 5918 -16102 6406 -16096
rect 5918 -16136 5930 -16102
rect 6394 -16136 6406 -16102
rect 5918 -16142 6406 -16136
rect 5614 -16230 5620 -16170
rect 5680 -16230 5686 -16170
rect 5616 -16334 5622 -16274
rect 5682 -16334 5688 -16274
rect 4898 -16626 5386 -16620
rect 4898 -16660 4910 -16626
rect 5374 -16660 5386 -16626
rect 4898 -16666 5386 -16660
rect 2566 -16766 2580 -16710
rect 2574 -17286 2580 -16766
rect 2614 -16766 2626 -16710
rect 3586 -16742 3598 -16710
rect 2614 -17286 2620 -16766
rect 3592 -17242 3598 -16742
rect 2574 -17298 2620 -17286
rect 3586 -17286 3598 -17242
rect 3632 -16742 3646 -16710
rect 4604 -16736 4616 -16710
rect 3632 -17242 3638 -16742
rect 3632 -17286 3646 -17242
rect 2862 -17336 3350 -17330
rect 2862 -17370 2874 -17336
rect 3338 -17370 3350 -17336
rect 2862 -17376 3350 -17370
rect 3586 -17438 3646 -17286
rect 4610 -17286 4616 -16736
rect 4650 -16736 4664 -16710
rect 5622 -16710 5682 -16334
rect 6122 -16620 6182 -16142
rect 6634 -16274 6694 -16052
rect 7666 -16052 7672 -15520
rect 7706 -15510 7718 -15476
rect 7706 -15520 7716 -15510
rect 8676 -15518 8690 -15476
rect 7706 -16052 7712 -15520
rect 8684 -16010 8690 -15518
rect 8676 -16052 8690 -16010
rect 8724 -15518 8736 -15476
rect 8724 -16010 8730 -15518
rect 9692 -15538 9708 -15476
rect 8724 -16052 8736 -16010
rect 9702 -16052 9708 -15538
rect 9742 -15516 9756 -15476
rect 10708 -15476 10768 -15018
rect 11230 -15068 11290 -14910
rect 11224 -15128 11230 -15068
rect 11290 -15128 11296 -15068
rect 11230 -15386 11290 -15128
rect 11730 -15174 11790 -14820
rect 12026 -14870 12514 -14864
rect 12026 -14904 12038 -14870
rect 12502 -14904 12514 -14870
rect 12026 -14910 12514 -14904
rect 12232 -15068 12292 -14910
rect 12744 -14958 12804 -14820
rect 13766 -14820 13780 -14772
rect 13814 -14278 13824 -14244
rect 13814 -14772 13820 -14278
rect 14782 -14298 14798 -14244
rect 14792 -14760 14798 -14298
rect 13814 -14820 13826 -14772
rect 13044 -14870 13532 -14864
rect 13044 -14904 13056 -14870
rect 13520 -14904 13532 -14870
rect 13044 -14910 13532 -14904
rect 12738 -15018 12744 -14958
rect 12804 -15018 12810 -14958
rect 12226 -15128 12232 -15068
rect 12292 -15128 12298 -15068
rect 11724 -15234 11730 -15174
rect 11790 -15234 11796 -15174
rect 11724 -15340 11730 -15280
rect 11790 -15340 11796 -15280
rect 11008 -15392 11496 -15386
rect 11008 -15426 11020 -15392
rect 11484 -15426 11496 -15392
rect 11008 -15432 11496 -15426
rect 11730 -15476 11790 -15340
rect 12232 -15386 12292 -15128
rect 12026 -15392 12514 -15386
rect 12026 -15426 12038 -15392
rect 12502 -15426 12514 -15392
rect 12026 -15432 12514 -15426
rect 12744 -15476 12804 -15018
rect 13258 -15068 13318 -14910
rect 13252 -15128 13258 -15068
rect 13318 -15128 13324 -15068
rect 13258 -15386 13318 -15128
rect 13766 -15174 13826 -14820
rect 14780 -14820 14798 -14760
rect 14832 -14298 14842 -14244
rect 15802 -14284 15816 -14244
rect 14832 -14760 14838 -14298
rect 15810 -14754 15816 -14284
rect 14832 -14820 14840 -14760
rect 15806 -14780 15816 -14754
rect 14062 -14870 14550 -14864
rect 14062 -14904 14074 -14870
rect 14538 -14904 14550 -14870
rect 14062 -14910 14550 -14904
rect 14276 -15068 14336 -14910
rect 14780 -14958 14840 -14820
rect 15804 -14820 15816 -14780
rect 15850 -14284 15862 -14244
rect 15850 -14754 15856 -14284
rect 16822 -14298 16834 -14244
rect 15850 -14820 15866 -14754
rect 16828 -14770 16834 -14298
rect 16818 -14820 16834 -14770
rect 16868 -14298 16882 -14244
rect 17844 -14244 17904 -14096
rect 18342 -14154 18402 -13986
rect 18134 -14160 18622 -14154
rect 18134 -14194 18146 -14160
rect 18610 -14194 18622 -14160
rect 18134 -14200 18622 -14194
rect 16868 -14770 16874 -14298
rect 17844 -14308 17852 -14244
rect 17846 -14764 17852 -14308
rect 16868 -14820 16878 -14770
rect 17838 -14820 17852 -14764
rect 17886 -14308 17904 -14244
rect 18858 -14244 18918 -13854
rect 19362 -13920 19422 -13914
rect 20376 -13920 20436 -13914
rect 19422 -13980 19424 -13974
rect 19362 -13986 19424 -13980
rect 20436 -13980 20438 -13974
rect 20376 -13986 20438 -13980
rect 19364 -14154 19424 -13986
rect 20378 -14154 20438 -13986
rect 19152 -14160 19640 -14154
rect 19152 -14194 19164 -14160
rect 19628 -14194 19640 -14160
rect 19152 -14200 19640 -14194
rect 20170 -14160 20658 -14154
rect 20170 -14194 20182 -14160
rect 20646 -14194 20658 -14160
rect 20170 -14200 20658 -14194
rect 19882 -14244 19928 -14232
rect 20892 -14244 20952 -13854
rect 21400 -13920 21460 -13914
rect 21398 -13980 21400 -13974
rect 21398 -13986 21460 -13980
rect 21398 -14154 21458 -13986
rect 21910 -14096 21916 -14036
rect 21976 -14096 21982 -14036
rect 23042 -14096 23048 -14036
rect 23108 -14096 23114 -14036
rect 21188 -14160 21676 -14154
rect 21188 -14194 21200 -14160
rect 21664 -14194 21676 -14160
rect 21188 -14200 21676 -14194
rect 21916 -14244 21976 -14096
rect 22206 -14160 22694 -14154
rect 22206 -14194 22218 -14160
rect 22682 -14194 22694 -14160
rect 22206 -14200 22694 -14194
rect 18858 -14304 18870 -14244
rect 17886 -14764 17892 -14308
rect 17886 -14766 17898 -14764
rect 17886 -14820 17900 -14766
rect 18864 -14784 18870 -14304
rect 18856 -14820 18870 -14784
rect 18904 -14304 18918 -14244
rect 19874 -14284 19888 -14244
rect 18904 -14784 18910 -14304
rect 19882 -14764 19888 -14284
rect 18904 -14820 18916 -14784
rect 15080 -14870 15568 -14864
rect 15080 -14904 15092 -14870
rect 15556 -14904 15568 -14870
rect 15080 -14910 15568 -14904
rect 14774 -15018 14780 -14958
rect 14840 -15018 14846 -14958
rect 14270 -15128 14276 -15068
rect 14336 -15128 14342 -15068
rect 13760 -15234 13766 -15174
rect 13826 -15234 13832 -15174
rect 13762 -15340 13768 -15280
rect 13828 -15340 13834 -15280
rect 13044 -15392 13532 -15386
rect 13044 -15426 13056 -15392
rect 13520 -15426 13532 -15392
rect 13044 -15432 13532 -15426
rect 13768 -15476 13828 -15340
rect 14276 -15386 14336 -15128
rect 14062 -15392 14550 -15386
rect 14062 -15426 14074 -15392
rect 14538 -15426 14550 -15392
rect 14062 -15432 14550 -15426
rect 14780 -15476 14840 -15018
rect 15284 -15068 15344 -14910
rect 15804 -15036 15864 -14820
rect 16296 -14864 16356 -14862
rect 16098 -14870 16586 -14864
rect 16098 -14904 16110 -14870
rect 16574 -14904 16586 -14870
rect 16098 -14910 16586 -14904
rect 15278 -15128 15284 -15068
rect 15344 -15128 15350 -15068
rect 15648 -15096 15864 -15036
rect 16296 -15068 16356 -14910
rect 16818 -14958 16878 -14820
rect 17846 -14832 17892 -14820
rect 17328 -14864 17388 -14862
rect 17116 -14870 17604 -14864
rect 17116 -14904 17128 -14870
rect 17592 -14904 17604 -14870
rect 17116 -14910 17604 -14904
rect 18134 -14870 18622 -14864
rect 18134 -14904 18146 -14870
rect 18610 -14904 18622 -14870
rect 18134 -14910 18622 -14904
rect 16812 -15018 16818 -14958
rect 16878 -15018 16884 -14958
rect 15284 -15386 15344 -15128
rect 15648 -15280 15708 -15096
rect 16290 -15128 16296 -15068
rect 16356 -15128 16362 -15068
rect 15796 -15234 15802 -15174
rect 15862 -15234 15868 -15174
rect 15642 -15340 15648 -15280
rect 15708 -15340 15714 -15280
rect 15080 -15392 15568 -15386
rect 15080 -15426 15092 -15392
rect 15556 -15426 15568 -15392
rect 15080 -15432 15568 -15426
rect 9742 -15538 9752 -15516
rect 10708 -15532 10726 -15476
rect 9742 -16052 9748 -15538
rect 10720 -16010 10726 -15532
rect 7666 -16064 7712 -16052
rect 8684 -16064 8730 -16052
rect 9702 -16064 9748 -16052
rect 10712 -16052 10726 -16010
rect 10760 -15532 10768 -15476
rect 11728 -15528 11744 -15476
rect 10760 -16010 10766 -15532
rect 10760 -16052 10772 -16010
rect 6936 -16102 7424 -16096
rect 6936 -16136 6948 -16102
rect 7412 -16136 7424 -16102
rect 6936 -16142 7424 -16136
rect 7954 -16102 8442 -16096
rect 7954 -16136 7966 -16102
rect 8430 -16136 8442 -16102
rect 7954 -16142 8442 -16136
rect 8972 -16102 9460 -16096
rect 8972 -16136 8984 -16102
rect 9448 -16136 9460 -16102
rect 8972 -16142 9460 -16136
rect 9990 -16102 10478 -16096
rect 9990 -16136 10002 -16102
rect 10466 -16136 10478 -16102
rect 9990 -16142 10478 -16136
rect 6628 -16334 6634 -16274
rect 6694 -16334 6700 -16274
rect 6634 -16568 6640 -16508
rect 6700 -16568 6706 -16508
rect 5916 -16626 6404 -16620
rect 5916 -16660 5928 -16626
rect 6392 -16660 6404 -16626
rect 5916 -16666 6404 -16660
rect 4650 -17286 4656 -16736
rect 5622 -16742 5634 -16710
rect 5628 -17246 5634 -16742
rect 4610 -17298 4656 -17286
rect 5620 -17286 5634 -17246
rect 5668 -16742 5682 -16710
rect 6640 -16710 6700 -16568
rect 7134 -16620 7194 -16142
rect 7648 -16334 7654 -16274
rect 7714 -16334 7720 -16274
rect 6934 -16626 7422 -16620
rect 6934 -16660 6946 -16626
rect 7410 -16660 7422 -16626
rect 6934 -16666 7422 -16660
rect 6640 -16740 6652 -16710
rect 5668 -17246 5674 -16742
rect 5668 -17286 5680 -17246
rect 3880 -17336 4368 -17330
rect 3880 -17370 3892 -17336
rect 4356 -17370 4368 -17336
rect 3880 -17376 4368 -17370
rect 4898 -17336 5386 -17330
rect 4898 -17370 4910 -17336
rect 5374 -17370 5386 -17336
rect 4898 -17376 5386 -17370
rect 2442 -17498 2448 -17438
rect 2508 -17498 2514 -17438
rect 3580 -17498 3586 -17438
rect 3646 -17498 3652 -17438
rect 2330 -17698 2336 -17638
rect 2396 -17698 2402 -17638
rect 2224 -17800 2230 -17740
rect 2290 -17800 2296 -17740
rect 2114 -21252 2120 -21192
rect 2180 -21252 2186 -21192
rect 2230 -21230 2290 -17800
rect 2336 -18874 2396 -17698
rect 2330 -18934 2336 -18874
rect 2396 -18934 2402 -18874
rect 1882 -21402 1888 -21342
rect 1948 -21402 1954 -21342
rect 2120 -24928 2180 -21252
rect 2224 -21290 2230 -21230
rect 2290 -21290 2296 -21230
rect 2230 -23720 2290 -21290
rect 2336 -23594 2396 -18934
rect 2448 -20212 2508 -17498
rect 3578 -17698 3584 -17638
rect 3644 -17698 3650 -17638
rect 3584 -17742 3644 -17698
rect 2568 -17802 3644 -17742
rect 2568 -17804 3132 -17802
rect 2568 -17944 2628 -17804
rect 3072 -17854 3132 -17804
rect 2862 -17860 3350 -17854
rect 2862 -17894 2874 -17860
rect 3338 -17894 3350 -17860
rect 2862 -17900 3350 -17894
rect 2568 -17976 2580 -17944
rect 2574 -18520 2580 -17976
rect 2614 -17976 2628 -17944
rect 3584 -17944 3644 -17802
rect 4088 -17854 4148 -17376
rect 4596 -17578 4602 -17518
rect 4662 -17578 4668 -17518
rect 3880 -17860 4368 -17854
rect 3880 -17894 3892 -17860
rect 4356 -17894 4368 -17860
rect 3880 -17900 4368 -17894
rect 2614 -18520 2620 -17976
rect 3584 -17980 3598 -17944
rect 2574 -18532 2620 -18520
rect 3592 -18520 3598 -17980
rect 3632 -17980 3644 -17944
rect 4602 -17944 4662 -17578
rect 5116 -17632 5176 -17376
rect 5620 -17414 5680 -17286
rect 6646 -17286 6652 -16740
rect 6686 -16740 6700 -16710
rect 7654 -16710 7714 -16334
rect 8160 -16620 8220 -16142
rect 8670 -16230 8676 -16170
rect 8736 -16230 8742 -16170
rect 7952 -16626 8440 -16620
rect 7952 -16660 7964 -16626
rect 8428 -16660 8440 -16626
rect 7952 -16666 8440 -16660
rect 6686 -17286 6692 -16740
rect 7654 -16754 7670 -16710
rect 7664 -17236 7670 -16754
rect 6646 -17298 6692 -17286
rect 7656 -17286 7670 -17236
rect 7704 -16754 7714 -16710
rect 8676 -16710 8736 -16230
rect 10712 -16274 10772 -16052
rect 11738 -16052 11744 -15528
rect 11778 -15520 11792 -15476
rect 11778 -15528 11788 -15520
rect 12744 -15524 12762 -15476
rect 11778 -16052 11784 -15528
rect 12756 -16004 12762 -15524
rect 11738 -16064 11784 -16052
rect 12750 -16052 12762 -16004
rect 12796 -15524 12804 -15476
rect 13764 -15516 13780 -15476
rect 12796 -16004 12802 -15524
rect 12796 -16052 12810 -16004
rect 11008 -16102 11496 -16096
rect 11008 -16136 11020 -16102
rect 11484 -16136 11496 -16102
rect 11008 -16142 11496 -16136
rect 12026 -16102 12514 -16096
rect 12026 -16136 12038 -16102
rect 12502 -16136 12514 -16102
rect 12026 -16142 12514 -16136
rect 12750 -16274 12810 -16052
rect 13774 -16052 13780 -15516
rect 13814 -15514 13830 -15476
rect 13814 -15516 13828 -15514
rect 13814 -16052 13820 -15516
rect 14780 -15522 14798 -15476
rect 14792 -15998 14798 -15522
rect 14780 -16052 14798 -15998
rect 14832 -15522 14840 -15476
rect 15802 -15476 15862 -15234
rect 16296 -15386 16356 -15128
rect 16098 -15392 16586 -15386
rect 16098 -15426 16110 -15392
rect 16574 -15426 16586 -15392
rect 16098 -15432 16586 -15426
rect 16818 -15476 16878 -15018
rect 17328 -15068 17388 -14910
rect 18342 -15068 18402 -14910
rect 18856 -14958 18916 -14820
rect 19872 -14820 19888 -14764
rect 19922 -14284 19934 -14244
rect 19922 -14764 19928 -14284
rect 19922 -14820 19932 -14764
rect 19152 -14870 19640 -14864
rect 19152 -14904 19164 -14870
rect 19628 -14904 19640 -14870
rect 19152 -14910 19640 -14904
rect 18850 -15018 18856 -14958
rect 18916 -15018 18922 -14958
rect 17322 -15128 17328 -15068
rect 17388 -15128 17394 -15068
rect 18336 -15128 18342 -15068
rect 18402 -15128 18408 -15068
rect 17328 -15386 17388 -15128
rect 17836 -15234 17842 -15174
rect 17902 -15234 17908 -15174
rect 17116 -15392 17604 -15386
rect 17116 -15426 17128 -15392
rect 17592 -15426 17604 -15392
rect 17116 -15432 17604 -15426
rect 17842 -15476 17902 -15234
rect 18342 -15386 18402 -15128
rect 18134 -15392 18622 -15386
rect 18134 -15426 18146 -15392
rect 18610 -15426 18622 -15392
rect 18134 -15432 18622 -15426
rect 14832 -15998 14838 -15522
rect 15802 -15528 15816 -15476
rect 14832 -16052 14840 -15998
rect 15810 -16052 15816 -15528
rect 15850 -15518 15866 -15476
rect 15850 -15528 15862 -15518
rect 15850 -16052 15856 -15528
rect 13774 -16064 13820 -16052
rect 14792 -16064 14838 -16052
rect 15810 -16064 15856 -16052
rect 16818 -16052 16834 -15476
rect 16868 -16052 16878 -15476
rect 17838 -15518 17852 -15476
rect 17842 -15538 17852 -15518
rect 13044 -16102 13532 -16096
rect 13044 -16136 13056 -16102
rect 13520 -16136 13532 -16102
rect 13044 -16142 13532 -16136
rect 14062 -16102 14550 -16096
rect 14062 -16136 14074 -16102
rect 14538 -16136 14550 -16102
rect 14062 -16142 14550 -16136
rect 15080 -16102 15568 -16096
rect 15080 -16136 15092 -16102
rect 15556 -16136 15568 -16102
rect 15080 -16142 15568 -16136
rect 16098 -16102 16586 -16096
rect 16098 -16136 16110 -16102
rect 16574 -16136 16586 -16102
rect 16098 -16142 16586 -16136
rect 14776 -16230 14782 -16170
rect 14842 -16230 14848 -16170
rect 10706 -16334 10712 -16274
rect 10772 -16334 10778 -16274
rect 12744 -16334 12750 -16274
rect 12810 -16334 12816 -16274
rect 9690 -16456 9696 -16396
rect 9756 -16456 9762 -16396
rect 11724 -16456 11730 -16396
rect 11790 -16456 11796 -16396
rect 13754 -16456 13760 -16396
rect 13820 -16456 13826 -16396
rect 8970 -16626 9458 -16620
rect 8970 -16660 8982 -16626
rect 9446 -16660 9458 -16626
rect 8970 -16666 9458 -16660
rect 7704 -17236 7710 -16754
rect 8676 -16772 8688 -16710
rect 7704 -17286 7716 -17236
rect 8682 -17250 8688 -16772
rect 5916 -17336 6404 -17330
rect 5916 -17370 5928 -17336
rect 6392 -17370 6404 -17336
rect 5916 -17376 6404 -17370
rect 6934 -17336 7422 -17330
rect 6934 -17370 6946 -17336
rect 7410 -17370 7422 -17336
rect 6934 -17376 7422 -17370
rect 5614 -17474 5620 -17414
rect 5680 -17474 5686 -17414
rect 5110 -17692 5116 -17632
rect 5176 -17692 5182 -17632
rect 5116 -17854 5176 -17692
rect 4898 -17860 5386 -17854
rect 4898 -17894 4910 -17860
rect 5374 -17894 5386 -17860
rect 4898 -17900 5386 -17894
rect 3632 -18520 3638 -17980
rect 4602 -17986 4616 -17944
rect 4610 -18462 4616 -17986
rect 3592 -18532 3638 -18520
rect 4604 -18520 4616 -18462
rect 4650 -17986 4662 -17944
rect 5620 -17944 5680 -17474
rect 6118 -17626 6178 -17376
rect 6636 -17578 6642 -17518
rect 6702 -17578 6708 -17518
rect 6118 -17632 6180 -17626
rect 6118 -17692 6120 -17632
rect 6118 -17698 6180 -17692
rect 6118 -17854 6178 -17698
rect 5916 -17860 6404 -17854
rect 5916 -17894 5928 -17860
rect 6392 -17894 6404 -17860
rect 5916 -17900 6404 -17894
rect 4650 -18462 4656 -17986
rect 5620 -17988 5634 -17944
rect 4650 -18520 4664 -18462
rect 5628 -18472 5634 -17988
rect 2862 -18570 3350 -18564
rect 2862 -18604 2874 -18570
rect 3338 -18604 3350 -18570
rect 2862 -18610 3350 -18604
rect 3880 -18570 4368 -18564
rect 3880 -18604 3892 -18570
rect 4356 -18604 4368 -18570
rect 3880 -18610 4368 -18604
rect 3578 -18730 3584 -18670
rect 3644 -18730 3650 -18670
rect 2862 -19092 3350 -19086
rect 2862 -19126 2874 -19092
rect 3338 -19126 3350 -19092
rect 2862 -19132 3350 -19126
rect 2574 -19176 2620 -19164
rect 2574 -19706 2580 -19176
rect 2564 -19752 2580 -19706
rect 2614 -19706 2620 -19176
rect 3584 -19176 3644 -18730
rect 4090 -18772 4150 -18610
rect 4084 -18832 4090 -18772
rect 4150 -18832 4156 -18772
rect 4604 -18974 4664 -18520
rect 5622 -18520 5634 -18472
rect 5668 -17988 5680 -17944
rect 6642 -17944 6702 -17578
rect 7134 -17626 7194 -17376
rect 7656 -17414 7716 -17286
rect 8674 -17286 8688 -17250
rect 8722 -16772 8736 -16710
rect 9696 -16710 9756 -16456
rect 9988 -16626 10476 -16620
rect 9988 -16660 10000 -16626
rect 10464 -16660 10476 -16626
rect 9988 -16666 10476 -16660
rect 11006 -16626 11494 -16620
rect 11006 -16660 11018 -16626
rect 11482 -16660 11494 -16626
rect 11006 -16666 11494 -16660
rect 9696 -16766 9706 -16710
rect 8722 -17250 8728 -16772
rect 8722 -17286 8734 -17250
rect 7952 -17336 8440 -17330
rect 7952 -17370 7964 -17336
rect 8428 -17370 8440 -17336
rect 7952 -17376 8440 -17370
rect 7650 -17474 7656 -17414
rect 7716 -17474 7722 -17414
rect 7132 -17632 7194 -17626
rect 7192 -17692 7194 -17632
rect 7132 -17698 7194 -17692
rect 7134 -17854 7194 -17698
rect 6934 -17860 7422 -17854
rect 6934 -17894 6946 -17860
rect 7410 -17894 7422 -17860
rect 6934 -17900 7422 -17894
rect 6642 -17986 6652 -17944
rect 5668 -18472 5674 -17988
rect 5668 -18520 5682 -18472
rect 4898 -18570 5386 -18564
rect 4898 -18604 4910 -18570
rect 5374 -18604 5386 -18570
rect 4898 -18610 5386 -18604
rect 5622 -18670 5682 -18520
rect 6646 -18520 6652 -17986
rect 6686 -17986 6702 -17944
rect 7656 -17944 7716 -17474
rect 8152 -17632 8212 -17376
rect 8674 -17518 8734 -17286
rect 9700 -17286 9706 -16766
rect 9740 -16766 9756 -16710
rect 10718 -16710 10764 -16698
rect 9740 -17286 9746 -16766
rect 10718 -17256 10724 -16710
rect 9700 -17298 9746 -17286
rect 10708 -17286 10724 -17256
rect 10758 -17256 10764 -16710
rect 11730 -16710 11790 -16456
rect 12024 -16626 12512 -16620
rect 12024 -16660 12036 -16626
rect 12500 -16660 12512 -16626
rect 12024 -16666 12512 -16660
rect 13042 -16626 13530 -16620
rect 13042 -16660 13054 -16626
rect 13518 -16660 13530 -16626
rect 13042 -16666 13530 -16660
rect 11730 -16760 11742 -16710
rect 10758 -17286 10768 -17256
rect 8970 -17336 9458 -17330
rect 8970 -17370 8982 -17336
rect 9446 -17370 9458 -17336
rect 8970 -17376 9458 -17370
rect 9988 -17336 10476 -17330
rect 9988 -17370 10000 -17336
rect 10464 -17370 10476 -17336
rect 9988 -17376 10476 -17370
rect 8668 -17578 8674 -17518
rect 8734 -17578 8740 -17518
rect 9164 -17574 9224 -17376
rect 10206 -17574 10266 -17376
rect 10708 -17518 10768 -17286
rect 11736 -17286 11742 -16760
rect 11776 -16760 11790 -16710
rect 12754 -16710 12800 -16698
rect 11776 -17286 11782 -16760
rect 12754 -17244 12760 -16710
rect 11736 -17298 11782 -17286
rect 12748 -17286 12760 -17244
rect 12794 -17244 12800 -16710
rect 13760 -16710 13820 -16456
rect 14060 -16626 14548 -16620
rect 14060 -16660 14072 -16626
rect 14536 -16660 14548 -16626
rect 14060 -16666 14548 -16660
rect 13760 -16754 13778 -16710
rect 12794 -17286 12808 -17244
rect 11006 -17336 11494 -17330
rect 11006 -17370 11018 -17336
rect 11482 -17370 11494 -17336
rect 11006 -17376 11494 -17370
rect 12024 -17336 12512 -17330
rect 12024 -17370 12036 -17336
rect 12500 -17370 12512 -17336
rect 12024 -17376 12512 -17370
rect 8668 -17690 8674 -17630
rect 8734 -17690 8740 -17630
rect 9164 -17634 10266 -17574
rect 10702 -17578 10708 -17518
rect 10768 -17578 10774 -17518
rect 8152 -17854 8212 -17692
rect 7952 -17860 8440 -17854
rect 7952 -17894 7964 -17860
rect 8428 -17894 8440 -17860
rect 7952 -17900 8440 -17894
rect 6686 -18520 6692 -17986
rect 7656 -17992 7670 -17944
rect 7664 -18470 7670 -17992
rect 6646 -18532 6692 -18520
rect 7658 -18520 7670 -18470
rect 7704 -17992 7716 -17944
rect 8674 -17944 8734 -17690
rect 9164 -17854 9224 -17634
rect 9686 -17800 9692 -17740
rect 9752 -17800 9758 -17740
rect 8970 -17860 9458 -17854
rect 8970 -17894 8982 -17860
rect 9446 -17894 9458 -17860
rect 8970 -17900 9458 -17894
rect 7704 -18470 7710 -17992
rect 8674 -18002 8688 -17944
rect 7704 -18520 7718 -18470
rect 5916 -18570 6404 -18564
rect 5916 -18604 5928 -18570
rect 6392 -18604 6404 -18570
rect 5916 -18610 6404 -18604
rect 6934 -18570 7422 -18564
rect 6934 -18604 6946 -18570
rect 7410 -18604 7422 -18570
rect 6934 -18610 7422 -18604
rect 5616 -18730 5622 -18670
rect 5682 -18730 5688 -18670
rect 5614 -18934 5620 -18874
rect 5680 -18934 5686 -18874
rect 6128 -18880 6188 -18610
rect 7150 -18880 7210 -18610
rect 7658 -18670 7718 -18520
rect 8682 -18520 8688 -18002
rect 8722 -18002 8734 -17944
rect 9692 -17944 9752 -17800
rect 10206 -17854 10266 -17634
rect 10704 -17690 10710 -17630
rect 10770 -17690 10776 -17630
rect 9988 -17860 10476 -17854
rect 9988 -17894 10000 -17860
rect 10464 -17894 10476 -17860
rect 9988 -17900 10476 -17894
rect 9692 -17990 9706 -17944
rect 8722 -18520 8728 -18002
rect 8682 -18532 8728 -18520
rect 9700 -18520 9706 -17990
rect 9740 -17990 9752 -17944
rect 10710 -17944 10770 -17690
rect 11206 -17854 11266 -17376
rect 11720 -17800 11726 -17740
rect 11786 -17800 11792 -17740
rect 11006 -17860 11494 -17854
rect 11006 -17894 11018 -17860
rect 11482 -17894 11494 -17860
rect 11006 -17900 11494 -17894
rect 9740 -18520 9746 -17990
rect 10710 -18012 10724 -17944
rect 9700 -18532 9746 -18520
rect 10718 -18520 10724 -18012
rect 10758 -18012 10770 -17944
rect 11726 -17944 11786 -17800
rect 12240 -17854 12300 -17376
rect 12748 -17518 12808 -17286
rect 13772 -17286 13778 -16754
rect 13812 -16754 13820 -16710
rect 14782 -16710 14842 -16230
rect 15304 -16620 15364 -16142
rect 15794 -16334 15800 -16274
rect 15860 -16334 15866 -16274
rect 15078 -16626 15566 -16620
rect 15078 -16660 15090 -16626
rect 15554 -16660 15566 -16626
rect 15078 -16666 15566 -16660
rect 13812 -17286 13818 -16754
rect 14782 -16762 14796 -16710
rect 14790 -17234 14796 -16762
rect 13772 -17298 13818 -17286
rect 14782 -17286 14796 -17234
rect 14830 -16762 14842 -16710
rect 15800 -16710 15860 -16334
rect 16306 -16620 16366 -16142
rect 16818 -16274 16878 -16052
rect 17846 -16052 17852 -15538
rect 17886 -15538 17902 -15476
rect 18856 -15476 18916 -15018
rect 19360 -15068 19420 -14910
rect 19354 -15128 19360 -15068
rect 19420 -15128 19426 -15068
rect 19360 -15386 19420 -15128
rect 19872 -15174 19932 -14820
rect 20892 -14820 20906 -14244
rect 20940 -14276 20954 -14244
rect 21912 -14272 21924 -14244
rect 20940 -14820 20952 -14276
rect 21916 -14308 21924 -14272
rect 21918 -14760 21924 -14308
rect 20170 -14870 20658 -14864
rect 20170 -14904 20182 -14870
rect 20646 -14904 20658 -14870
rect 20170 -14910 20658 -14904
rect 20384 -15068 20444 -14910
rect 20892 -14958 20952 -14820
rect 21912 -14820 21924 -14760
rect 21958 -14308 21976 -14244
rect 22936 -14244 22982 -14232
rect 21958 -14760 21964 -14308
rect 21958 -14820 21972 -14760
rect 22936 -14772 22942 -14244
rect 21188 -14870 21676 -14864
rect 21188 -14904 21200 -14870
rect 21664 -14904 21676 -14870
rect 21188 -14910 21676 -14904
rect 20886 -15018 20892 -14958
rect 20952 -15018 20958 -14958
rect 20378 -15128 20384 -15068
rect 20444 -15128 20450 -15068
rect 19866 -15234 19872 -15174
rect 19932 -15234 19938 -15174
rect 19866 -15338 19872 -15278
rect 19932 -15338 19938 -15278
rect 19152 -15392 19640 -15386
rect 19152 -15426 19164 -15392
rect 19628 -15426 19640 -15392
rect 19152 -15432 19640 -15426
rect 19352 -15444 19412 -15432
rect 19872 -15476 19932 -15338
rect 20384 -15386 20444 -15128
rect 20170 -15392 20658 -15386
rect 20170 -15426 20182 -15392
rect 20646 -15426 20658 -15392
rect 20170 -15432 20658 -15426
rect 18856 -15534 18870 -15476
rect 17886 -16052 17892 -15538
rect 18864 -16004 18870 -15534
rect 17846 -16064 17892 -16052
rect 18854 -16052 18870 -16004
rect 18904 -15534 18916 -15476
rect 19870 -15522 19888 -15476
rect 18904 -16004 18910 -15534
rect 19872 -15550 19888 -15522
rect 19882 -15998 19888 -15550
rect 18904 -16052 18914 -16004
rect 17116 -16102 17604 -16096
rect 17116 -16136 17128 -16102
rect 17592 -16136 17604 -16102
rect 17116 -16142 17604 -16136
rect 18134 -16102 18622 -16096
rect 18134 -16136 18146 -16102
rect 18610 -16136 18622 -16102
rect 18134 -16142 18622 -16136
rect 16812 -16334 16818 -16274
rect 16878 -16334 16884 -16274
rect 17318 -16620 17378 -16142
rect 17832 -16334 17838 -16274
rect 17898 -16334 17904 -16274
rect 16096 -16626 16584 -16620
rect 16096 -16660 16108 -16626
rect 16572 -16660 16584 -16626
rect 16096 -16666 16584 -16660
rect 17114 -16626 17602 -16620
rect 17114 -16660 17126 -16626
rect 17590 -16660 17602 -16626
rect 17114 -16666 17602 -16660
rect 15800 -16758 15814 -16710
rect 14830 -17234 14836 -16762
rect 14830 -17286 14842 -17234
rect 15808 -17254 15814 -16758
rect 13042 -17336 13530 -17330
rect 13042 -17370 13054 -17336
rect 13518 -17370 13530 -17336
rect 13042 -17376 13530 -17370
rect 14060 -17336 14548 -17330
rect 14060 -17370 14072 -17336
rect 14536 -17370 14548 -17336
rect 14060 -17376 14548 -17370
rect 12742 -17578 12748 -17518
rect 12808 -17578 12814 -17518
rect 13262 -17574 13322 -17376
rect 14270 -17574 14330 -17376
rect 14782 -17518 14842 -17286
rect 15800 -17286 15814 -17254
rect 15848 -16758 15860 -16710
rect 16826 -16710 16872 -16698
rect 15848 -17254 15854 -16758
rect 16826 -17250 16832 -16710
rect 15848 -17286 15860 -17254
rect 15078 -17336 15566 -17330
rect 15078 -17370 15090 -17336
rect 15554 -17370 15566 -17336
rect 15078 -17376 15566 -17370
rect 12740 -17690 12746 -17630
rect 12806 -17690 12812 -17630
rect 13262 -17634 14330 -17574
rect 14776 -17578 14782 -17518
rect 14842 -17578 14848 -17518
rect 14972 -17582 14978 -17522
rect 15038 -17582 15044 -17522
rect 12024 -17860 12512 -17854
rect 12024 -17894 12036 -17860
rect 12500 -17894 12512 -17860
rect 12024 -17900 12512 -17894
rect 11726 -17992 11742 -17944
rect 10758 -18520 10764 -18012
rect 10718 -18532 10764 -18520
rect 11736 -18520 11742 -17992
rect 11776 -17992 11786 -17944
rect 12746 -17944 12806 -17690
rect 13262 -17854 13322 -17634
rect 13760 -17800 13766 -17740
rect 13826 -17800 13832 -17740
rect 13042 -17860 13530 -17854
rect 13042 -17894 13054 -17860
rect 13518 -17894 13530 -17860
rect 13042 -17900 13530 -17894
rect 11776 -18520 11782 -17992
rect 12746 -17994 12760 -17944
rect 11736 -18532 11782 -18520
rect 12754 -18520 12760 -17994
rect 12794 -17994 12806 -17944
rect 13766 -17944 13826 -17800
rect 14270 -17854 14330 -17634
rect 14776 -17690 14782 -17630
rect 14842 -17690 14848 -17630
rect 14060 -17860 14548 -17854
rect 14060 -17894 14072 -17860
rect 14536 -17894 14548 -17860
rect 14060 -17900 14548 -17894
rect 13766 -17982 13778 -17944
rect 12794 -18520 12800 -17994
rect 13772 -18474 13778 -17982
rect 12754 -18532 12800 -18520
rect 13766 -18520 13778 -18474
rect 13812 -17982 13826 -17944
rect 14782 -17944 14842 -17690
rect 14978 -17740 15038 -17582
rect 15272 -17738 15332 -17376
rect 15800 -17414 15860 -17286
rect 16816 -17286 16832 -17250
rect 16866 -17250 16872 -16710
rect 17838 -16710 17898 -16334
rect 18352 -16620 18412 -16142
rect 18854 -16274 18914 -16052
rect 19876 -16052 19888 -15998
rect 19922 -15550 19932 -15476
rect 20892 -15476 20952 -15018
rect 21404 -15068 21464 -14910
rect 21912 -14968 21972 -14820
rect 22928 -14820 22942 -14772
rect 22976 -14772 22982 -14244
rect 22976 -14820 22988 -14772
rect 22206 -14870 22694 -14864
rect 22206 -14904 22218 -14870
rect 22682 -14904 22694 -14870
rect 22206 -14910 22694 -14904
rect 22422 -14968 22482 -14910
rect 22928 -14968 22988 -14820
rect 23048 -14968 23108 -14096
rect 21912 -15028 23108 -14968
rect 21398 -15128 21404 -15068
rect 21464 -15128 21470 -15068
rect 21404 -15386 21464 -15128
rect 21906 -15234 21912 -15174
rect 21972 -15234 21978 -15174
rect 21912 -15276 21972 -15234
rect 21912 -15336 22990 -15276
rect 23048 -15278 23108 -15028
rect 21188 -15392 21676 -15386
rect 21188 -15426 21200 -15392
rect 21664 -15426 21676 -15392
rect 21188 -15432 21676 -15426
rect 20892 -15502 20906 -15476
rect 19922 -15998 19928 -15550
rect 20900 -15994 20906 -15502
rect 19922 -16052 19936 -15998
rect 19152 -16102 19640 -16096
rect 19152 -16136 19164 -16102
rect 19628 -16136 19640 -16102
rect 19152 -16142 19640 -16136
rect 19876 -16170 19936 -16052
rect 20890 -16052 20906 -15994
rect 20940 -15502 20952 -15476
rect 21912 -15476 21972 -15336
rect 22398 -15386 22458 -15336
rect 22206 -15392 22694 -15386
rect 22206 -15426 22218 -15392
rect 22682 -15426 22694 -15392
rect 22206 -15432 22694 -15426
rect 22930 -15476 22990 -15336
rect 23042 -15338 23048 -15278
rect 23108 -15338 23114 -15278
rect 20940 -15994 20946 -15502
rect 21912 -15532 21924 -15476
rect 20940 -16052 20950 -15994
rect 20170 -16102 20658 -16096
rect 20170 -16136 20182 -16102
rect 20646 -16136 20658 -16102
rect 20170 -16142 20658 -16136
rect 19870 -16230 19876 -16170
rect 19936 -16230 19942 -16170
rect 20890 -16274 20950 -16052
rect 21918 -16052 21924 -15532
rect 21958 -15532 21972 -15476
rect 22926 -15512 22942 -15476
rect 22930 -15518 22942 -15512
rect 21958 -16052 21964 -15532
rect 22936 -16008 22942 -15518
rect 21918 -16064 21964 -16052
rect 22932 -16052 22942 -16008
rect 22976 -15518 22990 -15476
rect 22976 -16008 22982 -15518
rect 22976 -16052 22992 -16008
rect 21188 -16102 21676 -16096
rect 21188 -16136 21200 -16102
rect 21664 -16136 21676 -16102
rect 21188 -16142 21676 -16136
rect 22206 -16102 22694 -16096
rect 22206 -16136 22218 -16102
rect 22682 -16136 22694 -16102
rect 22206 -16142 22694 -16136
rect 18848 -16334 18854 -16274
rect 18914 -16334 18920 -16274
rect 20884 -16334 20890 -16274
rect 20950 -16334 20956 -16274
rect 21380 -16620 21440 -16142
rect 22932 -16178 22992 -16052
rect 22932 -16238 23222 -16178
rect 22418 -16544 22986 -16484
rect 22418 -16620 22478 -16544
rect 18132 -16626 18620 -16620
rect 18132 -16660 18144 -16626
rect 18608 -16660 18620 -16626
rect 18132 -16666 18620 -16660
rect 19150 -16626 19638 -16620
rect 19150 -16660 19162 -16626
rect 19626 -16660 19638 -16626
rect 19150 -16666 19638 -16660
rect 20168 -16626 20656 -16620
rect 20168 -16660 20180 -16626
rect 20644 -16660 20656 -16626
rect 20168 -16666 20656 -16660
rect 21186 -16626 21674 -16620
rect 21186 -16660 21198 -16626
rect 21662 -16660 21674 -16626
rect 21186 -16666 21674 -16660
rect 22204 -16626 22692 -16620
rect 22204 -16660 22216 -16626
rect 22680 -16660 22692 -16626
rect 22204 -16666 22692 -16660
rect 17838 -16768 17850 -16710
rect 17844 -17240 17850 -16768
rect 16866 -17286 16876 -17250
rect 16096 -17336 16584 -17330
rect 16096 -17370 16108 -17336
rect 16572 -17370 16584 -17336
rect 16096 -17376 16584 -17370
rect 15794 -17474 15800 -17414
rect 15860 -17474 15866 -17414
rect 14972 -17800 14978 -17740
rect 15038 -17800 15044 -17740
rect 15266 -17798 15272 -17738
rect 15332 -17798 15338 -17738
rect 15272 -17854 15332 -17798
rect 15078 -17860 15566 -17854
rect 15078 -17894 15090 -17860
rect 15554 -17894 15566 -17860
rect 15078 -17900 15566 -17894
rect 13812 -18474 13818 -17982
rect 14782 -17988 14796 -17944
rect 13812 -18520 13826 -18474
rect 7952 -18570 8440 -18564
rect 7952 -18604 7964 -18570
rect 8428 -18604 8440 -18570
rect 7952 -18610 8440 -18604
rect 8970 -18570 9458 -18564
rect 8970 -18604 8982 -18570
rect 9446 -18604 9458 -18570
rect 8970 -18610 9458 -18604
rect 9988 -18570 10476 -18564
rect 9988 -18604 10000 -18570
rect 10464 -18604 10476 -18570
rect 9988 -18610 10476 -18604
rect 11006 -18570 11494 -18564
rect 11006 -18604 11018 -18570
rect 11482 -18604 11494 -18570
rect 11006 -18610 11494 -18604
rect 12024 -18570 12512 -18564
rect 12024 -18604 12036 -18570
rect 12500 -18604 12512 -18570
rect 12024 -18610 12512 -18604
rect 13042 -18570 13530 -18564
rect 13042 -18604 13054 -18570
rect 13518 -18604 13530 -18570
rect 13042 -18610 13530 -18604
rect 7652 -18730 7658 -18670
rect 7718 -18730 7724 -18670
rect 4598 -19034 4604 -18974
rect 4664 -19034 4670 -18974
rect 3880 -19092 4368 -19086
rect 3880 -19126 3892 -19092
rect 4356 -19126 4368 -19092
rect 3880 -19132 4368 -19126
rect 3584 -19214 3598 -19176
rect 2614 -19752 2624 -19706
rect 3592 -19710 3598 -19214
rect 2564 -19914 2624 -19752
rect 3582 -19752 3598 -19710
rect 3632 -19214 3644 -19176
rect 4604 -19176 4664 -19034
rect 4898 -19092 5386 -19086
rect 4898 -19126 4910 -19092
rect 5374 -19126 5386 -19092
rect 4898 -19132 5386 -19126
rect 3632 -19710 3638 -19214
rect 4604 -19216 4616 -19176
rect 3632 -19752 3642 -19710
rect 2862 -19802 3350 -19796
rect 2862 -19836 2874 -19802
rect 3338 -19836 3350 -19802
rect 2862 -19842 3350 -19836
rect 3076 -19914 3136 -19842
rect 3582 -19914 3642 -19752
rect 4610 -19752 4616 -19216
rect 4650 -19216 4664 -19176
rect 5620 -19176 5680 -18934
rect 6122 -18940 6128 -18880
rect 6188 -18940 6194 -18880
rect 7144 -18940 7150 -18880
rect 7210 -18940 7216 -18880
rect 6632 -19034 6638 -18974
rect 6698 -19034 6704 -18974
rect 5916 -19092 6404 -19086
rect 5916 -19126 5928 -19092
rect 6392 -19126 6404 -19092
rect 5916 -19132 6404 -19126
rect 4650 -19752 4656 -19216
rect 5620 -19228 5634 -19176
rect 4610 -19764 4656 -19752
rect 5628 -19752 5634 -19228
rect 5668 -19228 5680 -19176
rect 6638 -19176 6698 -19034
rect 7150 -19086 7210 -18940
rect 6934 -19092 7422 -19086
rect 6934 -19126 6946 -19092
rect 7410 -19126 7422 -19092
rect 6934 -19132 7422 -19126
rect 6638 -19220 6652 -19176
rect 5668 -19752 5674 -19228
rect 6646 -19716 6652 -19220
rect 5628 -19764 5674 -19752
rect 6638 -19752 6652 -19716
rect 6686 -19220 6698 -19176
rect 7658 -19176 7718 -18730
rect 8164 -18880 8224 -18610
rect 9182 -18772 9242 -18610
rect 10202 -18660 10262 -18610
rect 11202 -18660 11262 -18610
rect 12240 -18660 12300 -18610
rect 13268 -18660 13328 -18610
rect 9684 -18730 9690 -18670
rect 9750 -18730 9756 -18670
rect 10202 -18720 13328 -18660
rect 9176 -18832 9182 -18772
rect 9242 -18832 9248 -18772
rect 8158 -18940 8164 -18880
rect 8224 -18940 8230 -18880
rect 9176 -18940 9182 -18880
rect 9242 -18940 9248 -18880
rect 8164 -19086 8224 -18940
rect 8668 -19034 8674 -18974
rect 8734 -19034 8740 -18974
rect 7952 -19092 8440 -19086
rect 7952 -19126 7964 -19092
rect 8428 -19126 8440 -19092
rect 7952 -19132 8440 -19126
rect 6686 -19716 6692 -19220
rect 6686 -19752 6698 -19716
rect 3880 -19802 4368 -19796
rect 3880 -19836 3892 -19802
rect 4356 -19836 4368 -19802
rect 3880 -19842 4368 -19836
rect 4898 -19802 5386 -19796
rect 4898 -19836 4910 -19802
rect 5374 -19836 5386 -19802
rect 4898 -19842 5386 -19836
rect 5916 -19802 6404 -19796
rect 5916 -19836 5928 -19802
rect 6392 -19836 6404 -19802
rect 5916 -19842 6404 -19836
rect 4086 -19898 4146 -19842
rect 2564 -19974 3642 -19914
rect 4080 -19958 4086 -19898
rect 4146 -19958 4152 -19898
rect 4990 -19958 4996 -19898
rect 5056 -19958 5062 -19898
rect 4080 -20174 4086 -20114
rect 4146 -20174 4152 -20114
rect 4086 -20180 4148 -20174
rect 2448 -20218 2510 -20212
rect 2448 -20278 2450 -20218
rect 2448 -20284 2510 -20278
rect 2448 -22462 2508 -20284
rect 4088 -20320 4148 -20180
rect 4996 -20320 5056 -19958
rect 5124 -20114 5184 -19842
rect 5992 -19958 5998 -19898
rect 6058 -19958 6064 -19898
rect 5124 -20180 5184 -20174
rect 5998 -20320 6058 -19958
rect 6138 -20114 6198 -19842
rect 6638 -20000 6698 -19752
rect 7658 -19752 7670 -19176
rect 7704 -19752 7718 -19176
rect 8674 -19176 8734 -19034
rect 9182 -19086 9242 -18940
rect 8970 -19092 9458 -19086
rect 8970 -19126 8982 -19092
rect 9446 -19126 9458 -19092
rect 8970 -19132 9458 -19126
rect 8674 -19212 8688 -19176
rect 6934 -19802 7422 -19796
rect 6934 -19836 6946 -19802
rect 7410 -19836 7422 -19802
rect 6934 -19842 7422 -19836
rect 7150 -19898 7210 -19842
rect 7144 -19958 7150 -19898
rect 7210 -19958 7216 -19898
rect 6632 -20060 6638 -20000
rect 6698 -20060 6704 -20000
rect 6132 -20174 6138 -20114
rect 6198 -20174 6204 -20114
rect 7150 -20320 7210 -19958
rect 2862 -20326 3350 -20320
rect 2862 -20360 2874 -20326
rect 3338 -20360 3350 -20326
rect 2862 -20366 3350 -20360
rect 3880 -20326 4368 -20320
rect 3880 -20360 3892 -20326
rect 4356 -20360 4368 -20326
rect 3880 -20366 4368 -20360
rect 4898 -20326 5386 -20320
rect 4898 -20360 4910 -20326
rect 5374 -20360 5386 -20326
rect 4898 -20366 5386 -20360
rect 5916 -20326 6404 -20320
rect 5916 -20360 5928 -20326
rect 6392 -20360 6404 -20326
rect 5916 -20366 6404 -20360
rect 6934 -20326 7422 -20320
rect 6934 -20360 6946 -20326
rect 7410 -20360 7422 -20326
rect 6934 -20366 7422 -20360
rect 2574 -20410 2620 -20398
rect 2574 -20948 2580 -20410
rect 2568 -20986 2580 -20948
rect 2614 -20948 2620 -20410
rect 3592 -20410 3638 -20398
rect 3592 -20948 3598 -20410
rect 2614 -20986 2628 -20948
rect 2568 -21116 2628 -20986
rect 3586 -20986 3598 -20948
rect 3632 -20948 3638 -20410
rect 4610 -20410 4656 -20398
rect 4610 -20936 4616 -20410
rect 3632 -20986 3646 -20948
rect 2862 -21036 3350 -21030
rect 2862 -21070 2874 -21036
rect 3338 -21070 3350 -21036
rect 2862 -21076 3350 -21070
rect 3066 -21116 3126 -21076
rect 3586 -21116 3646 -20986
rect 4602 -20986 4616 -20936
rect 4650 -20936 4656 -20410
rect 5628 -20410 5674 -20398
rect 5628 -20928 5634 -20410
rect 4650 -20986 4662 -20936
rect 3880 -21036 4368 -21030
rect 3880 -21070 3892 -21036
rect 4356 -21070 4368 -21036
rect 3880 -21076 4368 -21070
rect 2568 -21176 3646 -21116
rect 3586 -21230 3646 -21176
rect 4078 -21186 4084 -21126
rect 4144 -21186 4150 -21126
rect 3580 -21290 3586 -21230
rect 3646 -21290 3652 -21230
rect 3576 -21500 3582 -21440
rect 3642 -21500 3648 -21440
rect 2862 -21560 3350 -21554
rect 2862 -21594 2874 -21560
rect 3338 -21594 3350 -21560
rect 2862 -21600 3350 -21594
rect 2574 -21644 2620 -21632
rect 2574 -22186 2580 -21644
rect 2564 -22220 2580 -22186
rect 2614 -22186 2620 -21644
rect 3582 -21644 3642 -21500
rect 4084 -21554 4144 -21186
rect 4602 -21342 4662 -20986
rect 5620 -20986 5634 -20928
rect 5668 -20928 5674 -20410
rect 6646 -20410 6692 -20398
rect 5668 -20986 5680 -20928
rect 6646 -20940 6652 -20410
rect 4898 -21036 5386 -21030
rect 4898 -21070 4910 -21036
rect 5374 -21070 5386 -21036
rect 4898 -21076 5386 -21070
rect 5092 -21126 5152 -21076
rect 5086 -21186 5092 -21126
rect 5152 -21186 5158 -21126
rect 4596 -21402 4602 -21342
rect 4662 -21402 4668 -21342
rect 5620 -21440 5680 -20986
rect 6640 -20986 6652 -20940
rect 6686 -20940 6692 -20410
rect 7658 -20410 7718 -19752
rect 8682 -19752 8688 -19212
rect 8722 -19212 8734 -19176
rect 9690 -19176 9750 -18730
rect 10196 -18940 10202 -18880
rect 10262 -18940 10268 -18880
rect 13268 -18896 13328 -18720
rect 13766 -18786 13826 -18520
rect 14790 -18520 14796 -17988
rect 14830 -17988 14842 -17944
rect 15800 -17944 15860 -17474
rect 16302 -17732 16362 -17376
rect 16816 -17630 16876 -17286
rect 17836 -17286 17850 -17240
rect 17884 -16768 17898 -16710
rect 18862 -16710 18908 -16698
rect 17884 -17240 17890 -16768
rect 18862 -17230 18868 -16710
rect 17884 -17286 17896 -17240
rect 17114 -17336 17602 -17330
rect 17114 -17370 17126 -17336
rect 17590 -17370 17602 -17336
rect 17114 -17376 17602 -17370
rect 16810 -17690 16816 -17630
rect 16876 -17690 16882 -17630
rect 16300 -17738 16362 -17732
rect 16360 -17798 16362 -17738
rect 16300 -17804 16362 -17798
rect 16812 -17804 16818 -17744
rect 16878 -17804 16884 -17744
rect 16302 -17854 16362 -17804
rect 16096 -17860 16584 -17854
rect 16096 -17894 16108 -17860
rect 16572 -17894 16584 -17860
rect 16096 -17900 16584 -17894
rect 15800 -17988 15814 -17944
rect 14830 -18520 14836 -17988
rect 14790 -18532 14836 -18520
rect 15808 -18520 15814 -17988
rect 15848 -17988 15860 -17944
rect 16818 -17944 16878 -17804
rect 17326 -17854 17386 -17376
rect 17836 -17414 17896 -17286
rect 18854 -17286 18868 -17230
rect 18902 -17230 18908 -16710
rect 19880 -16710 19926 -16698
rect 18902 -17286 18914 -17230
rect 19880 -17242 19886 -16710
rect 18132 -17336 18620 -17330
rect 18132 -17370 18144 -17336
rect 18608 -17370 18620 -17336
rect 18132 -17376 18620 -17370
rect 17830 -17474 17836 -17414
rect 17896 -17474 17902 -17414
rect 17114 -17860 17602 -17854
rect 17114 -17894 17126 -17860
rect 17590 -17894 17602 -17860
rect 17114 -17900 17602 -17894
rect 16818 -17974 16832 -17944
rect 15848 -18520 15854 -17988
rect 16826 -18480 16832 -17974
rect 15808 -18532 15854 -18520
rect 16818 -18520 16832 -18480
rect 16866 -17974 16878 -17944
rect 17836 -17944 17896 -17474
rect 18352 -17854 18412 -17376
rect 18854 -17630 18914 -17286
rect 19870 -17286 19886 -17242
rect 19920 -17242 19926 -16710
rect 20898 -16710 20944 -16698
rect 20898 -17242 20904 -16710
rect 19920 -17286 19930 -17242
rect 19150 -17336 19638 -17330
rect 19150 -17370 19162 -17336
rect 19626 -17370 19638 -17336
rect 19150 -17376 19638 -17370
rect 18848 -17690 18854 -17630
rect 18914 -17690 18920 -17630
rect 19360 -17680 19420 -17376
rect 19870 -17522 19930 -17286
rect 20894 -17286 20904 -17242
rect 20938 -17242 20944 -16710
rect 21916 -16710 21962 -16698
rect 21916 -17236 21922 -16710
rect 20938 -17286 20954 -17242
rect 20168 -17336 20656 -17330
rect 20168 -17370 20180 -17336
rect 20644 -17370 20656 -17336
rect 20168 -17376 20656 -17370
rect 20376 -17520 20436 -17376
rect 19864 -17582 19870 -17522
rect 19930 -17582 19936 -17522
rect 20374 -17526 20436 -17520
rect 20434 -17586 20436 -17526
rect 20374 -17592 20436 -17586
rect 20376 -17680 20436 -17592
rect 20894 -17630 20954 -17286
rect 21910 -17286 21922 -17236
rect 21956 -17236 21962 -16710
rect 22926 -16710 22986 -16544
rect 23028 -16568 23034 -16508
rect 23094 -16568 23100 -16508
rect 23162 -16526 23222 -16238
rect 22926 -16738 22940 -16710
rect 22934 -17228 22940 -16738
rect 21956 -17286 21970 -17236
rect 21186 -17336 21674 -17330
rect 21186 -17370 21198 -17336
rect 21662 -17370 21674 -17336
rect 21186 -17376 21674 -17370
rect 19360 -17740 20436 -17680
rect 20888 -17690 20894 -17630
rect 20954 -17690 20960 -17630
rect 18848 -17804 18854 -17744
rect 18914 -17804 18920 -17744
rect 18132 -17860 18620 -17854
rect 18132 -17894 18144 -17860
rect 18608 -17894 18620 -17860
rect 18132 -17900 18620 -17894
rect 16866 -18480 16872 -17974
rect 17836 -17984 17850 -17944
rect 16866 -18520 16878 -18480
rect 17844 -18486 17850 -17984
rect 14060 -18570 14548 -18564
rect 14060 -18604 14072 -18570
rect 14536 -18604 14548 -18570
rect 14060 -18610 14548 -18604
rect 15078 -18570 15566 -18564
rect 15078 -18604 15090 -18570
rect 15554 -18604 15566 -18570
rect 15078 -18610 15566 -18604
rect 16096 -18570 16584 -18564
rect 16096 -18604 16108 -18570
rect 16572 -18604 16584 -18570
rect 16096 -18610 16584 -18604
rect 14272 -18658 14332 -18610
rect 13760 -18846 13766 -18786
rect 13826 -18846 13832 -18786
rect 14272 -18896 14332 -18718
rect 10202 -19086 10262 -18940
rect 13268 -18956 14332 -18896
rect 15796 -19044 15802 -18984
rect 15862 -19044 15868 -18984
rect 9988 -19092 10476 -19086
rect 9988 -19126 10000 -19092
rect 10464 -19126 10476 -19092
rect 9988 -19132 10476 -19126
rect 11006 -19092 11494 -19086
rect 11006 -19126 11018 -19092
rect 11482 -19126 11494 -19092
rect 11006 -19132 11494 -19126
rect 12024 -19092 12512 -19086
rect 12024 -19126 12036 -19092
rect 12500 -19126 12512 -19092
rect 12024 -19132 12512 -19126
rect 13042 -19092 13530 -19086
rect 13042 -19126 13054 -19092
rect 13518 -19126 13530 -19092
rect 13042 -19132 13530 -19126
rect 14060 -19092 14548 -19086
rect 14060 -19126 14072 -19092
rect 14536 -19126 14548 -19092
rect 14060 -19132 14548 -19126
rect 15078 -19092 15566 -19086
rect 15078 -19126 15090 -19092
rect 15554 -19126 15566 -19092
rect 15078 -19132 15566 -19126
rect 8722 -19752 8728 -19212
rect 9690 -19214 9706 -19176
rect 8682 -19764 8728 -19752
rect 9700 -19752 9706 -19214
rect 9740 -19214 9750 -19176
rect 10718 -19176 10764 -19164
rect 9740 -19752 9746 -19214
rect 10718 -19710 10724 -19176
rect 9700 -19764 9746 -19752
rect 10710 -19752 10724 -19710
rect 10758 -19710 10764 -19176
rect 11736 -19176 11782 -19164
rect 10758 -19752 10770 -19710
rect 11736 -19714 11742 -19176
rect 7952 -19802 8440 -19796
rect 7952 -19836 7964 -19802
rect 8428 -19836 8440 -19802
rect 7952 -19842 8440 -19836
rect 8970 -19802 9458 -19796
rect 8970 -19836 8982 -19802
rect 9446 -19836 9458 -19802
rect 8970 -19842 9458 -19836
rect 9988 -19802 10476 -19796
rect 9988 -19836 10000 -19802
rect 10464 -19836 10476 -19802
rect 9988 -19842 10476 -19836
rect 8160 -19898 8220 -19842
rect 9166 -19898 9226 -19842
rect 10210 -19898 10270 -19842
rect 10710 -19892 10770 -19752
rect 11730 -19752 11742 -19714
rect 11776 -19714 11782 -19176
rect 12754 -19176 12800 -19164
rect 11776 -19752 11790 -19714
rect 12754 -19720 12760 -19176
rect 11006 -19802 11494 -19796
rect 11006 -19836 11018 -19802
rect 11482 -19836 11494 -19802
rect 11006 -19842 11494 -19836
rect 8154 -19958 8160 -19898
rect 8220 -19958 8226 -19898
rect 9160 -19958 9166 -19898
rect 9226 -19958 9232 -19898
rect 10204 -19958 10210 -19898
rect 10270 -19958 10276 -19898
rect 10704 -19952 10710 -19892
rect 10770 -19952 10776 -19892
rect 8160 -20320 8220 -19958
rect 9158 -20174 9164 -20114
rect 9224 -20174 9230 -20114
rect 10198 -20174 10204 -20114
rect 10264 -20174 10270 -20114
rect 9164 -20320 9224 -20174
rect 9682 -20278 9688 -20218
rect 9748 -20278 9754 -20218
rect 7952 -20326 8440 -20320
rect 7952 -20360 7964 -20326
rect 8428 -20360 8440 -20326
rect 7952 -20366 8440 -20360
rect 8970 -20326 9458 -20320
rect 8970 -20360 8982 -20326
rect 9446 -20360 9458 -20326
rect 8970 -20366 9458 -20360
rect 7658 -20492 7670 -20410
rect 7664 -20940 7670 -20492
rect 6686 -20986 6700 -20940
rect 5916 -21036 6404 -21030
rect 5916 -21070 5928 -21036
rect 6392 -21070 6404 -21036
rect 5916 -21076 6404 -21070
rect 6106 -21126 6166 -21076
rect 6100 -21186 6106 -21126
rect 6166 -21186 6172 -21126
rect 6640 -21342 6700 -20986
rect 7660 -20986 7670 -20940
rect 7704 -20492 7718 -20410
rect 8682 -20410 8728 -20398
rect 7704 -20940 7710 -20492
rect 7704 -20986 7720 -20940
rect 8682 -20942 8688 -20410
rect 6934 -21036 7422 -21030
rect 6934 -21070 6946 -21036
rect 7410 -21070 7422 -21036
rect 6934 -21076 7422 -21070
rect 7144 -21126 7204 -21076
rect 7138 -21186 7144 -21126
rect 7204 -21186 7210 -21126
rect 6634 -21402 6640 -21342
rect 6700 -21402 6706 -21342
rect 5614 -21500 5620 -21440
rect 5680 -21500 5686 -21440
rect 7144 -21554 7204 -21186
rect 7660 -21440 7720 -20986
rect 8678 -20986 8688 -20942
rect 8722 -20942 8728 -20410
rect 9688 -20410 9748 -20278
rect 10204 -20320 10264 -20174
rect 9988 -20326 10476 -20320
rect 9988 -20360 10000 -20326
rect 10464 -20360 10476 -20326
rect 9988 -20366 10476 -20360
rect 9688 -20474 9706 -20410
rect 8722 -20986 8738 -20942
rect 7952 -21036 8440 -21030
rect 7952 -21070 7964 -21036
rect 8428 -21070 8440 -21036
rect 7952 -21076 8440 -21070
rect 8162 -21126 8222 -21076
rect 8678 -21120 8738 -20986
rect 9700 -20986 9706 -20474
rect 9740 -20474 9748 -20410
rect 10710 -20410 10770 -19952
rect 11218 -20114 11278 -19842
rect 11212 -20174 11218 -20114
rect 11278 -20174 11284 -20114
rect 11218 -20320 11278 -20174
rect 11730 -20218 11790 -19752
rect 12746 -19752 12760 -19720
rect 12794 -19720 12800 -19176
rect 13772 -19176 13818 -19164
rect 13772 -19718 13778 -19176
rect 12794 -19752 12806 -19720
rect 12024 -19802 12512 -19796
rect 12024 -19836 12036 -19802
rect 12500 -19836 12512 -19802
rect 12024 -19842 12512 -19836
rect 12226 -20114 12286 -19842
rect 12746 -19892 12806 -19752
rect 13768 -19752 13778 -19718
rect 13812 -19718 13818 -19176
rect 14790 -19176 14836 -19164
rect 13812 -19752 13828 -19718
rect 14790 -19720 14796 -19176
rect 13042 -19802 13530 -19796
rect 13042 -19836 13054 -19802
rect 13518 -19836 13530 -19802
rect 13042 -19842 13530 -19836
rect 12740 -19952 12746 -19892
rect 12806 -19952 12812 -19892
rect 13270 -20114 13330 -19842
rect 12220 -20174 12226 -20114
rect 12286 -20174 12292 -20114
rect 13264 -20174 13270 -20114
rect 13330 -20174 13336 -20114
rect 11724 -20278 11730 -20218
rect 11790 -20278 11796 -20218
rect 11006 -20326 11494 -20320
rect 11006 -20360 11018 -20326
rect 11482 -20360 11494 -20326
rect 11006 -20366 11494 -20360
rect 10710 -20446 10724 -20410
rect 9740 -20986 9746 -20474
rect 10718 -20928 10724 -20446
rect 9700 -20998 9746 -20986
rect 10714 -20986 10724 -20928
rect 10758 -20446 10770 -20410
rect 11730 -20410 11790 -20278
rect 12226 -20320 12286 -20174
rect 13270 -20320 13330 -20174
rect 13768 -20218 13828 -19752
rect 14782 -19752 14796 -19720
rect 14830 -19720 14836 -19176
rect 15802 -19176 15862 -19044
rect 16096 -19092 16584 -19086
rect 16096 -19126 16108 -19092
rect 16572 -19126 16584 -19092
rect 16096 -19132 16584 -19126
rect 14830 -19752 14842 -19720
rect 14060 -19802 14548 -19796
rect 14060 -19836 14072 -19802
rect 14536 -19836 14548 -19802
rect 14060 -19842 14548 -19836
rect 14260 -20114 14320 -19842
rect 14782 -19892 14842 -19752
rect 15802 -19752 15814 -19176
rect 15848 -19752 15862 -19176
rect 16818 -19176 16878 -18520
rect 17838 -18520 17850 -18486
rect 17884 -17984 17896 -17944
rect 18854 -17944 18914 -17804
rect 19360 -17854 19420 -17740
rect 20376 -17854 20436 -17740
rect 20886 -17804 20892 -17744
rect 20952 -17804 20958 -17744
rect 19150 -17860 19638 -17854
rect 19150 -17894 19162 -17860
rect 19626 -17894 19638 -17860
rect 19150 -17900 19638 -17894
rect 20168 -17860 20656 -17854
rect 20168 -17894 20180 -17860
rect 20644 -17894 20656 -17860
rect 20168 -17900 20656 -17894
rect 17884 -18486 17890 -17984
rect 18854 -17986 18868 -17944
rect 17884 -18520 17898 -18486
rect 17114 -18570 17602 -18564
rect 17114 -18604 17126 -18570
rect 17590 -18604 17602 -18570
rect 17114 -18610 17602 -18604
rect 17314 -18880 17374 -18610
rect 17308 -18940 17314 -18880
rect 17374 -18940 17380 -18880
rect 17314 -19086 17374 -18940
rect 17114 -19092 17602 -19086
rect 17114 -19126 17126 -19092
rect 17590 -19126 17602 -19092
rect 17114 -19132 17602 -19126
rect 16818 -19216 16832 -19176
rect 16826 -19720 16832 -19216
rect 15078 -19802 15566 -19796
rect 15078 -19836 15090 -19802
rect 15554 -19836 15566 -19802
rect 15078 -19842 15566 -19836
rect 14776 -19952 14782 -19892
rect 14842 -19952 14848 -19892
rect 15278 -20114 15338 -19842
rect 14254 -20174 14260 -20114
rect 14320 -20174 14326 -20114
rect 15272 -20174 15278 -20114
rect 15338 -20174 15344 -20114
rect 13762 -20278 13768 -20218
rect 13828 -20278 13834 -20218
rect 12024 -20326 12512 -20320
rect 12024 -20360 12036 -20326
rect 12500 -20360 12512 -20326
rect 12024 -20366 12512 -20360
rect 13042 -20326 13530 -20320
rect 13042 -20360 13054 -20326
rect 13518 -20360 13530 -20326
rect 13042 -20366 13530 -20360
rect 10758 -20928 10764 -20446
rect 11730 -20448 11742 -20410
rect 10758 -20986 10774 -20928
rect 8970 -21036 9458 -21030
rect 8970 -21070 8982 -21036
rect 9446 -21070 9458 -21036
rect 8970 -21076 9458 -21070
rect 9988 -21036 10476 -21030
rect 9988 -21070 10000 -21036
rect 10464 -21070 10476 -21036
rect 9988 -21076 10476 -21070
rect 10714 -21120 10774 -20986
rect 11736 -20986 11742 -20448
rect 11776 -20448 11790 -20410
rect 12754 -20410 12800 -20398
rect 11776 -20986 11782 -20448
rect 12754 -20936 12760 -20410
rect 11736 -20998 11782 -20986
rect 12746 -20986 12760 -20936
rect 12794 -20936 12800 -20410
rect 13768 -20410 13828 -20278
rect 14260 -20320 14320 -20174
rect 15802 -20218 15862 -19752
rect 16820 -19752 16832 -19720
rect 16866 -19216 16878 -19176
rect 17838 -19176 17898 -18520
rect 18862 -18520 18868 -17986
rect 18902 -17986 18914 -17944
rect 19880 -17944 19926 -17932
rect 18902 -18520 18908 -17986
rect 19880 -18462 19886 -17944
rect 18862 -18532 18908 -18520
rect 19872 -18520 19886 -18462
rect 19920 -18462 19926 -17944
rect 20892 -17944 20952 -17804
rect 21394 -17854 21454 -17376
rect 21910 -17414 21970 -17286
rect 22928 -17286 22940 -17228
rect 22974 -16738 22986 -16710
rect 22974 -17228 22980 -16738
rect 22974 -17286 22988 -17228
rect 22204 -17336 22692 -17330
rect 22204 -17370 22216 -17336
rect 22680 -17370 22692 -17336
rect 22204 -17376 22692 -17370
rect 22928 -17396 22988 -17286
rect 21904 -17474 21910 -17414
rect 21970 -17474 21976 -17414
rect 22922 -17456 22928 -17396
rect 22988 -17456 22994 -17396
rect 21910 -17692 21970 -17474
rect 21910 -17752 22984 -17692
rect 23034 -17744 23094 -16568
rect 23156 -16586 23162 -16526
rect 23222 -16586 23228 -16526
rect 23528 -17526 23588 -13640
rect 23522 -17586 23528 -17526
rect 23588 -17586 23594 -17526
rect 23272 -17690 23278 -17630
rect 23338 -17690 23344 -17630
rect 21186 -17860 21674 -17854
rect 21186 -17894 21198 -17860
rect 21662 -17894 21674 -17860
rect 21186 -17900 21674 -17894
rect 20892 -17986 20904 -17944
rect 19920 -18520 19932 -18462
rect 18344 -18564 18404 -18562
rect 18132 -18570 18620 -18564
rect 18132 -18604 18144 -18570
rect 18608 -18604 18620 -18570
rect 18132 -18610 18620 -18604
rect 19150 -18570 19638 -18564
rect 19150 -18604 19162 -18570
rect 19626 -18604 19638 -18570
rect 19150 -18610 19638 -18604
rect 18344 -18880 18404 -18610
rect 19366 -18658 19426 -18610
rect 19360 -18718 19366 -18658
rect 19426 -18718 19432 -18658
rect 19498 -18714 19504 -18654
rect 19564 -18714 19570 -18654
rect 19504 -18880 19564 -18714
rect 19872 -18880 19932 -18520
rect 20898 -18520 20904 -17986
rect 20938 -17986 20952 -17944
rect 21910 -17944 21970 -17752
rect 22414 -17854 22474 -17752
rect 22204 -17860 22692 -17854
rect 22204 -17894 22216 -17860
rect 22680 -17894 22692 -17860
rect 22204 -17900 22692 -17894
rect 21910 -17978 21922 -17944
rect 20938 -18520 20944 -17986
rect 21916 -18480 21922 -17978
rect 20898 -18532 20944 -18520
rect 21910 -18520 21922 -18480
rect 21956 -17978 21970 -17944
rect 22924 -17944 22984 -17752
rect 23028 -17804 23034 -17744
rect 23094 -17804 23100 -17744
rect 22924 -17968 22940 -17944
rect 21956 -18480 21962 -17978
rect 21956 -18520 21970 -18480
rect 20168 -18570 20656 -18564
rect 20168 -18604 20180 -18570
rect 20644 -18604 20656 -18570
rect 20168 -18610 20656 -18604
rect 21186 -18570 21674 -18564
rect 21186 -18604 21198 -18570
rect 21662 -18604 21674 -18570
rect 21186 -18610 21674 -18604
rect 21392 -18654 21452 -18610
rect 20380 -18714 20386 -18654
rect 20446 -18714 20452 -18654
rect 21386 -18714 21392 -18654
rect 21452 -18714 21458 -18654
rect 21910 -18658 21970 -18520
rect 22934 -18520 22940 -17968
rect 22974 -17968 22984 -17944
rect 22974 -18520 22980 -17968
rect 22934 -18532 22980 -18520
rect 22204 -18570 22692 -18564
rect 22204 -18604 22216 -18570
rect 22680 -18604 22692 -18570
rect 22204 -18610 22692 -18604
rect 18338 -18940 18344 -18880
rect 18404 -18940 18410 -18880
rect 19498 -18940 19504 -18880
rect 19564 -18940 19570 -18880
rect 19866 -18940 19872 -18880
rect 19932 -18940 19938 -18880
rect 18344 -19086 18404 -18940
rect 19504 -19086 19564 -18940
rect 19872 -18984 19932 -18940
rect 19866 -19044 19872 -18984
rect 19932 -19044 19938 -18984
rect 20386 -19086 20446 -18714
rect 21904 -18718 21910 -18658
rect 21970 -18718 21976 -18658
rect 21904 -18846 21910 -18786
rect 21970 -18846 21976 -18786
rect 20882 -19042 20888 -18982
rect 20948 -19042 20954 -18982
rect 18132 -19092 18620 -19086
rect 18132 -19126 18144 -19092
rect 18608 -19126 18620 -19092
rect 18132 -19132 18620 -19126
rect 19150 -19092 19638 -19086
rect 19150 -19126 19162 -19092
rect 19626 -19126 19638 -19092
rect 19150 -19132 19638 -19126
rect 20168 -19092 20656 -19086
rect 20168 -19126 20180 -19092
rect 20644 -19126 20656 -19092
rect 20168 -19132 20656 -19126
rect 20386 -19134 20446 -19132
rect 16866 -19720 16872 -19216
rect 17838 -19222 17850 -19176
rect 17844 -19708 17850 -19222
rect 16866 -19752 16880 -19720
rect 16096 -19802 16584 -19796
rect 16096 -19836 16108 -19802
rect 16572 -19836 16584 -19802
rect 16096 -19842 16584 -19836
rect 16312 -20114 16372 -19842
rect 16820 -19892 16880 -19752
rect 17836 -19752 17850 -19708
rect 17884 -19222 17898 -19176
rect 18862 -19176 18908 -19164
rect 17884 -19708 17890 -19222
rect 17884 -19752 17896 -19708
rect 18862 -19712 18868 -19176
rect 17114 -19802 17602 -19796
rect 17114 -19836 17126 -19802
rect 17590 -19836 17602 -19802
rect 17114 -19842 17602 -19836
rect 16814 -19952 16820 -19892
rect 16880 -19952 16886 -19892
rect 16806 -20060 16812 -20000
rect 16872 -20060 16878 -20000
rect 16306 -20174 16312 -20114
rect 16372 -20174 16378 -20114
rect 15796 -20278 15802 -20218
rect 15862 -20278 15868 -20218
rect 16308 -20282 16314 -20222
rect 16374 -20282 16380 -20222
rect 16314 -20320 16374 -20282
rect 14060 -20326 14548 -20320
rect 14060 -20360 14072 -20326
rect 14536 -20360 14548 -20326
rect 14060 -20366 14548 -20360
rect 15078 -20326 15566 -20320
rect 15078 -20360 15090 -20326
rect 15554 -20360 15566 -20326
rect 15078 -20366 15566 -20360
rect 16096 -20326 16584 -20320
rect 16096 -20360 16108 -20326
rect 16572 -20360 16584 -20326
rect 16096 -20366 16584 -20360
rect 13768 -20446 13778 -20410
rect 12794 -20986 12806 -20936
rect 11006 -21036 11494 -21030
rect 11006 -21070 11018 -21036
rect 11482 -21070 11494 -21036
rect 11006 -21076 11494 -21070
rect 12024 -21036 12512 -21030
rect 12024 -21070 12036 -21036
rect 12500 -21070 12512 -21036
rect 12024 -21076 12512 -21070
rect 12746 -21120 12806 -20986
rect 13772 -20986 13778 -20446
rect 13812 -20446 13828 -20410
rect 14790 -20410 14836 -20398
rect 13812 -20986 13818 -20446
rect 14790 -20924 14796 -20410
rect 13772 -20998 13818 -20986
rect 14780 -20986 14796 -20924
rect 14830 -20924 14836 -20410
rect 15808 -20410 15854 -20398
rect 14830 -20986 14840 -20924
rect 15808 -20944 15814 -20410
rect 13042 -21036 13530 -21030
rect 13042 -21070 13054 -21036
rect 13518 -21070 13530 -21036
rect 13042 -21076 13530 -21070
rect 14060 -21036 14548 -21030
rect 14060 -21070 14072 -21036
rect 14536 -21070 14548 -21036
rect 14060 -21076 14548 -21070
rect 14780 -21120 14840 -20986
rect 15802 -20986 15814 -20944
rect 15848 -20944 15854 -20410
rect 16812 -20410 16872 -20060
rect 17336 -20222 17396 -19842
rect 17836 -20216 17896 -19752
rect 18856 -19752 18868 -19712
rect 18902 -19712 18908 -19176
rect 19880 -19176 19926 -19164
rect 19880 -19708 19886 -19176
rect 18902 -19752 18916 -19712
rect 18132 -19802 18620 -19796
rect 18132 -19836 18144 -19802
rect 18608 -19836 18620 -19802
rect 18132 -19842 18620 -19836
rect 17330 -20282 17336 -20222
rect 17396 -20282 17402 -20222
rect 17830 -20276 17836 -20216
rect 17896 -20276 17902 -20216
rect 17336 -20320 17396 -20282
rect 17114 -20326 17602 -20320
rect 17114 -20360 17126 -20326
rect 17590 -20360 17602 -20326
rect 17114 -20366 17602 -20360
rect 16812 -20446 16832 -20410
rect 15848 -20986 15862 -20944
rect 15078 -21036 15566 -21030
rect 15078 -21070 15090 -21036
rect 15554 -21070 15566 -21036
rect 15078 -21076 15566 -21070
rect 8156 -21186 8162 -21126
rect 8222 -21186 8228 -21126
rect 8672 -21180 8678 -21120
rect 8738 -21180 8744 -21120
rect 12740 -21180 12746 -21120
rect 12806 -21180 12812 -21120
rect 14774 -21180 14780 -21120
rect 14840 -21180 14846 -21120
rect 7654 -21500 7660 -21440
rect 7720 -21500 7726 -21440
rect 3880 -21560 4368 -21554
rect 3880 -21594 3892 -21560
rect 4356 -21594 4368 -21560
rect 3880 -21600 4368 -21594
rect 4898 -21560 5386 -21554
rect 4898 -21594 4910 -21560
rect 5374 -21594 5386 -21560
rect 4898 -21600 5386 -21594
rect 5916 -21560 6404 -21554
rect 5916 -21594 5928 -21560
rect 6392 -21594 6404 -21560
rect 5916 -21600 6404 -21594
rect 6934 -21560 7422 -21554
rect 6934 -21594 6946 -21560
rect 7410 -21594 7422 -21560
rect 6934 -21600 7422 -21594
rect 3582 -21698 3598 -21644
rect 2614 -22220 2624 -22186
rect 3592 -22190 3598 -21698
rect 2564 -22352 2624 -22220
rect 3588 -22220 3598 -22190
rect 3632 -21698 3642 -21644
rect 4610 -21644 4656 -21632
rect 3632 -22190 3638 -21698
rect 4610 -22174 4616 -21644
rect 3632 -22220 3648 -22190
rect 2862 -22270 3350 -22264
rect 2862 -22304 2874 -22270
rect 3338 -22304 3350 -22270
rect 2862 -22310 3350 -22304
rect 3084 -22352 3144 -22310
rect 3588 -22352 3648 -22220
rect 4602 -22220 4616 -22174
rect 4650 -22174 4656 -21644
rect 5628 -21644 5674 -21632
rect 4650 -22220 4662 -22174
rect 5628 -22190 5634 -21644
rect 3880 -22270 4368 -22264
rect 3880 -22304 3892 -22270
rect 4356 -22304 4368 -22270
rect 3880 -22310 4368 -22304
rect 2564 -22412 3648 -22352
rect 2442 -22522 2448 -22462
rect 2508 -22522 2514 -22462
rect 3588 -22558 3648 -22412
rect 2564 -22618 3648 -22558
rect 2564 -22876 2624 -22618
rect 3076 -22786 3136 -22618
rect 3588 -22678 3648 -22618
rect 3582 -22738 3588 -22678
rect 3648 -22738 3654 -22678
rect 2862 -22792 3350 -22786
rect 2862 -22826 2874 -22792
rect 3338 -22826 3350 -22792
rect 2862 -22832 3350 -22826
rect 2564 -22912 2580 -22876
rect 2574 -23452 2580 -22912
rect 2614 -22912 2624 -22876
rect 3588 -22876 3648 -22738
rect 4080 -22786 4140 -22310
rect 4602 -22364 4662 -22220
rect 5620 -22220 5634 -22190
rect 5668 -22190 5674 -21644
rect 6646 -21644 6692 -21632
rect 6646 -22178 6652 -21644
rect 5668 -22220 5680 -22190
rect 4898 -22270 5386 -22264
rect 4898 -22304 4910 -22270
rect 5374 -22304 5386 -22270
rect 4898 -22310 5386 -22304
rect 4596 -22424 4602 -22364
rect 4662 -22424 4668 -22364
rect 4600 -22618 4606 -22558
rect 4666 -22618 4672 -22558
rect 3880 -22792 4368 -22786
rect 3880 -22826 3892 -22792
rect 4356 -22826 4368 -22792
rect 3880 -22832 4368 -22826
rect 2614 -23452 2620 -22912
rect 3588 -22916 3598 -22876
rect 2574 -23464 2620 -23452
rect 3592 -23452 3598 -22916
rect 3632 -22916 3648 -22876
rect 4606 -22876 4666 -22618
rect 5100 -22622 5160 -22310
rect 5620 -22462 5680 -22220
rect 6638 -22220 6652 -22178
rect 6686 -22178 6692 -21644
rect 7660 -21644 7720 -21500
rect 8162 -21554 8222 -21186
rect 7952 -21560 8440 -21554
rect 7952 -21594 7964 -21560
rect 8428 -21594 8440 -21560
rect 7952 -21600 8440 -21594
rect 7660 -21674 7670 -21644
rect 7664 -22156 7670 -21674
rect 6686 -22220 6698 -22178
rect 5916 -22270 6404 -22264
rect 5916 -22304 5928 -22270
rect 6392 -22304 6404 -22270
rect 5916 -22310 6404 -22304
rect 5614 -22522 5620 -22462
rect 5680 -22522 5686 -22462
rect 6134 -22622 6194 -22310
rect 6638 -22364 6698 -22220
rect 7656 -22220 7670 -22156
rect 7704 -21674 7720 -21644
rect 8678 -21644 8738 -21180
rect 10714 -21186 10774 -21180
rect 11724 -21290 11730 -21230
rect 11790 -21290 11796 -21230
rect 13760 -21290 13766 -21230
rect 13826 -21290 13832 -21230
rect 10706 -21402 10712 -21342
rect 10772 -21402 10778 -21342
rect 9690 -21500 9696 -21440
rect 9756 -21500 9762 -21440
rect 8970 -21560 9458 -21554
rect 8970 -21594 8982 -21560
rect 9446 -21594 9458 -21560
rect 8970 -21600 9458 -21594
rect 7704 -22156 7710 -21674
rect 8678 -21686 8688 -21644
rect 7704 -22220 7716 -22156
rect 8682 -22180 8688 -21686
rect 6934 -22270 7422 -22264
rect 6934 -22304 6946 -22270
rect 7410 -22304 7422 -22270
rect 6934 -22310 7422 -22304
rect 6632 -22424 6638 -22364
rect 6698 -22424 6704 -22364
rect 7144 -22462 7204 -22310
rect 7138 -22522 7144 -22462
rect 7204 -22522 7210 -22462
rect 6636 -22618 6642 -22558
rect 6702 -22618 6708 -22558
rect 5100 -22682 6194 -22622
rect 5100 -22786 5160 -22682
rect 6134 -22786 6194 -22682
rect 4898 -22792 5386 -22786
rect 4898 -22826 4910 -22792
rect 5374 -22826 5386 -22792
rect 4898 -22832 5386 -22826
rect 5916 -22792 6404 -22786
rect 5916 -22826 5928 -22792
rect 6392 -22826 6404 -22792
rect 5916 -22832 6404 -22826
rect 3632 -23452 3638 -22916
rect 4606 -22920 4616 -22876
rect 3592 -23464 3638 -23452
rect 4610 -23452 4616 -22920
rect 4650 -22920 4666 -22876
rect 5628 -22876 5674 -22864
rect 4650 -23452 4656 -22920
rect 5628 -23410 5634 -22876
rect 4610 -23464 4656 -23452
rect 5620 -23452 5634 -23410
rect 5668 -23410 5674 -22876
rect 6642 -22876 6702 -22618
rect 7144 -22786 7204 -22522
rect 7656 -22678 7716 -22220
rect 8676 -22220 8688 -22180
rect 8722 -21686 8738 -21644
rect 9696 -21644 9756 -21500
rect 9988 -21560 10476 -21554
rect 9988 -21594 10000 -21560
rect 10464 -21594 10476 -21560
rect 9988 -21600 10476 -21594
rect 9696 -21680 9706 -21644
rect 8722 -22180 8728 -21686
rect 8722 -22220 8736 -22180
rect 9700 -22186 9706 -21680
rect 7952 -22270 8440 -22264
rect 7952 -22304 7964 -22270
rect 8428 -22304 8440 -22270
rect 7952 -22310 8440 -22304
rect 8166 -22462 8226 -22310
rect 8676 -22364 8736 -22220
rect 9690 -22220 9706 -22186
rect 9740 -21680 9756 -21644
rect 10712 -21644 10772 -21402
rect 11006 -21560 11494 -21554
rect 11006 -21594 11018 -21560
rect 11482 -21594 11494 -21560
rect 11006 -21600 11494 -21594
rect 10712 -21670 10724 -21644
rect 9740 -22186 9746 -21680
rect 10718 -22164 10724 -21670
rect 9740 -22220 9750 -22186
rect 8970 -22270 9458 -22264
rect 8970 -22304 8982 -22270
rect 9446 -22304 9458 -22270
rect 8970 -22310 9458 -22304
rect 8670 -22424 8676 -22364
rect 8736 -22424 8742 -22364
rect 9190 -22456 9250 -22310
rect 7650 -22738 7656 -22678
rect 7716 -22738 7722 -22678
rect 6934 -22792 7422 -22786
rect 6934 -22826 6946 -22792
rect 7410 -22826 7422 -22792
rect 6934 -22832 7422 -22826
rect 6642 -22928 6652 -22876
rect 5668 -23452 5680 -23410
rect 2862 -23502 3350 -23496
rect 2862 -23536 2874 -23502
rect 3338 -23536 3350 -23502
rect 2862 -23542 3350 -23536
rect 3880 -23502 4368 -23496
rect 3880 -23536 3892 -23502
rect 4356 -23536 4368 -23502
rect 3880 -23542 4368 -23536
rect 4898 -23502 5386 -23496
rect 4898 -23536 4910 -23502
rect 5374 -23536 5386 -23502
rect 4898 -23542 5386 -23536
rect 2330 -23654 2336 -23594
rect 2396 -23654 2402 -23594
rect 2224 -23780 2230 -23720
rect 2290 -23780 2296 -23720
rect 2564 -23960 3644 -23900
rect 2564 -24110 2624 -23960
rect 3072 -24020 3132 -23960
rect 2862 -24026 3350 -24020
rect 2862 -24060 2874 -24026
rect 3338 -24060 3350 -24026
rect 2862 -24066 3350 -24060
rect 2564 -24166 2580 -24110
rect 2574 -24686 2580 -24166
rect 2614 -24166 2624 -24110
rect 3584 -24110 3644 -23960
rect 4082 -24020 4142 -23542
rect 5620 -23720 5680 -23452
rect 6646 -23452 6652 -22928
rect 6686 -22928 6702 -22876
rect 7656 -22876 7716 -22738
rect 8166 -22786 8226 -22522
rect 9188 -22462 9250 -22456
rect 9248 -22522 9250 -22462
rect 9188 -22528 9250 -22522
rect 8664 -22618 8670 -22558
rect 8730 -22618 8736 -22558
rect 7952 -22792 8440 -22786
rect 7952 -22826 7964 -22792
rect 8428 -22826 8440 -22792
rect 7952 -22832 8440 -22826
rect 7656 -22916 7670 -22876
rect 6686 -23452 6692 -22928
rect 7664 -23398 7670 -22916
rect 6646 -23464 6692 -23452
rect 7658 -23452 7670 -23398
rect 7704 -22916 7716 -22876
rect 8670 -22876 8730 -22618
rect 9190 -22786 9250 -22528
rect 9690 -22678 9750 -22220
rect 10708 -22220 10724 -22164
rect 10758 -21670 10772 -21644
rect 11730 -21644 11790 -21290
rect 12024 -21560 12512 -21554
rect 12024 -21594 12036 -21560
rect 12500 -21594 12512 -21560
rect 12024 -21600 12512 -21594
rect 13042 -21560 13530 -21554
rect 13042 -21594 13054 -21560
rect 13518 -21594 13530 -21560
rect 13042 -21600 13530 -21594
rect 10758 -22164 10764 -21670
rect 11730 -21676 11742 -21644
rect 10758 -22220 10768 -22164
rect 9988 -22270 10476 -22264
rect 9988 -22304 10000 -22270
rect 10464 -22304 10476 -22270
rect 9988 -22310 10476 -22304
rect 10192 -22462 10252 -22310
rect 10538 -22344 10598 -22338
rect 10708 -22344 10768 -22220
rect 11736 -22220 11742 -21676
rect 11776 -21676 11790 -21644
rect 12754 -21644 12800 -21632
rect 11776 -22220 11782 -21676
rect 12754 -22150 12760 -21644
rect 11736 -22232 11782 -22220
rect 12750 -22220 12760 -22150
rect 12794 -22150 12800 -21644
rect 13766 -21644 13826 -21290
rect 15308 -21328 15368 -21076
rect 15802 -21118 15862 -20986
rect 16826 -20986 16832 -20446
rect 16866 -20986 16872 -20410
rect 17836 -20410 17896 -20276
rect 18314 -20320 18374 -19842
rect 18856 -19892 18916 -19752
rect 19870 -19752 19886 -19708
rect 19920 -19708 19926 -19176
rect 20888 -19176 20948 -19042
rect 21186 -19092 21674 -19086
rect 21186 -19126 21198 -19092
rect 21662 -19126 21674 -19092
rect 21186 -19132 21674 -19126
rect 20888 -19226 20904 -19176
rect 19920 -19752 19930 -19708
rect 20898 -19724 20904 -19226
rect 19150 -19802 19638 -19796
rect 19150 -19836 19162 -19802
rect 19626 -19836 19638 -19802
rect 19150 -19842 19638 -19836
rect 18850 -19952 18856 -19892
rect 18916 -19952 18922 -19892
rect 18846 -20060 18852 -20000
rect 18912 -20060 18918 -20000
rect 18132 -20326 18620 -20320
rect 18132 -20360 18144 -20326
rect 18608 -20360 18620 -20326
rect 18132 -20366 18620 -20360
rect 17836 -20504 17850 -20410
rect 17844 -20944 17850 -20504
rect 16826 -20998 16872 -20986
rect 17836 -20986 17850 -20944
rect 17884 -20504 17896 -20410
rect 18852 -20410 18912 -20060
rect 19338 -20174 19344 -20114
rect 19404 -20174 19410 -20114
rect 19344 -20320 19404 -20174
rect 19870 -20216 19930 -19752
rect 20894 -19752 20904 -19724
rect 20938 -19226 20948 -19176
rect 21910 -19176 21970 -18846
rect 22204 -19092 22692 -19086
rect 22204 -19126 22216 -19092
rect 22680 -19126 22692 -19092
rect 22204 -19132 22692 -19126
rect 20938 -19724 20944 -19226
rect 21910 -19228 21922 -19176
rect 21916 -19724 21922 -19228
rect 20938 -19752 20954 -19724
rect 20168 -19802 20656 -19796
rect 20168 -19836 20180 -19802
rect 20644 -19836 20656 -19802
rect 20168 -19842 20656 -19836
rect 20894 -19892 20954 -19752
rect 21910 -19752 21922 -19724
rect 21956 -19228 21970 -19176
rect 22934 -19176 22980 -19164
rect 21956 -19724 21962 -19228
rect 22934 -19718 22940 -19176
rect 21956 -19752 21970 -19724
rect 21186 -19802 21674 -19796
rect 21186 -19836 21198 -19802
rect 21662 -19836 21674 -19802
rect 21186 -19842 21674 -19836
rect 20888 -19952 20894 -19892
rect 20954 -19952 20960 -19892
rect 20884 -20060 20890 -20000
rect 20950 -20060 20956 -20000
rect 20376 -20174 20382 -20114
rect 20442 -20174 20448 -20114
rect 19864 -20276 19870 -20216
rect 19930 -20276 19936 -20216
rect 20382 -20320 20442 -20174
rect 19150 -20326 19638 -20320
rect 19150 -20360 19162 -20326
rect 19626 -20360 19638 -20326
rect 19150 -20366 19638 -20360
rect 20168 -20326 20656 -20320
rect 20168 -20360 20180 -20326
rect 20644 -20360 20656 -20326
rect 20168 -20366 20656 -20360
rect 18852 -20476 18868 -20410
rect 17884 -20944 17890 -20504
rect 17884 -20986 17896 -20944
rect 16096 -21036 16584 -21030
rect 16096 -21070 16108 -21036
rect 16572 -21070 16584 -21036
rect 16096 -21076 16584 -21070
rect 17114 -21036 17602 -21030
rect 17114 -21070 17126 -21036
rect 17590 -21070 17602 -21036
rect 17114 -21076 17602 -21070
rect 15796 -21178 15802 -21118
rect 15862 -21178 15868 -21118
rect 16150 -21178 16156 -21118
rect 16216 -21178 16222 -21118
rect 15792 -21290 15798 -21230
rect 15858 -21290 15864 -21230
rect 15302 -21388 15308 -21328
rect 15368 -21388 15374 -21328
rect 14060 -21560 14548 -21554
rect 14060 -21594 14072 -21560
rect 14536 -21594 14548 -21560
rect 14060 -21600 14548 -21594
rect 15078 -21560 15566 -21554
rect 15078 -21594 15090 -21560
rect 15554 -21594 15566 -21560
rect 15078 -21600 15566 -21594
rect 13766 -21682 13778 -21644
rect 12794 -22220 12810 -22150
rect 11006 -22270 11494 -22264
rect 11006 -22304 11018 -22270
rect 11482 -22304 11494 -22270
rect 11006 -22310 11494 -22304
rect 12024 -22270 12512 -22264
rect 12024 -22304 12036 -22270
rect 12500 -22304 12512 -22270
rect 12024 -22310 12512 -22304
rect 10702 -22404 10708 -22344
rect 10768 -22404 10774 -22344
rect 10186 -22522 10192 -22462
rect 10252 -22522 10258 -22462
rect 9684 -22738 9690 -22678
rect 9750 -22738 9756 -22678
rect 8970 -22792 9458 -22786
rect 8970 -22826 8982 -22792
rect 9446 -22826 9458 -22792
rect 8970 -22832 9458 -22826
rect 7704 -23398 7710 -22916
rect 8670 -22936 8688 -22876
rect 7704 -23452 7718 -23398
rect 5916 -23502 6404 -23496
rect 5916 -23536 5928 -23502
rect 6392 -23536 6404 -23502
rect 5916 -23542 6404 -23536
rect 6934 -23502 7422 -23496
rect 6934 -23536 6946 -23502
rect 7410 -23536 7422 -23502
rect 6934 -23542 7422 -23536
rect 6140 -23708 6200 -23542
rect 5614 -23780 5620 -23720
rect 5680 -23780 5686 -23720
rect 6134 -23768 6140 -23708
rect 6200 -23768 6206 -23708
rect 4596 -23882 4602 -23822
rect 4662 -23882 4668 -23822
rect 6632 -23882 6638 -23822
rect 6698 -23882 6704 -23822
rect 3880 -24026 4368 -24020
rect 3880 -24060 3892 -24026
rect 4356 -24060 4368 -24026
rect 3880 -24066 4368 -24060
rect 2614 -24686 2620 -24166
rect 2574 -24698 2620 -24686
rect 3584 -24686 3598 -24110
rect 3632 -24686 3644 -24110
rect 4602 -24110 4662 -23882
rect 5614 -23986 5620 -23926
rect 5680 -23986 5686 -23926
rect 4898 -24026 5386 -24020
rect 4898 -24060 4910 -24026
rect 5374 -24060 5386 -24026
rect 4898 -24066 5386 -24060
rect 4602 -24170 4616 -24110
rect 4610 -24650 4616 -24170
rect 2862 -24736 3350 -24730
rect 2862 -24770 2874 -24736
rect 3338 -24770 3350 -24736
rect 2862 -24776 3350 -24770
rect 2442 -24884 2448 -24824
rect 2508 -24884 2514 -24824
rect 2114 -24988 2120 -24928
rect 2180 -24988 2186 -24928
rect 2448 -25154 2508 -24884
rect 3584 -24928 3644 -24686
rect 4604 -24686 4616 -24650
rect 4650 -24170 4662 -24110
rect 5620 -24110 5680 -23986
rect 5916 -24026 6404 -24020
rect 5916 -24060 5928 -24026
rect 6392 -24060 6404 -24026
rect 5916 -24066 6404 -24060
rect 5620 -24164 5634 -24110
rect 4650 -24650 4656 -24170
rect 5628 -24646 5634 -24164
rect 4650 -24686 4664 -24650
rect 3880 -24736 4368 -24730
rect 3880 -24770 3892 -24736
rect 4356 -24770 4368 -24736
rect 3880 -24776 4368 -24770
rect 3578 -24988 3584 -24928
rect 3644 -24988 3650 -24928
rect 4092 -25034 4152 -24776
rect 4086 -25094 4092 -25034
rect 4152 -25094 4158 -25034
rect 2448 -25214 3648 -25154
rect 1064 -26048 1070 -25988
rect 1130 -26048 1136 -25988
rect 2448 -26066 2508 -25214
rect 2568 -25342 2628 -25214
rect 3054 -25252 3114 -25214
rect 2862 -25258 3350 -25252
rect 2862 -25292 2874 -25258
rect 3338 -25292 3350 -25258
rect 2862 -25298 3350 -25292
rect 2568 -25414 2580 -25342
rect 2574 -25918 2580 -25414
rect 2614 -25414 2628 -25342
rect 3588 -25342 3648 -25214
rect 4092 -25252 4152 -25094
rect 4604 -25144 4664 -24686
rect 5618 -24686 5634 -24646
rect 5668 -24164 5680 -24110
rect 6638 -24110 6698 -23882
rect 7140 -24020 7200 -23542
rect 7658 -23822 7718 -23452
rect 8682 -23452 8688 -22936
rect 8722 -22936 8730 -22876
rect 9690 -22876 9750 -22738
rect 10192 -22786 10252 -22522
rect 10538 -22558 10598 -22404
rect 10532 -22618 10538 -22558
rect 10598 -22618 10604 -22558
rect 10708 -22612 10714 -22552
rect 10774 -22612 10780 -22552
rect 9988 -22792 10476 -22786
rect 9988 -22826 10000 -22792
rect 10464 -22826 10476 -22792
rect 9988 -22832 10476 -22826
rect 9690 -22916 9706 -22876
rect 8722 -23452 8728 -22936
rect 9700 -23386 9706 -22916
rect 8682 -23464 8728 -23452
rect 9694 -23452 9706 -23386
rect 9740 -22916 9750 -22876
rect 10714 -22876 10774 -22612
rect 11230 -22614 11290 -22310
rect 12244 -22450 12304 -22310
rect 12750 -22344 12810 -22220
rect 13772 -22220 13778 -21682
rect 13812 -21682 13826 -21644
rect 14790 -21644 14836 -21632
rect 13812 -22220 13818 -21682
rect 14790 -22150 14796 -21644
rect 13772 -22232 13818 -22220
rect 14782 -22220 14796 -22150
rect 14830 -22150 14836 -21644
rect 15798 -21644 15858 -21290
rect 16156 -21436 16216 -21178
rect 16346 -21328 16406 -21076
rect 17322 -21328 17382 -21076
rect 16340 -21388 16346 -21328
rect 16406 -21388 16412 -21328
rect 17316 -21388 17322 -21328
rect 17382 -21388 17388 -21328
rect 17836 -21440 17896 -20986
rect 18862 -20986 18868 -20476
rect 18902 -20476 18912 -20410
rect 19880 -20410 19926 -20398
rect 18902 -20986 18908 -20476
rect 19880 -20942 19886 -20410
rect 18862 -20998 18908 -20986
rect 19874 -20986 19886 -20942
rect 19920 -20942 19926 -20410
rect 20890 -20410 20950 -20060
rect 21408 -20114 21468 -19842
rect 21910 -19934 21970 -19752
rect 22924 -19752 22940 -19718
rect 22974 -19718 22980 -19176
rect 22974 -19752 22984 -19718
rect 22204 -19802 22692 -19796
rect 22204 -19836 22216 -19802
rect 22680 -19836 22692 -19802
rect 22204 -19842 22692 -19836
rect 22418 -19934 22478 -19842
rect 22924 -19934 22984 -19752
rect 21910 -19994 22984 -19934
rect 21402 -20174 21408 -20114
rect 21468 -20174 21474 -20114
rect 21906 -20276 21912 -20216
rect 21972 -20276 21978 -20216
rect 21186 -20326 21674 -20320
rect 21186 -20360 21198 -20326
rect 21662 -20360 21674 -20326
rect 21186 -20366 21674 -20360
rect 20890 -20462 20904 -20410
rect 20898 -20936 20904 -20462
rect 19920 -20986 19934 -20942
rect 18132 -21036 18620 -21030
rect 18132 -21070 18144 -21036
rect 18608 -21070 18620 -21036
rect 18132 -21076 18620 -21070
rect 19150 -21036 19638 -21030
rect 19150 -21070 19162 -21036
rect 19626 -21070 19638 -21036
rect 19150 -21076 19638 -21070
rect 18338 -21328 18398 -21076
rect 19874 -21118 19934 -20986
rect 20892 -20986 20904 -20936
rect 20938 -20462 20950 -20410
rect 21912 -20410 21972 -20276
rect 22204 -20326 22692 -20320
rect 22204 -20360 22216 -20326
rect 22680 -20360 22692 -20326
rect 22204 -20366 22692 -20360
rect 21912 -20444 21922 -20410
rect 20938 -20936 20944 -20462
rect 20938 -20986 20952 -20936
rect 21916 -20942 21922 -20444
rect 20168 -21036 20656 -21030
rect 20168 -21070 20180 -21036
rect 20644 -21070 20656 -21036
rect 20168 -21076 20656 -21070
rect 19868 -21178 19874 -21118
rect 19934 -21178 19940 -21118
rect 18332 -21388 18338 -21328
rect 18398 -21388 18404 -21328
rect 20358 -21388 20364 -21328
rect 20424 -21388 20430 -21328
rect 16156 -21502 16216 -21496
rect 17830 -21500 17836 -21440
rect 17896 -21500 17902 -21440
rect 19866 -21500 19872 -21440
rect 19932 -21500 19938 -21440
rect 16096 -21560 16584 -21554
rect 16096 -21594 16108 -21560
rect 16572 -21594 16584 -21560
rect 16096 -21600 16584 -21594
rect 17114 -21560 17602 -21554
rect 17114 -21594 17126 -21560
rect 17590 -21594 17602 -21560
rect 17114 -21600 17602 -21594
rect 15798 -21686 15814 -21644
rect 14830 -22220 14842 -22150
rect 13042 -22270 13530 -22264
rect 13042 -22304 13054 -22270
rect 13518 -22304 13530 -22270
rect 13042 -22310 13530 -22304
rect 14060 -22270 14548 -22264
rect 14060 -22304 14072 -22270
rect 14536 -22304 14548 -22270
rect 14060 -22310 14548 -22304
rect 12744 -22404 12750 -22344
rect 12810 -22404 12816 -22344
rect 13266 -22450 13326 -22310
rect 14280 -22450 14340 -22310
rect 14782 -22344 14842 -22220
rect 15808 -22220 15814 -21686
rect 15848 -21686 15858 -21644
rect 16826 -21644 16872 -21632
rect 15848 -22220 15854 -21686
rect 16826 -22184 16832 -21644
rect 15808 -22232 15854 -22220
rect 16822 -22220 16832 -22184
rect 16866 -22184 16872 -21644
rect 17836 -21644 17896 -21500
rect 18132 -21560 18620 -21554
rect 18132 -21594 18144 -21560
rect 18608 -21594 18620 -21560
rect 18132 -21600 18620 -21594
rect 19150 -21560 19638 -21554
rect 19150 -21594 19162 -21560
rect 19626 -21594 19638 -21560
rect 19150 -21600 19638 -21594
rect 17836 -21682 17850 -21644
rect 17844 -22168 17850 -21682
rect 16866 -22220 16882 -22184
rect 15078 -22270 15566 -22264
rect 15078 -22304 15090 -22270
rect 15554 -22304 15566 -22270
rect 15078 -22310 15566 -22304
rect 16096 -22270 16584 -22264
rect 16096 -22304 16108 -22270
rect 16572 -22304 16584 -22270
rect 16096 -22310 16584 -22304
rect 14776 -22404 14782 -22344
rect 14842 -22404 14848 -22344
rect 15282 -22350 15342 -22310
rect 16308 -22350 16368 -22310
rect 16822 -22344 16882 -22220
rect 17840 -22220 17850 -22168
rect 17884 -21682 17896 -21644
rect 18862 -21644 18908 -21632
rect 17884 -22168 17890 -21682
rect 17884 -22220 17900 -22168
rect 18862 -22176 18868 -21644
rect 17114 -22270 17602 -22264
rect 17114 -22304 17126 -22270
rect 17590 -22304 17602 -22270
rect 17114 -22310 17602 -22304
rect 15282 -22410 16368 -22350
rect 16816 -22404 16822 -22344
rect 16882 -22404 16888 -22344
rect 15282 -22450 15342 -22410
rect 12244 -22510 15342 -22450
rect 15794 -22502 15800 -22442
rect 15860 -22502 15866 -22442
rect 12244 -22614 12304 -22510
rect 12736 -22612 12742 -22552
rect 12802 -22612 12808 -22552
rect 11230 -22674 12304 -22614
rect 11230 -22786 11290 -22674
rect 12244 -22786 12304 -22674
rect 11006 -22792 11494 -22786
rect 11006 -22826 11018 -22792
rect 11482 -22826 11494 -22792
rect 11006 -22832 11494 -22826
rect 12024 -22792 12512 -22786
rect 12024 -22826 12036 -22792
rect 12500 -22826 12512 -22792
rect 12024 -22832 12512 -22826
rect 9740 -23386 9746 -22916
rect 10714 -22920 10724 -22876
rect 9740 -23452 9754 -23386
rect 10718 -23394 10724 -22920
rect 7952 -23502 8440 -23496
rect 7952 -23536 7964 -23502
rect 8428 -23536 8440 -23502
rect 7952 -23542 8440 -23536
rect 8970 -23502 9458 -23496
rect 8970 -23536 8982 -23502
rect 9446 -23536 9458 -23502
rect 8970 -23542 9458 -23536
rect 7652 -23882 7658 -23822
rect 7718 -23882 7724 -23822
rect 8162 -24020 8222 -23542
rect 8668 -23882 8674 -23822
rect 8734 -23882 8740 -23822
rect 6934 -24026 7422 -24020
rect 6934 -24060 6946 -24026
rect 7410 -24060 7422 -24026
rect 6934 -24066 7422 -24060
rect 7952 -24026 8440 -24020
rect 7952 -24060 7964 -24026
rect 8428 -24060 8440 -24026
rect 7952 -24066 8440 -24060
rect 6638 -24160 6652 -24110
rect 5668 -24646 5674 -24164
rect 5668 -24686 5678 -24646
rect 6646 -24662 6652 -24160
rect 4898 -24736 5386 -24730
rect 4898 -24770 4910 -24736
rect 5374 -24770 5386 -24736
rect 4898 -24776 5386 -24770
rect 5112 -25034 5172 -24776
rect 5618 -24824 5678 -24686
rect 6640 -24686 6652 -24662
rect 6686 -24160 6698 -24110
rect 7664 -24110 7710 -24098
rect 6686 -24662 6692 -24160
rect 6686 -24686 6700 -24662
rect 7664 -24672 7670 -24110
rect 5916 -24736 6404 -24730
rect 5916 -24770 5928 -24736
rect 6392 -24770 6404 -24736
rect 5916 -24776 6404 -24770
rect 5612 -24884 5618 -24824
rect 5678 -24884 5684 -24824
rect 5618 -24988 5624 -24928
rect 5684 -24988 5690 -24928
rect 5106 -25094 5112 -25034
rect 5172 -25094 5178 -25034
rect 4598 -25204 4604 -25144
rect 4664 -25204 4670 -25144
rect 3880 -25258 4368 -25252
rect 3880 -25292 3892 -25258
rect 4356 -25292 4368 -25258
rect 3880 -25298 4368 -25292
rect 2614 -25918 2620 -25414
rect 3588 -25418 3598 -25342
rect 3592 -25870 3598 -25418
rect 2574 -25930 2620 -25918
rect 3584 -25918 3598 -25870
rect 3632 -25418 3648 -25342
rect 4604 -25342 4664 -25204
rect 5112 -25252 5172 -25094
rect 4898 -25258 5386 -25252
rect 4898 -25292 4910 -25258
rect 5374 -25292 5386 -25258
rect 4898 -25298 5386 -25292
rect 3632 -25870 3638 -25418
rect 3632 -25918 3644 -25870
rect 2862 -25968 3350 -25962
rect 2862 -26002 2874 -25968
rect 3338 -26002 3350 -25968
rect 2862 -26008 3350 -26002
rect 3584 -26066 3644 -25918
rect 4604 -25918 4616 -25342
rect 4650 -25918 4664 -25342
rect 5624 -25342 5684 -24988
rect 6136 -25034 6196 -24776
rect 6130 -25094 6136 -25034
rect 6196 -25094 6202 -25034
rect 6136 -25252 6196 -25094
rect 6640 -25144 6700 -24686
rect 7654 -24686 7670 -24672
rect 7704 -24672 7710 -24110
rect 8674 -24110 8734 -23882
rect 9174 -24020 9234 -23542
rect 9694 -23822 9754 -23452
rect 10706 -23452 10724 -23394
rect 10758 -22920 10774 -22876
rect 11736 -22876 11782 -22864
rect 10758 -23394 10764 -22920
rect 10758 -23452 10766 -23394
rect 11736 -23400 11742 -22876
rect 9988 -23502 10476 -23496
rect 9988 -23536 10000 -23502
rect 10464 -23536 10476 -23502
rect 9988 -23542 10476 -23536
rect 9688 -23882 9694 -23822
rect 9754 -23882 9760 -23822
rect 10204 -24020 10264 -23542
rect 10706 -23654 10766 -23452
rect 11724 -23452 11742 -23400
rect 11776 -23400 11782 -22876
rect 12742 -22876 12802 -22612
rect 13266 -22786 13326 -22510
rect 14280 -22786 14340 -22510
rect 14780 -22612 14786 -22552
rect 14846 -22612 14852 -22552
rect 13042 -22792 13530 -22786
rect 13042 -22826 13054 -22792
rect 13518 -22826 13530 -22792
rect 13042 -22832 13530 -22826
rect 14060 -22792 14548 -22786
rect 14060 -22826 14072 -22792
rect 14536 -22826 14548 -22792
rect 14060 -22832 14548 -22826
rect 12742 -22920 12760 -22876
rect 11776 -23452 11784 -23400
rect 11006 -23502 11494 -23496
rect 11006 -23536 11018 -23502
rect 11482 -23536 11494 -23502
rect 11006 -23542 11494 -23536
rect 10556 -23714 10766 -23654
rect 11220 -23708 11280 -23542
rect 11724 -23594 11784 -23452
rect 12754 -23452 12760 -22920
rect 12794 -22920 12802 -22876
rect 13772 -22876 13818 -22864
rect 12794 -23452 12800 -22920
rect 13772 -23400 13778 -22876
rect 12754 -23464 12800 -23452
rect 13766 -23452 13778 -23400
rect 13812 -23400 13818 -22876
rect 14786 -22876 14846 -22612
rect 15282 -22786 15342 -22510
rect 15078 -22792 15566 -22786
rect 15078 -22826 15090 -22792
rect 15554 -22826 15566 -22792
rect 15078 -22832 15566 -22826
rect 14786 -22924 14796 -22876
rect 13812 -23452 13826 -23400
rect 12024 -23502 12512 -23496
rect 12024 -23536 12036 -23502
rect 12500 -23536 12512 -23502
rect 12024 -23542 12512 -23536
rect 13042 -23502 13530 -23496
rect 13042 -23536 13054 -23502
rect 13518 -23536 13530 -23502
rect 13042 -23542 13530 -23536
rect 13766 -23594 13826 -23452
rect 14790 -23452 14796 -22924
rect 14830 -22924 14846 -22876
rect 15800 -22876 15860 -22502
rect 16308 -22786 16368 -22410
rect 16808 -22612 16814 -22552
rect 16874 -22612 16880 -22552
rect 16096 -22792 16584 -22786
rect 16096 -22826 16108 -22792
rect 16572 -22826 16584 -22792
rect 16096 -22832 16584 -22826
rect 15800 -22912 15814 -22876
rect 14830 -23452 14836 -22924
rect 15808 -23408 15814 -22912
rect 14790 -23464 14836 -23452
rect 15802 -23452 15814 -23408
rect 15848 -22912 15860 -22876
rect 16814 -22876 16874 -22612
rect 17328 -22786 17388 -22310
rect 17840 -22678 17900 -22220
rect 18852 -22220 18868 -22176
rect 18902 -22176 18908 -21644
rect 19872 -21644 19932 -21500
rect 20364 -21554 20424 -21388
rect 20168 -21560 20656 -21554
rect 20168 -21594 20180 -21560
rect 20644 -21594 20656 -21560
rect 20168 -21600 20656 -21594
rect 19872 -21702 19886 -21644
rect 18902 -22220 18912 -22176
rect 19880 -22180 19886 -21702
rect 18132 -22270 18620 -22264
rect 18132 -22304 18144 -22270
rect 18608 -22304 18620 -22270
rect 18132 -22310 18620 -22304
rect 17834 -22738 17840 -22678
rect 17900 -22738 17906 -22678
rect 17114 -22792 17602 -22786
rect 17114 -22826 17126 -22792
rect 17590 -22826 17602 -22792
rect 17114 -22832 17602 -22826
rect 15848 -23408 15854 -22912
rect 16814 -22924 16832 -22876
rect 15848 -23452 15862 -23408
rect 16826 -23412 16832 -22924
rect 14060 -23502 14548 -23496
rect 14060 -23536 14072 -23502
rect 14536 -23536 14548 -23502
rect 14060 -23542 14548 -23536
rect 15078 -23502 15566 -23496
rect 15078 -23536 15090 -23502
rect 15554 -23536 15566 -23502
rect 15078 -23542 15566 -23536
rect 15802 -23594 15862 -23452
rect 16816 -23452 16832 -23412
rect 16866 -22924 16874 -22876
rect 17840 -22876 17900 -22738
rect 18344 -22786 18404 -22310
rect 18852 -22552 18912 -22220
rect 19870 -22220 19886 -22180
rect 19920 -21702 19932 -21644
rect 20892 -21644 20952 -20986
rect 21908 -20986 21922 -20942
rect 21956 -20444 21972 -20410
rect 22934 -20410 22980 -20398
rect 21956 -20942 21962 -20444
rect 21956 -20986 21968 -20942
rect 22934 -20956 22940 -20410
rect 21186 -21036 21674 -21030
rect 21186 -21070 21198 -21036
rect 21662 -21070 21674 -21036
rect 21186 -21076 21674 -21070
rect 21394 -21328 21454 -21076
rect 21908 -21168 21968 -20986
rect 22924 -20986 22940 -20956
rect 22974 -20956 22980 -20410
rect 22974 -20986 22984 -20956
rect 22204 -21036 22692 -21030
rect 22204 -21070 22216 -21036
rect 22680 -21070 22692 -21036
rect 22204 -21076 22692 -21070
rect 22414 -21168 22474 -21076
rect 22924 -21168 22984 -20986
rect 21908 -21228 22984 -21168
rect 21388 -21388 21394 -21328
rect 21454 -21388 21460 -21328
rect 21908 -21440 21968 -21228
rect 21902 -21500 21908 -21440
rect 21968 -21500 21974 -21440
rect 21186 -21560 21674 -21554
rect 21186 -21594 21198 -21560
rect 21662 -21594 21674 -21560
rect 21186 -21600 21674 -21594
rect 22204 -21560 22692 -21554
rect 22204 -21594 22216 -21560
rect 22680 -21594 22692 -21560
rect 22204 -21600 22692 -21594
rect 20892 -21686 20904 -21644
rect 19920 -22180 19926 -21702
rect 20898 -22166 20904 -21686
rect 19920 -22220 19930 -22180
rect 19150 -22270 19638 -22264
rect 19150 -22304 19162 -22270
rect 19626 -22304 19638 -22270
rect 19150 -22310 19638 -22304
rect 18846 -22612 18852 -22552
rect 18912 -22612 18918 -22552
rect 19378 -22786 19438 -22310
rect 19870 -22678 19930 -22220
rect 20892 -22220 20904 -22166
rect 20938 -21686 20952 -21644
rect 21916 -21644 21962 -21632
rect 20938 -22166 20944 -21686
rect 20938 -22220 20952 -22166
rect 21916 -22174 21922 -21644
rect 20168 -22270 20656 -22264
rect 20168 -22304 20180 -22270
rect 20644 -22304 20656 -22270
rect 20168 -22310 20656 -22304
rect 20396 -22676 20456 -22310
rect 20892 -22552 20952 -22220
rect 21906 -22220 21922 -22174
rect 21956 -22174 21962 -21644
rect 22934 -21644 22980 -21632
rect 21956 -22220 21966 -22174
rect 22934 -22192 22940 -21644
rect 21186 -22270 21674 -22264
rect 21186 -22304 21198 -22270
rect 21662 -22304 21674 -22270
rect 21186 -22310 21674 -22304
rect 21410 -22548 21470 -22310
rect 21906 -22346 21966 -22220
rect 22926 -22220 22940 -22192
rect 22974 -22192 22980 -21644
rect 22974 -22220 22986 -22192
rect 22204 -22270 22692 -22264
rect 22204 -22304 22216 -22270
rect 22680 -22304 22692 -22270
rect 22204 -22310 22692 -22304
rect 22412 -22344 22472 -22310
rect 22926 -22344 22986 -22220
rect 22412 -22346 22986 -22344
rect 21906 -22406 22986 -22346
rect 21906 -22442 21966 -22406
rect 21900 -22502 21906 -22442
rect 21966 -22502 21972 -22442
rect 20886 -22612 20892 -22552
rect 20952 -22612 20958 -22552
rect 21404 -22608 21410 -22548
rect 21470 -22608 21476 -22548
rect 22916 -22608 22922 -22548
rect 22982 -22608 22988 -22548
rect 19864 -22738 19870 -22678
rect 19930 -22738 19936 -22678
rect 18132 -22792 18620 -22786
rect 18132 -22826 18144 -22792
rect 18608 -22826 18620 -22792
rect 18132 -22832 18620 -22826
rect 19150 -22792 19638 -22786
rect 19150 -22826 19162 -22792
rect 19626 -22826 19638 -22792
rect 19150 -22832 19638 -22826
rect 17840 -22922 17850 -22876
rect 16866 -23412 16872 -22924
rect 17844 -23392 17850 -22922
rect 16866 -23452 16876 -23412
rect 16096 -23502 16584 -23496
rect 16096 -23536 16108 -23502
rect 16572 -23536 16584 -23502
rect 16096 -23542 16584 -23536
rect 11718 -23654 11724 -23594
rect 11784 -23654 11790 -23594
rect 13760 -23654 13766 -23594
rect 13826 -23654 13832 -23594
rect 15796 -23654 15802 -23594
rect 15862 -23654 15868 -23594
rect 16308 -23704 16368 -23542
rect 16816 -23602 16876 -23452
rect 17838 -23452 17850 -23392
rect 17884 -22922 17900 -22876
rect 18862 -22876 18908 -22864
rect 17884 -23392 17890 -22922
rect 17884 -23452 17898 -23392
rect 18862 -23408 18868 -22876
rect 17114 -23502 17602 -23496
rect 17114 -23536 17126 -23502
rect 17590 -23536 17602 -23502
rect 17114 -23542 17602 -23536
rect 16816 -23662 17022 -23602
rect 10556 -23926 10616 -23714
rect 11214 -23768 11220 -23708
rect 11280 -23768 11286 -23708
rect 16302 -23764 16308 -23704
rect 16368 -23764 16374 -23704
rect 10706 -23882 10712 -23822
rect 10772 -23882 10778 -23822
rect 12736 -23882 12742 -23822
rect 12802 -23882 12808 -23822
rect 14774 -23882 14780 -23822
rect 14840 -23882 14846 -23822
rect 16810 -23882 16816 -23822
rect 16876 -23882 16882 -23822
rect 10550 -23986 10556 -23926
rect 10616 -23986 10622 -23926
rect 8970 -24026 9458 -24020
rect 8970 -24060 8982 -24026
rect 9446 -24060 9458 -24026
rect 8970 -24066 9458 -24060
rect 9988 -24026 10476 -24020
rect 9988 -24060 10000 -24026
rect 10464 -24060 10476 -24026
rect 9988 -24066 10476 -24060
rect 8674 -24592 8688 -24110
rect 8682 -24666 8688 -24592
rect 7704 -24686 7714 -24672
rect 6934 -24736 7422 -24730
rect 6934 -24770 6946 -24736
rect 7410 -24770 7422 -24736
rect 6934 -24776 7422 -24770
rect 7154 -25034 7214 -24776
rect 7654 -24928 7714 -24686
rect 8678 -24686 8688 -24666
rect 8722 -24592 8734 -24110
rect 9700 -24110 9746 -24098
rect 8722 -24666 8728 -24592
rect 9700 -24660 9706 -24110
rect 8722 -24686 8738 -24666
rect 7952 -24736 8440 -24730
rect 7952 -24770 7964 -24736
rect 8428 -24770 8440 -24736
rect 7952 -24776 8440 -24770
rect 7648 -24988 7654 -24928
rect 7714 -24988 7720 -24928
rect 8168 -25034 8228 -24776
rect 7148 -25094 7154 -25034
rect 7214 -25094 7220 -25034
rect 8162 -25094 8168 -25034
rect 8228 -25094 8234 -25034
rect 6634 -25204 6640 -25144
rect 6700 -25204 6706 -25144
rect 5916 -25258 6404 -25252
rect 5916 -25292 5928 -25258
rect 6392 -25292 6404 -25258
rect 5916 -25298 6404 -25292
rect 5624 -25356 5634 -25342
rect 3880 -25968 4368 -25962
rect 3880 -26002 3892 -25968
rect 4356 -26002 4368 -25968
rect 3880 -26008 4368 -26002
rect 2442 -26126 2448 -26066
rect 2508 -26126 2514 -26066
rect 3578 -26126 3584 -26066
rect 3644 -26126 3650 -26066
rect 4096 -26174 4156 -26008
rect 4090 -26234 4096 -26174
rect 4156 -26234 4162 -26174
rect 4604 -26430 4664 -25918
rect 5628 -25918 5634 -25356
rect 5668 -25356 5684 -25342
rect 6640 -25342 6700 -25204
rect 7154 -25252 7214 -25094
rect 8168 -25252 8228 -25094
rect 8678 -25144 8738 -24686
rect 9694 -24686 9706 -24660
rect 9740 -24660 9746 -24110
rect 10712 -24110 10772 -23882
rect 11006 -24026 11494 -24020
rect 11006 -24060 11018 -24026
rect 11482 -24060 11494 -24026
rect 11006 -24066 11494 -24060
rect 12024 -24026 12512 -24020
rect 12024 -24060 12036 -24026
rect 12500 -24060 12512 -24026
rect 12024 -24066 12512 -24060
rect 11736 -24110 11782 -24098
rect 12742 -24110 12802 -23882
rect 13042 -24026 13530 -24020
rect 13042 -24060 13054 -24026
rect 13518 -24060 13530 -24026
rect 13042 -24066 13530 -24060
rect 14060 -24026 14548 -24020
rect 14060 -24060 14072 -24026
rect 14536 -24060 14548 -24026
rect 14060 -24066 14548 -24060
rect 13772 -24110 13818 -24098
rect 14780 -24110 14840 -23882
rect 15078 -24026 15566 -24020
rect 15078 -24060 15090 -24026
rect 15554 -24060 15566 -24026
rect 15078 -24066 15566 -24060
rect 16096 -24026 16584 -24020
rect 16096 -24060 16108 -24026
rect 16572 -24060 16584 -24026
rect 16096 -24066 16584 -24060
rect 10712 -24166 10724 -24110
rect 9740 -24686 9754 -24660
rect 10718 -24662 10724 -24166
rect 8970 -24736 9458 -24730
rect 8970 -24770 8982 -24736
rect 9446 -24770 9458 -24736
rect 8970 -24776 9458 -24770
rect 9200 -25034 9260 -24776
rect 9694 -24928 9754 -24686
rect 10716 -24686 10724 -24662
rect 10758 -24166 10772 -24110
rect 11730 -24146 11742 -24110
rect 10758 -24662 10764 -24166
rect 11736 -24634 11742 -24146
rect 10758 -24686 10776 -24662
rect 9988 -24736 10476 -24730
rect 9988 -24770 10000 -24736
rect 10464 -24770 10476 -24736
rect 9988 -24776 10476 -24770
rect 9842 -24882 9848 -24822
rect 9908 -24882 9914 -24822
rect 9688 -24988 9694 -24928
rect 9754 -24988 9760 -24928
rect 9194 -25094 9200 -25034
rect 9260 -25094 9266 -25034
rect 9848 -25066 9908 -24882
rect 10212 -25034 10272 -24776
rect 8672 -25204 8678 -25144
rect 8738 -25204 8744 -25144
rect 6934 -25258 7422 -25252
rect 6934 -25292 6946 -25258
rect 7410 -25292 7422 -25258
rect 6934 -25298 7422 -25292
rect 7952 -25258 8440 -25252
rect 7952 -25292 7964 -25258
rect 8428 -25292 8440 -25258
rect 7952 -25298 8440 -25292
rect 5668 -25918 5674 -25356
rect 5628 -25930 5674 -25918
rect 6640 -25918 6652 -25342
rect 6686 -25918 6700 -25342
rect 7664 -25342 7710 -25330
rect 7664 -25876 7670 -25342
rect 4898 -25968 5386 -25962
rect 4898 -26002 4910 -25968
rect 5374 -26002 5386 -25968
rect 4898 -26008 5386 -26002
rect 5916 -25968 6404 -25962
rect 5916 -26002 5928 -25968
rect 6392 -26002 6404 -25968
rect 5916 -26008 6404 -26002
rect 5110 -26174 5170 -26008
rect 5110 -26240 5170 -26234
rect 6132 -26174 6192 -26008
rect 6132 -26240 6192 -26234
rect 6640 -26430 6700 -25918
rect 7654 -25918 7670 -25876
rect 7704 -25876 7710 -25342
rect 8678 -25342 8738 -25204
rect 9200 -25252 9260 -25094
rect 9692 -25126 9908 -25066
rect 10206 -25094 10212 -25034
rect 10272 -25094 10278 -25034
rect 8970 -25258 9458 -25252
rect 8970 -25292 8982 -25258
rect 9446 -25292 9458 -25258
rect 8970 -25298 9458 -25292
rect 7704 -25918 7714 -25876
rect 6934 -25968 7422 -25962
rect 6934 -26002 6946 -25968
rect 7410 -26002 7422 -25968
rect 6934 -26008 7422 -26002
rect 7144 -26168 7204 -26008
rect 7654 -26066 7714 -25918
rect 8678 -25918 8688 -25342
rect 8722 -25918 8738 -25342
rect 9692 -25342 9752 -25126
rect 10212 -25252 10272 -25094
rect 10716 -25144 10776 -24686
rect 11726 -24686 11742 -24634
rect 11776 -24146 11790 -24110
rect 11776 -24634 11782 -24146
rect 12742 -24160 12760 -24110
rect 11776 -24686 11786 -24634
rect 12754 -24656 12760 -24160
rect 11006 -24736 11494 -24730
rect 11006 -24770 11018 -24736
rect 11482 -24770 11494 -24736
rect 11006 -24776 11494 -24770
rect 11220 -25034 11280 -24776
rect 11726 -24822 11786 -24686
rect 12752 -24686 12760 -24656
rect 12794 -24160 12802 -24110
rect 13766 -24142 13778 -24110
rect 12794 -24656 12800 -24160
rect 13772 -24646 13778 -24142
rect 12794 -24686 12812 -24656
rect 12024 -24736 12512 -24730
rect 12024 -24770 12036 -24736
rect 12500 -24770 12512 -24736
rect 12024 -24776 12512 -24770
rect 11720 -24882 11726 -24822
rect 11786 -24882 11792 -24822
rect 11724 -24988 11730 -24928
rect 11790 -24988 11796 -24928
rect 11214 -25094 11220 -25034
rect 11280 -25094 11286 -25034
rect 10710 -25204 10716 -25144
rect 10776 -25204 10782 -25144
rect 9988 -25258 10476 -25252
rect 9988 -25292 10000 -25258
rect 10464 -25292 10476 -25258
rect 9988 -25298 10476 -25292
rect 9692 -25368 9706 -25342
rect 7952 -25968 8440 -25962
rect 7952 -26002 7964 -25968
rect 8428 -26002 8440 -25968
rect 7952 -26008 8440 -26002
rect 7648 -26126 7654 -26066
rect 7714 -26126 7720 -26066
rect 8170 -26168 8230 -26008
rect 7144 -26174 7206 -26168
rect 7144 -26180 7146 -26174
rect 8170 -26174 8232 -26168
rect 8170 -26180 8172 -26174
rect 7146 -26240 7206 -26234
rect 8172 -26240 8232 -26234
rect 8678 -26430 8738 -25918
rect 9700 -25918 9706 -25368
rect 9740 -25368 9752 -25342
rect 10716 -25342 10776 -25204
rect 11220 -25252 11280 -25094
rect 11006 -25258 11494 -25252
rect 11006 -25292 11018 -25258
rect 11482 -25292 11494 -25258
rect 11006 -25298 11494 -25292
rect 9740 -25918 9746 -25368
rect 9700 -25930 9746 -25918
rect 10716 -25918 10724 -25342
rect 10758 -25918 10776 -25342
rect 11730 -25342 11790 -24988
rect 12238 -25034 12298 -24776
rect 12232 -25094 12238 -25034
rect 12298 -25094 12304 -25034
rect 12238 -25252 12298 -25094
rect 12752 -25144 12812 -24686
rect 13764 -24686 13778 -24646
rect 13812 -24142 13826 -24110
rect 13812 -24646 13818 -24142
rect 14780 -24154 14796 -24110
rect 13812 -24686 13824 -24646
rect 14790 -24662 14796 -24154
rect 13042 -24736 13530 -24730
rect 13042 -24770 13054 -24736
rect 13518 -24770 13530 -24736
rect 13042 -24776 13530 -24770
rect 13264 -25034 13324 -24776
rect 13764 -24822 13824 -24686
rect 14788 -24686 14796 -24662
rect 14830 -24154 14840 -24110
rect 15808 -24110 15854 -24098
rect 14830 -24662 14836 -24154
rect 15808 -24640 15814 -24110
rect 14830 -24686 14848 -24662
rect 14060 -24736 14548 -24730
rect 14060 -24770 14072 -24736
rect 14536 -24770 14548 -24736
rect 14060 -24776 14548 -24770
rect 13758 -24882 13764 -24822
rect 13824 -24882 13830 -24822
rect 13760 -24988 13766 -24928
rect 13826 -24988 13832 -24928
rect 13258 -25094 13264 -25034
rect 13324 -25094 13330 -25034
rect 12746 -25204 12752 -25144
rect 12812 -25204 12818 -25144
rect 12024 -25258 12512 -25252
rect 12024 -25292 12036 -25258
rect 12500 -25292 12512 -25258
rect 12024 -25298 12512 -25292
rect 11730 -25368 11742 -25342
rect 8970 -25968 9458 -25962
rect 8970 -26002 8982 -25968
rect 9446 -26002 9458 -25968
rect 8970 -26008 9458 -26002
rect 9988 -25968 10476 -25962
rect 9988 -26002 10000 -25968
rect 10464 -26002 10476 -25968
rect 9988 -26008 10476 -26002
rect 9184 -26174 9244 -26008
rect 9184 -26240 9244 -26234
rect 10220 -26174 10280 -26008
rect 10220 -26240 10280 -26234
rect 10716 -26430 10776 -25918
rect 11736 -25918 11742 -25368
rect 11776 -25368 11790 -25342
rect 12752 -25342 12812 -25204
rect 13264 -25252 13324 -25094
rect 13042 -25258 13530 -25252
rect 13042 -25292 13054 -25258
rect 13518 -25292 13530 -25258
rect 13042 -25298 13530 -25292
rect 11776 -25918 11782 -25368
rect 11736 -25930 11782 -25918
rect 12752 -25918 12760 -25342
rect 12794 -25918 12812 -25342
rect 13766 -25342 13826 -24988
rect 14266 -25034 14326 -24776
rect 14260 -25094 14266 -25034
rect 14326 -25094 14332 -25034
rect 14266 -25252 14326 -25094
rect 14788 -25144 14848 -24686
rect 15800 -24686 15814 -24640
rect 15848 -24640 15854 -24110
rect 16816 -24110 16876 -23882
rect 16962 -23926 17022 -23662
rect 16956 -23986 16962 -23926
rect 17022 -23986 17028 -23926
rect 17326 -24020 17386 -23542
rect 17838 -23822 17898 -23452
rect 18856 -23452 18868 -23408
rect 18902 -23408 18908 -22876
rect 19870 -22876 19930 -22738
rect 20396 -22786 20456 -22736
rect 21410 -22786 21470 -22608
rect 21904 -22736 21910 -22676
rect 21970 -22736 21976 -22676
rect 20168 -22792 20656 -22786
rect 20168 -22826 20180 -22792
rect 20644 -22826 20656 -22792
rect 20168 -22832 20656 -22826
rect 21186 -22792 21674 -22786
rect 21186 -22826 21198 -22792
rect 21662 -22826 21674 -22792
rect 21186 -22832 21674 -22826
rect 19870 -22922 19886 -22876
rect 19880 -23404 19886 -22922
rect 18902 -23452 18916 -23408
rect 18132 -23502 18620 -23496
rect 18132 -23536 18144 -23502
rect 18608 -23536 18620 -23502
rect 18132 -23542 18620 -23536
rect 17832 -23882 17838 -23822
rect 17898 -23882 17904 -23822
rect 18346 -24020 18406 -23542
rect 18856 -23594 18916 -23452
rect 19872 -23452 19886 -23404
rect 19920 -22922 19930 -22876
rect 20898 -22876 20944 -22864
rect 21910 -22876 21970 -22736
rect 22204 -22792 22692 -22786
rect 22204 -22826 22216 -22792
rect 22680 -22826 22692 -22792
rect 22204 -22832 22692 -22826
rect 19920 -23404 19926 -22922
rect 19920 -23452 19932 -23404
rect 20898 -23408 20904 -22876
rect 19150 -23502 19638 -23496
rect 19150 -23536 19162 -23502
rect 19626 -23536 19638 -23502
rect 19150 -23542 19638 -23536
rect 18850 -23654 18856 -23594
rect 18916 -23654 18922 -23594
rect 18852 -23882 18858 -23822
rect 18918 -23882 18924 -23822
rect 17114 -24026 17602 -24020
rect 17114 -24060 17126 -24026
rect 17590 -24060 17602 -24026
rect 17114 -24066 17602 -24060
rect 18132 -24026 18620 -24020
rect 18132 -24060 18144 -24026
rect 18608 -24060 18620 -24026
rect 18132 -24066 18620 -24060
rect 16816 -24154 16832 -24110
rect 15848 -24686 15860 -24640
rect 16826 -24660 16832 -24154
rect 15078 -24736 15566 -24730
rect 15078 -24770 15090 -24736
rect 15554 -24770 15566 -24736
rect 15078 -24776 15566 -24770
rect 15286 -25034 15346 -24776
rect 15628 -24882 15634 -24822
rect 15694 -24882 15700 -24822
rect 15280 -25094 15286 -25034
rect 15346 -25094 15352 -25034
rect 15634 -25074 15694 -24882
rect 15800 -24928 15860 -24686
rect 16820 -24686 16832 -24660
rect 16866 -24154 16876 -24110
rect 17844 -24110 17890 -24098
rect 16866 -24660 16872 -24154
rect 17844 -24646 17850 -24110
rect 16866 -24686 16880 -24660
rect 16096 -24736 16584 -24730
rect 16096 -24770 16108 -24736
rect 16572 -24770 16584 -24736
rect 16096 -24776 16584 -24770
rect 15794 -24988 15800 -24928
rect 15860 -24988 15866 -24928
rect 16306 -25034 16366 -24776
rect 14782 -25204 14788 -25144
rect 14848 -25204 14854 -25144
rect 14060 -25258 14548 -25252
rect 14060 -25292 14072 -25258
rect 14536 -25292 14548 -25258
rect 14060 -25298 14548 -25292
rect 13766 -25378 13778 -25342
rect 11006 -25968 11494 -25962
rect 11006 -26002 11018 -25968
rect 11482 -26002 11494 -25968
rect 11006 -26008 11494 -26002
rect 12024 -25968 12512 -25962
rect 12024 -26002 12036 -25968
rect 12500 -26002 12512 -25968
rect 12024 -26008 12512 -26002
rect 11226 -26174 11286 -26008
rect 12240 -26174 12300 -26008
rect 12234 -26234 12240 -26174
rect 12300 -26234 12306 -26174
rect 11226 -26240 11286 -26234
rect 12752 -26430 12812 -25918
rect 13772 -25918 13778 -25378
rect 13812 -25378 13826 -25342
rect 14788 -25342 14848 -25204
rect 15286 -25252 15346 -25094
rect 15634 -25134 15860 -25074
rect 16300 -25094 16306 -25034
rect 16366 -25094 16372 -25034
rect 15078 -25258 15566 -25252
rect 15078 -25292 15090 -25258
rect 15554 -25292 15566 -25258
rect 15078 -25298 15566 -25292
rect 13812 -25918 13818 -25378
rect 13772 -25930 13818 -25918
rect 14788 -25918 14796 -25342
rect 14830 -25918 14848 -25342
rect 15800 -25342 15860 -25134
rect 16306 -25252 16366 -25094
rect 16820 -25144 16880 -24686
rect 17840 -24686 17850 -24646
rect 17884 -24646 17890 -24110
rect 18858 -24110 18918 -23882
rect 19360 -24020 19420 -23542
rect 19872 -23822 19932 -23452
rect 20888 -23452 20904 -23408
rect 20938 -23408 20944 -22876
rect 21908 -22910 21922 -22876
rect 21910 -22920 21922 -22910
rect 20938 -23452 20948 -23408
rect 20168 -23502 20656 -23496
rect 20168 -23536 20180 -23502
rect 20644 -23536 20656 -23502
rect 20168 -23542 20656 -23536
rect 19866 -23882 19872 -23822
rect 19932 -23882 19938 -23822
rect 19866 -23986 19872 -23926
rect 19932 -23986 19938 -23926
rect 19150 -24026 19638 -24020
rect 19150 -24060 19162 -24026
rect 19626 -24060 19638 -24026
rect 19150 -24066 19638 -24060
rect 19368 -24070 19428 -24066
rect 18858 -24176 18868 -24110
rect 18862 -24640 18868 -24176
rect 17884 -24686 17900 -24646
rect 17114 -24736 17602 -24730
rect 17114 -24770 17126 -24736
rect 17590 -24770 17602 -24736
rect 17114 -24776 17602 -24770
rect 17332 -25034 17392 -24776
rect 17840 -24928 17900 -24686
rect 18852 -24686 18868 -24640
rect 18902 -24176 18918 -24110
rect 19872 -24110 19932 -23986
rect 20396 -24020 20456 -23542
rect 20888 -23594 20948 -23452
rect 21916 -23452 21922 -22920
rect 21956 -22920 21970 -22876
rect 22922 -22876 22982 -22608
rect 21956 -23452 21962 -22920
rect 22922 -22930 22940 -22876
rect 21916 -23464 21962 -23452
rect 22934 -23452 22940 -22930
rect 22974 -22914 22986 -22876
rect 22974 -22930 22982 -22914
rect 22974 -23452 22980 -22930
rect 22934 -23464 22980 -23452
rect 21186 -23502 21674 -23496
rect 21186 -23536 21198 -23502
rect 21662 -23536 21674 -23502
rect 21186 -23542 21674 -23536
rect 22204 -23502 22692 -23496
rect 22204 -23536 22216 -23502
rect 22680 -23536 22692 -23502
rect 22204 -23542 22692 -23536
rect 20882 -23654 20888 -23594
rect 20948 -23654 20954 -23594
rect 21408 -23704 21468 -23542
rect 22416 -23704 22476 -23542
rect 23034 -23594 23094 -17804
rect 23156 -18718 23162 -18658
rect 23222 -18718 23228 -18658
rect 23162 -20216 23222 -18718
rect 23278 -18982 23338 -17690
rect 23394 -18940 23400 -18880
rect 23460 -18940 23466 -18880
rect 23272 -19042 23278 -18982
rect 23338 -19042 23344 -18982
rect 23156 -20276 23162 -20216
rect 23222 -20276 23228 -20216
rect 23152 -21178 23158 -21118
rect 23218 -21178 23224 -21118
rect 23158 -22442 23218 -21178
rect 23278 -22344 23338 -19042
rect 23272 -22404 23278 -22344
rect 23338 -22404 23344 -22344
rect 23152 -22502 23158 -22442
rect 23218 -22502 23224 -22442
rect 23028 -23654 23034 -23594
rect 23094 -23654 23100 -23594
rect 21402 -23764 21408 -23704
rect 21468 -23764 21474 -23704
rect 22410 -23764 22416 -23704
rect 22476 -23764 22482 -23704
rect 23278 -23820 23338 -22404
rect 23400 -22676 23460 -18940
rect 23528 -20108 23588 -17586
rect 23526 -20114 23588 -20108
rect 23586 -20174 23588 -20114
rect 23526 -20180 23588 -20174
rect 23528 -22548 23588 -20180
rect 23522 -22608 23528 -22548
rect 23588 -22608 23594 -22548
rect 23394 -22736 23400 -22676
rect 23460 -22736 23466 -22676
rect 23650 -23704 23710 -12776
rect 23756 -16586 23762 -16526
rect 23822 -16586 23828 -16526
rect 23644 -23764 23650 -23704
rect 23710 -23764 23716 -23704
rect 20888 -23882 20894 -23822
rect 20954 -23882 20960 -23822
rect 21910 -23880 23338 -23820
rect 20168 -24026 20656 -24020
rect 20168 -24060 20180 -24026
rect 20644 -24060 20656 -24026
rect 20168 -24066 20656 -24060
rect 19872 -24156 19886 -24110
rect 18902 -24640 18908 -24176
rect 18902 -24686 18912 -24640
rect 18132 -24736 18620 -24730
rect 18132 -24770 18144 -24736
rect 18608 -24770 18620 -24736
rect 18132 -24776 18620 -24770
rect 17834 -24988 17840 -24928
rect 17900 -24988 17906 -24928
rect 18350 -25034 18410 -24776
rect 17326 -25094 17332 -25034
rect 17392 -25094 17398 -25034
rect 18344 -25094 18350 -25034
rect 18410 -25094 18416 -25034
rect 16814 -25204 16820 -25144
rect 16880 -25204 16886 -25144
rect 16096 -25258 16584 -25252
rect 16096 -25292 16108 -25258
rect 16572 -25292 16584 -25258
rect 16096 -25298 16584 -25292
rect 15800 -25378 15814 -25342
rect 13042 -25968 13530 -25962
rect 13042 -26002 13054 -25968
rect 13518 -26002 13530 -25968
rect 13042 -26008 13530 -26002
rect 14060 -25968 14548 -25962
rect 14060 -26002 14072 -25968
rect 14536 -26002 14548 -25968
rect 14060 -26008 14548 -26002
rect 13256 -26174 13316 -26008
rect 14266 -26168 14326 -26008
rect 13256 -26240 13316 -26234
rect 14264 -26174 14326 -26168
rect 14324 -26180 14326 -26174
rect 14264 -26240 14324 -26234
rect 14788 -26430 14848 -25918
rect 15808 -25918 15814 -25378
rect 15848 -25378 15860 -25342
rect 16820 -25342 16880 -25204
rect 17332 -25252 17392 -25094
rect 18350 -25252 18410 -25094
rect 18852 -25144 18912 -24686
rect 19880 -24686 19886 -24156
rect 19920 -24156 19932 -24110
rect 20894 -24110 20954 -23882
rect 21186 -24026 21674 -24020
rect 21186 -24060 21198 -24026
rect 21662 -24060 21674 -24026
rect 21186 -24066 21674 -24060
rect 19920 -24686 19926 -24156
rect 20894 -24170 20904 -24110
rect 20898 -24662 20904 -24170
rect 19880 -24698 19926 -24686
rect 20892 -24686 20904 -24662
rect 20938 -24170 20954 -24110
rect 21910 -24110 21970 -23880
rect 22408 -24020 22468 -23880
rect 22204 -24026 22692 -24020
rect 22204 -24060 22216 -24026
rect 22680 -24060 22692 -24026
rect 22204 -24066 22692 -24060
rect 20938 -24662 20944 -24170
rect 20938 -24686 20952 -24662
rect 19150 -24736 19638 -24730
rect 19150 -24770 19162 -24736
rect 19626 -24770 19638 -24736
rect 19150 -24776 19638 -24770
rect 20168 -24736 20656 -24730
rect 20168 -24770 20180 -24736
rect 20644 -24770 20656 -24736
rect 20168 -24776 20656 -24770
rect 19364 -25034 19424 -24776
rect 19864 -24988 19870 -24928
rect 19930 -24988 19936 -24928
rect 19358 -25094 19364 -25034
rect 19424 -25094 19430 -25034
rect 18846 -25204 18852 -25144
rect 18912 -25204 18918 -25144
rect 17114 -25258 17602 -25252
rect 17114 -25292 17126 -25258
rect 17590 -25292 17602 -25258
rect 17114 -25298 17602 -25292
rect 18132 -25258 18620 -25252
rect 18132 -25292 18144 -25258
rect 18608 -25292 18620 -25258
rect 18132 -25298 18620 -25292
rect 15848 -25918 15854 -25378
rect 15808 -25930 15854 -25918
rect 16820 -25918 16832 -25342
rect 16866 -25918 16880 -25342
rect 17844 -25342 17890 -25330
rect 17844 -25866 17850 -25342
rect 16304 -25962 16364 -25960
rect 15078 -25968 15566 -25962
rect 15078 -26002 15090 -25968
rect 15554 -26002 15566 -25968
rect 15078 -26008 15566 -26002
rect 16096 -25968 16584 -25962
rect 16096 -26002 16108 -25968
rect 16572 -26002 16584 -25968
rect 16096 -26008 16584 -26002
rect 15282 -26168 15342 -26008
rect 15280 -26174 15342 -26168
rect 15340 -26180 15342 -26174
rect 16304 -26174 16364 -26008
rect 15280 -26240 15340 -26234
rect 16304 -26240 16364 -26234
rect 16820 -26430 16880 -25918
rect 17834 -25918 17850 -25866
rect 17884 -25866 17890 -25342
rect 18852 -25342 18912 -25204
rect 19364 -25252 19424 -25094
rect 19150 -25258 19638 -25252
rect 19150 -25292 19162 -25258
rect 19626 -25292 19638 -25258
rect 19150 -25298 19638 -25292
rect 17884 -25918 17894 -25866
rect 17114 -25968 17602 -25962
rect 17114 -26002 17126 -25968
rect 17590 -26002 17602 -25968
rect 17114 -26008 17602 -26002
rect 17326 -26174 17386 -26008
rect 17834 -26066 17894 -25918
rect 18852 -25918 18868 -25342
rect 18902 -25918 18912 -25342
rect 19870 -25342 19930 -24988
rect 20378 -25034 20438 -24776
rect 20372 -25094 20378 -25034
rect 20438 -25094 20444 -25034
rect 20378 -25252 20438 -25094
rect 20892 -25144 20952 -24686
rect 21910 -24686 21922 -24110
rect 21956 -24686 21970 -24110
rect 22924 -24110 22984 -23880
rect 23048 -23986 23054 -23926
rect 23114 -23986 23120 -23926
rect 22924 -24164 22940 -24110
rect 21186 -24736 21674 -24730
rect 21186 -24770 21198 -24736
rect 21662 -24770 21674 -24736
rect 21186 -24776 21674 -24770
rect 21400 -25034 21460 -24776
rect 21910 -24822 21970 -24686
rect 22934 -24686 22940 -24164
rect 22974 -24164 22984 -24110
rect 22974 -24686 22980 -24164
rect 22934 -24698 22980 -24686
rect 22204 -24736 22692 -24730
rect 22204 -24770 22216 -24736
rect 22680 -24770 22692 -24736
rect 22204 -24776 22692 -24770
rect 21904 -24882 21910 -24822
rect 21970 -24882 21976 -24822
rect 21904 -24988 21910 -24928
rect 21970 -24988 21976 -24928
rect 21394 -25094 21400 -25034
rect 21460 -25094 21466 -25034
rect 20886 -25204 20892 -25144
rect 20952 -25204 20958 -25144
rect 20168 -25258 20656 -25252
rect 20168 -25292 20180 -25258
rect 20644 -25292 20656 -25258
rect 20168 -25298 20656 -25292
rect 19870 -25386 19886 -25342
rect 18132 -25968 18620 -25962
rect 18132 -26002 18144 -25968
rect 18608 -26002 18620 -25968
rect 18132 -26008 18620 -26002
rect 17828 -26126 17834 -26066
rect 17894 -26126 17900 -26066
rect 18346 -26168 18406 -26008
rect 18346 -26174 18408 -26168
rect 18346 -26180 18348 -26174
rect 17326 -26240 17386 -26234
rect 18348 -26240 18408 -26234
rect 18852 -26430 18912 -25918
rect 19880 -25918 19886 -25386
rect 19920 -25386 19930 -25342
rect 20892 -25342 20952 -25204
rect 21400 -25252 21460 -25094
rect 21910 -25144 21970 -24988
rect 21910 -25204 22988 -25144
rect 21186 -25258 21674 -25252
rect 21186 -25292 21198 -25258
rect 21662 -25292 21674 -25258
rect 21186 -25298 21674 -25292
rect 19920 -25918 19926 -25386
rect 19880 -25930 19926 -25918
rect 20892 -25918 20904 -25342
rect 20938 -25918 20952 -25342
rect 21910 -25342 21970 -25204
rect 22426 -25252 22486 -25204
rect 22204 -25258 22692 -25252
rect 22204 -25292 22216 -25258
rect 22680 -25292 22692 -25258
rect 22204 -25298 22692 -25292
rect 21910 -25350 21922 -25342
rect 19368 -25962 19428 -25960
rect 19150 -25968 19638 -25962
rect 19150 -26002 19162 -25968
rect 19626 -26002 19638 -25968
rect 19150 -26008 19638 -26002
rect 20168 -25968 20656 -25962
rect 20168 -26002 20180 -25968
rect 20644 -26002 20656 -25968
rect 20168 -26008 20656 -26002
rect 19368 -26168 19428 -26008
rect 20382 -26168 20442 -26008
rect 19366 -26174 19428 -26168
rect 19426 -26180 19428 -26174
rect 20380 -26174 20442 -26168
rect 19366 -26240 19426 -26234
rect 20440 -26180 20442 -26174
rect 20380 -26240 20440 -26234
rect 20892 -26430 20952 -25918
rect 21916 -25918 21922 -25350
rect 21956 -25350 21970 -25342
rect 22928 -25342 22988 -25204
rect 21956 -25918 21962 -25350
rect 22928 -25360 22940 -25342
rect 21916 -25930 21962 -25918
rect 22934 -25918 22940 -25360
rect 22974 -25360 22988 -25342
rect 22974 -25918 22980 -25360
rect 22934 -25930 22980 -25918
rect 21402 -25962 21462 -25960
rect 21186 -25968 21674 -25962
rect 21186 -26002 21198 -25968
rect 21662 -26002 21674 -25968
rect 21186 -26008 21674 -26002
rect 22204 -25968 22692 -25962
rect 22204 -26002 22216 -25968
rect 22680 -26002 22692 -25968
rect 22204 -26008 22692 -26002
rect 21402 -26168 21462 -26008
rect 23054 -26066 23114 -23986
rect 23762 -24928 23822 -16586
rect 23756 -24988 23762 -24928
rect 23822 -24988 23828 -24928
rect 23048 -26126 23054 -26066
rect 23114 -26126 23120 -26066
rect 21402 -26174 21464 -26168
rect 21402 -26180 21404 -26174
rect 21404 -26240 21464 -26234
rect 24816 -26330 24822 -12070
rect 24922 -26330 24928 -12070
rect -8118 -26476 -7968 -26430
rect -7922 -26476 -4748 -26430
rect -4688 -26476 1704 -26430
rect 1764 -26476 23806 -26430
rect 23866 -26476 23968 -26430
rect -8118 -26630 -8072 -26476
rect 23928 -26630 23968 -26476
rect -8118 -26676 23968 -26630
rect -11616 -27116 -11606 -26816
rect 24206 -27116 24216 -26816
rect 24816 -27116 24928 -26330
rect -12328 -27122 24928 -27116
rect -12328 -27222 -12222 -27122
rect 24822 -27222 24928 -27122
rect -12328 -27228 24928 -27222
<< via1 >>
rect 484 3916 1084 4216
rect 24116 3916 24716 4216
rect 4061 3620 20846 3834
rect 7986 1858 8046 1918
rect 9068 1858 9128 1918
rect 10026 1858 10086 1918
rect 8512 1612 8572 1672
rect 10548 1612 10608 1672
rect 6330 680 6390 740
rect 7494 680 7554 740
rect 6200 476 6260 536
rect 4192 -1708 4252 -1648
rect 7494 476 7554 536
rect 13090 1858 13150 1918
rect 14108 1858 14168 1918
rect 12586 1614 12646 1674
rect 9530 576 9590 636
rect 7980 -674 8040 -614
rect 15132 1858 15192 1918
rect 16144 1858 16204 1918
rect 14616 1614 14676 1674
rect 11566 576 11626 636
rect 16658 1616 16718 1676
rect 13604 680 13664 740
rect 13600 476 13660 536
rect 10036 -458 10096 -398
rect 10546 -458 10606 -398
rect 9528 -560 9592 -496
rect 9018 -674 9078 -614
rect 10030 -674 10090 -614
rect 6330 -1994 6390 -1934
rect 6686 -4402 6746 -4342
rect 6560 -5012 6620 -4952
rect 3676 -5966 3736 -5906
rect 3784 -6078 3844 -6018
rect 2014 -7000 2074 -6940
rect 4698 -5966 4758 -5906
rect 4568 -6078 4628 -6018
rect 3174 -7110 3234 -7050
rect 5208 -7000 5268 -6940
rect 1888 -8088 1948 -8028
rect 3690 -8034 3750 -7974
rect 3796 -8134 3856 -8074
rect 6360 -7110 6420 -7050
rect 4700 -8034 4760 -7974
rect 6552 -7238 6612 -7178
rect 4582 -8134 4642 -8074
rect 1402 -9144 1462 -9084
rect 1542 -9320 1602 -9260
rect 2442 -9494 2502 -9434
rect 6802 -5012 6862 -4952
rect 7488 -1848 7552 -1784
rect 7312 -1994 7372 -1934
rect 11404 -560 11468 -496
rect 17668 1616 17728 1676
rect 19202 1858 19262 1918
rect 20214 1858 20274 1918
rect 18690 1616 18750 1676
rect 15638 680 15698 740
rect 15636 476 15696 536
rect 16138 476 16198 536
rect 12580 -458 12640 -398
rect 11040 -666 11100 -606
rect 12064 -666 12124 -606
rect 8510 -1596 8570 -1536
rect 9526 -1710 9590 -1646
rect 13092 -666 13152 -606
rect 21232 1858 21292 1918
rect 20726 1616 20786 1676
rect 17672 576 17732 636
rect 17158 476 17218 536
rect 14618 -460 14678 -400
rect 10546 -1596 10606 -1536
rect 11068 -1596 11128 -1536
rect 11566 -1596 11626 -1536
rect 18184 476 18244 536
rect 19706 576 19766 636
rect 18690 472 18750 532
rect 19204 472 19264 532
rect 19708 472 19768 532
rect 20214 472 20274 532
rect 20734 472 20794 532
rect 15638 -558 15698 -498
rect 21746 680 21806 740
rect 22996 680 23056 740
rect 16654 -460 16714 -400
rect 17154 -460 17214 -400
rect 17668 -460 17728 -400
rect 18192 -460 18252 -400
rect 18690 -460 18750 -400
rect 19192 -460 19252 -400
rect 12040 -1600 12100 -1540
rect 7428 -2100 7488 -2040
rect 7990 -2100 8050 -2040
rect 9032 -2100 9092 -2040
rect 10032 -2100 10092 -2040
rect 12580 -1538 12640 -1536
rect 12548 -1596 12640 -1538
rect 13040 -1596 13100 -1536
rect 12548 -1598 12608 -1596
rect 13598 -1852 13662 -1788
rect 14084 -1594 14144 -1534
rect 13194 -2100 13254 -2040
rect 14616 -1596 14676 -1536
rect 19706 -462 19766 -402
rect 20214 -462 20274 -402
rect 20724 -462 20784 -402
rect 19196 -674 19256 -614
rect 20208 -674 20268 -614
rect 16128 -1594 16188 -1534
rect 15634 -1994 15698 -1930
rect 14204 -2100 14264 -2040
rect 15146 -2100 15206 -2040
rect 16654 -1540 16714 -1538
rect 16622 -1598 16714 -1540
rect 16622 -1600 16682 -1598
rect 17150 -1604 17210 -1544
rect 17638 -1542 17698 -1540
rect 17638 -1600 17732 -1542
rect 17672 -1602 17732 -1600
rect 21746 -558 21806 -498
rect 21210 -674 21270 -614
rect 18150 -1604 18210 -1544
rect 18690 -1600 18750 -1540
rect 20724 -1600 20784 -1540
rect 19706 -1710 19770 -1646
rect 22992 -1848 23056 -1784
rect 21740 -1994 21800 -1934
rect 7542 -2302 7602 -2242
rect 10720 -2302 10780 -2242
rect 8686 -3238 8746 -3178
rect 9190 -3346 9250 -3286
rect 10720 -3238 10780 -3178
rect 10212 -3346 10272 -3286
rect 11230 -3346 11290 -3286
rect 8682 -4270 8742 -4210
rect 9188 -4404 9248 -4344
rect 14788 -2302 14848 -2242
rect 12762 -3238 12822 -3178
rect 12254 -3346 12314 -3286
rect 13268 -3346 13328 -3286
rect 10202 -4408 10262 -4348
rect 11234 -4400 11294 -4340
rect 14788 -3238 14848 -3178
rect 14286 -3346 14346 -3286
rect 15296 -3346 15356 -3286
rect 12762 -4270 12822 -4210
rect 12232 -4400 12292 -4340
rect 13276 -4400 13336 -4340
rect 18864 -2302 18924 -2242
rect 16830 -3238 16890 -3178
rect 16318 -3346 16378 -3286
rect 17332 -3346 17392 -3286
rect 14280 -4404 14340 -4344
rect 15296 -4404 15356 -4344
rect 14080 -4612 14140 -4552
rect 7312 -4930 7372 -4870
rect 8478 -4930 8538 -4870
rect 7044 -5976 7104 -5916
rect 6802 -7134 6862 -7074
rect 6798 -7348 6858 -7288
rect 6686 -8390 6746 -8330
rect 1282 -9644 1342 -9584
rect 7180 -6074 7240 -6014
rect 7044 -9648 7104 -9588
rect 10514 -4930 10574 -4870
rect 11022 -4934 11086 -4870
rect 9496 -5878 9556 -5818
rect 22060 -2302 22120 -2242
rect 18866 -3238 18926 -3178
rect 18364 -3346 18424 -3286
rect 19374 -3346 19434 -3286
rect 16830 -4270 16890 -4210
rect 16300 -4404 16360 -4344
rect 17332 -4400 17392 -4340
rect 15816 -4612 15876 -4552
rect 15096 -4812 15160 -4748
rect 20902 -3238 20962 -3178
rect 20396 -3346 20456 -3286
rect 18348 -4404 18408 -4344
rect 19376 -4404 19436 -4344
rect 20898 -4270 20958 -4210
rect 20396 -4404 20456 -4344
rect 22854 -4402 22914 -4342
rect 21714 -4628 21774 -4568
rect 19160 -4812 19224 -4748
rect 20184 -4812 20248 -4748
rect 21196 -4812 21260 -4748
rect 15098 -4934 15162 -4870
rect 11532 -5878 11592 -5818
rect 11874 -5876 11934 -5816
rect 9496 -6074 9556 -6014
rect 10516 -6072 10576 -6012
rect 8482 -6184 8542 -6124
rect 10516 -6184 10576 -6124
rect 7464 -7348 7524 -7288
rect 14588 -5876 14648 -5816
rect 18660 -4930 18720 -4870
rect 20694 -4930 20754 -4870
rect 15606 -6072 15666 -6012
rect 13572 -6186 13632 -6126
rect 15606 -6186 15666 -6126
rect 9498 -7238 9558 -7178
rect 9498 -7442 9558 -7382
rect 11534 -7238 11594 -7178
rect 11532 -7340 11592 -7280
rect 11532 -7442 11592 -7382
rect 8480 -8390 8540 -8330
rect 7312 -8598 7372 -8538
rect 9494 -8700 9554 -8640
rect 13568 -7134 13628 -7074
rect 10516 -8390 10576 -8330
rect 10516 -8498 10576 -8438
rect 14588 -7134 14648 -7074
rect 14588 -7440 14648 -7380
rect 18662 -6186 18722 -6126
rect 15606 -7440 15666 -7380
rect 19676 -5878 19736 -5818
rect 20696 -6186 20756 -6126
rect 21712 -5878 21772 -5818
rect 16624 -7134 16684 -7074
rect 16622 -7440 16682 -7380
rect 11534 -8382 11594 -8322
rect 13336 -8382 13396 -8322
rect 11528 -8700 11588 -8640
rect 11732 -8712 11792 -8652
rect 8476 -9648 8536 -9588
rect 13570 -8388 13630 -8328
rect 18658 -7238 18718 -7178
rect 19526 -7120 19586 -7060
rect 19674 -7230 19734 -7170
rect 19526 -7440 19586 -7380
rect 19678 -7438 19738 -7378
rect 15606 -8388 15666 -8328
rect 15604 -8498 15664 -8438
rect 10512 -9648 10572 -9588
rect 7180 -9778 7240 -9718
rect 2336 -9906 2396 -9846
rect 2216 -10024 2276 -9964
rect 15094 -8712 15154 -8652
rect 20694 -7340 20754 -7280
rect 23290 -4270 23350 -4210
rect 22996 -4630 23056 -4570
rect 23138 -4930 23198 -4870
rect 22978 -6072 23038 -6012
rect 21714 -7230 21774 -7170
rect 22854 -7230 22914 -7170
rect 21712 -7438 21772 -7378
rect 16110 -8712 16170 -8652
rect 18660 -8386 18720 -8326
rect 19170 -8712 19230 -8652
rect 19682 -8700 19742 -8640
rect 20696 -8386 20756 -8326
rect 22978 -7438 23038 -7378
rect 22854 -8498 22914 -8438
rect 21716 -8700 21776 -8640
rect 18664 -9648 18724 -9588
rect 20700 -9648 20760 -9588
rect 11534 -9918 11594 -9858
rect 23290 -6186 23350 -6126
rect 23138 -9918 23198 -9858
rect 1770 -10142 1830 -10082
rect -13630 -10670 -2866 -10378
rect 1888 -11418 1948 -11358
rect 2216 -11408 2276 -11348
rect 1282 -11554 1342 -11494
rect 1402 -11552 1462 -11492
rect 1542 -11534 1602 -11474
rect 1770 -11518 1830 -11458
rect 1150 -11682 1210 -11622
rect -1562 -12280 -1502 -12220
rect -36 -12414 24 -12354
rect 1150 -18882 1210 -18822
rect -3398 -19808 -3338 -19748
rect -9508 -19954 -9448 -19894
rect -5428 -19954 -5368 -19894
rect -10662 -20082 -10602 -20022
rect -7984 -20082 -7924 -20022
rect -6952 -20082 -6892 -20022
rect -9004 -21044 -8944 -20984
rect -9504 -21148 -9444 -21088
rect -7980 -21044 -7920 -20984
rect -8486 -21252 -8426 -21192
rect -10662 -22314 -10602 -22254
rect -3892 -20082 -3832 -20022
rect -6948 -21044 -6888 -20984
rect -7468 -21148 -7408 -21088
rect -1368 -19954 -1308 -19894
rect 816 -19954 876 -19894
rect -2896 -20082 -2836 -20022
rect -5948 -21044 -5888 -20984
rect -4928 -21044 -4868 -20984
rect -5432 -21148 -5372 -21088
rect -6450 -21252 -6390 -21192
rect -9012 -22314 -8952 -22254
rect -7474 -22194 -7414 -22134
rect -3908 -21044 -3848 -20984
rect -4418 -21252 -4358 -21192
rect -5942 -22314 -5882 -22254
rect -2898 -21044 -2838 -20984
rect -3398 -21148 -3338 -21088
rect -1884 -21044 -1824 -20984
rect -866 -21044 -806 -20984
rect -1362 -21148 -1302 -21088
rect -2384 -21252 -2324 -21192
rect -4934 -22314 -4874 -22254
rect -8486 -23258 -8426 -23198
rect -9500 -23366 -9440 -23306
rect -9006 -23478 -8946 -23418
rect -7464 -23366 -7404 -23306
rect -7982 -23478 -7922 -23418
rect -3398 -22194 -3338 -22134
rect -6450 -23258 -6390 -23198
rect -6950 -23478 -6890 -23418
rect -340 -21252 -280 -21192
rect -1872 -22314 -1812 -22254
rect 936 -21044 996 -20984
rect 816 -22194 876 -22134
rect -846 -22314 -786 -22254
rect -4418 -23258 -4358 -23198
rect -5428 -23366 -5368 -23306
rect -5950 -23478 -5890 -23418
rect -4930 -23478 -4870 -23418
rect -3394 -23366 -3334 -23306
rect -3910 -23478 -3850 -23418
rect -10662 -24440 -10602 -24380
rect -7992 -24440 -7932 -24380
rect -6960 -24440 -6900 -24380
rect -2900 -23478 -2840 -23418
rect -2384 -23258 -2324 -23198
rect -340 -23258 -280 -23198
rect -1358 -23366 -1298 -23306
rect -1886 -23478 -1826 -23418
rect -868 -23478 -808 -23418
rect -3900 -24440 -3840 -24380
rect -2904 -24440 -2844 -24380
rect 936 -23478 996 -23418
rect -9506 -24570 -9446 -24510
rect -5426 -24570 -5366 -24510
rect -1366 -24570 -1306 -24510
rect 816 -24570 876 -24510
rect -8028 -25936 -7968 -25876
rect -5990 -25936 -5930 -25876
rect -3954 -25936 -3894 -25876
rect -7010 -26048 -6950 -25988
rect -1918 -25936 -1858 -25876
rect -2936 -26048 -2876 -25988
rect 1282 -19954 1342 -19894
rect 1402 -20082 1462 -20022
rect 1660 -11672 1720 -11612
rect 1770 -12414 1830 -12354
rect 2336 -11416 2396 -11356
rect 2216 -12280 2276 -12220
rect 2012 -13638 2072 -13578
rect 1886 -15340 1946 -15280
rect 1660 -17800 1720 -17740
rect 1542 -21044 1602 -20984
rect 2224 -13974 2284 -13914
rect 2120 -15234 2180 -15174
rect 2012 -16334 2072 -16274
rect 2442 -11552 2502 -11492
rect 13254 -11902 13314 -11842
rect 18358 -11902 18418 -11842
rect 22418 -11908 22478 -11848
rect 3586 -13638 3646 -13578
rect 4600 -13854 4660 -13794
rect 6640 -13854 6700 -13794
rect 8680 -13854 8740 -13794
rect 10710 -13854 10770 -13794
rect 12750 -13854 12810 -13794
rect 14782 -13854 14842 -13794
rect 16822 -13854 16882 -13794
rect 18858 -13854 18918 -13794
rect 20892 -13854 20952 -13794
rect 2568 -13974 2628 -13914
rect 4092 -13980 4152 -13920
rect 2442 -14096 2502 -14036
rect 5106 -13980 5166 -13920
rect 6128 -13980 6188 -13920
rect 7142 -13980 7202 -13920
rect 8168 -13980 8228 -13920
rect 7656 -14096 7716 -14036
rect 9180 -13980 9240 -13920
rect 10216 -13980 10276 -13920
rect 11222 -13980 11282 -13920
rect 12236 -13980 12296 -13920
rect 4604 -15018 4664 -14958
rect 4096 -15128 4156 -15068
rect 3586 -15234 3646 -15174
rect 2572 -15340 2632 -15280
rect 3070 -15340 3130 -15280
rect 3582 -15340 3642 -15280
rect 5118 -15128 5178 -15068
rect 6644 -15018 6704 -14958
rect 6132 -15128 6192 -15068
rect 5626 -15234 5686 -15174
rect 8676 -15018 8736 -14958
rect 7146 -15128 7206 -15068
rect 8164 -15128 8224 -15068
rect 7656 -15234 7716 -15174
rect 2442 -16230 2502 -16170
rect 2566 -16334 2626 -16274
rect 4086 -16334 4146 -16274
rect 4598 -16334 4658 -16274
rect 2336 -16456 2396 -16396
rect 2224 -16570 2284 -16510
rect 3072 -16570 3132 -16510
rect 4604 -16568 4664 -16508
rect 9190 -15128 9250 -15068
rect 13252 -13980 13312 -13920
rect 14260 -13980 14320 -13920
rect 15276 -13980 15336 -13920
rect 16300 -13980 16360 -13920
rect 17322 -13980 17382 -13920
rect 18344 -13980 18404 -13920
rect 17844 -14096 17904 -14036
rect 10708 -15018 10768 -14958
rect 9696 -15234 9756 -15174
rect 10210 -15128 10270 -15068
rect 9862 -15340 9922 -15280
rect 5620 -16230 5680 -16170
rect 5622 -16334 5682 -16274
rect 11230 -15128 11290 -15068
rect 12744 -15018 12804 -14958
rect 12232 -15128 12292 -15068
rect 11730 -15234 11790 -15174
rect 11730 -15340 11790 -15280
rect 13258 -15128 13318 -15068
rect 19362 -13980 19422 -13920
rect 20376 -13980 20436 -13920
rect 21400 -13980 21460 -13920
rect 21916 -14096 21976 -14036
rect 23048 -14096 23108 -14036
rect 14780 -15018 14840 -14958
rect 14276 -15128 14336 -15068
rect 13766 -15234 13826 -15174
rect 13768 -15340 13828 -15280
rect 15284 -15128 15344 -15068
rect 16818 -15018 16878 -14958
rect 16296 -15128 16356 -15068
rect 15802 -15234 15862 -15174
rect 15648 -15340 15708 -15280
rect 6634 -16334 6694 -16274
rect 6640 -16568 6700 -16508
rect 7654 -16334 7714 -16274
rect 2448 -17498 2508 -17438
rect 3586 -17498 3646 -17438
rect 2336 -17698 2396 -17638
rect 2230 -17800 2290 -17740
rect 2120 -21252 2180 -21192
rect 2336 -18934 2396 -18874
rect 1888 -21402 1948 -21342
rect 2230 -21290 2290 -21230
rect 3584 -17698 3644 -17638
rect 4602 -17578 4662 -17518
rect 8676 -16230 8736 -16170
rect 18856 -15018 18916 -14958
rect 17328 -15128 17388 -15068
rect 18342 -15128 18402 -15068
rect 17842 -15234 17902 -15174
rect 14782 -16230 14842 -16170
rect 10712 -16334 10772 -16274
rect 12750 -16334 12810 -16274
rect 9696 -16456 9756 -16396
rect 11730 -16456 11790 -16396
rect 13760 -16456 13820 -16396
rect 5620 -17474 5680 -17414
rect 5116 -17692 5176 -17632
rect 6642 -17578 6702 -17518
rect 6120 -17692 6180 -17632
rect 3584 -18730 3644 -18670
rect 4090 -18832 4150 -18772
rect 7656 -17474 7716 -17414
rect 7132 -17692 7192 -17632
rect 8674 -17578 8734 -17518
rect 8152 -17692 8212 -17632
rect 8674 -17690 8734 -17630
rect 10708 -17578 10768 -17518
rect 9692 -17800 9752 -17740
rect 5622 -18730 5682 -18670
rect 5620 -18934 5680 -18874
rect 10710 -17690 10770 -17630
rect 11726 -17800 11786 -17740
rect 15800 -16334 15860 -16274
rect 19360 -15128 19420 -15068
rect 20892 -15018 20952 -14958
rect 20384 -15128 20444 -15068
rect 19872 -15234 19932 -15174
rect 19872 -15338 19932 -15278
rect 16818 -16334 16878 -16274
rect 17838 -16334 17898 -16274
rect 12748 -17578 12808 -17518
rect 12746 -17690 12806 -17630
rect 14782 -17578 14842 -17518
rect 14978 -17582 15038 -17522
rect 13766 -17800 13826 -17740
rect 14782 -17690 14842 -17630
rect 21404 -15128 21464 -15068
rect 21912 -15234 21972 -15174
rect 23048 -15338 23108 -15278
rect 19876 -16230 19936 -16170
rect 18854 -16334 18914 -16274
rect 20890 -16334 20950 -16274
rect 15800 -17474 15860 -17414
rect 14978 -17800 15038 -17740
rect 15272 -17798 15332 -17738
rect 7658 -18730 7718 -18670
rect 4604 -19034 4664 -18974
rect 6128 -18940 6188 -18880
rect 7150 -18940 7210 -18880
rect 6638 -19034 6698 -18974
rect 9690 -18730 9750 -18670
rect 9182 -18832 9242 -18772
rect 8164 -18940 8224 -18880
rect 9182 -18940 9242 -18880
rect 8674 -19034 8734 -18974
rect 4086 -19958 4146 -19898
rect 4996 -19958 5056 -19898
rect 4086 -20174 4146 -20114
rect 2450 -20278 2510 -20218
rect 5998 -19958 6058 -19898
rect 5124 -20174 5184 -20114
rect 7150 -19958 7210 -19898
rect 6638 -20060 6698 -20000
rect 6138 -20174 6198 -20114
rect 4084 -21186 4144 -21126
rect 3586 -21290 3646 -21230
rect 3582 -21500 3642 -21440
rect 5092 -21186 5152 -21126
rect 4602 -21402 4662 -21342
rect 10202 -18940 10262 -18880
rect 16816 -17690 16876 -17630
rect 16300 -17798 16360 -17738
rect 16818 -17804 16878 -17744
rect 17836 -17474 17896 -17414
rect 18854 -17690 18914 -17630
rect 19870 -17582 19930 -17522
rect 20374 -17586 20434 -17526
rect 23034 -16568 23094 -16508
rect 20894 -17690 20954 -17630
rect 18854 -17804 18914 -17744
rect 14272 -18718 14332 -18658
rect 13766 -18846 13826 -18786
rect 15802 -19044 15862 -18984
rect 8160 -19958 8220 -19898
rect 9166 -19958 9226 -19898
rect 10210 -19958 10270 -19898
rect 10710 -19952 10770 -19892
rect 9164 -20174 9224 -20114
rect 10204 -20174 10264 -20114
rect 9688 -20278 9748 -20218
rect 6106 -21186 6166 -21126
rect 7144 -21186 7204 -21126
rect 6640 -21402 6700 -21342
rect 5620 -21500 5680 -21440
rect 11218 -20174 11278 -20114
rect 12746 -19952 12806 -19892
rect 12226 -20174 12286 -20114
rect 13270 -20174 13330 -20114
rect 11730 -20278 11790 -20218
rect 20892 -17804 20952 -17744
rect 17314 -18940 17374 -18880
rect 14782 -19952 14842 -19892
rect 14260 -20174 14320 -20114
rect 15278 -20174 15338 -20114
rect 13768 -20278 13828 -20218
rect 21910 -17474 21970 -17414
rect 22928 -17456 22988 -17396
rect 23162 -16586 23222 -16526
rect 23528 -17586 23588 -17526
rect 23278 -17690 23338 -17630
rect 19366 -18718 19426 -18658
rect 19504 -18714 19564 -18654
rect 23034 -17804 23094 -17744
rect 20386 -18714 20446 -18654
rect 21392 -18714 21452 -18654
rect 18344 -18940 18404 -18880
rect 19504 -18940 19564 -18880
rect 19872 -18940 19932 -18880
rect 19872 -19044 19932 -18984
rect 21910 -18718 21970 -18658
rect 21910 -18846 21970 -18786
rect 20888 -19042 20948 -18982
rect 16820 -19952 16880 -19892
rect 16812 -20060 16872 -20000
rect 16312 -20174 16372 -20114
rect 15802 -20278 15862 -20218
rect 16314 -20282 16374 -20222
rect 17336 -20282 17396 -20222
rect 17836 -20276 17896 -20216
rect 8162 -21186 8222 -21126
rect 8678 -21180 8738 -21120
rect 10714 -21180 10774 -21120
rect 12746 -21180 12806 -21120
rect 14780 -21180 14840 -21120
rect 7660 -21500 7720 -21440
rect 2448 -22522 2508 -22462
rect 3588 -22738 3648 -22678
rect 4602 -22424 4662 -22364
rect 4606 -22618 4666 -22558
rect 5620 -22522 5680 -22462
rect 11730 -21290 11790 -21230
rect 13766 -21290 13826 -21230
rect 10712 -21402 10772 -21342
rect 9696 -21500 9756 -21440
rect 6638 -22424 6698 -22364
rect 7144 -22522 7204 -22462
rect 6642 -22618 6702 -22558
rect 8676 -22424 8736 -22364
rect 8166 -22522 8226 -22462
rect 7656 -22738 7716 -22678
rect 2336 -23654 2396 -23594
rect 2230 -23780 2290 -23720
rect 9188 -22522 9248 -22462
rect 8670 -22618 8730 -22558
rect 18856 -19952 18916 -19892
rect 18852 -20060 18912 -20000
rect 19344 -20174 19404 -20114
rect 20894 -19952 20954 -19892
rect 20890 -20060 20950 -20000
rect 20382 -20174 20442 -20114
rect 19870 -20276 19930 -20216
rect 15802 -21178 15862 -21118
rect 16156 -21178 16216 -21118
rect 15798 -21290 15858 -21230
rect 15308 -21388 15368 -21328
rect 10538 -22404 10598 -22344
rect 10708 -22404 10768 -22344
rect 10192 -22522 10252 -22462
rect 9690 -22738 9750 -22678
rect 5620 -23780 5680 -23720
rect 6140 -23768 6200 -23708
rect 4602 -23882 4662 -23822
rect 6638 -23882 6698 -23822
rect 5620 -23986 5680 -23926
rect 2448 -24884 2508 -24824
rect 2120 -24988 2180 -24928
rect 3584 -24988 3644 -24928
rect 4092 -25094 4152 -25034
rect 1070 -26048 1130 -25988
rect 10538 -22618 10598 -22558
rect 10714 -22612 10774 -22552
rect 16346 -21388 16406 -21328
rect 17322 -21388 17382 -21328
rect 16156 -21496 16216 -21436
rect 21408 -20174 21468 -20114
rect 21912 -20276 21972 -20216
rect 19874 -21178 19934 -21118
rect 18338 -21388 18398 -21328
rect 20364 -21388 20424 -21328
rect 17836 -21500 17896 -21440
rect 19872 -21500 19932 -21440
rect 12750 -22404 12810 -22344
rect 14782 -22404 14842 -22344
rect 16822 -22404 16882 -22344
rect 15800 -22502 15860 -22442
rect 12742 -22612 12802 -22552
rect 7658 -23882 7718 -23822
rect 8674 -23882 8734 -23822
rect 5618 -24884 5678 -24824
rect 5624 -24988 5684 -24928
rect 5112 -25094 5172 -25034
rect 4604 -25204 4664 -25144
rect 6136 -25094 6196 -25034
rect 9694 -23882 9754 -23822
rect 14786 -22612 14846 -22552
rect 16814 -22612 16874 -22552
rect 17840 -22738 17900 -22678
rect 21394 -21388 21454 -21328
rect 21908 -21500 21968 -21440
rect 18852 -22612 18912 -22552
rect 21906 -22502 21966 -22442
rect 20892 -22612 20952 -22552
rect 21410 -22608 21470 -22548
rect 22922 -22608 22982 -22548
rect 19870 -22738 19930 -22678
rect 20396 -22736 20456 -22676
rect 11724 -23654 11784 -23594
rect 13766 -23654 13826 -23594
rect 15802 -23654 15862 -23594
rect 11220 -23768 11280 -23708
rect 16308 -23764 16368 -23704
rect 10712 -23882 10772 -23822
rect 12742 -23882 12802 -23822
rect 14780 -23882 14840 -23822
rect 16816 -23882 16876 -23822
rect 10556 -23986 10616 -23926
rect 7654 -24988 7714 -24928
rect 7154 -25094 7214 -25034
rect 8168 -25094 8228 -25034
rect 6640 -25204 6700 -25144
rect 2448 -26126 2508 -26066
rect 3584 -26126 3644 -26066
rect 4096 -26234 4156 -26174
rect 9848 -24882 9908 -24822
rect 9694 -24988 9754 -24928
rect 9200 -25094 9260 -25034
rect 8678 -25204 8738 -25144
rect 5110 -26234 5170 -26174
rect 6132 -26234 6192 -26174
rect 10212 -25094 10272 -25034
rect 11726 -24882 11786 -24822
rect 11730 -24988 11790 -24928
rect 11220 -25094 11280 -25034
rect 10716 -25204 10776 -25144
rect 7654 -26126 7714 -26066
rect 7146 -26234 7206 -26174
rect 8172 -26234 8232 -26174
rect 12238 -25094 12298 -25034
rect 13764 -24882 13824 -24822
rect 13766 -24988 13826 -24928
rect 13264 -25094 13324 -25034
rect 12752 -25204 12812 -25144
rect 9184 -26234 9244 -26174
rect 10220 -26234 10280 -26174
rect 14266 -25094 14326 -25034
rect 16962 -23986 17022 -23926
rect 21910 -22736 21970 -22676
rect 17838 -23882 17898 -23822
rect 18856 -23654 18916 -23594
rect 18858 -23882 18918 -23822
rect 15634 -24882 15694 -24822
rect 15286 -25094 15346 -25034
rect 15800 -24988 15860 -24928
rect 14788 -25204 14848 -25144
rect 11226 -26234 11286 -26174
rect 12240 -26234 12300 -26174
rect 16306 -25094 16366 -25034
rect 19872 -23882 19932 -23822
rect 19872 -23986 19932 -23926
rect 20888 -23654 20948 -23594
rect 23162 -18718 23222 -18658
rect 23400 -18940 23460 -18880
rect 23278 -19042 23338 -18982
rect 23162 -20276 23222 -20216
rect 23158 -21178 23218 -21118
rect 23278 -22404 23338 -22344
rect 23158 -22502 23218 -22442
rect 23034 -23654 23094 -23594
rect 21408 -23764 21468 -23704
rect 22416 -23764 22476 -23704
rect 23526 -20174 23586 -20114
rect 23528 -22608 23588 -22548
rect 23400 -22736 23460 -22676
rect 23762 -16586 23822 -16526
rect 23650 -23764 23710 -23704
rect 20894 -23882 20954 -23822
rect 17840 -24988 17900 -24928
rect 17332 -25094 17392 -25034
rect 18350 -25094 18410 -25034
rect 16820 -25204 16880 -25144
rect 13256 -26234 13316 -26174
rect 14264 -26234 14324 -26174
rect 19870 -24988 19930 -24928
rect 19364 -25094 19424 -25034
rect 18852 -25204 18912 -25144
rect 15280 -26234 15340 -26174
rect 16304 -26234 16364 -26174
rect 20378 -25094 20438 -25034
rect 23054 -23986 23114 -23926
rect 21910 -24882 21970 -24822
rect 21910 -24988 21970 -24928
rect 21400 -25094 21460 -25034
rect 20892 -25204 20952 -25144
rect 17834 -26126 17894 -26066
rect 17326 -26234 17386 -26174
rect 18348 -26234 18408 -26174
rect 19366 -26234 19426 -26174
rect 20380 -26234 20440 -26174
rect 23762 -24988 23822 -24928
rect 23054 -26126 23114 -26066
rect 21404 -26234 21464 -26174
rect -8072 -26630 23928 -26476
rect -12216 -27116 -11616 -26816
rect 24216 -27116 24816 -26816
<< metal2 >>
rect 484 4216 1084 4226
rect 484 3906 1084 3916
rect 24116 4216 24716 4226
rect 24116 3906 24716 3916
rect 3998 3834 20878 3866
rect 3998 3620 4061 3834
rect 20846 3620 20878 3834
rect 3998 3600 20878 3620
rect 3998 3598 8352 3600
rect 7986 1918 8046 1924
rect 9068 1918 9128 1924
rect 10026 1918 10086 1924
rect 13090 1918 13150 1924
rect 14108 1918 14168 1924
rect 15132 1918 15192 1924
rect 16144 1918 16204 1924
rect 19202 1918 19262 1924
rect 20214 1918 20274 1924
rect 21232 1918 21292 1924
rect 8046 1858 9068 1918
rect 9128 1858 10026 1918
rect 10086 1858 13090 1918
rect 13150 1858 14108 1918
rect 14168 1858 15132 1918
rect 15192 1858 16144 1918
rect 16204 1858 19202 1918
rect 19262 1858 20214 1918
rect 20274 1858 21232 1918
rect 7986 1852 8046 1858
rect 9068 1852 9128 1858
rect 10026 1852 10086 1858
rect 13090 1852 13150 1858
rect 14108 1852 14168 1858
rect 15132 1852 15192 1858
rect 16144 1852 16204 1858
rect 19202 1852 19262 1858
rect 20214 1852 20274 1858
rect 21232 1852 21292 1858
rect 8512 1672 8572 1678
rect 10548 1672 10608 1678
rect 12586 1674 12646 1680
rect 14616 1674 14676 1680
rect 16658 1676 16718 1682
rect 17668 1676 17728 1682
rect 18690 1676 18750 1682
rect 20726 1676 20786 1682
rect 8572 1612 10548 1672
rect 10608 1614 12586 1672
rect 12646 1614 14616 1674
rect 14676 1616 16658 1674
rect 16718 1616 17668 1676
rect 17728 1616 18690 1676
rect 18750 1616 20726 1676
rect 14676 1614 16856 1616
rect 10608 1612 12768 1614
rect 8512 1606 8572 1612
rect 10548 1606 10608 1612
rect 12586 1608 12646 1612
rect 14616 1608 14676 1614
rect 16658 1610 16718 1614
rect 17668 1610 17728 1616
rect 18690 1610 18750 1616
rect 20726 1610 20786 1616
rect 6330 740 6390 746
rect 7494 740 7554 746
rect 13604 740 13664 746
rect 6390 680 7494 740
rect 7554 680 13604 740
rect 6330 674 6390 680
rect 7494 674 7554 680
rect 13604 674 13664 680
rect 15638 740 15698 746
rect 21746 740 21806 746
rect 22996 740 23056 746
rect 15698 680 21746 740
rect 21806 680 22996 740
rect 15638 674 15698 680
rect 21746 674 21806 680
rect 22996 674 23056 680
rect 9530 636 9590 642
rect 11566 636 11626 642
rect 17672 636 17732 642
rect 19706 636 19766 642
rect 9590 576 11566 636
rect 11626 628 12044 636
rect 12260 628 17672 636
rect 11626 582 17672 628
rect 11626 578 14060 582
rect 11626 576 13034 578
rect 13272 576 14060 578
rect 14276 576 17672 582
rect 17732 576 19706 636
rect 9530 570 9590 576
rect 11566 570 11626 576
rect 17672 570 17732 576
rect 19706 570 19766 576
rect 6200 536 6260 542
rect 7494 536 7554 542
rect 13600 536 13660 542
rect 15636 536 15696 542
rect 6260 476 7494 536
rect 7554 476 13600 536
rect 13660 476 15636 536
rect 6200 470 6260 476
rect 7494 470 7554 476
rect 13600 470 13660 476
rect 15636 470 15696 476
rect 16138 536 16198 542
rect 17158 536 17218 542
rect 18184 536 18244 542
rect 16198 476 17158 536
rect 17218 476 18184 536
rect 16138 470 16198 476
rect 17158 470 17218 476
rect 18184 470 18244 476
rect 18690 532 18750 538
rect 19204 532 19264 538
rect 19708 532 19768 538
rect 20214 532 20274 538
rect 18750 472 19204 532
rect 19264 472 19708 532
rect 19768 472 20214 532
rect 20274 472 20734 532
rect 20794 472 20800 532
rect 18690 466 18750 472
rect 19204 466 19264 472
rect 19708 466 19768 472
rect 20214 466 20274 472
rect 10546 -398 10606 -392
rect 12580 -398 12640 -392
rect 14618 -398 14678 -394
rect 10030 -458 10036 -398
rect 10096 -458 10546 -398
rect 10606 -458 12580 -398
rect 12640 -400 14822 -398
rect 16654 -400 16714 -394
rect 17154 -400 17214 -394
rect 17668 -400 17728 -394
rect 18192 -400 18252 -394
rect 18690 -400 18750 -394
rect 19192 -400 19252 -394
rect 12640 -458 14618 -400
rect 10546 -464 10606 -458
rect 12580 -464 12640 -458
rect 14678 -460 16654 -400
rect 16714 -460 17154 -400
rect 17214 -460 17668 -400
rect 17728 -460 18192 -400
rect 18252 -460 18690 -400
rect 18750 -460 19192 -400
rect 19252 -402 19560 -400
rect 19706 -402 19766 -396
rect 20214 -402 20274 -396
rect 20724 -402 20784 -396
rect 19252 -460 19706 -402
rect 14618 -466 14678 -460
rect 16654 -466 16714 -460
rect 17154 -466 17214 -460
rect 17668 -466 17728 -460
rect 18192 -466 18252 -460
rect 18589 -462 19104 -460
rect 18690 -466 18750 -462
rect 19192 -466 19252 -460
rect 19354 -462 19706 -460
rect 19766 -462 20214 -402
rect 20274 -462 20724 -402
rect 19706 -468 19766 -462
rect 20214 -468 20274 -462
rect 20724 -468 20784 -462
rect 9528 -496 9592 -490
rect 11404 -496 11468 -490
rect 9592 -560 11404 -496
rect 9528 -566 9592 -560
rect 11404 -566 11468 -560
rect 15638 -498 15698 -492
rect 21746 -498 21806 -492
rect 15698 -558 21746 -498
rect 15638 -564 15698 -558
rect 21746 -564 21806 -558
rect 11040 -606 11100 -600
rect 12064 -606 12124 -600
rect 13092 -606 13152 -600
rect 9018 -614 9078 -608
rect 10030 -614 10090 -608
rect 7974 -674 7980 -614
rect 8040 -674 9018 -614
rect 9078 -674 10030 -614
rect 11100 -666 12064 -606
rect 12124 -666 13092 -606
rect 11040 -672 11100 -666
rect 12064 -672 12124 -666
rect 13092 -672 13152 -666
rect 19196 -614 19256 -608
rect 20208 -614 20268 -608
rect 21210 -614 21270 -608
rect 9018 -680 9078 -674
rect 10030 -680 10090 -674
rect 19256 -674 20208 -614
rect 20268 -674 21210 -614
rect 19196 -680 19256 -674
rect 20208 -680 20268 -674
rect 21210 -680 21270 -674
rect 8510 -1536 8570 -1530
rect 10546 -1536 10606 -1530
rect 11068 -1536 11128 -1530
rect 11566 -1536 11626 -1530
rect 12580 -1536 12640 -1530
rect 13040 -1536 13100 -1530
rect 14078 -1536 14084 -1534
rect 8570 -1596 10546 -1536
rect 10606 -1596 11068 -1536
rect 11128 -1596 11566 -1536
rect 11626 -1538 12580 -1536
rect 11626 -1540 12548 -1538
rect 11626 -1596 12040 -1540
rect 8510 -1602 8570 -1596
rect 10546 -1602 10606 -1596
rect 11068 -1602 11128 -1596
rect 11566 -1602 11626 -1596
rect 12034 -1600 12040 -1596
rect 12100 -1596 12548 -1540
rect 12640 -1596 13040 -1536
rect 13100 -1594 14084 -1536
rect 14144 -1536 14150 -1534
rect 14616 -1536 14676 -1530
rect 16122 -1536 16128 -1534
rect 14144 -1594 14616 -1536
rect 13100 -1596 14616 -1594
rect 14676 -1594 16128 -1536
rect 16188 -1536 16194 -1534
rect 16188 -1538 16500 -1536
rect 16654 -1538 16714 -1532
rect 18690 -1538 18750 -1534
rect 16188 -1540 16654 -1538
rect 16714 -1540 18878 -1538
rect 20724 -1540 20784 -1534
rect 16188 -1594 16622 -1540
rect 14676 -1596 16622 -1594
rect 12100 -1600 12106 -1596
rect 12542 -1598 12548 -1596
rect 12608 -1598 12640 -1596
rect 12580 -1602 12640 -1598
rect 13040 -1602 13100 -1596
rect 14616 -1602 14676 -1596
rect 14760 -1598 16086 -1596
rect 16292 -1598 16622 -1596
rect 16714 -1544 17638 -1540
rect 17698 -1542 18690 -1540
rect 16714 -1598 17150 -1544
rect 16616 -1600 16622 -1598
rect 16682 -1600 16714 -1598
rect 16654 -1604 16714 -1600
rect 17144 -1604 17150 -1598
rect 17210 -1598 17638 -1544
rect 17210 -1604 17216 -1598
rect 17632 -1600 17638 -1598
rect 17732 -1544 18690 -1542
rect 17732 -1598 18150 -1544
rect 17666 -1602 17672 -1600
rect 17732 -1602 17738 -1598
rect 18144 -1604 18150 -1598
rect 18210 -1598 18690 -1544
rect 18210 -1604 18216 -1598
rect 18750 -1600 20724 -1540
rect 18690 -1606 18750 -1600
rect 20724 -1606 20784 -1600
rect 4192 -1646 4252 -1642
rect 9526 -1646 9590 -1640
rect 19706 -1646 19770 -1640
rect 4190 -1648 9526 -1646
rect 4190 -1708 4192 -1648
rect 4252 -1708 9526 -1648
rect 4190 -1710 9526 -1708
rect 9590 -1710 19706 -1646
rect 4192 -1714 4252 -1710
rect 9526 -1716 9590 -1710
rect 19706 -1716 19770 -1710
rect 7488 -1784 7552 -1778
rect 7552 -1788 22992 -1784
rect 7552 -1848 13598 -1788
rect 7488 -1854 7552 -1848
rect 13592 -1852 13598 -1848
rect 13662 -1848 22992 -1788
rect 23056 -1848 23062 -1784
rect 13662 -1852 13668 -1848
rect 6330 -1934 6390 -1928
rect 15634 -1930 15698 -1924
rect 6390 -1994 7312 -1934
rect 7372 -1994 15634 -1934
rect 21740 -1934 21800 -1928
rect 15698 -1994 21740 -1934
rect 6330 -2000 6390 -1994
rect 15634 -2000 15698 -1994
rect 21740 -2000 21800 -1994
rect 7428 -2040 7488 -2034
rect 7990 -2040 8050 -2034
rect 9032 -2040 9092 -2034
rect 10032 -2040 10092 -2034
rect 13194 -2040 13254 -2034
rect 14204 -2040 14264 -2034
rect 15146 -2040 15206 -2034
rect 7488 -2100 7990 -2040
rect 8050 -2100 9032 -2040
rect 9092 -2100 10032 -2040
rect 10092 -2100 13194 -2040
rect 13254 -2100 14204 -2040
rect 14264 -2100 15146 -2040
rect 7428 -2106 7488 -2100
rect 7990 -2106 8050 -2100
rect 9032 -2106 9092 -2100
rect 10032 -2106 10092 -2100
rect 13194 -2106 13254 -2100
rect 14204 -2106 14264 -2100
rect 15146 -2106 15206 -2100
rect 7542 -2242 7602 -2236
rect 10720 -2242 10780 -2236
rect 14788 -2242 14848 -2236
rect 18864 -2242 18924 -2236
rect 22060 -2242 22120 -2236
rect 7602 -2302 10720 -2242
rect 10780 -2302 14788 -2242
rect 14848 -2302 18864 -2242
rect 18924 -2302 22060 -2242
rect 7542 -2308 7602 -2302
rect 10720 -2308 10780 -2302
rect 14788 -2308 14848 -2302
rect 18864 -2308 18924 -2302
rect 22060 -2308 22120 -2302
rect 8686 -3178 8746 -3172
rect 10720 -3178 10780 -3172
rect 12762 -3178 12822 -3172
rect 14788 -3178 14848 -3172
rect 16830 -3178 16890 -3172
rect 18866 -3178 18926 -3172
rect 20902 -3178 20962 -3172
rect 8746 -3238 10720 -3178
rect 10780 -3238 12762 -3178
rect 12822 -3238 14788 -3178
rect 14848 -3238 16830 -3178
rect 16890 -3238 18866 -3178
rect 18926 -3238 20902 -3178
rect 8686 -3244 8746 -3238
rect 10720 -3244 10780 -3238
rect 12762 -3244 12822 -3238
rect 14788 -3244 14848 -3238
rect 16830 -3244 16890 -3238
rect 18866 -3244 18926 -3238
rect 20902 -3244 20962 -3238
rect 9190 -3286 9250 -3280
rect 9250 -3346 10212 -3286
rect 10272 -3346 11230 -3286
rect 11290 -3346 12254 -3286
rect 12314 -3346 13268 -3286
rect 13328 -3346 14286 -3286
rect 14346 -3346 15296 -3286
rect 15356 -3346 16318 -3286
rect 16378 -3346 17332 -3286
rect 17392 -3346 18364 -3286
rect 18424 -3346 19374 -3286
rect 19434 -3346 20396 -3286
rect 20456 -3346 20462 -3286
rect 9190 -3352 9250 -3346
rect 8682 -4210 8742 -4204
rect 12762 -4210 12822 -4204
rect 16830 -4210 16890 -4204
rect 20898 -4210 20958 -4204
rect 23290 -4210 23350 -4204
rect 1150 -4270 8682 -4210
rect 8742 -4270 12762 -4210
rect 12822 -4270 16830 -4210
rect 16890 -4270 20898 -4210
rect 20958 -4270 23290 -4210
rect -13992 -10378 -2722 -10122
rect -13992 -10670 -13630 -10378
rect -2778 -10670 -2722 -10378
rect -13992 -10978 -2722 -10670
rect -13992 -11300 -1640 -10978
rect 1150 -11622 1210 -4270
rect 8682 -4276 8742 -4270
rect 12762 -4276 12822 -4270
rect 16830 -4276 16890 -4270
rect 20898 -4276 20958 -4270
rect 23290 -4276 23350 -4270
rect 6686 -4342 6746 -4336
rect 11228 -4342 11234 -4340
rect 6746 -4344 11234 -4342
rect 6746 -4402 9188 -4344
rect 6686 -4408 6746 -4402
rect 9182 -4404 9188 -4402
rect 9248 -4348 11234 -4344
rect 9248 -4402 10202 -4348
rect 9248 -4404 9254 -4402
rect 10196 -4408 10202 -4402
rect 10262 -4400 11234 -4348
rect 11294 -4342 11300 -4340
rect 12226 -4342 12232 -4340
rect 11294 -4400 12232 -4342
rect 12292 -4342 12298 -4340
rect 13270 -4342 13276 -4340
rect 12292 -4400 13276 -4342
rect 13336 -4342 13342 -4340
rect 17326 -4342 17332 -4340
rect 13336 -4344 17332 -4342
rect 13336 -4400 14280 -4344
rect 10262 -4402 14280 -4400
rect 10262 -4408 10268 -4402
rect 14274 -4404 14280 -4402
rect 14340 -4402 15296 -4344
rect 14340 -4404 14346 -4402
rect 15290 -4404 15296 -4402
rect 15356 -4402 16300 -4344
rect 15356 -4404 15362 -4402
rect 16294 -4404 16300 -4402
rect 16360 -4400 17332 -4344
rect 17392 -4342 17398 -4340
rect 22854 -4342 22914 -4336
rect 17392 -4344 22854 -4342
rect 17392 -4400 18348 -4344
rect 16360 -4402 18348 -4400
rect 16360 -4404 16366 -4402
rect 18342 -4404 18348 -4402
rect 18408 -4402 19376 -4344
rect 18408 -4404 18414 -4402
rect 19370 -4404 19376 -4402
rect 19436 -4402 20396 -4344
rect 19436 -4404 19442 -4402
rect 20390 -4404 20396 -4402
rect 20456 -4402 22854 -4344
rect 20456 -4404 20462 -4402
rect 22854 -4408 22914 -4402
rect 14080 -4552 14140 -4546
rect 14140 -4612 15816 -4552
rect 15876 -4612 15882 -4552
rect 21714 -4566 21774 -4562
rect 21712 -4568 23056 -4566
rect 14080 -4618 14140 -4612
rect 21712 -4628 21714 -4568
rect 21774 -4570 23056 -4568
rect 21774 -4628 22996 -4570
rect 21712 -4630 22996 -4628
rect 23056 -4630 23062 -4570
rect 21714 -4634 21774 -4630
rect 15096 -4748 15160 -4742
rect 19160 -4748 19224 -4742
rect 20184 -4748 20248 -4742
rect 21196 -4748 21260 -4742
rect 15160 -4812 19160 -4748
rect 19224 -4812 20184 -4748
rect 20248 -4812 21196 -4748
rect 15096 -4818 15160 -4812
rect 19160 -4818 19224 -4812
rect 20184 -4818 20248 -4812
rect 21196 -4818 21260 -4812
rect 7312 -4870 7372 -4864
rect 8478 -4870 8538 -4864
rect 10514 -4870 10574 -4864
rect 7372 -4930 8478 -4870
rect 8538 -4930 10514 -4870
rect 7312 -4936 7372 -4930
rect 8478 -4936 8538 -4930
rect 10514 -4936 10574 -4930
rect 11022 -4870 11086 -4864
rect 15098 -4870 15162 -4864
rect 11086 -4934 15098 -4870
rect 11022 -4940 11086 -4934
rect 15098 -4940 15162 -4934
rect 18660 -4870 18720 -4864
rect 20694 -4870 20754 -4864
rect 23138 -4870 23198 -4864
rect 18720 -4930 20694 -4870
rect 20754 -4930 23138 -4870
rect 18660 -4936 18720 -4930
rect 20694 -4936 20754 -4930
rect 23138 -4936 23198 -4930
rect 6560 -4952 6620 -4946
rect 6802 -4952 6862 -4946
rect 6620 -5012 6802 -4952
rect 6560 -5018 6620 -5012
rect 6802 -5018 6862 -5012
rect 9496 -5818 9556 -5812
rect 11532 -5818 11592 -5812
rect 9556 -5878 11532 -5818
rect 9496 -5884 9556 -5878
rect 11532 -5884 11592 -5878
rect 11874 -5816 11934 -5810
rect 14588 -5816 14648 -5810
rect 11934 -5876 14588 -5816
rect 11874 -5882 11934 -5876
rect 14588 -5882 14648 -5876
rect 19676 -5818 19736 -5812
rect 21712 -5818 21772 -5812
rect 19736 -5878 21712 -5818
rect 19676 -5884 19736 -5878
rect 3676 -5906 3736 -5900
rect 4698 -5906 4758 -5900
rect 3736 -5966 4698 -5906
rect 3676 -5972 3736 -5966
rect 4698 -5972 4758 -5966
rect 7044 -5916 7104 -5910
rect 19784 -5916 19844 -5878
rect 21712 -5884 21772 -5878
rect 7104 -5976 19844 -5916
rect 7044 -5982 7104 -5976
rect 3784 -6018 3844 -6012
rect 4568 -6018 4628 -6012
rect 3844 -6078 4568 -6018
rect 3784 -6084 3844 -6078
rect 4568 -6084 4628 -6078
rect 7180 -6014 7240 -6008
rect 9496 -6014 9556 -6008
rect 7240 -6074 9496 -6014
rect 7180 -6080 7240 -6074
rect 9496 -6080 9556 -6074
rect 10516 -6012 10576 -6006
rect 15606 -6012 15666 -6006
rect 22978 -6012 23038 -6006
rect 10576 -6072 15606 -6012
rect 15666 -6072 22978 -6012
rect 10516 -6078 10576 -6072
rect 15606 -6078 15666 -6072
rect 22978 -6078 23038 -6072
rect 8482 -6124 8542 -6118
rect 10516 -6124 10576 -6118
rect 8542 -6184 10516 -6124
rect 8482 -6190 8542 -6184
rect 10516 -6190 10576 -6184
rect 13572 -6126 13632 -6120
rect 15606 -6126 15666 -6120
rect 13632 -6186 15606 -6126
rect 13572 -6192 13632 -6186
rect 15606 -6192 15666 -6186
rect 18662 -6126 18722 -6120
rect 20696 -6124 20756 -6120
rect 20628 -6126 20756 -6124
rect 23290 -6126 23350 -6120
rect 18722 -6186 20696 -6126
rect 20756 -6186 23290 -6126
rect 18662 -6192 18722 -6186
rect 20628 -6188 20756 -6186
rect 20696 -6192 20756 -6188
rect 23290 -6192 23350 -6186
rect 2014 -6940 2074 -6934
rect 5208 -6940 5268 -6934
rect 2074 -7000 5208 -6940
rect 2014 -7006 2074 -7000
rect 5208 -7006 5268 -7000
rect 3174 -7050 3234 -7044
rect 6360 -7050 6420 -7044
rect 3234 -7110 6360 -7050
rect 19526 -7060 19586 -7054
rect 3174 -7116 3234 -7110
rect 6360 -7116 6420 -7110
rect 6802 -7074 6862 -7068
rect 13568 -7074 13628 -7068
rect 14588 -7074 14648 -7068
rect 16624 -7074 16684 -7068
rect 6862 -7134 13568 -7074
rect 13628 -7134 14588 -7074
rect 14648 -7134 16624 -7074
rect 19586 -7120 23948 -7060
rect 19526 -7126 19586 -7120
rect 6802 -7140 6862 -7134
rect 13568 -7140 13628 -7134
rect 14588 -7140 14648 -7134
rect 16624 -7140 16684 -7134
rect 19674 -7170 19734 -7164
rect 21714 -7170 21774 -7164
rect 22854 -7170 22914 -7164
rect 6552 -7178 6612 -7172
rect 11534 -7178 11594 -7172
rect 18658 -7178 18718 -7172
rect 6612 -7238 9498 -7178
rect 9558 -7238 11534 -7178
rect 11594 -7238 18658 -7178
rect 19734 -7230 21714 -7170
rect 21774 -7230 22854 -7170
rect 19674 -7236 19734 -7230
rect 21714 -7236 21774 -7230
rect 22854 -7236 22914 -7230
rect 6552 -7244 6612 -7238
rect 11534 -7244 11594 -7238
rect 18658 -7244 18718 -7238
rect 11532 -7280 11592 -7274
rect 20694 -7280 20754 -7274
rect 6798 -7288 6858 -7282
rect 7464 -7288 7524 -7282
rect 6858 -7348 7464 -7288
rect 11592 -7340 20694 -7280
rect 11532 -7346 11592 -7340
rect 20694 -7346 20754 -7340
rect 6798 -7354 6858 -7348
rect 7464 -7354 7524 -7348
rect 9498 -7382 9558 -7376
rect 11532 -7382 11592 -7376
rect 9558 -7442 11532 -7382
rect 9498 -7448 9558 -7442
rect 11532 -7448 11592 -7442
rect 14588 -7380 14648 -7374
rect 15606 -7380 15666 -7374
rect 16622 -7380 16682 -7374
rect 19526 -7380 19586 -7374
rect 14648 -7440 15606 -7380
rect 15666 -7440 16622 -7380
rect 16682 -7440 19526 -7380
rect 14588 -7446 14648 -7440
rect 15606 -7446 15666 -7440
rect 16622 -7446 16682 -7440
rect 19526 -7446 19586 -7440
rect 19678 -7378 19738 -7372
rect 21712 -7378 21772 -7372
rect 22978 -7378 23038 -7372
rect 19738 -7438 21712 -7378
rect 21772 -7438 22978 -7378
rect 23038 -7438 23820 -7378
rect 19678 -7444 19738 -7438
rect 21712 -7444 21772 -7438
rect 22978 -7444 23038 -7438
rect 3690 -7974 3750 -7968
rect 4700 -7974 4760 -7968
rect 1882 -8088 1888 -8028
rect 1948 -8088 1954 -8028
rect 3750 -8034 4700 -7974
rect 3690 -8040 3750 -8034
rect 4700 -8040 4760 -8034
rect 3796 -8074 3856 -8068
rect 4582 -8074 4642 -8068
rect 1396 -9144 1402 -9084
rect 1462 -9144 1468 -9084
rect 1276 -9644 1282 -9584
rect 1342 -9644 1348 -9584
rect 1282 -11494 1342 -9644
rect 1282 -11560 1342 -11554
rect 1402 -11492 1462 -9144
rect 1536 -9320 1542 -9260
rect 1602 -9320 1608 -9260
rect 1542 -11474 1602 -9320
rect 1764 -10142 1770 -10082
rect 1830 -10142 1836 -10082
rect 1770 -11458 1830 -10142
rect 1888 -11358 1948 -8088
rect 3856 -8134 4582 -8074
rect 3796 -8140 3856 -8134
rect 4582 -8140 4642 -8134
rect 11534 -8322 11594 -8316
rect 13336 -8322 13396 -8316
rect 6686 -8330 6746 -8324
rect 8480 -8330 8540 -8324
rect 10516 -8330 10576 -8324
rect 6746 -8390 8480 -8330
rect 8540 -8390 10516 -8330
rect 11594 -8382 13336 -8322
rect 11534 -8388 11594 -8382
rect 13336 -8388 13396 -8382
rect 13570 -8328 13630 -8322
rect 15606 -8328 15666 -8322
rect 13630 -8388 15606 -8328
rect 6686 -8396 6746 -8390
rect 2436 -9494 2442 -9434
rect 2502 -9494 2508 -9434
rect 2330 -9906 2336 -9846
rect 2396 -9906 2402 -9846
rect 2210 -10024 2216 -9964
rect 2276 -10024 2282 -9964
rect 2216 -11348 2276 -10024
rect 2336 -10940 2396 -9906
rect 2319 -10949 2409 -10940
rect 2319 -11048 2409 -11039
rect 1882 -11418 1888 -11358
rect 1948 -11418 1954 -11358
rect 2336 -11356 2396 -11048
rect 2216 -11414 2276 -11408
rect 2330 -11416 2336 -11356
rect 2396 -11416 2402 -11356
rect 2442 -11492 2502 -9494
rect 1770 -11524 1830 -11518
rect 1542 -11540 1602 -11534
rect 2436 -11552 2442 -11492
rect 2502 -11552 2508 -11492
rect 1402 -11558 1462 -11552
rect 1660 -11612 1720 -11606
rect 6914 -11612 6974 -8390
rect 8480 -8396 8540 -8390
rect 10516 -8396 10576 -8390
rect 13570 -8394 13630 -8388
rect 15606 -8394 15666 -8388
rect 18660 -8326 18720 -8320
rect 20696 -8326 20756 -8320
rect 18720 -8386 20696 -8326
rect 18660 -8392 18720 -8386
rect 20696 -8392 20756 -8386
rect 10516 -8438 10576 -8432
rect 15604 -8438 15664 -8432
rect 22854 -8438 22914 -8432
rect 10576 -8498 15604 -8438
rect 15664 -8498 22854 -8438
rect 10516 -8504 10576 -8498
rect 15604 -8504 15664 -8498
rect 22854 -8504 22914 -8498
rect 7312 -8538 7372 -8532
rect 7372 -8598 19896 -8538
rect 7312 -8604 7372 -8598
rect 9494 -8640 9554 -8634
rect 11528 -8640 11588 -8634
rect 9554 -8700 11528 -8640
rect 19682 -8640 19742 -8634
rect 19836 -8640 19896 -8598
rect 21716 -8640 21776 -8634
rect 9494 -8706 9554 -8700
rect 11528 -8706 11588 -8700
rect 11732 -8652 11792 -8646
rect 11792 -8712 15094 -8652
rect 15154 -8712 16110 -8652
rect 16170 -8712 19170 -8652
rect 19230 -8712 19236 -8652
rect 19742 -8700 21716 -8640
rect 19682 -8706 19742 -8700
rect 21716 -8706 21776 -8700
rect 11732 -8718 11792 -8712
rect 7044 -9588 7104 -9582
rect 8476 -9588 8536 -9582
rect 10512 -9588 10572 -9582
rect 7104 -9648 8476 -9588
rect 8536 -9648 10512 -9588
rect 7044 -9654 7104 -9648
rect 8476 -9654 8536 -9648
rect 10512 -9654 10572 -9648
rect 18664 -9588 18724 -9582
rect 20700 -9588 20760 -9582
rect 18724 -9648 20700 -9588
rect 18664 -9654 18724 -9648
rect 7180 -9718 7240 -9712
rect 18794 -9718 18854 -9648
rect 20700 -9654 20760 -9648
rect 7240 -9778 18854 -9718
rect 7180 -9784 7240 -9778
rect 11534 -9858 11594 -9852
rect 23138 -9858 23198 -9852
rect 11594 -9918 23138 -9858
rect 11534 -9924 11594 -9918
rect 1720 -11672 6974 -11612
rect 1660 -11678 1720 -11672
rect 1150 -11688 1210 -11682
rect 13254 -11842 13314 -9918
rect 13254 -11908 13314 -11902
rect 18358 -11842 18418 -9918
rect 22418 -11848 22478 -9918
rect 23138 -9924 23198 -9918
rect 18358 -11908 18418 -11902
rect 22412 -11908 22418 -11848
rect 22478 -11908 22484 -11848
rect -1562 -12220 -1502 -12214
rect 2216 -12220 2276 -12214
rect -1502 -12280 2216 -12220
rect -1562 -12286 -1502 -12280
rect 2216 -12286 2276 -12280
rect -36 -12354 24 -12348
rect 1770 -12354 1830 -12348
rect 24 -12414 1770 -12354
rect -36 -12420 24 -12414
rect 1770 -12420 1830 -12414
rect 2012 -13578 2072 -13572
rect 2072 -13638 3586 -13578
rect 3646 -13638 3652 -13578
rect 2012 -13644 2072 -13638
rect 4600 -13794 4660 -13788
rect 6640 -13794 6700 -13788
rect 8680 -13794 8740 -13788
rect 10710 -13794 10770 -13788
rect 12750 -13794 12810 -13788
rect 14782 -13794 14842 -13788
rect 16822 -13794 16882 -13788
rect 18858 -13794 18918 -13788
rect 20892 -13794 20952 -13788
rect 4660 -13854 6640 -13794
rect 6700 -13854 8680 -13794
rect 8740 -13854 10710 -13794
rect 10770 -13854 12750 -13794
rect 12810 -13854 14782 -13794
rect 14842 -13854 16822 -13794
rect 16882 -13854 18858 -13794
rect 18918 -13854 20892 -13794
rect 4600 -13860 4660 -13854
rect 6640 -13860 6700 -13854
rect 8680 -13860 8740 -13854
rect 10710 -13860 10770 -13854
rect 12750 -13860 12810 -13854
rect 14782 -13860 14842 -13854
rect 16822 -13860 16882 -13854
rect 18858 -13860 18918 -13854
rect 20892 -13860 20952 -13854
rect 2224 -13914 2284 -13908
rect 2568 -13914 2628 -13908
rect 2284 -13974 2568 -13914
rect 2224 -13980 2284 -13974
rect 2568 -13980 2628 -13974
rect 4092 -13920 4152 -13914
rect 12236 -13920 12296 -13914
rect 4152 -13980 5106 -13920
rect 5166 -13980 6128 -13920
rect 6188 -13980 7142 -13920
rect 7202 -13980 8168 -13920
rect 8228 -13980 9180 -13920
rect 9240 -13980 10216 -13920
rect 10276 -13980 11222 -13920
rect 11282 -13980 12236 -13920
rect 12296 -13980 13252 -13920
rect 13312 -13980 14260 -13920
rect 14320 -13980 15276 -13920
rect 15336 -13980 16300 -13920
rect 16360 -13980 17322 -13920
rect 17382 -13980 18344 -13920
rect 18404 -13980 19362 -13920
rect 19422 -13980 20376 -13920
rect 20436 -13980 21400 -13920
rect 21460 -13980 21466 -13920
rect 4092 -13986 4152 -13980
rect 12236 -13986 12296 -13980
rect 2442 -14036 2502 -14030
rect 7656 -14036 7716 -14030
rect 17844 -14036 17904 -14030
rect 21916 -14036 21976 -14030
rect 23048 -14036 23108 -14030
rect 2502 -14096 7656 -14036
rect 7716 -14096 17844 -14036
rect 17904 -14096 21916 -14036
rect 21976 -14096 23048 -14036
rect 2442 -14102 2502 -14096
rect 7656 -14102 7716 -14096
rect 17844 -14102 17904 -14096
rect 21916 -14102 21976 -14096
rect 23048 -14102 23108 -14096
rect 4604 -14958 4664 -14952
rect 6644 -14958 6704 -14952
rect 8676 -14958 8736 -14952
rect 10708 -14958 10768 -14952
rect 12744 -14958 12804 -14952
rect 14780 -14958 14840 -14952
rect 16818 -14958 16878 -14952
rect 18856 -14958 18916 -14952
rect 20892 -14958 20952 -14952
rect 4664 -15018 6644 -14958
rect 6704 -15018 8676 -14958
rect 8736 -15018 10708 -14958
rect 10768 -15018 12744 -14958
rect 12804 -15018 14780 -14958
rect 14840 -15018 16818 -14958
rect 16878 -15018 18856 -14958
rect 18916 -15018 20892 -14958
rect 4604 -15024 4664 -15018
rect 6644 -15024 6704 -15018
rect 8676 -15024 8736 -15018
rect 10708 -15024 10768 -15018
rect 12744 -15024 12804 -15018
rect 14780 -15024 14840 -15018
rect 16818 -15024 16878 -15018
rect 18856 -15024 18916 -15018
rect 20892 -15024 20952 -15018
rect 4096 -15068 4156 -15062
rect 5118 -15068 5178 -15062
rect 6132 -15068 6192 -15062
rect 7146 -15068 7206 -15062
rect 8164 -15068 8224 -15062
rect 9190 -15068 9250 -15062
rect 10210 -15068 10270 -15062
rect 11230 -15068 11290 -15062
rect 12232 -15068 12292 -15062
rect 13258 -15068 13318 -15062
rect 14276 -15068 14336 -15062
rect 15284 -15068 15344 -15062
rect 16296 -15068 16356 -15062
rect 17328 -15068 17388 -15062
rect 18342 -15068 18402 -15062
rect 19360 -15068 19420 -15062
rect 20384 -15068 20444 -15062
rect 21404 -15068 21464 -15062
rect 4156 -15128 5118 -15068
rect 5178 -15128 6132 -15068
rect 6192 -15128 7146 -15068
rect 7206 -15128 8164 -15068
rect 8224 -15128 9190 -15068
rect 9250 -15128 10210 -15068
rect 10270 -15128 11230 -15068
rect 11290 -15128 12232 -15068
rect 12292 -15128 13258 -15068
rect 13318 -15128 14276 -15068
rect 14336 -15128 15284 -15068
rect 15344 -15128 16296 -15068
rect 16356 -15128 17328 -15068
rect 17388 -15128 18342 -15068
rect 18402 -15128 19360 -15068
rect 19420 -15128 20384 -15068
rect 20444 -15128 21404 -15068
rect 4096 -15134 4156 -15128
rect 5118 -15134 5178 -15128
rect 6132 -15134 6192 -15128
rect 7146 -15134 7206 -15128
rect 8164 -15134 8224 -15128
rect 9190 -15134 9250 -15128
rect 10210 -15134 10270 -15128
rect 11230 -15134 11290 -15128
rect 12232 -15134 12292 -15128
rect 13258 -15134 13318 -15128
rect 14276 -15134 14336 -15128
rect 15284 -15134 15344 -15128
rect 16296 -15134 16356 -15128
rect 17328 -15134 17388 -15128
rect 18342 -15134 18402 -15128
rect 19360 -15134 19420 -15128
rect 20384 -15134 20444 -15128
rect 21404 -15134 21464 -15128
rect 2120 -15174 2180 -15168
rect 3586 -15174 3646 -15168
rect 5626 -15174 5686 -15168
rect 7656 -15174 7716 -15168
rect 9696 -15174 9756 -15168
rect 11730 -15174 11790 -15168
rect 13766 -15174 13826 -15168
rect 15802 -15174 15862 -15168
rect 17842 -15174 17902 -15168
rect 19872 -15174 19932 -15168
rect 21912 -15174 21972 -15168
rect 2180 -15234 3586 -15174
rect 3646 -15234 5626 -15174
rect 5686 -15234 7656 -15174
rect 7716 -15234 9696 -15174
rect 9756 -15234 11730 -15174
rect 11790 -15234 13766 -15174
rect 13826 -15234 15802 -15174
rect 15862 -15234 17842 -15174
rect 17902 -15234 19872 -15174
rect 19932 -15234 21912 -15174
rect 2120 -15240 2180 -15234
rect 3586 -15240 3646 -15234
rect 5626 -15240 5686 -15234
rect 7656 -15240 7716 -15234
rect 9696 -15240 9756 -15234
rect 11730 -15240 11790 -15234
rect 13766 -15240 13826 -15234
rect 15802 -15240 15862 -15234
rect 17842 -15240 17902 -15234
rect 19872 -15240 19932 -15234
rect 21912 -15240 21972 -15234
rect 2572 -15280 2632 -15274
rect 3070 -15280 3130 -15274
rect 3582 -15280 3642 -15274
rect 9862 -15280 9922 -15274
rect 11730 -15280 11790 -15274
rect 13768 -15280 13828 -15274
rect 15648 -15280 15708 -15274
rect 1880 -15340 1886 -15280
rect 1946 -15340 2572 -15280
rect 2632 -15340 3070 -15280
rect 3130 -15340 3582 -15280
rect 3642 -15340 9862 -15280
rect 9922 -15340 11730 -15280
rect 11790 -15340 13768 -15280
rect 13828 -15340 15648 -15280
rect 2572 -15346 2632 -15340
rect 3070 -15346 3130 -15340
rect 3582 -15346 3642 -15340
rect 9862 -15346 9922 -15340
rect 11730 -15346 11790 -15340
rect 13768 -15346 13828 -15340
rect 15648 -15346 15708 -15340
rect 19872 -15278 19932 -15272
rect 23048 -15278 23108 -15272
rect 19932 -15338 23048 -15278
rect 19872 -15344 19932 -15338
rect 23048 -15344 23108 -15338
rect 2442 -16170 2502 -16164
rect 5620 -16170 5680 -16164
rect 8676 -16170 8736 -16164
rect 14782 -16170 14842 -16164
rect 19876 -16170 19936 -16164
rect 2502 -16230 5620 -16170
rect 5680 -16230 8676 -16170
rect 8736 -16230 14782 -16170
rect 14842 -16230 19876 -16170
rect 2442 -16236 2502 -16230
rect 5620 -16236 5680 -16230
rect 8676 -16236 8736 -16230
rect 14782 -16236 14842 -16230
rect 19876 -16236 19936 -16230
rect 2012 -16274 2072 -16268
rect 2566 -16274 2626 -16268
rect 4086 -16274 4146 -16268
rect 2072 -16334 2566 -16274
rect 2626 -16334 4086 -16274
rect 2012 -16340 2072 -16334
rect 2566 -16340 2626 -16334
rect 4086 -16340 4146 -16334
rect 4598 -16274 4658 -16268
rect 5622 -16274 5682 -16268
rect 6634 -16274 6694 -16268
rect 7654 -16274 7714 -16268
rect 10712 -16274 10772 -16268
rect 12750 -16274 12810 -16268
rect 15800 -16274 15860 -16268
rect 16818 -16274 16878 -16268
rect 17838 -16274 17898 -16268
rect 18854 -16274 18914 -16268
rect 20890 -16274 20950 -16268
rect 4658 -16334 5622 -16274
rect 5682 -16334 6634 -16274
rect 6694 -16334 7654 -16274
rect 7714 -16334 10712 -16274
rect 10772 -16334 12750 -16274
rect 12810 -16334 15800 -16274
rect 15860 -16334 16818 -16274
rect 16878 -16334 17838 -16274
rect 17898 -16334 18854 -16274
rect 18914 -16334 20890 -16274
rect 4598 -16340 4658 -16334
rect 5622 -16340 5682 -16334
rect 6634 -16340 6694 -16334
rect 7654 -16340 7714 -16334
rect 10712 -16340 10772 -16334
rect 12750 -16340 12810 -16334
rect 15800 -16340 15860 -16334
rect 16818 -16340 16878 -16334
rect 17838 -16340 17898 -16334
rect 18854 -16340 18914 -16334
rect 20890 -16340 20950 -16334
rect 2336 -16396 2396 -16390
rect 9696 -16396 9756 -16390
rect 11730 -16396 11790 -16390
rect 13760 -16396 13820 -16390
rect 23760 -16396 23820 -7438
rect 2396 -16456 9696 -16396
rect 9756 -16456 11730 -16396
rect 11790 -16456 13760 -16396
rect 13820 -16456 23820 -16396
rect 2336 -16462 2396 -16456
rect 9696 -16462 9756 -16456
rect 11730 -16462 11790 -16456
rect 13760 -16462 13820 -16456
rect 2224 -16510 2284 -16504
rect 3072 -16510 3132 -16504
rect 2284 -16570 3072 -16510
rect 2224 -16576 2284 -16570
rect 3072 -16576 3132 -16570
rect 4604 -16508 4664 -16502
rect 6640 -16508 6700 -16502
rect 23034 -16508 23094 -16502
rect 4664 -16568 6640 -16508
rect 6700 -16568 23034 -16508
rect 4604 -16574 4664 -16568
rect 6640 -16574 6700 -16568
rect 23034 -16574 23094 -16568
rect 23162 -16526 23222 -16520
rect 23762 -16526 23822 -16520
rect 23222 -16586 23762 -16526
rect 23162 -16592 23222 -16586
rect 23762 -16592 23822 -16586
rect 22928 -17396 22988 -17390
rect 23888 -17396 23948 -7120
rect 5620 -17414 5680 -17408
rect 7656 -17414 7716 -17408
rect 15800 -17414 15860 -17408
rect 17836 -17414 17896 -17408
rect 21910 -17414 21970 -17408
rect 2448 -17438 2508 -17432
rect 3586 -17438 3646 -17432
rect 2508 -17498 3586 -17438
rect 3646 -17498 4468 -17438
rect 5680 -17474 7656 -17414
rect 7716 -17474 15800 -17414
rect 15860 -17474 17836 -17414
rect 17896 -17474 21910 -17414
rect 22988 -17456 23948 -17396
rect 22928 -17462 22988 -17456
rect 5620 -17480 5680 -17474
rect 7656 -17480 7716 -17474
rect 15800 -17480 15860 -17474
rect 17836 -17480 17896 -17474
rect 21910 -17480 21970 -17474
rect 2448 -17504 2508 -17498
rect 3586 -17504 3646 -17498
rect 2336 -17638 2396 -17632
rect 3584 -17638 3644 -17632
rect 2396 -17698 3584 -17638
rect 4408 -17634 4468 -17498
rect 4602 -17518 4662 -17512
rect 6642 -17518 6702 -17512
rect 8674 -17518 8734 -17512
rect 10708 -17518 10768 -17512
rect 12748 -17518 12808 -17512
rect 14782 -17518 14842 -17512
rect 4662 -17578 6642 -17518
rect 6702 -17578 8674 -17518
rect 8734 -17578 10708 -17518
rect 10768 -17578 12748 -17518
rect 12808 -17578 14782 -17518
rect 4602 -17584 4662 -17578
rect 6642 -17584 6702 -17578
rect 8674 -17584 8734 -17578
rect 10708 -17584 10768 -17578
rect 12748 -17584 12808 -17578
rect 14782 -17584 14842 -17578
rect 14978 -17522 15038 -17516
rect 19870 -17522 19930 -17516
rect 15038 -17582 19870 -17522
rect 23528 -17526 23588 -17520
rect 14978 -17588 15038 -17582
rect 19870 -17588 19930 -17582
rect 20368 -17586 20374 -17526
rect 20434 -17586 23528 -17526
rect 23528 -17592 23588 -17586
rect 5116 -17632 5176 -17626
rect 8674 -17630 8734 -17624
rect 10710 -17630 10770 -17624
rect 12746 -17630 12806 -17624
rect 14782 -17630 14842 -17624
rect 16816 -17630 16876 -17624
rect 18854 -17630 18914 -17624
rect 20894 -17630 20954 -17624
rect 23278 -17630 23338 -17624
rect 4408 -17692 5116 -17634
rect 5176 -17692 6120 -17632
rect 6180 -17692 7132 -17632
rect 7192 -17692 8152 -17632
rect 8212 -17692 8218 -17632
rect 8734 -17690 10710 -17630
rect 10770 -17690 12746 -17630
rect 12806 -17690 14782 -17630
rect 14842 -17690 16816 -17630
rect 16876 -17690 18854 -17630
rect 18914 -17690 20894 -17630
rect 20954 -17690 23278 -17630
rect 4408 -17694 5458 -17692
rect 5116 -17698 5176 -17694
rect 8674 -17696 8734 -17690
rect 10710 -17696 10770 -17690
rect 12746 -17696 12806 -17690
rect 14782 -17696 14842 -17690
rect 16816 -17696 16876 -17690
rect 18854 -17696 18914 -17690
rect 20894 -17696 20954 -17690
rect 23278 -17696 23338 -17690
rect 2336 -17704 2396 -17698
rect 3584 -17704 3644 -17698
rect 1660 -17740 1720 -17734
rect 2230 -17740 2290 -17734
rect 9692 -17740 9752 -17734
rect 11726 -17740 11786 -17734
rect 13766 -17740 13826 -17734
rect 14978 -17740 15038 -17734
rect 1720 -17800 2230 -17740
rect 2290 -17800 9692 -17740
rect 9752 -17800 11726 -17740
rect 11786 -17800 13766 -17740
rect 13826 -17800 14978 -17740
rect 1660 -17806 1720 -17800
rect 2230 -17806 2290 -17800
rect 9692 -17806 9752 -17800
rect 11726 -17806 11786 -17800
rect 13766 -17806 13826 -17800
rect 14978 -17806 15038 -17800
rect 15272 -17738 15332 -17732
rect 15332 -17798 16300 -17738
rect 16360 -17798 16366 -17738
rect 16818 -17744 16878 -17738
rect 18854 -17744 18914 -17738
rect 20892 -17744 20952 -17738
rect 23034 -17744 23094 -17738
rect 15272 -17804 15332 -17798
rect 16878 -17804 18854 -17744
rect 18914 -17804 20892 -17744
rect 20952 -17804 23034 -17744
rect 16818 -17810 16878 -17804
rect 18854 -17810 18914 -17804
rect 20892 -17810 20952 -17804
rect 23034 -17810 23094 -17804
rect 19366 -18658 19426 -18652
rect 3584 -18670 3644 -18664
rect 5622 -18670 5682 -18664
rect 7658 -18670 7718 -18664
rect 9690 -18670 9750 -18664
rect 3644 -18730 5622 -18670
rect 5682 -18730 7658 -18670
rect 7718 -18730 9690 -18670
rect 14266 -18718 14272 -18658
rect 14332 -18718 19366 -18658
rect 19366 -18724 19426 -18718
rect 19504 -18654 19564 -18648
rect 20386 -18654 20446 -18648
rect 21392 -18654 21452 -18648
rect 19564 -18714 20386 -18654
rect 20446 -18714 21392 -18654
rect 19504 -18720 19564 -18714
rect 20386 -18720 20446 -18714
rect 21392 -18720 21452 -18714
rect 21910 -18658 21970 -18652
rect 23162 -18658 23222 -18652
rect 21970 -18718 23162 -18658
rect 21910 -18724 21970 -18718
rect 23162 -18724 23222 -18718
rect 3584 -18736 3644 -18730
rect 5622 -18736 5682 -18730
rect 7658 -18736 7718 -18730
rect 9690 -18736 9750 -18730
rect 4090 -18772 4150 -18766
rect 9182 -18772 9242 -18766
rect 1150 -18822 1210 -18816
rect 4150 -18832 9182 -18772
rect 4090 -18838 4150 -18832
rect 9182 -18838 9242 -18832
rect 13766 -18786 13826 -18780
rect 21910 -18786 21970 -18780
rect 13826 -18846 21910 -18786
rect 13766 -18852 13826 -18846
rect 21910 -18852 21970 -18846
rect -3398 -19748 -3338 -19742
rect 1150 -19748 1210 -18882
rect 2336 -18874 2396 -18868
rect 5620 -18874 5680 -18868
rect 2396 -18934 5620 -18874
rect 2336 -18940 2396 -18934
rect 5620 -18940 5680 -18934
rect 6128 -18880 6188 -18874
rect 7150 -18880 7210 -18874
rect 8164 -18880 8224 -18874
rect 9182 -18880 9242 -18874
rect 10202 -18880 10262 -18874
rect 17314 -18880 17374 -18874
rect 18344 -18880 18404 -18874
rect 19504 -18880 19564 -18874
rect 6188 -18940 7150 -18880
rect 7210 -18940 8164 -18880
rect 8224 -18940 9182 -18880
rect 9242 -18940 10202 -18880
rect 10262 -18940 17314 -18880
rect 17374 -18940 18344 -18880
rect 18404 -18940 19504 -18880
rect 6128 -18946 6188 -18940
rect 7150 -18946 7210 -18940
rect 8164 -18946 8224 -18940
rect 9182 -18946 9242 -18940
rect 10202 -18946 10262 -18940
rect 17314 -18946 17374 -18940
rect 18344 -18946 18404 -18940
rect 19504 -18946 19564 -18940
rect 19872 -18880 19932 -18874
rect 23400 -18880 23460 -18874
rect 19932 -18940 23400 -18880
rect 19872 -18946 19932 -18940
rect 23400 -18946 23460 -18940
rect 4604 -18974 4664 -18968
rect 6638 -18974 6698 -18968
rect 8674 -18974 8734 -18968
rect 4664 -19034 6638 -18974
rect 6698 -19034 8674 -18974
rect 4604 -19040 4664 -19034
rect 6638 -19040 6698 -19034
rect 8674 -19040 8734 -19034
rect 15802 -18984 15862 -18978
rect 19872 -18984 19932 -18978
rect 15862 -19044 19872 -18984
rect 15802 -19050 15862 -19044
rect 19872 -19050 19932 -19044
rect 20888 -18982 20948 -18976
rect 23278 -18982 23338 -18976
rect 20948 -19042 23278 -18982
rect 20888 -19048 20948 -19042
rect 23278 -19048 23338 -19042
rect -3338 -19808 1210 -19748
rect -3398 -19814 -3338 -19808
rect -5428 -19894 -5368 -19888
rect -1368 -19894 -1308 -19888
rect 816 -19894 876 -19888
rect 1282 -19894 1342 -19888
rect 10710 -19892 10770 -19886
rect 12746 -19892 12806 -19886
rect 14782 -19892 14842 -19886
rect 16820 -19892 16880 -19886
rect -9514 -19954 -9508 -19894
rect -9448 -19954 -5428 -19894
rect -5368 -19954 -1368 -19894
rect -1308 -19954 816 -19894
rect 876 -19954 1282 -19894
rect -5428 -19960 -5368 -19954
rect -1368 -19960 -1308 -19954
rect 816 -19960 876 -19954
rect 1282 -19960 1342 -19954
rect 4086 -19898 4146 -19892
rect 4996 -19898 5056 -19892
rect 5998 -19898 6058 -19892
rect 7150 -19898 7210 -19892
rect 8160 -19898 8220 -19892
rect 9166 -19898 9226 -19892
rect 10210 -19898 10270 -19892
rect 4146 -19958 4996 -19898
rect 5056 -19958 5998 -19898
rect 6058 -19958 7150 -19898
rect 7210 -19958 8160 -19898
rect 8220 -19958 9166 -19898
rect 9226 -19958 10210 -19898
rect 10770 -19952 12746 -19892
rect 12806 -19952 14782 -19892
rect 14842 -19952 16820 -19892
rect 10710 -19958 10770 -19952
rect 12746 -19958 12806 -19952
rect 14782 -19958 14842 -19952
rect 16820 -19958 16880 -19952
rect 18856 -19892 18916 -19886
rect 20894 -19892 20954 -19886
rect 18916 -19952 20894 -19892
rect 18856 -19958 18916 -19952
rect 20894 -19958 20954 -19952
rect 4086 -19964 4146 -19958
rect 4996 -19964 5056 -19958
rect 5998 -19964 6058 -19958
rect 7150 -19964 7210 -19958
rect 8160 -19964 8220 -19958
rect 9166 -19964 9226 -19958
rect 10210 -19964 10270 -19958
rect 6638 -20000 6698 -19994
rect 16812 -20000 16872 -19994
rect 18852 -20000 18912 -19994
rect 20890 -20000 20950 -19994
rect -10662 -20022 -10602 -20016
rect -7984 -20022 -7924 -20016
rect -6952 -20022 -6892 -20016
rect -3892 -20022 -3832 -20016
rect -2896 -20022 -2836 -20016
rect 1402 -20022 1462 -20016
rect -10602 -20082 -7984 -20022
rect -7924 -20082 -6952 -20022
rect -6892 -20082 -3892 -20022
rect -3832 -20082 -2896 -20022
rect -2836 -20082 1402 -20022
rect 6698 -20060 16812 -20000
rect 16872 -20060 18852 -20000
rect 18912 -20060 20890 -20000
rect 6638 -20066 6698 -20060
rect 16812 -20066 16872 -20060
rect 18852 -20066 18912 -20060
rect 20890 -20066 20950 -20060
rect -10662 -20088 -10602 -20082
rect -7984 -20088 -7924 -20082
rect -6952 -20088 -6892 -20082
rect -3892 -20088 -3832 -20082
rect -2896 -20088 -2836 -20082
rect 1402 -20088 1462 -20082
rect 4086 -20114 4146 -20108
rect 6138 -20114 6198 -20108
rect 9164 -20114 9224 -20108
rect 10204 -20114 10264 -20108
rect 11218 -20114 11278 -20108
rect 12226 -20114 12286 -20108
rect 13270 -20114 13330 -20108
rect 14260 -20114 14320 -20108
rect 15278 -20114 15338 -20108
rect 16312 -20114 16372 -20108
rect 19344 -20114 19404 -20108
rect 20382 -20114 20442 -20108
rect 21408 -20114 21468 -20108
rect 4146 -20174 5124 -20114
rect 5184 -20174 6138 -20114
rect 6198 -20174 9164 -20114
rect 9224 -20174 10204 -20114
rect 10264 -20174 11218 -20114
rect 11278 -20174 12226 -20114
rect 12286 -20174 13270 -20114
rect 13330 -20174 14260 -20114
rect 14320 -20174 15278 -20114
rect 15338 -20174 16312 -20114
rect 16372 -20174 19344 -20114
rect 19404 -20174 20382 -20114
rect 20442 -20174 21408 -20114
rect 21468 -20174 23526 -20114
rect 23586 -20174 23592 -20114
rect 4086 -20180 4146 -20174
rect 6138 -20180 6198 -20174
rect 9164 -20180 9224 -20174
rect 10204 -20180 10264 -20174
rect 11218 -20180 11278 -20174
rect 12226 -20180 12286 -20174
rect 13270 -20180 13330 -20174
rect 14260 -20180 14320 -20174
rect 15278 -20180 15338 -20174
rect 16312 -20180 16372 -20174
rect 19344 -20180 19404 -20174
rect 20382 -20180 20442 -20174
rect 21408 -20180 21468 -20174
rect 9688 -20218 9748 -20212
rect 11730 -20218 11790 -20212
rect 13768 -20218 13828 -20212
rect 15802 -20218 15862 -20212
rect 17836 -20216 17896 -20210
rect 19870 -20216 19930 -20210
rect 21912 -20216 21972 -20210
rect 23162 -20216 23222 -20210
rect 2444 -20278 2450 -20218
rect 2510 -20278 9688 -20218
rect 9748 -20278 11730 -20218
rect 11790 -20278 13768 -20218
rect 13828 -20278 15802 -20218
rect 9688 -20284 9748 -20278
rect 11730 -20284 11790 -20278
rect 13768 -20284 13828 -20278
rect 15802 -20284 15862 -20278
rect 16314 -20222 16374 -20216
rect 17336 -20222 17396 -20216
rect 16374 -20282 17336 -20222
rect 17896 -20276 19870 -20216
rect 19930 -20276 21912 -20216
rect 21972 -20276 23162 -20216
rect 17836 -20282 17896 -20276
rect 19870 -20282 19930 -20276
rect 21912 -20282 21972 -20276
rect 23162 -20282 23222 -20276
rect 16314 -20288 16374 -20282
rect 17336 -20288 17396 -20282
rect -9004 -20984 -8944 -20978
rect -7980 -20984 -7920 -20978
rect -6948 -20984 -6888 -20978
rect -5948 -20984 -5888 -20978
rect -4928 -20984 -4868 -20978
rect -3908 -20984 -3848 -20978
rect -1884 -20984 -1824 -20978
rect 936 -20984 996 -20978
rect 1542 -20984 1602 -20978
rect -8944 -21044 -7980 -20984
rect -7920 -21044 -6948 -20984
rect -6888 -21044 -5948 -20984
rect -5888 -21044 -4928 -20984
rect -4868 -21044 -3908 -20984
rect -3848 -21044 -2898 -20984
rect -2838 -21044 -1884 -20984
rect -1824 -21044 -866 -20984
rect -806 -21044 936 -20984
rect 996 -21044 1542 -20984
rect -9004 -21050 -8944 -21044
rect -7980 -21050 -7920 -21044
rect -6948 -21050 -6888 -21044
rect -5948 -21050 -5888 -21044
rect -4928 -21050 -4868 -21044
rect -3908 -21050 -3848 -21044
rect -1884 -21050 -1824 -21044
rect 936 -21050 996 -21044
rect 1542 -21050 1602 -21044
rect -9504 -21088 -9444 -21082
rect -7468 -21088 -7408 -21082
rect -5432 -21088 -5372 -21082
rect -3398 -21088 -3338 -21082
rect -1362 -21088 -1302 -21082
rect -9444 -21148 -7468 -21088
rect -7408 -21148 -5432 -21088
rect -5372 -21148 -3398 -21088
rect -3338 -21148 -1362 -21088
rect 8678 -21120 8738 -21114
rect 12746 -21120 12806 -21114
rect 14780 -21120 14840 -21114
rect -9504 -21154 -9444 -21148
rect -7468 -21154 -7408 -21148
rect -5432 -21154 -5372 -21148
rect -3398 -21154 -3338 -21148
rect -1362 -21154 -1302 -21148
rect 4084 -21126 4144 -21120
rect 5092 -21126 5152 -21120
rect 6106 -21126 6166 -21120
rect 7144 -21126 7204 -21120
rect 8162 -21126 8222 -21120
rect 4144 -21186 5092 -21126
rect 5152 -21186 6106 -21126
rect 6166 -21186 7144 -21126
rect 7204 -21186 8162 -21126
rect 8738 -21180 10714 -21120
rect 10774 -21180 12746 -21120
rect 12806 -21180 14780 -21120
rect 8678 -21186 8738 -21180
rect 12746 -21186 12806 -21180
rect 14780 -21186 14840 -21180
rect 15802 -21118 15862 -21112
rect 16156 -21118 16216 -21112
rect 15862 -21178 16156 -21118
rect 15802 -21184 15862 -21178
rect 16156 -21184 16216 -21178
rect 19874 -21118 19934 -21112
rect 23158 -21118 23218 -21112
rect 19934 -21178 23158 -21118
rect 19874 -21184 19934 -21178
rect 23158 -21184 23218 -21178
rect -4418 -21192 -4358 -21186
rect 2120 -21192 2180 -21186
rect 4084 -21192 4144 -21186
rect 5092 -21192 5152 -21186
rect 6106 -21192 6166 -21186
rect 7144 -21192 7204 -21186
rect 8162 -21192 8222 -21186
rect -8492 -21252 -8486 -21192
rect -8426 -21252 -6450 -21192
rect -6390 -21252 -4418 -21192
rect -4358 -21252 -2384 -21192
rect -2324 -21252 -340 -21192
rect -280 -21252 2120 -21192
rect -4418 -21258 -4358 -21252
rect 2120 -21258 2180 -21252
rect 2230 -21230 2290 -21224
rect 3586 -21230 3646 -21224
rect 11730 -21230 11790 -21224
rect 13766 -21230 13826 -21224
rect 15798 -21230 15858 -21224
rect 2290 -21290 3586 -21230
rect 3646 -21290 11730 -21230
rect 11790 -21290 13766 -21230
rect 13826 -21290 15798 -21230
rect 2230 -21296 2290 -21290
rect 3586 -21296 3646 -21290
rect 11730 -21296 11790 -21290
rect 13766 -21296 13826 -21290
rect 15798 -21296 15858 -21290
rect 15308 -21328 15368 -21322
rect 16346 -21328 16406 -21322
rect 17322 -21328 17382 -21322
rect 18338 -21328 18398 -21322
rect 20364 -21328 20424 -21322
rect 21394 -21328 21454 -21322
rect 1888 -21342 1948 -21336
rect 4602 -21342 4662 -21336
rect 6640 -21342 6700 -21336
rect 10712 -21342 10772 -21336
rect 1948 -21402 4602 -21342
rect 4662 -21402 6640 -21342
rect 6700 -21402 10712 -21342
rect 15368 -21388 16346 -21328
rect 16406 -21388 17322 -21328
rect 17382 -21388 18338 -21328
rect 18398 -21388 20364 -21328
rect 20424 -21388 21394 -21328
rect 15308 -21394 15368 -21388
rect 16346 -21394 16406 -21388
rect 17322 -21394 17382 -21388
rect 18338 -21394 18398 -21388
rect 20364 -21394 20424 -21388
rect 21394 -21394 21454 -21388
rect 1888 -21408 1948 -21402
rect 4602 -21408 4662 -21402
rect 6640 -21408 6700 -21402
rect 10712 -21408 10772 -21402
rect 3582 -21440 3642 -21434
rect 5620 -21440 5680 -21434
rect 7660 -21440 7720 -21434
rect 9696 -21440 9756 -21434
rect 15800 -21440 15860 -21434
rect 16150 -21440 16156 -21436
rect 3642 -21500 5620 -21440
rect 5680 -21500 7660 -21440
rect 7720 -21500 9696 -21440
rect 9756 -21496 16156 -21440
rect 16216 -21440 16222 -21436
rect 17836 -21440 17896 -21434
rect 19872 -21440 19932 -21434
rect 21908 -21440 21968 -21434
rect 16216 -21496 17836 -21440
rect 9756 -21500 17836 -21496
rect 17896 -21500 19872 -21440
rect 19932 -21500 21908 -21440
rect 3582 -21506 3642 -21500
rect 5620 -21506 5680 -21500
rect 7660 -21506 7720 -21500
rect 9696 -21506 9756 -21500
rect 15800 -21506 15860 -21500
rect 17836 -21506 17896 -21500
rect 19872 -21506 19932 -21500
rect 21908 -21506 21968 -21500
rect -7474 -22134 -7414 -22128
rect -3398 -22134 -3338 -22128
rect 816 -22134 876 -22128
rect -7414 -22194 -3398 -22134
rect -3338 -22194 816 -22134
rect -7474 -22200 -7414 -22194
rect -3398 -22200 -3338 -22194
rect 816 -22200 876 -22194
rect -10662 -22254 -10602 -22248
rect -9012 -22254 -8952 -22248
rect -5942 -22254 -5882 -22248
rect -4934 -22254 -4874 -22248
rect -1872 -22254 -1812 -22248
rect -846 -22254 -786 -22248
rect -10602 -22314 -9012 -22254
rect -8952 -22314 -5942 -22254
rect -5882 -22314 -4934 -22254
rect -4874 -22314 -1872 -22254
rect -1812 -22314 -846 -22254
rect -10662 -22320 -10602 -22314
rect -9012 -22320 -8952 -22314
rect -5942 -22320 -5882 -22314
rect -4934 -22320 -4874 -22314
rect -1872 -22320 -1812 -22314
rect -846 -22320 -786 -22314
rect 10708 -22344 10768 -22338
rect 12750 -22344 12810 -22338
rect 14782 -22344 14842 -22338
rect 16822 -22344 16882 -22338
rect 23278 -22344 23338 -22338
rect 4602 -22364 4662 -22358
rect 6638 -22364 6698 -22358
rect 8676 -22364 8736 -22358
rect 4662 -22424 6638 -22364
rect 6698 -22424 8676 -22364
rect 10532 -22404 10538 -22344
rect 10598 -22404 10708 -22344
rect 10768 -22404 12750 -22344
rect 12810 -22404 14782 -22344
rect 14842 -22404 16822 -22344
rect 16882 -22404 23278 -22344
rect 10708 -22410 10768 -22404
rect 12750 -22410 12810 -22404
rect 14782 -22410 14842 -22404
rect 16822 -22410 16882 -22404
rect 23278 -22410 23338 -22404
rect 4602 -22430 4662 -22424
rect 6638 -22430 6698 -22424
rect 8676 -22430 8736 -22424
rect 15800 -22442 15860 -22436
rect 21906 -22442 21966 -22436
rect 23158 -22442 23218 -22436
rect 2448 -22462 2508 -22456
rect 5620 -22462 5680 -22456
rect 2508 -22522 5620 -22462
rect 2448 -22528 2508 -22522
rect 5620 -22528 5680 -22522
rect 7144 -22462 7204 -22456
rect 10192 -22462 10252 -22456
rect 7204 -22522 8166 -22462
rect 8226 -22522 9188 -22462
rect 9248 -22522 10192 -22462
rect 15860 -22502 21906 -22442
rect 21966 -22502 23158 -22442
rect 15800 -22508 15860 -22502
rect 21906 -22508 21966 -22502
rect 23158 -22508 23218 -22502
rect 7144 -22528 7204 -22522
rect 10192 -22528 10252 -22522
rect 10714 -22552 10774 -22546
rect 12742 -22552 12802 -22546
rect 14786 -22552 14846 -22546
rect 16814 -22552 16874 -22546
rect 18852 -22552 18912 -22546
rect 20892 -22552 20952 -22546
rect 4606 -22558 4666 -22552
rect 6642 -22558 6702 -22552
rect 8670 -22558 8730 -22552
rect 10538 -22558 10598 -22552
rect 4666 -22618 6642 -22558
rect 6702 -22618 8670 -22558
rect 8730 -22618 10538 -22558
rect 10774 -22612 12742 -22552
rect 12802 -22612 14786 -22552
rect 14846 -22612 16814 -22552
rect 16874 -22612 18852 -22552
rect 18912 -22612 20892 -22552
rect 10714 -22618 10774 -22612
rect 12742 -22618 12802 -22612
rect 14786 -22618 14846 -22612
rect 16814 -22618 16874 -22612
rect 18852 -22618 18912 -22612
rect 20892 -22618 20952 -22612
rect 21410 -22548 21470 -22542
rect 22922 -22548 22982 -22542
rect 23528 -22548 23588 -22542
rect 21470 -22608 22922 -22548
rect 22982 -22608 23528 -22548
rect 21410 -22614 21470 -22608
rect 22922 -22614 22982 -22608
rect 23528 -22614 23588 -22608
rect 4606 -22624 4666 -22618
rect 6642 -22624 6702 -22618
rect 8670 -22624 8730 -22618
rect 10538 -22624 10598 -22618
rect 3588 -22678 3648 -22672
rect 7656 -22678 7716 -22672
rect 9690 -22678 9750 -22672
rect 17840 -22678 17900 -22672
rect 19870 -22678 19930 -22672
rect 21910 -22676 21970 -22670
rect 23400 -22676 23460 -22670
rect 3648 -22738 7656 -22678
rect 7716 -22738 9690 -22678
rect 9750 -22738 17840 -22678
rect 17900 -22738 19870 -22678
rect 20390 -22736 20396 -22676
rect 20456 -22736 21910 -22676
rect 21970 -22736 23400 -22676
rect 3588 -22744 3648 -22738
rect 7656 -22744 7716 -22738
rect 9690 -22744 9750 -22738
rect 17840 -22744 17900 -22738
rect 19870 -22744 19930 -22738
rect 21910 -22742 21970 -22736
rect 23400 -22742 23460 -22736
rect -340 -23198 -280 -23192
rect -8492 -23258 -8486 -23198
rect -8426 -23258 -6450 -23198
rect -6390 -23258 -4418 -23198
rect -4358 -23258 -2384 -23198
rect -2324 -23258 -340 -23198
rect -340 -23264 -280 -23258
rect -9500 -23306 -9440 -23300
rect -7464 -23306 -7404 -23300
rect -5428 -23306 -5368 -23300
rect -3394 -23306 -3334 -23300
rect -1358 -23306 -1298 -23300
rect -9440 -23366 -7464 -23306
rect -7404 -23366 -5428 -23306
rect -5368 -23366 -3394 -23306
rect -3334 -23366 -1358 -23306
rect -9500 -23372 -9440 -23366
rect -7464 -23372 -7404 -23366
rect -5428 -23372 -5368 -23366
rect -3394 -23372 -3334 -23366
rect -1358 -23372 -1298 -23366
rect -9006 -23418 -8946 -23412
rect -7982 -23418 -7922 -23412
rect -6950 -23418 -6890 -23412
rect -5950 -23418 -5890 -23412
rect -4930 -23418 -4870 -23412
rect -3910 -23418 -3850 -23412
rect -1886 -23418 -1826 -23412
rect 936 -23418 996 -23412
rect -8946 -23478 -7982 -23418
rect -7922 -23478 -6950 -23418
rect -6890 -23478 -5950 -23418
rect -5890 -23478 -4930 -23418
rect -4870 -23478 -3910 -23418
rect -3850 -23478 -2900 -23418
rect -2840 -23478 -1886 -23418
rect -1826 -23478 -868 -23418
rect -808 -23478 936 -23418
rect -9006 -23484 -8946 -23478
rect -7982 -23484 -7922 -23478
rect -6950 -23484 -6890 -23478
rect -5950 -23484 -5890 -23478
rect -4930 -23484 -4870 -23478
rect -3910 -23484 -3850 -23478
rect -1886 -23484 -1826 -23478
rect 936 -23484 996 -23478
rect 2336 -23594 2396 -23588
rect 11724 -23594 11784 -23588
rect 13766 -23594 13826 -23588
rect 15802 -23594 15862 -23588
rect 2396 -23654 11724 -23594
rect 11784 -23654 13766 -23594
rect 13826 -23654 15802 -23594
rect 2336 -23660 2396 -23654
rect 11724 -23660 11784 -23654
rect 13766 -23660 13826 -23654
rect 15802 -23660 15862 -23654
rect 18856 -23594 18916 -23588
rect 20888 -23594 20948 -23588
rect 23034 -23594 23094 -23588
rect 18916 -23654 20888 -23594
rect 20948 -23654 23034 -23594
rect 18856 -23660 18916 -23654
rect 20888 -23660 20948 -23654
rect 23034 -23660 23094 -23654
rect 6140 -23708 6200 -23702
rect 11220 -23708 11280 -23702
rect 2230 -23720 2290 -23714
rect 5620 -23720 5680 -23714
rect 2290 -23780 5620 -23720
rect 6200 -23768 11220 -23708
rect 6140 -23774 6200 -23768
rect 11220 -23774 11280 -23768
rect 16308 -23704 16368 -23698
rect 21408 -23704 21468 -23698
rect 16368 -23764 21408 -23704
rect 16308 -23770 16368 -23764
rect 21408 -23770 21468 -23764
rect 22416 -23704 22476 -23698
rect 23650 -23704 23710 -23698
rect 22476 -23764 23650 -23704
rect 22416 -23770 22476 -23764
rect 23650 -23770 23710 -23764
rect 2230 -23786 2290 -23780
rect 5620 -23786 5680 -23780
rect 4602 -23822 4662 -23816
rect 6638 -23822 6698 -23816
rect 7658 -23822 7718 -23816
rect 8674 -23822 8734 -23816
rect 9694 -23822 9754 -23816
rect 10712 -23822 10772 -23816
rect 12742 -23822 12802 -23816
rect 14780 -23822 14840 -23816
rect 16816 -23822 16876 -23816
rect 17838 -23822 17898 -23816
rect 18858 -23822 18918 -23816
rect 19872 -23822 19932 -23816
rect 20894 -23822 20954 -23816
rect 4662 -23882 6638 -23822
rect 6698 -23882 7658 -23822
rect 7718 -23882 8674 -23822
rect 8734 -23882 9694 -23822
rect 9754 -23882 10712 -23822
rect 10772 -23882 12742 -23822
rect 12802 -23882 14780 -23822
rect 14840 -23882 16816 -23822
rect 16876 -23882 17838 -23822
rect 17898 -23882 18858 -23822
rect 18918 -23882 19872 -23822
rect 19932 -23882 20894 -23822
rect 4602 -23888 4662 -23882
rect 6638 -23888 6698 -23882
rect 7658 -23888 7718 -23882
rect 8674 -23888 8734 -23882
rect 9694 -23888 9754 -23882
rect 10712 -23888 10772 -23882
rect 12742 -23888 12802 -23882
rect 14780 -23888 14840 -23882
rect 16816 -23888 16876 -23882
rect 17838 -23888 17898 -23882
rect 18858 -23888 18918 -23882
rect 19872 -23888 19932 -23882
rect 20894 -23888 20954 -23882
rect 5620 -23926 5680 -23920
rect 10556 -23926 10616 -23920
rect 16962 -23926 17022 -23920
rect 19872 -23926 19932 -23920
rect 23054 -23926 23114 -23920
rect 5680 -23986 10556 -23926
rect 10616 -23986 16962 -23926
rect 17022 -23986 19872 -23926
rect 19932 -23986 23054 -23926
rect 5620 -23992 5680 -23986
rect 10556 -23992 10616 -23986
rect 16962 -23992 17022 -23986
rect 19872 -23992 19932 -23986
rect 23054 -23992 23114 -23986
rect -10662 -24380 -10602 -24374
rect -7992 -24380 -7932 -24374
rect -6960 -24380 -6900 -24374
rect -3900 -24380 -3840 -24374
rect -2904 -24380 -2844 -24374
rect -10602 -24440 -7992 -24380
rect -7932 -24440 -6960 -24380
rect -6900 -24440 -3900 -24380
rect -3840 -24440 -2904 -24380
rect -10662 -24446 -10602 -24440
rect -7992 -24446 -7932 -24440
rect -6960 -24446 -6900 -24440
rect -3900 -24446 -3840 -24440
rect -2904 -24446 -2844 -24440
rect -5426 -24510 -5366 -24504
rect -1366 -24510 -1306 -24504
rect 816 -24510 876 -24504
rect -9512 -24570 -9506 -24510
rect -9446 -24570 -5426 -24510
rect -5366 -24570 -1366 -24510
rect -1306 -24570 816 -24510
rect -5426 -24576 -5366 -24570
rect -1366 -24576 -1306 -24570
rect 816 -24576 876 -24570
rect 2448 -24824 2508 -24818
rect 5618 -24824 5678 -24818
rect 2508 -24884 5618 -24824
rect 2448 -24890 2508 -24884
rect 5618 -24890 5678 -24884
rect 9848 -24822 9908 -24816
rect 11726 -24822 11786 -24816
rect 13764 -24822 13824 -24816
rect 15634 -24822 15694 -24816
rect 21910 -24822 21970 -24816
rect 9908 -24882 11726 -24822
rect 11786 -24882 13764 -24822
rect 13824 -24882 15634 -24822
rect 15694 -24882 21910 -24822
rect 9848 -24888 9908 -24882
rect 11726 -24888 11786 -24882
rect 13764 -24888 13824 -24882
rect 15634 -24888 15694 -24882
rect 21910 -24888 21970 -24882
rect 2120 -24928 2180 -24922
rect 3584 -24928 3644 -24922
rect 5624 -24928 5684 -24922
rect 7654 -24928 7714 -24922
rect 9694 -24928 9754 -24922
rect 11730 -24928 11790 -24922
rect 13766 -24928 13826 -24922
rect 15800 -24928 15860 -24922
rect 17840 -24928 17900 -24922
rect 19870 -24928 19930 -24922
rect 21910 -24928 21970 -24922
rect 23762 -24928 23822 -24922
rect 2180 -24988 3584 -24928
rect 3644 -24988 5624 -24928
rect 5684 -24988 7654 -24928
rect 7714 -24988 9694 -24928
rect 9754 -24988 11730 -24928
rect 11790 -24988 13766 -24928
rect 13826 -24988 15800 -24928
rect 15860 -24988 17840 -24928
rect 17900 -24988 19870 -24928
rect 19930 -24988 21910 -24928
rect 21970 -24988 23762 -24928
rect 2120 -24994 2180 -24988
rect 3584 -24994 3644 -24988
rect 5624 -24994 5684 -24988
rect 7654 -24994 7714 -24988
rect 9694 -24994 9754 -24988
rect 11730 -24994 11790 -24988
rect 13766 -24994 13826 -24988
rect 15800 -24994 15860 -24988
rect 17840 -24994 17900 -24988
rect 19870 -24994 19930 -24988
rect 21910 -24994 21970 -24988
rect 23762 -24994 23822 -24988
rect 4092 -25034 4152 -25028
rect 5112 -25034 5172 -25028
rect 6136 -25034 6196 -25028
rect 7154 -25034 7214 -25028
rect 8168 -25034 8228 -25028
rect 9200 -25034 9260 -25028
rect 10212 -25034 10272 -25028
rect 11220 -25034 11280 -25028
rect 12238 -25034 12298 -25028
rect 13264 -25034 13324 -25028
rect 14266 -25034 14326 -25028
rect 15286 -25034 15346 -25028
rect 16306 -25034 16366 -25028
rect 17332 -25034 17392 -25028
rect 18350 -25034 18410 -25028
rect 19364 -25034 19424 -25028
rect 20378 -25034 20438 -25028
rect 21400 -25034 21460 -25028
rect 4152 -25094 5112 -25034
rect 5172 -25094 6136 -25034
rect 6196 -25094 7154 -25034
rect 7214 -25094 8168 -25034
rect 8228 -25094 9200 -25034
rect 9260 -25094 10212 -25034
rect 10272 -25094 11220 -25034
rect 11280 -25094 12238 -25034
rect 12298 -25094 13264 -25034
rect 13324 -25094 14266 -25034
rect 14326 -25094 15286 -25034
rect 15346 -25094 16306 -25034
rect 16366 -25094 17332 -25034
rect 17392 -25094 18350 -25034
rect 18410 -25094 19364 -25034
rect 19424 -25094 20378 -25034
rect 20438 -25094 21400 -25034
rect 4092 -25100 4152 -25094
rect 5112 -25100 5172 -25094
rect 6136 -25100 6196 -25094
rect 7154 -25100 7214 -25094
rect 8168 -25100 8228 -25094
rect 9200 -25100 9260 -25094
rect 10212 -25100 10272 -25094
rect 11220 -25100 11280 -25094
rect 12238 -25100 12298 -25094
rect 13264 -25100 13324 -25094
rect 14266 -25100 14326 -25094
rect 15286 -25100 15346 -25094
rect 16306 -25100 16366 -25094
rect 17332 -25100 17392 -25094
rect 18350 -25100 18410 -25094
rect 19364 -25100 19424 -25094
rect 20378 -25100 20438 -25094
rect 21400 -25100 21460 -25094
rect 4604 -25144 4664 -25138
rect 6640 -25144 6700 -25138
rect 8678 -25144 8738 -25138
rect 10716 -25144 10776 -25138
rect 12752 -25144 12812 -25138
rect 14788 -25144 14848 -25138
rect 16820 -25144 16880 -25138
rect 18852 -25144 18912 -25138
rect 20892 -25144 20952 -25138
rect 4664 -25204 6640 -25144
rect 6700 -25204 8678 -25144
rect 8738 -25204 10716 -25144
rect 10776 -25204 12752 -25144
rect 12812 -25204 14788 -25144
rect 14848 -25204 16820 -25144
rect 16880 -25204 18852 -25144
rect 18912 -25204 20892 -25144
rect 4604 -25210 4664 -25204
rect 6640 -25210 6700 -25204
rect 8678 -25210 8738 -25204
rect 10716 -25210 10776 -25204
rect 12752 -25210 12812 -25204
rect 14788 -25210 14848 -25204
rect 16820 -25210 16880 -25204
rect 18852 -25210 18912 -25204
rect 20892 -25210 20952 -25204
rect -8028 -25876 -7968 -25870
rect -5990 -25876 -5930 -25870
rect -3954 -25876 -3894 -25870
rect -1918 -25876 -1858 -25870
rect -7968 -25936 -5990 -25876
rect -5930 -25936 -3954 -25876
rect -3894 -25936 -1918 -25876
rect -8028 -25942 -7968 -25936
rect -5990 -25942 -5930 -25936
rect -3954 -25942 -3894 -25936
rect -1918 -25942 -1858 -25936
rect -7010 -25988 -6950 -25982
rect -2936 -25988 -2876 -25982
rect 1070 -25988 1130 -25982
rect -6950 -26048 -2936 -25988
rect -2876 -26048 1070 -25988
rect -7010 -26054 -6950 -26048
rect -2936 -26054 -2876 -26048
rect 1070 -26054 1130 -26048
rect 2448 -26066 2508 -26060
rect 3584 -26066 3644 -26060
rect 7654 -26066 7714 -26060
rect 17834 -26066 17894 -26060
rect 23054 -26066 23114 -26060
rect 2508 -26126 3584 -26066
rect 3644 -26126 7654 -26066
rect 7714 -26126 17834 -26066
rect 17894 -26126 23054 -26066
rect 2448 -26132 2508 -26126
rect 3584 -26132 3644 -26126
rect 7654 -26132 7714 -26126
rect 17834 -26132 17894 -26126
rect 23054 -26132 23114 -26126
rect 4096 -26174 4156 -26168
rect 12240 -26174 12300 -26168
rect 4156 -26234 5110 -26174
rect 5170 -26234 6132 -26174
rect 6192 -26234 7146 -26174
rect 7206 -26234 8172 -26174
rect 8232 -26234 9184 -26174
rect 9244 -26234 10220 -26174
rect 10280 -26234 11226 -26174
rect 11286 -26234 12240 -26174
rect 12300 -26234 13256 -26174
rect 13316 -26234 14264 -26174
rect 14324 -26234 15280 -26174
rect 15340 -26234 16304 -26174
rect 16364 -26234 17326 -26174
rect 17386 -26234 18348 -26174
rect 18408 -26234 19366 -26174
rect 19426 -26234 20380 -26174
rect 20440 -26234 21404 -26174
rect 21464 -26234 21470 -26174
rect 4096 -26240 4156 -26234
rect 12240 -26240 12300 -26234
rect -8118 -26476 23968 -26430
rect -8118 -26630 -8072 -26476
rect 23928 -26630 23968 -26476
rect -8118 -26676 23968 -26630
rect -12216 -26816 -11616 -26806
rect -12216 -27126 -11616 -27116
rect 24216 -26816 24816 -26806
rect 24216 -27126 24816 -27116
<< via2 >>
rect 484 3916 1084 4216
rect 24116 3916 24716 4216
rect 4061 3620 20846 3834
rect -13630 -10670 -2866 -10378
rect -2866 -10670 -2778 -10378
rect 2319 -11039 2409 -10949
rect -8072 -26630 23928 -26476
rect -12216 -27116 -11616 -26816
rect 24216 -27116 24816 -26816
<< metal3 >>
rect 474 4216 1094 4221
rect 474 3916 484 4216
rect 1084 3916 1094 4216
rect 474 3911 1094 3916
rect 24106 4216 24726 4221
rect 24106 3916 24116 4216
rect 24716 3916 24726 4216
rect 24106 3911 24726 3916
rect 3998 3834 20878 3866
rect 3998 3620 4061 3834
rect 20846 3620 20878 3834
rect 3998 3600 20878 3620
rect 3998 3598 8352 3600
rect -15168 2940 -128 3086
rect -15168 2930 -974 2940
rect -15168 2240 -15016 2930
rect -14320 2242 -974 2930
rect -284 2242 -128 2940
rect -14320 2240 -128 2242
rect -15168 1910 -128 2240
rect -15168 -10752 -13986 1910
rect -13698 -9290 -1792 1650
rect -1428 -9290 -128 1910
rect -13698 -10378 -128 -9290
rect -2778 -10670 -128 -10378
rect -2866 -10752 -128 -10670
rect -15168 -10978 -128 -10752
rect 2315 -10944 2413 -10939
rect 2314 -10945 2414 -10944
rect -15168 -11078 -1626 -10978
rect 2314 -11043 2315 -10945
rect 2413 -11043 2414 -10945
rect 2314 -11044 2414 -11043
rect 2315 -11049 2413 -11044
rect -15168 -11760 -15014 -11078
rect -14680 -11760 -1626 -11078
rect -15168 -11916 -1626 -11760
rect -8118 -26476 23968 -26430
rect -8118 -26630 -8072 -26476
rect 23928 -26630 23968 -26476
rect -8118 -26676 23968 -26630
rect -12226 -26816 -11606 -26811
rect -12226 -27116 -12216 -26816
rect -11616 -27116 -11606 -26816
rect -12226 -27121 -11606 -27116
rect 24206 -26816 24826 -26811
rect 24206 -27116 24216 -26816
rect 24816 -27116 24826 -26816
rect 24206 -27121 24826 -27116
<< via3 >>
rect 484 3916 1084 4216
rect 24116 3916 24716 4216
rect 4061 3620 20846 3834
rect -15016 2240 -14320 2930
rect -974 2242 -284 2940
rect -13986 1650 -1428 1910
rect -13986 -10378 -13698 1650
rect -1792 -9290 -1428 1650
rect -13986 -10670 -13630 -10378
rect -13630 -10670 -2866 -10378
rect -13986 -10752 -2866 -10670
rect 2315 -10949 2413 -10945
rect 2315 -11039 2319 -10949
rect 2319 -11039 2409 -10949
rect 2409 -11039 2413 -10949
rect 2315 -11043 2413 -11039
rect -15014 -11760 -14680 -11078
rect -8072 -26630 23928 -26476
rect -12216 -27116 -11616 -26816
rect 24216 -27116 24816 -26816
<< mimcap >>
rect -13982 2936 -7782 2986
rect -13982 2636 -8132 2936
rect -7832 2636 -7782 2936
rect -13982 2586 -7782 2636
rect -7582 2936 -1382 2986
rect -7582 2636 -1732 2936
rect -1432 2636 -1382 2936
rect -7582 2586 -1382 2636
rect -15068 1854 -14268 1904
rect -15068 -3846 -14618 1854
rect -14318 -3846 -14268 1854
rect -1024 1854 -224 1904
rect -13128 936 -7928 986
rect -13128 -3764 -8278 936
rect -7978 -3764 -7928 936
rect -13128 -3814 -7928 -3764
rect -7528 936 -2328 986
rect -7528 -3764 -2678 936
rect -2378 -3764 -2328 936
rect -7528 -3814 -2328 -3764
rect -15068 -3896 -14268 -3846
rect -1024 -3846 -574 1854
rect -274 -3846 -224 1854
rect -1024 -3896 -224 -3846
rect -15068 -4638 -14268 -4588
rect -15068 -10338 -14618 -4638
rect -14318 -10338 -14268 -4638
rect -13128 -4664 -7928 -4614
rect -13128 -9364 -8278 -4664
rect -7978 -9364 -7928 -4664
rect -13128 -9414 -7928 -9364
rect -7528 -4664 -2328 -4614
rect -7528 -9364 -2678 -4664
rect -2378 -9364 -2328 -4664
rect -7528 -9414 -2328 -9364
rect -1024 -4638 -224 -4588
rect -15068 -10388 -14268 -10338
rect -1024 -10338 -574 -4638
rect -274 -10338 -224 -4638
rect -1024 -10388 -224 -10338
rect -14482 -11064 -8282 -11014
rect -14482 -11364 -8632 -11064
rect -8332 -11364 -8282 -11064
rect -14482 -11414 -8282 -11364
rect -8082 -11064 -1882 -11014
rect -8082 -11364 -2232 -11064
rect -1932 -11364 -1882 -11064
rect -8082 -11414 -1882 -11364
<< mimcapcontact >>
rect -8132 2636 -7832 2936
rect -1732 2636 -1432 2936
rect -14618 -3846 -14318 1854
rect -8278 -3764 -7978 936
rect -2678 -3764 -2378 936
rect -574 -3846 -274 1854
rect -14618 -10338 -14318 -4638
rect -8278 -9364 -7978 -4664
rect -2678 -9364 -2378 -4664
rect -574 -10338 -274 -4638
rect -8632 -11364 -8332 -11064
rect -2232 -11364 -1932 -11064
<< metal4 >>
rect -15168 4216 25000 4400
rect -15168 3916 484 4216
rect 1084 3916 24116 4216
rect 24716 3916 25000 4216
rect -15168 3834 25000 3916
rect -15168 3620 4061 3834
rect 20846 3620 25000 3834
rect -15168 3600 25000 3620
rect -15168 2940 -128 3086
rect -15168 2936 -974 2940
rect -15168 2930 -8132 2936
rect -15168 2240 -15016 2930
rect -14320 2636 -8132 2930
rect -7832 2636 -1732 2936
rect -1432 2636 -974 2936
rect -14320 2242 -974 2636
rect -284 2242 -128 2940
rect -14320 2240 -128 2242
rect -15168 1910 -128 2240
rect -15168 1854 -13986 1910
rect -15168 -3846 -14618 1854
rect -14318 -3846 -13986 1854
rect -1428 1854 -128 1910
rect -15168 -4638 -13986 -3846
rect -15168 -10338 -14618 -4638
rect -14318 -10338 -13986 -4638
rect -15168 -10752 -13986 -10338
rect -13228 936 -2228 1086
rect -13228 -3764 -8278 936
rect -7978 -3764 -2678 936
rect -2378 -3764 -2228 936
rect -13228 -4664 -2228 -3764
rect -13228 -9364 -8278 -4664
rect -7978 -9364 -2678 -4664
rect -2378 -9364 -2228 -4664
rect -13228 -9816 -2228 -9364
rect -1428 -3846 -574 1854
rect -274 -3846 -128 1854
rect -1428 -4638 -128 -3846
rect -1428 -9436 -574 -4638
rect -13228 -9913 -1327 -9816
rect -13228 -9914 -2228 -9913
rect -13498 -10378 -2722 -10296
rect -2834 -10752 -2722 -10378
rect -15168 -10838 -2722 -10752
rect -15166 -10978 -2722 -10838
rect -15166 -11064 -1722 -10978
rect -15166 -11078 -8632 -11064
rect -15166 -11760 -15014 -11078
rect -14680 -11364 -8632 -11078
rect -8332 -11364 -2232 -11064
rect -1932 -11364 -1722 -11064
rect -14680 -11760 -1722 -11364
rect -1424 -11400 -1327 -9913
rect -1058 -10338 -574 -9436
rect -274 -10338 -128 -4638
rect -1058 -10848 -128 -10338
rect 226 -10945 2414 -10944
rect 226 -11043 2315 -10945
rect 2413 -11043 2414 -10945
rect 226 -11044 2414 -11043
rect 226 -11400 326 -11044
rect -1424 -11500 326 -11400
rect -15166 -11916 -1722 -11760
rect -15168 -26476 25000 -26400
rect -15168 -26630 -8072 -26476
rect 23928 -26630 25000 -26476
rect -15168 -26816 25000 -26630
rect -15168 -27116 -12216 -26816
rect -11616 -27116 24216 -26816
rect 24816 -27116 25000 -26816
rect -15168 -27200 25000 -27116
<< via4 >>
rect -15016 2240 -14320 2930
rect -974 2242 -284 2940
rect -13986 1650 -1428 1910
rect -13986 -10378 -13698 1650
rect -13698 1446 -1792 1650
rect -13698 -10378 -13498 1446
rect -1884 -9290 -1792 1446
rect -1792 -9290 -1428 1650
rect -1884 -9436 -1428 -9290
rect -13986 -10752 -2866 -10378
rect -2866 -10752 -2834 -10378
rect -15014 -11760 -14680 -11078
<< mimcap2 >>
rect -13982 2536 -8182 2986
rect -13982 2236 -13932 2536
rect -8232 2236 -8182 2536
rect -13982 2186 -8182 2236
rect -7582 2536 -1782 2986
rect -7582 2236 -7532 2536
rect -1832 2236 -1782 2536
rect -7582 2186 -1782 2236
rect -15068 -3946 -14668 1904
rect -15068 -4246 -15018 -3946
rect -14718 -4246 -14668 -3946
rect -13128 -3864 -8328 986
rect -13128 -4164 -13078 -3864
rect -8378 -4164 -8328 -3864
rect -13128 -4214 -8328 -4164
rect -7528 -3864 -2728 986
rect -7528 -4164 -7478 -3864
rect -2778 -4164 -2728 -3864
rect -7528 -4214 -2728 -4164
rect -1024 -3946 -624 1904
rect -15068 -4296 -14668 -4246
rect -1024 -4246 -974 -3946
rect -674 -4246 -624 -3946
rect -1024 -4296 -624 -4246
rect -15068 -10438 -14668 -4588
rect -13128 -9464 -8328 -4614
rect -13128 -9764 -13078 -9464
rect -8378 -9764 -8328 -9464
rect -13128 -9814 -8328 -9764
rect -7528 -9464 -2728 -4614
rect -7528 -9764 -7478 -9464
rect -2778 -9764 -2728 -9464
rect -7528 -9814 -2728 -9764
rect -15068 -10738 -15018 -10438
rect -14718 -10738 -14668 -10438
rect -15068 -10788 -14668 -10738
rect -1024 -10438 -624 -4588
rect -1024 -10724 -974 -10438
rect -674 -10724 -624 -10438
rect -1024 -10788 -624 -10724
rect -14482 -11464 -8682 -11014
rect -14482 -11764 -14432 -11464
rect -8732 -11764 -8682 -11464
rect -14482 -11814 -8682 -11764
rect -8082 -11464 -2282 -11014
rect -8082 -11764 -8032 -11464
rect -2332 -11764 -2282 -11464
rect -8082 -11814 -2282 -11764
<< mimcap2contact >>
rect -13932 2236 -8232 2536
rect -7532 2236 -1832 2536
rect -15018 -4246 -14718 -3946
rect -13078 -4164 -8378 -3864
rect -7478 -4164 -2778 -3864
rect -974 -4246 -674 -3946
rect -13078 -9764 -8378 -9464
rect -7478 -9764 -2778 -9464
rect -15018 -10738 -14718 -10438
rect -974 -10724 -674 -10438
rect -14432 -11764 -8732 -11464
rect -8032 -11764 -2332 -11464
<< metal5 >>
rect -15168 2940 -128 3086
rect -15168 2930 -974 2940
rect -15168 2240 -15016 2930
rect -14320 2536 -974 2930
rect -14320 2240 -13932 2536
rect -15168 2236 -13932 2240
rect -8232 2236 -7532 2536
rect -1832 2242 -974 2536
rect -284 2242 -128 2940
rect -1832 2236 -128 2242
rect -15168 1910 -128 2236
rect -15168 -3946 -13986 1910
rect -15168 -4246 -15018 -3946
rect -14718 -4246 -13986 -3946
rect -15168 -10438 -13986 -4246
rect -13498 -3864 -1884 1446
rect -13498 -4164 -13078 -3864
rect -8378 -4164 -7478 -3864
rect -2778 -4164 -1884 -3864
rect -13498 -9436 -1884 -4164
rect -1428 -3946 -128 1910
rect -1428 -4246 -974 -3946
rect -674 -4246 -128 -3946
rect -1428 -9436 -128 -4246
rect -13498 -9464 -128 -9436
rect -13498 -9764 -13078 -9464
rect -8378 -9764 -7478 -9464
rect -2778 -9518 -128 -9464
rect -2778 -9764 -2726 -9518
rect -13498 -10378 -2726 -9764
rect -15168 -10738 -15018 -10438
rect -14718 -10738 -13986 -10438
rect -15168 -10752 -13986 -10738
rect -2834 -10752 -2726 -10378
rect -15168 -10982 -2726 -10752
rect -1072 -10438 -128 -9518
rect -1072 -10724 -974 -10438
rect -674 -10724 -128 -10438
rect -1072 -10764 -128 -10724
rect -15168 -11078 -1828 -10982
rect -15168 -11760 -15014 -11078
rect -14680 -11464 -1828 -11078
rect -14680 -11760 -14432 -11464
rect -15168 -11764 -14432 -11760
rect -8732 -11764 -8032 -11464
rect -2332 -11764 -1828 -11464
rect -15168 -11916 -1828 -11764
<< labels >>
flabel metal1 -8078 -12352 -8078 -12352 1 FreeSans 480 0 0 0 vbias1
flabel metal1 -6206 -19026 -6206 -19026 1 FreeSans 480 0 0 0 vbias2
flabel metal1 23180 -19318 23204 -19288 1 FreeSans 480 0 0 0 VSS
port 6 n ground bidirectional
flabel metal1 23556 -18470 23556 -18470 1 FreeSans 480 0 0 0 vbias3
flabel metal1 23300 -18264 23300 -18264 1 FreeSans 480 0 0 0 vcascnm
flabel metal1 23436 -22496 23436 -22496 1 FreeSans 480 0 0 0 vbias4
flabel metal1 2138 -18102 2166 -18072 1 FreeSans 480 0 0 0 vtail_cascn
flabel metal1 2456 -14760 2488 -14720 1 FreeSans 480 0 0 0 vcascnp
flabel metal1 3322 -11898 3412 -11868 1 FreeSans 480 0 0 0 M8d
flabel metal1 2244 -18362 2282 -18326 1 FreeSans 480 0 0 0 vmirror
flabel metal1 22938 -16630 22974 -16600 1 FreeSans 480 0 0 0 M16d
flabel metal1 -10646 -21540 -10618 -21496 1 FreeSans 480 0 0 0 vip
port 1 n
flabel metal1 954 -21536 986 -21498 1 FreeSans 480 0 0 0 vim
port 2 n
flabel metal1 -5202 -24966 -5106 -24930 1 FreeSans 480 0 0 0 ibiasn
port 4 n
flabel metal1 -52 -22240 -4 -22216 1 FreeSans 480 0 0 0 vtail_cascn
flabel metal4 -10920 -26744 -10894 -26722 1 FreeSans 3200 0 0 0 VSS
flabel metal2 -6564 -19934 -6516 -19918 1 FreeSans 480 0 0 0 vcascpp
flabel metal1 -9488 -22168 -9456 -22140 1 FreeSans 480 0 0 0 vcascpm
flabel metal4 -11704 3910 -11678 4004 1 FreeSans 3200 0 0 0 VDD
port 5 n power bidirectional
flabel metal4 594 -11002 614 -10982 1 FreeSans 480 0 0 0 vo
port 3 n
flabel metal1 22608 -8372 22614 -8354 1 FreeSans 480 0 0 0 vo
flabel metal1 7498 -1550 7530 -1518 1 FreeSans 480 0 0 0 M9d
flabel metal1 2932 -5008 3004 -4978 1 FreeSans 480 0 0 0 vcascnm
flabel metal1 5656 -5000 5698 -4978 1 FreeSans 480 0 0 0 vcascnp
flabel metal1 4210 -5038 4236 -5000 1 FreeSans 480 0 0 0 vtail_cascp
flabel metal1 3698 -9046 3728 -9020 1 FreeSans 480 0 0 0 vip
flabel metal1 4706 -9050 4736 -9016 1 FreeSans 480 0 0 0 vim
flabel metal2 20172 -4390 20234 -4362 1 FreeSans 480 0 0 0 vmirror
flabel metal1 16210 -2186 16262 -2160 1 FreeSans 480 0 0 0 VDD
flabel metal2 10446 -3228 10514 -3198 1 FreeSans 480 0 0 0 vcascpp
flabel metal2 10670 -4260 10722 -4226 1 FreeSans 480 0 0 0 vcascpm
flabel metal2 8324 1884 8324 1884 1 FreeSans 480 0 0 0 vbias1
flabel metal2 9302 1622 9332 1650 1 FreeSans 480 0 0 0 VDD
flabel metal1 6346 610 6380 632 1 FreeSans 480 0 0 0 M7d
flabel metal2 7734 486 7792 522 1 FreeSans 480 0 0 0 M13d
flabel metal2 9760 -1694 9838 -1660 1 FreeSans 480 0 0 0 vtail_cascp
flabel metal1 17510 -5860 17546 -5832 1 FreeSans 480 0 0 0 VDD
flabel metal2 11866 -9908 11920 -9874 1 FreeSans 480 0 0 0 M8d
flabel metal2 12290 -4920 12372 -4888 1 FreeSans 480 0 0 0 vbias2
flabel metal2 16840 -7430 16902 -7400 1 FreeSans 480 0 0 0 M16d
flabel metal2 16432 -7118 16496 -7086 1 FreeSans 480 0 0 0 M13d
flabel metal1 7324 -5080 7364 -5046 1 FreeSans 480 0 0 0 M7d
flabel metal2 22394 -7218 22456 -7186 1 FreeSans 480 0 0 0 vmirror
flabel metal2 20508 -7328 20558 -7292 1 FreeSans 480 0 0 0 vcascpm
flabel metal2 20560 -8376 20652 -8344 1 FreeSans 480 0 0 0 vcascpp
flabel metal2 7618 -6048 7618 -6048 1 FreeSans 480 0 0 0 vbias1
flabel metal2 7488 -9634 7544 -9600 1 FreeSans 480 0 0 0 M9d
<< end >>
