magic
tech sky130A
magscale 1 2
timestamp 1624494425
<< error_p >>
rect 5 65 71 66
rect 0 1 6 65
rect 5 0 71 1
<< metal3 >>
rect 0 1 6 65
rect 70 1 76 65
<< via3 >>
rect 6 1 70 65
<< metal4 >>
rect 5 65 71 66
rect 5 1 6 65
rect 70 1 71 65
rect 5 0 71 1
<< properties >>
string FIXED_BBOX 0 0 76 66
<< end >>
