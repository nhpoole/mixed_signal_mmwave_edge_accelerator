magic
tech sky130A
timestamp 1626065694
<< checkpaint >>
rect -798 -1038 798 1038
<< metal4 >>
rect -168 379 168 408
rect -168 -379 -139 379
rect 139 -379 168 379
rect -168 -408 168 -379
<< via4 >>
rect -139 -379 139 379
<< metal5 >>
rect -168 379 168 408
rect -168 -379 -139 379
rect 139 -379 168 379
rect -168 -408 168 -379
<< end >>
