magic
tech sky130A
timestamp 1625948044
<< metal2 >>
rect -61 14 61 24
rect -61 -14 -54 14
rect -26 -14 -14 14
rect 14 -14 26 14
rect 54 -14 61 14
rect -61 -24 61 -14
<< via2 >>
rect -54 -14 -26 14
rect -14 -14 14 14
rect 26 -14 54 14
<< metal3 >>
rect -61 14 61 24
rect -61 -14 -54 14
rect -26 -14 -14 14
rect 14 -14 26 14
rect 54 -14 61 14
rect -61 -24 61 -14
<< end >>
