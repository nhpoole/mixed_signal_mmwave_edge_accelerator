magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect -1610 -1560 1609 1560
<< metal3 >>
rect -350 272 349 300
rect -350 208 265 272
rect 329 208 349 272
rect -350 192 349 208
rect -350 128 265 192
rect 329 128 349 192
rect -350 112 349 128
rect -350 48 265 112
rect 329 48 349 112
rect -350 32 349 48
rect -350 -32 265 32
rect 329 -32 349 32
rect -350 -48 349 -32
rect -350 -112 265 -48
rect 329 -112 349 -48
rect -350 -128 349 -112
rect -350 -192 265 -128
rect 329 -192 349 -128
rect -350 -208 349 -192
rect -350 -272 265 -208
rect 329 -272 349 -208
rect -350 -300 349 -272
<< via3 >>
rect 265 208 329 272
rect 265 128 329 192
rect 265 48 329 112
rect 265 -32 329 32
rect 265 -112 329 -48
rect 265 -192 329 -128
rect 265 -272 329 -208
<< mimcap >>
rect -250 152 150 200
rect -250 -152 -202 152
rect 102 -152 150 152
rect -250 -200 150 -152
<< mimcapcontact >>
rect -202 -152 102 152
<< metal4 >>
rect 249 272 345 288
rect 249 208 265 272
rect 329 208 345 272
rect 249 192 345 208
rect -211 152 111 161
rect -211 -152 -202 152
rect 102 -152 111 152
rect -211 -161 111 -152
rect 249 128 265 192
rect 329 128 345 192
rect 249 112 345 128
rect 249 48 265 112
rect 329 48 345 112
rect 249 32 345 48
rect 249 -32 265 32
rect 329 -32 345 32
rect 249 -48 345 -32
rect 249 -112 265 -48
rect 329 -112 345 -48
rect 249 -128 345 -112
rect 249 -192 265 -128
rect 329 -192 345 -128
rect 249 -208 345 -192
rect 249 -272 265 -208
rect 329 -272 345 -208
rect 249 -288 345 -272
<< properties >>
string FIXED_BBOX -350 -300 250 300
<< end >>
