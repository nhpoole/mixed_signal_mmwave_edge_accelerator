magic
tech sky130A
timestamp 1626065694
<< checkpaint >>
rect -677 -654 677 654
<< metal2 >>
rect -47 14 47 24
rect -47 -14 -34 14
rect -6 -14 6 14
rect 34 -14 47 14
rect -47 -24 47 -14
<< via2 >>
rect -34 -14 -6 14
rect 6 -14 34 14
<< metal3 >>
rect -47 14 47 24
rect -47 -14 -34 14
rect -6 -14 6 14
rect 34 -14 47 14
rect -47 -24 47 -14
<< end >>
