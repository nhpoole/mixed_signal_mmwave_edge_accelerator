magic
tech sky130A
magscale 1 2
timestamp 1621821863
<< nwell >>
rect -3323 -900 3323 900
<< pmoshvt >>
rect -3229 -800 -29 800
rect 29 -800 3229 800
<< pdiff >>
rect -3287 788 -3229 800
rect -3287 -788 -3275 788
rect -3241 -788 -3229 788
rect -3287 -800 -3229 -788
rect -29 788 29 800
rect -29 -788 -17 788
rect 17 -788 29 788
rect -29 -800 29 -788
rect 3229 788 3287 800
rect 3229 -788 3241 788
rect 3275 -788 3287 788
rect 3229 -800 3287 -788
<< pdiffc >>
rect -3275 -788 -3241 788
rect -17 -788 17 788
rect 3241 -788 3275 788
<< poly >>
rect -2595 881 -663 897
rect -2595 864 -2579 881
rect -3229 847 -2579 864
rect -679 864 -663 881
rect 663 881 2595 897
rect 663 864 679 881
rect -679 847 -29 864
rect -3229 800 -29 847
rect 29 847 679 864
rect 2579 864 2595 881
rect 2579 847 3229 864
rect 29 800 3229 847
rect -3229 -847 -29 -800
rect -3229 -864 -2579 -847
rect -2595 -881 -2579 -864
rect -679 -864 -29 -847
rect 29 -847 3229 -800
rect 29 -864 679 -847
rect -679 -881 -663 -864
rect -2595 -897 -663 -881
rect 663 -881 679 -864
rect 2579 -864 3229 -847
rect 2579 -881 2595 -864
rect 663 -897 2595 -881
<< polycont >>
rect -2579 847 -679 881
rect 679 847 2579 881
rect -2579 -881 -679 -847
rect 679 -881 2579 -847
<< locali >>
rect -2595 847 -2579 881
rect -679 847 -663 881
rect 663 847 679 881
rect 2579 847 2595 881
rect -3275 788 -3241 804
rect -3275 -804 -3241 -788
rect -17 788 17 804
rect -17 -804 17 -788
rect 3241 788 3275 804
rect 3241 -804 3275 -788
rect -2595 -881 -2579 -847
rect -679 -881 -663 -847
rect 663 -881 679 -847
rect 2579 -881 2595 -847
<< viali >>
rect -2421 847 -837 881
rect 837 847 2421 881
rect -3275 -788 -3241 788
rect -17 -788 17 788
rect 3241 -788 3275 788
rect -2421 -881 -837 -847
rect 837 -881 2421 -847
<< metal1 >>
rect -2433 881 -825 887
rect -2433 847 -2421 881
rect -837 847 -825 881
rect -2433 841 -825 847
rect 825 881 2433 887
rect 825 847 837 881
rect 2421 847 2433 881
rect 825 841 2433 847
rect -3281 788 -3235 800
rect -3281 -788 -3275 788
rect -3241 -788 -3235 788
rect -3281 -800 -3235 -788
rect -23 788 23 800
rect -23 -788 -17 788
rect 17 -788 23 788
rect -23 -800 23 -788
rect 3235 788 3281 800
rect 3235 -788 3241 788
rect 3275 -788 3281 788
rect 3235 -800 3281 -788
rect -2433 -847 -825 -841
rect -2433 -881 -2421 -847
rect -837 -881 -825 -847
rect -2433 -887 -825 -881
rect 825 -847 2433 -841
rect 825 -881 837 -847
rect 2421 -881 2433 -847
rect 825 -887 2433 -881
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_hvt
string parameters w 8 l 16 m 1 nf 2 diffcov 100 polycov 60 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
