magic
tech sky130A
timestamp 1626486988
<< checkpaint >>
rect -630 -630 726 726
<< metal1 >>
rect 0 3 3 93
rect 93 3 96 93
<< via1 >>
rect 3 3 93 93
<< metal2 >>
rect 3 93 93 96
rect 3 0 93 3
<< properties >>
string FIXED_BBOX 0 0 96 96
<< end >>
