magic
tech sky130A
magscale 1 2
timestamp 1624494425
<< nwell >>
rect -36 679 4832 1471
<< poly >>
rect 114 740 144 907
rect 81 674 144 740
rect 114 507 144 674
<< locali >>
rect 0 1397 4796 1431
rect 62 1130 96 1397
rect 274 1130 308 1397
rect 490 1130 524 1397
rect 706 1130 740 1397
rect 922 1130 956 1397
rect 1138 1130 1172 1397
rect 1354 1130 1388 1397
rect 1570 1130 1604 1397
rect 1786 1130 1820 1397
rect 2002 1130 2036 1397
rect 2218 1130 2252 1397
rect 2434 1130 2468 1397
rect 2650 1130 2684 1397
rect 2866 1130 2900 1397
rect 3082 1130 3116 1397
rect 3298 1130 3332 1397
rect 3514 1130 3548 1397
rect 3730 1130 3764 1397
rect 3946 1130 3980 1397
rect 4162 1130 4196 1397
rect 4378 1130 4412 1397
rect 4590 1130 4624 1397
rect 4694 1322 4728 1397
rect 64 674 98 740
rect 2326 724 2360 1096
rect 2326 690 2377 724
rect 2326 318 2360 690
rect 62 17 96 218
rect 274 17 308 218
rect 490 17 524 218
rect 706 17 740 218
rect 922 17 956 218
rect 1138 17 1172 218
rect 1354 17 1388 218
rect 1570 17 1604 218
rect 1786 17 1820 218
rect 2002 17 2036 218
rect 2218 17 2252 218
rect 2434 17 2468 218
rect 2650 17 2684 218
rect 2866 17 2900 218
rect 3082 17 3116 218
rect 3298 17 3332 218
rect 3514 17 3548 218
rect 3730 17 3764 218
rect 3946 17 3980 218
rect 4162 17 4196 218
rect 4378 17 4412 218
rect 4590 17 4624 218
rect 4694 17 4728 92
rect 0 -17 4796 17
use nmos_m42_w2_000_sli_dli_da_p  nmos_m42_w2_000_sli_dli_da_p_0
timestamp 1624494425
transform 1 0 54 0 1 51
box -26 -26 4604 456
use pmos_m42_w2_000_sli_dli_da_p  pmos_m42_w2_000_sli_dli_da_p_0
timestamp 1624494425
transform 1 0 54 0 1 963
box -59 -56 4637 454
use contact_15  contact_15_0
timestamp 1624494425
transform 1 0 48 0 1 674
box 0 0 66 66
use contact_28  contact_28_0
timestamp 1624494425
transform 1 0 4686 0 1 51
box -26 -26 76 108
use contact_27  contact_27_0
timestamp 1624494425
transform 1 0 4686 0 1 1281
box -59 -43 109 125
<< labels >>
rlabel locali s 81 707 81 707 4 A
rlabel locali s 2360 707 2360 707 4 Z
rlabel locali s 2398 0 2398 0 4 gnd
rlabel locali s 2398 1414 2398 1414 4 vdd
<< properties >>
string FIXED_BBOX 0 0 4796 1414
<< end >>
