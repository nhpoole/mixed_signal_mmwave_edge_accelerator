* Stimulus file.

.param vdd=1.8 Itail=10u vcmdes=1.1 vincm=1.1 vsig=0 Wp=1 Wn_diff=8 Wpcm=1 Wncm=8 Wn_bias=1 Lp=1 Ln_diff=1
+   Lpcm=1 Lncm=1 Ln_bias=4

vdd VDD GND 'vdd'
vip vip GND dc 'vincm+vsig' ac 1 0
vim vim GND dc 'vincm-vsig'
vocm vocm GND 'vcmdes'

*.options savecurrents
.save all
+ @m.xm1.msky130_fd_pr__nfet_01v8_lvt[id]
+ @m.xm1.msky130_fd_pr__nfet_01v8_lvt[vth]
+ @m.xm2.msky130_fd_pr__nfet_01v8_lvt[id]
+ @m.xm2.msky130_fd_pr__nfet_01v8_lvt[vth]
+ @m.xm3.msky130_fd_pr__nfet_01v8[id]
+ @m.xm3.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm4.msky130_fd_pr__pfet_01v8[id]
+ @m.xm4.msky130_fd_pr__pfet_01v8[vth]
+ @m.xm5.msky130_fd_pr__pfet_01v8[id]
+ @m.xm5.msky130_fd_pr__pfet_01v8[vth]
+ @m.xm6.msky130_fd_pr__pfet_01v8[id]
+ @m.xm6.msky130_fd_pr__pfet_01v8[vth]
+ @m.xm7.msky130_fd_pr__nfet_01v8[id]
+ @m.xm7.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm8.msky130_fd_pr__pfet_01v8[id]
+ @m.xm8.msky130_fd_pr__pfet_01v8[vth]
+ @m.xm9.msky130_fd_pr__pfet_01v8[id]
+ @m.xm9.msky130_fd_pr__pfet_01v8[vth]
+ @m.xm10.msky130_fd_pr__nfet_01v8[id]
+ @m.xm10.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm11.msky130_fd_pr__pfet_01v8[id]
+ @m.xm11.msky130_fd_pr__pfet_01v8[vth]
+ @m.xm12.msky130_fd_pr__nfet_01v8[id]
+ @m.xm12.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm13.msky130_fd_pr__nfet_01v8[id]
+ @m.xm13.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm14.msky130_fd_pr__nfet_01v8[id]
+ @m.xm14.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm15.msky130_fd_pr__nfet_01v8[id]
+ @m.xm15.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm16.msky130_fd_pr__nfet_01v8[id]
+ @m.xm16.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm16.msky130_fd_pr__nfet_01v8[cgg]
+ @m.xm17.msky130_fd_pr__nfet_01v8[id]
+ @m.xm17.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm18.msky130_fd_pr__nfet_01v8[id]
+ @m.xm18.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm18.msky130_fd_pr__nfet_01v8[cgg]
+ @m.xm19.msky130_fd_pr__nfet_01v8[id]
+ @m.xm19.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm56.msky130_fd_pr__pfet_01v8[id]
+ @m.xm56.msky130_fd_pr__pfet_01v8[vth]

*.op
*.print all
*write gm_c_stage_op.raw

* Control Block 1
*.control
*    op
*    print all
*    *ac dec 100 0.1 1g
*    noise v(vop, vom) vip dec 100 1 100k
*    run
*    *write gm_c_stage_ac.raw
*    *setplot noise1
*    *write gm_c_stage_noise1.raw v(onoise_spectrum) v(inoise_spectrum)
*    setplot noise2
*    write gm_c_stage_noise2.raw v(onoise_total) v(inoise_total)
*    quit
*.endc

* Control Block 2
.ac dec 100 0.1 1g
*.noise v(vop, vom) vip dec 100 1 100k
.control
    let incm = 0.4
    while incm < 1.6
        set incm = $&incm
        alter @vip[dc]=$incm
        alter @vim[dc]=$incm
        run
        write gm_c_stage_ac_{$incm}.raw
        *setplot noise1
        *write gm_c_stage_noise1_{$incm}.raw v(onoise_spectrum) v(inoise_spectrum)
        *setplot noise2
        *write gm_c_stage_noise2_{$incm}.raw v(onoise_total) v(inoise_total)
        let incm = incm + 0.1
    end
    alter @vip[dc]=0.7
    alter @vim[dc]=0.7
    op
    print all
    quit
.endc

* Control Block 3
*.ac dec 100 0.1 1g
*.control
*    let temperature = -40
*    while temperature < 130
*        set temp = $&temperature
*        run
*        write gm_c_stage_ac_temp_{$temp}.raw
*        let temperature = temperature + 10
*    end
*    quit
*.endc

* Control Block 4
*.ac dec 100 0.1 1g
*.control
*    let supply = 1.62
*    while supply < 2
*        alterparam vdd = {$&supply}
*        reset
*        run
*        write gm_c_stage_ac_vdd_{$&supply}.raw
*        let supply = supply + 0.04
*    end
*    quit
*.endc

