magic
tech sky130A
magscale 1 2
timestamp 1626065694
<< checkpaint >>
rect -13660 -28508 26260 3060
<< nwell >>
rect 342 -8918 24858 1758
<< pwell >>
rect -12348 -11304 24948 -11152
rect -12348 -27096 -12196 -11304
rect 2544 -12344 23014 -11692
rect -9222 -18864 50 -12486
rect 2544 -13578 23014 -12926
rect 2544 -14810 23014 -14158
rect 2542 -16044 23012 -15392
rect 2542 -17278 23012 -16626
rect 2542 -18510 23012 -17858
rect -2362 -19848 -72 -19596
rect 2542 -19744 23012 -19092
rect -2362 -20680 -72 -20428
rect 2542 -20978 23012 -20326
rect -9443 -22407 -3225 -21755
rect -2448 -22406 940 -21754
rect 2542 -22210 23012 -21558
rect -9444 -23520 -3226 -22868
rect -2448 -23518 940 -22866
rect 2542 -23444 23012 -22792
rect -9443 -24631 -3225 -23979
rect -2450 -24630 938 -23978
rect 2542 -24678 23012 -24026
rect -9444 -25744 -3226 -25092
rect -2450 -25740 938 -25088
rect 2542 -25910 23012 -25258
rect 24796 -27096 24948 -11304
rect -12348 -27248 24948 -27096
<< nmos >>
rect 2628 -12318 3588 -11718
rect 3646 -12318 4606 -11718
rect 4664 -12318 5624 -11718
rect 5682 -12318 6642 -11718
rect 6700 -12318 7660 -11718
rect 7718 -12318 8678 -11718
rect 8736 -12318 9696 -11718
rect 9754 -12318 10714 -11718
rect 10772 -12318 11732 -11718
rect 11790 -12318 12750 -11718
rect 12808 -12318 13768 -11718
rect 13826 -12318 14786 -11718
rect 14844 -12318 15804 -11718
rect 15862 -12318 16822 -11718
rect 16880 -12318 17840 -11718
rect 17898 -12318 18858 -11718
rect 18916 -12318 19876 -11718
rect 19934 -12318 20894 -11718
rect 20952 -12318 21912 -11718
rect 21970 -12318 22930 -11718
rect 2628 -13552 3588 -12952
rect 3646 -13552 4606 -12952
rect 4664 -13552 5624 -12952
rect 5682 -13552 6642 -12952
rect 6700 -13552 7660 -12952
rect 7718 -13552 8678 -12952
rect 8736 -13552 9696 -12952
rect 9754 -13552 10714 -12952
rect 10772 -13552 11732 -12952
rect 11790 -13552 12750 -12952
rect 12808 -13552 13768 -12952
rect 13826 -13552 14786 -12952
rect 14844 -13552 15804 -12952
rect 15862 -13552 16822 -12952
rect 16880 -13552 17840 -12952
rect 17898 -13552 18858 -12952
rect 18916 -13552 19876 -12952
rect 19934 -13552 20894 -12952
rect 20952 -13552 21912 -12952
rect 21970 -13552 22930 -12952
rect 2628 -14784 3588 -14184
rect 3646 -14784 4606 -14184
rect 4664 -14784 5624 -14184
rect 5682 -14784 6642 -14184
rect 6700 -14784 7660 -14184
rect 7718 -14784 8678 -14184
rect 8736 -14784 9696 -14184
rect 9754 -14784 10714 -14184
rect 10772 -14784 11732 -14184
rect 11790 -14784 12750 -14184
rect 12808 -14784 13768 -14184
rect 13826 -14784 14786 -14184
rect 14844 -14784 15804 -14184
rect 15862 -14784 16822 -14184
rect 16880 -14784 17840 -14184
rect 17898 -14784 18858 -14184
rect 18916 -14784 19876 -14184
rect 19934 -14784 20894 -14184
rect 20952 -14784 21912 -14184
rect 21970 -14784 22930 -14184
rect 2626 -16018 3586 -15418
rect 3644 -16018 4604 -15418
rect 4662 -16018 5622 -15418
rect 5680 -16018 6640 -15418
rect 6698 -16018 7658 -15418
rect 7716 -16018 8676 -15418
rect 8734 -16018 9694 -15418
rect 9752 -16018 10712 -15418
rect 10770 -16018 11730 -15418
rect 11788 -16018 12748 -15418
rect 12806 -16018 13766 -15418
rect 13824 -16018 14784 -15418
rect 14842 -16018 15802 -15418
rect 15860 -16018 16820 -15418
rect 16878 -16018 17838 -15418
rect 17896 -16018 18856 -15418
rect 18914 -16018 19874 -15418
rect 19932 -16018 20892 -15418
rect 20950 -16018 21910 -15418
rect 21968 -16018 22928 -15418
rect 2626 -17252 3586 -16652
rect 3644 -17252 4604 -16652
rect 4662 -17252 5622 -16652
rect 5680 -17252 6640 -16652
rect 6698 -17252 7658 -16652
rect 7716 -17252 8676 -16652
rect 8734 -17252 9694 -16652
rect 9752 -17252 10712 -16652
rect 10770 -17252 11730 -16652
rect 11788 -17252 12748 -16652
rect 12806 -17252 13766 -16652
rect 13824 -17252 14784 -16652
rect 14842 -17252 15802 -16652
rect 15860 -17252 16820 -16652
rect 16878 -17252 17838 -16652
rect 17896 -17252 18856 -16652
rect 18914 -17252 19874 -16652
rect 19932 -17252 20892 -16652
rect 20950 -17252 21910 -16652
rect 21968 -17252 22928 -16652
rect 2626 -18484 3586 -17884
rect 3644 -18484 4604 -17884
rect 4662 -18484 5622 -17884
rect 5680 -18484 6640 -17884
rect 6698 -18484 7658 -17884
rect 7716 -18484 8676 -17884
rect 8734 -18484 9694 -17884
rect 9752 -18484 10712 -17884
rect 10770 -18484 11730 -17884
rect 11788 -18484 12748 -17884
rect 12806 -18484 13766 -17884
rect 13824 -18484 14784 -17884
rect 14842 -18484 15802 -17884
rect 15860 -18484 16820 -17884
rect 16878 -18484 17838 -17884
rect 17896 -18484 18856 -17884
rect 18914 -18484 19874 -17884
rect 19932 -18484 20892 -17884
rect 20950 -18484 21910 -17884
rect 21968 -18484 22928 -17884
rect 2626 -19718 3586 -19118
rect 3644 -19718 4604 -19118
rect 4662 -19718 5622 -19118
rect 5680 -19718 6640 -19118
rect 6698 -19718 7658 -19118
rect 7716 -19718 8676 -19118
rect 8734 -19718 9694 -19118
rect 9752 -19718 10712 -19118
rect 10770 -19718 11730 -19118
rect 11788 -19718 12748 -19118
rect 12806 -19718 13766 -19118
rect 13824 -19718 14784 -19118
rect 14842 -19718 15802 -19118
rect 15860 -19718 16820 -19118
rect 16878 -19718 17838 -19118
rect 17896 -19718 18856 -19118
rect 18914 -19718 19874 -19118
rect 19932 -19718 20892 -19118
rect 20950 -19718 21910 -19118
rect 21968 -19718 22928 -19118
rect 2626 -20952 3586 -20352
rect 3644 -20952 4604 -20352
rect 4662 -20952 5622 -20352
rect 5680 -20952 6640 -20352
rect 6698 -20952 7658 -20352
rect 7716 -20952 8676 -20352
rect 8734 -20952 9694 -20352
rect 9752 -20952 10712 -20352
rect 10770 -20952 11730 -20352
rect 11788 -20952 12748 -20352
rect 12806 -20952 13766 -20352
rect 13824 -20952 14784 -20352
rect 14842 -20952 15802 -20352
rect 15860 -20952 16820 -20352
rect 16878 -20952 17838 -20352
rect 17896 -20952 18856 -20352
rect 18914 -20952 19874 -20352
rect 19932 -20952 20892 -20352
rect 20950 -20952 21910 -20352
rect 21968 -20952 22928 -20352
rect -9359 -22381 -8399 -21781
rect -8341 -22381 -7381 -21781
rect -7323 -22381 -6363 -21781
rect -6305 -22381 -5345 -21781
rect -5287 -22381 -4327 -21781
rect -4269 -22381 -3309 -21781
rect 2626 -22184 3586 -21584
rect 3644 -22184 4604 -21584
rect 4662 -22184 5622 -21584
rect 5680 -22184 6640 -21584
rect 6698 -22184 7658 -21584
rect 7716 -22184 8676 -21584
rect 8734 -22184 9694 -21584
rect 9752 -22184 10712 -21584
rect 10770 -22184 11730 -21584
rect 11788 -22184 12748 -21584
rect 12806 -22184 13766 -21584
rect 13824 -22184 14784 -21584
rect 14842 -22184 15802 -21584
rect 15860 -22184 16820 -21584
rect 16878 -22184 17838 -21584
rect 17896 -22184 18856 -21584
rect 18914 -22184 19874 -21584
rect 19932 -22184 20892 -21584
rect 20950 -22184 21910 -21584
rect 21968 -22184 22928 -21584
rect -9360 -23494 -8400 -22894
rect -8342 -23494 -7382 -22894
rect -7324 -23494 -6364 -22894
rect -6306 -23494 -5346 -22894
rect -5288 -23494 -4328 -22894
rect -4270 -23494 -3310 -22894
rect 2626 -23418 3586 -22818
rect 3644 -23418 4604 -22818
rect 4662 -23418 5622 -22818
rect 5680 -23418 6640 -22818
rect 6698 -23418 7658 -22818
rect 7716 -23418 8676 -22818
rect 8734 -23418 9694 -22818
rect 9752 -23418 10712 -22818
rect 10770 -23418 11730 -22818
rect 11788 -23418 12748 -22818
rect 12806 -23418 13766 -22818
rect 13824 -23418 14784 -22818
rect 14842 -23418 15802 -22818
rect 15860 -23418 16820 -22818
rect 16878 -23418 17838 -22818
rect 17896 -23418 18856 -22818
rect 18914 -23418 19874 -22818
rect 19932 -23418 20892 -22818
rect 20950 -23418 21910 -22818
rect 21968 -23418 22928 -22818
rect -9359 -24605 -8399 -24005
rect -8341 -24605 -7381 -24005
rect -7323 -24605 -6363 -24005
rect -6305 -24605 -5345 -24005
rect -5287 -24605 -4327 -24005
rect -4269 -24605 -3309 -24005
rect 2626 -24652 3586 -24052
rect 3644 -24652 4604 -24052
rect 4662 -24652 5622 -24052
rect 5680 -24652 6640 -24052
rect 6698 -24652 7658 -24052
rect 7716 -24652 8676 -24052
rect 8734 -24652 9694 -24052
rect 9752 -24652 10712 -24052
rect 10770 -24652 11730 -24052
rect 11788 -24652 12748 -24052
rect 12806 -24652 13766 -24052
rect 13824 -24652 14784 -24052
rect 14842 -24652 15802 -24052
rect 15860 -24652 16820 -24052
rect 16878 -24652 17838 -24052
rect 17896 -24652 18856 -24052
rect 18914 -24652 19874 -24052
rect 19932 -24652 20892 -24052
rect 20950 -24652 21910 -24052
rect 21968 -24652 22928 -24052
rect -9360 -25718 -8400 -25118
rect -8342 -25718 -7382 -25118
rect -7324 -25718 -6364 -25118
rect -6306 -25718 -5346 -25118
rect -5288 -25718 -4328 -25118
rect -4270 -25718 -3310 -25118
rect 2626 -25884 3586 -25284
rect 3644 -25884 4604 -25284
rect 4662 -25884 5622 -25284
rect 5680 -25884 6640 -25284
rect 6698 -25884 7658 -25284
rect 7716 -25884 8676 -25284
rect 8734 -25884 9694 -25284
rect 9752 -25884 10712 -25284
rect 10770 -25884 11730 -25284
rect 11788 -25884 12748 -25284
rect 12806 -25884 13766 -25284
rect 13824 -25884 14784 -25284
rect 14842 -25884 15802 -25284
rect 15860 -25884 16820 -25284
rect 16878 -25884 17838 -25284
rect 17896 -25884 18856 -25284
rect 18914 -25884 19874 -25284
rect 19932 -25884 20892 -25284
rect 20950 -25884 21910 -25284
rect 21968 -25884 22928 -25284
<< pmos >>
rect 3672 -5090 3832 -4690
rect 3890 -5090 4050 -4690
rect 4108 -5090 4268 -4690
rect 4326 -5090 4486 -4690
rect 4544 -5090 4704 -4690
rect 4762 -5090 4922 -4690
rect 4980 -5090 5140 -4690
rect 5198 -5090 5358 -4690
rect 5416 -5090 5576 -4690
rect 5634 -5090 5794 -4690
rect 3672 -6028 3832 -5628
rect 3890 -6028 4050 -5628
rect 4108 -6028 4268 -5628
rect 4326 -6028 4486 -5628
rect 4544 -6028 4704 -5628
rect 4762 -6028 4922 -5628
rect 4980 -6028 5140 -5628
rect 5198 -6028 5358 -5628
rect 5416 -6028 5576 -5628
rect 5634 -6028 5794 -5628
rect 3672 -6966 3832 -6566
rect 3890 -6966 4050 -6566
rect 4108 -6966 4268 -6566
rect 4326 -6966 4486 -6566
rect 4544 -6966 4704 -6566
rect 4762 -6966 4922 -6566
rect 4980 -6966 5140 -6566
rect 5198 -6966 5358 -6566
rect 5416 -6966 5576 -6566
rect 5634 -6966 5794 -6566
rect 3672 -7904 3832 -7504
rect 3890 -7904 4050 -7504
rect 4108 -7904 4268 -7504
rect 4326 -7904 4486 -7504
rect 4544 -7904 4704 -7504
rect 4762 -7904 4922 -7504
rect 4980 -7904 5140 -7504
rect 5198 -7904 5358 -7504
rect 5416 -7904 5576 -7504
rect 5634 -7904 5794 -7504
<< nmoslvt >>
rect -9138 -13112 -8178 -12512
rect -8120 -13112 -7160 -12512
rect -7102 -13112 -6142 -12512
rect -6084 -13112 -5124 -12512
rect -5066 -13112 -4106 -12512
rect -4048 -13112 -3088 -12512
rect -3030 -13112 -2070 -12512
rect -2012 -13112 -1052 -12512
rect -994 -13112 -34 -12512
rect -9138 -13930 -8178 -13330
rect -8120 -13930 -7160 -13330
rect -7102 -13930 -6142 -13330
rect -6084 -13930 -5124 -13330
rect -5066 -13930 -4106 -13330
rect -4048 -13930 -3088 -13330
rect -3030 -13930 -2070 -13330
rect -2012 -13930 -1052 -13330
rect -994 -13930 -34 -13330
rect -9138 -14748 -8178 -14148
rect -8120 -14748 -7160 -14148
rect -7102 -14748 -6142 -14148
rect -6084 -14748 -5124 -14148
rect -5066 -14748 -4106 -14148
rect -4048 -14748 -3088 -14148
rect -3030 -14748 -2070 -14148
rect -2012 -14748 -1052 -14148
rect -994 -14748 -34 -14148
rect -9138 -15566 -8178 -14966
rect -8120 -15566 -7160 -14966
rect -7102 -15566 -6142 -14966
rect -6084 -15566 -5124 -14966
rect -5066 -15566 -4106 -14966
rect -4048 -15566 -3088 -14966
rect -3030 -15566 -2070 -14966
rect -2012 -15566 -1052 -14966
rect -994 -15566 -34 -14966
rect -9138 -16384 -8178 -15784
rect -8120 -16384 -7160 -15784
rect -7102 -16384 -6142 -15784
rect -6084 -16384 -5124 -15784
rect -5066 -16384 -4106 -15784
rect -4048 -16384 -3088 -15784
rect -3030 -16384 -2070 -15784
rect -2012 -16384 -1052 -15784
rect -994 -16384 -34 -15784
rect -9138 -17202 -8178 -16602
rect -8120 -17202 -7160 -16602
rect -7102 -17202 -6142 -16602
rect -6084 -17202 -5124 -16602
rect -5066 -17202 -4106 -16602
rect -4048 -17202 -3088 -16602
rect -3030 -17202 -2070 -16602
rect -2012 -17202 -1052 -16602
rect -994 -17202 -34 -16602
rect -9138 -18020 -8178 -17420
rect -8120 -18020 -7160 -17420
rect -7102 -18020 -6142 -17420
rect -6084 -18020 -5124 -17420
rect -5066 -18020 -4106 -17420
rect -4048 -18020 -3088 -17420
rect -3030 -18020 -2070 -17420
rect -2012 -18020 -1052 -17420
rect -994 -18020 -34 -17420
rect -9138 -18838 -8178 -18238
rect -8120 -18838 -7160 -18238
rect -7102 -18838 -6142 -18238
rect -6084 -18838 -5124 -18238
rect -5066 -18838 -4106 -18238
rect -4048 -18838 -3088 -18238
rect -3030 -18838 -2070 -18238
rect -2012 -18838 -1052 -18238
rect -994 -18838 -34 -18238
rect -2278 -19822 -2118 -19622
rect -2060 -19822 -1900 -19622
rect -1842 -19822 -1682 -19622
rect -1624 -19822 -1464 -19622
rect -1406 -19822 -1246 -19622
rect -1188 -19822 -1028 -19622
rect -970 -19822 -810 -19622
rect -752 -19822 -592 -19622
rect -534 -19822 -374 -19622
rect -316 -19822 -156 -19622
rect -2278 -20654 -2118 -20454
rect -2060 -20654 -1900 -20454
rect -1842 -20654 -1682 -20454
rect -1624 -20654 -1464 -20454
rect -1406 -20654 -1246 -20454
rect -1188 -20654 -1028 -20454
rect -970 -20654 -810 -20454
rect -752 -20654 -592 -20454
rect -534 -20654 -374 -20454
rect -316 -20654 -156 -20454
rect -2364 -22380 -2124 -21780
rect -2066 -22380 -1826 -21780
rect -1768 -22380 -1528 -21780
rect -1470 -22380 -1230 -21780
rect -1172 -22380 -932 -21780
rect -874 -22380 -634 -21780
rect -576 -22380 -336 -21780
rect -278 -22380 -38 -21780
rect 20 -22380 260 -21780
rect 318 -22380 558 -21780
rect 616 -22380 856 -21780
rect -2364 -23492 -2124 -22892
rect -2066 -23492 -1826 -22892
rect -1768 -23492 -1528 -22892
rect -1470 -23492 -1230 -22892
rect -1172 -23492 -932 -22892
rect -874 -23492 -634 -22892
rect -576 -23492 -336 -22892
rect -278 -23492 -38 -22892
rect 20 -23492 260 -22892
rect 318 -23492 558 -22892
rect 616 -23492 856 -22892
rect -2366 -24604 -2126 -24004
rect -2068 -24604 -1828 -24004
rect -1770 -24604 -1530 -24004
rect -1472 -24604 -1232 -24004
rect -1174 -24604 -934 -24004
rect -876 -24604 -636 -24004
rect -578 -24604 -338 -24004
rect -280 -24604 -40 -24004
rect 18 -24604 258 -24004
rect 316 -24604 556 -24004
rect 614 -24604 854 -24004
rect -2366 -25714 -2126 -25114
rect -2068 -25714 -1828 -25114
rect -1770 -25714 -1530 -25114
rect -1472 -25714 -1232 -25114
rect -1174 -25714 -934 -25114
rect -876 -25714 -636 -25114
rect -578 -25714 -338 -25114
rect -280 -25714 -40 -25114
rect 18 -25714 258 -25114
rect 316 -25714 556 -25114
rect 614 -25714 854 -25114
<< ndiff >>
rect 2570 -11763 2628 -11718
rect 2570 -11797 2582 -11763
rect 2616 -11797 2628 -11763
rect 2570 -11831 2628 -11797
rect 2570 -11865 2582 -11831
rect 2616 -11865 2628 -11831
rect 2570 -11899 2628 -11865
rect 2570 -11933 2582 -11899
rect 2616 -11933 2628 -11899
rect 2570 -11967 2628 -11933
rect 2570 -12001 2582 -11967
rect 2616 -12001 2628 -11967
rect 2570 -12035 2628 -12001
rect 2570 -12069 2582 -12035
rect 2616 -12069 2628 -12035
rect 2570 -12103 2628 -12069
rect 2570 -12137 2582 -12103
rect 2616 -12137 2628 -12103
rect 2570 -12171 2628 -12137
rect 2570 -12205 2582 -12171
rect 2616 -12205 2628 -12171
rect 2570 -12239 2628 -12205
rect 2570 -12273 2582 -12239
rect 2616 -12273 2628 -12239
rect 2570 -12318 2628 -12273
rect 3588 -11763 3646 -11718
rect 3588 -11797 3600 -11763
rect 3634 -11797 3646 -11763
rect 3588 -11831 3646 -11797
rect 3588 -11865 3600 -11831
rect 3634 -11865 3646 -11831
rect 3588 -11899 3646 -11865
rect 3588 -11933 3600 -11899
rect 3634 -11933 3646 -11899
rect 3588 -11967 3646 -11933
rect 3588 -12001 3600 -11967
rect 3634 -12001 3646 -11967
rect 3588 -12035 3646 -12001
rect 3588 -12069 3600 -12035
rect 3634 -12069 3646 -12035
rect 3588 -12103 3646 -12069
rect 3588 -12137 3600 -12103
rect 3634 -12137 3646 -12103
rect 3588 -12171 3646 -12137
rect 3588 -12205 3600 -12171
rect 3634 -12205 3646 -12171
rect 3588 -12239 3646 -12205
rect 3588 -12273 3600 -12239
rect 3634 -12273 3646 -12239
rect 3588 -12318 3646 -12273
rect 4606 -11763 4664 -11718
rect 4606 -11797 4618 -11763
rect 4652 -11797 4664 -11763
rect 4606 -11831 4664 -11797
rect 4606 -11865 4618 -11831
rect 4652 -11865 4664 -11831
rect 4606 -11899 4664 -11865
rect 4606 -11933 4618 -11899
rect 4652 -11933 4664 -11899
rect 4606 -11967 4664 -11933
rect 4606 -12001 4618 -11967
rect 4652 -12001 4664 -11967
rect 4606 -12035 4664 -12001
rect 4606 -12069 4618 -12035
rect 4652 -12069 4664 -12035
rect 4606 -12103 4664 -12069
rect 4606 -12137 4618 -12103
rect 4652 -12137 4664 -12103
rect 4606 -12171 4664 -12137
rect 4606 -12205 4618 -12171
rect 4652 -12205 4664 -12171
rect 4606 -12239 4664 -12205
rect 4606 -12273 4618 -12239
rect 4652 -12273 4664 -12239
rect 4606 -12318 4664 -12273
rect 5624 -11763 5682 -11718
rect 5624 -11797 5636 -11763
rect 5670 -11797 5682 -11763
rect 5624 -11831 5682 -11797
rect 5624 -11865 5636 -11831
rect 5670 -11865 5682 -11831
rect 5624 -11899 5682 -11865
rect 5624 -11933 5636 -11899
rect 5670 -11933 5682 -11899
rect 5624 -11967 5682 -11933
rect 5624 -12001 5636 -11967
rect 5670 -12001 5682 -11967
rect 5624 -12035 5682 -12001
rect 5624 -12069 5636 -12035
rect 5670 -12069 5682 -12035
rect 5624 -12103 5682 -12069
rect 5624 -12137 5636 -12103
rect 5670 -12137 5682 -12103
rect 5624 -12171 5682 -12137
rect 5624 -12205 5636 -12171
rect 5670 -12205 5682 -12171
rect 5624 -12239 5682 -12205
rect 5624 -12273 5636 -12239
rect 5670 -12273 5682 -12239
rect 5624 -12318 5682 -12273
rect 6642 -11763 6700 -11718
rect 6642 -11797 6654 -11763
rect 6688 -11797 6700 -11763
rect 6642 -11831 6700 -11797
rect 6642 -11865 6654 -11831
rect 6688 -11865 6700 -11831
rect 6642 -11899 6700 -11865
rect 6642 -11933 6654 -11899
rect 6688 -11933 6700 -11899
rect 6642 -11967 6700 -11933
rect 6642 -12001 6654 -11967
rect 6688 -12001 6700 -11967
rect 6642 -12035 6700 -12001
rect 6642 -12069 6654 -12035
rect 6688 -12069 6700 -12035
rect 6642 -12103 6700 -12069
rect 6642 -12137 6654 -12103
rect 6688 -12137 6700 -12103
rect 6642 -12171 6700 -12137
rect 6642 -12205 6654 -12171
rect 6688 -12205 6700 -12171
rect 6642 -12239 6700 -12205
rect 6642 -12273 6654 -12239
rect 6688 -12273 6700 -12239
rect 6642 -12318 6700 -12273
rect 7660 -11763 7718 -11718
rect 7660 -11797 7672 -11763
rect 7706 -11797 7718 -11763
rect 7660 -11831 7718 -11797
rect 7660 -11865 7672 -11831
rect 7706 -11865 7718 -11831
rect 7660 -11899 7718 -11865
rect 7660 -11933 7672 -11899
rect 7706 -11933 7718 -11899
rect 7660 -11967 7718 -11933
rect 7660 -12001 7672 -11967
rect 7706 -12001 7718 -11967
rect 7660 -12035 7718 -12001
rect 7660 -12069 7672 -12035
rect 7706 -12069 7718 -12035
rect 7660 -12103 7718 -12069
rect 7660 -12137 7672 -12103
rect 7706 -12137 7718 -12103
rect 7660 -12171 7718 -12137
rect 7660 -12205 7672 -12171
rect 7706 -12205 7718 -12171
rect 7660 -12239 7718 -12205
rect 7660 -12273 7672 -12239
rect 7706 -12273 7718 -12239
rect 7660 -12318 7718 -12273
rect 8678 -11763 8736 -11718
rect 8678 -11797 8690 -11763
rect 8724 -11797 8736 -11763
rect 8678 -11831 8736 -11797
rect 8678 -11865 8690 -11831
rect 8724 -11865 8736 -11831
rect 8678 -11899 8736 -11865
rect 8678 -11933 8690 -11899
rect 8724 -11933 8736 -11899
rect 8678 -11967 8736 -11933
rect 8678 -12001 8690 -11967
rect 8724 -12001 8736 -11967
rect 8678 -12035 8736 -12001
rect 8678 -12069 8690 -12035
rect 8724 -12069 8736 -12035
rect 8678 -12103 8736 -12069
rect 8678 -12137 8690 -12103
rect 8724 -12137 8736 -12103
rect 8678 -12171 8736 -12137
rect 8678 -12205 8690 -12171
rect 8724 -12205 8736 -12171
rect 8678 -12239 8736 -12205
rect 8678 -12273 8690 -12239
rect 8724 -12273 8736 -12239
rect 8678 -12318 8736 -12273
rect 9696 -11763 9754 -11718
rect 9696 -11797 9708 -11763
rect 9742 -11797 9754 -11763
rect 9696 -11831 9754 -11797
rect 9696 -11865 9708 -11831
rect 9742 -11865 9754 -11831
rect 9696 -11899 9754 -11865
rect 9696 -11933 9708 -11899
rect 9742 -11933 9754 -11899
rect 9696 -11967 9754 -11933
rect 9696 -12001 9708 -11967
rect 9742 -12001 9754 -11967
rect 9696 -12035 9754 -12001
rect 9696 -12069 9708 -12035
rect 9742 -12069 9754 -12035
rect 9696 -12103 9754 -12069
rect 9696 -12137 9708 -12103
rect 9742 -12137 9754 -12103
rect 9696 -12171 9754 -12137
rect 9696 -12205 9708 -12171
rect 9742 -12205 9754 -12171
rect 9696 -12239 9754 -12205
rect 9696 -12273 9708 -12239
rect 9742 -12273 9754 -12239
rect 9696 -12318 9754 -12273
rect 10714 -11763 10772 -11718
rect 10714 -11797 10726 -11763
rect 10760 -11797 10772 -11763
rect 10714 -11831 10772 -11797
rect 10714 -11865 10726 -11831
rect 10760 -11865 10772 -11831
rect 10714 -11899 10772 -11865
rect 10714 -11933 10726 -11899
rect 10760 -11933 10772 -11899
rect 10714 -11967 10772 -11933
rect 10714 -12001 10726 -11967
rect 10760 -12001 10772 -11967
rect 10714 -12035 10772 -12001
rect 10714 -12069 10726 -12035
rect 10760 -12069 10772 -12035
rect 10714 -12103 10772 -12069
rect 10714 -12137 10726 -12103
rect 10760 -12137 10772 -12103
rect 10714 -12171 10772 -12137
rect 10714 -12205 10726 -12171
rect 10760 -12205 10772 -12171
rect 10714 -12239 10772 -12205
rect 10714 -12273 10726 -12239
rect 10760 -12273 10772 -12239
rect 10714 -12318 10772 -12273
rect 11732 -11763 11790 -11718
rect 11732 -11797 11744 -11763
rect 11778 -11797 11790 -11763
rect 11732 -11831 11790 -11797
rect 11732 -11865 11744 -11831
rect 11778 -11865 11790 -11831
rect 11732 -11899 11790 -11865
rect 11732 -11933 11744 -11899
rect 11778 -11933 11790 -11899
rect 11732 -11967 11790 -11933
rect 11732 -12001 11744 -11967
rect 11778 -12001 11790 -11967
rect 11732 -12035 11790 -12001
rect 11732 -12069 11744 -12035
rect 11778 -12069 11790 -12035
rect 11732 -12103 11790 -12069
rect 11732 -12137 11744 -12103
rect 11778 -12137 11790 -12103
rect 11732 -12171 11790 -12137
rect 11732 -12205 11744 -12171
rect 11778 -12205 11790 -12171
rect 11732 -12239 11790 -12205
rect 11732 -12273 11744 -12239
rect 11778 -12273 11790 -12239
rect 11732 -12318 11790 -12273
rect 12750 -11763 12808 -11718
rect 12750 -11797 12762 -11763
rect 12796 -11797 12808 -11763
rect 12750 -11831 12808 -11797
rect 12750 -11865 12762 -11831
rect 12796 -11865 12808 -11831
rect 12750 -11899 12808 -11865
rect 12750 -11933 12762 -11899
rect 12796 -11933 12808 -11899
rect 12750 -11967 12808 -11933
rect 12750 -12001 12762 -11967
rect 12796 -12001 12808 -11967
rect 12750 -12035 12808 -12001
rect 12750 -12069 12762 -12035
rect 12796 -12069 12808 -12035
rect 12750 -12103 12808 -12069
rect 12750 -12137 12762 -12103
rect 12796 -12137 12808 -12103
rect 12750 -12171 12808 -12137
rect 12750 -12205 12762 -12171
rect 12796 -12205 12808 -12171
rect 12750 -12239 12808 -12205
rect 12750 -12273 12762 -12239
rect 12796 -12273 12808 -12239
rect 12750 -12318 12808 -12273
rect 13768 -11763 13826 -11718
rect 13768 -11797 13780 -11763
rect 13814 -11797 13826 -11763
rect 13768 -11831 13826 -11797
rect 13768 -11865 13780 -11831
rect 13814 -11865 13826 -11831
rect 13768 -11899 13826 -11865
rect 13768 -11933 13780 -11899
rect 13814 -11933 13826 -11899
rect 13768 -11967 13826 -11933
rect 13768 -12001 13780 -11967
rect 13814 -12001 13826 -11967
rect 13768 -12035 13826 -12001
rect 13768 -12069 13780 -12035
rect 13814 -12069 13826 -12035
rect 13768 -12103 13826 -12069
rect 13768 -12137 13780 -12103
rect 13814 -12137 13826 -12103
rect 13768 -12171 13826 -12137
rect 13768 -12205 13780 -12171
rect 13814 -12205 13826 -12171
rect 13768 -12239 13826 -12205
rect 13768 -12273 13780 -12239
rect 13814 -12273 13826 -12239
rect 13768 -12318 13826 -12273
rect 14786 -11763 14844 -11718
rect 14786 -11797 14798 -11763
rect 14832 -11797 14844 -11763
rect 14786 -11831 14844 -11797
rect 14786 -11865 14798 -11831
rect 14832 -11865 14844 -11831
rect 14786 -11899 14844 -11865
rect 14786 -11933 14798 -11899
rect 14832 -11933 14844 -11899
rect 14786 -11967 14844 -11933
rect 14786 -12001 14798 -11967
rect 14832 -12001 14844 -11967
rect 14786 -12035 14844 -12001
rect 14786 -12069 14798 -12035
rect 14832 -12069 14844 -12035
rect 14786 -12103 14844 -12069
rect 14786 -12137 14798 -12103
rect 14832 -12137 14844 -12103
rect 14786 -12171 14844 -12137
rect 14786 -12205 14798 -12171
rect 14832 -12205 14844 -12171
rect 14786 -12239 14844 -12205
rect 14786 -12273 14798 -12239
rect 14832 -12273 14844 -12239
rect 14786 -12318 14844 -12273
rect 15804 -11763 15862 -11718
rect 15804 -11797 15816 -11763
rect 15850 -11797 15862 -11763
rect 15804 -11831 15862 -11797
rect 15804 -11865 15816 -11831
rect 15850 -11865 15862 -11831
rect 15804 -11899 15862 -11865
rect 15804 -11933 15816 -11899
rect 15850 -11933 15862 -11899
rect 15804 -11967 15862 -11933
rect 15804 -12001 15816 -11967
rect 15850 -12001 15862 -11967
rect 15804 -12035 15862 -12001
rect 15804 -12069 15816 -12035
rect 15850 -12069 15862 -12035
rect 15804 -12103 15862 -12069
rect 15804 -12137 15816 -12103
rect 15850 -12137 15862 -12103
rect 15804 -12171 15862 -12137
rect 15804 -12205 15816 -12171
rect 15850 -12205 15862 -12171
rect 15804 -12239 15862 -12205
rect 15804 -12273 15816 -12239
rect 15850 -12273 15862 -12239
rect 15804 -12318 15862 -12273
rect 16822 -11763 16880 -11718
rect 16822 -11797 16834 -11763
rect 16868 -11797 16880 -11763
rect 16822 -11831 16880 -11797
rect 16822 -11865 16834 -11831
rect 16868 -11865 16880 -11831
rect 16822 -11899 16880 -11865
rect 16822 -11933 16834 -11899
rect 16868 -11933 16880 -11899
rect 16822 -11967 16880 -11933
rect 16822 -12001 16834 -11967
rect 16868 -12001 16880 -11967
rect 16822 -12035 16880 -12001
rect 16822 -12069 16834 -12035
rect 16868 -12069 16880 -12035
rect 16822 -12103 16880 -12069
rect 16822 -12137 16834 -12103
rect 16868 -12137 16880 -12103
rect 16822 -12171 16880 -12137
rect 16822 -12205 16834 -12171
rect 16868 -12205 16880 -12171
rect 16822 -12239 16880 -12205
rect 16822 -12273 16834 -12239
rect 16868 -12273 16880 -12239
rect 16822 -12318 16880 -12273
rect 17840 -11763 17898 -11718
rect 17840 -11797 17852 -11763
rect 17886 -11797 17898 -11763
rect 17840 -11831 17898 -11797
rect 17840 -11865 17852 -11831
rect 17886 -11865 17898 -11831
rect 17840 -11899 17898 -11865
rect 17840 -11933 17852 -11899
rect 17886 -11933 17898 -11899
rect 17840 -11967 17898 -11933
rect 17840 -12001 17852 -11967
rect 17886 -12001 17898 -11967
rect 17840 -12035 17898 -12001
rect 17840 -12069 17852 -12035
rect 17886 -12069 17898 -12035
rect 17840 -12103 17898 -12069
rect 17840 -12137 17852 -12103
rect 17886 -12137 17898 -12103
rect 17840 -12171 17898 -12137
rect 17840 -12205 17852 -12171
rect 17886 -12205 17898 -12171
rect 17840 -12239 17898 -12205
rect 17840 -12273 17852 -12239
rect 17886 -12273 17898 -12239
rect 17840 -12318 17898 -12273
rect 18858 -11763 18916 -11718
rect 18858 -11797 18870 -11763
rect 18904 -11797 18916 -11763
rect 18858 -11831 18916 -11797
rect 18858 -11865 18870 -11831
rect 18904 -11865 18916 -11831
rect 18858 -11899 18916 -11865
rect 18858 -11933 18870 -11899
rect 18904 -11933 18916 -11899
rect 18858 -11967 18916 -11933
rect 18858 -12001 18870 -11967
rect 18904 -12001 18916 -11967
rect 18858 -12035 18916 -12001
rect 18858 -12069 18870 -12035
rect 18904 -12069 18916 -12035
rect 18858 -12103 18916 -12069
rect 18858 -12137 18870 -12103
rect 18904 -12137 18916 -12103
rect 18858 -12171 18916 -12137
rect 18858 -12205 18870 -12171
rect 18904 -12205 18916 -12171
rect 18858 -12239 18916 -12205
rect 18858 -12273 18870 -12239
rect 18904 -12273 18916 -12239
rect 18858 -12318 18916 -12273
rect 19876 -11763 19934 -11718
rect 19876 -11797 19888 -11763
rect 19922 -11797 19934 -11763
rect 19876 -11831 19934 -11797
rect 19876 -11865 19888 -11831
rect 19922 -11865 19934 -11831
rect 19876 -11899 19934 -11865
rect 19876 -11933 19888 -11899
rect 19922 -11933 19934 -11899
rect 19876 -11967 19934 -11933
rect 19876 -12001 19888 -11967
rect 19922 -12001 19934 -11967
rect 19876 -12035 19934 -12001
rect 19876 -12069 19888 -12035
rect 19922 -12069 19934 -12035
rect 19876 -12103 19934 -12069
rect 19876 -12137 19888 -12103
rect 19922 -12137 19934 -12103
rect 19876 -12171 19934 -12137
rect 19876 -12205 19888 -12171
rect 19922 -12205 19934 -12171
rect 19876 -12239 19934 -12205
rect 19876 -12273 19888 -12239
rect 19922 -12273 19934 -12239
rect 19876 -12318 19934 -12273
rect 20894 -11763 20952 -11718
rect 20894 -11797 20906 -11763
rect 20940 -11797 20952 -11763
rect 20894 -11831 20952 -11797
rect 20894 -11865 20906 -11831
rect 20940 -11865 20952 -11831
rect 20894 -11899 20952 -11865
rect 20894 -11933 20906 -11899
rect 20940 -11933 20952 -11899
rect 20894 -11967 20952 -11933
rect 20894 -12001 20906 -11967
rect 20940 -12001 20952 -11967
rect 20894 -12035 20952 -12001
rect 20894 -12069 20906 -12035
rect 20940 -12069 20952 -12035
rect 20894 -12103 20952 -12069
rect 20894 -12137 20906 -12103
rect 20940 -12137 20952 -12103
rect 20894 -12171 20952 -12137
rect 20894 -12205 20906 -12171
rect 20940 -12205 20952 -12171
rect 20894 -12239 20952 -12205
rect 20894 -12273 20906 -12239
rect 20940 -12273 20952 -12239
rect 20894 -12318 20952 -12273
rect 21912 -11763 21970 -11718
rect 21912 -11797 21924 -11763
rect 21958 -11797 21970 -11763
rect 21912 -11831 21970 -11797
rect 21912 -11865 21924 -11831
rect 21958 -11865 21970 -11831
rect 21912 -11899 21970 -11865
rect 21912 -11933 21924 -11899
rect 21958 -11933 21970 -11899
rect 21912 -11967 21970 -11933
rect 21912 -12001 21924 -11967
rect 21958 -12001 21970 -11967
rect 21912 -12035 21970 -12001
rect 21912 -12069 21924 -12035
rect 21958 -12069 21970 -12035
rect 21912 -12103 21970 -12069
rect 21912 -12137 21924 -12103
rect 21958 -12137 21970 -12103
rect 21912 -12171 21970 -12137
rect 21912 -12205 21924 -12171
rect 21958 -12205 21970 -12171
rect 21912 -12239 21970 -12205
rect 21912 -12273 21924 -12239
rect 21958 -12273 21970 -12239
rect 21912 -12318 21970 -12273
rect 22930 -11763 22988 -11718
rect 22930 -11797 22942 -11763
rect 22976 -11797 22988 -11763
rect 22930 -11831 22988 -11797
rect 22930 -11865 22942 -11831
rect 22976 -11865 22988 -11831
rect 22930 -11899 22988 -11865
rect 22930 -11933 22942 -11899
rect 22976 -11933 22988 -11899
rect 22930 -11967 22988 -11933
rect 22930 -12001 22942 -11967
rect 22976 -12001 22988 -11967
rect 22930 -12035 22988 -12001
rect 22930 -12069 22942 -12035
rect 22976 -12069 22988 -12035
rect 22930 -12103 22988 -12069
rect 22930 -12137 22942 -12103
rect 22976 -12137 22988 -12103
rect 22930 -12171 22988 -12137
rect 22930 -12205 22942 -12171
rect 22976 -12205 22988 -12171
rect 22930 -12239 22988 -12205
rect 22930 -12273 22942 -12239
rect 22976 -12273 22988 -12239
rect 22930 -12318 22988 -12273
rect -9196 -12557 -9138 -12512
rect -9196 -12591 -9184 -12557
rect -9150 -12591 -9138 -12557
rect -9196 -12625 -9138 -12591
rect -9196 -12659 -9184 -12625
rect -9150 -12659 -9138 -12625
rect -9196 -12693 -9138 -12659
rect -9196 -12727 -9184 -12693
rect -9150 -12727 -9138 -12693
rect -9196 -12761 -9138 -12727
rect -9196 -12795 -9184 -12761
rect -9150 -12795 -9138 -12761
rect -9196 -12829 -9138 -12795
rect -9196 -12863 -9184 -12829
rect -9150 -12863 -9138 -12829
rect -9196 -12897 -9138 -12863
rect -9196 -12931 -9184 -12897
rect -9150 -12931 -9138 -12897
rect -9196 -12965 -9138 -12931
rect -9196 -12999 -9184 -12965
rect -9150 -12999 -9138 -12965
rect -9196 -13033 -9138 -12999
rect -9196 -13067 -9184 -13033
rect -9150 -13067 -9138 -13033
rect -9196 -13112 -9138 -13067
rect -8178 -12557 -8120 -12512
rect -8178 -12591 -8166 -12557
rect -8132 -12591 -8120 -12557
rect -8178 -12625 -8120 -12591
rect -8178 -12659 -8166 -12625
rect -8132 -12659 -8120 -12625
rect -8178 -12693 -8120 -12659
rect -8178 -12727 -8166 -12693
rect -8132 -12727 -8120 -12693
rect -8178 -12761 -8120 -12727
rect -8178 -12795 -8166 -12761
rect -8132 -12795 -8120 -12761
rect -8178 -12829 -8120 -12795
rect -8178 -12863 -8166 -12829
rect -8132 -12863 -8120 -12829
rect -8178 -12897 -8120 -12863
rect -8178 -12931 -8166 -12897
rect -8132 -12931 -8120 -12897
rect -8178 -12965 -8120 -12931
rect -8178 -12999 -8166 -12965
rect -8132 -12999 -8120 -12965
rect -8178 -13033 -8120 -12999
rect -8178 -13067 -8166 -13033
rect -8132 -13067 -8120 -13033
rect -8178 -13112 -8120 -13067
rect -7160 -12557 -7102 -12512
rect -7160 -12591 -7148 -12557
rect -7114 -12591 -7102 -12557
rect -7160 -12625 -7102 -12591
rect -7160 -12659 -7148 -12625
rect -7114 -12659 -7102 -12625
rect -7160 -12693 -7102 -12659
rect -7160 -12727 -7148 -12693
rect -7114 -12727 -7102 -12693
rect -7160 -12761 -7102 -12727
rect -7160 -12795 -7148 -12761
rect -7114 -12795 -7102 -12761
rect -7160 -12829 -7102 -12795
rect -7160 -12863 -7148 -12829
rect -7114 -12863 -7102 -12829
rect -7160 -12897 -7102 -12863
rect -7160 -12931 -7148 -12897
rect -7114 -12931 -7102 -12897
rect -7160 -12965 -7102 -12931
rect -7160 -12999 -7148 -12965
rect -7114 -12999 -7102 -12965
rect -7160 -13033 -7102 -12999
rect -7160 -13067 -7148 -13033
rect -7114 -13067 -7102 -13033
rect -7160 -13112 -7102 -13067
rect -6142 -12557 -6084 -12512
rect -6142 -12591 -6130 -12557
rect -6096 -12591 -6084 -12557
rect -6142 -12625 -6084 -12591
rect -6142 -12659 -6130 -12625
rect -6096 -12659 -6084 -12625
rect -6142 -12693 -6084 -12659
rect -6142 -12727 -6130 -12693
rect -6096 -12727 -6084 -12693
rect -6142 -12761 -6084 -12727
rect -6142 -12795 -6130 -12761
rect -6096 -12795 -6084 -12761
rect -6142 -12829 -6084 -12795
rect -6142 -12863 -6130 -12829
rect -6096 -12863 -6084 -12829
rect -6142 -12897 -6084 -12863
rect -6142 -12931 -6130 -12897
rect -6096 -12931 -6084 -12897
rect -6142 -12965 -6084 -12931
rect -6142 -12999 -6130 -12965
rect -6096 -12999 -6084 -12965
rect -6142 -13033 -6084 -12999
rect -6142 -13067 -6130 -13033
rect -6096 -13067 -6084 -13033
rect -6142 -13112 -6084 -13067
rect -5124 -12557 -5066 -12512
rect -5124 -12591 -5112 -12557
rect -5078 -12591 -5066 -12557
rect -5124 -12625 -5066 -12591
rect -5124 -12659 -5112 -12625
rect -5078 -12659 -5066 -12625
rect -5124 -12693 -5066 -12659
rect -5124 -12727 -5112 -12693
rect -5078 -12727 -5066 -12693
rect -5124 -12761 -5066 -12727
rect -5124 -12795 -5112 -12761
rect -5078 -12795 -5066 -12761
rect -5124 -12829 -5066 -12795
rect -5124 -12863 -5112 -12829
rect -5078 -12863 -5066 -12829
rect -5124 -12897 -5066 -12863
rect -5124 -12931 -5112 -12897
rect -5078 -12931 -5066 -12897
rect -5124 -12965 -5066 -12931
rect -5124 -12999 -5112 -12965
rect -5078 -12999 -5066 -12965
rect -5124 -13033 -5066 -12999
rect -5124 -13067 -5112 -13033
rect -5078 -13067 -5066 -13033
rect -5124 -13112 -5066 -13067
rect -4106 -12557 -4048 -12512
rect -4106 -12591 -4094 -12557
rect -4060 -12591 -4048 -12557
rect -4106 -12625 -4048 -12591
rect -4106 -12659 -4094 -12625
rect -4060 -12659 -4048 -12625
rect -4106 -12693 -4048 -12659
rect -4106 -12727 -4094 -12693
rect -4060 -12727 -4048 -12693
rect -4106 -12761 -4048 -12727
rect -4106 -12795 -4094 -12761
rect -4060 -12795 -4048 -12761
rect -4106 -12829 -4048 -12795
rect -4106 -12863 -4094 -12829
rect -4060 -12863 -4048 -12829
rect -4106 -12897 -4048 -12863
rect -4106 -12931 -4094 -12897
rect -4060 -12931 -4048 -12897
rect -4106 -12965 -4048 -12931
rect -4106 -12999 -4094 -12965
rect -4060 -12999 -4048 -12965
rect -4106 -13033 -4048 -12999
rect -4106 -13067 -4094 -13033
rect -4060 -13067 -4048 -13033
rect -4106 -13112 -4048 -13067
rect -3088 -12557 -3030 -12512
rect -3088 -12591 -3076 -12557
rect -3042 -12591 -3030 -12557
rect -3088 -12625 -3030 -12591
rect -3088 -12659 -3076 -12625
rect -3042 -12659 -3030 -12625
rect -3088 -12693 -3030 -12659
rect -3088 -12727 -3076 -12693
rect -3042 -12727 -3030 -12693
rect -3088 -12761 -3030 -12727
rect -3088 -12795 -3076 -12761
rect -3042 -12795 -3030 -12761
rect -3088 -12829 -3030 -12795
rect -3088 -12863 -3076 -12829
rect -3042 -12863 -3030 -12829
rect -3088 -12897 -3030 -12863
rect -3088 -12931 -3076 -12897
rect -3042 -12931 -3030 -12897
rect -3088 -12965 -3030 -12931
rect -3088 -12999 -3076 -12965
rect -3042 -12999 -3030 -12965
rect -3088 -13033 -3030 -12999
rect -3088 -13067 -3076 -13033
rect -3042 -13067 -3030 -13033
rect -3088 -13112 -3030 -13067
rect -2070 -12557 -2012 -12512
rect -2070 -12591 -2058 -12557
rect -2024 -12591 -2012 -12557
rect -2070 -12625 -2012 -12591
rect -2070 -12659 -2058 -12625
rect -2024 -12659 -2012 -12625
rect -2070 -12693 -2012 -12659
rect -2070 -12727 -2058 -12693
rect -2024 -12727 -2012 -12693
rect -2070 -12761 -2012 -12727
rect -2070 -12795 -2058 -12761
rect -2024 -12795 -2012 -12761
rect -2070 -12829 -2012 -12795
rect -2070 -12863 -2058 -12829
rect -2024 -12863 -2012 -12829
rect -2070 -12897 -2012 -12863
rect -2070 -12931 -2058 -12897
rect -2024 -12931 -2012 -12897
rect -2070 -12965 -2012 -12931
rect -2070 -12999 -2058 -12965
rect -2024 -12999 -2012 -12965
rect -2070 -13033 -2012 -12999
rect -2070 -13067 -2058 -13033
rect -2024 -13067 -2012 -13033
rect -2070 -13112 -2012 -13067
rect -1052 -12557 -994 -12512
rect -1052 -12591 -1040 -12557
rect -1006 -12591 -994 -12557
rect -1052 -12625 -994 -12591
rect -1052 -12659 -1040 -12625
rect -1006 -12659 -994 -12625
rect -1052 -12693 -994 -12659
rect -1052 -12727 -1040 -12693
rect -1006 -12727 -994 -12693
rect -1052 -12761 -994 -12727
rect -1052 -12795 -1040 -12761
rect -1006 -12795 -994 -12761
rect -1052 -12829 -994 -12795
rect -1052 -12863 -1040 -12829
rect -1006 -12863 -994 -12829
rect -1052 -12897 -994 -12863
rect -1052 -12931 -1040 -12897
rect -1006 -12931 -994 -12897
rect -1052 -12965 -994 -12931
rect -1052 -12999 -1040 -12965
rect -1006 -12999 -994 -12965
rect -1052 -13033 -994 -12999
rect -1052 -13067 -1040 -13033
rect -1006 -13067 -994 -13033
rect -1052 -13112 -994 -13067
rect -34 -12557 24 -12512
rect -34 -12591 -22 -12557
rect 12 -12591 24 -12557
rect -34 -12625 24 -12591
rect -34 -12659 -22 -12625
rect 12 -12659 24 -12625
rect -34 -12693 24 -12659
rect -34 -12727 -22 -12693
rect 12 -12727 24 -12693
rect -34 -12761 24 -12727
rect -34 -12795 -22 -12761
rect 12 -12795 24 -12761
rect -34 -12829 24 -12795
rect -34 -12863 -22 -12829
rect 12 -12863 24 -12829
rect -34 -12897 24 -12863
rect -34 -12931 -22 -12897
rect 12 -12931 24 -12897
rect -34 -12965 24 -12931
rect -34 -12999 -22 -12965
rect 12 -12999 24 -12965
rect -34 -13033 24 -12999
rect -34 -13067 -22 -13033
rect 12 -13067 24 -13033
rect -34 -13112 24 -13067
rect 2570 -12997 2628 -12952
rect 2570 -13031 2582 -12997
rect 2616 -13031 2628 -12997
rect 2570 -13065 2628 -13031
rect 2570 -13099 2582 -13065
rect 2616 -13099 2628 -13065
rect 2570 -13133 2628 -13099
rect 2570 -13167 2582 -13133
rect 2616 -13167 2628 -13133
rect 2570 -13201 2628 -13167
rect 2570 -13235 2582 -13201
rect 2616 -13235 2628 -13201
rect 2570 -13269 2628 -13235
rect 2570 -13303 2582 -13269
rect 2616 -13303 2628 -13269
rect -9196 -13375 -9138 -13330
rect -9196 -13409 -9184 -13375
rect -9150 -13409 -9138 -13375
rect -9196 -13443 -9138 -13409
rect -9196 -13477 -9184 -13443
rect -9150 -13477 -9138 -13443
rect -9196 -13511 -9138 -13477
rect -9196 -13545 -9184 -13511
rect -9150 -13545 -9138 -13511
rect -9196 -13579 -9138 -13545
rect -9196 -13613 -9184 -13579
rect -9150 -13613 -9138 -13579
rect -9196 -13647 -9138 -13613
rect -9196 -13681 -9184 -13647
rect -9150 -13681 -9138 -13647
rect -9196 -13715 -9138 -13681
rect -9196 -13749 -9184 -13715
rect -9150 -13749 -9138 -13715
rect -9196 -13783 -9138 -13749
rect -9196 -13817 -9184 -13783
rect -9150 -13817 -9138 -13783
rect -9196 -13851 -9138 -13817
rect -9196 -13885 -9184 -13851
rect -9150 -13885 -9138 -13851
rect -9196 -13930 -9138 -13885
rect -8178 -13375 -8120 -13330
rect -8178 -13409 -8166 -13375
rect -8132 -13409 -8120 -13375
rect -8178 -13443 -8120 -13409
rect -8178 -13477 -8166 -13443
rect -8132 -13477 -8120 -13443
rect -8178 -13511 -8120 -13477
rect -8178 -13545 -8166 -13511
rect -8132 -13545 -8120 -13511
rect -8178 -13579 -8120 -13545
rect -8178 -13613 -8166 -13579
rect -8132 -13613 -8120 -13579
rect -8178 -13647 -8120 -13613
rect -8178 -13681 -8166 -13647
rect -8132 -13681 -8120 -13647
rect -8178 -13715 -8120 -13681
rect -8178 -13749 -8166 -13715
rect -8132 -13749 -8120 -13715
rect -8178 -13783 -8120 -13749
rect -8178 -13817 -8166 -13783
rect -8132 -13817 -8120 -13783
rect -8178 -13851 -8120 -13817
rect -8178 -13885 -8166 -13851
rect -8132 -13885 -8120 -13851
rect -8178 -13930 -8120 -13885
rect -7160 -13375 -7102 -13330
rect -7160 -13409 -7148 -13375
rect -7114 -13409 -7102 -13375
rect -7160 -13443 -7102 -13409
rect -7160 -13477 -7148 -13443
rect -7114 -13477 -7102 -13443
rect -7160 -13511 -7102 -13477
rect -7160 -13545 -7148 -13511
rect -7114 -13545 -7102 -13511
rect -7160 -13579 -7102 -13545
rect -7160 -13613 -7148 -13579
rect -7114 -13613 -7102 -13579
rect -7160 -13647 -7102 -13613
rect -7160 -13681 -7148 -13647
rect -7114 -13681 -7102 -13647
rect -7160 -13715 -7102 -13681
rect -7160 -13749 -7148 -13715
rect -7114 -13749 -7102 -13715
rect -7160 -13783 -7102 -13749
rect -7160 -13817 -7148 -13783
rect -7114 -13817 -7102 -13783
rect -7160 -13851 -7102 -13817
rect -7160 -13885 -7148 -13851
rect -7114 -13885 -7102 -13851
rect -7160 -13930 -7102 -13885
rect -6142 -13375 -6084 -13330
rect -6142 -13409 -6130 -13375
rect -6096 -13409 -6084 -13375
rect -6142 -13443 -6084 -13409
rect -6142 -13477 -6130 -13443
rect -6096 -13477 -6084 -13443
rect -6142 -13511 -6084 -13477
rect -6142 -13545 -6130 -13511
rect -6096 -13545 -6084 -13511
rect -6142 -13579 -6084 -13545
rect -6142 -13613 -6130 -13579
rect -6096 -13613 -6084 -13579
rect -6142 -13647 -6084 -13613
rect -6142 -13681 -6130 -13647
rect -6096 -13681 -6084 -13647
rect -6142 -13715 -6084 -13681
rect -6142 -13749 -6130 -13715
rect -6096 -13749 -6084 -13715
rect -6142 -13783 -6084 -13749
rect -6142 -13817 -6130 -13783
rect -6096 -13817 -6084 -13783
rect -6142 -13851 -6084 -13817
rect -6142 -13885 -6130 -13851
rect -6096 -13885 -6084 -13851
rect -6142 -13930 -6084 -13885
rect -5124 -13375 -5066 -13330
rect -5124 -13409 -5112 -13375
rect -5078 -13409 -5066 -13375
rect -5124 -13443 -5066 -13409
rect -5124 -13477 -5112 -13443
rect -5078 -13477 -5066 -13443
rect -5124 -13511 -5066 -13477
rect -5124 -13545 -5112 -13511
rect -5078 -13545 -5066 -13511
rect -5124 -13579 -5066 -13545
rect -5124 -13613 -5112 -13579
rect -5078 -13613 -5066 -13579
rect -5124 -13647 -5066 -13613
rect -5124 -13681 -5112 -13647
rect -5078 -13681 -5066 -13647
rect -5124 -13715 -5066 -13681
rect -5124 -13749 -5112 -13715
rect -5078 -13749 -5066 -13715
rect -5124 -13783 -5066 -13749
rect -5124 -13817 -5112 -13783
rect -5078 -13817 -5066 -13783
rect -5124 -13851 -5066 -13817
rect -5124 -13885 -5112 -13851
rect -5078 -13885 -5066 -13851
rect -5124 -13930 -5066 -13885
rect -4106 -13375 -4048 -13330
rect -4106 -13409 -4094 -13375
rect -4060 -13409 -4048 -13375
rect -4106 -13443 -4048 -13409
rect -4106 -13477 -4094 -13443
rect -4060 -13477 -4048 -13443
rect -4106 -13511 -4048 -13477
rect -4106 -13545 -4094 -13511
rect -4060 -13545 -4048 -13511
rect -4106 -13579 -4048 -13545
rect -4106 -13613 -4094 -13579
rect -4060 -13613 -4048 -13579
rect -4106 -13647 -4048 -13613
rect -4106 -13681 -4094 -13647
rect -4060 -13681 -4048 -13647
rect -4106 -13715 -4048 -13681
rect -4106 -13749 -4094 -13715
rect -4060 -13749 -4048 -13715
rect -4106 -13783 -4048 -13749
rect -4106 -13817 -4094 -13783
rect -4060 -13817 -4048 -13783
rect -4106 -13851 -4048 -13817
rect -4106 -13885 -4094 -13851
rect -4060 -13885 -4048 -13851
rect -4106 -13930 -4048 -13885
rect -3088 -13375 -3030 -13330
rect -3088 -13409 -3076 -13375
rect -3042 -13409 -3030 -13375
rect -3088 -13443 -3030 -13409
rect -3088 -13477 -3076 -13443
rect -3042 -13477 -3030 -13443
rect -3088 -13511 -3030 -13477
rect -3088 -13545 -3076 -13511
rect -3042 -13545 -3030 -13511
rect -3088 -13579 -3030 -13545
rect -3088 -13613 -3076 -13579
rect -3042 -13613 -3030 -13579
rect -3088 -13647 -3030 -13613
rect -3088 -13681 -3076 -13647
rect -3042 -13681 -3030 -13647
rect -3088 -13715 -3030 -13681
rect -3088 -13749 -3076 -13715
rect -3042 -13749 -3030 -13715
rect -3088 -13783 -3030 -13749
rect -3088 -13817 -3076 -13783
rect -3042 -13817 -3030 -13783
rect -3088 -13851 -3030 -13817
rect -3088 -13885 -3076 -13851
rect -3042 -13885 -3030 -13851
rect -3088 -13930 -3030 -13885
rect -2070 -13375 -2012 -13330
rect -2070 -13409 -2058 -13375
rect -2024 -13409 -2012 -13375
rect -2070 -13443 -2012 -13409
rect -2070 -13477 -2058 -13443
rect -2024 -13477 -2012 -13443
rect -2070 -13511 -2012 -13477
rect -2070 -13545 -2058 -13511
rect -2024 -13545 -2012 -13511
rect -2070 -13579 -2012 -13545
rect -2070 -13613 -2058 -13579
rect -2024 -13613 -2012 -13579
rect -2070 -13647 -2012 -13613
rect -2070 -13681 -2058 -13647
rect -2024 -13681 -2012 -13647
rect -2070 -13715 -2012 -13681
rect -2070 -13749 -2058 -13715
rect -2024 -13749 -2012 -13715
rect -2070 -13783 -2012 -13749
rect -2070 -13817 -2058 -13783
rect -2024 -13817 -2012 -13783
rect -2070 -13851 -2012 -13817
rect -2070 -13885 -2058 -13851
rect -2024 -13885 -2012 -13851
rect -2070 -13930 -2012 -13885
rect -1052 -13375 -994 -13330
rect -1052 -13409 -1040 -13375
rect -1006 -13409 -994 -13375
rect -1052 -13443 -994 -13409
rect -1052 -13477 -1040 -13443
rect -1006 -13477 -994 -13443
rect -1052 -13511 -994 -13477
rect -1052 -13545 -1040 -13511
rect -1006 -13545 -994 -13511
rect -1052 -13579 -994 -13545
rect -1052 -13613 -1040 -13579
rect -1006 -13613 -994 -13579
rect -1052 -13647 -994 -13613
rect -1052 -13681 -1040 -13647
rect -1006 -13681 -994 -13647
rect -1052 -13715 -994 -13681
rect -1052 -13749 -1040 -13715
rect -1006 -13749 -994 -13715
rect -1052 -13783 -994 -13749
rect -1052 -13817 -1040 -13783
rect -1006 -13817 -994 -13783
rect -1052 -13851 -994 -13817
rect -1052 -13885 -1040 -13851
rect -1006 -13885 -994 -13851
rect -1052 -13930 -994 -13885
rect -34 -13375 24 -13330
rect -34 -13409 -22 -13375
rect 12 -13409 24 -13375
rect -34 -13443 24 -13409
rect -34 -13477 -22 -13443
rect 12 -13477 24 -13443
rect -34 -13511 24 -13477
rect -34 -13545 -22 -13511
rect 12 -13545 24 -13511
rect -34 -13579 24 -13545
rect 2570 -13337 2628 -13303
rect 2570 -13371 2582 -13337
rect 2616 -13371 2628 -13337
rect 2570 -13405 2628 -13371
rect 2570 -13439 2582 -13405
rect 2616 -13439 2628 -13405
rect 2570 -13473 2628 -13439
rect 2570 -13507 2582 -13473
rect 2616 -13507 2628 -13473
rect 2570 -13552 2628 -13507
rect 3588 -12997 3646 -12952
rect 3588 -13031 3600 -12997
rect 3634 -13031 3646 -12997
rect 3588 -13065 3646 -13031
rect 3588 -13099 3600 -13065
rect 3634 -13099 3646 -13065
rect 3588 -13133 3646 -13099
rect 3588 -13167 3600 -13133
rect 3634 -13167 3646 -13133
rect 3588 -13201 3646 -13167
rect 3588 -13235 3600 -13201
rect 3634 -13235 3646 -13201
rect 3588 -13269 3646 -13235
rect 3588 -13303 3600 -13269
rect 3634 -13303 3646 -13269
rect 3588 -13337 3646 -13303
rect 3588 -13371 3600 -13337
rect 3634 -13371 3646 -13337
rect 3588 -13405 3646 -13371
rect 3588 -13439 3600 -13405
rect 3634 -13439 3646 -13405
rect 3588 -13473 3646 -13439
rect 3588 -13507 3600 -13473
rect 3634 -13507 3646 -13473
rect 3588 -13552 3646 -13507
rect 4606 -12997 4664 -12952
rect 4606 -13031 4618 -12997
rect 4652 -13031 4664 -12997
rect 4606 -13065 4664 -13031
rect 4606 -13099 4618 -13065
rect 4652 -13099 4664 -13065
rect 4606 -13133 4664 -13099
rect 4606 -13167 4618 -13133
rect 4652 -13167 4664 -13133
rect 4606 -13201 4664 -13167
rect 4606 -13235 4618 -13201
rect 4652 -13235 4664 -13201
rect 4606 -13269 4664 -13235
rect 4606 -13303 4618 -13269
rect 4652 -13303 4664 -13269
rect 4606 -13337 4664 -13303
rect 4606 -13371 4618 -13337
rect 4652 -13371 4664 -13337
rect 4606 -13405 4664 -13371
rect 4606 -13439 4618 -13405
rect 4652 -13439 4664 -13405
rect 4606 -13473 4664 -13439
rect 4606 -13507 4618 -13473
rect 4652 -13507 4664 -13473
rect 4606 -13552 4664 -13507
rect 5624 -12997 5682 -12952
rect 5624 -13031 5636 -12997
rect 5670 -13031 5682 -12997
rect 5624 -13065 5682 -13031
rect 5624 -13099 5636 -13065
rect 5670 -13099 5682 -13065
rect 5624 -13133 5682 -13099
rect 5624 -13167 5636 -13133
rect 5670 -13167 5682 -13133
rect 5624 -13201 5682 -13167
rect 5624 -13235 5636 -13201
rect 5670 -13235 5682 -13201
rect 5624 -13269 5682 -13235
rect 5624 -13303 5636 -13269
rect 5670 -13303 5682 -13269
rect 5624 -13337 5682 -13303
rect 5624 -13371 5636 -13337
rect 5670 -13371 5682 -13337
rect 5624 -13405 5682 -13371
rect 5624 -13439 5636 -13405
rect 5670 -13439 5682 -13405
rect 5624 -13473 5682 -13439
rect 5624 -13507 5636 -13473
rect 5670 -13507 5682 -13473
rect 5624 -13552 5682 -13507
rect 6642 -12997 6700 -12952
rect 6642 -13031 6654 -12997
rect 6688 -13031 6700 -12997
rect 6642 -13065 6700 -13031
rect 6642 -13099 6654 -13065
rect 6688 -13099 6700 -13065
rect 6642 -13133 6700 -13099
rect 6642 -13167 6654 -13133
rect 6688 -13167 6700 -13133
rect 6642 -13201 6700 -13167
rect 6642 -13235 6654 -13201
rect 6688 -13235 6700 -13201
rect 6642 -13269 6700 -13235
rect 6642 -13303 6654 -13269
rect 6688 -13303 6700 -13269
rect 6642 -13337 6700 -13303
rect 6642 -13371 6654 -13337
rect 6688 -13371 6700 -13337
rect 6642 -13405 6700 -13371
rect 6642 -13439 6654 -13405
rect 6688 -13439 6700 -13405
rect 6642 -13473 6700 -13439
rect 6642 -13507 6654 -13473
rect 6688 -13507 6700 -13473
rect 6642 -13552 6700 -13507
rect 7660 -12997 7718 -12952
rect 7660 -13031 7672 -12997
rect 7706 -13031 7718 -12997
rect 7660 -13065 7718 -13031
rect 7660 -13099 7672 -13065
rect 7706 -13099 7718 -13065
rect 7660 -13133 7718 -13099
rect 7660 -13167 7672 -13133
rect 7706 -13167 7718 -13133
rect 7660 -13201 7718 -13167
rect 7660 -13235 7672 -13201
rect 7706 -13235 7718 -13201
rect 7660 -13269 7718 -13235
rect 7660 -13303 7672 -13269
rect 7706 -13303 7718 -13269
rect 7660 -13337 7718 -13303
rect 7660 -13371 7672 -13337
rect 7706 -13371 7718 -13337
rect 7660 -13405 7718 -13371
rect 7660 -13439 7672 -13405
rect 7706 -13439 7718 -13405
rect 7660 -13473 7718 -13439
rect 7660 -13507 7672 -13473
rect 7706 -13507 7718 -13473
rect 7660 -13552 7718 -13507
rect 8678 -12997 8736 -12952
rect 8678 -13031 8690 -12997
rect 8724 -13031 8736 -12997
rect 8678 -13065 8736 -13031
rect 8678 -13099 8690 -13065
rect 8724 -13099 8736 -13065
rect 8678 -13133 8736 -13099
rect 8678 -13167 8690 -13133
rect 8724 -13167 8736 -13133
rect 8678 -13201 8736 -13167
rect 8678 -13235 8690 -13201
rect 8724 -13235 8736 -13201
rect 8678 -13269 8736 -13235
rect 8678 -13303 8690 -13269
rect 8724 -13303 8736 -13269
rect 8678 -13337 8736 -13303
rect 8678 -13371 8690 -13337
rect 8724 -13371 8736 -13337
rect 8678 -13405 8736 -13371
rect 8678 -13439 8690 -13405
rect 8724 -13439 8736 -13405
rect 8678 -13473 8736 -13439
rect 8678 -13507 8690 -13473
rect 8724 -13507 8736 -13473
rect 8678 -13552 8736 -13507
rect 9696 -12997 9754 -12952
rect 9696 -13031 9708 -12997
rect 9742 -13031 9754 -12997
rect 9696 -13065 9754 -13031
rect 9696 -13099 9708 -13065
rect 9742 -13099 9754 -13065
rect 9696 -13133 9754 -13099
rect 9696 -13167 9708 -13133
rect 9742 -13167 9754 -13133
rect 9696 -13201 9754 -13167
rect 9696 -13235 9708 -13201
rect 9742 -13235 9754 -13201
rect 9696 -13269 9754 -13235
rect 9696 -13303 9708 -13269
rect 9742 -13303 9754 -13269
rect 9696 -13337 9754 -13303
rect 9696 -13371 9708 -13337
rect 9742 -13371 9754 -13337
rect 9696 -13405 9754 -13371
rect 9696 -13439 9708 -13405
rect 9742 -13439 9754 -13405
rect 9696 -13473 9754 -13439
rect 9696 -13507 9708 -13473
rect 9742 -13507 9754 -13473
rect 9696 -13552 9754 -13507
rect 10714 -12997 10772 -12952
rect 10714 -13031 10726 -12997
rect 10760 -13031 10772 -12997
rect 10714 -13065 10772 -13031
rect 10714 -13099 10726 -13065
rect 10760 -13099 10772 -13065
rect 10714 -13133 10772 -13099
rect 10714 -13167 10726 -13133
rect 10760 -13167 10772 -13133
rect 10714 -13201 10772 -13167
rect 10714 -13235 10726 -13201
rect 10760 -13235 10772 -13201
rect 10714 -13269 10772 -13235
rect 10714 -13303 10726 -13269
rect 10760 -13303 10772 -13269
rect 10714 -13337 10772 -13303
rect 10714 -13371 10726 -13337
rect 10760 -13371 10772 -13337
rect 10714 -13405 10772 -13371
rect 10714 -13439 10726 -13405
rect 10760 -13439 10772 -13405
rect 10714 -13473 10772 -13439
rect 10714 -13507 10726 -13473
rect 10760 -13507 10772 -13473
rect 10714 -13552 10772 -13507
rect 11732 -12997 11790 -12952
rect 11732 -13031 11744 -12997
rect 11778 -13031 11790 -12997
rect 11732 -13065 11790 -13031
rect 11732 -13099 11744 -13065
rect 11778 -13099 11790 -13065
rect 11732 -13133 11790 -13099
rect 11732 -13167 11744 -13133
rect 11778 -13167 11790 -13133
rect 11732 -13201 11790 -13167
rect 11732 -13235 11744 -13201
rect 11778 -13235 11790 -13201
rect 11732 -13269 11790 -13235
rect 11732 -13303 11744 -13269
rect 11778 -13303 11790 -13269
rect 11732 -13337 11790 -13303
rect 11732 -13371 11744 -13337
rect 11778 -13371 11790 -13337
rect 11732 -13405 11790 -13371
rect 11732 -13439 11744 -13405
rect 11778 -13439 11790 -13405
rect 11732 -13473 11790 -13439
rect 11732 -13507 11744 -13473
rect 11778 -13507 11790 -13473
rect 11732 -13552 11790 -13507
rect 12750 -12997 12808 -12952
rect 12750 -13031 12762 -12997
rect 12796 -13031 12808 -12997
rect 12750 -13065 12808 -13031
rect 12750 -13099 12762 -13065
rect 12796 -13099 12808 -13065
rect 12750 -13133 12808 -13099
rect 12750 -13167 12762 -13133
rect 12796 -13167 12808 -13133
rect 12750 -13201 12808 -13167
rect 12750 -13235 12762 -13201
rect 12796 -13235 12808 -13201
rect 12750 -13269 12808 -13235
rect 12750 -13303 12762 -13269
rect 12796 -13303 12808 -13269
rect 12750 -13337 12808 -13303
rect 12750 -13371 12762 -13337
rect 12796 -13371 12808 -13337
rect 12750 -13405 12808 -13371
rect 12750 -13439 12762 -13405
rect 12796 -13439 12808 -13405
rect 12750 -13473 12808 -13439
rect 12750 -13507 12762 -13473
rect 12796 -13507 12808 -13473
rect 12750 -13552 12808 -13507
rect 13768 -12997 13826 -12952
rect 13768 -13031 13780 -12997
rect 13814 -13031 13826 -12997
rect 13768 -13065 13826 -13031
rect 13768 -13099 13780 -13065
rect 13814 -13099 13826 -13065
rect 13768 -13133 13826 -13099
rect 13768 -13167 13780 -13133
rect 13814 -13167 13826 -13133
rect 13768 -13201 13826 -13167
rect 13768 -13235 13780 -13201
rect 13814 -13235 13826 -13201
rect 13768 -13269 13826 -13235
rect 13768 -13303 13780 -13269
rect 13814 -13303 13826 -13269
rect 13768 -13337 13826 -13303
rect 13768 -13371 13780 -13337
rect 13814 -13371 13826 -13337
rect 13768 -13405 13826 -13371
rect 13768 -13439 13780 -13405
rect 13814 -13439 13826 -13405
rect 13768 -13473 13826 -13439
rect 13768 -13507 13780 -13473
rect 13814 -13507 13826 -13473
rect 13768 -13552 13826 -13507
rect 14786 -12997 14844 -12952
rect 14786 -13031 14798 -12997
rect 14832 -13031 14844 -12997
rect 14786 -13065 14844 -13031
rect 14786 -13099 14798 -13065
rect 14832 -13099 14844 -13065
rect 14786 -13133 14844 -13099
rect 14786 -13167 14798 -13133
rect 14832 -13167 14844 -13133
rect 14786 -13201 14844 -13167
rect 14786 -13235 14798 -13201
rect 14832 -13235 14844 -13201
rect 14786 -13269 14844 -13235
rect 14786 -13303 14798 -13269
rect 14832 -13303 14844 -13269
rect 14786 -13337 14844 -13303
rect 14786 -13371 14798 -13337
rect 14832 -13371 14844 -13337
rect 14786 -13405 14844 -13371
rect 14786 -13439 14798 -13405
rect 14832 -13439 14844 -13405
rect 14786 -13473 14844 -13439
rect 14786 -13507 14798 -13473
rect 14832 -13507 14844 -13473
rect 14786 -13552 14844 -13507
rect 15804 -12997 15862 -12952
rect 15804 -13031 15816 -12997
rect 15850 -13031 15862 -12997
rect 15804 -13065 15862 -13031
rect 15804 -13099 15816 -13065
rect 15850 -13099 15862 -13065
rect 15804 -13133 15862 -13099
rect 15804 -13167 15816 -13133
rect 15850 -13167 15862 -13133
rect 15804 -13201 15862 -13167
rect 15804 -13235 15816 -13201
rect 15850 -13235 15862 -13201
rect 15804 -13269 15862 -13235
rect 15804 -13303 15816 -13269
rect 15850 -13303 15862 -13269
rect 15804 -13337 15862 -13303
rect 15804 -13371 15816 -13337
rect 15850 -13371 15862 -13337
rect 15804 -13405 15862 -13371
rect 15804 -13439 15816 -13405
rect 15850 -13439 15862 -13405
rect 15804 -13473 15862 -13439
rect 15804 -13507 15816 -13473
rect 15850 -13507 15862 -13473
rect 15804 -13552 15862 -13507
rect 16822 -12997 16880 -12952
rect 16822 -13031 16834 -12997
rect 16868 -13031 16880 -12997
rect 16822 -13065 16880 -13031
rect 16822 -13099 16834 -13065
rect 16868 -13099 16880 -13065
rect 16822 -13133 16880 -13099
rect 16822 -13167 16834 -13133
rect 16868 -13167 16880 -13133
rect 16822 -13201 16880 -13167
rect 16822 -13235 16834 -13201
rect 16868 -13235 16880 -13201
rect 16822 -13269 16880 -13235
rect 16822 -13303 16834 -13269
rect 16868 -13303 16880 -13269
rect 16822 -13337 16880 -13303
rect 16822 -13371 16834 -13337
rect 16868 -13371 16880 -13337
rect 16822 -13405 16880 -13371
rect 16822 -13439 16834 -13405
rect 16868 -13439 16880 -13405
rect 16822 -13473 16880 -13439
rect 16822 -13507 16834 -13473
rect 16868 -13507 16880 -13473
rect 16822 -13552 16880 -13507
rect 17840 -12997 17898 -12952
rect 17840 -13031 17852 -12997
rect 17886 -13031 17898 -12997
rect 17840 -13065 17898 -13031
rect 17840 -13099 17852 -13065
rect 17886 -13099 17898 -13065
rect 17840 -13133 17898 -13099
rect 17840 -13167 17852 -13133
rect 17886 -13167 17898 -13133
rect 17840 -13201 17898 -13167
rect 17840 -13235 17852 -13201
rect 17886 -13235 17898 -13201
rect 17840 -13269 17898 -13235
rect 17840 -13303 17852 -13269
rect 17886 -13303 17898 -13269
rect 17840 -13337 17898 -13303
rect 17840 -13371 17852 -13337
rect 17886 -13371 17898 -13337
rect 17840 -13405 17898 -13371
rect 17840 -13439 17852 -13405
rect 17886 -13439 17898 -13405
rect 17840 -13473 17898 -13439
rect 17840 -13507 17852 -13473
rect 17886 -13507 17898 -13473
rect 17840 -13552 17898 -13507
rect 18858 -12997 18916 -12952
rect 18858 -13031 18870 -12997
rect 18904 -13031 18916 -12997
rect 18858 -13065 18916 -13031
rect 18858 -13099 18870 -13065
rect 18904 -13099 18916 -13065
rect 18858 -13133 18916 -13099
rect 18858 -13167 18870 -13133
rect 18904 -13167 18916 -13133
rect 18858 -13201 18916 -13167
rect 18858 -13235 18870 -13201
rect 18904 -13235 18916 -13201
rect 18858 -13269 18916 -13235
rect 18858 -13303 18870 -13269
rect 18904 -13303 18916 -13269
rect 18858 -13337 18916 -13303
rect 18858 -13371 18870 -13337
rect 18904 -13371 18916 -13337
rect 18858 -13405 18916 -13371
rect 18858 -13439 18870 -13405
rect 18904 -13439 18916 -13405
rect 18858 -13473 18916 -13439
rect 18858 -13507 18870 -13473
rect 18904 -13507 18916 -13473
rect 18858 -13552 18916 -13507
rect 19876 -12997 19934 -12952
rect 19876 -13031 19888 -12997
rect 19922 -13031 19934 -12997
rect 19876 -13065 19934 -13031
rect 19876 -13099 19888 -13065
rect 19922 -13099 19934 -13065
rect 19876 -13133 19934 -13099
rect 19876 -13167 19888 -13133
rect 19922 -13167 19934 -13133
rect 19876 -13201 19934 -13167
rect 19876 -13235 19888 -13201
rect 19922 -13235 19934 -13201
rect 19876 -13269 19934 -13235
rect 19876 -13303 19888 -13269
rect 19922 -13303 19934 -13269
rect 19876 -13337 19934 -13303
rect 19876 -13371 19888 -13337
rect 19922 -13371 19934 -13337
rect 19876 -13405 19934 -13371
rect 19876 -13439 19888 -13405
rect 19922 -13439 19934 -13405
rect 19876 -13473 19934 -13439
rect 19876 -13507 19888 -13473
rect 19922 -13507 19934 -13473
rect 19876 -13552 19934 -13507
rect 20894 -12997 20952 -12952
rect 20894 -13031 20906 -12997
rect 20940 -13031 20952 -12997
rect 20894 -13065 20952 -13031
rect 20894 -13099 20906 -13065
rect 20940 -13099 20952 -13065
rect 20894 -13133 20952 -13099
rect 20894 -13167 20906 -13133
rect 20940 -13167 20952 -13133
rect 20894 -13201 20952 -13167
rect 20894 -13235 20906 -13201
rect 20940 -13235 20952 -13201
rect 20894 -13269 20952 -13235
rect 20894 -13303 20906 -13269
rect 20940 -13303 20952 -13269
rect 20894 -13337 20952 -13303
rect 20894 -13371 20906 -13337
rect 20940 -13371 20952 -13337
rect 20894 -13405 20952 -13371
rect 20894 -13439 20906 -13405
rect 20940 -13439 20952 -13405
rect 20894 -13473 20952 -13439
rect 20894 -13507 20906 -13473
rect 20940 -13507 20952 -13473
rect 20894 -13552 20952 -13507
rect 21912 -12997 21970 -12952
rect 21912 -13031 21924 -12997
rect 21958 -13031 21970 -12997
rect 21912 -13065 21970 -13031
rect 21912 -13099 21924 -13065
rect 21958 -13099 21970 -13065
rect 21912 -13133 21970 -13099
rect 21912 -13167 21924 -13133
rect 21958 -13167 21970 -13133
rect 21912 -13201 21970 -13167
rect 21912 -13235 21924 -13201
rect 21958 -13235 21970 -13201
rect 21912 -13269 21970 -13235
rect 21912 -13303 21924 -13269
rect 21958 -13303 21970 -13269
rect 21912 -13337 21970 -13303
rect 21912 -13371 21924 -13337
rect 21958 -13371 21970 -13337
rect 21912 -13405 21970 -13371
rect 21912 -13439 21924 -13405
rect 21958 -13439 21970 -13405
rect 21912 -13473 21970 -13439
rect 21912 -13507 21924 -13473
rect 21958 -13507 21970 -13473
rect 21912 -13552 21970 -13507
rect 22930 -12997 22988 -12952
rect 22930 -13031 22942 -12997
rect 22976 -13031 22988 -12997
rect 22930 -13065 22988 -13031
rect 22930 -13099 22942 -13065
rect 22976 -13099 22988 -13065
rect 22930 -13133 22988 -13099
rect 22930 -13167 22942 -13133
rect 22976 -13167 22988 -13133
rect 22930 -13201 22988 -13167
rect 22930 -13235 22942 -13201
rect 22976 -13235 22988 -13201
rect 22930 -13269 22988 -13235
rect 22930 -13303 22942 -13269
rect 22976 -13303 22988 -13269
rect 22930 -13337 22988 -13303
rect 22930 -13371 22942 -13337
rect 22976 -13371 22988 -13337
rect 22930 -13405 22988 -13371
rect 22930 -13439 22942 -13405
rect 22976 -13439 22988 -13405
rect 22930 -13473 22988 -13439
rect 22930 -13507 22942 -13473
rect 22976 -13507 22988 -13473
rect 22930 -13552 22988 -13507
rect -34 -13613 -22 -13579
rect 12 -13613 24 -13579
rect -34 -13647 24 -13613
rect -34 -13681 -22 -13647
rect 12 -13681 24 -13647
rect -34 -13715 24 -13681
rect -34 -13749 -22 -13715
rect 12 -13749 24 -13715
rect -34 -13783 24 -13749
rect -34 -13817 -22 -13783
rect 12 -13817 24 -13783
rect -34 -13851 24 -13817
rect -34 -13885 -22 -13851
rect 12 -13885 24 -13851
rect -34 -13930 24 -13885
rect -9196 -14193 -9138 -14148
rect -9196 -14227 -9184 -14193
rect -9150 -14227 -9138 -14193
rect -9196 -14261 -9138 -14227
rect -9196 -14295 -9184 -14261
rect -9150 -14295 -9138 -14261
rect -9196 -14329 -9138 -14295
rect -9196 -14363 -9184 -14329
rect -9150 -14363 -9138 -14329
rect -9196 -14397 -9138 -14363
rect -9196 -14431 -9184 -14397
rect -9150 -14431 -9138 -14397
rect -9196 -14465 -9138 -14431
rect -9196 -14499 -9184 -14465
rect -9150 -14499 -9138 -14465
rect -9196 -14533 -9138 -14499
rect -9196 -14567 -9184 -14533
rect -9150 -14567 -9138 -14533
rect -9196 -14601 -9138 -14567
rect -9196 -14635 -9184 -14601
rect -9150 -14635 -9138 -14601
rect -9196 -14669 -9138 -14635
rect -9196 -14703 -9184 -14669
rect -9150 -14703 -9138 -14669
rect -9196 -14748 -9138 -14703
rect -8178 -14193 -8120 -14148
rect -8178 -14227 -8166 -14193
rect -8132 -14227 -8120 -14193
rect -8178 -14261 -8120 -14227
rect -8178 -14295 -8166 -14261
rect -8132 -14295 -8120 -14261
rect -8178 -14329 -8120 -14295
rect -8178 -14363 -8166 -14329
rect -8132 -14363 -8120 -14329
rect -8178 -14397 -8120 -14363
rect -8178 -14431 -8166 -14397
rect -8132 -14431 -8120 -14397
rect -8178 -14465 -8120 -14431
rect -8178 -14499 -8166 -14465
rect -8132 -14499 -8120 -14465
rect -8178 -14533 -8120 -14499
rect -8178 -14567 -8166 -14533
rect -8132 -14567 -8120 -14533
rect -8178 -14601 -8120 -14567
rect -8178 -14635 -8166 -14601
rect -8132 -14635 -8120 -14601
rect -8178 -14669 -8120 -14635
rect -8178 -14703 -8166 -14669
rect -8132 -14703 -8120 -14669
rect -8178 -14748 -8120 -14703
rect -7160 -14193 -7102 -14148
rect -7160 -14227 -7148 -14193
rect -7114 -14227 -7102 -14193
rect -7160 -14261 -7102 -14227
rect -7160 -14295 -7148 -14261
rect -7114 -14295 -7102 -14261
rect -7160 -14329 -7102 -14295
rect -7160 -14363 -7148 -14329
rect -7114 -14363 -7102 -14329
rect -7160 -14397 -7102 -14363
rect -7160 -14431 -7148 -14397
rect -7114 -14431 -7102 -14397
rect -7160 -14465 -7102 -14431
rect -7160 -14499 -7148 -14465
rect -7114 -14499 -7102 -14465
rect -7160 -14533 -7102 -14499
rect -7160 -14567 -7148 -14533
rect -7114 -14567 -7102 -14533
rect -7160 -14601 -7102 -14567
rect -7160 -14635 -7148 -14601
rect -7114 -14635 -7102 -14601
rect -7160 -14669 -7102 -14635
rect -7160 -14703 -7148 -14669
rect -7114 -14703 -7102 -14669
rect -7160 -14748 -7102 -14703
rect -6142 -14193 -6084 -14148
rect -6142 -14227 -6130 -14193
rect -6096 -14227 -6084 -14193
rect -6142 -14261 -6084 -14227
rect -6142 -14295 -6130 -14261
rect -6096 -14295 -6084 -14261
rect -6142 -14329 -6084 -14295
rect -6142 -14363 -6130 -14329
rect -6096 -14363 -6084 -14329
rect -6142 -14397 -6084 -14363
rect -6142 -14431 -6130 -14397
rect -6096 -14431 -6084 -14397
rect -6142 -14465 -6084 -14431
rect -6142 -14499 -6130 -14465
rect -6096 -14499 -6084 -14465
rect -6142 -14533 -6084 -14499
rect -6142 -14567 -6130 -14533
rect -6096 -14567 -6084 -14533
rect -6142 -14601 -6084 -14567
rect -6142 -14635 -6130 -14601
rect -6096 -14635 -6084 -14601
rect -6142 -14669 -6084 -14635
rect -6142 -14703 -6130 -14669
rect -6096 -14703 -6084 -14669
rect -6142 -14748 -6084 -14703
rect -5124 -14193 -5066 -14148
rect -5124 -14227 -5112 -14193
rect -5078 -14227 -5066 -14193
rect -5124 -14261 -5066 -14227
rect -5124 -14295 -5112 -14261
rect -5078 -14295 -5066 -14261
rect -5124 -14329 -5066 -14295
rect -5124 -14363 -5112 -14329
rect -5078 -14363 -5066 -14329
rect -5124 -14397 -5066 -14363
rect -5124 -14431 -5112 -14397
rect -5078 -14431 -5066 -14397
rect -5124 -14465 -5066 -14431
rect -5124 -14499 -5112 -14465
rect -5078 -14499 -5066 -14465
rect -5124 -14533 -5066 -14499
rect -5124 -14567 -5112 -14533
rect -5078 -14567 -5066 -14533
rect -5124 -14601 -5066 -14567
rect -5124 -14635 -5112 -14601
rect -5078 -14635 -5066 -14601
rect -5124 -14669 -5066 -14635
rect -5124 -14703 -5112 -14669
rect -5078 -14703 -5066 -14669
rect -5124 -14748 -5066 -14703
rect -4106 -14193 -4048 -14148
rect -4106 -14227 -4094 -14193
rect -4060 -14227 -4048 -14193
rect -4106 -14261 -4048 -14227
rect -4106 -14295 -4094 -14261
rect -4060 -14295 -4048 -14261
rect -4106 -14329 -4048 -14295
rect -4106 -14363 -4094 -14329
rect -4060 -14363 -4048 -14329
rect -4106 -14397 -4048 -14363
rect -4106 -14431 -4094 -14397
rect -4060 -14431 -4048 -14397
rect -4106 -14465 -4048 -14431
rect -4106 -14499 -4094 -14465
rect -4060 -14499 -4048 -14465
rect -4106 -14533 -4048 -14499
rect -4106 -14567 -4094 -14533
rect -4060 -14567 -4048 -14533
rect -4106 -14601 -4048 -14567
rect -4106 -14635 -4094 -14601
rect -4060 -14635 -4048 -14601
rect -4106 -14669 -4048 -14635
rect -4106 -14703 -4094 -14669
rect -4060 -14703 -4048 -14669
rect -4106 -14748 -4048 -14703
rect -3088 -14193 -3030 -14148
rect -3088 -14227 -3076 -14193
rect -3042 -14227 -3030 -14193
rect -3088 -14261 -3030 -14227
rect -3088 -14295 -3076 -14261
rect -3042 -14295 -3030 -14261
rect -3088 -14329 -3030 -14295
rect -3088 -14363 -3076 -14329
rect -3042 -14363 -3030 -14329
rect -3088 -14397 -3030 -14363
rect -3088 -14431 -3076 -14397
rect -3042 -14431 -3030 -14397
rect -3088 -14465 -3030 -14431
rect -3088 -14499 -3076 -14465
rect -3042 -14499 -3030 -14465
rect -3088 -14533 -3030 -14499
rect -3088 -14567 -3076 -14533
rect -3042 -14567 -3030 -14533
rect -3088 -14601 -3030 -14567
rect -3088 -14635 -3076 -14601
rect -3042 -14635 -3030 -14601
rect -3088 -14669 -3030 -14635
rect -3088 -14703 -3076 -14669
rect -3042 -14703 -3030 -14669
rect -3088 -14748 -3030 -14703
rect -2070 -14193 -2012 -14148
rect -2070 -14227 -2058 -14193
rect -2024 -14227 -2012 -14193
rect -2070 -14261 -2012 -14227
rect -2070 -14295 -2058 -14261
rect -2024 -14295 -2012 -14261
rect -2070 -14329 -2012 -14295
rect -2070 -14363 -2058 -14329
rect -2024 -14363 -2012 -14329
rect -2070 -14397 -2012 -14363
rect -2070 -14431 -2058 -14397
rect -2024 -14431 -2012 -14397
rect -2070 -14465 -2012 -14431
rect -2070 -14499 -2058 -14465
rect -2024 -14499 -2012 -14465
rect -2070 -14533 -2012 -14499
rect -2070 -14567 -2058 -14533
rect -2024 -14567 -2012 -14533
rect -2070 -14601 -2012 -14567
rect -2070 -14635 -2058 -14601
rect -2024 -14635 -2012 -14601
rect -2070 -14669 -2012 -14635
rect -2070 -14703 -2058 -14669
rect -2024 -14703 -2012 -14669
rect -2070 -14748 -2012 -14703
rect -1052 -14193 -994 -14148
rect -1052 -14227 -1040 -14193
rect -1006 -14227 -994 -14193
rect -1052 -14261 -994 -14227
rect -1052 -14295 -1040 -14261
rect -1006 -14295 -994 -14261
rect -1052 -14329 -994 -14295
rect -1052 -14363 -1040 -14329
rect -1006 -14363 -994 -14329
rect -1052 -14397 -994 -14363
rect -1052 -14431 -1040 -14397
rect -1006 -14431 -994 -14397
rect -1052 -14465 -994 -14431
rect -1052 -14499 -1040 -14465
rect -1006 -14499 -994 -14465
rect -1052 -14533 -994 -14499
rect -1052 -14567 -1040 -14533
rect -1006 -14567 -994 -14533
rect -1052 -14601 -994 -14567
rect -1052 -14635 -1040 -14601
rect -1006 -14635 -994 -14601
rect -1052 -14669 -994 -14635
rect -1052 -14703 -1040 -14669
rect -1006 -14703 -994 -14669
rect -1052 -14748 -994 -14703
rect -34 -14193 24 -14148
rect -34 -14227 -22 -14193
rect 12 -14227 24 -14193
rect -34 -14261 24 -14227
rect -34 -14295 -22 -14261
rect 12 -14295 24 -14261
rect -34 -14329 24 -14295
rect -34 -14363 -22 -14329
rect 12 -14363 24 -14329
rect -34 -14397 24 -14363
rect -34 -14431 -22 -14397
rect 12 -14431 24 -14397
rect -34 -14465 24 -14431
rect -34 -14499 -22 -14465
rect 12 -14499 24 -14465
rect -34 -14533 24 -14499
rect -34 -14567 -22 -14533
rect 12 -14567 24 -14533
rect -34 -14601 24 -14567
rect -34 -14635 -22 -14601
rect 12 -14635 24 -14601
rect -34 -14669 24 -14635
rect -34 -14703 -22 -14669
rect 12 -14703 24 -14669
rect -34 -14748 24 -14703
rect 2570 -14229 2628 -14184
rect 2570 -14263 2582 -14229
rect 2616 -14263 2628 -14229
rect 2570 -14297 2628 -14263
rect 2570 -14331 2582 -14297
rect 2616 -14331 2628 -14297
rect 2570 -14365 2628 -14331
rect 2570 -14399 2582 -14365
rect 2616 -14399 2628 -14365
rect 2570 -14433 2628 -14399
rect 2570 -14467 2582 -14433
rect 2616 -14467 2628 -14433
rect 2570 -14501 2628 -14467
rect 2570 -14535 2582 -14501
rect 2616 -14535 2628 -14501
rect 2570 -14569 2628 -14535
rect 2570 -14603 2582 -14569
rect 2616 -14603 2628 -14569
rect 2570 -14637 2628 -14603
rect 2570 -14671 2582 -14637
rect 2616 -14671 2628 -14637
rect 2570 -14705 2628 -14671
rect 2570 -14739 2582 -14705
rect 2616 -14739 2628 -14705
rect 2570 -14784 2628 -14739
rect 3588 -14229 3646 -14184
rect 3588 -14263 3600 -14229
rect 3634 -14263 3646 -14229
rect 3588 -14297 3646 -14263
rect 3588 -14331 3600 -14297
rect 3634 -14331 3646 -14297
rect 3588 -14365 3646 -14331
rect 3588 -14399 3600 -14365
rect 3634 -14399 3646 -14365
rect 3588 -14433 3646 -14399
rect 3588 -14467 3600 -14433
rect 3634 -14467 3646 -14433
rect 3588 -14501 3646 -14467
rect 3588 -14535 3600 -14501
rect 3634 -14535 3646 -14501
rect 3588 -14569 3646 -14535
rect 3588 -14603 3600 -14569
rect 3634 -14603 3646 -14569
rect 3588 -14637 3646 -14603
rect 3588 -14671 3600 -14637
rect 3634 -14671 3646 -14637
rect 3588 -14705 3646 -14671
rect 3588 -14739 3600 -14705
rect 3634 -14739 3646 -14705
rect 3588 -14784 3646 -14739
rect 4606 -14229 4664 -14184
rect 4606 -14263 4618 -14229
rect 4652 -14263 4664 -14229
rect 4606 -14297 4664 -14263
rect 4606 -14331 4618 -14297
rect 4652 -14331 4664 -14297
rect 4606 -14365 4664 -14331
rect 4606 -14399 4618 -14365
rect 4652 -14399 4664 -14365
rect 4606 -14433 4664 -14399
rect 4606 -14467 4618 -14433
rect 4652 -14467 4664 -14433
rect 4606 -14501 4664 -14467
rect 4606 -14535 4618 -14501
rect 4652 -14535 4664 -14501
rect 4606 -14569 4664 -14535
rect 4606 -14603 4618 -14569
rect 4652 -14603 4664 -14569
rect 4606 -14637 4664 -14603
rect 4606 -14671 4618 -14637
rect 4652 -14671 4664 -14637
rect 4606 -14705 4664 -14671
rect 4606 -14739 4618 -14705
rect 4652 -14739 4664 -14705
rect 4606 -14784 4664 -14739
rect 5624 -14229 5682 -14184
rect 5624 -14263 5636 -14229
rect 5670 -14263 5682 -14229
rect 5624 -14297 5682 -14263
rect 5624 -14331 5636 -14297
rect 5670 -14331 5682 -14297
rect 5624 -14365 5682 -14331
rect 5624 -14399 5636 -14365
rect 5670 -14399 5682 -14365
rect 5624 -14433 5682 -14399
rect 5624 -14467 5636 -14433
rect 5670 -14467 5682 -14433
rect 5624 -14501 5682 -14467
rect 5624 -14535 5636 -14501
rect 5670 -14535 5682 -14501
rect 5624 -14569 5682 -14535
rect 5624 -14603 5636 -14569
rect 5670 -14603 5682 -14569
rect 5624 -14637 5682 -14603
rect 5624 -14671 5636 -14637
rect 5670 -14671 5682 -14637
rect 5624 -14705 5682 -14671
rect 5624 -14739 5636 -14705
rect 5670 -14739 5682 -14705
rect 5624 -14784 5682 -14739
rect 6642 -14229 6700 -14184
rect 6642 -14263 6654 -14229
rect 6688 -14263 6700 -14229
rect 6642 -14297 6700 -14263
rect 6642 -14331 6654 -14297
rect 6688 -14331 6700 -14297
rect 6642 -14365 6700 -14331
rect 6642 -14399 6654 -14365
rect 6688 -14399 6700 -14365
rect 6642 -14433 6700 -14399
rect 6642 -14467 6654 -14433
rect 6688 -14467 6700 -14433
rect 6642 -14501 6700 -14467
rect 6642 -14535 6654 -14501
rect 6688 -14535 6700 -14501
rect 6642 -14569 6700 -14535
rect 6642 -14603 6654 -14569
rect 6688 -14603 6700 -14569
rect 6642 -14637 6700 -14603
rect 6642 -14671 6654 -14637
rect 6688 -14671 6700 -14637
rect 6642 -14705 6700 -14671
rect 6642 -14739 6654 -14705
rect 6688 -14739 6700 -14705
rect 6642 -14784 6700 -14739
rect 7660 -14229 7718 -14184
rect 7660 -14263 7672 -14229
rect 7706 -14263 7718 -14229
rect 7660 -14297 7718 -14263
rect 7660 -14331 7672 -14297
rect 7706 -14331 7718 -14297
rect 7660 -14365 7718 -14331
rect 7660 -14399 7672 -14365
rect 7706 -14399 7718 -14365
rect 7660 -14433 7718 -14399
rect 7660 -14467 7672 -14433
rect 7706 -14467 7718 -14433
rect 7660 -14501 7718 -14467
rect 7660 -14535 7672 -14501
rect 7706 -14535 7718 -14501
rect 7660 -14569 7718 -14535
rect 7660 -14603 7672 -14569
rect 7706 -14603 7718 -14569
rect 7660 -14637 7718 -14603
rect 7660 -14671 7672 -14637
rect 7706 -14671 7718 -14637
rect 7660 -14705 7718 -14671
rect 7660 -14739 7672 -14705
rect 7706 -14739 7718 -14705
rect 7660 -14784 7718 -14739
rect 8678 -14229 8736 -14184
rect 8678 -14263 8690 -14229
rect 8724 -14263 8736 -14229
rect 8678 -14297 8736 -14263
rect 8678 -14331 8690 -14297
rect 8724 -14331 8736 -14297
rect 8678 -14365 8736 -14331
rect 8678 -14399 8690 -14365
rect 8724 -14399 8736 -14365
rect 8678 -14433 8736 -14399
rect 8678 -14467 8690 -14433
rect 8724 -14467 8736 -14433
rect 8678 -14501 8736 -14467
rect 8678 -14535 8690 -14501
rect 8724 -14535 8736 -14501
rect 8678 -14569 8736 -14535
rect 8678 -14603 8690 -14569
rect 8724 -14603 8736 -14569
rect 8678 -14637 8736 -14603
rect 8678 -14671 8690 -14637
rect 8724 -14671 8736 -14637
rect 8678 -14705 8736 -14671
rect 8678 -14739 8690 -14705
rect 8724 -14739 8736 -14705
rect 8678 -14784 8736 -14739
rect 9696 -14229 9754 -14184
rect 9696 -14263 9708 -14229
rect 9742 -14263 9754 -14229
rect 9696 -14297 9754 -14263
rect 9696 -14331 9708 -14297
rect 9742 -14331 9754 -14297
rect 9696 -14365 9754 -14331
rect 9696 -14399 9708 -14365
rect 9742 -14399 9754 -14365
rect 9696 -14433 9754 -14399
rect 9696 -14467 9708 -14433
rect 9742 -14467 9754 -14433
rect 9696 -14501 9754 -14467
rect 9696 -14535 9708 -14501
rect 9742 -14535 9754 -14501
rect 9696 -14569 9754 -14535
rect 9696 -14603 9708 -14569
rect 9742 -14603 9754 -14569
rect 9696 -14637 9754 -14603
rect 9696 -14671 9708 -14637
rect 9742 -14671 9754 -14637
rect 9696 -14705 9754 -14671
rect 9696 -14739 9708 -14705
rect 9742 -14739 9754 -14705
rect 9696 -14784 9754 -14739
rect 10714 -14229 10772 -14184
rect 10714 -14263 10726 -14229
rect 10760 -14263 10772 -14229
rect 10714 -14297 10772 -14263
rect 10714 -14331 10726 -14297
rect 10760 -14331 10772 -14297
rect 10714 -14365 10772 -14331
rect 10714 -14399 10726 -14365
rect 10760 -14399 10772 -14365
rect 10714 -14433 10772 -14399
rect 10714 -14467 10726 -14433
rect 10760 -14467 10772 -14433
rect 10714 -14501 10772 -14467
rect 10714 -14535 10726 -14501
rect 10760 -14535 10772 -14501
rect 10714 -14569 10772 -14535
rect 10714 -14603 10726 -14569
rect 10760 -14603 10772 -14569
rect 10714 -14637 10772 -14603
rect 10714 -14671 10726 -14637
rect 10760 -14671 10772 -14637
rect 10714 -14705 10772 -14671
rect 10714 -14739 10726 -14705
rect 10760 -14739 10772 -14705
rect 10714 -14784 10772 -14739
rect 11732 -14229 11790 -14184
rect 11732 -14263 11744 -14229
rect 11778 -14263 11790 -14229
rect 11732 -14297 11790 -14263
rect 11732 -14331 11744 -14297
rect 11778 -14331 11790 -14297
rect 11732 -14365 11790 -14331
rect 11732 -14399 11744 -14365
rect 11778 -14399 11790 -14365
rect 11732 -14433 11790 -14399
rect 11732 -14467 11744 -14433
rect 11778 -14467 11790 -14433
rect 11732 -14501 11790 -14467
rect 11732 -14535 11744 -14501
rect 11778 -14535 11790 -14501
rect 11732 -14569 11790 -14535
rect 11732 -14603 11744 -14569
rect 11778 -14603 11790 -14569
rect 11732 -14637 11790 -14603
rect 11732 -14671 11744 -14637
rect 11778 -14671 11790 -14637
rect 11732 -14705 11790 -14671
rect 11732 -14739 11744 -14705
rect 11778 -14739 11790 -14705
rect 11732 -14784 11790 -14739
rect 12750 -14229 12808 -14184
rect 12750 -14263 12762 -14229
rect 12796 -14263 12808 -14229
rect 12750 -14297 12808 -14263
rect 12750 -14331 12762 -14297
rect 12796 -14331 12808 -14297
rect 12750 -14365 12808 -14331
rect 12750 -14399 12762 -14365
rect 12796 -14399 12808 -14365
rect 12750 -14433 12808 -14399
rect 12750 -14467 12762 -14433
rect 12796 -14467 12808 -14433
rect 12750 -14501 12808 -14467
rect 12750 -14535 12762 -14501
rect 12796 -14535 12808 -14501
rect 12750 -14569 12808 -14535
rect 12750 -14603 12762 -14569
rect 12796 -14603 12808 -14569
rect 12750 -14637 12808 -14603
rect 12750 -14671 12762 -14637
rect 12796 -14671 12808 -14637
rect 12750 -14705 12808 -14671
rect 12750 -14739 12762 -14705
rect 12796 -14739 12808 -14705
rect 12750 -14784 12808 -14739
rect 13768 -14229 13826 -14184
rect 13768 -14263 13780 -14229
rect 13814 -14263 13826 -14229
rect 13768 -14297 13826 -14263
rect 13768 -14331 13780 -14297
rect 13814 -14331 13826 -14297
rect 13768 -14365 13826 -14331
rect 13768 -14399 13780 -14365
rect 13814 -14399 13826 -14365
rect 13768 -14433 13826 -14399
rect 13768 -14467 13780 -14433
rect 13814 -14467 13826 -14433
rect 13768 -14501 13826 -14467
rect 13768 -14535 13780 -14501
rect 13814 -14535 13826 -14501
rect 13768 -14569 13826 -14535
rect 13768 -14603 13780 -14569
rect 13814 -14603 13826 -14569
rect 13768 -14637 13826 -14603
rect 13768 -14671 13780 -14637
rect 13814 -14671 13826 -14637
rect 13768 -14705 13826 -14671
rect 13768 -14739 13780 -14705
rect 13814 -14739 13826 -14705
rect 13768 -14784 13826 -14739
rect 14786 -14229 14844 -14184
rect 14786 -14263 14798 -14229
rect 14832 -14263 14844 -14229
rect 14786 -14297 14844 -14263
rect 14786 -14331 14798 -14297
rect 14832 -14331 14844 -14297
rect 14786 -14365 14844 -14331
rect 14786 -14399 14798 -14365
rect 14832 -14399 14844 -14365
rect 14786 -14433 14844 -14399
rect 14786 -14467 14798 -14433
rect 14832 -14467 14844 -14433
rect 14786 -14501 14844 -14467
rect 14786 -14535 14798 -14501
rect 14832 -14535 14844 -14501
rect 14786 -14569 14844 -14535
rect 14786 -14603 14798 -14569
rect 14832 -14603 14844 -14569
rect 14786 -14637 14844 -14603
rect 14786 -14671 14798 -14637
rect 14832 -14671 14844 -14637
rect 14786 -14705 14844 -14671
rect 14786 -14739 14798 -14705
rect 14832 -14739 14844 -14705
rect 14786 -14784 14844 -14739
rect 15804 -14229 15862 -14184
rect 15804 -14263 15816 -14229
rect 15850 -14263 15862 -14229
rect 15804 -14297 15862 -14263
rect 15804 -14331 15816 -14297
rect 15850 -14331 15862 -14297
rect 15804 -14365 15862 -14331
rect 15804 -14399 15816 -14365
rect 15850 -14399 15862 -14365
rect 15804 -14433 15862 -14399
rect 15804 -14467 15816 -14433
rect 15850 -14467 15862 -14433
rect 15804 -14501 15862 -14467
rect 15804 -14535 15816 -14501
rect 15850 -14535 15862 -14501
rect 15804 -14569 15862 -14535
rect 15804 -14603 15816 -14569
rect 15850 -14603 15862 -14569
rect 15804 -14637 15862 -14603
rect 15804 -14671 15816 -14637
rect 15850 -14671 15862 -14637
rect 15804 -14705 15862 -14671
rect 15804 -14739 15816 -14705
rect 15850 -14739 15862 -14705
rect 15804 -14784 15862 -14739
rect 16822 -14229 16880 -14184
rect 16822 -14263 16834 -14229
rect 16868 -14263 16880 -14229
rect 16822 -14297 16880 -14263
rect 16822 -14331 16834 -14297
rect 16868 -14331 16880 -14297
rect 16822 -14365 16880 -14331
rect 16822 -14399 16834 -14365
rect 16868 -14399 16880 -14365
rect 16822 -14433 16880 -14399
rect 16822 -14467 16834 -14433
rect 16868 -14467 16880 -14433
rect 16822 -14501 16880 -14467
rect 16822 -14535 16834 -14501
rect 16868 -14535 16880 -14501
rect 16822 -14569 16880 -14535
rect 16822 -14603 16834 -14569
rect 16868 -14603 16880 -14569
rect 16822 -14637 16880 -14603
rect 16822 -14671 16834 -14637
rect 16868 -14671 16880 -14637
rect 16822 -14705 16880 -14671
rect 16822 -14739 16834 -14705
rect 16868 -14739 16880 -14705
rect 16822 -14784 16880 -14739
rect 17840 -14229 17898 -14184
rect 17840 -14263 17852 -14229
rect 17886 -14263 17898 -14229
rect 17840 -14297 17898 -14263
rect 17840 -14331 17852 -14297
rect 17886 -14331 17898 -14297
rect 17840 -14365 17898 -14331
rect 17840 -14399 17852 -14365
rect 17886 -14399 17898 -14365
rect 17840 -14433 17898 -14399
rect 17840 -14467 17852 -14433
rect 17886 -14467 17898 -14433
rect 17840 -14501 17898 -14467
rect 17840 -14535 17852 -14501
rect 17886 -14535 17898 -14501
rect 17840 -14569 17898 -14535
rect 17840 -14603 17852 -14569
rect 17886 -14603 17898 -14569
rect 17840 -14637 17898 -14603
rect 17840 -14671 17852 -14637
rect 17886 -14671 17898 -14637
rect 17840 -14705 17898 -14671
rect 17840 -14739 17852 -14705
rect 17886 -14739 17898 -14705
rect 17840 -14784 17898 -14739
rect 18858 -14229 18916 -14184
rect 18858 -14263 18870 -14229
rect 18904 -14263 18916 -14229
rect 18858 -14297 18916 -14263
rect 18858 -14331 18870 -14297
rect 18904 -14331 18916 -14297
rect 18858 -14365 18916 -14331
rect 18858 -14399 18870 -14365
rect 18904 -14399 18916 -14365
rect 18858 -14433 18916 -14399
rect 18858 -14467 18870 -14433
rect 18904 -14467 18916 -14433
rect 18858 -14501 18916 -14467
rect 18858 -14535 18870 -14501
rect 18904 -14535 18916 -14501
rect 18858 -14569 18916 -14535
rect 18858 -14603 18870 -14569
rect 18904 -14603 18916 -14569
rect 18858 -14637 18916 -14603
rect 18858 -14671 18870 -14637
rect 18904 -14671 18916 -14637
rect 18858 -14705 18916 -14671
rect 18858 -14739 18870 -14705
rect 18904 -14739 18916 -14705
rect 18858 -14784 18916 -14739
rect 19876 -14229 19934 -14184
rect 19876 -14263 19888 -14229
rect 19922 -14263 19934 -14229
rect 19876 -14297 19934 -14263
rect 19876 -14331 19888 -14297
rect 19922 -14331 19934 -14297
rect 19876 -14365 19934 -14331
rect 19876 -14399 19888 -14365
rect 19922 -14399 19934 -14365
rect 19876 -14433 19934 -14399
rect 19876 -14467 19888 -14433
rect 19922 -14467 19934 -14433
rect 19876 -14501 19934 -14467
rect 19876 -14535 19888 -14501
rect 19922 -14535 19934 -14501
rect 19876 -14569 19934 -14535
rect 19876 -14603 19888 -14569
rect 19922 -14603 19934 -14569
rect 19876 -14637 19934 -14603
rect 19876 -14671 19888 -14637
rect 19922 -14671 19934 -14637
rect 19876 -14705 19934 -14671
rect 19876 -14739 19888 -14705
rect 19922 -14739 19934 -14705
rect 19876 -14784 19934 -14739
rect 20894 -14229 20952 -14184
rect 20894 -14263 20906 -14229
rect 20940 -14263 20952 -14229
rect 20894 -14297 20952 -14263
rect 20894 -14331 20906 -14297
rect 20940 -14331 20952 -14297
rect 20894 -14365 20952 -14331
rect 20894 -14399 20906 -14365
rect 20940 -14399 20952 -14365
rect 20894 -14433 20952 -14399
rect 20894 -14467 20906 -14433
rect 20940 -14467 20952 -14433
rect 20894 -14501 20952 -14467
rect 20894 -14535 20906 -14501
rect 20940 -14535 20952 -14501
rect 20894 -14569 20952 -14535
rect 20894 -14603 20906 -14569
rect 20940 -14603 20952 -14569
rect 20894 -14637 20952 -14603
rect 20894 -14671 20906 -14637
rect 20940 -14671 20952 -14637
rect 20894 -14705 20952 -14671
rect 20894 -14739 20906 -14705
rect 20940 -14739 20952 -14705
rect 20894 -14784 20952 -14739
rect 21912 -14229 21970 -14184
rect 21912 -14263 21924 -14229
rect 21958 -14263 21970 -14229
rect 21912 -14297 21970 -14263
rect 21912 -14331 21924 -14297
rect 21958 -14331 21970 -14297
rect 21912 -14365 21970 -14331
rect 21912 -14399 21924 -14365
rect 21958 -14399 21970 -14365
rect 21912 -14433 21970 -14399
rect 21912 -14467 21924 -14433
rect 21958 -14467 21970 -14433
rect 21912 -14501 21970 -14467
rect 21912 -14535 21924 -14501
rect 21958 -14535 21970 -14501
rect 21912 -14569 21970 -14535
rect 21912 -14603 21924 -14569
rect 21958 -14603 21970 -14569
rect 21912 -14637 21970 -14603
rect 21912 -14671 21924 -14637
rect 21958 -14671 21970 -14637
rect 21912 -14705 21970 -14671
rect 21912 -14739 21924 -14705
rect 21958 -14739 21970 -14705
rect 21912 -14784 21970 -14739
rect 22930 -14229 22988 -14184
rect 22930 -14263 22942 -14229
rect 22976 -14263 22988 -14229
rect 22930 -14297 22988 -14263
rect 22930 -14331 22942 -14297
rect 22976 -14331 22988 -14297
rect 22930 -14365 22988 -14331
rect 22930 -14399 22942 -14365
rect 22976 -14399 22988 -14365
rect 22930 -14433 22988 -14399
rect 22930 -14467 22942 -14433
rect 22976 -14467 22988 -14433
rect 22930 -14501 22988 -14467
rect 22930 -14535 22942 -14501
rect 22976 -14535 22988 -14501
rect 22930 -14569 22988 -14535
rect 22930 -14603 22942 -14569
rect 22976 -14603 22988 -14569
rect 22930 -14637 22988 -14603
rect 22930 -14671 22942 -14637
rect 22976 -14671 22988 -14637
rect 22930 -14705 22988 -14671
rect 22930 -14739 22942 -14705
rect 22976 -14739 22988 -14705
rect 22930 -14784 22988 -14739
rect -9196 -15011 -9138 -14966
rect -9196 -15045 -9184 -15011
rect -9150 -15045 -9138 -15011
rect -9196 -15079 -9138 -15045
rect -9196 -15113 -9184 -15079
rect -9150 -15113 -9138 -15079
rect -9196 -15147 -9138 -15113
rect -9196 -15181 -9184 -15147
rect -9150 -15181 -9138 -15147
rect -9196 -15215 -9138 -15181
rect -9196 -15249 -9184 -15215
rect -9150 -15249 -9138 -15215
rect -9196 -15283 -9138 -15249
rect -9196 -15317 -9184 -15283
rect -9150 -15317 -9138 -15283
rect -9196 -15351 -9138 -15317
rect -9196 -15385 -9184 -15351
rect -9150 -15385 -9138 -15351
rect -9196 -15419 -9138 -15385
rect -9196 -15453 -9184 -15419
rect -9150 -15453 -9138 -15419
rect -9196 -15487 -9138 -15453
rect -9196 -15521 -9184 -15487
rect -9150 -15521 -9138 -15487
rect -9196 -15566 -9138 -15521
rect -8178 -15011 -8120 -14966
rect -8178 -15045 -8166 -15011
rect -8132 -15045 -8120 -15011
rect -8178 -15079 -8120 -15045
rect -8178 -15113 -8166 -15079
rect -8132 -15113 -8120 -15079
rect -8178 -15147 -8120 -15113
rect -8178 -15181 -8166 -15147
rect -8132 -15181 -8120 -15147
rect -8178 -15215 -8120 -15181
rect -8178 -15249 -8166 -15215
rect -8132 -15249 -8120 -15215
rect -8178 -15283 -8120 -15249
rect -8178 -15317 -8166 -15283
rect -8132 -15317 -8120 -15283
rect -8178 -15351 -8120 -15317
rect -8178 -15385 -8166 -15351
rect -8132 -15385 -8120 -15351
rect -8178 -15419 -8120 -15385
rect -8178 -15453 -8166 -15419
rect -8132 -15453 -8120 -15419
rect -8178 -15487 -8120 -15453
rect -8178 -15521 -8166 -15487
rect -8132 -15521 -8120 -15487
rect -8178 -15566 -8120 -15521
rect -7160 -15011 -7102 -14966
rect -7160 -15045 -7148 -15011
rect -7114 -15045 -7102 -15011
rect -7160 -15079 -7102 -15045
rect -7160 -15113 -7148 -15079
rect -7114 -15113 -7102 -15079
rect -7160 -15147 -7102 -15113
rect -7160 -15181 -7148 -15147
rect -7114 -15181 -7102 -15147
rect -7160 -15215 -7102 -15181
rect -7160 -15249 -7148 -15215
rect -7114 -15249 -7102 -15215
rect -7160 -15283 -7102 -15249
rect -7160 -15317 -7148 -15283
rect -7114 -15317 -7102 -15283
rect -7160 -15351 -7102 -15317
rect -7160 -15385 -7148 -15351
rect -7114 -15385 -7102 -15351
rect -7160 -15419 -7102 -15385
rect -7160 -15453 -7148 -15419
rect -7114 -15453 -7102 -15419
rect -7160 -15487 -7102 -15453
rect -7160 -15521 -7148 -15487
rect -7114 -15521 -7102 -15487
rect -7160 -15566 -7102 -15521
rect -6142 -15011 -6084 -14966
rect -6142 -15045 -6130 -15011
rect -6096 -15045 -6084 -15011
rect -6142 -15079 -6084 -15045
rect -6142 -15113 -6130 -15079
rect -6096 -15113 -6084 -15079
rect -6142 -15147 -6084 -15113
rect -6142 -15181 -6130 -15147
rect -6096 -15181 -6084 -15147
rect -6142 -15215 -6084 -15181
rect -6142 -15249 -6130 -15215
rect -6096 -15249 -6084 -15215
rect -6142 -15283 -6084 -15249
rect -6142 -15317 -6130 -15283
rect -6096 -15317 -6084 -15283
rect -6142 -15351 -6084 -15317
rect -6142 -15385 -6130 -15351
rect -6096 -15385 -6084 -15351
rect -6142 -15419 -6084 -15385
rect -6142 -15453 -6130 -15419
rect -6096 -15453 -6084 -15419
rect -6142 -15487 -6084 -15453
rect -6142 -15521 -6130 -15487
rect -6096 -15521 -6084 -15487
rect -6142 -15566 -6084 -15521
rect -5124 -15011 -5066 -14966
rect -5124 -15045 -5112 -15011
rect -5078 -15045 -5066 -15011
rect -5124 -15079 -5066 -15045
rect -5124 -15113 -5112 -15079
rect -5078 -15113 -5066 -15079
rect -5124 -15147 -5066 -15113
rect -5124 -15181 -5112 -15147
rect -5078 -15181 -5066 -15147
rect -5124 -15215 -5066 -15181
rect -5124 -15249 -5112 -15215
rect -5078 -15249 -5066 -15215
rect -5124 -15283 -5066 -15249
rect -5124 -15317 -5112 -15283
rect -5078 -15317 -5066 -15283
rect -5124 -15351 -5066 -15317
rect -5124 -15385 -5112 -15351
rect -5078 -15385 -5066 -15351
rect -5124 -15419 -5066 -15385
rect -5124 -15453 -5112 -15419
rect -5078 -15453 -5066 -15419
rect -5124 -15487 -5066 -15453
rect -5124 -15521 -5112 -15487
rect -5078 -15521 -5066 -15487
rect -5124 -15566 -5066 -15521
rect -4106 -15011 -4048 -14966
rect -4106 -15045 -4094 -15011
rect -4060 -15045 -4048 -15011
rect -4106 -15079 -4048 -15045
rect -4106 -15113 -4094 -15079
rect -4060 -15113 -4048 -15079
rect -4106 -15147 -4048 -15113
rect -4106 -15181 -4094 -15147
rect -4060 -15181 -4048 -15147
rect -4106 -15215 -4048 -15181
rect -4106 -15249 -4094 -15215
rect -4060 -15249 -4048 -15215
rect -4106 -15283 -4048 -15249
rect -4106 -15317 -4094 -15283
rect -4060 -15317 -4048 -15283
rect -4106 -15351 -4048 -15317
rect -4106 -15385 -4094 -15351
rect -4060 -15385 -4048 -15351
rect -4106 -15419 -4048 -15385
rect -4106 -15453 -4094 -15419
rect -4060 -15453 -4048 -15419
rect -4106 -15487 -4048 -15453
rect -4106 -15521 -4094 -15487
rect -4060 -15521 -4048 -15487
rect -4106 -15566 -4048 -15521
rect -3088 -15011 -3030 -14966
rect -3088 -15045 -3076 -15011
rect -3042 -15045 -3030 -15011
rect -3088 -15079 -3030 -15045
rect -3088 -15113 -3076 -15079
rect -3042 -15113 -3030 -15079
rect -3088 -15147 -3030 -15113
rect -3088 -15181 -3076 -15147
rect -3042 -15181 -3030 -15147
rect -3088 -15215 -3030 -15181
rect -3088 -15249 -3076 -15215
rect -3042 -15249 -3030 -15215
rect -3088 -15283 -3030 -15249
rect -3088 -15317 -3076 -15283
rect -3042 -15317 -3030 -15283
rect -3088 -15351 -3030 -15317
rect -3088 -15385 -3076 -15351
rect -3042 -15385 -3030 -15351
rect -3088 -15419 -3030 -15385
rect -3088 -15453 -3076 -15419
rect -3042 -15453 -3030 -15419
rect -3088 -15487 -3030 -15453
rect -3088 -15521 -3076 -15487
rect -3042 -15521 -3030 -15487
rect -3088 -15566 -3030 -15521
rect -2070 -15011 -2012 -14966
rect -2070 -15045 -2058 -15011
rect -2024 -15045 -2012 -15011
rect -2070 -15079 -2012 -15045
rect -2070 -15113 -2058 -15079
rect -2024 -15113 -2012 -15079
rect -2070 -15147 -2012 -15113
rect -2070 -15181 -2058 -15147
rect -2024 -15181 -2012 -15147
rect -2070 -15215 -2012 -15181
rect -2070 -15249 -2058 -15215
rect -2024 -15249 -2012 -15215
rect -2070 -15283 -2012 -15249
rect -2070 -15317 -2058 -15283
rect -2024 -15317 -2012 -15283
rect -2070 -15351 -2012 -15317
rect -2070 -15385 -2058 -15351
rect -2024 -15385 -2012 -15351
rect -2070 -15419 -2012 -15385
rect -2070 -15453 -2058 -15419
rect -2024 -15453 -2012 -15419
rect -2070 -15487 -2012 -15453
rect -2070 -15521 -2058 -15487
rect -2024 -15521 -2012 -15487
rect -2070 -15566 -2012 -15521
rect -1052 -15011 -994 -14966
rect -1052 -15045 -1040 -15011
rect -1006 -15045 -994 -15011
rect -1052 -15079 -994 -15045
rect -1052 -15113 -1040 -15079
rect -1006 -15113 -994 -15079
rect -1052 -15147 -994 -15113
rect -1052 -15181 -1040 -15147
rect -1006 -15181 -994 -15147
rect -1052 -15215 -994 -15181
rect -1052 -15249 -1040 -15215
rect -1006 -15249 -994 -15215
rect -1052 -15283 -994 -15249
rect -1052 -15317 -1040 -15283
rect -1006 -15317 -994 -15283
rect -1052 -15351 -994 -15317
rect -1052 -15385 -1040 -15351
rect -1006 -15385 -994 -15351
rect -1052 -15419 -994 -15385
rect -1052 -15453 -1040 -15419
rect -1006 -15453 -994 -15419
rect -1052 -15487 -994 -15453
rect -1052 -15521 -1040 -15487
rect -1006 -15521 -994 -15487
rect -1052 -15566 -994 -15521
rect -34 -15011 24 -14966
rect -34 -15045 -22 -15011
rect 12 -15045 24 -15011
rect -34 -15079 24 -15045
rect -34 -15113 -22 -15079
rect 12 -15113 24 -15079
rect -34 -15147 24 -15113
rect -34 -15181 -22 -15147
rect 12 -15181 24 -15147
rect -34 -15215 24 -15181
rect -34 -15249 -22 -15215
rect 12 -15249 24 -15215
rect -34 -15283 24 -15249
rect -34 -15317 -22 -15283
rect 12 -15317 24 -15283
rect -34 -15351 24 -15317
rect -34 -15385 -22 -15351
rect 12 -15385 24 -15351
rect -34 -15419 24 -15385
rect -34 -15453 -22 -15419
rect 12 -15453 24 -15419
rect -34 -15487 24 -15453
rect -34 -15521 -22 -15487
rect 12 -15521 24 -15487
rect -34 -15566 24 -15521
rect 2568 -15463 2626 -15418
rect 2568 -15497 2580 -15463
rect 2614 -15497 2626 -15463
rect 2568 -15531 2626 -15497
rect 2568 -15565 2580 -15531
rect 2614 -15565 2626 -15531
rect 2568 -15599 2626 -15565
rect 2568 -15633 2580 -15599
rect 2614 -15633 2626 -15599
rect 2568 -15667 2626 -15633
rect 2568 -15701 2580 -15667
rect 2614 -15701 2626 -15667
rect 2568 -15735 2626 -15701
rect 2568 -15769 2580 -15735
rect 2614 -15769 2626 -15735
rect -9196 -15829 -9138 -15784
rect -9196 -15863 -9184 -15829
rect -9150 -15863 -9138 -15829
rect -9196 -15897 -9138 -15863
rect -9196 -15931 -9184 -15897
rect -9150 -15931 -9138 -15897
rect -9196 -15965 -9138 -15931
rect -9196 -15999 -9184 -15965
rect -9150 -15999 -9138 -15965
rect -9196 -16033 -9138 -15999
rect -9196 -16067 -9184 -16033
rect -9150 -16067 -9138 -16033
rect -9196 -16101 -9138 -16067
rect -9196 -16135 -9184 -16101
rect -9150 -16135 -9138 -16101
rect -9196 -16169 -9138 -16135
rect -9196 -16203 -9184 -16169
rect -9150 -16203 -9138 -16169
rect -9196 -16237 -9138 -16203
rect -9196 -16271 -9184 -16237
rect -9150 -16271 -9138 -16237
rect -9196 -16305 -9138 -16271
rect -9196 -16339 -9184 -16305
rect -9150 -16339 -9138 -16305
rect -9196 -16384 -9138 -16339
rect -8178 -15829 -8120 -15784
rect -8178 -15863 -8166 -15829
rect -8132 -15863 -8120 -15829
rect -8178 -15897 -8120 -15863
rect -8178 -15931 -8166 -15897
rect -8132 -15931 -8120 -15897
rect -8178 -15965 -8120 -15931
rect -8178 -15999 -8166 -15965
rect -8132 -15999 -8120 -15965
rect -8178 -16033 -8120 -15999
rect -8178 -16067 -8166 -16033
rect -8132 -16067 -8120 -16033
rect -8178 -16101 -8120 -16067
rect -8178 -16135 -8166 -16101
rect -8132 -16135 -8120 -16101
rect -8178 -16169 -8120 -16135
rect -8178 -16203 -8166 -16169
rect -8132 -16203 -8120 -16169
rect -8178 -16237 -8120 -16203
rect -8178 -16271 -8166 -16237
rect -8132 -16271 -8120 -16237
rect -8178 -16305 -8120 -16271
rect -8178 -16339 -8166 -16305
rect -8132 -16339 -8120 -16305
rect -8178 -16384 -8120 -16339
rect -7160 -15829 -7102 -15784
rect -7160 -15863 -7148 -15829
rect -7114 -15863 -7102 -15829
rect -7160 -15897 -7102 -15863
rect -7160 -15931 -7148 -15897
rect -7114 -15931 -7102 -15897
rect -7160 -15965 -7102 -15931
rect -7160 -15999 -7148 -15965
rect -7114 -15999 -7102 -15965
rect -7160 -16033 -7102 -15999
rect -7160 -16067 -7148 -16033
rect -7114 -16067 -7102 -16033
rect -7160 -16101 -7102 -16067
rect -7160 -16135 -7148 -16101
rect -7114 -16135 -7102 -16101
rect -7160 -16169 -7102 -16135
rect -7160 -16203 -7148 -16169
rect -7114 -16203 -7102 -16169
rect -7160 -16237 -7102 -16203
rect -7160 -16271 -7148 -16237
rect -7114 -16271 -7102 -16237
rect -7160 -16305 -7102 -16271
rect -7160 -16339 -7148 -16305
rect -7114 -16339 -7102 -16305
rect -7160 -16384 -7102 -16339
rect -6142 -15829 -6084 -15784
rect -6142 -15863 -6130 -15829
rect -6096 -15863 -6084 -15829
rect -6142 -15897 -6084 -15863
rect -6142 -15931 -6130 -15897
rect -6096 -15931 -6084 -15897
rect -6142 -15965 -6084 -15931
rect -6142 -15999 -6130 -15965
rect -6096 -15999 -6084 -15965
rect -6142 -16033 -6084 -15999
rect -6142 -16067 -6130 -16033
rect -6096 -16067 -6084 -16033
rect -6142 -16101 -6084 -16067
rect -6142 -16135 -6130 -16101
rect -6096 -16135 -6084 -16101
rect -6142 -16169 -6084 -16135
rect -6142 -16203 -6130 -16169
rect -6096 -16203 -6084 -16169
rect -6142 -16237 -6084 -16203
rect -6142 -16271 -6130 -16237
rect -6096 -16271 -6084 -16237
rect -6142 -16305 -6084 -16271
rect -6142 -16339 -6130 -16305
rect -6096 -16339 -6084 -16305
rect -6142 -16384 -6084 -16339
rect -5124 -15829 -5066 -15784
rect -5124 -15863 -5112 -15829
rect -5078 -15863 -5066 -15829
rect -5124 -15897 -5066 -15863
rect -5124 -15931 -5112 -15897
rect -5078 -15931 -5066 -15897
rect -5124 -15965 -5066 -15931
rect -5124 -15999 -5112 -15965
rect -5078 -15999 -5066 -15965
rect -5124 -16033 -5066 -15999
rect -5124 -16067 -5112 -16033
rect -5078 -16067 -5066 -16033
rect -5124 -16101 -5066 -16067
rect -5124 -16135 -5112 -16101
rect -5078 -16135 -5066 -16101
rect -5124 -16169 -5066 -16135
rect -5124 -16203 -5112 -16169
rect -5078 -16203 -5066 -16169
rect -5124 -16237 -5066 -16203
rect -5124 -16271 -5112 -16237
rect -5078 -16271 -5066 -16237
rect -5124 -16305 -5066 -16271
rect -5124 -16339 -5112 -16305
rect -5078 -16339 -5066 -16305
rect -5124 -16384 -5066 -16339
rect -4106 -15829 -4048 -15784
rect -4106 -15863 -4094 -15829
rect -4060 -15863 -4048 -15829
rect -4106 -15897 -4048 -15863
rect -4106 -15931 -4094 -15897
rect -4060 -15931 -4048 -15897
rect -4106 -15965 -4048 -15931
rect -4106 -15999 -4094 -15965
rect -4060 -15999 -4048 -15965
rect -4106 -16033 -4048 -15999
rect -4106 -16067 -4094 -16033
rect -4060 -16067 -4048 -16033
rect -4106 -16101 -4048 -16067
rect -4106 -16135 -4094 -16101
rect -4060 -16135 -4048 -16101
rect -4106 -16169 -4048 -16135
rect -4106 -16203 -4094 -16169
rect -4060 -16203 -4048 -16169
rect -4106 -16237 -4048 -16203
rect -4106 -16271 -4094 -16237
rect -4060 -16271 -4048 -16237
rect -4106 -16305 -4048 -16271
rect -4106 -16339 -4094 -16305
rect -4060 -16339 -4048 -16305
rect -4106 -16384 -4048 -16339
rect -3088 -15829 -3030 -15784
rect -3088 -15863 -3076 -15829
rect -3042 -15863 -3030 -15829
rect -3088 -15897 -3030 -15863
rect -3088 -15931 -3076 -15897
rect -3042 -15931 -3030 -15897
rect -3088 -15965 -3030 -15931
rect -3088 -15999 -3076 -15965
rect -3042 -15999 -3030 -15965
rect -3088 -16033 -3030 -15999
rect -3088 -16067 -3076 -16033
rect -3042 -16067 -3030 -16033
rect -3088 -16101 -3030 -16067
rect -3088 -16135 -3076 -16101
rect -3042 -16135 -3030 -16101
rect -3088 -16169 -3030 -16135
rect -3088 -16203 -3076 -16169
rect -3042 -16203 -3030 -16169
rect -3088 -16237 -3030 -16203
rect -3088 -16271 -3076 -16237
rect -3042 -16271 -3030 -16237
rect -3088 -16305 -3030 -16271
rect -3088 -16339 -3076 -16305
rect -3042 -16339 -3030 -16305
rect -3088 -16384 -3030 -16339
rect -2070 -15829 -2012 -15784
rect -2070 -15863 -2058 -15829
rect -2024 -15863 -2012 -15829
rect -2070 -15897 -2012 -15863
rect -2070 -15931 -2058 -15897
rect -2024 -15931 -2012 -15897
rect -2070 -15965 -2012 -15931
rect -2070 -15999 -2058 -15965
rect -2024 -15999 -2012 -15965
rect -2070 -16033 -2012 -15999
rect -2070 -16067 -2058 -16033
rect -2024 -16067 -2012 -16033
rect -2070 -16101 -2012 -16067
rect -2070 -16135 -2058 -16101
rect -2024 -16135 -2012 -16101
rect -2070 -16169 -2012 -16135
rect -2070 -16203 -2058 -16169
rect -2024 -16203 -2012 -16169
rect -2070 -16237 -2012 -16203
rect -2070 -16271 -2058 -16237
rect -2024 -16271 -2012 -16237
rect -2070 -16305 -2012 -16271
rect -2070 -16339 -2058 -16305
rect -2024 -16339 -2012 -16305
rect -2070 -16384 -2012 -16339
rect -1052 -15829 -994 -15784
rect -1052 -15863 -1040 -15829
rect -1006 -15863 -994 -15829
rect -1052 -15897 -994 -15863
rect -1052 -15931 -1040 -15897
rect -1006 -15931 -994 -15897
rect -1052 -15965 -994 -15931
rect -1052 -15999 -1040 -15965
rect -1006 -15999 -994 -15965
rect -1052 -16033 -994 -15999
rect -1052 -16067 -1040 -16033
rect -1006 -16067 -994 -16033
rect -1052 -16101 -994 -16067
rect -1052 -16135 -1040 -16101
rect -1006 -16135 -994 -16101
rect -1052 -16169 -994 -16135
rect -1052 -16203 -1040 -16169
rect -1006 -16203 -994 -16169
rect -1052 -16237 -994 -16203
rect -1052 -16271 -1040 -16237
rect -1006 -16271 -994 -16237
rect -1052 -16305 -994 -16271
rect -1052 -16339 -1040 -16305
rect -1006 -16339 -994 -16305
rect -1052 -16384 -994 -16339
rect -34 -15829 24 -15784
rect -34 -15863 -22 -15829
rect 12 -15863 24 -15829
rect -34 -15897 24 -15863
rect -34 -15931 -22 -15897
rect 12 -15931 24 -15897
rect -34 -15965 24 -15931
rect -34 -15999 -22 -15965
rect 12 -15999 24 -15965
rect -34 -16033 24 -15999
rect 2568 -15803 2626 -15769
rect 2568 -15837 2580 -15803
rect 2614 -15837 2626 -15803
rect 2568 -15871 2626 -15837
rect 2568 -15905 2580 -15871
rect 2614 -15905 2626 -15871
rect 2568 -15939 2626 -15905
rect 2568 -15973 2580 -15939
rect 2614 -15973 2626 -15939
rect 2568 -16018 2626 -15973
rect 3586 -15463 3644 -15418
rect 3586 -15497 3598 -15463
rect 3632 -15497 3644 -15463
rect 3586 -15531 3644 -15497
rect 3586 -15565 3598 -15531
rect 3632 -15565 3644 -15531
rect 3586 -15599 3644 -15565
rect 3586 -15633 3598 -15599
rect 3632 -15633 3644 -15599
rect 3586 -15667 3644 -15633
rect 3586 -15701 3598 -15667
rect 3632 -15701 3644 -15667
rect 3586 -15735 3644 -15701
rect 3586 -15769 3598 -15735
rect 3632 -15769 3644 -15735
rect 3586 -15803 3644 -15769
rect 3586 -15837 3598 -15803
rect 3632 -15837 3644 -15803
rect 3586 -15871 3644 -15837
rect 3586 -15905 3598 -15871
rect 3632 -15905 3644 -15871
rect 3586 -15939 3644 -15905
rect 3586 -15973 3598 -15939
rect 3632 -15973 3644 -15939
rect 3586 -16018 3644 -15973
rect 4604 -15463 4662 -15418
rect 4604 -15497 4616 -15463
rect 4650 -15497 4662 -15463
rect 4604 -15531 4662 -15497
rect 4604 -15565 4616 -15531
rect 4650 -15565 4662 -15531
rect 4604 -15599 4662 -15565
rect 4604 -15633 4616 -15599
rect 4650 -15633 4662 -15599
rect 4604 -15667 4662 -15633
rect 4604 -15701 4616 -15667
rect 4650 -15701 4662 -15667
rect 4604 -15735 4662 -15701
rect 4604 -15769 4616 -15735
rect 4650 -15769 4662 -15735
rect 4604 -15803 4662 -15769
rect 4604 -15837 4616 -15803
rect 4650 -15837 4662 -15803
rect 4604 -15871 4662 -15837
rect 4604 -15905 4616 -15871
rect 4650 -15905 4662 -15871
rect 4604 -15939 4662 -15905
rect 4604 -15973 4616 -15939
rect 4650 -15973 4662 -15939
rect 4604 -16018 4662 -15973
rect 5622 -15463 5680 -15418
rect 5622 -15497 5634 -15463
rect 5668 -15497 5680 -15463
rect 5622 -15531 5680 -15497
rect 5622 -15565 5634 -15531
rect 5668 -15565 5680 -15531
rect 5622 -15599 5680 -15565
rect 5622 -15633 5634 -15599
rect 5668 -15633 5680 -15599
rect 5622 -15667 5680 -15633
rect 5622 -15701 5634 -15667
rect 5668 -15701 5680 -15667
rect 5622 -15735 5680 -15701
rect 5622 -15769 5634 -15735
rect 5668 -15769 5680 -15735
rect 5622 -15803 5680 -15769
rect 5622 -15837 5634 -15803
rect 5668 -15837 5680 -15803
rect 5622 -15871 5680 -15837
rect 5622 -15905 5634 -15871
rect 5668 -15905 5680 -15871
rect 5622 -15939 5680 -15905
rect 5622 -15973 5634 -15939
rect 5668 -15973 5680 -15939
rect 5622 -16018 5680 -15973
rect 6640 -15463 6698 -15418
rect 6640 -15497 6652 -15463
rect 6686 -15497 6698 -15463
rect 6640 -15531 6698 -15497
rect 6640 -15565 6652 -15531
rect 6686 -15565 6698 -15531
rect 6640 -15599 6698 -15565
rect 6640 -15633 6652 -15599
rect 6686 -15633 6698 -15599
rect 6640 -15667 6698 -15633
rect 6640 -15701 6652 -15667
rect 6686 -15701 6698 -15667
rect 6640 -15735 6698 -15701
rect 6640 -15769 6652 -15735
rect 6686 -15769 6698 -15735
rect 6640 -15803 6698 -15769
rect 6640 -15837 6652 -15803
rect 6686 -15837 6698 -15803
rect 6640 -15871 6698 -15837
rect 6640 -15905 6652 -15871
rect 6686 -15905 6698 -15871
rect 6640 -15939 6698 -15905
rect 6640 -15973 6652 -15939
rect 6686 -15973 6698 -15939
rect 6640 -16018 6698 -15973
rect 7658 -15463 7716 -15418
rect 7658 -15497 7670 -15463
rect 7704 -15497 7716 -15463
rect 7658 -15531 7716 -15497
rect 7658 -15565 7670 -15531
rect 7704 -15565 7716 -15531
rect 7658 -15599 7716 -15565
rect 7658 -15633 7670 -15599
rect 7704 -15633 7716 -15599
rect 7658 -15667 7716 -15633
rect 7658 -15701 7670 -15667
rect 7704 -15701 7716 -15667
rect 7658 -15735 7716 -15701
rect 7658 -15769 7670 -15735
rect 7704 -15769 7716 -15735
rect 7658 -15803 7716 -15769
rect 7658 -15837 7670 -15803
rect 7704 -15837 7716 -15803
rect 7658 -15871 7716 -15837
rect 7658 -15905 7670 -15871
rect 7704 -15905 7716 -15871
rect 7658 -15939 7716 -15905
rect 7658 -15973 7670 -15939
rect 7704 -15973 7716 -15939
rect 7658 -16018 7716 -15973
rect 8676 -15463 8734 -15418
rect 8676 -15497 8688 -15463
rect 8722 -15497 8734 -15463
rect 8676 -15531 8734 -15497
rect 8676 -15565 8688 -15531
rect 8722 -15565 8734 -15531
rect 8676 -15599 8734 -15565
rect 8676 -15633 8688 -15599
rect 8722 -15633 8734 -15599
rect 8676 -15667 8734 -15633
rect 8676 -15701 8688 -15667
rect 8722 -15701 8734 -15667
rect 8676 -15735 8734 -15701
rect 8676 -15769 8688 -15735
rect 8722 -15769 8734 -15735
rect 8676 -15803 8734 -15769
rect 8676 -15837 8688 -15803
rect 8722 -15837 8734 -15803
rect 8676 -15871 8734 -15837
rect 8676 -15905 8688 -15871
rect 8722 -15905 8734 -15871
rect 8676 -15939 8734 -15905
rect 8676 -15973 8688 -15939
rect 8722 -15973 8734 -15939
rect 8676 -16018 8734 -15973
rect 9694 -15463 9752 -15418
rect 9694 -15497 9706 -15463
rect 9740 -15497 9752 -15463
rect 9694 -15531 9752 -15497
rect 9694 -15565 9706 -15531
rect 9740 -15565 9752 -15531
rect 9694 -15599 9752 -15565
rect 9694 -15633 9706 -15599
rect 9740 -15633 9752 -15599
rect 9694 -15667 9752 -15633
rect 9694 -15701 9706 -15667
rect 9740 -15701 9752 -15667
rect 9694 -15735 9752 -15701
rect 9694 -15769 9706 -15735
rect 9740 -15769 9752 -15735
rect 9694 -15803 9752 -15769
rect 9694 -15837 9706 -15803
rect 9740 -15837 9752 -15803
rect 9694 -15871 9752 -15837
rect 9694 -15905 9706 -15871
rect 9740 -15905 9752 -15871
rect 9694 -15939 9752 -15905
rect 9694 -15973 9706 -15939
rect 9740 -15973 9752 -15939
rect 9694 -16018 9752 -15973
rect 10712 -15463 10770 -15418
rect 10712 -15497 10724 -15463
rect 10758 -15497 10770 -15463
rect 10712 -15531 10770 -15497
rect 10712 -15565 10724 -15531
rect 10758 -15565 10770 -15531
rect 10712 -15599 10770 -15565
rect 10712 -15633 10724 -15599
rect 10758 -15633 10770 -15599
rect 10712 -15667 10770 -15633
rect 10712 -15701 10724 -15667
rect 10758 -15701 10770 -15667
rect 10712 -15735 10770 -15701
rect 10712 -15769 10724 -15735
rect 10758 -15769 10770 -15735
rect 10712 -15803 10770 -15769
rect 10712 -15837 10724 -15803
rect 10758 -15837 10770 -15803
rect 10712 -15871 10770 -15837
rect 10712 -15905 10724 -15871
rect 10758 -15905 10770 -15871
rect 10712 -15939 10770 -15905
rect 10712 -15973 10724 -15939
rect 10758 -15973 10770 -15939
rect 10712 -16018 10770 -15973
rect 11730 -15463 11788 -15418
rect 11730 -15497 11742 -15463
rect 11776 -15497 11788 -15463
rect 11730 -15531 11788 -15497
rect 11730 -15565 11742 -15531
rect 11776 -15565 11788 -15531
rect 11730 -15599 11788 -15565
rect 11730 -15633 11742 -15599
rect 11776 -15633 11788 -15599
rect 11730 -15667 11788 -15633
rect 11730 -15701 11742 -15667
rect 11776 -15701 11788 -15667
rect 11730 -15735 11788 -15701
rect 11730 -15769 11742 -15735
rect 11776 -15769 11788 -15735
rect 11730 -15803 11788 -15769
rect 11730 -15837 11742 -15803
rect 11776 -15837 11788 -15803
rect 11730 -15871 11788 -15837
rect 11730 -15905 11742 -15871
rect 11776 -15905 11788 -15871
rect 11730 -15939 11788 -15905
rect 11730 -15973 11742 -15939
rect 11776 -15973 11788 -15939
rect 11730 -16018 11788 -15973
rect 12748 -15463 12806 -15418
rect 12748 -15497 12760 -15463
rect 12794 -15497 12806 -15463
rect 12748 -15531 12806 -15497
rect 12748 -15565 12760 -15531
rect 12794 -15565 12806 -15531
rect 12748 -15599 12806 -15565
rect 12748 -15633 12760 -15599
rect 12794 -15633 12806 -15599
rect 12748 -15667 12806 -15633
rect 12748 -15701 12760 -15667
rect 12794 -15701 12806 -15667
rect 12748 -15735 12806 -15701
rect 12748 -15769 12760 -15735
rect 12794 -15769 12806 -15735
rect 12748 -15803 12806 -15769
rect 12748 -15837 12760 -15803
rect 12794 -15837 12806 -15803
rect 12748 -15871 12806 -15837
rect 12748 -15905 12760 -15871
rect 12794 -15905 12806 -15871
rect 12748 -15939 12806 -15905
rect 12748 -15973 12760 -15939
rect 12794 -15973 12806 -15939
rect 12748 -16018 12806 -15973
rect 13766 -15463 13824 -15418
rect 13766 -15497 13778 -15463
rect 13812 -15497 13824 -15463
rect 13766 -15531 13824 -15497
rect 13766 -15565 13778 -15531
rect 13812 -15565 13824 -15531
rect 13766 -15599 13824 -15565
rect 13766 -15633 13778 -15599
rect 13812 -15633 13824 -15599
rect 13766 -15667 13824 -15633
rect 13766 -15701 13778 -15667
rect 13812 -15701 13824 -15667
rect 13766 -15735 13824 -15701
rect 13766 -15769 13778 -15735
rect 13812 -15769 13824 -15735
rect 13766 -15803 13824 -15769
rect 13766 -15837 13778 -15803
rect 13812 -15837 13824 -15803
rect 13766 -15871 13824 -15837
rect 13766 -15905 13778 -15871
rect 13812 -15905 13824 -15871
rect 13766 -15939 13824 -15905
rect 13766 -15973 13778 -15939
rect 13812 -15973 13824 -15939
rect 13766 -16018 13824 -15973
rect 14784 -15463 14842 -15418
rect 14784 -15497 14796 -15463
rect 14830 -15497 14842 -15463
rect 14784 -15531 14842 -15497
rect 14784 -15565 14796 -15531
rect 14830 -15565 14842 -15531
rect 14784 -15599 14842 -15565
rect 14784 -15633 14796 -15599
rect 14830 -15633 14842 -15599
rect 14784 -15667 14842 -15633
rect 14784 -15701 14796 -15667
rect 14830 -15701 14842 -15667
rect 14784 -15735 14842 -15701
rect 14784 -15769 14796 -15735
rect 14830 -15769 14842 -15735
rect 14784 -15803 14842 -15769
rect 14784 -15837 14796 -15803
rect 14830 -15837 14842 -15803
rect 14784 -15871 14842 -15837
rect 14784 -15905 14796 -15871
rect 14830 -15905 14842 -15871
rect 14784 -15939 14842 -15905
rect 14784 -15973 14796 -15939
rect 14830 -15973 14842 -15939
rect 14784 -16018 14842 -15973
rect 15802 -15463 15860 -15418
rect 15802 -15497 15814 -15463
rect 15848 -15497 15860 -15463
rect 15802 -15531 15860 -15497
rect 15802 -15565 15814 -15531
rect 15848 -15565 15860 -15531
rect 15802 -15599 15860 -15565
rect 15802 -15633 15814 -15599
rect 15848 -15633 15860 -15599
rect 15802 -15667 15860 -15633
rect 15802 -15701 15814 -15667
rect 15848 -15701 15860 -15667
rect 15802 -15735 15860 -15701
rect 15802 -15769 15814 -15735
rect 15848 -15769 15860 -15735
rect 15802 -15803 15860 -15769
rect 15802 -15837 15814 -15803
rect 15848 -15837 15860 -15803
rect 15802 -15871 15860 -15837
rect 15802 -15905 15814 -15871
rect 15848 -15905 15860 -15871
rect 15802 -15939 15860 -15905
rect 15802 -15973 15814 -15939
rect 15848 -15973 15860 -15939
rect 15802 -16018 15860 -15973
rect 16820 -15463 16878 -15418
rect 16820 -15497 16832 -15463
rect 16866 -15497 16878 -15463
rect 16820 -15531 16878 -15497
rect 16820 -15565 16832 -15531
rect 16866 -15565 16878 -15531
rect 16820 -15599 16878 -15565
rect 16820 -15633 16832 -15599
rect 16866 -15633 16878 -15599
rect 16820 -15667 16878 -15633
rect 16820 -15701 16832 -15667
rect 16866 -15701 16878 -15667
rect 16820 -15735 16878 -15701
rect 16820 -15769 16832 -15735
rect 16866 -15769 16878 -15735
rect 16820 -15803 16878 -15769
rect 16820 -15837 16832 -15803
rect 16866 -15837 16878 -15803
rect 16820 -15871 16878 -15837
rect 16820 -15905 16832 -15871
rect 16866 -15905 16878 -15871
rect 16820 -15939 16878 -15905
rect 16820 -15973 16832 -15939
rect 16866 -15973 16878 -15939
rect 16820 -16018 16878 -15973
rect 17838 -15463 17896 -15418
rect 17838 -15497 17850 -15463
rect 17884 -15497 17896 -15463
rect 17838 -15531 17896 -15497
rect 17838 -15565 17850 -15531
rect 17884 -15565 17896 -15531
rect 17838 -15599 17896 -15565
rect 17838 -15633 17850 -15599
rect 17884 -15633 17896 -15599
rect 17838 -15667 17896 -15633
rect 17838 -15701 17850 -15667
rect 17884 -15701 17896 -15667
rect 17838 -15735 17896 -15701
rect 17838 -15769 17850 -15735
rect 17884 -15769 17896 -15735
rect 17838 -15803 17896 -15769
rect 17838 -15837 17850 -15803
rect 17884 -15837 17896 -15803
rect 17838 -15871 17896 -15837
rect 17838 -15905 17850 -15871
rect 17884 -15905 17896 -15871
rect 17838 -15939 17896 -15905
rect 17838 -15973 17850 -15939
rect 17884 -15973 17896 -15939
rect 17838 -16018 17896 -15973
rect 18856 -15463 18914 -15418
rect 18856 -15497 18868 -15463
rect 18902 -15497 18914 -15463
rect 18856 -15531 18914 -15497
rect 18856 -15565 18868 -15531
rect 18902 -15565 18914 -15531
rect 18856 -15599 18914 -15565
rect 18856 -15633 18868 -15599
rect 18902 -15633 18914 -15599
rect 18856 -15667 18914 -15633
rect 18856 -15701 18868 -15667
rect 18902 -15701 18914 -15667
rect 18856 -15735 18914 -15701
rect 18856 -15769 18868 -15735
rect 18902 -15769 18914 -15735
rect 18856 -15803 18914 -15769
rect 18856 -15837 18868 -15803
rect 18902 -15837 18914 -15803
rect 18856 -15871 18914 -15837
rect 18856 -15905 18868 -15871
rect 18902 -15905 18914 -15871
rect 18856 -15939 18914 -15905
rect 18856 -15973 18868 -15939
rect 18902 -15973 18914 -15939
rect 18856 -16018 18914 -15973
rect 19874 -15463 19932 -15418
rect 19874 -15497 19886 -15463
rect 19920 -15497 19932 -15463
rect 19874 -15531 19932 -15497
rect 19874 -15565 19886 -15531
rect 19920 -15565 19932 -15531
rect 19874 -15599 19932 -15565
rect 19874 -15633 19886 -15599
rect 19920 -15633 19932 -15599
rect 19874 -15667 19932 -15633
rect 19874 -15701 19886 -15667
rect 19920 -15701 19932 -15667
rect 19874 -15735 19932 -15701
rect 19874 -15769 19886 -15735
rect 19920 -15769 19932 -15735
rect 19874 -15803 19932 -15769
rect 19874 -15837 19886 -15803
rect 19920 -15837 19932 -15803
rect 19874 -15871 19932 -15837
rect 19874 -15905 19886 -15871
rect 19920 -15905 19932 -15871
rect 19874 -15939 19932 -15905
rect 19874 -15973 19886 -15939
rect 19920 -15973 19932 -15939
rect 19874 -16018 19932 -15973
rect 20892 -15463 20950 -15418
rect 20892 -15497 20904 -15463
rect 20938 -15497 20950 -15463
rect 20892 -15531 20950 -15497
rect 20892 -15565 20904 -15531
rect 20938 -15565 20950 -15531
rect 20892 -15599 20950 -15565
rect 20892 -15633 20904 -15599
rect 20938 -15633 20950 -15599
rect 20892 -15667 20950 -15633
rect 20892 -15701 20904 -15667
rect 20938 -15701 20950 -15667
rect 20892 -15735 20950 -15701
rect 20892 -15769 20904 -15735
rect 20938 -15769 20950 -15735
rect 20892 -15803 20950 -15769
rect 20892 -15837 20904 -15803
rect 20938 -15837 20950 -15803
rect 20892 -15871 20950 -15837
rect 20892 -15905 20904 -15871
rect 20938 -15905 20950 -15871
rect 20892 -15939 20950 -15905
rect 20892 -15973 20904 -15939
rect 20938 -15973 20950 -15939
rect 20892 -16018 20950 -15973
rect 21910 -15463 21968 -15418
rect 21910 -15497 21922 -15463
rect 21956 -15497 21968 -15463
rect 21910 -15531 21968 -15497
rect 21910 -15565 21922 -15531
rect 21956 -15565 21968 -15531
rect 21910 -15599 21968 -15565
rect 21910 -15633 21922 -15599
rect 21956 -15633 21968 -15599
rect 21910 -15667 21968 -15633
rect 21910 -15701 21922 -15667
rect 21956 -15701 21968 -15667
rect 21910 -15735 21968 -15701
rect 21910 -15769 21922 -15735
rect 21956 -15769 21968 -15735
rect 21910 -15803 21968 -15769
rect 21910 -15837 21922 -15803
rect 21956 -15837 21968 -15803
rect 21910 -15871 21968 -15837
rect 21910 -15905 21922 -15871
rect 21956 -15905 21968 -15871
rect 21910 -15939 21968 -15905
rect 21910 -15973 21922 -15939
rect 21956 -15973 21968 -15939
rect 21910 -16018 21968 -15973
rect 22928 -15463 22986 -15418
rect 22928 -15497 22940 -15463
rect 22974 -15497 22986 -15463
rect 22928 -15531 22986 -15497
rect 22928 -15565 22940 -15531
rect 22974 -15565 22986 -15531
rect 22928 -15599 22986 -15565
rect 22928 -15633 22940 -15599
rect 22974 -15633 22986 -15599
rect 22928 -15667 22986 -15633
rect 22928 -15701 22940 -15667
rect 22974 -15701 22986 -15667
rect 22928 -15735 22986 -15701
rect 22928 -15769 22940 -15735
rect 22974 -15769 22986 -15735
rect 22928 -15803 22986 -15769
rect 22928 -15837 22940 -15803
rect 22974 -15837 22986 -15803
rect 22928 -15871 22986 -15837
rect 22928 -15905 22940 -15871
rect 22974 -15905 22986 -15871
rect 22928 -15939 22986 -15905
rect 22928 -15973 22940 -15939
rect 22974 -15973 22986 -15939
rect 22928 -16018 22986 -15973
rect -34 -16067 -22 -16033
rect 12 -16067 24 -16033
rect -34 -16101 24 -16067
rect -34 -16135 -22 -16101
rect 12 -16135 24 -16101
rect -34 -16169 24 -16135
rect -34 -16203 -22 -16169
rect 12 -16203 24 -16169
rect -34 -16237 24 -16203
rect -34 -16271 -22 -16237
rect 12 -16271 24 -16237
rect -34 -16305 24 -16271
rect -34 -16339 -22 -16305
rect 12 -16339 24 -16305
rect -34 -16384 24 -16339
rect -9196 -16647 -9138 -16602
rect -9196 -16681 -9184 -16647
rect -9150 -16681 -9138 -16647
rect -9196 -16715 -9138 -16681
rect -9196 -16749 -9184 -16715
rect -9150 -16749 -9138 -16715
rect -9196 -16783 -9138 -16749
rect -9196 -16817 -9184 -16783
rect -9150 -16817 -9138 -16783
rect -9196 -16851 -9138 -16817
rect -9196 -16885 -9184 -16851
rect -9150 -16885 -9138 -16851
rect -9196 -16919 -9138 -16885
rect -9196 -16953 -9184 -16919
rect -9150 -16953 -9138 -16919
rect -9196 -16987 -9138 -16953
rect -9196 -17021 -9184 -16987
rect -9150 -17021 -9138 -16987
rect -9196 -17055 -9138 -17021
rect -9196 -17089 -9184 -17055
rect -9150 -17089 -9138 -17055
rect -9196 -17123 -9138 -17089
rect -9196 -17157 -9184 -17123
rect -9150 -17157 -9138 -17123
rect -9196 -17202 -9138 -17157
rect -8178 -16647 -8120 -16602
rect -8178 -16681 -8166 -16647
rect -8132 -16681 -8120 -16647
rect -8178 -16715 -8120 -16681
rect -8178 -16749 -8166 -16715
rect -8132 -16749 -8120 -16715
rect -8178 -16783 -8120 -16749
rect -8178 -16817 -8166 -16783
rect -8132 -16817 -8120 -16783
rect -8178 -16851 -8120 -16817
rect -8178 -16885 -8166 -16851
rect -8132 -16885 -8120 -16851
rect -8178 -16919 -8120 -16885
rect -8178 -16953 -8166 -16919
rect -8132 -16953 -8120 -16919
rect -8178 -16987 -8120 -16953
rect -8178 -17021 -8166 -16987
rect -8132 -17021 -8120 -16987
rect -8178 -17055 -8120 -17021
rect -8178 -17089 -8166 -17055
rect -8132 -17089 -8120 -17055
rect -8178 -17123 -8120 -17089
rect -8178 -17157 -8166 -17123
rect -8132 -17157 -8120 -17123
rect -8178 -17202 -8120 -17157
rect -7160 -16647 -7102 -16602
rect -7160 -16681 -7148 -16647
rect -7114 -16681 -7102 -16647
rect -7160 -16715 -7102 -16681
rect -7160 -16749 -7148 -16715
rect -7114 -16749 -7102 -16715
rect -7160 -16783 -7102 -16749
rect -7160 -16817 -7148 -16783
rect -7114 -16817 -7102 -16783
rect -7160 -16851 -7102 -16817
rect -7160 -16885 -7148 -16851
rect -7114 -16885 -7102 -16851
rect -7160 -16919 -7102 -16885
rect -7160 -16953 -7148 -16919
rect -7114 -16953 -7102 -16919
rect -7160 -16987 -7102 -16953
rect -7160 -17021 -7148 -16987
rect -7114 -17021 -7102 -16987
rect -7160 -17055 -7102 -17021
rect -7160 -17089 -7148 -17055
rect -7114 -17089 -7102 -17055
rect -7160 -17123 -7102 -17089
rect -7160 -17157 -7148 -17123
rect -7114 -17157 -7102 -17123
rect -7160 -17202 -7102 -17157
rect -6142 -16647 -6084 -16602
rect -6142 -16681 -6130 -16647
rect -6096 -16681 -6084 -16647
rect -6142 -16715 -6084 -16681
rect -6142 -16749 -6130 -16715
rect -6096 -16749 -6084 -16715
rect -6142 -16783 -6084 -16749
rect -6142 -16817 -6130 -16783
rect -6096 -16817 -6084 -16783
rect -6142 -16851 -6084 -16817
rect -6142 -16885 -6130 -16851
rect -6096 -16885 -6084 -16851
rect -6142 -16919 -6084 -16885
rect -6142 -16953 -6130 -16919
rect -6096 -16953 -6084 -16919
rect -6142 -16987 -6084 -16953
rect -6142 -17021 -6130 -16987
rect -6096 -17021 -6084 -16987
rect -6142 -17055 -6084 -17021
rect -6142 -17089 -6130 -17055
rect -6096 -17089 -6084 -17055
rect -6142 -17123 -6084 -17089
rect -6142 -17157 -6130 -17123
rect -6096 -17157 -6084 -17123
rect -6142 -17202 -6084 -17157
rect -5124 -16647 -5066 -16602
rect -5124 -16681 -5112 -16647
rect -5078 -16681 -5066 -16647
rect -5124 -16715 -5066 -16681
rect -5124 -16749 -5112 -16715
rect -5078 -16749 -5066 -16715
rect -5124 -16783 -5066 -16749
rect -5124 -16817 -5112 -16783
rect -5078 -16817 -5066 -16783
rect -5124 -16851 -5066 -16817
rect -5124 -16885 -5112 -16851
rect -5078 -16885 -5066 -16851
rect -5124 -16919 -5066 -16885
rect -5124 -16953 -5112 -16919
rect -5078 -16953 -5066 -16919
rect -5124 -16987 -5066 -16953
rect -5124 -17021 -5112 -16987
rect -5078 -17021 -5066 -16987
rect -5124 -17055 -5066 -17021
rect -5124 -17089 -5112 -17055
rect -5078 -17089 -5066 -17055
rect -5124 -17123 -5066 -17089
rect -5124 -17157 -5112 -17123
rect -5078 -17157 -5066 -17123
rect -5124 -17202 -5066 -17157
rect -4106 -16647 -4048 -16602
rect -4106 -16681 -4094 -16647
rect -4060 -16681 -4048 -16647
rect -4106 -16715 -4048 -16681
rect -4106 -16749 -4094 -16715
rect -4060 -16749 -4048 -16715
rect -4106 -16783 -4048 -16749
rect -4106 -16817 -4094 -16783
rect -4060 -16817 -4048 -16783
rect -4106 -16851 -4048 -16817
rect -4106 -16885 -4094 -16851
rect -4060 -16885 -4048 -16851
rect -4106 -16919 -4048 -16885
rect -4106 -16953 -4094 -16919
rect -4060 -16953 -4048 -16919
rect -4106 -16987 -4048 -16953
rect -4106 -17021 -4094 -16987
rect -4060 -17021 -4048 -16987
rect -4106 -17055 -4048 -17021
rect -4106 -17089 -4094 -17055
rect -4060 -17089 -4048 -17055
rect -4106 -17123 -4048 -17089
rect -4106 -17157 -4094 -17123
rect -4060 -17157 -4048 -17123
rect -4106 -17202 -4048 -17157
rect -3088 -16647 -3030 -16602
rect -3088 -16681 -3076 -16647
rect -3042 -16681 -3030 -16647
rect -3088 -16715 -3030 -16681
rect -3088 -16749 -3076 -16715
rect -3042 -16749 -3030 -16715
rect -3088 -16783 -3030 -16749
rect -3088 -16817 -3076 -16783
rect -3042 -16817 -3030 -16783
rect -3088 -16851 -3030 -16817
rect -3088 -16885 -3076 -16851
rect -3042 -16885 -3030 -16851
rect -3088 -16919 -3030 -16885
rect -3088 -16953 -3076 -16919
rect -3042 -16953 -3030 -16919
rect -3088 -16987 -3030 -16953
rect -3088 -17021 -3076 -16987
rect -3042 -17021 -3030 -16987
rect -3088 -17055 -3030 -17021
rect -3088 -17089 -3076 -17055
rect -3042 -17089 -3030 -17055
rect -3088 -17123 -3030 -17089
rect -3088 -17157 -3076 -17123
rect -3042 -17157 -3030 -17123
rect -3088 -17202 -3030 -17157
rect -2070 -16647 -2012 -16602
rect -2070 -16681 -2058 -16647
rect -2024 -16681 -2012 -16647
rect -2070 -16715 -2012 -16681
rect -2070 -16749 -2058 -16715
rect -2024 -16749 -2012 -16715
rect -2070 -16783 -2012 -16749
rect -2070 -16817 -2058 -16783
rect -2024 -16817 -2012 -16783
rect -2070 -16851 -2012 -16817
rect -2070 -16885 -2058 -16851
rect -2024 -16885 -2012 -16851
rect -2070 -16919 -2012 -16885
rect -2070 -16953 -2058 -16919
rect -2024 -16953 -2012 -16919
rect -2070 -16987 -2012 -16953
rect -2070 -17021 -2058 -16987
rect -2024 -17021 -2012 -16987
rect -2070 -17055 -2012 -17021
rect -2070 -17089 -2058 -17055
rect -2024 -17089 -2012 -17055
rect -2070 -17123 -2012 -17089
rect -2070 -17157 -2058 -17123
rect -2024 -17157 -2012 -17123
rect -2070 -17202 -2012 -17157
rect -1052 -16647 -994 -16602
rect -1052 -16681 -1040 -16647
rect -1006 -16681 -994 -16647
rect -1052 -16715 -994 -16681
rect -1052 -16749 -1040 -16715
rect -1006 -16749 -994 -16715
rect -1052 -16783 -994 -16749
rect -1052 -16817 -1040 -16783
rect -1006 -16817 -994 -16783
rect -1052 -16851 -994 -16817
rect -1052 -16885 -1040 -16851
rect -1006 -16885 -994 -16851
rect -1052 -16919 -994 -16885
rect -1052 -16953 -1040 -16919
rect -1006 -16953 -994 -16919
rect -1052 -16987 -994 -16953
rect -1052 -17021 -1040 -16987
rect -1006 -17021 -994 -16987
rect -1052 -17055 -994 -17021
rect -1052 -17089 -1040 -17055
rect -1006 -17089 -994 -17055
rect -1052 -17123 -994 -17089
rect -1052 -17157 -1040 -17123
rect -1006 -17157 -994 -17123
rect -1052 -17202 -994 -17157
rect -34 -16647 24 -16602
rect -34 -16681 -22 -16647
rect 12 -16681 24 -16647
rect -34 -16715 24 -16681
rect -34 -16749 -22 -16715
rect 12 -16749 24 -16715
rect -34 -16783 24 -16749
rect -34 -16817 -22 -16783
rect 12 -16817 24 -16783
rect -34 -16851 24 -16817
rect -34 -16885 -22 -16851
rect 12 -16885 24 -16851
rect -34 -16919 24 -16885
rect -34 -16953 -22 -16919
rect 12 -16953 24 -16919
rect -34 -16987 24 -16953
rect -34 -17021 -22 -16987
rect 12 -17021 24 -16987
rect -34 -17055 24 -17021
rect -34 -17089 -22 -17055
rect 12 -17089 24 -17055
rect -34 -17123 24 -17089
rect -34 -17157 -22 -17123
rect 12 -17157 24 -17123
rect -34 -17202 24 -17157
rect 2568 -16697 2626 -16652
rect 2568 -16731 2580 -16697
rect 2614 -16731 2626 -16697
rect 2568 -16765 2626 -16731
rect 2568 -16799 2580 -16765
rect 2614 -16799 2626 -16765
rect 2568 -16833 2626 -16799
rect 2568 -16867 2580 -16833
rect 2614 -16867 2626 -16833
rect 2568 -16901 2626 -16867
rect 2568 -16935 2580 -16901
rect 2614 -16935 2626 -16901
rect 2568 -16969 2626 -16935
rect 2568 -17003 2580 -16969
rect 2614 -17003 2626 -16969
rect 2568 -17037 2626 -17003
rect 2568 -17071 2580 -17037
rect 2614 -17071 2626 -17037
rect 2568 -17105 2626 -17071
rect 2568 -17139 2580 -17105
rect 2614 -17139 2626 -17105
rect 2568 -17173 2626 -17139
rect 2568 -17207 2580 -17173
rect 2614 -17207 2626 -17173
rect 2568 -17252 2626 -17207
rect 3586 -16697 3644 -16652
rect 3586 -16731 3598 -16697
rect 3632 -16731 3644 -16697
rect 3586 -16765 3644 -16731
rect 3586 -16799 3598 -16765
rect 3632 -16799 3644 -16765
rect 3586 -16833 3644 -16799
rect 3586 -16867 3598 -16833
rect 3632 -16867 3644 -16833
rect 3586 -16901 3644 -16867
rect 3586 -16935 3598 -16901
rect 3632 -16935 3644 -16901
rect 3586 -16969 3644 -16935
rect 3586 -17003 3598 -16969
rect 3632 -17003 3644 -16969
rect 3586 -17037 3644 -17003
rect 3586 -17071 3598 -17037
rect 3632 -17071 3644 -17037
rect 3586 -17105 3644 -17071
rect 3586 -17139 3598 -17105
rect 3632 -17139 3644 -17105
rect 3586 -17173 3644 -17139
rect 3586 -17207 3598 -17173
rect 3632 -17207 3644 -17173
rect 3586 -17252 3644 -17207
rect 4604 -16697 4662 -16652
rect 4604 -16731 4616 -16697
rect 4650 -16731 4662 -16697
rect 4604 -16765 4662 -16731
rect 4604 -16799 4616 -16765
rect 4650 -16799 4662 -16765
rect 4604 -16833 4662 -16799
rect 4604 -16867 4616 -16833
rect 4650 -16867 4662 -16833
rect 4604 -16901 4662 -16867
rect 4604 -16935 4616 -16901
rect 4650 -16935 4662 -16901
rect 4604 -16969 4662 -16935
rect 4604 -17003 4616 -16969
rect 4650 -17003 4662 -16969
rect 4604 -17037 4662 -17003
rect 4604 -17071 4616 -17037
rect 4650 -17071 4662 -17037
rect 4604 -17105 4662 -17071
rect 4604 -17139 4616 -17105
rect 4650 -17139 4662 -17105
rect 4604 -17173 4662 -17139
rect 4604 -17207 4616 -17173
rect 4650 -17207 4662 -17173
rect 4604 -17252 4662 -17207
rect 5622 -16697 5680 -16652
rect 5622 -16731 5634 -16697
rect 5668 -16731 5680 -16697
rect 5622 -16765 5680 -16731
rect 5622 -16799 5634 -16765
rect 5668 -16799 5680 -16765
rect 5622 -16833 5680 -16799
rect 5622 -16867 5634 -16833
rect 5668 -16867 5680 -16833
rect 5622 -16901 5680 -16867
rect 5622 -16935 5634 -16901
rect 5668 -16935 5680 -16901
rect 5622 -16969 5680 -16935
rect 5622 -17003 5634 -16969
rect 5668 -17003 5680 -16969
rect 5622 -17037 5680 -17003
rect 5622 -17071 5634 -17037
rect 5668 -17071 5680 -17037
rect 5622 -17105 5680 -17071
rect 5622 -17139 5634 -17105
rect 5668 -17139 5680 -17105
rect 5622 -17173 5680 -17139
rect 5622 -17207 5634 -17173
rect 5668 -17207 5680 -17173
rect 5622 -17252 5680 -17207
rect 6640 -16697 6698 -16652
rect 6640 -16731 6652 -16697
rect 6686 -16731 6698 -16697
rect 6640 -16765 6698 -16731
rect 6640 -16799 6652 -16765
rect 6686 -16799 6698 -16765
rect 6640 -16833 6698 -16799
rect 6640 -16867 6652 -16833
rect 6686 -16867 6698 -16833
rect 6640 -16901 6698 -16867
rect 6640 -16935 6652 -16901
rect 6686 -16935 6698 -16901
rect 6640 -16969 6698 -16935
rect 6640 -17003 6652 -16969
rect 6686 -17003 6698 -16969
rect 6640 -17037 6698 -17003
rect 6640 -17071 6652 -17037
rect 6686 -17071 6698 -17037
rect 6640 -17105 6698 -17071
rect 6640 -17139 6652 -17105
rect 6686 -17139 6698 -17105
rect 6640 -17173 6698 -17139
rect 6640 -17207 6652 -17173
rect 6686 -17207 6698 -17173
rect 6640 -17252 6698 -17207
rect 7658 -16697 7716 -16652
rect 7658 -16731 7670 -16697
rect 7704 -16731 7716 -16697
rect 7658 -16765 7716 -16731
rect 7658 -16799 7670 -16765
rect 7704 -16799 7716 -16765
rect 7658 -16833 7716 -16799
rect 7658 -16867 7670 -16833
rect 7704 -16867 7716 -16833
rect 7658 -16901 7716 -16867
rect 7658 -16935 7670 -16901
rect 7704 -16935 7716 -16901
rect 7658 -16969 7716 -16935
rect 7658 -17003 7670 -16969
rect 7704 -17003 7716 -16969
rect 7658 -17037 7716 -17003
rect 7658 -17071 7670 -17037
rect 7704 -17071 7716 -17037
rect 7658 -17105 7716 -17071
rect 7658 -17139 7670 -17105
rect 7704 -17139 7716 -17105
rect 7658 -17173 7716 -17139
rect 7658 -17207 7670 -17173
rect 7704 -17207 7716 -17173
rect 7658 -17252 7716 -17207
rect 8676 -16697 8734 -16652
rect 8676 -16731 8688 -16697
rect 8722 -16731 8734 -16697
rect 8676 -16765 8734 -16731
rect 8676 -16799 8688 -16765
rect 8722 -16799 8734 -16765
rect 8676 -16833 8734 -16799
rect 8676 -16867 8688 -16833
rect 8722 -16867 8734 -16833
rect 8676 -16901 8734 -16867
rect 8676 -16935 8688 -16901
rect 8722 -16935 8734 -16901
rect 8676 -16969 8734 -16935
rect 8676 -17003 8688 -16969
rect 8722 -17003 8734 -16969
rect 8676 -17037 8734 -17003
rect 8676 -17071 8688 -17037
rect 8722 -17071 8734 -17037
rect 8676 -17105 8734 -17071
rect 8676 -17139 8688 -17105
rect 8722 -17139 8734 -17105
rect 8676 -17173 8734 -17139
rect 8676 -17207 8688 -17173
rect 8722 -17207 8734 -17173
rect 8676 -17252 8734 -17207
rect 9694 -16697 9752 -16652
rect 9694 -16731 9706 -16697
rect 9740 -16731 9752 -16697
rect 9694 -16765 9752 -16731
rect 9694 -16799 9706 -16765
rect 9740 -16799 9752 -16765
rect 9694 -16833 9752 -16799
rect 9694 -16867 9706 -16833
rect 9740 -16867 9752 -16833
rect 9694 -16901 9752 -16867
rect 9694 -16935 9706 -16901
rect 9740 -16935 9752 -16901
rect 9694 -16969 9752 -16935
rect 9694 -17003 9706 -16969
rect 9740 -17003 9752 -16969
rect 9694 -17037 9752 -17003
rect 9694 -17071 9706 -17037
rect 9740 -17071 9752 -17037
rect 9694 -17105 9752 -17071
rect 9694 -17139 9706 -17105
rect 9740 -17139 9752 -17105
rect 9694 -17173 9752 -17139
rect 9694 -17207 9706 -17173
rect 9740 -17207 9752 -17173
rect 9694 -17252 9752 -17207
rect 10712 -16697 10770 -16652
rect 10712 -16731 10724 -16697
rect 10758 -16731 10770 -16697
rect 10712 -16765 10770 -16731
rect 10712 -16799 10724 -16765
rect 10758 -16799 10770 -16765
rect 10712 -16833 10770 -16799
rect 10712 -16867 10724 -16833
rect 10758 -16867 10770 -16833
rect 10712 -16901 10770 -16867
rect 10712 -16935 10724 -16901
rect 10758 -16935 10770 -16901
rect 10712 -16969 10770 -16935
rect 10712 -17003 10724 -16969
rect 10758 -17003 10770 -16969
rect 10712 -17037 10770 -17003
rect 10712 -17071 10724 -17037
rect 10758 -17071 10770 -17037
rect 10712 -17105 10770 -17071
rect 10712 -17139 10724 -17105
rect 10758 -17139 10770 -17105
rect 10712 -17173 10770 -17139
rect 10712 -17207 10724 -17173
rect 10758 -17207 10770 -17173
rect 10712 -17252 10770 -17207
rect 11730 -16697 11788 -16652
rect 11730 -16731 11742 -16697
rect 11776 -16731 11788 -16697
rect 11730 -16765 11788 -16731
rect 11730 -16799 11742 -16765
rect 11776 -16799 11788 -16765
rect 11730 -16833 11788 -16799
rect 11730 -16867 11742 -16833
rect 11776 -16867 11788 -16833
rect 11730 -16901 11788 -16867
rect 11730 -16935 11742 -16901
rect 11776 -16935 11788 -16901
rect 11730 -16969 11788 -16935
rect 11730 -17003 11742 -16969
rect 11776 -17003 11788 -16969
rect 11730 -17037 11788 -17003
rect 11730 -17071 11742 -17037
rect 11776 -17071 11788 -17037
rect 11730 -17105 11788 -17071
rect 11730 -17139 11742 -17105
rect 11776 -17139 11788 -17105
rect 11730 -17173 11788 -17139
rect 11730 -17207 11742 -17173
rect 11776 -17207 11788 -17173
rect 11730 -17252 11788 -17207
rect 12748 -16697 12806 -16652
rect 12748 -16731 12760 -16697
rect 12794 -16731 12806 -16697
rect 12748 -16765 12806 -16731
rect 12748 -16799 12760 -16765
rect 12794 -16799 12806 -16765
rect 12748 -16833 12806 -16799
rect 12748 -16867 12760 -16833
rect 12794 -16867 12806 -16833
rect 12748 -16901 12806 -16867
rect 12748 -16935 12760 -16901
rect 12794 -16935 12806 -16901
rect 12748 -16969 12806 -16935
rect 12748 -17003 12760 -16969
rect 12794 -17003 12806 -16969
rect 12748 -17037 12806 -17003
rect 12748 -17071 12760 -17037
rect 12794 -17071 12806 -17037
rect 12748 -17105 12806 -17071
rect 12748 -17139 12760 -17105
rect 12794 -17139 12806 -17105
rect 12748 -17173 12806 -17139
rect 12748 -17207 12760 -17173
rect 12794 -17207 12806 -17173
rect 12748 -17252 12806 -17207
rect 13766 -16697 13824 -16652
rect 13766 -16731 13778 -16697
rect 13812 -16731 13824 -16697
rect 13766 -16765 13824 -16731
rect 13766 -16799 13778 -16765
rect 13812 -16799 13824 -16765
rect 13766 -16833 13824 -16799
rect 13766 -16867 13778 -16833
rect 13812 -16867 13824 -16833
rect 13766 -16901 13824 -16867
rect 13766 -16935 13778 -16901
rect 13812 -16935 13824 -16901
rect 13766 -16969 13824 -16935
rect 13766 -17003 13778 -16969
rect 13812 -17003 13824 -16969
rect 13766 -17037 13824 -17003
rect 13766 -17071 13778 -17037
rect 13812 -17071 13824 -17037
rect 13766 -17105 13824 -17071
rect 13766 -17139 13778 -17105
rect 13812 -17139 13824 -17105
rect 13766 -17173 13824 -17139
rect 13766 -17207 13778 -17173
rect 13812 -17207 13824 -17173
rect 13766 -17252 13824 -17207
rect 14784 -16697 14842 -16652
rect 14784 -16731 14796 -16697
rect 14830 -16731 14842 -16697
rect 14784 -16765 14842 -16731
rect 14784 -16799 14796 -16765
rect 14830 -16799 14842 -16765
rect 14784 -16833 14842 -16799
rect 14784 -16867 14796 -16833
rect 14830 -16867 14842 -16833
rect 14784 -16901 14842 -16867
rect 14784 -16935 14796 -16901
rect 14830 -16935 14842 -16901
rect 14784 -16969 14842 -16935
rect 14784 -17003 14796 -16969
rect 14830 -17003 14842 -16969
rect 14784 -17037 14842 -17003
rect 14784 -17071 14796 -17037
rect 14830 -17071 14842 -17037
rect 14784 -17105 14842 -17071
rect 14784 -17139 14796 -17105
rect 14830 -17139 14842 -17105
rect 14784 -17173 14842 -17139
rect 14784 -17207 14796 -17173
rect 14830 -17207 14842 -17173
rect 14784 -17252 14842 -17207
rect 15802 -16697 15860 -16652
rect 15802 -16731 15814 -16697
rect 15848 -16731 15860 -16697
rect 15802 -16765 15860 -16731
rect 15802 -16799 15814 -16765
rect 15848 -16799 15860 -16765
rect 15802 -16833 15860 -16799
rect 15802 -16867 15814 -16833
rect 15848 -16867 15860 -16833
rect 15802 -16901 15860 -16867
rect 15802 -16935 15814 -16901
rect 15848 -16935 15860 -16901
rect 15802 -16969 15860 -16935
rect 15802 -17003 15814 -16969
rect 15848 -17003 15860 -16969
rect 15802 -17037 15860 -17003
rect 15802 -17071 15814 -17037
rect 15848 -17071 15860 -17037
rect 15802 -17105 15860 -17071
rect 15802 -17139 15814 -17105
rect 15848 -17139 15860 -17105
rect 15802 -17173 15860 -17139
rect 15802 -17207 15814 -17173
rect 15848 -17207 15860 -17173
rect 15802 -17252 15860 -17207
rect 16820 -16697 16878 -16652
rect 16820 -16731 16832 -16697
rect 16866 -16731 16878 -16697
rect 16820 -16765 16878 -16731
rect 16820 -16799 16832 -16765
rect 16866 -16799 16878 -16765
rect 16820 -16833 16878 -16799
rect 16820 -16867 16832 -16833
rect 16866 -16867 16878 -16833
rect 16820 -16901 16878 -16867
rect 16820 -16935 16832 -16901
rect 16866 -16935 16878 -16901
rect 16820 -16969 16878 -16935
rect 16820 -17003 16832 -16969
rect 16866 -17003 16878 -16969
rect 16820 -17037 16878 -17003
rect 16820 -17071 16832 -17037
rect 16866 -17071 16878 -17037
rect 16820 -17105 16878 -17071
rect 16820 -17139 16832 -17105
rect 16866 -17139 16878 -17105
rect 16820 -17173 16878 -17139
rect 16820 -17207 16832 -17173
rect 16866 -17207 16878 -17173
rect 16820 -17252 16878 -17207
rect 17838 -16697 17896 -16652
rect 17838 -16731 17850 -16697
rect 17884 -16731 17896 -16697
rect 17838 -16765 17896 -16731
rect 17838 -16799 17850 -16765
rect 17884 -16799 17896 -16765
rect 17838 -16833 17896 -16799
rect 17838 -16867 17850 -16833
rect 17884 -16867 17896 -16833
rect 17838 -16901 17896 -16867
rect 17838 -16935 17850 -16901
rect 17884 -16935 17896 -16901
rect 17838 -16969 17896 -16935
rect 17838 -17003 17850 -16969
rect 17884 -17003 17896 -16969
rect 17838 -17037 17896 -17003
rect 17838 -17071 17850 -17037
rect 17884 -17071 17896 -17037
rect 17838 -17105 17896 -17071
rect 17838 -17139 17850 -17105
rect 17884 -17139 17896 -17105
rect 17838 -17173 17896 -17139
rect 17838 -17207 17850 -17173
rect 17884 -17207 17896 -17173
rect 17838 -17252 17896 -17207
rect 18856 -16697 18914 -16652
rect 18856 -16731 18868 -16697
rect 18902 -16731 18914 -16697
rect 18856 -16765 18914 -16731
rect 18856 -16799 18868 -16765
rect 18902 -16799 18914 -16765
rect 18856 -16833 18914 -16799
rect 18856 -16867 18868 -16833
rect 18902 -16867 18914 -16833
rect 18856 -16901 18914 -16867
rect 18856 -16935 18868 -16901
rect 18902 -16935 18914 -16901
rect 18856 -16969 18914 -16935
rect 18856 -17003 18868 -16969
rect 18902 -17003 18914 -16969
rect 18856 -17037 18914 -17003
rect 18856 -17071 18868 -17037
rect 18902 -17071 18914 -17037
rect 18856 -17105 18914 -17071
rect 18856 -17139 18868 -17105
rect 18902 -17139 18914 -17105
rect 18856 -17173 18914 -17139
rect 18856 -17207 18868 -17173
rect 18902 -17207 18914 -17173
rect 18856 -17252 18914 -17207
rect 19874 -16697 19932 -16652
rect 19874 -16731 19886 -16697
rect 19920 -16731 19932 -16697
rect 19874 -16765 19932 -16731
rect 19874 -16799 19886 -16765
rect 19920 -16799 19932 -16765
rect 19874 -16833 19932 -16799
rect 19874 -16867 19886 -16833
rect 19920 -16867 19932 -16833
rect 19874 -16901 19932 -16867
rect 19874 -16935 19886 -16901
rect 19920 -16935 19932 -16901
rect 19874 -16969 19932 -16935
rect 19874 -17003 19886 -16969
rect 19920 -17003 19932 -16969
rect 19874 -17037 19932 -17003
rect 19874 -17071 19886 -17037
rect 19920 -17071 19932 -17037
rect 19874 -17105 19932 -17071
rect 19874 -17139 19886 -17105
rect 19920 -17139 19932 -17105
rect 19874 -17173 19932 -17139
rect 19874 -17207 19886 -17173
rect 19920 -17207 19932 -17173
rect 19874 -17252 19932 -17207
rect 20892 -16697 20950 -16652
rect 20892 -16731 20904 -16697
rect 20938 -16731 20950 -16697
rect 20892 -16765 20950 -16731
rect 20892 -16799 20904 -16765
rect 20938 -16799 20950 -16765
rect 20892 -16833 20950 -16799
rect 20892 -16867 20904 -16833
rect 20938 -16867 20950 -16833
rect 20892 -16901 20950 -16867
rect 20892 -16935 20904 -16901
rect 20938 -16935 20950 -16901
rect 20892 -16969 20950 -16935
rect 20892 -17003 20904 -16969
rect 20938 -17003 20950 -16969
rect 20892 -17037 20950 -17003
rect 20892 -17071 20904 -17037
rect 20938 -17071 20950 -17037
rect 20892 -17105 20950 -17071
rect 20892 -17139 20904 -17105
rect 20938 -17139 20950 -17105
rect 20892 -17173 20950 -17139
rect 20892 -17207 20904 -17173
rect 20938 -17207 20950 -17173
rect 20892 -17252 20950 -17207
rect 21910 -16697 21968 -16652
rect 21910 -16731 21922 -16697
rect 21956 -16731 21968 -16697
rect 21910 -16765 21968 -16731
rect 21910 -16799 21922 -16765
rect 21956 -16799 21968 -16765
rect 21910 -16833 21968 -16799
rect 21910 -16867 21922 -16833
rect 21956 -16867 21968 -16833
rect 21910 -16901 21968 -16867
rect 21910 -16935 21922 -16901
rect 21956 -16935 21968 -16901
rect 21910 -16969 21968 -16935
rect 21910 -17003 21922 -16969
rect 21956 -17003 21968 -16969
rect 21910 -17037 21968 -17003
rect 21910 -17071 21922 -17037
rect 21956 -17071 21968 -17037
rect 21910 -17105 21968 -17071
rect 21910 -17139 21922 -17105
rect 21956 -17139 21968 -17105
rect 21910 -17173 21968 -17139
rect 21910 -17207 21922 -17173
rect 21956 -17207 21968 -17173
rect 21910 -17252 21968 -17207
rect 22928 -16697 22986 -16652
rect 22928 -16731 22940 -16697
rect 22974 -16731 22986 -16697
rect 22928 -16765 22986 -16731
rect 22928 -16799 22940 -16765
rect 22974 -16799 22986 -16765
rect 22928 -16833 22986 -16799
rect 22928 -16867 22940 -16833
rect 22974 -16867 22986 -16833
rect 22928 -16901 22986 -16867
rect 22928 -16935 22940 -16901
rect 22974 -16935 22986 -16901
rect 22928 -16969 22986 -16935
rect 22928 -17003 22940 -16969
rect 22974 -17003 22986 -16969
rect 22928 -17037 22986 -17003
rect 22928 -17071 22940 -17037
rect 22974 -17071 22986 -17037
rect 22928 -17105 22986 -17071
rect 22928 -17139 22940 -17105
rect 22974 -17139 22986 -17105
rect 22928 -17173 22986 -17139
rect 22928 -17207 22940 -17173
rect 22974 -17207 22986 -17173
rect 22928 -17252 22986 -17207
rect -9196 -17465 -9138 -17420
rect -9196 -17499 -9184 -17465
rect -9150 -17499 -9138 -17465
rect -9196 -17533 -9138 -17499
rect -9196 -17567 -9184 -17533
rect -9150 -17567 -9138 -17533
rect -9196 -17601 -9138 -17567
rect -9196 -17635 -9184 -17601
rect -9150 -17635 -9138 -17601
rect -9196 -17669 -9138 -17635
rect -9196 -17703 -9184 -17669
rect -9150 -17703 -9138 -17669
rect -9196 -17737 -9138 -17703
rect -9196 -17771 -9184 -17737
rect -9150 -17771 -9138 -17737
rect -9196 -17805 -9138 -17771
rect -9196 -17839 -9184 -17805
rect -9150 -17839 -9138 -17805
rect -9196 -17873 -9138 -17839
rect -9196 -17907 -9184 -17873
rect -9150 -17907 -9138 -17873
rect -9196 -17941 -9138 -17907
rect -9196 -17975 -9184 -17941
rect -9150 -17975 -9138 -17941
rect -9196 -18020 -9138 -17975
rect -8178 -17465 -8120 -17420
rect -8178 -17499 -8166 -17465
rect -8132 -17499 -8120 -17465
rect -8178 -17533 -8120 -17499
rect -8178 -17567 -8166 -17533
rect -8132 -17567 -8120 -17533
rect -8178 -17601 -8120 -17567
rect -8178 -17635 -8166 -17601
rect -8132 -17635 -8120 -17601
rect -8178 -17669 -8120 -17635
rect -8178 -17703 -8166 -17669
rect -8132 -17703 -8120 -17669
rect -8178 -17737 -8120 -17703
rect -8178 -17771 -8166 -17737
rect -8132 -17771 -8120 -17737
rect -8178 -17805 -8120 -17771
rect -8178 -17839 -8166 -17805
rect -8132 -17839 -8120 -17805
rect -8178 -17873 -8120 -17839
rect -8178 -17907 -8166 -17873
rect -8132 -17907 -8120 -17873
rect -8178 -17941 -8120 -17907
rect -8178 -17975 -8166 -17941
rect -8132 -17975 -8120 -17941
rect -8178 -18020 -8120 -17975
rect -7160 -17465 -7102 -17420
rect -7160 -17499 -7148 -17465
rect -7114 -17499 -7102 -17465
rect -7160 -17533 -7102 -17499
rect -7160 -17567 -7148 -17533
rect -7114 -17567 -7102 -17533
rect -7160 -17601 -7102 -17567
rect -7160 -17635 -7148 -17601
rect -7114 -17635 -7102 -17601
rect -7160 -17669 -7102 -17635
rect -7160 -17703 -7148 -17669
rect -7114 -17703 -7102 -17669
rect -7160 -17737 -7102 -17703
rect -7160 -17771 -7148 -17737
rect -7114 -17771 -7102 -17737
rect -7160 -17805 -7102 -17771
rect -7160 -17839 -7148 -17805
rect -7114 -17839 -7102 -17805
rect -7160 -17873 -7102 -17839
rect -7160 -17907 -7148 -17873
rect -7114 -17907 -7102 -17873
rect -7160 -17941 -7102 -17907
rect -7160 -17975 -7148 -17941
rect -7114 -17975 -7102 -17941
rect -7160 -18020 -7102 -17975
rect -6142 -17465 -6084 -17420
rect -6142 -17499 -6130 -17465
rect -6096 -17499 -6084 -17465
rect -6142 -17533 -6084 -17499
rect -6142 -17567 -6130 -17533
rect -6096 -17567 -6084 -17533
rect -6142 -17601 -6084 -17567
rect -6142 -17635 -6130 -17601
rect -6096 -17635 -6084 -17601
rect -6142 -17669 -6084 -17635
rect -6142 -17703 -6130 -17669
rect -6096 -17703 -6084 -17669
rect -6142 -17737 -6084 -17703
rect -6142 -17771 -6130 -17737
rect -6096 -17771 -6084 -17737
rect -6142 -17805 -6084 -17771
rect -6142 -17839 -6130 -17805
rect -6096 -17839 -6084 -17805
rect -6142 -17873 -6084 -17839
rect -6142 -17907 -6130 -17873
rect -6096 -17907 -6084 -17873
rect -6142 -17941 -6084 -17907
rect -6142 -17975 -6130 -17941
rect -6096 -17975 -6084 -17941
rect -6142 -18020 -6084 -17975
rect -5124 -17465 -5066 -17420
rect -5124 -17499 -5112 -17465
rect -5078 -17499 -5066 -17465
rect -5124 -17533 -5066 -17499
rect -5124 -17567 -5112 -17533
rect -5078 -17567 -5066 -17533
rect -5124 -17601 -5066 -17567
rect -5124 -17635 -5112 -17601
rect -5078 -17635 -5066 -17601
rect -5124 -17669 -5066 -17635
rect -5124 -17703 -5112 -17669
rect -5078 -17703 -5066 -17669
rect -5124 -17737 -5066 -17703
rect -5124 -17771 -5112 -17737
rect -5078 -17771 -5066 -17737
rect -5124 -17805 -5066 -17771
rect -5124 -17839 -5112 -17805
rect -5078 -17839 -5066 -17805
rect -5124 -17873 -5066 -17839
rect -5124 -17907 -5112 -17873
rect -5078 -17907 -5066 -17873
rect -5124 -17941 -5066 -17907
rect -5124 -17975 -5112 -17941
rect -5078 -17975 -5066 -17941
rect -5124 -18020 -5066 -17975
rect -4106 -17465 -4048 -17420
rect -4106 -17499 -4094 -17465
rect -4060 -17499 -4048 -17465
rect -4106 -17533 -4048 -17499
rect -4106 -17567 -4094 -17533
rect -4060 -17567 -4048 -17533
rect -4106 -17601 -4048 -17567
rect -4106 -17635 -4094 -17601
rect -4060 -17635 -4048 -17601
rect -4106 -17669 -4048 -17635
rect -4106 -17703 -4094 -17669
rect -4060 -17703 -4048 -17669
rect -4106 -17737 -4048 -17703
rect -4106 -17771 -4094 -17737
rect -4060 -17771 -4048 -17737
rect -4106 -17805 -4048 -17771
rect -4106 -17839 -4094 -17805
rect -4060 -17839 -4048 -17805
rect -4106 -17873 -4048 -17839
rect -4106 -17907 -4094 -17873
rect -4060 -17907 -4048 -17873
rect -4106 -17941 -4048 -17907
rect -4106 -17975 -4094 -17941
rect -4060 -17975 -4048 -17941
rect -4106 -18020 -4048 -17975
rect -3088 -17465 -3030 -17420
rect -3088 -17499 -3076 -17465
rect -3042 -17499 -3030 -17465
rect -3088 -17533 -3030 -17499
rect -3088 -17567 -3076 -17533
rect -3042 -17567 -3030 -17533
rect -3088 -17601 -3030 -17567
rect -3088 -17635 -3076 -17601
rect -3042 -17635 -3030 -17601
rect -3088 -17669 -3030 -17635
rect -3088 -17703 -3076 -17669
rect -3042 -17703 -3030 -17669
rect -3088 -17737 -3030 -17703
rect -3088 -17771 -3076 -17737
rect -3042 -17771 -3030 -17737
rect -3088 -17805 -3030 -17771
rect -3088 -17839 -3076 -17805
rect -3042 -17839 -3030 -17805
rect -3088 -17873 -3030 -17839
rect -3088 -17907 -3076 -17873
rect -3042 -17907 -3030 -17873
rect -3088 -17941 -3030 -17907
rect -3088 -17975 -3076 -17941
rect -3042 -17975 -3030 -17941
rect -3088 -18020 -3030 -17975
rect -2070 -17465 -2012 -17420
rect -2070 -17499 -2058 -17465
rect -2024 -17499 -2012 -17465
rect -2070 -17533 -2012 -17499
rect -2070 -17567 -2058 -17533
rect -2024 -17567 -2012 -17533
rect -2070 -17601 -2012 -17567
rect -2070 -17635 -2058 -17601
rect -2024 -17635 -2012 -17601
rect -2070 -17669 -2012 -17635
rect -2070 -17703 -2058 -17669
rect -2024 -17703 -2012 -17669
rect -2070 -17737 -2012 -17703
rect -2070 -17771 -2058 -17737
rect -2024 -17771 -2012 -17737
rect -2070 -17805 -2012 -17771
rect -2070 -17839 -2058 -17805
rect -2024 -17839 -2012 -17805
rect -2070 -17873 -2012 -17839
rect -2070 -17907 -2058 -17873
rect -2024 -17907 -2012 -17873
rect -2070 -17941 -2012 -17907
rect -2070 -17975 -2058 -17941
rect -2024 -17975 -2012 -17941
rect -2070 -18020 -2012 -17975
rect -1052 -17465 -994 -17420
rect -1052 -17499 -1040 -17465
rect -1006 -17499 -994 -17465
rect -1052 -17533 -994 -17499
rect -1052 -17567 -1040 -17533
rect -1006 -17567 -994 -17533
rect -1052 -17601 -994 -17567
rect -1052 -17635 -1040 -17601
rect -1006 -17635 -994 -17601
rect -1052 -17669 -994 -17635
rect -1052 -17703 -1040 -17669
rect -1006 -17703 -994 -17669
rect -1052 -17737 -994 -17703
rect -1052 -17771 -1040 -17737
rect -1006 -17771 -994 -17737
rect -1052 -17805 -994 -17771
rect -1052 -17839 -1040 -17805
rect -1006 -17839 -994 -17805
rect -1052 -17873 -994 -17839
rect -1052 -17907 -1040 -17873
rect -1006 -17907 -994 -17873
rect -1052 -17941 -994 -17907
rect -1052 -17975 -1040 -17941
rect -1006 -17975 -994 -17941
rect -1052 -18020 -994 -17975
rect -34 -17465 24 -17420
rect -34 -17499 -22 -17465
rect 12 -17499 24 -17465
rect -34 -17533 24 -17499
rect -34 -17567 -22 -17533
rect 12 -17567 24 -17533
rect -34 -17601 24 -17567
rect -34 -17635 -22 -17601
rect 12 -17635 24 -17601
rect -34 -17669 24 -17635
rect -34 -17703 -22 -17669
rect 12 -17703 24 -17669
rect -34 -17737 24 -17703
rect -34 -17771 -22 -17737
rect 12 -17771 24 -17737
rect -34 -17805 24 -17771
rect -34 -17839 -22 -17805
rect 12 -17839 24 -17805
rect -34 -17873 24 -17839
rect -34 -17907 -22 -17873
rect 12 -17907 24 -17873
rect -34 -17941 24 -17907
rect -34 -17975 -22 -17941
rect 12 -17975 24 -17941
rect -34 -18020 24 -17975
rect 2568 -17929 2626 -17884
rect 2568 -17963 2580 -17929
rect 2614 -17963 2626 -17929
rect 2568 -17997 2626 -17963
rect 2568 -18031 2580 -17997
rect 2614 -18031 2626 -17997
rect 2568 -18065 2626 -18031
rect 2568 -18099 2580 -18065
rect 2614 -18099 2626 -18065
rect 2568 -18133 2626 -18099
rect 2568 -18167 2580 -18133
rect 2614 -18167 2626 -18133
rect 2568 -18201 2626 -18167
rect 2568 -18235 2580 -18201
rect 2614 -18235 2626 -18201
rect -9196 -18283 -9138 -18238
rect -9196 -18317 -9184 -18283
rect -9150 -18317 -9138 -18283
rect -9196 -18351 -9138 -18317
rect -9196 -18385 -9184 -18351
rect -9150 -18385 -9138 -18351
rect -9196 -18419 -9138 -18385
rect -9196 -18453 -9184 -18419
rect -9150 -18453 -9138 -18419
rect -9196 -18487 -9138 -18453
rect -9196 -18521 -9184 -18487
rect -9150 -18521 -9138 -18487
rect -9196 -18555 -9138 -18521
rect -9196 -18589 -9184 -18555
rect -9150 -18589 -9138 -18555
rect -9196 -18623 -9138 -18589
rect -9196 -18657 -9184 -18623
rect -9150 -18657 -9138 -18623
rect -9196 -18691 -9138 -18657
rect -9196 -18725 -9184 -18691
rect -9150 -18725 -9138 -18691
rect -9196 -18759 -9138 -18725
rect -9196 -18793 -9184 -18759
rect -9150 -18793 -9138 -18759
rect -9196 -18838 -9138 -18793
rect -8178 -18283 -8120 -18238
rect -8178 -18317 -8166 -18283
rect -8132 -18317 -8120 -18283
rect -8178 -18351 -8120 -18317
rect -8178 -18385 -8166 -18351
rect -8132 -18385 -8120 -18351
rect -8178 -18419 -8120 -18385
rect -8178 -18453 -8166 -18419
rect -8132 -18453 -8120 -18419
rect -8178 -18487 -8120 -18453
rect -8178 -18521 -8166 -18487
rect -8132 -18521 -8120 -18487
rect -8178 -18555 -8120 -18521
rect -8178 -18589 -8166 -18555
rect -8132 -18589 -8120 -18555
rect -8178 -18623 -8120 -18589
rect -8178 -18657 -8166 -18623
rect -8132 -18657 -8120 -18623
rect -8178 -18691 -8120 -18657
rect -8178 -18725 -8166 -18691
rect -8132 -18725 -8120 -18691
rect -8178 -18759 -8120 -18725
rect -8178 -18793 -8166 -18759
rect -8132 -18793 -8120 -18759
rect -8178 -18838 -8120 -18793
rect -7160 -18283 -7102 -18238
rect -7160 -18317 -7148 -18283
rect -7114 -18317 -7102 -18283
rect -7160 -18351 -7102 -18317
rect -7160 -18385 -7148 -18351
rect -7114 -18385 -7102 -18351
rect -7160 -18419 -7102 -18385
rect -7160 -18453 -7148 -18419
rect -7114 -18453 -7102 -18419
rect -7160 -18487 -7102 -18453
rect -7160 -18521 -7148 -18487
rect -7114 -18521 -7102 -18487
rect -7160 -18555 -7102 -18521
rect -7160 -18589 -7148 -18555
rect -7114 -18589 -7102 -18555
rect -7160 -18623 -7102 -18589
rect -7160 -18657 -7148 -18623
rect -7114 -18657 -7102 -18623
rect -7160 -18691 -7102 -18657
rect -7160 -18725 -7148 -18691
rect -7114 -18725 -7102 -18691
rect -7160 -18759 -7102 -18725
rect -7160 -18793 -7148 -18759
rect -7114 -18793 -7102 -18759
rect -7160 -18838 -7102 -18793
rect -6142 -18283 -6084 -18238
rect -6142 -18317 -6130 -18283
rect -6096 -18317 -6084 -18283
rect -6142 -18351 -6084 -18317
rect -6142 -18385 -6130 -18351
rect -6096 -18385 -6084 -18351
rect -6142 -18419 -6084 -18385
rect -6142 -18453 -6130 -18419
rect -6096 -18453 -6084 -18419
rect -6142 -18487 -6084 -18453
rect -6142 -18521 -6130 -18487
rect -6096 -18521 -6084 -18487
rect -6142 -18555 -6084 -18521
rect -6142 -18589 -6130 -18555
rect -6096 -18589 -6084 -18555
rect -6142 -18623 -6084 -18589
rect -6142 -18657 -6130 -18623
rect -6096 -18657 -6084 -18623
rect -6142 -18691 -6084 -18657
rect -6142 -18725 -6130 -18691
rect -6096 -18725 -6084 -18691
rect -6142 -18759 -6084 -18725
rect -6142 -18793 -6130 -18759
rect -6096 -18793 -6084 -18759
rect -6142 -18838 -6084 -18793
rect -5124 -18283 -5066 -18238
rect -5124 -18317 -5112 -18283
rect -5078 -18317 -5066 -18283
rect -5124 -18351 -5066 -18317
rect -5124 -18385 -5112 -18351
rect -5078 -18385 -5066 -18351
rect -5124 -18419 -5066 -18385
rect -5124 -18453 -5112 -18419
rect -5078 -18453 -5066 -18419
rect -5124 -18487 -5066 -18453
rect -5124 -18521 -5112 -18487
rect -5078 -18521 -5066 -18487
rect -5124 -18555 -5066 -18521
rect -5124 -18589 -5112 -18555
rect -5078 -18589 -5066 -18555
rect -5124 -18623 -5066 -18589
rect -5124 -18657 -5112 -18623
rect -5078 -18657 -5066 -18623
rect -5124 -18691 -5066 -18657
rect -5124 -18725 -5112 -18691
rect -5078 -18725 -5066 -18691
rect -5124 -18759 -5066 -18725
rect -5124 -18793 -5112 -18759
rect -5078 -18793 -5066 -18759
rect -5124 -18838 -5066 -18793
rect -4106 -18283 -4048 -18238
rect -4106 -18317 -4094 -18283
rect -4060 -18317 -4048 -18283
rect -4106 -18351 -4048 -18317
rect -4106 -18385 -4094 -18351
rect -4060 -18385 -4048 -18351
rect -4106 -18419 -4048 -18385
rect -4106 -18453 -4094 -18419
rect -4060 -18453 -4048 -18419
rect -4106 -18487 -4048 -18453
rect -4106 -18521 -4094 -18487
rect -4060 -18521 -4048 -18487
rect -4106 -18555 -4048 -18521
rect -4106 -18589 -4094 -18555
rect -4060 -18589 -4048 -18555
rect -4106 -18623 -4048 -18589
rect -4106 -18657 -4094 -18623
rect -4060 -18657 -4048 -18623
rect -4106 -18691 -4048 -18657
rect -4106 -18725 -4094 -18691
rect -4060 -18725 -4048 -18691
rect -4106 -18759 -4048 -18725
rect -4106 -18793 -4094 -18759
rect -4060 -18793 -4048 -18759
rect -4106 -18838 -4048 -18793
rect -3088 -18283 -3030 -18238
rect -3088 -18317 -3076 -18283
rect -3042 -18317 -3030 -18283
rect -3088 -18351 -3030 -18317
rect -3088 -18385 -3076 -18351
rect -3042 -18385 -3030 -18351
rect -3088 -18419 -3030 -18385
rect -3088 -18453 -3076 -18419
rect -3042 -18453 -3030 -18419
rect -3088 -18487 -3030 -18453
rect -3088 -18521 -3076 -18487
rect -3042 -18521 -3030 -18487
rect -3088 -18555 -3030 -18521
rect -3088 -18589 -3076 -18555
rect -3042 -18589 -3030 -18555
rect -3088 -18623 -3030 -18589
rect -3088 -18657 -3076 -18623
rect -3042 -18657 -3030 -18623
rect -3088 -18691 -3030 -18657
rect -3088 -18725 -3076 -18691
rect -3042 -18725 -3030 -18691
rect -3088 -18759 -3030 -18725
rect -3088 -18793 -3076 -18759
rect -3042 -18793 -3030 -18759
rect -3088 -18838 -3030 -18793
rect -2070 -18283 -2012 -18238
rect -2070 -18317 -2058 -18283
rect -2024 -18317 -2012 -18283
rect -2070 -18351 -2012 -18317
rect -2070 -18385 -2058 -18351
rect -2024 -18385 -2012 -18351
rect -2070 -18419 -2012 -18385
rect -2070 -18453 -2058 -18419
rect -2024 -18453 -2012 -18419
rect -2070 -18487 -2012 -18453
rect -2070 -18521 -2058 -18487
rect -2024 -18521 -2012 -18487
rect -2070 -18555 -2012 -18521
rect -2070 -18589 -2058 -18555
rect -2024 -18589 -2012 -18555
rect -2070 -18623 -2012 -18589
rect -2070 -18657 -2058 -18623
rect -2024 -18657 -2012 -18623
rect -2070 -18691 -2012 -18657
rect -2070 -18725 -2058 -18691
rect -2024 -18725 -2012 -18691
rect -2070 -18759 -2012 -18725
rect -2070 -18793 -2058 -18759
rect -2024 -18793 -2012 -18759
rect -2070 -18838 -2012 -18793
rect -1052 -18283 -994 -18238
rect -1052 -18317 -1040 -18283
rect -1006 -18317 -994 -18283
rect -1052 -18351 -994 -18317
rect -1052 -18385 -1040 -18351
rect -1006 -18385 -994 -18351
rect -1052 -18419 -994 -18385
rect -1052 -18453 -1040 -18419
rect -1006 -18453 -994 -18419
rect -1052 -18487 -994 -18453
rect -1052 -18521 -1040 -18487
rect -1006 -18521 -994 -18487
rect -1052 -18555 -994 -18521
rect -1052 -18589 -1040 -18555
rect -1006 -18589 -994 -18555
rect -1052 -18623 -994 -18589
rect -1052 -18657 -1040 -18623
rect -1006 -18657 -994 -18623
rect -1052 -18691 -994 -18657
rect -1052 -18725 -1040 -18691
rect -1006 -18725 -994 -18691
rect -1052 -18759 -994 -18725
rect -1052 -18793 -1040 -18759
rect -1006 -18793 -994 -18759
rect -1052 -18838 -994 -18793
rect -34 -18283 24 -18238
rect -34 -18317 -22 -18283
rect 12 -18317 24 -18283
rect -34 -18351 24 -18317
rect -34 -18385 -22 -18351
rect 12 -18385 24 -18351
rect -34 -18419 24 -18385
rect -34 -18453 -22 -18419
rect 12 -18453 24 -18419
rect -34 -18487 24 -18453
rect 2568 -18269 2626 -18235
rect 2568 -18303 2580 -18269
rect 2614 -18303 2626 -18269
rect 2568 -18337 2626 -18303
rect 2568 -18371 2580 -18337
rect 2614 -18371 2626 -18337
rect 2568 -18405 2626 -18371
rect 2568 -18439 2580 -18405
rect 2614 -18439 2626 -18405
rect 2568 -18484 2626 -18439
rect 3586 -17929 3644 -17884
rect 3586 -17963 3598 -17929
rect 3632 -17963 3644 -17929
rect 3586 -17997 3644 -17963
rect 3586 -18031 3598 -17997
rect 3632 -18031 3644 -17997
rect 3586 -18065 3644 -18031
rect 3586 -18099 3598 -18065
rect 3632 -18099 3644 -18065
rect 3586 -18133 3644 -18099
rect 3586 -18167 3598 -18133
rect 3632 -18167 3644 -18133
rect 3586 -18201 3644 -18167
rect 3586 -18235 3598 -18201
rect 3632 -18235 3644 -18201
rect 3586 -18269 3644 -18235
rect 3586 -18303 3598 -18269
rect 3632 -18303 3644 -18269
rect 3586 -18337 3644 -18303
rect 3586 -18371 3598 -18337
rect 3632 -18371 3644 -18337
rect 3586 -18405 3644 -18371
rect 3586 -18439 3598 -18405
rect 3632 -18439 3644 -18405
rect 3586 -18484 3644 -18439
rect 4604 -17929 4662 -17884
rect 4604 -17963 4616 -17929
rect 4650 -17963 4662 -17929
rect 4604 -17997 4662 -17963
rect 4604 -18031 4616 -17997
rect 4650 -18031 4662 -17997
rect 4604 -18065 4662 -18031
rect 4604 -18099 4616 -18065
rect 4650 -18099 4662 -18065
rect 4604 -18133 4662 -18099
rect 4604 -18167 4616 -18133
rect 4650 -18167 4662 -18133
rect 4604 -18201 4662 -18167
rect 4604 -18235 4616 -18201
rect 4650 -18235 4662 -18201
rect 4604 -18269 4662 -18235
rect 4604 -18303 4616 -18269
rect 4650 -18303 4662 -18269
rect 4604 -18337 4662 -18303
rect 4604 -18371 4616 -18337
rect 4650 -18371 4662 -18337
rect 4604 -18405 4662 -18371
rect 4604 -18439 4616 -18405
rect 4650 -18439 4662 -18405
rect 4604 -18484 4662 -18439
rect 5622 -17929 5680 -17884
rect 5622 -17963 5634 -17929
rect 5668 -17963 5680 -17929
rect 5622 -17997 5680 -17963
rect 5622 -18031 5634 -17997
rect 5668 -18031 5680 -17997
rect 5622 -18065 5680 -18031
rect 5622 -18099 5634 -18065
rect 5668 -18099 5680 -18065
rect 5622 -18133 5680 -18099
rect 5622 -18167 5634 -18133
rect 5668 -18167 5680 -18133
rect 5622 -18201 5680 -18167
rect 5622 -18235 5634 -18201
rect 5668 -18235 5680 -18201
rect 5622 -18269 5680 -18235
rect 5622 -18303 5634 -18269
rect 5668 -18303 5680 -18269
rect 5622 -18337 5680 -18303
rect 5622 -18371 5634 -18337
rect 5668 -18371 5680 -18337
rect 5622 -18405 5680 -18371
rect 5622 -18439 5634 -18405
rect 5668 -18439 5680 -18405
rect 5622 -18484 5680 -18439
rect 6640 -17929 6698 -17884
rect 6640 -17963 6652 -17929
rect 6686 -17963 6698 -17929
rect 6640 -17997 6698 -17963
rect 6640 -18031 6652 -17997
rect 6686 -18031 6698 -17997
rect 6640 -18065 6698 -18031
rect 6640 -18099 6652 -18065
rect 6686 -18099 6698 -18065
rect 6640 -18133 6698 -18099
rect 6640 -18167 6652 -18133
rect 6686 -18167 6698 -18133
rect 6640 -18201 6698 -18167
rect 6640 -18235 6652 -18201
rect 6686 -18235 6698 -18201
rect 6640 -18269 6698 -18235
rect 6640 -18303 6652 -18269
rect 6686 -18303 6698 -18269
rect 6640 -18337 6698 -18303
rect 6640 -18371 6652 -18337
rect 6686 -18371 6698 -18337
rect 6640 -18405 6698 -18371
rect 6640 -18439 6652 -18405
rect 6686 -18439 6698 -18405
rect 6640 -18484 6698 -18439
rect 7658 -17929 7716 -17884
rect 7658 -17963 7670 -17929
rect 7704 -17963 7716 -17929
rect 7658 -17997 7716 -17963
rect 7658 -18031 7670 -17997
rect 7704 -18031 7716 -17997
rect 7658 -18065 7716 -18031
rect 7658 -18099 7670 -18065
rect 7704 -18099 7716 -18065
rect 7658 -18133 7716 -18099
rect 7658 -18167 7670 -18133
rect 7704 -18167 7716 -18133
rect 7658 -18201 7716 -18167
rect 7658 -18235 7670 -18201
rect 7704 -18235 7716 -18201
rect 7658 -18269 7716 -18235
rect 7658 -18303 7670 -18269
rect 7704 -18303 7716 -18269
rect 7658 -18337 7716 -18303
rect 7658 -18371 7670 -18337
rect 7704 -18371 7716 -18337
rect 7658 -18405 7716 -18371
rect 7658 -18439 7670 -18405
rect 7704 -18439 7716 -18405
rect 7658 -18484 7716 -18439
rect 8676 -17929 8734 -17884
rect 8676 -17963 8688 -17929
rect 8722 -17963 8734 -17929
rect 8676 -17997 8734 -17963
rect 8676 -18031 8688 -17997
rect 8722 -18031 8734 -17997
rect 8676 -18065 8734 -18031
rect 8676 -18099 8688 -18065
rect 8722 -18099 8734 -18065
rect 8676 -18133 8734 -18099
rect 8676 -18167 8688 -18133
rect 8722 -18167 8734 -18133
rect 8676 -18201 8734 -18167
rect 8676 -18235 8688 -18201
rect 8722 -18235 8734 -18201
rect 8676 -18269 8734 -18235
rect 8676 -18303 8688 -18269
rect 8722 -18303 8734 -18269
rect 8676 -18337 8734 -18303
rect 8676 -18371 8688 -18337
rect 8722 -18371 8734 -18337
rect 8676 -18405 8734 -18371
rect 8676 -18439 8688 -18405
rect 8722 -18439 8734 -18405
rect 8676 -18484 8734 -18439
rect 9694 -17929 9752 -17884
rect 9694 -17963 9706 -17929
rect 9740 -17963 9752 -17929
rect 9694 -17997 9752 -17963
rect 9694 -18031 9706 -17997
rect 9740 -18031 9752 -17997
rect 9694 -18065 9752 -18031
rect 9694 -18099 9706 -18065
rect 9740 -18099 9752 -18065
rect 9694 -18133 9752 -18099
rect 9694 -18167 9706 -18133
rect 9740 -18167 9752 -18133
rect 9694 -18201 9752 -18167
rect 9694 -18235 9706 -18201
rect 9740 -18235 9752 -18201
rect 9694 -18269 9752 -18235
rect 9694 -18303 9706 -18269
rect 9740 -18303 9752 -18269
rect 9694 -18337 9752 -18303
rect 9694 -18371 9706 -18337
rect 9740 -18371 9752 -18337
rect 9694 -18405 9752 -18371
rect 9694 -18439 9706 -18405
rect 9740 -18439 9752 -18405
rect 9694 -18484 9752 -18439
rect 10712 -17929 10770 -17884
rect 10712 -17963 10724 -17929
rect 10758 -17963 10770 -17929
rect 10712 -17997 10770 -17963
rect 10712 -18031 10724 -17997
rect 10758 -18031 10770 -17997
rect 10712 -18065 10770 -18031
rect 10712 -18099 10724 -18065
rect 10758 -18099 10770 -18065
rect 10712 -18133 10770 -18099
rect 10712 -18167 10724 -18133
rect 10758 -18167 10770 -18133
rect 10712 -18201 10770 -18167
rect 10712 -18235 10724 -18201
rect 10758 -18235 10770 -18201
rect 10712 -18269 10770 -18235
rect 10712 -18303 10724 -18269
rect 10758 -18303 10770 -18269
rect 10712 -18337 10770 -18303
rect 10712 -18371 10724 -18337
rect 10758 -18371 10770 -18337
rect 10712 -18405 10770 -18371
rect 10712 -18439 10724 -18405
rect 10758 -18439 10770 -18405
rect 10712 -18484 10770 -18439
rect 11730 -17929 11788 -17884
rect 11730 -17963 11742 -17929
rect 11776 -17963 11788 -17929
rect 11730 -17997 11788 -17963
rect 11730 -18031 11742 -17997
rect 11776 -18031 11788 -17997
rect 11730 -18065 11788 -18031
rect 11730 -18099 11742 -18065
rect 11776 -18099 11788 -18065
rect 11730 -18133 11788 -18099
rect 11730 -18167 11742 -18133
rect 11776 -18167 11788 -18133
rect 11730 -18201 11788 -18167
rect 11730 -18235 11742 -18201
rect 11776 -18235 11788 -18201
rect 11730 -18269 11788 -18235
rect 11730 -18303 11742 -18269
rect 11776 -18303 11788 -18269
rect 11730 -18337 11788 -18303
rect 11730 -18371 11742 -18337
rect 11776 -18371 11788 -18337
rect 11730 -18405 11788 -18371
rect 11730 -18439 11742 -18405
rect 11776 -18439 11788 -18405
rect 11730 -18484 11788 -18439
rect 12748 -17929 12806 -17884
rect 12748 -17963 12760 -17929
rect 12794 -17963 12806 -17929
rect 12748 -17997 12806 -17963
rect 12748 -18031 12760 -17997
rect 12794 -18031 12806 -17997
rect 12748 -18065 12806 -18031
rect 12748 -18099 12760 -18065
rect 12794 -18099 12806 -18065
rect 12748 -18133 12806 -18099
rect 12748 -18167 12760 -18133
rect 12794 -18167 12806 -18133
rect 12748 -18201 12806 -18167
rect 12748 -18235 12760 -18201
rect 12794 -18235 12806 -18201
rect 12748 -18269 12806 -18235
rect 12748 -18303 12760 -18269
rect 12794 -18303 12806 -18269
rect 12748 -18337 12806 -18303
rect 12748 -18371 12760 -18337
rect 12794 -18371 12806 -18337
rect 12748 -18405 12806 -18371
rect 12748 -18439 12760 -18405
rect 12794 -18439 12806 -18405
rect 12748 -18484 12806 -18439
rect 13766 -17929 13824 -17884
rect 13766 -17963 13778 -17929
rect 13812 -17963 13824 -17929
rect 13766 -17997 13824 -17963
rect 13766 -18031 13778 -17997
rect 13812 -18031 13824 -17997
rect 13766 -18065 13824 -18031
rect 13766 -18099 13778 -18065
rect 13812 -18099 13824 -18065
rect 13766 -18133 13824 -18099
rect 13766 -18167 13778 -18133
rect 13812 -18167 13824 -18133
rect 13766 -18201 13824 -18167
rect 13766 -18235 13778 -18201
rect 13812 -18235 13824 -18201
rect 13766 -18269 13824 -18235
rect 13766 -18303 13778 -18269
rect 13812 -18303 13824 -18269
rect 13766 -18337 13824 -18303
rect 13766 -18371 13778 -18337
rect 13812 -18371 13824 -18337
rect 13766 -18405 13824 -18371
rect 13766 -18439 13778 -18405
rect 13812 -18439 13824 -18405
rect 13766 -18484 13824 -18439
rect 14784 -17929 14842 -17884
rect 14784 -17963 14796 -17929
rect 14830 -17963 14842 -17929
rect 14784 -17997 14842 -17963
rect 14784 -18031 14796 -17997
rect 14830 -18031 14842 -17997
rect 14784 -18065 14842 -18031
rect 14784 -18099 14796 -18065
rect 14830 -18099 14842 -18065
rect 14784 -18133 14842 -18099
rect 14784 -18167 14796 -18133
rect 14830 -18167 14842 -18133
rect 14784 -18201 14842 -18167
rect 14784 -18235 14796 -18201
rect 14830 -18235 14842 -18201
rect 14784 -18269 14842 -18235
rect 14784 -18303 14796 -18269
rect 14830 -18303 14842 -18269
rect 14784 -18337 14842 -18303
rect 14784 -18371 14796 -18337
rect 14830 -18371 14842 -18337
rect 14784 -18405 14842 -18371
rect 14784 -18439 14796 -18405
rect 14830 -18439 14842 -18405
rect 14784 -18484 14842 -18439
rect 15802 -17929 15860 -17884
rect 15802 -17963 15814 -17929
rect 15848 -17963 15860 -17929
rect 15802 -17997 15860 -17963
rect 15802 -18031 15814 -17997
rect 15848 -18031 15860 -17997
rect 15802 -18065 15860 -18031
rect 15802 -18099 15814 -18065
rect 15848 -18099 15860 -18065
rect 15802 -18133 15860 -18099
rect 15802 -18167 15814 -18133
rect 15848 -18167 15860 -18133
rect 15802 -18201 15860 -18167
rect 15802 -18235 15814 -18201
rect 15848 -18235 15860 -18201
rect 15802 -18269 15860 -18235
rect 15802 -18303 15814 -18269
rect 15848 -18303 15860 -18269
rect 15802 -18337 15860 -18303
rect 15802 -18371 15814 -18337
rect 15848 -18371 15860 -18337
rect 15802 -18405 15860 -18371
rect 15802 -18439 15814 -18405
rect 15848 -18439 15860 -18405
rect 15802 -18484 15860 -18439
rect 16820 -17929 16878 -17884
rect 16820 -17963 16832 -17929
rect 16866 -17963 16878 -17929
rect 16820 -17997 16878 -17963
rect 16820 -18031 16832 -17997
rect 16866 -18031 16878 -17997
rect 16820 -18065 16878 -18031
rect 16820 -18099 16832 -18065
rect 16866 -18099 16878 -18065
rect 16820 -18133 16878 -18099
rect 16820 -18167 16832 -18133
rect 16866 -18167 16878 -18133
rect 16820 -18201 16878 -18167
rect 16820 -18235 16832 -18201
rect 16866 -18235 16878 -18201
rect 16820 -18269 16878 -18235
rect 16820 -18303 16832 -18269
rect 16866 -18303 16878 -18269
rect 16820 -18337 16878 -18303
rect 16820 -18371 16832 -18337
rect 16866 -18371 16878 -18337
rect 16820 -18405 16878 -18371
rect 16820 -18439 16832 -18405
rect 16866 -18439 16878 -18405
rect 16820 -18484 16878 -18439
rect 17838 -17929 17896 -17884
rect 17838 -17963 17850 -17929
rect 17884 -17963 17896 -17929
rect 17838 -17997 17896 -17963
rect 17838 -18031 17850 -17997
rect 17884 -18031 17896 -17997
rect 17838 -18065 17896 -18031
rect 17838 -18099 17850 -18065
rect 17884 -18099 17896 -18065
rect 17838 -18133 17896 -18099
rect 17838 -18167 17850 -18133
rect 17884 -18167 17896 -18133
rect 17838 -18201 17896 -18167
rect 17838 -18235 17850 -18201
rect 17884 -18235 17896 -18201
rect 17838 -18269 17896 -18235
rect 17838 -18303 17850 -18269
rect 17884 -18303 17896 -18269
rect 17838 -18337 17896 -18303
rect 17838 -18371 17850 -18337
rect 17884 -18371 17896 -18337
rect 17838 -18405 17896 -18371
rect 17838 -18439 17850 -18405
rect 17884 -18439 17896 -18405
rect 17838 -18484 17896 -18439
rect 18856 -17929 18914 -17884
rect 18856 -17963 18868 -17929
rect 18902 -17963 18914 -17929
rect 18856 -17997 18914 -17963
rect 18856 -18031 18868 -17997
rect 18902 -18031 18914 -17997
rect 18856 -18065 18914 -18031
rect 18856 -18099 18868 -18065
rect 18902 -18099 18914 -18065
rect 18856 -18133 18914 -18099
rect 18856 -18167 18868 -18133
rect 18902 -18167 18914 -18133
rect 18856 -18201 18914 -18167
rect 18856 -18235 18868 -18201
rect 18902 -18235 18914 -18201
rect 18856 -18269 18914 -18235
rect 18856 -18303 18868 -18269
rect 18902 -18303 18914 -18269
rect 18856 -18337 18914 -18303
rect 18856 -18371 18868 -18337
rect 18902 -18371 18914 -18337
rect 18856 -18405 18914 -18371
rect 18856 -18439 18868 -18405
rect 18902 -18439 18914 -18405
rect 18856 -18484 18914 -18439
rect 19874 -17929 19932 -17884
rect 19874 -17963 19886 -17929
rect 19920 -17963 19932 -17929
rect 19874 -17997 19932 -17963
rect 19874 -18031 19886 -17997
rect 19920 -18031 19932 -17997
rect 19874 -18065 19932 -18031
rect 19874 -18099 19886 -18065
rect 19920 -18099 19932 -18065
rect 19874 -18133 19932 -18099
rect 19874 -18167 19886 -18133
rect 19920 -18167 19932 -18133
rect 19874 -18201 19932 -18167
rect 19874 -18235 19886 -18201
rect 19920 -18235 19932 -18201
rect 19874 -18269 19932 -18235
rect 19874 -18303 19886 -18269
rect 19920 -18303 19932 -18269
rect 19874 -18337 19932 -18303
rect 19874 -18371 19886 -18337
rect 19920 -18371 19932 -18337
rect 19874 -18405 19932 -18371
rect 19874 -18439 19886 -18405
rect 19920 -18439 19932 -18405
rect 19874 -18484 19932 -18439
rect 20892 -17929 20950 -17884
rect 20892 -17963 20904 -17929
rect 20938 -17963 20950 -17929
rect 20892 -17997 20950 -17963
rect 20892 -18031 20904 -17997
rect 20938 -18031 20950 -17997
rect 20892 -18065 20950 -18031
rect 20892 -18099 20904 -18065
rect 20938 -18099 20950 -18065
rect 20892 -18133 20950 -18099
rect 20892 -18167 20904 -18133
rect 20938 -18167 20950 -18133
rect 20892 -18201 20950 -18167
rect 20892 -18235 20904 -18201
rect 20938 -18235 20950 -18201
rect 20892 -18269 20950 -18235
rect 20892 -18303 20904 -18269
rect 20938 -18303 20950 -18269
rect 20892 -18337 20950 -18303
rect 20892 -18371 20904 -18337
rect 20938 -18371 20950 -18337
rect 20892 -18405 20950 -18371
rect 20892 -18439 20904 -18405
rect 20938 -18439 20950 -18405
rect 20892 -18484 20950 -18439
rect 21910 -17929 21968 -17884
rect 21910 -17963 21922 -17929
rect 21956 -17963 21968 -17929
rect 21910 -17997 21968 -17963
rect 21910 -18031 21922 -17997
rect 21956 -18031 21968 -17997
rect 21910 -18065 21968 -18031
rect 21910 -18099 21922 -18065
rect 21956 -18099 21968 -18065
rect 21910 -18133 21968 -18099
rect 21910 -18167 21922 -18133
rect 21956 -18167 21968 -18133
rect 21910 -18201 21968 -18167
rect 21910 -18235 21922 -18201
rect 21956 -18235 21968 -18201
rect 21910 -18269 21968 -18235
rect 21910 -18303 21922 -18269
rect 21956 -18303 21968 -18269
rect 21910 -18337 21968 -18303
rect 21910 -18371 21922 -18337
rect 21956 -18371 21968 -18337
rect 21910 -18405 21968 -18371
rect 21910 -18439 21922 -18405
rect 21956 -18439 21968 -18405
rect 21910 -18484 21968 -18439
rect 22928 -17929 22986 -17884
rect 22928 -17963 22940 -17929
rect 22974 -17963 22986 -17929
rect 22928 -17997 22986 -17963
rect 22928 -18031 22940 -17997
rect 22974 -18031 22986 -17997
rect 22928 -18065 22986 -18031
rect 22928 -18099 22940 -18065
rect 22974 -18099 22986 -18065
rect 22928 -18133 22986 -18099
rect 22928 -18167 22940 -18133
rect 22974 -18167 22986 -18133
rect 22928 -18201 22986 -18167
rect 22928 -18235 22940 -18201
rect 22974 -18235 22986 -18201
rect 22928 -18269 22986 -18235
rect 22928 -18303 22940 -18269
rect 22974 -18303 22986 -18269
rect 22928 -18337 22986 -18303
rect 22928 -18371 22940 -18337
rect 22974 -18371 22986 -18337
rect 22928 -18405 22986 -18371
rect 22928 -18439 22940 -18405
rect 22974 -18439 22986 -18405
rect 22928 -18484 22986 -18439
rect -34 -18521 -22 -18487
rect 12 -18521 24 -18487
rect -34 -18555 24 -18521
rect -34 -18589 -22 -18555
rect 12 -18589 24 -18555
rect -34 -18623 24 -18589
rect -34 -18657 -22 -18623
rect 12 -18657 24 -18623
rect -34 -18691 24 -18657
rect -34 -18725 -22 -18691
rect 12 -18725 24 -18691
rect -34 -18759 24 -18725
rect -34 -18793 -22 -18759
rect 12 -18793 24 -18759
rect -34 -18838 24 -18793
rect 2568 -19163 2626 -19118
rect 2568 -19197 2580 -19163
rect 2614 -19197 2626 -19163
rect 2568 -19231 2626 -19197
rect 2568 -19265 2580 -19231
rect 2614 -19265 2626 -19231
rect 2568 -19299 2626 -19265
rect 2568 -19333 2580 -19299
rect 2614 -19333 2626 -19299
rect 2568 -19367 2626 -19333
rect 2568 -19401 2580 -19367
rect 2614 -19401 2626 -19367
rect 2568 -19435 2626 -19401
rect 2568 -19469 2580 -19435
rect 2614 -19469 2626 -19435
rect 2568 -19503 2626 -19469
rect 2568 -19537 2580 -19503
rect 2614 -19537 2626 -19503
rect 2568 -19571 2626 -19537
rect 2568 -19605 2580 -19571
rect 2614 -19605 2626 -19571
rect -2336 -19637 -2278 -19622
rect -2336 -19671 -2324 -19637
rect -2290 -19671 -2278 -19637
rect -2336 -19705 -2278 -19671
rect -2336 -19739 -2324 -19705
rect -2290 -19739 -2278 -19705
rect -2336 -19773 -2278 -19739
rect -2336 -19807 -2324 -19773
rect -2290 -19807 -2278 -19773
rect -2336 -19822 -2278 -19807
rect -2118 -19637 -2060 -19622
rect -2118 -19671 -2106 -19637
rect -2072 -19671 -2060 -19637
rect -2118 -19705 -2060 -19671
rect -2118 -19739 -2106 -19705
rect -2072 -19739 -2060 -19705
rect -2118 -19773 -2060 -19739
rect -2118 -19807 -2106 -19773
rect -2072 -19807 -2060 -19773
rect -2118 -19822 -2060 -19807
rect -1900 -19637 -1842 -19622
rect -1900 -19671 -1888 -19637
rect -1854 -19671 -1842 -19637
rect -1900 -19705 -1842 -19671
rect -1900 -19739 -1888 -19705
rect -1854 -19739 -1842 -19705
rect -1900 -19773 -1842 -19739
rect -1900 -19807 -1888 -19773
rect -1854 -19807 -1842 -19773
rect -1900 -19822 -1842 -19807
rect -1682 -19637 -1624 -19622
rect -1682 -19671 -1670 -19637
rect -1636 -19671 -1624 -19637
rect -1682 -19705 -1624 -19671
rect -1682 -19739 -1670 -19705
rect -1636 -19739 -1624 -19705
rect -1682 -19773 -1624 -19739
rect -1682 -19807 -1670 -19773
rect -1636 -19807 -1624 -19773
rect -1682 -19822 -1624 -19807
rect -1464 -19637 -1406 -19622
rect -1464 -19671 -1452 -19637
rect -1418 -19671 -1406 -19637
rect -1464 -19705 -1406 -19671
rect -1464 -19739 -1452 -19705
rect -1418 -19739 -1406 -19705
rect -1464 -19773 -1406 -19739
rect -1464 -19807 -1452 -19773
rect -1418 -19807 -1406 -19773
rect -1464 -19822 -1406 -19807
rect -1246 -19637 -1188 -19622
rect -1246 -19671 -1234 -19637
rect -1200 -19671 -1188 -19637
rect -1246 -19705 -1188 -19671
rect -1246 -19739 -1234 -19705
rect -1200 -19739 -1188 -19705
rect -1246 -19773 -1188 -19739
rect -1246 -19807 -1234 -19773
rect -1200 -19807 -1188 -19773
rect -1246 -19822 -1188 -19807
rect -1028 -19637 -970 -19622
rect -1028 -19671 -1016 -19637
rect -982 -19671 -970 -19637
rect -1028 -19705 -970 -19671
rect -1028 -19739 -1016 -19705
rect -982 -19739 -970 -19705
rect -1028 -19773 -970 -19739
rect -1028 -19807 -1016 -19773
rect -982 -19807 -970 -19773
rect -1028 -19822 -970 -19807
rect -810 -19637 -752 -19622
rect -810 -19671 -798 -19637
rect -764 -19671 -752 -19637
rect -810 -19705 -752 -19671
rect -810 -19739 -798 -19705
rect -764 -19739 -752 -19705
rect -810 -19773 -752 -19739
rect -810 -19807 -798 -19773
rect -764 -19807 -752 -19773
rect -810 -19822 -752 -19807
rect -592 -19637 -534 -19622
rect -592 -19671 -580 -19637
rect -546 -19671 -534 -19637
rect -592 -19705 -534 -19671
rect -592 -19739 -580 -19705
rect -546 -19739 -534 -19705
rect -592 -19773 -534 -19739
rect -592 -19807 -580 -19773
rect -546 -19807 -534 -19773
rect -592 -19822 -534 -19807
rect -374 -19637 -316 -19622
rect -374 -19671 -362 -19637
rect -328 -19671 -316 -19637
rect -374 -19705 -316 -19671
rect -374 -19739 -362 -19705
rect -328 -19739 -316 -19705
rect -374 -19773 -316 -19739
rect -374 -19807 -362 -19773
rect -328 -19807 -316 -19773
rect -374 -19822 -316 -19807
rect -156 -19637 -98 -19622
rect -156 -19671 -144 -19637
rect -110 -19671 -98 -19637
rect -156 -19705 -98 -19671
rect -156 -19739 -144 -19705
rect -110 -19739 -98 -19705
rect 2568 -19639 2626 -19605
rect 2568 -19673 2580 -19639
rect 2614 -19673 2626 -19639
rect 2568 -19718 2626 -19673
rect 3586 -19163 3644 -19118
rect 3586 -19197 3598 -19163
rect 3632 -19197 3644 -19163
rect 3586 -19231 3644 -19197
rect 3586 -19265 3598 -19231
rect 3632 -19265 3644 -19231
rect 3586 -19299 3644 -19265
rect 3586 -19333 3598 -19299
rect 3632 -19333 3644 -19299
rect 3586 -19367 3644 -19333
rect 3586 -19401 3598 -19367
rect 3632 -19401 3644 -19367
rect 3586 -19435 3644 -19401
rect 3586 -19469 3598 -19435
rect 3632 -19469 3644 -19435
rect 3586 -19503 3644 -19469
rect 3586 -19537 3598 -19503
rect 3632 -19537 3644 -19503
rect 3586 -19571 3644 -19537
rect 3586 -19605 3598 -19571
rect 3632 -19605 3644 -19571
rect 3586 -19639 3644 -19605
rect 3586 -19673 3598 -19639
rect 3632 -19673 3644 -19639
rect 3586 -19718 3644 -19673
rect 4604 -19163 4662 -19118
rect 4604 -19197 4616 -19163
rect 4650 -19197 4662 -19163
rect 4604 -19231 4662 -19197
rect 4604 -19265 4616 -19231
rect 4650 -19265 4662 -19231
rect 4604 -19299 4662 -19265
rect 4604 -19333 4616 -19299
rect 4650 -19333 4662 -19299
rect 4604 -19367 4662 -19333
rect 4604 -19401 4616 -19367
rect 4650 -19401 4662 -19367
rect 4604 -19435 4662 -19401
rect 4604 -19469 4616 -19435
rect 4650 -19469 4662 -19435
rect 4604 -19503 4662 -19469
rect 4604 -19537 4616 -19503
rect 4650 -19537 4662 -19503
rect 4604 -19571 4662 -19537
rect 4604 -19605 4616 -19571
rect 4650 -19605 4662 -19571
rect 4604 -19639 4662 -19605
rect 4604 -19673 4616 -19639
rect 4650 -19673 4662 -19639
rect 4604 -19718 4662 -19673
rect 5622 -19163 5680 -19118
rect 5622 -19197 5634 -19163
rect 5668 -19197 5680 -19163
rect 5622 -19231 5680 -19197
rect 5622 -19265 5634 -19231
rect 5668 -19265 5680 -19231
rect 5622 -19299 5680 -19265
rect 5622 -19333 5634 -19299
rect 5668 -19333 5680 -19299
rect 5622 -19367 5680 -19333
rect 5622 -19401 5634 -19367
rect 5668 -19401 5680 -19367
rect 5622 -19435 5680 -19401
rect 5622 -19469 5634 -19435
rect 5668 -19469 5680 -19435
rect 5622 -19503 5680 -19469
rect 5622 -19537 5634 -19503
rect 5668 -19537 5680 -19503
rect 5622 -19571 5680 -19537
rect 5622 -19605 5634 -19571
rect 5668 -19605 5680 -19571
rect 5622 -19639 5680 -19605
rect 5622 -19673 5634 -19639
rect 5668 -19673 5680 -19639
rect 5622 -19718 5680 -19673
rect 6640 -19163 6698 -19118
rect 6640 -19197 6652 -19163
rect 6686 -19197 6698 -19163
rect 6640 -19231 6698 -19197
rect 6640 -19265 6652 -19231
rect 6686 -19265 6698 -19231
rect 6640 -19299 6698 -19265
rect 6640 -19333 6652 -19299
rect 6686 -19333 6698 -19299
rect 6640 -19367 6698 -19333
rect 6640 -19401 6652 -19367
rect 6686 -19401 6698 -19367
rect 6640 -19435 6698 -19401
rect 6640 -19469 6652 -19435
rect 6686 -19469 6698 -19435
rect 6640 -19503 6698 -19469
rect 6640 -19537 6652 -19503
rect 6686 -19537 6698 -19503
rect 6640 -19571 6698 -19537
rect 6640 -19605 6652 -19571
rect 6686 -19605 6698 -19571
rect 6640 -19639 6698 -19605
rect 6640 -19673 6652 -19639
rect 6686 -19673 6698 -19639
rect 6640 -19718 6698 -19673
rect 7658 -19163 7716 -19118
rect 7658 -19197 7670 -19163
rect 7704 -19197 7716 -19163
rect 7658 -19231 7716 -19197
rect 7658 -19265 7670 -19231
rect 7704 -19265 7716 -19231
rect 7658 -19299 7716 -19265
rect 7658 -19333 7670 -19299
rect 7704 -19333 7716 -19299
rect 7658 -19367 7716 -19333
rect 7658 -19401 7670 -19367
rect 7704 -19401 7716 -19367
rect 7658 -19435 7716 -19401
rect 7658 -19469 7670 -19435
rect 7704 -19469 7716 -19435
rect 7658 -19503 7716 -19469
rect 7658 -19537 7670 -19503
rect 7704 -19537 7716 -19503
rect 7658 -19571 7716 -19537
rect 7658 -19605 7670 -19571
rect 7704 -19605 7716 -19571
rect 7658 -19639 7716 -19605
rect 7658 -19673 7670 -19639
rect 7704 -19673 7716 -19639
rect 7658 -19718 7716 -19673
rect 8676 -19163 8734 -19118
rect 8676 -19197 8688 -19163
rect 8722 -19197 8734 -19163
rect 8676 -19231 8734 -19197
rect 8676 -19265 8688 -19231
rect 8722 -19265 8734 -19231
rect 8676 -19299 8734 -19265
rect 8676 -19333 8688 -19299
rect 8722 -19333 8734 -19299
rect 8676 -19367 8734 -19333
rect 8676 -19401 8688 -19367
rect 8722 -19401 8734 -19367
rect 8676 -19435 8734 -19401
rect 8676 -19469 8688 -19435
rect 8722 -19469 8734 -19435
rect 8676 -19503 8734 -19469
rect 8676 -19537 8688 -19503
rect 8722 -19537 8734 -19503
rect 8676 -19571 8734 -19537
rect 8676 -19605 8688 -19571
rect 8722 -19605 8734 -19571
rect 8676 -19639 8734 -19605
rect 8676 -19673 8688 -19639
rect 8722 -19673 8734 -19639
rect 8676 -19718 8734 -19673
rect 9694 -19163 9752 -19118
rect 9694 -19197 9706 -19163
rect 9740 -19197 9752 -19163
rect 9694 -19231 9752 -19197
rect 9694 -19265 9706 -19231
rect 9740 -19265 9752 -19231
rect 9694 -19299 9752 -19265
rect 9694 -19333 9706 -19299
rect 9740 -19333 9752 -19299
rect 9694 -19367 9752 -19333
rect 9694 -19401 9706 -19367
rect 9740 -19401 9752 -19367
rect 9694 -19435 9752 -19401
rect 9694 -19469 9706 -19435
rect 9740 -19469 9752 -19435
rect 9694 -19503 9752 -19469
rect 9694 -19537 9706 -19503
rect 9740 -19537 9752 -19503
rect 9694 -19571 9752 -19537
rect 9694 -19605 9706 -19571
rect 9740 -19605 9752 -19571
rect 9694 -19639 9752 -19605
rect 9694 -19673 9706 -19639
rect 9740 -19673 9752 -19639
rect 9694 -19718 9752 -19673
rect 10712 -19163 10770 -19118
rect 10712 -19197 10724 -19163
rect 10758 -19197 10770 -19163
rect 10712 -19231 10770 -19197
rect 10712 -19265 10724 -19231
rect 10758 -19265 10770 -19231
rect 10712 -19299 10770 -19265
rect 10712 -19333 10724 -19299
rect 10758 -19333 10770 -19299
rect 10712 -19367 10770 -19333
rect 10712 -19401 10724 -19367
rect 10758 -19401 10770 -19367
rect 10712 -19435 10770 -19401
rect 10712 -19469 10724 -19435
rect 10758 -19469 10770 -19435
rect 10712 -19503 10770 -19469
rect 10712 -19537 10724 -19503
rect 10758 -19537 10770 -19503
rect 10712 -19571 10770 -19537
rect 10712 -19605 10724 -19571
rect 10758 -19605 10770 -19571
rect 10712 -19639 10770 -19605
rect 10712 -19673 10724 -19639
rect 10758 -19673 10770 -19639
rect 10712 -19718 10770 -19673
rect 11730 -19163 11788 -19118
rect 11730 -19197 11742 -19163
rect 11776 -19197 11788 -19163
rect 11730 -19231 11788 -19197
rect 11730 -19265 11742 -19231
rect 11776 -19265 11788 -19231
rect 11730 -19299 11788 -19265
rect 11730 -19333 11742 -19299
rect 11776 -19333 11788 -19299
rect 11730 -19367 11788 -19333
rect 11730 -19401 11742 -19367
rect 11776 -19401 11788 -19367
rect 11730 -19435 11788 -19401
rect 11730 -19469 11742 -19435
rect 11776 -19469 11788 -19435
rect 11730 -19503 11788 -19469
rect 11730 -19537 11742 -19503
rect 11776 -19537 11788 -19503
rect 11730 -19571 11788 -19537
rect 11730 -19605 11742 -19571
rect 11776 -19605 11788 -19571
rect 11730 -19639 11788 -19605
rect 11730 -19673 11742 -19639
rect 11776 -19673 11788 -19639
rect 11730 -19718 11788 -19673
rect 12748 -19163 12806 -19118
rect 12748 -19197 12760 -19163
rect 12794 -19197 12806 -19163
rect 12748 -19231 12806 -19197
rect 12748 -19265 12760 -19231
rect 12794 -19265 12806 -19231
rect 12748 -19299 12806 -19265
rect 12748 -19333 12760 -19299
rect 12794 -19333 12806 -19299
rect 12748 -19367 12806 -19333
rect 12748 -19401 12760 -19367
rect 12794 -19401 12806 -19367
rect 12748 -19435 12806 -19401
rect 12748 -19469 12760 -19435
rect 12794 -19469 12806 -19435
rect 12748 -19503 12806 -19469
rect 12748 -19537 12760 -19503
rect 12794 -19537 12806 -19503
rect 12748 -19571 12806 -19537
rect 12748 -19605 12760 -19571
rect 12794 -19605 12806 -19571
rect 12748 -19639 12806 -19605
rect 12748 -19673 12760 -19639
rect 12794 -19673 12806 -19639
rect 12748 -19718 12806 -19673
rect 13766 -19163 13824 -19118
rect 13766 -19197 13778 -19163
rect 13812 -19197 13824 -19163
rect 13766 -19231 13824 -19197
rect 13766 -19265 13778 -19231
rect 13812 -19265 13824 -19231
rect 13766 -19299 13824 -19265
rect 13766 -19333 13778 -19299
rect 13812 -19333 13824 -19299
rect 13766 -19367 13824 -19333
rect 13766 -19401 13778 -19367
rect 13812 -19401 13824 -19367
rect 13766 -19435 13824 -19401
rect 13766 -19469 13778 -19435
rect 13812 -19469 13824 -19435
rect 13766 -19503 13824 -19469
rect 13766 -19537 13778 -19503
rect 13812 -19537 13824 -19503
rect 13766 -19571 13824 -19537
rect 13766 -19605 13778 -19571
rect 13812 -19605 13824 -19571
rect 13766 -19639 13824 -19605
rect 13766 -19673 13778 -19639
rect 13812 -19673 13824 -19639
rect 13766 -19718 13824 -19673
rect 14784 -19163 14842 -19118
rect 14784 -19197 14796 -19163
rect 14830 -19197 14842 -19163
rect 14784 -19231 14842 -19197
rect 14784 -19265 14796 -19231
rect 14830 -19265 14842 -19231
rect 14784 -19299 14842 -19265
rect 14784 -19333 14796 -19299
rect 14830 -19333 14842 -19299
rect 14784 -19367 14842 -19333
rect 14784 -19401 14796 -19367
rect 14830 -19401 14842 -19367
rect 14784 -19435 14842 -19401
rect 14784 -19469 14796 -19435
rect 14830 -19469 14842 -19435
rect 14784 -19503 14842 -19469
rect 14784 -19537 14796 -19503
rect 14830 -19537 14842 -19503
rect 14784 -19571 14842 -19537
rect 14784 -19605 14796 -19571
rect 14830 -19605 14842 -19571
rect 14784 -19639 14842 -19605
rect 14784 -19673 14796 -19639
rect 14830 -19673 14842 -19639
rect 14784 -19718 14842 -19673
rect 15802 -19163 15860 -19118
rect 15802 -19197 15814 -19163
rect 15848 -19197 15860 -19163
rect 15802 -19231 15860 -19197
rect 15802 -19265 15814 -19231
rect 15848 -19265 15860 -19231
rect 15802 -19299 15860 -19265
rect 15802 -19333 15814 -19299
rect 15848 -19333 15860 -19299
rect 15802 -19367 15860 -19333
rect 15802 -19401 15814 -19367
rect 15848 -19401 15860 -19367
rect 15802 -19435 15860 -19401
rect 15802 -19469 15814 -19435
rect 15848 -19469 15860 -19435
rect 15802 -19503 15860 -19469
rect 15802 -19537 15814 -19503
rect 15848 -19537 15860 -19503
rect 15802 -19571 15860 -19537
rect 15802 -19605 15814 -19571
rect 15848 -19605 15860 -19571
rect 15802 -19639 15860 -19605
rect 15802 -19673 15814 -19639
rect 15848 -19673 15860 -19639
rect 15802 -19718 15860 -19673
rect 16820 -19163 16878 -19118
rect 16820 -19197 16832 -19163
rect 16866 -19197 16878 -19163
rect 16820 -19231 16878 -19197
rect 16820 -19265 16832 -19231
rect 16866 -19265 16878 -19231
rect 16820 -19299 16878 -19265
rect 16820 -19333 16832 -19299
rect 16866 -19333 16878 -19299
rect 16820 -19367 16878 -19333
rect 16820 -19401 16832 -19367
rect 16866 -19401 16878 -19367
rect 16820 -19435 16878 -19401
rect 16820 -19469 16832 -19435
rect 16866 -19469 16878 -19435
rect 16820 -19503 16878 -19469
rect 16820 -19537 16832 -19503
rect 16866 -19537 16878 -19503
rect 16820 -19571 16878 -19537
rect 16820 -19605 16832 -19571
rect 16866 -19605 16878 -19571
rect 16820 -19639 16878 -19605
rect 16820 -19673 16832 -19639
rect 16866 -19673 16878 -19639
rect 16820 -19718 16878 -19673
rect 17838 -19163 17896 -19118
rect 17838 -19197 17850 -19163
rect 17884 -19197 17896 -19163
rect 17838 -19231 17896 -19197
rect 17838 -19265 17850 -19231
rect 17884 -19265 17896 -19231
rect 17838 -19299 17896 -19265
rect 17838 -19333 17850 -19299
rect 17884 -19333 17896 -19299
rect 17838 -19367 17896 -19333
rect 17838 -19401 17850 -19367
rect 17884 -19401 17896 -19367
rect 17838 -19435 17896 -19401
rect 17838 -19469 17850 -19435
rect 17884 -19469 17896 -19435
rect 17838 -19503 17896 -19469
rect 17838 -19537 17850 -19503
rect 17884 -19537 17896 -19503
rect 17838 -19571 17896 -19537
rect 17838 -19605 17850 -19571
rect 17884 -19605 17896 -19571
rect 17838 -19639 17896 -19605
rect 17838 -19673 17850 -19639
rect 17884 -19673 17896 -19639
rect 17838 -19718 17896 -19673
rect 18856 -19163 18914 -19118
rect 18856 -19197 18868 -19163
rect 18902 -19197 18914 -19163
rect 18856 -19231 18914 -19197
rect 18856 -19265 18868 -19231
rect 18902 -19265 18914 -19231
rect 18856 -19299 18914 -19265
rect 18856 -19333 18868 -19299
rect 18902 -19333 18914 -19299
rect 18856 -19367 18914 -19333
rect 18856 -19401 18868 -19367
rect 18902 -19401 18914 -19367
rect 18856 -19435 18914 -19401
rect 18856 -19469 18868 -19435
rect 18902 -19469 18914 -19435
rect 18856 -19503 18914 -19469
rect 18856 -19537 18868 -19503
rect 18902 -19537 18914 -19503
rect 18856 -19571 18914 -19537
rect 18856 -19605 18868 -19571
rect 18902 -19605 18914 -19571
rect 18856 -19639 18914 -19605
rect 18856 -19673 18868 -19639
rect 18902 -19673 18914 -19639
rect 18856 -19718 18914 -19673
rect 19874 -19163 19932 -19118
rect 19874 -19197 19886 -19163
rect 19920 -19197 19932 -19163
rect 19874 -19231 19932 -19197
rect 19874 -19265 19886 -19231
rect 19920 -19265 19932 -19231
rect 19874 -19299 19932 -19265
rect 19874 -19333 19886 -19299
rect 19920 -19333 19932 -19299
rect 19874 -19367 19932 -19333
rect 19874 -19401 19886 -19367
rect 19920 -19401 19932 -19367
rect 19874 -19435 19932 -19401
rect 19874 -19469 19886 -19435
rect 19920 -19469 19932 -19435
rect 19874 -19503 19932 -19469
rect 19874 -19537 19886 -19503
rect 19920 -19537 19932 -19503
rect 19874 -19571 19932 -19537
rect 19874 -19605 19886 -19571
rect 19920 -19605 19932 -19571
rect 19874 -19639 19932 -19605
rect 19874 -19673 19886 -19639
rect 19920 -19673 19932 -19639
rect 19874 -19718 19932 -19673
rect 20892 -19163 20950 -19118
rect 20892 -19197 20904 -19163
rect 20938 -19197 20950 -19163
rect 20892 -19231 20950 -19197
rect 20892 -19265 20904 -19231
rect 20938 -19265 20950 -19231
rect 20892 -19299 20950 -19265
rect 20892 -19333 20904 -19299
rect 20938 -19333 20950 -19299
rect 20892 -19367 20950 -19333
rect 20892 -19401 20904 -19367
rect 20938 -19401 20950 -19367
rect 20892 -19435 20950 -19401
rect 20892 -19469 20904 -19435
rect 20938 -19469 20950 -19435
rect 20892 -19503 20950 -19469
rect 20892 -19537 20904 -19503
rect 20938 -19537 20950 -19503
rect 20892 -19571 20950 -19537
rect 20892 -19605 20904 -19571
rect 20938 -19605 20950 -19571
rect 20892 -19639 20950 -19605
rect 20892 -19673 20904 -19639
rect 20938 -19673 20950 -19639
rect 20892 -19718 20950 -19673
rect 21910 -19163 21968 -19118
rect 21910 -19197 21922 -19163
rect 21956 -19197 21968 -19163
rect 21910 -19231 21968 -19197
rect 21910 -19265 21922 -19231
rect 21956 -19265 21968 -19231
rect 21910 -19299 21968 -19265
rect 21910 -19333 21922 -19299
rect 21956 -19333 21968 -19299
rect 21910 -19367 21968 -19333
rect 21910 -19401 21922 -19367
rect 21956 -19401 21968 -19367
rect 21910 -19435 21968 -19401
rect 21910 -19469 21922 -19435
rect 21956 -19469 21968 -19435
rect 21910 -19503 21968 -19469
rect 21910 -19537 21922 -19503
rect 21956 -19537 21968 -19503
rect 21910 -19571 21968 -19537
rect 21910 -19605 21922 -19571
rect 21956 -19605 21968 -19571
rect 21910 -19639 21968 -19605
rect 21910 -19673 21922 -19639
rect 21956 -19673 21968 -19639
rect 21910 -19718 21968 -19673
rect 22928 -19163 22986 -19118
rect 22928 -19197 22940 -19163
rect 22974 -19197 22986 -19163
rect 22928 -19231 22986 -19197
rect 22928 -19265 22940 -19231
rect 22974 -19265 22986 -19231
rect 22928 -19299 22986 -19265
rect 22928 -19333 22940 -19299
rect 22974 -19333 22986 -19299
rect 22928 -19367 22986 -19333
rect 22928 -19401 22940 -19367
rect 22974 -19401 22986 -19367
rect 22928 -19435 22986 -19401
rect 22928 -19469 22940 -19435
rect 22974 -19469 22986 -19435
rect 22928 -19503 22986 -19469
rect 22928 -19537 22940 -19503
rect 22974 -19537 22986 -19503
rect 22928 -19571 22986 -19537
rect 22928 -19605 22940 -19571
rect 22974 -19605 22986 -19571
rect 22928 -19639 22986 -19605
rect 22928 -19673 22940 -19639
rect 22974 -19673 22986 -19639
rect 22928 -19718 22986 -19673
rect -156 -19773 -98 -19739
rect -156 -19807 -144 -19773
rect -110 -19807 -98 -19773
rect -156 -19822 -98 -19807
rect 2568 -20397 2626 -20352
rect 2568 -20431 2580 -20397
rect 2614 -20431 2626 -20397
rect -2336 -20469 -2278 -20454
rect -2336 -20503 -2324 -20469
rect -2290 -20503 -2278 -20469
rect -2336 -20537 -2278 -20503
rect -2336 -20571 -2324 -20537
rect -2290 -20571 -2278 -20537
rect -2336 -20605 -2278 -20571
rect -2336 -20639 -2324 -20605
rect -2290 -20639 -2278 -20605
rect -2336 -20654 -2278 -20639
rect -2118 -20469 -2060 -20454
rect -2118 -20503 -2106 -20469
rect -2072 -20503 -2060 -20469
rect -2118 -20537 -2060 -20503
rect -2118 -20571 -2106 -20537
rect -2072 -20571 -2060 -20537
rect -2118 -20605 -2060 -20571
rect -2118 -20639 -2106 -20605
rect -2072 -20639 -2060 -20605
rect -2118 -20654 -2060 -20639
rect -1900 -20469 -1842 -20454
rect -1900 -20503 -1888 -20469
rect -1854 -20503 -1842 -20469
rect -1900 -20537 -1842 -20503
rect -1900 -20571 -1888 -20537
rect -1854 -20571 -1842 -20537
rect -1900 -20605 -1842 -20571
rect -1900 -20639 -1888 -20605
rect -1854 -20639 -1842 -20605
rect -1900 -20654 -1842 -20639
rect -1682 -20469 -1624 -20454
rect -1682 -20503 -1670 -20469
rect -1636 -20503 -1624 -20469
rect -1682 -20537 -1624 -20503
rect -1682 -20571 -1670 -20537
rect -1636 -20571 -1624 -20537
rect -1682 -20605 -1624 -20571
rect -1682 -20639 -1670 -20605
rect -1636 -20639 -1624 -20605
rect -1682 -20654 -1624 -20639
rect -1464 -20469 -1406 -20454
rect -1464 -20503 -1452 -20469
rect -1418 -20503 -1406 -20469
rect -1464 -20537 -1406 -20503
rect -1464 -20571 -1452 -20537
rect -1418 -20571 -1406 -20537
rect -1464 -20605 -1406 -20571
rect -1464 -20639 -1452 -20605
rect -1418 -20639 -1406 -20605
rect -1464 -20654 -1406 -20639
rect -1246 -20469 -1188 -20454
rect -1246 -20503 -1234 -20469
rect -1200 -20503 -1188 -20469
rect -1246 -20537 -1188 -20503
rect -1246 -20571 -1234 -20537
rect -1200 -20571 -1188 -20537
rect -1246 -20605 -1188 -20571
rect -1246 -20639 -1234 -20605
rect -1200 -20639 -1188 -20605
rect -1246 -20654 -1188 -20639
rect -1028 -20469 -970 -20454
rect -1028 -20503 -1016 -20469
rect -982 -20503 -970 -20469
rect -1028 -20537 -970 -20503
rect -1028 -20571 -1016 -20537
rect -982 -20571 -970 -20537
rect -1028 -20605 -970 -20571
rect -1028 -20639 -1016 -20605
rect -982 -20639 -970 -20605
rect -1028 -20654 -970 -20639
rect -810 -20469 -752 -20454
rect -810 -20503 -798 -20469
rect -764 -20503 -752 -20469
rect -810 -20537 -752 -20503
rect -810 -20571 -798 -20537
rect -764 -20571 -752 -20537
rect -810 -20605 -752 -20571
rect -810 -20639 -798 -20605
rect -764 -20639 -752 -20605
rect -810 -20654 -752 -20639
rect -592 -20469 -534 -20454
rect -592 -20503 -580 -20469
rect -546 -20503 -534 -20469
rect -592 -20537 -534 -20503
rect -592 -20571 -580 -20537
rect -546 -20571 -534 -20537
rect -592 -20605 -534 -20571
rect -592 -20639 -580 -20605
rect -546 -20639 -534 -20605
rect -592 -20654 -534 -20639
rect -374 -20469 -316 -20454
rect -374 -20503 -362 -20469
rect -328 -20503 -316 -20469
rect -374 -20537 -316 -20503
rect -374 -20571 -362 -20537
rect -328 -20571 -316 -20537
rect -374 -20605 -316 -20571
rect -374 -20639 -362 -20605
rect -328 -20639 -316 -20605
rect -374 -20654 -316 -20639
rect -156 -20469 -98 -20454
rect -156 -20503 -144 -20469
rect -110 -20503 -98 -20469
rect -156 -20537 -98 -20503
rect -156 -20571 -144 -20537
rect -110 -20571 -98 -20537
rect -156 -20605 -98 -20571
rect -156 -20639 -144 -20605
rect -110 -20639 -98 -20605
rect -156 -20654 -98 -20639
rect 2568 -20465 2626 -20431
rect 2568 -20499 2580 -20465
rect 2614 -20499 2626 -20465
rect 2568 -20533 2626 -20499
rect 2568 -20567 2580 -20533
rect 2614 -20567 2626 -20533
rect 2568 -20601 2626 -20567
rect 2568 -20635 2580 -20601
rect 2614 -20635 2626 -20601
rect 2568 -20669 2626 -20635
rect 2568 -20703 2580 -20669
rect 2614 -20703 2626 -20669
rect 2568 -20737 2626 -20703
rect 2568 -20771 2580 -20737
rect 2614 -20771 2626 -20737
rect 2568 -20805 2626 -20771
rect 2568 -20839 2580 -20805
rect 2614 -20839 2626 -20805
rect 2568 -20873 2626 -20839
rect 2568 -20907 2580 -20873
rect 2614 -20907 2626 -20873
rect 2568 -20952 2626 -20907
rect 3586 -20397 3644 -20352
rect 3586 -20431 3598 -20397
rect 3632 -20431 3644 -20397
rect 3586 -20465 3644 -20431
rect 3586 -20499 3598 -20465
rect 3632 -20499 3644 -20465
rect 3586 -20533 3644 -20499
rect 3586 -20567 3598 -20533
rect 3632 -20567 3644 -20533
rect 3586 -20601 3644 -20567
rect 3586 -20635 3598 -20601
rect 3632 -20635 3644 -20601
rect 3586 -20669 3644 -20635
rect 3586 -20703 3598 -20669
rect 3632 -20703 3644 -20669
rect 3586 -20737 3644 -20703
rect 3586 -20771 3598 -20737
rect 3632 -20771 3644 -20737
rect 3586 -20805 3644 -20771
rect 3586 -20839 3598 -20805
rect 3632 -20839 3644 -20805
rect 3586 -20873 3644 -20839
rect 3586 -20907 3598 -20873
rect 3632 -20907 3644 -20873
rect 3586 -20952 3644 -20907
rect 4604 -20397 4662 -20352
rect 4604 -20431 4616 -20397
rect 4650 -20431 4662 -20397
rect 4604 -20465 4662 -20431
rect 4604 -20499 4616 -20465
rect 4650 -20499 4662 -20465
rect 4604 -20533 4662 -20499
rect 4604 -20567 4616 -20533
rect 4650 -20567 4662 -20533
rect 4604 -20601 4662 -20567
rect 4604 -20635 4616 -20601
rect 4650 -20635 4662 -20601
rect 4604 -20669 4662 -20635
rect 4604 -20703 4616 -20669
rect 4650 -20703 4662 -20669
rect 4604 -20737 4662 -20703
rect 4604 -20771 4616 -20737
rect 4650 -20771 4662 -20737
rect 4604 -20805 4662 -20771
rect 4604 -20839 4616 -20805
rect 4650 -20839 4662 -20805
rect 4604 -20873 4662 -20839
rect 4604 -20907 4616 -20873
rect 4650 -20907 4662 -20873
rect 4604 -20952 4662 -20907
rect 5622 -20397 5680 -20352
rect 5622 -20431 5634 -20397
rect 5668 -20431 5680 -20397
rect 5622 -20465 5680 -20431
rect 5622 -20499 5634 -20465
rect 5668 -20499 5680 -20465
rect 5622 -20533 5680 -20499
rect 5622 -20567 5634 -20533
rect 5668 -20567 5680 -20533
rect 5622 -20601 5680 -20567
rect 5622 -20635 5634 -20601
rect 5668 -20635 5680 -20601
rect 5622 -20669 5680 -20635
rect 5622 -20703 5634 -20669
rect 5668 -20703 5680 -20669
rect 5622 -20737 5680 -20703
rect 5622 -20771 5634 -20737
rect 5668 -20771 5680 -20737
rect 5622 -20805 5680 -20771
rect 5622 -20839 5634 -20805
rect 5668 -20839 5680 -20805
rect 5622 -20873 5680 -20839
rect 5622 -20907 5634 -20873
rect 5668 -20907 5680 -20873
rect 5622 -20952 5680 -20907
rect 6640 -20397 6698 -20352
rect 6640 -20431 6652 -20397
rect 6686 -20431 6698 -20397
rect 6640 -20465 6698 -20431
rect 6640 -20499 6652 -20465
rect 6686 -20499 6698 -20465
rect 6640 -20533 6698 -20499
rect 6640 -20567 6652 -20533
rect 6686 -20567 6698 -20533
rect 6640 -20601 6698 -20567
rect 6640 -20635 6652 -20601
rect 6686 -20635 6698 -20601
rect 6640 -20669 6698 -20635
rect 6640 -20703 6652 -20669
rect 6686 -20703 6698 -20669
rect 6640 -20737 6698 -20703
rect 6640 -20771 6652 -20737
rect 6686 -20771 6698 -20737
rect 6640 -20805 6698 -20771
rect 6640 -20839 6652 -20805
rect 6686 -20839 6698 -20805
rect 6640 -20873 6698 -20839
rect 6640 -20907 6652 -20873
rect 6686 -20907 6698 -20873
rect 6640 -20952 6698 -20907
rect 7658 -20397 7716 -20352
rect 7658 -20431 7670 -20397
rect 7704 -20431 7716 -20397
rect 7658 -20465 7716 -20431
rect 7658 -20499 7670 -20465
rect 7704 -20499 7716 -20465
rect 7658 -20533 7716 -20499
rect 7658 -20567 7670 -20533
rect 7704 -20567 7716 -20533
rect 7658 -20601 7716 -20567
rect 7658 -20635 7670 -20601
rect 7704 -20635 7716 -20601
rect 7658 -20669 7716 -20635
rect 7658 -20703 7670 -20669
rect 7704 -20703 7716 -20669
rect 7658 -20737 7716 -20703
rect 7658 -20771 7670 -20737
rect 7704 -20771 7716 -20737
rect 7658 -20805 7716 -20771
rect 7658 -20839 7670 -20805
rect 7704 -20839 7716 -20805
rect 7658 -20873 7716 -20839
rect 7658 -20907 7670 -20873
rect 7704 -20907 7716 -20873
rect 7658 -20952 7716 -20907
rect 8676 -20397 8734 -20352
rect 8676 -20431 8688 -20397
rect 8722 -20431 8734 -20397
rect 8676 -20465 8734 -20431
rect 8676 -20499 8688 -20465
rect 8722 -20499 8734 -20465
rect 8676 -20533 8734 -20499
rect 8676 -20567 8688 -20533
rect 8722 -20567 8734 -20533
rect 8676 -20601 8734 -20567
rect 8676 -20635 8688 -20601
rect 8722 -20635 8734 -20601
rect 8676 -20669 8734 -20635
rect 8676 -20703 8688 -20669
rect 8722 -20703 8734 -20669
rect 8676 -20737 8734 -20703
rect 8676 -20771 8688 -20737
rect 8722 -20771 8734 -20737
rect 8676 -20805 8734 -20771
rect 8676 -20839 8688 -20805
rect 8722 -20839 8734 -20805
rect 8676 -20873 8734 -20839
rect 8676 -20907 8688 -20873
rect 8722 -20907 8734 -20873
rect 8676 -20952 8734 -20907
rect 9694 -20397 9752 -20352
rect 9694 -20431 9706 -20397
rect 9740 -20431 9752 -20397
rect 9694 -20465 9752 -20431
rect 9694 -20499 9706 -20465
rect 9740 -20499 9752 -20465
rect 9694 -20533 9752 -20499
rect 9694 -20567 9706 -20533
rect 9740 -20567 9752 -20533
rect 9694 -20601 9752 -20567
rect 9694 -20635 9706 -20601
rect 9740 -20635 9752 -20601
rect 9694 -20669 9752 -20635
rect 9694 -20703 9706 -20669
rect 9740 -20703 9752 -20669
rect 9694 -20737 9752 -20703
rect 9694 -20771 9706 -20737
rect 9740 -20771 9752 -20737
rect 9694 -20805 9752 -20771
rect 9694 -20839 9706 -20805
rect 9740 -20839 9752 -20805
rect 9694 -20873 9752 -20839
rect 9694 -20907 9706 -20873
rect 9740 -20907 9752 -20873
rect 9694 -20952 9752 -20907
rect 10712 -20397 10770 -20352
rect 10712 -20431 10724 -20397
rect 10758 -20431 10770 -20397
rect 10712 -20465 10770 -20431
rect 10712 -20499 10724 -20465
rect 10758 -20499 10770 -20465
rect 10712 -20533 10770 -20499
rect 10712 -20567 10724 -20533
rect 10758 -20567 10770 -20533
rect 10712 -20601 10770 -20567
rect 10712 -20635 10724 -20601
rect 10758 -20635 10770 -20601
rect 10712 -20669 10770 -20635
rect 10712 -20703 10724 -20669
rect 10758 -20703 10770 -20669
rect 10712 -20737 10770 -20703
rect 10712 -20771 10724 -20737
rect 10758 -20771 10770 -20737
rect 10712 -20805 10770 -20771
rect 10712 -20839 10724 -20805
rect 10758 -20839 10770 -20805
rect 10712 -20873 10770 -20839
rect 10712 -20907 10724 -20873
rect 10758 -20907 10770 -20873
rect 10712 -20952 10770 -20907
rect 11730 -20397 11788 -20352
rect 11730 -20431 11742 -20397
rect 11776 -20431 11788 -20397
rect 11730 -20465 11788 -20431
rect 11730 -20499 11742 -20465
rect 11776 -20499 11788 -20465
rect 11730 -20533 11788 -20499
rect 11730 -20567 11742 -20533
rect 11776 -20567 11788 -20533
rect 11730 -20601 11788 -20567
rect 11730 -20635 11742 -20601
rect 11776 -20635 11788 -20601
rect 11730 -20669 11788 -20635
rect 11730 -20703 11742 -20669
rect 11776 -20703 11788 -20669
rect 11730 -20737 11788 -20703
rect 11730 -20771 11742 -20737
rect 11776 -20771 11788 -20737
rect 11730 -20805 11788 -20771
rect 11730 -20839 11742 -20805
rect 11776 -20839 11788 -20805
rect 11730 -20873 11788 -20839
rect 11730 -20907 11742 -20873
rect 11776 -20907 11788 -20873
rect 11730 -20952 11788 -20907
rect 12748 -20397 12806 -20352
rect 12748 -20431 12760 -20397
rect 12794 -20431 12806 -20397
rect 12748 -20465 12806 -20431
rect 12748 -20499 12760 -20465
rect 12794 -20499 12806 -20465
rect 12748 -20533 12806 -20499
rect 12748 -20567 12760 -20533
rect 12794 -20567 12806 -20533
rect 12748 -20601 12806 -20567
rect 12748 -20635 12760 -20601
rect 12794 -20635 12806 -20601
rect 12748 -20669 12806 -20635
rect 12748 -20703 12760 -20669
rect 12794 -20703 12806 -20669
rect 12748 -20737 12806 -20703
rect 12748 -20771 12760 -20737
rect 12794 -20771 12806 -20737
rect 12748 -20805 12806 -20771
rect 12748 -20839 12760 -20805
rect 12794 -20839 12806 -20805
rect 12748 -20873 12806 -20839
rect 12748 -20907 12760 -20873
rect 12794 -20907 12806 -20873
rect 12748 -20952 12806 -20907
rect 13766 -20397 13824 -20352
rect 13766 -20431 13778 -20397
rect 13812 -20431 13824 -20397
rect 13766 -20465 13824 -20431
rect 13766 -20499 13778 -20465
rect 13812 -20499 13824 -20465
rect 13766 -20533 13824 -20499
rect 13766 -20567 13778 -20533
rect 13812 -20567 13824 -20533
rect 13766 -20601 13824 -20567
rect 13766 -20635 13778 -20601
rect 13812 -20635 13824 -20601
rect 13766 -20669 13824 -20635
rect 13766 -20703 13778 -20669
rect 13812 -20703 13824 -20669
rect 13766 -20737 13824 -20703
rect 13766 -20771 13778 -20737
rect 13812 -20771 13824 -20737
rect 13766 -20805 13824 -20771
rect 13766 -20839 13778 -20805
rect 13812 -20839 13824 -20805
rect 13766 -20873 13824 -20839
rect 13766 -20907 13778 -20873
rect 13812 -20907 13824 -20873
rect 13766 -20952 13824 -20907
rect 14784 -20397 14842 -20352
rect 14784 -20431 14796 -20397
rect 14830 -20431 14842 -20397
rect 14784 -20465 14842 -20431
rect 14784 -20499 14796 -20465
rect 14830 -20499 14842 -20465
rect 14784 -20533 14842 -20499
rect 14784 -20567 14796 -20533
rect 14830 -20567 14842 -20533
rect 14784 -20601 14842 -20567
rect 14784 -20635 14796 -20601
rect 14830 -20635 14842 -20601
rect 14784 -20669 14842 -20635
rect 14784 -20703 14796 -20669
rect 14830 -20703 14842 -20669
rect 14784 -20737 14842 -20703
rect 14784 -20771 14796 -20737
rect 14830 -20771 14842 -20737
rect 14784 -20805 14842 -20771
rect 14784 -20839 14796 -20805
rect 14830 -20839 14842 -20805
rect 14784 -20873 14842 -20839
rect 14784 -20907 14796 -20873
rect 14830 -20907 14842 -20873
rect 14784 -20952 14842 -20907
rect 15802 -20397 15860 -20352
rect 15802 -20431 15814 -20397
rect 15848 -20431 15860 -20397
rect 15802 -20465 15860 -20431
rect 15802 -20499 15814 -20465
rect 15848 -20499 15860 -20465
rect 15802 -20533 15860 -20499
rect 15802 -20567 15814 -20533
rect 15848 -20567 15860 -20533
rect 15802 -20601 15860 -20567
rect 15802 -20635 15814 -20601
rect 15848 -20635 15860 -20601
rect 15802 -20669 15860 -20635
rect 15802 -20703 15814 -20669
rect 15848 -20703 15860 -20669
rect 15802 -20737 15860 -20703
rect 15802 -20771 15814 -20737
rect 15848 -20771 15860 -20737
rect 15802 -20805 15860 -20771
rect 15802 -20839 15814 -20805
rect 15848 -20839 15860 -20805
rect 15802 -20873 15860 -20839
rect 15802 -20907 15814 -20873
rect 15848 -20907 15860 -20873
rect 15802 -20952 15860 -20907
rect 16820 -20397 16878 -20352
rect 16820 -20431 16832 -20397
rect 16866 -20431 16878 -20397
rect 16820 -20465 16878 -20431
rect 16820 -20499 16832 -20465
rect 16866 -20499 16878 -20465
rect 16820 -20533 16878 -20499
rect 16820 -20567 16832 -20533
rect 16866 -20567 16878 -20533
rect 16820 -20601 16878 -20567
rect 16820 -20635 16832 -20601
rect 16866 -20635 16878 -20601
rect 16820 -20669 16878 -20635
rect 16820 -20703 16832 -20669
rect 16866 -20703 16878 -20669
rect 16820 -20737 16878 -20703
rect 16820 -20771 16832 -20737
rect 16866 -20771 16878 -20737
rect 16820 -20805 16878 -20771
rect 16820 -20839 16832 -20805
rect 16866 -20839 16878 -20805
rect 16820 -20873 16878 -20839
rect 16820 -20907 16832 -20873
rect 16866 -20907 16878 -20873
rect 16820 -20952 16878 -20907
rect 17838 -20397 17896 -20352
rect 17838 -20431 17850 -20397
rect 17884 -20431 17896 -20397
rect 17838 -20465 17896 -20431
rect 17838 -20499 17850 -20465
rect 17884 -20499 17896 -20465
rect 17838 -20533 17896 -20499
rect 17838 -20567 17850 -20533
rect 17884 -20567 17896 -20533
rect 17838 -20601 17896 -20567
rect 17838 -20635 17850 -20601
rect 17884 -20635 17896 -20601
rect 17838 -20669 17896 -20635
rect 17838 -20703 17850 -20669
rect 17884 -20703 17896 -20669
rect 17838 -20737 17896 -20703
rect 17838 -20771 17850 -20737
rect 17884 -20771 17896 -20737
rect 17838 -20805 17896 -20771
rect 17838 -20839 17850 -20805
rect 17884 -20839 17896 -20805
rect 17838 -20873 17896 -20839
rect 17838 -20907 17850 -20873
rect 17884 -20907 17896 -20873
rect 17838 -20952 17896 -20907
rect 18856 -20397 18914 -20352
rect 18856 -20431 18868 -20397
rect 18902 -20431 18914 -20397
rect 18856 -20465 18914 -20431
rect 18856 -20499 18868 -20465
rect 18902 -20499 18914 -20465
rect 18856 -20533 18914 -20499
rect 18856 -20567 18868 -20533
rect 18902 -20567 18914 -20533
rect 18856 -20601 18914 -20567
rect 18856 -20635 18868 -20601
rect 18902 -20635 18914 -20601
rect 18856 -20669 18914 -20635
rect 18856 -20703 18868 -20669
rect 18902 -20703 18914 -20669
rect 18856 -20737 18914 -20703
rect 18856 -20771 18868 -20737
rect 18902 -20771 18914 -20737
rect 18856 -20805 18914 -20771
rect 18856 -20839 18868 -20805
rect 18902 -20839 18914 -20805
rect 18856 -20873 18914 -20839
rect 18856 -20907 18868 -20873
rect 18902 -20907 18914 -20873
rect 18856 -20952 18914 -20907
rect 19874 -20397 19932 -20352
rect 19874 -20431 19886 -20397
rect 19920 -20431 19932 -20397
rect 19874 -20465 19932 -20431
rect 19874 -20499 19886 -20465
rect 19920 -20499 19932 -20465
rect 19874 -20533 19932 -20499
rect 19874 -20567 19886 -20533
rect 19920 -20567 19932 -20533
rect 19874 -20601 19932 -20567
rect 19874 -20635 19886 -20601
rect 19920 -20635 19932 -20601
rect 19874 -20669 19932 -20635
rect 19874 -20703 19886 -20669
rect 19920 -20703 19932 -20669
rect 19874 -20737 19932 -20703
rect 19874 -20771 19886 -20737
rect 19920 -20771 19932 -20737
rect 19874 -20805 19932 -20771
rect 19874 -20839 19886 -20805
rect 19920 -20839 19932 -20805
rect 19874 -20873 19932 -20839
rect 19874 -20907 19886 -20873
rect 19920 -20907 19932 -20873
rect 19874 -20952 19932 -20907
rect 20892 -20397 20950 -20352
rect 20892 -20431 20904 -20397
rect 20938 -20431 20950 -20397
rect 20892 -20465 20950 -20431
rect 20892 -20499 20904 -20465
rect 20938 -20499 20950 -20465
rect 20892 -20533 20950 -20499
rect 20892 -20567 20904 -20533
rect 20938 -20567 20950 -20533
rect 20892 -20601 20950 -20567
rect 20892 -20635 20904 -20601
rect 20938 -20635 20950 -20601
rect 20892 -20669 20950 -20635
rect 20892 -20703 20904 -20669
rect 20938 -20703 20950 -20669
rect 20892 -20737 20950 -20703
rect 20892 -20771 20904 -20737
rect 20938 -20771 20950 -20737
rect 20892 -20805 20950 -20771
rect 20892 -20839 20904 -20805
rect 20938 -20839 20950 -20805
rect 20892 -20873 20950 -20839
rect 20892 -20907 20904 -20873
rect 20938 -20907 20950 -20873
rect 20892 -20952 20950 -20907
rect 21910 -20397 21968 -20352
rect 21910 -20431 21922 -20397
rect 21956 -20431 21968 -20397
rect 21910 -20465 21968 -20431
rect 21910 -20499 21922 -20465
rect 21956 -20499 21968 -20465
rect 21910 -20533 21968 -20499
rect 21910 -20567 21922 -20533
rect 21956 -20567 21968 -20533
rect 21910 -20601 21968 -20567
rect 21910 -20635 21922 -20601
rect 21956 -20635 21968 -20601
rect 21910 -20669 21968 -20635
rect 21910 -20703 21922 -20669
rect 21956 -20703 21968 -20669
rect 21910 -20737 21968 -20703
rect 21910 -20771 21922 -20737
rect 21956 -20771 21968 -20737
rect 21910 -20805 21968 -20771
rect 21910 -20839 21922 -20805
rect 21956 -20839 21968 -20805
rect 21910 -20873 21968 -20839
rect 21910 -20907 21922 -20873
rect 21956 -20907 21968 -20873
rect 21910 -20952 21968 -20907
rect 22928 -20397 22986 -20352
rect 22928 -20431 22940 -20397
rect 22974 -20431 22986 -20397
rect 22928 -20465 22986 -20431
rect 22928 -20499 22940 -20465
rect 22974 -20499 22986 -20465
rect 22928 -20533 22986 -20499
rect 22928 -20567 22940 -20533
rect 22974 -20567 22986 -20533
rect 22928 -20601 22986 -20567
rect 22928 -20635 22940 -20601
rect 22974 -20635 22986 -20601
rect 22928 -20669 22986 -20635
rect 22928 -20703 22940 -20669
rect 22974 -20703 22986 -20669
rect 22928 -20737 22986 -20703
rect 22928 -20771 22940 -20737
rect 22974 -20771 22986 -20737
rect 22928 -20805 22986 -20771
rect 22928 -20839 22940 -20805
rect 22974 -20839 22986 -20805
rect 22928 -20873 22986 -20839
rect 22928 -20907 22940 -20873
rect 22974 -20907 22986 -20873
rect 22928 -20952 22986 -20907
rect 2568 -21629 2626 -21584
rect 2568 -21663 2580 -21629
rect 2614 -21663 2626 -21629
rect 2568 -21697 2626 -21663
rect 2568 -21731 2580 -21697
rect 2614 -21731 2626 -21697
rect 2568 -21765 2626 -21731
rect -9417 -21826 -9359 -21781
rect -9417 -21860 -9405 -21826
rect -9371 -21860 -9359 -21826
rect -9417 -21894 -9359 -21860
rect -9417 -21928 -9405 -21894
rect -9371 -21928 -9359 -21894
rect -9417 -21962 -9359 -21928
rect -9417 -21996 -9405 -21962
rect -9371 -21996 -9359 -21962
rect -9417 -22030 -9359 -21996
rect -9417 -22064 -9405 -22030
rect -9371 -22064 -9359 -22030
rect -9417 -22098 -9359 -22064
rect -9417 -22132 -9405 -22098
rect -9371 -22132 -9359 -22098
rect -9417 -22166 -9359 -22132
rect -9417 -22200 -9405 -22166
rect -9371 -22200 -9359 -22166
rect -9417 -22234 -9359 -22200
rect -9417 -22268 -9405 -22234
rect -9371 -22268 -9359 -22234
rect -9417 -22302 -9359 -22268
rect -9417 -22336 -9405 -22302
rect -9371 -22336 -9359 -22302
rect -9417 -22381 -9359 -22336
rect -8399 -21826 -8341 -21781
rect -8399 -21860 -8387 -21826
rect -8353 -21860 -8341 -21826
rect -8399 -21894 -8341 -21860
rect -8399 -21928 -8387 -21894
rect -8353 -21928 -8341 -21894
rect -8399 -21962 -8341 -21928
rect -8399 -21996 -8387 -21962
rect -8353 -21996 -8341 -21962
rect -8399 -22030 -8341 -21996
rect -8399 -22064 -8387 -22030
rect -8353 -22064 -8341 -22030
rect -8399 -22098 -8341 -22064
rect -8399 -22132 -8387 -22098
rect -8353 -22132 -8341 -22098
rect -8399 -22166 -8341 -22132
rect -8399 -22200 -8387 -22166
rect -8353 -22200 -8341 -22166
rect -8399 -22234 -8341 -22200
rect -8399 -22268 -8387 -22234
rect -8353 -22268 -8341 -22234
rect -8399 -22302 -8341 -22268
rect -8399 -22336 -8387 -22302
rect -8353 -22336 -8341 -22302
rect -8399 -22381 -8341 -22336
rect -7381 -21826 -7323 -21781
rect -7381 -21860 -7369 -21826
rect -7335 -21860 -7323 -21826
rect -7381 -21894 -7323 -21860
rect -7381 -21928 -7369 -21894
rect -7335 -21928 -7323 -21894
rect -7381 -21962 -7323 -21928
rect -7381 -21996 -7369 -21962
rect -7335 -21996 -7323 -21962
rect -7381 -22030 -7323 -21996
rect -7381 -22064 -7369 -22030
rect -7335 -22064 -7323 -22030
rect -7381 -22098 -7323 -22064
rect -7381 -22132 -7369 -22098
rect -7335 -22132 -7323 -22098
rect -7381 -22166 -7323 -22132
rect -7381 -22200 -7369 -22166
rect -7335 -22200 -7323 -22166
rect -7381 -22234 -7323 -22200
rect -7381 -22268 -7369 -22234
rect -7335 -22268 -7323 -22234
rect -7381 -22302 -7323 -22268
rect -7381 -22336 -7369 -22302
rect -7335 -22336 -7323 -22302
rect -7381 -22381 -7323 -22336
rect -6363 -21826 -6305 -21781
rect -6363 -21860 -6351 -21826
rect -6317 -21860 -6305 -21826
rect -6363 -21894 -6305 -21860
rect -6363 -21928 -6351 -21894
rect -6317 -21928 -6305 -21894
rect -6363 -21962 -6305 -21928
rect -6363 -21996 -6351 -21962
rect -6317 -21996 -6305 -21962
rect -6363 -22030 -6305 -21996
rect -6363 -22064 -6351 -22030
rect -6317 -22064 -6305 -22030
rect -6363 -22098 -6305 -22064
rect -6363 -22132 -6351 -22098
rect -6317 -22132 -6305 -22098
rect -6363 -22166 -6305 -22132
rect -6363 -22200 -6351 -22166
rect -6317 -22200 -6305 -22166
rect -6363 -22234 -6305 -22200
rect -6363 -22268 -6351 -22234
rect -6317 -22268 -6305 -22234
rect -6363 -22302 -6305 -22268
rect -6363 -22336 -6351 -22302
rect -6317 -22336 -6305 -22302
rect -6363 -22381 -6305 -22336
rect -5345 -21826 -5287 -21781
rect -5345 -21860 -5333 -21826
rect -5299 -21860 -5287 -21826
rect -5345 -21894 -5287 -21860
rect -5345 -21928 -5333 -21894
rect -5299 -21928 -5287 -21894
rect -5345 -21962 -5287 -21928
rect -5345 -21996 -5333 -21962
rect -5299 -21996 -5287 -21962
rect -5345 -22030 -5287 -21996
rect -5345 -22064 -5333 -22030
rect -5299 -22064 -5287 -22030
rect -5345 -22098 -5287 -22064
rect -5345 -22132 -5333 -22098
rect -5299 -22132 -5287 -22098
rect -5345 -22166 -5287 -22132
rect -5345 -22200 -5333 -22166
rect -5299 -22200 -5287 -22166
rect -5345 -22234 -5287 -22200
rect -5345 -22268 -5333 -22234
rect -5299 -22268 -5287 -22234
rect -5345 -22302 -5287 -22268
rect -5345 -22336 -5333 -22302
rect -5299 -22336 -5287 -22302
rect -5345 -22381 -5287 -22336
rect -4327 -21826 -4269 -21781
rect -4327 -21860 -4315 -21826
rect -4281 -21860 -4269 -21826
rect -4327 -21894 -4269 -21860
rect -4327 -21928 -4315 -21894
rect -4281 -21928 -4269 -21894
rect -4327 -21962 -4269 -21928
rect -4327 -21996 -4315 -21962
rect -4281 -21996 -4269 -21962
rect -4327 -22030 -4269 -21996
rect -4327 -22064 -4315 -22030
rect -4281 -22064 -4269 -22030
rect -4327 -22098 -4269 -22064
rect -4327 -22132 -4315 -22098
rect -4281 -22132 -4269 -22098
rect -4327 -22166 -4269 -22132
rect -4327 -22200 -4315 -22166
rect -4281 -22200 -4269 -22166
rect -4327 -22234 -4269 -22200
rect -4327 -22268 -4315 -22234
rect -4281 -22268 -4269 -22234
rect -4327 -22302 -4269 -22268
rect -4327 -22336 -4315 -22302
rect -4281 -22336 -4269 -22302
rect -4327 -22381 -4269 -22336
rect -3309 -21826 -3251 -21781
rect -3309 -21860 -3297 -21826
rect -3263 -21860 -3251 -21826
rect -3309 -21894 -3251 -21860
rect -3309 -21928 -3297 -21894
rect -3263 -21928 -3251 -21894
rect -3309 -21962 -3251 -21928
rect -3309 -21996 -3297 -21962
rect -3263 -21996 -3251 -21962
rect -3309 -22030 -3251 -21996
rect -3309 -22064 -3297 -22030
rect -3263 -22064 -3251 -22030
rect -3309 -22098 -3251 -22064
rect -3309 -22132 -3297 -22098
rect -3263 -22132 -3251 -22098
rect -3309 -22166 -3251 -22132
rect -3309 -22200 -3297 -22166
rect -3263 -22200 -3251 -22166
rect -3309 -22234 -3251 -22200
rect -3309 -22268 -3297 -22234
rect -3263 -22268 -3251 -22234
rect -3309 -22302 -3251 -22268
rect -3309 -22336 -3297 -22302
rect -3263 -22336 -3251 -22302
rect -3309 -22381 -3251 -22336
rect -2422 -21825 -2364 -21780
rect -2422 -21859 -2410 -21825
rect -2376 -21859 -2364 -21825
rect -2422 -21893 -2364 -21859
rect -2422 -21927 -2410 -21893
rect -2376 -21927 -2364 -21893
rect -2422 -21961 -2364 -21927
rect -2422 -21995 -2410 -21961
rect -2376 -21995 -2364 -21961
rect -2422 -22029 -2364 -21995
rect -2422 -22063 -2410 -22029
rect -2376 -22063 -2364 -22029
rect -2422 -22097 -2364 -22063
rect -2422 -22131 -2410 -22097
rect -2376 -22131 -2364 -22097
rect -2422 -22165 -2364 -22131
rect -2422 -22199 -2410 -22165
rect -2376 -22199 -2364 -22165
rect -2422 -22233 -2364 -22199
rect -2422 -22267 -2410 -22233
rect -2376 -22267 -2364 -22233
rect -2422 -22301 -2364 -22267
rect -2422 -22335 -2410 -22301
rect -2376 -22335 -2364 -22301
rect -2422 -22380 -2364 -22335
rect -2124 -21825 -2066 -21780
rect -2124 -21859 -2112 -21825
rect -2078 -21859 -2066 -21825
rect -2124 -21893 -2066 -21859
rect -2124 -21927 -2112 -21893
rect -2078 -21927 -2066 -21893
rect -2124 -21961 -2066 -21927
rect -2124 -21995 -2112 -21961
rect -2078 -21995 -2066 -21961
rect -2124 -22029 -2066 -21995
rect -2124 -22063 -2112 -22029
rect -2078 -22063 -2066 -22029
rect -2124 -22097 -2066 -22063
rect -2124 -22131 -2112 -22097
rect -2078 -22131 -2066 -22097
rect -2124 -22165 -2066 -22131
rect -2124 -22199 -2112 -22165
rect -2078 -22199 -2066 -22165
rect -2124 -22233 -2066 -22199
rect -2124 -22267 -2112 -22233
rect -2078 -22267 -2066 -22233
rect -2124 -22301 -2066 -22267
rect -2124 -22335 -2112 -22301
rect -2078 -22335 -2066 -22301
rect -2124 -22380 -2066 -22335
rect -1826 -21825 -1768 -21780
rect -1826 -21859 -1814 -21825
rect -1780 -21859 -1768 -21825
rect -1826 -21893 -1768 -21859
rect -1826 -21927 -1814 -21893
rect -1780 -21927 -1768 -21893
rect -1826 -21961 -1768 -21927
rect -1826 -21995 -1814 -21961
rect -1780 -21995 -1768 -21961
rect -1826 -22029 -1768 -21995
rect -1826 -22063 -1814 -22029
rect -1780 -22063 -1768 -22029
rect -1826 -22097 -1768 -22063
rect -1826 -22131 -1814 -22097
rect -1780 -22131 -1768 -22097
rect -1826 -22165 -1768 -22131
rect -1826 -22199 -1814 -22165
rect -1780 -22199 -1768 -22165
rect -1826 -22233 -1768 -22199
rect -1826 -22267 -1814 -22233
rect -1780 -22267 -1768 -22233
rect -1826 -22301 -1768 -22267
rect -1826 -22335 -1814 -22301
rect -1780 -22335 -1768 -22301
rect -1826 -22380 -1768 -22335
rect -1528 -21825 -1470 -21780
rect -1528 -21859 -1516 -21825
rect -1482 -21859 -1470 -21825
rect -1528 -21893 -1470 -21859
rect -1528 -21927 -1516 -21893
rect -1482 -21927 -1470 -21893
rect -1528 -21961 -1470 -21927
rect -1528 -21995 -1516 -21961
rect -1482 -21995 -1470 -21961
rect -1528 -22029 -1470 -21995
rect -1528 -22063 -1516 -22029
rect -1482 -22063 -1470 -22029
rect -1528 -22097 -1470 -22063
rect -1528 -22131 -1516 -22097
rect -1482 -22131 -1470 -22097
rect -1528 -22165 -1470 -22131
rect -1528 -22199 -1516 -22165
rect -1482 -22199 -1470 -22165
rect -1528 -22233 -1470 -22199
rect -1528 -22267 -1516 -22233
rect -1482 -22267 -1470 -22233
rect -1528 -22301 -1470 -22267
rect -1528 -22335 -1516 -22301
rect -1482 -22335 -1470 -22301
rect -1528 -22380 -1470 -22335
rect -1230 -21825 -1172 -21780
rect -1230 -21859 -1218 -21825
rect -1184 -21859 -1172 -21825
rect -1230 -21893 -1172 -21859
rect -1230 -21927 -1218 -21893
rect -1184 -21927 -1172 -21893
rect -1230 -21961 -1172 -21927
rect -1230 -21995 -1218 -21961
rect -1184 -21995 -1172 -21961
rect -1230 -22029 -1172 -21995
rect -1230 -22063 -1218 -22029
rect -1184 -22063 -1172 -22029
rect -1230 -22097 -1172 -22063
rect -1230 -22131 -1218 -22097
rect -1184 -22131 -1172 -22097
rect -1230 -22165 -1172 -22131
rect -1230 -22199 -1218 -22165
rect -1184 -22199 -1172 -22165
rect -1230 -22233 -1172 -22199
rect -1230 -22267 -1218 -22233
rect -1184 -22267 -1172 -22233
rect -1230 -22301 -1172 -22267
rect -1230 -22335 -1218 -22301
rect -1184 -22335 -1172 -22301
rect -1230 -22380 -1172 -22335
rect -932 -21825 -874 -21780
rect -932 -21859 -920 -21825
rect -886 -21859 -874 -21825
rect -932 -21893 -874 -21859
rect -932 -21927 -920 -21893
rect -886 -21927 -874 -21893
rect -932 -21961 -874 -21927
rect -932 -21995 -920 -21961
rect -886 -21995 -874 -21961
rect -932 -22029 -874 -21995
rect -932 -22063 -920 -22029
rect -886 -22063 -874 -22029
rect -932 -22097 -874 -22063
rect -932 -22131 -920 -22097
rect -886 -22131 -874 -22097
rect -932 -22165 -874 -22131
rect -932 -22199 -920 -22165
rect -886 -22199 -874 -22165
rect -932 -22233 -874 -22199
rect -932 -22267 -920 -22233
rect -886 -22267 -874 -22233
rect -932 -22301 -874 -22267
rect -932 -22335 -920 -22301
rect -886 -22335 -874 -22301
rect -932 -22380 -874 -22335
rect -634 -21825 -576 -21780
rect -634 -21859 -622 -21825
rect -588 -21859 -576 -21825
rect -634 -21893 -576 -21859
rect -634 -21927 -622 -21893
rect -588 -21927 -576 -21893
rect -634 -21961 -576 -21927
rect -634 -21995 -622 -21961
rect -588 -21995 -576 -21961
rect -634 -22029 -576 -21995
rect -634 -22063 -622 -22029
rect -588 -22063 -576 -22029
rect -634 -22097 -576 -22063
rect -634 -22131 -622 -22097
rect -588 -22131 -576 -22097
rect -634 -22165 -576 -22131
rect -634 -22199 -622 -22165
rect -588 -22199 -576 -22165
rect -634 -22233 -576 -22199
rect -634 -22267 -622 -22233
rect -588 -22267 -576 -22233
rect -634 -22301 -576 -22267
rect -634 -22335 -622 -22301
rect -588 -22335 -576 -22301
rect -634 -22380 -576 -22335
rect -336 -21825 -278 -21780
rect -336 -21859 -324 -21825
rect -290 -21859 -278 -21825
rect -336 -21893 -278 -21859
rect -336 -21927 -324 -21893
rect -290 -21927 -278 -21893
rect -336 -21961 -278 -21927
rect -336 -21995 -324 -21961
rect -290 -21995 -278 -21961
rect -336 -22029 -278 -21995
rect -336 -22063 -324 -22029
rect -290 -22063 -278 -22029
rect -336 -22097 -278 -22063
rect -336 -22131 -324 -22097
rect -290 -22131 -278 -22097
rect -336 -22165 -278 -22131
rect -336 -22199 -324 -22165
rect -290 -22199 -278 -22165
rect -336 -22233 -278 -22199
rect -336 -22267 -324 -22233
rect -290 -22267 -278 -22233
rect -336 -22301 -278 -22267
rect -336 -22335 -324 -22301
rect -290 -22335 -278 -22301
rect -336 -22380 -278 -22335
rect -38 -21825 20 -21780
rect -38 -21859 -26 -21825
rect 8 -21859 20 -21825
rect -38 -21893 20 -21859
rect -38 -21927 -26 -21893
rect 8 -21927 20 -21893
rect -38 -21961 20 -21927
rect -38 -21995 -26 -21961
rect 8 -21995 20 -21961
rect -38 -22029 20 -21995
rect -38 -22063 -26 -22029
rect 8 -22063 20 -22029
rect -38 -22097 20 -22063
rect -38 -22131 -26 -22097
rect 8 -22131 20 -22097
rect -38 -22165 20 -22131
rect -38 -22199 -26 -22165
rect 8 -22199 20 -22165
rect -38 -22233 20 -22199
rect -38 -22267 -26 -22233
rect 8 -22267 20 -22233
rect -38 -22301 20 -22267
rect -38 -22335 -26 -22301
rect 8 -22335 20 -22301
rect -38 -22380 20 -22335
rect 260 -21825 318 -21780
rect 260 -21859 272 -21825
rect 306 -21859 318 -21825
rect 260 -21893 318 -21859
rect 260 -21927 272 -21893
rect 306 -21927 318 -21893
rect 260 -21961 318 -21927
rect 260 -21995 272 -21961
rect 306 -21995 318 -21961
rect 260 -22029 318 -21995
rect 260 -22063 272 -22029
rect 306 -22063 318 -22029
rect 260 -22097 318 -22063
rect 260 -22131 272 -22097
rect 306 -22131 318 -22097
rect 260 -22165 318 -22131
rect 260 -22199 272 -22165
rect 306 -22199 318 -22165
rect 260 -22233 318 -22199
rect 260 -22267 272 -22233
rect 306 -22267 318 -22233
rect 260 -22301 318 -22267
rect 260 -22335 272 -22301
rect 306 -22335 318 -22301
rect 260 -22380 318 -22335
rect 558 -21825 616 -21780
rect 558 -21859 570 -21825
rect 604 -21859 616 -21825
rect 558 -21893 616 -21859
rect 558 -21927 570 -21893
rect 604 -21927 616 -21893
rect 558 -21961 616 -21927
rect 558 -21995 570 -21961
rect 604 -21995 616 -21961
rect 558 -22029 616 -21995
rect 558 -22063 570 -22029
rect 604 -22063 616 -22029
rect 558 -22097 616 -22063
rect 558 -22131 570 -22097
rect 604 -22131 616 -22097
rect 558 -22165 616 -22131
rect 558 -22199 570 -22165
rect 604 -22199 616 -22165
rect 558 -22233 616 -22199
rect 558 -22267 570 -22233
rect 604 -22267 616 -22233
rect 558 -22301 616 -22267
rect 558 -22335 570 -22301
rect 604 -22335 616 -22301
rect 558 -22380 616 -22335
rect 856 -21825 914 -21780
rect 856 -21859 868 -21825
rect 902 -21859 914 -21825
rect 856 -21893 914 -21859
rect 856 -21927 868 -21893
rect 902 -21927 914 -21893
rect 856 -21961 914 -21927
rect 856 -21995 868 -21961
rect 902 -21995 914 -21961
rect 856 -22029 914 -21995
rect 856 -22063 868 -22029
rect 902 -22063 914 -22029
rect 856 -22097 914 -22063
rect 856 -22131 868 -22097
rect 902 -22131 914 -22097
rect 856 -22165 914 -22131
rect 856 -22199 868 -22165
rect 902 -22199 914 -22165
rect 2568 -21799 2580 -21765
rect 2614 -21799 2626 -21765
rect 2568 -21833 2626 -21799
rect 2568 -21867 2580 -21833
rect 2614 -21867 2626 -21833
rect 2568 -21901 2626 -21867
rect 2568 -21935 2580 -21901
rect 2614 -21935 2626 -21901
rect 2568 -21969 2626 -21935
rect 2568 -22003 2580 -21969
rect 2614 -22003 2626 -21969
rect 2568 -22037 2626 -22003
rect 2568 -22071 2580 -22037
rect 2614 -22071 2626 -22037
rect 2568 -22105 2626 -22071
rect 2568 -22139 2580 -22105
rect 2614 -22139 2626 -22105
rect 2568 -22184 2626 -22139
rect 3586 -21629 3644 -21584
rect 3586 -21663 3598 -21629
rect 3632 -21663 3644 -21629
rect 3586 -21697 3644 -21663
rect 3586 -21731 3598 -21697
rect 3632 -21731 3644 -21697
rect 3586 -21765 3644 -21731
rect 3586 -21799 3598 -21765
rect 3632 -21799 3644 -21765
rect 3586 -21833 3644 -21799
rect 3586 -21867 3598 -21833
rect 3632 -21867 3644 -21833
rect 3586 -21901 3644 -21867
rect 3586 -21935 3598 -21901
rect 3632 -21935 3644 -21901
rect 3586 -21969 3644 -21935
rect 3586 -22003 3598 -21969
rect 3632 -22003 3644 -21969
rect 3586 -22037 3644 -22003
rect 3586 -22071 3598 -22037
rect 3632 -22071 3644 -22037
rect 3586 -22105 3644 -22071
rect 3586 -22139 3598 -22105
rect 3632 -22139 3644 -22105
rect 3586 -22184 3644 -22139
rect 4604 -21629 4662 -21584
rect 4604 -21663 4616 -21629
rect 4650 -21663 4662 -21629
rect 4604 -21697 4662 -21663
rect 4604 -21731 4616 -21697
rect 4650 -21731 4662 -21697
rect 4604 -21765 4662 -21731
rect 4604 -21799 4616 -21765
rect 4650 -21799 4662 -21765
rect 4604 -21833 4662 -21799
rect 4604 -21867 4616 -21833
rect 4650 -21867 4662 -21833
rect 4604 -21901 4662 -21867
rect 4604 -21935 4616 -21901
rect 4650 -21935 4662 -21901
rect 4604 -21969 4662 -21935
rect 4604 -22003 4616 -21969
rect 4650 -22003 4662 -21969
rect 4604 -22037 4662 -22003
rect 4604 -22071 4616 -22037
rect 4650 -22071 4662 -22037
rect 4604 -22105 4662 -22071
rect 4604 -22139 4616 -22105
rect 4650 -22139 4662 -22105
rect 4604 -22184 4662 -22139
rect 5622 -21629 5680 -21584
rect 5622 -21663 5634 -21629
rect 5668 -21663 5680 -21629
rect 5622 -21697 5680 -21663
rect 5622 -21731 5634 -21697
rect 5668 -21731 5680 -21697
rect 5622 -21765 5680 -21731
rect 5622 -21799 5634 -21765
rect 5668 -21799 5680 -21765
rect 5622 -21833 5680 -21799
rect 5622 -21867 5634 -21833
rect 5668 -21867 5680 -21833
rect 5622 -21901 5680 -21867
rect 5622 -21935 5634 -21901
rect 5668 -21935 5680 -21901
rect 5622 -21969 5680 -21935
rect 5622 -22003 5634 -21969
rect 5668 -22003 5680 -21969
rect 5622 -22037 5680 -22003
rect 5622 -22071 5634 -22037
rect 5668 -22071 5680 -22037
rect 5622 -22105 5680 -22071
rect 5622 -22139 5634 -22105
rect 5668 -22139 5680 -22105
rect 5622 -22184 5680 -22139
rect 6640 -21629 6698 -21584
rect 6640 -21663 6652 -21629
rect 6686 -21663 6698 -21629
rect 6640 -21697 6698 -21663
rect 6640 -21731 6652 -21697
rect 6686 -21731 6698 -21697
rect 6640 -21765 6698 -21731
rect 6640 -21799 6652 -21765
rect 6686 -21799 6698 -21765
rect 6640 -21833 6698 -21799
rect 6640 -21867 6652 -21833
rect 6686 -21867 6698 -21833
rect 6640 -21901 6698 -21867
rect 6640 -21935 6652 -21901
rect 6686 -21935 6698 -21901
rect 6640 -21969 6698 -21935
rect 6640 -22003 6652 -21969
rect 6686 -22003 6698 -21969
rect 6640 -22037 6698 -22003
rect 6640 -22071 6652 -22037
rect 6686 -22071 6698 -22037
rect 6640 -22105 6698 -22071
rect 6640 -22139 6652 -22105
rect 6686 -22139 6698 -22105
rect 6640 -22184 6698 -22139
rect 7658 -21629 7716 -21584
rect 7658 -21663 7670 -21629
rect 7704 -21663 7716 -21629
rect 7658 -21697 7716 -21663
rect 7658 -21731 7670 -21697
rect 7704 -21731 7716 -21697
rect 7658 -21765 7716 -21731
rect 7658 -21799 7670 -21765
rect 7704 -21799 7716 -21765
rect 7658 -21833 7716 -21799
rect 7658 -21867 7670 -21833
rect 7704 -21867 7716 -21833
rect 7658 -21901 7716 -21867
rect 7658 -21935 7670 -21901
rect 7704 -21935 7716 -21901
rect 7658 -21969 7716 -21935
rect 7658 -22003 7670 -21969
rect 7704 -22003 7716 -21969
rect 7658 -22037 7716 -22003
rect 7658 -22071 7670 -22037
rect 7704 -22071 7716 -22037
rect 7658 -22105 7716 -22071
rect 7658 -22139 7670 -22105
rect 7704 -22139 7716 -22105
rect 7658 -22184 7716 -22139
rect 8676 -21629 8734 -21584
rect 8676 -21663 8688 -21629
rect 8722 -21663 8734 -21629
rect 8676 -21697 8734 -21663
rect 8676 -21731 8688 -21697
rect 8722 -21731 8734 -21697
rect 8676 -21765 8734 -21731
rect 8676 -21799 8688 -21765
rect 8722 -21799 8734 -21765
rect 8676 -21833 8734 -21799
rect 8676 -21867 8688 -21833
rect 8722 -21867 8734 -21833
rect 8676 -21901 8734 -21867
rect 8676 -21935 8688 -21901
rect 8722 -21935 8734 -21901
rect 8676 -21969 8734 -21935
rect 8676 -22003 8688 -21969
rect 8722 -22003 8734 -21969
rect 8676 -22037 8734 -22003
rect 8676 -22071 8688 -22037
rect 8722 -22071 8734 -22037
rect 8676 -22105 8734 -22071
rect 8676 -22139 8688 -22105
rect 8722 -22139 8734 -22105
rect 8676 -22184 8734 -22139
rect 9694 -21629 9752 -21584
rect 9694 -21663 9706 -21629
rect 9740 -21663 9752 -21629
rect 9694 -21697 9752 -21663
rect 9694 -21731 9706 -21697
rect 9740 -21731 9752 -21697
rect 9694 -21765 9752 -21731
rect 9694 -21799 9706 -21765
rect 9740 -21799 9752 -21765
rect 9694 -21833 9752 -21799
rect 9694 -21867 9706 -21833
rect 9740 -21867 9752 -21833
rect 9694 -21901 9752 -21867
rect 9694 -21935 9706 -21901
rect 9740 -21935 9752 -21901
rect 9694 -21969 9752 -21935
rect 9694 -22003 9706 -21969
rect 9740 -22003 9752 -21969
rect 9694 -22037 9752 -22003
rect 9694 -22071 9706 -22037
rect 9740 -22071 9752 -22037
rect 9694 -22105 9752 -22071
rect 9694 -22139 9706 -22105
rect 9740 -22139 9752 -22105
rect 9694 -22184 9752 -22139
rect 10712 -21629 10770 -21584
rect 10712 -21663 10724 -21629
rect 10758 -21663 10770 -21629
rect 10712 -21697 10770 -21663
rect 10712 -21731 10724 -21697
rect 10758 -21731 10770 -21697
rect 10712 -21765 10770 -21731
rect 10712 -21799 10724 -21765
rect 10758 -21799 10770 -21765
rect 10712 -21833 10770 -21799
rect 10712 -21867 10724 -21833
rect 10758 -21867 10770 -21833
rect 10712 -21901 10770 -21867
rect 10712 -21935 10724 -21901
rect 10758 -21935 10770 -21901
rect 10712 -21969 10770 -21935
rect 10712 -22003 10724 -21969
rect 10758 -22003 10770 -21969
rect 10712 -22037 10770 -22003
rect 10712 -22071 10724 -22037
rect 10758 -22071 10770 -22037
rect 10712 -22105 10770 -22071
rect 10712 -22139 10724 -22105
rect 10758 -22139 10770 -22105
rect 10712 -22184 10770 -22139
rect 11730 -21629 11788 -21584
rect 11730 -21663 11742 -21629
rect 11776 -21663 11788 -21629
rect 11730 -21697 11788 -21663
rect 11730 -21731 11742 -21697
rect 11776 -21731 11788 -21697
rect 11730 -21765 11788 -21731
rect 11730 -21799 11742 -21765
rect 11776 -21799 11788 -21765
rect 11730 -21833 11788 -21799
rect 11730 -21867 11742 -21833
rect 11776 -21867 11788 -21833
rect 11730 -21901 11788 -21867
rect 11730 -21935 11742 -21901
rect 11776 -21935 11788 -21901
rect 11730 -21969 11788 -21935
rect 11730 -22003 11742 -21969
rect 11776 -22003 11788 -21969
rect 11730 -22037 11788 -22003
rect 11730 -22071 11742 -22037
rect 11776 -22071 11788 -22037
rect 11730 -22105 11788 -22071
rect 11730 -22139 11742 -22105
rect 11776 -22139 11788 -22105
rect 11730 -22184 11788 -22139
rect 12748 -21629 12806 -21584
rect 12748 -21663 12760 -21629
rect 12794 -21663 12806 -21629
rect 12748 -21697 12806 -21663
rect 12748 -21731 12760 -21697
rect 12794 -21731 12806 -21697
rect 12748 -21765 12806 -21731
rect 12748 -21799 12760 -21765
rect 12794 -21799 12806 -21765
rect 12748 -21833 12806 -21799
rect 12748 -21867 12760 -21833
rect 12794 -21867 12806 -21833
rect 12748 -21901 12806 -21867
rect 12748 -21935 12760 -21901
rect 12794 -21935 12806 -21901
rect 12748 -21969 12806 -21935
rect 12748 -22003 12760 -21969
rect 12794 -22003 12806 -21969
rect 12748 -22037 12806 -22003
rect 12748 -22071 12760 -22037
rect 12794 -22071 12806 -22037
rect 12748 -22105 12806 -22071
rect 12748 -22139 12760 -22105
rect 12794 -22139 12806 -22105
rect 12748 -22184 12806 -22139
rect 13766 -21629 13824 -21584
rect 13766 -21663 13778 -21629
rect 13812 -21663 13824 -21629
rect 13766 -21697 13824 -21663
rect 13766 -21731 13778 -21697
rect 13812 -21731 13824 -21697
rect 13766 -21765 13824 -21731
rect 13766 -21799 13778 -21765
rect 13812 -21799 13824 -21765
rect 13766 -21833 13824 -21799
rect 13766 -21867 13778 -21833
rect 13812 -21867 13824 -21833
rect 13766 -21901 13824 -21867
rect 13766 -21935 13778 -21901
rect 13812 -21935 13824 -21901
rect 13766 -21969 13824 -21935
rect 13766 -22003 13778 -21969
rect 13812 -22003 13824 -21969
rect 13766 -22037 13824 -22003
rect 13766 -22071 13778 -22037
rect 13812 -22071 13824 -22037
rect 13766 -22105 13824 -22071
rect 13766 -22139 13778 -22105
rect 13812 -22139 13824 -22105
rect 13766 -22184 13824 -22139
rect 14784 -21629 14842 -21584
rect 14784 -21663 14796 -21629
rect 14830 -21663 14842 -21629
rect 14784 -21697 14842 -21663
rect 14784 -21731 14796 -21697
rect 14830 -21731 14842 -21697
rect 14784 -21765 14842 -21731
rect 14784 -21799 14796 -21765
rect 14830 -21799 14842 -21765
rect 14784 -21833 14842 -21799
rect 14784 -21867 14796 -21833
rect 14830 -21867 14842 -21833
rect 14784 -21901 14842 -21867
rect 14784 -21935 14796 -21901
rect 14830 -21935 14842 -21901
rect 14784 -21969 14842 -21935
rect 14784 -22003 14796 -21969
rect 14830 -22003 14842 -21969
rect 14784 -22037 14842 -22003
rect 14784 -22071 14796 -22037
rect 14830 -22071 14842 -22037
rect 14784 -22105 14842 -22071
rect 14784 -22139 14796 -22105
rect 14830 -22139 14842 -22105
rect 14784 -22184 14842 -22139
rect 15802 -21629 15860 -21584
rect 15802 -21663 15814 -21629
rect 15848 -21663 15860 -21629
rect 15802 -21697 15860 -21663
rect 15802 -21731 15814 -21697
rect 15848 -21731 15860 -21697
rect 15802 -21765 15860 -21731
rect 15802 -21799 15814 -21765
rect 15848 -21799 15860 -21765
rect 15802 -21833 15860 -21799
rect 15802 -21867 15814 -21833
rect 15848 -21867 15860 -21833
rect 15802 -21901 15860 -21867
rect 15802 -21935 15814 -21901
rect 15848 -21935 15860 -21901
rect 15802 -21969 15860 -21935
rect 15802 -22003 15814 -21969
rect 15848 -22003 15860 -21969
rect 15802 -22037 15860 -22003
rect 15802 -22071 15814 -22037
rect 15848 -22071 15860 -22037
rect 15802 -22105 15860 -22071
rect 15802 -22139 15814 -22105
rect 15848 -22139 15860 -22105
rect 15802 -22184 15860 -22139
rect 16820 -21629 16878 -21584
rect 16820 -21663 16832 -21629
rect 16866 -21663 16878 -21629
rect 16820 -21697 16878 -21663
rect 16820 -21731 16832 -21697
rect 16866 -21731 16878 -21697
rect 16820 -21765 16878 -21731
rect 16820 -21799 16832 -21765
rect 16866 -21799 16878 -21765
rect 16820 -21833 16878 -21799
rect 16820 -21867 16832 -21833
rect 16866 -21867 16878 -21833
rect 16820 -21901 16878 -21867
rect 16820 -21935 16832 -21901
rect 16866 -21935 16878 -21901
rect 16820 -21969 16878 -21935
rect 16820 -22003 16832 -21969
rect 16866 -22003 16878 -21969
rect 16820 -22037 16878 -22003
rect 16820 -22071 16832 -22037
rect 16866 -22071 16878 -22037
rect 16820 -22105 16878 -22071
rect 16820 -22139 16832 -22105
rect 16866 -22139 16878 -22105
rect 16820 -22184 16878 -22139
rect 17838 -21629 17896 -21584
rect 17838 -21663 17850 -21629
rect 17884 -21663 17896 -21629
rect 17838 -21697 17896 -21663
rect 17838 -21731 17850 -21697
rect 17884 -21731 17896 -21697
rect 17838 -21765 17896 -21731
rect 17838 -21799 17850 -21765
rect 17884 -21799 17896 -21765
rect 17838 -21833 17896 -21799
rect 17838 -21867 17850 -21833
rect 17884 -21867 17896 -21833
rect 17838 -21901 17896 -21867
rect 17838 -21935 17850 -21901
rect 17884 -21935 17896 -21901
rect 17838 -21969 17896 -21935
rect 17838 -22003 17850 -21969
rect 17884 -22003 17896 -21969
rect 17838 -22037 17896 -22003
rect 17838 -22071 17850 -22037
rect 17884 -22071 17896 -22037
rect 17838 -22105 17896 -22071
rect 17838 -22139 17850 -22105
rect 17884 -22139 17896 -22105
rect 17838 -22184 17896 -22139
rect 18856 -21629 18914 -21584
rect 18856 -21663 18868 -21629
rect 18902 -21663 18914 -21629
rect 18856 -21697 18914 -21663
rect 18856 -21731 18868 -21697
rect 18902 -21731 18914 -21697
rect 18856 -21765 18914 -21731
rect 18856 -21799 18868 -21765
rect 18902 -21799 18914 -21765
rect 18856 -21833 18914 -21799
rect 18856 -21867 18868 -21833
rect 18902 -21867 18914 -21833
rect 18856 -21901 18914 -21867
rect 18856 -21935 18868 -21901
rect 18902 -21935 18914 -21901
rect 18856 -21969 18914 -21935
rect 18856 -22003 18868 -21969
rect 18902 -22003 18914 -21969
rect 18856 -22037 18914 -22003
rect 18856 -22071 18868 -22037
rect 18902 -22071 18914 -22037
rect 18856 -22105 18914 -22071
rect 18856 -22139 18868 -22105
rect 18902 -22139 18914 -22105
rect 18856 -22184 18914 -22139
rect 19874 -21629 19932 -21584
rect 19874 -21663 19886 -21629
rect 19920 -21663 19932 -21629
rect 19874 -21697 19932 -21663
rect 19874 -21731 19886 -21697
rect 19920 -21731 19932 -21697
rect 19874 -21765 19932 -21731
rect 19874 -21799 19886 -21765
rect 19920 -21799 19932 -21765
rect 19874 -21833 19932 -21799
rect 19874 -21867 19886 -21833
rect 19920 -21867 19932 -21833
rect 19874 -21901 19932 -21867
rect 19874 -21935 19886 -21901
rect 19920 -21935 19932 -21901
rect 19874 -21969 19932 -21935
rect 19874 -22003 19886 -21969
rect 19920 -22003 19932 -21969
rect 19874 -22037 19932 -22003
rect 19874 -22071 19886 -22037
rect 19920 -22071 19932 -22037
rect 19874 -22105 19932 -22071
rect 19874 -22139 19886 -22105
rect 19920 -22139 19932 -22105
rect 19874 -22184 19932 -22139
rect 20892 -21629 20950 -21584
rect 20892 -21663 20904 -21629
rect 20938 -21663 20950 -21629
rect 20892 -21697 20950 -21663
rect 20892 -21731 20904 -21697
rect 20938 -21731 20950 -21697
rect 20892 -21765 20950 -21731
rect 20892 -21799 20904 -21765
rect 20938 -21799 20950 -21765
rect 20892 -21833 20950 -21799
rect 20892 -21867 20904 -21833
rect 20938 -21867 20950 -21833
rect 20892 -21901 20950 -21867
rect 20892 -21935 20904 -21901
rect 20938 -21935 20950 -21901
rect 20892 -21969 20950 -21935
rect 20892 -22003 20904 -21969
rect 20938 -22003 20950 -21969
rect 20892 -22037 20950 -22003
rect 20892 -22071 20904 -22037
rect 20938 -22071 20950 -22037
rect 20892 -22105 20950 -22071
rect 20892 -22139 20904 -22105
rect 20938 -22139 20950 -22105
rect 20892 -22184 20950 -22139
rect 21910 -21629 21968 -21584
rect 21910 -21663 21922 -21629
rect 21956 -21663 21968 -21629
rect 21910 -21697 21968 -21663
rect 21910 -21731 21922 -21697
rect 21956 -21731 21968 -21697
rect 21910 -21765 21968 -21731
rect 21910 -21799 21922 -21765
rect 21956 -21799 21968 -21765
rect 21910 -21833 21968 -21799
rect 21910 -21867 21922 -21833
rect 21956 -21867 21968 -21833
rect 21910 -21901 21968 -21867
rect 21910 -21935 21922 -21901
rect 21956 -21935 21968 -21901
rect 21910 -21969 21968 -21935
rect 21910 -22003 21922 -21969
rect 21956 -22003 21968 -21969
rect 21910 -22037 21968 -22003
rect 21910 -22071 21922 -22037
rect 21956 -22071 21968 -22037
rect 21910 -22105 21968 -22071
rect 21910 -22139 21922 -22105
rect 21956 -22139 21968 -22105
rect 21910 -22184 21968 -22139
rect 22928 -21629 22986 -21584
rect 22928 -21663 22940 -21629
rect 22974 -21663 22986 -21629
rect 22928 -21697 22986 -21663
rect 22928 -21731 22940 -21697
rect 22974 -21731 22986 -21697
rect 22928 -21765 22986 -21731
rect 22928 -21799 22940 -21765
rect 22974 -21799 22986 -21765
rect 22928 -21833 22986 -21799
rect 22928 -21867 22940 -21833
rect 22974 -21867 22986 -21833
rect 22928 -21901 22986 -21867
rect 22928 -21935 22940 -21901
rect 22974 -21935 22986 -21901
rect 22928 -21969 22986 -21935
rect 22928 -22003 22940 -21969
rect 22974 -22003 22986 -21969
rect 22928 -22037 22986 -22003
rect 22928 -22071 22940 -22037
rect 22974 -22071 22986 -22037
rect 22928 -22105 22986 -22071
rect 22928 -22139 22940 -22105
rect 22974 -22139 22986 -22105
rect 22928 -22184 22986 -22139
rect 856 -22233 914 -22199
rect 856 -22267 868 -22233
rect 902 -22267 914 -22233
rect 856 -22301 914 -22267
rect 856 -22335 868 -22301
rect 902 -22335 914 -22301
rect 856 -22380 914 -22335
rect 2568 -22863 2626 -22818
rect -9418 -22939 -9360 -22894
rect -9418 -22973 -9406 -22939
rect -9372 -22973 -9360 -22939
rect -9418 -23007 -9360 -22973
rect -9418 -23041 -9406 -23007
rect -9372 -23041 -9360 -23007
rect -9418 -23075 -9360 -23041
rect -9418 -23109 -9406 -23075
rect -9372 -23109 -9360 -23075
rect -9418 -23143 -9360 -23109
rect -9418 -23177 -9406 -23143
rect -9372 -23177 -9360 -23143
rect -9418 -23211 -9360 -23177
rect -9418 -23245 -9406 -23211
rect -9372 -23245 -9360 -23211
rect -9418 -23279 -9360 -23245
rect -9418 -23313 -9406 -23279
rect -9372 -23313 -9360 -23279
rect -9418 -23347 -9360 -23313
rect -9418 -23381 -9406 -23347
rect -9372 -23381 -9360 -23347
rect -9418 -23415 -9360 -23381
rect -9418 -23449 -9406 -23415
rect -9372 -23449 -9360 -23415
rect -9418 -23494 -9360 -23449
rect -8400 -22939 -8342 -22894
rect -8400 -22973 -8388 -22939
rect -8354 -22973 -8342 -22939
rect -8400 -23007 -8342 -22973
rect -8400 -23041 -8388 -23007
rect -8354 -23041 -8342 -23007
rect -8400 -23075 -8342 -23041
rect -8400 -23109 -8388 -23075
rect -8354 -23109 -8342 -23075
rect -8400 -23143 -8342 -23109
rect -8400 -23177 -8388 -23143
rect -8354 -23177 -8342 -23143
rect -8400 -23211 -8342 -23177
rect -8400 -23245 -8388 -23211
rect -8354 -23245 -8342 -23211
rect -8400 -23279 -8342 -23245
rect -8400 -23313 -8388 -23279
rect -8354 -23313 -8342 -23279
rect -8400 -23347 -8342 -23313
rect -8400 -23381 -8388 -23347
rect -8354 -23381 -8342 -23347
rect -8400 -23415 -8342 -23381
rect -8400 -23449 -8388 -23415
rect -8354 -23449 -8342 -23415
rect -8400 -23494 -8342 -23449
rect -7382 -22939 -7324 -22894
rect -7382 -22973 -7370 -22939
rect -7336 -22973 -7324 -22939
rect -7382 -23007 -7324 -22973
rect -7382 -23041 -7370 -23007
rect -7336 -23041 -7324 -23007
rect -7382 -23075 -7324 -23041
rect -7382 -23109 -7370 -23075
rect -7336 -23109 -7324 -23075
rect -7382 -23143 -7324 -23109
rect -7382 -23177 -7370 -23143
rect -7336 -23177 -7324 -23143
rect -7382 -23211 -7324 -23177
rect -7382 -23245 -7370 -23211
rect -7336 -23245 -7324 -23211
rect -7382 -23279 -7324 -23245
rect -7382 -23313 -7370 -23279
rect -7336 -23313 -7324 -23279
rect -7382 -23347 -7324 -23313
rect -7382 -23381 -7370 -23347
rect -7336 -23381 -7324 -23347
rect -7382 -23415 -7324 -23381
rect -7382 -23449 -7370 -23415
rect -7336 -23449 -7324 -23415
rect -7382 -23494 -7324 -23449
rect -6364 -22939 -6306 -22894
rect -6364 -22973 -6352 -22939
rect -6318 -22973 -6306 -22939
rect -6364 -23007 -6306 -22973
rect -6364 -23041 -6352 -23007
rect -6318 -23041 -6306 -23007
rect -6364 -23075 -6306 -23041
rect -6364 -23109 -6352 -23075
rect -6318 -23109 -6306 -23075
rect -6364 -23143 -6306 -23109
rect -6364 -23177 -6352 -23143
rect -6318 -23177 -6306 -23143
rect -6364 -23211 -6306 -23177
rect -6364 -23245 -6352 -23211
rect -6318 -23245 -6306 -23211
rect -6364 -23279 -6306 -23245
rect -6364 -23313 -6352 -23279
rect -6318 -23313 -6306 -23279
rect -6364 -23347 -6306 -23313
rect -6364 -23381 -6352 -23347
rect -6318 -23381 -6306 -23347
rect -6364 -23415 -6306 -23381
rect -6364 -23449 -6352 -23415
rect -6318 -23449 -6306 -23415
rect -6364 -23494 -6306 -23449
rect -5346 -22939 -5288 -22894
rect -5346 -22973 -5334 -22939
rect -5300 -22973 -5288 -22939
rect -5346 -23007 -5288 -22973
rect -5346 -23041 -5334 -23007
rect -5300 -23041 -5288 -23007
rect -5346 -23075 -5288 -23041
rect -5346 -23109 -5334 -23075
rect -5300 -23109 -5288 -23075
rect -5346 -23143 -5288 -23109
rect -5346 -23177 -5334 -23143
rect -5300 -23177 -5288 -23143
rect -5346 -23211 -5288 -23177
rect -5346 -23245 -5334 -23211
rect -5300 -23245 -5288 -23211
rect -5346 -23279 -5288 -23245
rect -5346 -23313 -5334 -23279
rect -5300 -23313 -5288 -23279
rect -5346 -23347 -5288 -23313
rect -5346 -23381 -5334 -23347
rect -5300 -23381 -5288 -23347
rect -5346 -23415 -5288 -23381
rect -5346 -23449 -5334 -23415
rect -5300 -23449 -5288 -23415
rect -5346 -23494 -5288 -23449
rect -4328 -22939 -4270 -22894
rect -4328 -22973 -4316 -22939
rect -4282 -22973 -4270 -22939
rect -4328 -23007 -4270 -22973
rect -4328 -23041 -4316 -23007
rect -4282 -23041 -4270 -23007
rect -4328 -23075 -4270 -23041
rect -4328 -23109 -4316 -23075
rect -4282 -23109 -4270 -23075
rect -4328 -23143 -4270 -23109
rect -4328 -23177 -4316 -23143
rect -4282 -23177 -4270 -23143
rect -4328 -23211 -4270 -23177
rect -4328 -23245 -4316 -23211
rect -4282 -23245 -4270 -23211
rect -4328 -23279 -4270 -23245
rect -4328 -23313 -4316 -23279
rect -4282 -23313 -4270 -23279
rect -4328 -23347 -4270 -23313
rect -4328 -23381 -4316 -23347
rect -4282 -23381 -4270 -23347
rect -4328 -23415 -4270 -23381
rect -4328 -23449 -4316 -23415
rect -4282 -23449 -4270 -23415
rect -4328 -23494 -4270 -23449
rect -3310 -22939 -3252 -22894
rect -3310 -22973 -3298 -22939
rect -3264 -22973 -3252 -22939
rect -3310 -23007 -3252 -22973
rect -3310 -23041 -3298 -23007
rect -3264 -23041 -3252 -23007
rect -3310 -23075 -3252 -23041
rect -3310 -23109 -3298 -23075
rect -3264 -23109 -3252 -23075
rect -3310 -23143 -3252 -23109
rect -3310 -23177 -3298 -23143
rect -3264 -23177 -3252 -23143
rect -3310 -23211 -3252 -23177
rect -3310 -23245 -3298 -23211
rect -3264 -23245 -3252 -23211
rect -3310 -23279 -3252 -23245
rect -3310 -23313 -3298 -23279
rect -3264 -23313 -3252 -23279
rect -3310 -23347 -3252 -23313
rect -3310 -23381 -3298 -23347
rect -3264 -23381 -3252 -23347
rect -3310 -23415 -3252 -23381
rect -3310 -23449 -3298 -23415
rect -3264 -23449 -3252 -23415
rect -3310 -23494 -3252 -23449
rect -2422 -22937 -2364 -22892
rect -2422 -22971 -2410 -22937
rect -2376 -22971 -2364 -22937
rect -2422 -23005 -2364 -22971
rect -2422 -23039 -2410 -23005
rect -2376 -23039 -2364 -23005
rect -2422 -23073 -2364 -23039
rect -2422 -23107 -2410 -23073
rect -2376 -23107 -2364 -23073
rect -2422 -23141 -2364 -23107
rect -2422 -23175 -2410 -23141
rect -2376 -23175 -2364 -23141
rect -2422 -23209 -2364 -23175
rect -2422 -23243 -2410 -23209
rect -2376 -23243 -2364 -23209
rect -2422 -23277 -2364 -23243
rect -2422 -23311 -2410 -23277
rect -2376 -23311 -2364 -23277
rect -2422 -23345 -2364 -23311
rect -2422 -23379 -2410 -23345
rect -2376 -23379 -2364 -23345
rect -2422 -23413 -2364 -23379
rect -2422 -23447 -2410 -23413
rect -2376 -23447 -2364 -23413
rect -2422 -23492 -2364 -23447
rect -2124 -22937 -2066 -22892
rect -2124 -22971 -2112 -22937
rect -2078 -22971 -2066 -22937
rect -2124 -23005 -2066 -22971
rect -2124 -23039 -2112 -23005
rect -2078 -23039 -2066 -23005
rect -2124 -23073 -2066 -23039
rect -2124 -23107 -2112 -23073
rect -2078 -23107 -2066 -23073
rect -2124 -23141 -2066 -23107
rect -2124 -23175 -2112 -23141
rect -2078 -23175 -2066 -23141
rect -2124 -23209 -2066 -23175
rect -2124 -23243 -2112 -23209
rect -2078 -23243 -2066 -23209
rect -2124 -23277 -2066 -23243
rect -2124 -23311 -2112 -23277
rect -2078 -23311 -2066 -23277
rect -2124 -23345 -2066 -23311
rect -2124 -23379 -2112 -23345
rect -2078 -23379 -2066 -23345
rect -2124 -23413 -2066 -23379
rect -2124 -23447 -2112 -23413
rect -2078 -23447 -2066 -23413
rect -2124 -23492 -2066 -23447
rect -1826 -22937 -1768 -22892
rect -1826 -22971 -1814 -22937
rect -1780 -22971 -1768 -22937
rect -1826 -23005 -1768 -22971
rect -1826 -23039 -1814 -23005
rect -1780 -23039 -1768 -23005
rect -1826 -23073 -1768 -23039
rect -1826 -23107 -1814 -23073
rect -1780 -23107 -1768 -23073
rect -1826 -23141 -1768 -23107
rect -1826 -23175 -1814 -23141
rect -1780 -23175 -1768 -23141
rect -1826 -23209 -1768 -23175
rect -1826 -23243 -1814 -23209
rect -1780 -23243 -1768 -23209
rect -1826 -23277 -1768 -23243
rect -1826 -23311 -1814 -23277
rect -1780 -23311 -1768 -23277
rect -1826 -23345 -1768 -23311
rect -1826 -23379 -1814 -23345
rect -1780 -23379 -1768 -23345
rect -1826 -23413 -1768 -23379
rect -1826 -23447 -1814 -23413
rect -1780 -23447 -1768 -23413
rect -1826 -23492 -1768 -23447
rect -1528 -22937 -1470 -22892
rect -1528 -22971 -1516 -22937
rect -1482 -22971 -1470 -22937
rect -1528 -23005 -1470 -22971
rect -1528 -23039 -1516 -23005
rect -1482 -23039 -1470 -23005
rect -1528 -23073 -1470 -23039
rect -1528 -23107 -1516 -23073
rect -1482 -23107 -1470 -23073
rect -1528 -23141 -1470 -23107
rect -1528 -23175 -1516 -23141
rect -1482 -23175 -1470 -23141
rect -1528 -23209 -1470 -23175
rect -1528 -23243 -1516 -23209
rect -1482 -23243 -1470 -23209
rect -1528 -23277 -1470 -23243
rect -1528 -23311 -1516 -23277
rect -1482 -23311 -1470 -23277
rect -1528 -23345 -1470 -23311
rect -1528 -23379 -1516 -23345
rect -1482 -23379 -1470 -23345
rect -1528 -23413 -1470 -23379
rect -1528 -23447 -1516 -23413
rect -1482 -23447 -1470 -23413
rect -1528 -23492 -1470 -23447
rect -1230 -22937 -1172 -22892
rect -1230 -22971 -1218 -22937
rect -1184 -22971 -1172 -22937
rect -1230 -23005 -1172 -22971
rect -1230 -23039 -1218 -23005
rect -1184 -23039 -1172 -23005
rect -1230 -23073 -1172 -23039
rect -1230 -23107 -1218 -23073
rect -1184 -23107 -1172 -23073
rect -1230 -23141 -1172 -23107
rect -1230 -23175 -1218 -23141
rect -1184 -23175 -1172 -23141
rect -1230 -23209 -1172 -23175
rect -1230 -23243 -1218 -23209
rect -1184 -23243 -1172 -23209
rect -1230 -23277 -1172 -23243
rect -1230 -23311 -1218 -23277
rect -1184 -23311 -1172 -23277
rect -1230 -23345 -1172 -23311
rect -1230 -23379 -1218 -23345
rect -1184 -23379 -1172 -23345
rect -1230 -23413 -1172 -23379
rect -1230 -23447 -1218 -23413
rect -1184 -23447 -1172 -23413
rect -1230 -23492 -1172 -23447
rect -932 -22937 -874 -22892
rect -932 -22971 -920 -22937
rect -886 -22971 -874 -22937
rect -932 -23005 -874 -22971
rect -932 -23039 -920 -23005
rect -886 -23039 -874 -23005
rect -932 -23073 -874 -23039
rect -932 -23107 -920 -23073
rect -886 -23107 -874 -23073
rect -932 -23141 -874 -23107
rect -932 -23175 -920 -23141
rect -886 -23175 -874 -23141
rect -932 -23209 -874 -23175
rect -932 -23243 -920 -23209
rect -886 -23243 -874 -23209
rect -932 -23277 -874 -23243
rect -932 -23311 -920 -23277
rect -886 -23311 -874 -23277
rect -932 -23345 -874 -23311
rect -932 -23379 -920 -23345
rect -886 -23379 -874 -23345
rect -932 -23413 -874 -23379
rect -932 -23447 -920 -23413
rect -886 -23447 -874 -23413
rect -932 -23492 -874 -23447
rect -634 -22937 -576 -22892
rect -634 -22971 -622 -22937
rect -588 -22971 -576 -22937
rect -634 -23005 -576 -22971
rect -634 -23039 -622 -23005
rect -588 -23039 -576 -23005
rect -634 -23073 -576 -23039
rect -634 -23107 -622 -23073
rect -588 -23107 -576 -23073
rect -634 -23141 -576 -23107
rect -634 -23175 -622 -23141
rect -588 -23175 -576 -23141
rect -634 -23209 -576 -23175
rect -634 -23243 -622 -23209
rect -588 -23243 -576 -23209
rect -634 -23277 -576 -23243
rect -634 -23311 -622 -23277
rect -588 -23311 -576 -23277
rect -634 -23345 -576 -23311
rect -634 -23379 -622 -23345
rect -588 -23379 -576 -23345
rect -634 -23413 -576 -23379
rect -634 -23447 -622 -23413
rect -588 -23447 -576 -23413
rect -634 -23492 -576 -23447
rect -336 -22937 -278 -22892
rect -336 -22971 -324 -22937
rect -290 -22971 -278 -22937
rect -336 -23005 -278 -22971
rect -336 -23039 -324 -23005
rect -290 -23039 -278 -23005
rect -336 -23073 -278 -23039
rect -336 -23107 -324 -23073
rect -290 -23107 -278 -23073
rect -336 -23141 -278 -23107
rect -336 -23175 -324 -23141
rect -290 -23175 -278 -23141
rect -336 -23209 -278 -23175
rect -336 -23243 -324 -23209
rect -290 -23243 -278 -23209
rect -336 -23277 -278 -23243
rect -336 -23311 -324 -23277
rect -290 -23311 -278 -23277
rect -336 -23345 -278 -23311
rect -336 -23379 -324 -23345
rect -290 -23379 -278 -23345
rect -336 -23413 -278 -23379
rect -336 -23447 -324 -23413
rect -290 -23447 -278 -23413
rect -336 -23492 -278 -23447
rect -38 -22937 20 -22892
rect -38 -22971 -26 -22937
rect 8 -22971 20 -22937
rect -38 -23005 20 -22971
rect -38 -23039 -26 -23005
rect 8 -23039 20 -23005
rect -38 -23073 20 -23039
rect -38 -23107 -26 -23073
rect 8 -23107 20 -23073
rect -38 -23141 20 -23107
rect -38 -23175 -26 -23141
rect 8 -23175 20 -23141
rect -38 -23209 20 -23175
rect -38 -23243 -26 -23209
rect 8 -23243 20 -23209
rect -38 -23277 20 -23243
rect -38 -23311 -26 -23277
rect 8 -23311 20 -23277
rect -38 -23345 20 -23311
rect -38 -23379 -26 -23345
rect 8 -23379 20 -23345
rect -38 -23413 20 -23379
rect -38 -23447 -26 -23413
rect 8 -23447 20 -23413
rect -38 -23492 20 -23447
rect 260 -22937 318 -22892
rect 260 -22971 272 -22937
rect 306 -22971 318 -22937
rect 260 -23005 318 -22971
rect 260 -23039 272 -23005
rect 306 -23039 318 -23005
rect 260 -23073 318 -23039
rect 260 -23107 272 -23073
rect 306 -23107 318 -23073
rect 260 -23141 318 -23107
rect 260 -23175 272 -23141
rect 306 -23175 318 -23141
rect 260 -23209 318 -23175
rect 260 -23243 272 -23209
rect 306 -23243 318 -23209
rect 260 -23277 318 -23243
rect 260 -23311 272 -23277
rect 306 -23311 318 -23277
rect 260 -23345 318 -23311
rect 260 -23379 272 -23345
rect 306 -23379 318 -23345
rect 260 -23413 318 -23379
rect 260 -23447 272 -23413
rect 306 -23447 318 -23413
rect 260 -23492 318 -23447
rect 558 -22937 616 -22892
rect 558 -22971 570 -22937
rect 604 -22971 616 -22937
rect 558 -23005 616 -22971
rect 558 -23039 570 -23005
rect 604 -23039 616 -23005
rect 558 -23073 616 -23039
rect 558 -23107 570 -23073
rect 604 -23107 616 -23073
rect 558 -23141 616 -23107
rect 558 -23175 570 -23141
rect 604 -23175 616 -23141
rect 558 -23209 616 -23175
rect 558 -23243 570 -23209
rect 604 -23243 616 -23209
rect 558 -23277 616 -23243
rect 558 -23311 570 -23277
rect 604 -23311 616 -23277
rect 558 -23345 616 -23311
rect 558 -23379 570 -23345
rect 604 -23379 616 -23345
rect 558 -23413 616 -23379
rect 558 -23447 570 -23413
rect 604 -23447 616 -23413
rect 558 -23492 616 -23447
rect 856 -22937 914 -22892
rect 856 -22971 868 -22937
rect 902 -22971 914 -22937
rect 856 -23005 914 -22971
rect 856 -23039 868 -23005
rect 902 -23039 914 -23005
rect 856 -23073 914 -23039
rect 856 -23107 868 -23073
rect 902 -23107 914 -23073
rect 856 -23141 914 -23107
rect 856 -23175 868 -23141
rect 902 -23175 914 -23141
rect 856 -23209 914 -23175
rect 856 -23243 868 -23209
rect 902 -23243 914 -23209
rect 856 -23277 914 -23243
rect 856 -23311 868 -23277
rect 902 -23311 914 -23277
rect 856 -23345 914 -23311
rect 856 -23379 868 -23345
rect 902 -23379 914 -23345
rect 856 -23413 914 -23379
rect 856 -23447 868 -23413
rect 902 -23447 914 -23413
rect 2568 -22897 2580 -22863
rect 2614 -22897 2626 -22863
rect 2568 -22931 2626 -22897
rect 2568 -22965 2580 -22931
rect 2614 -22965 2626 -22931
rect 2568 -22999 2626 -22965
rect 2568 -23033 2580 -22999
rect 2614 -23033 2626 -22999
rect 2568 -23067 2626 -23033
rect 2568 -23101 2580 -23067
rect 2614 -23101 2626 -23067
rect 2568 -23135 2626 -23101
rect 2568 -23169 2580 -23135
rect 2614 -23169 2626 -23135
rect 2568 -23203 2626 -23169
rect 2568 -23237 2580 -23203
rect 2614 -23237 2626 -23203
rect 2568 -23271 2626 -23237
rect 2568 -23305 2580 -23271
rect 2614 -23305 2626 -23271
rect 2568 -23339 2626 -23305
rect 2568 -23373 2580 -23339
rect 2614 -23373 2626 -23339
rect 2568 -23418 2626 -23373
rect 3586 -22863 3644 -22818
rect 3586 -22897 3598 -22863
rect 3632 -22897 3644 -22863
rect 3586 -22931 3644 -22897
rect 3586 -22965 3598 -22931
rect 3632 -22965 3644 -22931
rect 3586 -22999 3644 -22965
rect 3586 -23033 3598 -22999
rect 3632 -23033 3644 -22999
rect 3586 -23067 3644 -23033
rect 3586 -23101 3598 -23067
rect 3632 -23101 3644 -23067
rect 3586 -23135 3644 -23101
rect 3586 -23169 3598 -23135
rect 3632 -23169 3644 -23135
rect 3586 -23203 3644 -23169
rect 3586 -23237 3598 -23203
rect 3632 -23237 3644 -23203
rect 3586 -23271 3644 -23237
rect 3586 -23305 3598 -23271
rect 3632 -23305 3644 -23271
rect 3586 -23339 3644 -23305
rect 3586 -23373 3598 -23339
rect 3632 -23373 3644 -23339
rect 3586 -23418 3644 -23373
rect 4604 -22863 4662 -22818
rect 4604 -22897 4616 -22863
rect 4650 -22897 4662 -22863
rect 4604 -22931 4662 -22897
rect 4604 -22965 4616 -22931
rect 4650 -22965 4662 -22931
rect 4604 -22999 4662 -22965
rect 4604 -23033 4616 -22999
rect 4650 -23033 4662 -22999
rect 4604 -23067 4662 -23033
rect 4604 -23101 4616 -23067
rect 4650 -23101 4662 -23067
rect 4604 -23135 4662 -23101
rect 4604 -23169 4616 -23135
rect 4650 -23169 4662 -23135
rect 4604 -23203 4662 -23169
rect 4604 -23237 4616 -23203
rect 4650 -23237 4662 -23203
rect 4604 -23271 4662 -23237
rect 4604 -23305 4616 -23271
rect 4650 -23305 4662 -23271
rect 4604 -23339 4662 -23305
rect 4604 -23373 4616 -23339
rect 4650 -23373 4662 -23339
rect 4604 -23418 4662 -23373
rect 5622 -22863 5680 -22818
rect 5622 -22897 5634 -22863
rect 5668 -22897 5680 -22863
rect 5622 -22931 5680 -22897
rect 5622 -22965 5634 -22931
rect 5668 -22965 5680 -22931
rect 5622 -22999 5680 -22965
rect 5622 -23033 5634 -22999
rect 5668 -23033 5680 -22999
rect 5622 -23067 5680 -23033
rect 5622 -23101 5634 -23067
rect 5668 -23101 5680 -23067
rect 5622 -23135 5680 -23101
rect 5622 -23169 5634 -23135
rect 5668 -23169 5680 -23135
rect 5622 -23203 5680 -23169
rect 5622 -23237 5634 -23203
rect 5668 -23237 5680 -23203
rect 5622 -23271 5680 -23237
rect 5622 -23305 5634 -23271
rect 5668 -23305 5680 -23271
rect 5622 -23339 5680 -23305
rect 5622 -23373 5634 -23339
rect 5668 -23373 5680 -23339
rect 5622 -23418 5680 -23373
rect 6640 -22863 6698 -22818
rect 6640 -22897 6652 -22863
rect 6686 -22897 6698 -22863
rect 6640 -22931 6698 -22897
rect 6640 -22965 6652 -22931
rect 6686 -22965 6698 -22931
rect 6640 -22999 6698 -22965
rect 6640 -23033 6652 -22999
rect 6686 -23033 6698 -22999
rect 6640 -23067 6698 -23033
rect 6640 -23101 6652 -23067
rect 6686 -23101 6698 -23067
rect 6640 -23135 6698 -23101
rect 6640 -23169 6652 -23135
rect 6686 -23169 6698 -23135
rect 6640 -23203 6698 -23169
rect 6640 -23237 6652 -23203
rect 6686 -23237 6698 -23203
rect 6640 -23271 6698 -23237
rect 6640 -23305 6652 -23271
rect 6686 -23305 6698 -23271
rect 6640 -23339 6698 -23305
rect 6640 -23373 6652 -23339
rect 6686 -23373 6698 -23339
rect 6640 -23418 6698 -23373
rect 7658 -22863 7716 -22818
rect 7658 -22897 7670 -22863
rect 7704 -22897 7716 -22863
rect 7658 -22931 7716 -22897
rect 7658 -22965 7670 -22931
rect 7704 -22965 7716 -22931
rect 7658 -22999 7716 -22965
rect 7658 -23033 7670 -22999
rect 7704 -23033 7716 -22999
rect 7658 -23067 7716 -23033
rect 7658 -23101 7670 -23067
rect 7704 -23101 7716 -23067
rect 7658 -23135 7716 -23101
rect 7658 -23169 7670 -23135
rect 7704 -23169 7716 -23135
rect 7658 -23203 7716 -23169
rect 7658 -23237 7670 -23203
rect 7704 -23237 7716 -23203
rect 7658 -23271 7716 -23237
rect 7658 -23305 7670 -23271
rect 7704 -23305 7716 -23271
rect 7658 -23339 7716 -23305
rect 7658 -23373 7670 -23339
rect 7704 -23373 7716 -23339
rect 7658 -23418 7716 -23373
rect 8676 -22863 8734 -22818
rect 8676 -22897 8688 -22863
rect 8722 -22897 8734 -22863
rect 8676 -22931 8734 -22897
rect 8676 -22965 8688 -22931
rect 8722 -22965 8734 -22931
rect 8676 -22999 8734 -22965
rect 8676 -23033 8688 -22999
rect 8722 -23033 8734 -22999
rect 8676 -23067 8734 -23033
rect 8676 -23101 8688 -23067
rect 8722 -23101 8734 -23067
rect 8676 -23135 8734 -23101
rect 8676 -23169 8688 -23135
rect 8722 -23169 8734 -23135
rect 8676 -23203 8734 -23169
rect 8676 -23237 8688 -23203
rect 8722 -23237 8734 -23203
rect 8676 -23271 8734 -23237
rect 8676 -23305 8688 -23271
rect 8722 -23305 8734 -23271
rect 8676 -23339 8734 -23305
rect 8676 -23373 8688 -23339
rect 8722 -23373 8734 -23339
rect 8676 -23418 8734 -23373
rect 9694 -22863 9752 -22818
rect 9694 -22897 9706 -22863
rect 9740 -22897 9752 -22863
rect 9694 -22931 9752 -22897
rect 9694 -22965 9706 -22931
rect 9740 -22965 9752 -22931
rect 9694 -22999 9752 -22965
rect 9694 -23033 9706 -22999
rect 9740 -23033 9752 -22999
rect 9694 -23067 9752 -23033
rect 9694 -23101 9706 -23067
rect 9740 -23101 9752 -23067
rect 9694 -23135 9752 -23101
rect 9694 -23169 9706 -23135
rect 9740 -23169 9752 -23135
rect 9694 -23203 9752 -23169
rect 9694 -23237 9706 -23203
rect 9740 -23237 9752 -23203
rect 9694 -23271 9752 -23237
rect 9694 -23305 9706 -23271
rect 9740 -23305 9752 -23271
rect 9694 -23339 9752 -23305
rect 9694 -23373 9706 -23339
rect 9740 -23373 9752 -23339
rect 9694 -23418 9752 -23373
rect 10712 -22863 10770 -22818
rect 10712 -22897 10724 -22863
rect 10758 -22897 10770 -22863
rect 10712 -22931 10770 -22897
rect 10712 -22965 10724 -22931
rect 10758 -22965 10770 -22931
rect 10712 -22999 10770 -22965
rect 10712 -23033 10724 -22999
rect 10758 -23033 10770 -22999
rect 10712 -23067 10770 -23033
rect 10712 -23101 10724 -23067
rect 10758 -23101 10770 -23067
rect 10712 -23135 10770 -23101
rect 10712 -23169 10724 -23135
rect 10758 -23169 10770 -23135
rect 10712 -23203 10770 -23169
rect 10712 -23237 10724 -23203
rect 10758 -23237 10770 -23203
rect 10712 -23271 10770 -23237
rect 10712 -23305 10724 -23271
rect 10758 -23305 10770 -23271
rect 10712 -23339 10770 -23305
rect 10712 -23373 10724 -23339
rect 10758 -23373 10770 -23339
rect 10712 -23418 10770 -23373
rect 11730 -22863 11788 -22818
rect 11730 -22897 11742 -22863
rect 11776 -22897 11788 -22863
rect 11730 -22931 11788 -22897
rect 11730 -22965 11742 -22931
rect 11776 -22965 11788 -22931
rect 11730 -22999 11788 -22965
rect 11730 -23033 11742 -22999
rect 11776 -23033 11788 -22999
rect 11730 -23067 11788 -23033
rect 11730 -23101 11742 -23067
rect 11776 -23101 11788 -23067
rect 11730 -23135 11788 -23101
rect 11730 -23169 11742 -23135
rect 11776 -23169 11788 -23135
rect 11730 -23203 11788 -23169
rect 11730 -23237 11742 -23203
rect 11776 -23237 11788 -23203
rect 11730 -23271 11788 -23237
rect 11730 -23305 11742 -23271
rect 11776 -23305 11788 -23271
rect 11730 -23339 11788 -23305
rect 11730 -23373 11742 -23339
rect 11776 -23373 11788 -23339
rect 11730 -23418 11788 -23373
rect 12748 -22863 12806 -22818
rect 12748 -22897 12760 -22863
rect 12794 -22897 12806 -22863
rect 12748 -22931 12806 -22897
rect 12748 -22965 12760 -22931
rect 12794 -22965 12806 -22931
rect 12748 -22999 12806 -22965
rect 12748 -23033 12760 -22999
rect 12794 -23033 12806 -22999
rect 12748 -23067 12806 -23033
rect 12748 -23101 12760 -23067
rect 12794 -23101 12806 -23067
rect 12748 -23135 12806 -23101
rect 12748 -23169 12760 -23135
rect 12794 -23169 12806 -23135
rect 12748 -23203 12806 -23169
rect 12748 -23237 12760 -23203
rect 12794 -23237 12806 -23203
rect 12748 -23271 12806 -23237
rect 12748 -23305 12760 -23271
rect 12794 -23305 12806 -23271
rect 12748 -23339 12806 -23305
rect 12748 -23373 12760 -23339
rect 12794 -23373 12806 -23339
rect 12748 -23418 12806 -23373
rect 13766 -22863 13824 -22818
rect 13766 -22897 13778 -22863
rect 13812 -22897 13824 -22863
rect 13766 -22931 13824 -22897
rect 13766 -22965 13778 -22931
rect 13812 -22965 13824 -22931
rect 13766 -22999 13824 -22965
rect 13766 -23033 13778 -22999
rect 13812 -23033 13824 -22999
rect 13766 -23067 13824 -23033
rect 13766 -23101 13778 -23067
rect 13812 -23101 13824 -23067
rect 13766 -23135 13824 -23101
rect 13766 -23169 13778 -23135
rect 13812 -23169 13824 -23135
rect 13766 -23203 13824 -23169
rect 13766 -23237 13778 -23203
rect 13812 -23237 13824 -23203
rect 13766 -23271 13824 -23237
rect 13766 -23305 13778 -23271
rect 13812 -23305 13824 -23271
rect 13766 -23339 13824 -23305
rect 13766 -23373 13778 -23339
rect 13812 -23373 13824 -23339
rect 13766 -23418 13824 -23373
rect 14784 -22863 14842 -22818
rect 14784 -22897 14796 -22863
rect 14830 -22897 14842 -22863
rect 14784 -22931 14842 -22897
rect 14784 -22965 14796 -22931
rect 14830 -22965 14842 -22931
rect 14784 -22999 14842 -22965
rect 14784 -23033 14796 -22999
rect 14830 -23033 14842 -22999
rect 14784 -23067 14842 -23033
rect 14784 -23101 14796 -23067
rect 14830 -23101 14842 -23067
rect 14784 -23135 14842 -23101
rect 14784 -23169 14796 -23135
rect 14830 -23169 14842 -23135
rect 14784 -23203 14842 -23169
rect 14784 -23237 14796 -23203
rect 14830 -23237 14842 -23203
rect 14784 -23271 14842 -23237
rect 14784 -23305 14796 -23271
rect 14830 -23305 14842 -23271
rect 14784 -23339 14842 -23305
rect 14784 -23373 14796 -23339
rect 14830 -23373 14842 -23339
rect 14784 -23418 14842 -23373
rect 15802 -22863 15860 -22818
rect 15802 -22897 15814 -22863
rect 15848 -22897 15860 -22863
rect 15802 -22931 15860 -22897
rect 15802 -22965 15814 -22931
rect 15848 -22965 15860 -22931
rect 15802 -22999 15860 -22965
rect 15802 -23033 15814 -22999
rect 15848 -23033 15860 -22999
rect 15802 -23067 15860 -23033
rect 15802 -23101 15814 -23067
rect 15848 -23101 15860 -23067
rect 15802 -23135 15860 -23101
rect 15802 -23169 15814 -23135
rect 15848 -23169 15860 -23135
rect 15802 -23203 15860 -23169
rect 15802 -23237 15814 -23203
rect 15848 -23237 15860 -23203
rect 15802 -23271 15860 -23237
rect 15802 -23305 15814 -23271
rect 15848 -23305 15860 -23271
rect 15802 -23339 15860 -23305
rect 15802 -23373 15814 -23339
rect 15848 -23373 15860 -23339
rect 15802 -23418 15860 -23373
rect 16820 -22863 16878 -22818
rect 16820 -22897 16832 -22863
rect 16866 -22897 16878 -22863
rect 16820 -22931 16878 -22897
rect 16820 -22965 16832 -22931
rect 16866 -22965 16878 -22931
rect 16820 -22999 16878 -22965
rect 16820 -23033 16832 -22999
rect 16866 -23033 16878 -22999
rect 16820 -23067 16878 -23033
rect 16820 -23101 16832 -23067
rect 16866 -23101 16878 -23067
rect 16820 -23135 16878 -23101
rect 16820 -23169 16832 -23135
rect 16866 -23169 16878 -23135
rect 16820 -23203 16878 -23169
rect 16820 -23237 16832 -23203
rect 16866 -23237 16878 -23203
rect 16820 -23271 16878 -23237
rect 16820 -23305 16832 -23271
rect 16866 -23305 16878 -23271
rect 16820 -23339 16878 -23305
rect 16820 -23373 16832 -23339
rect 16866 -23373 16878 -23339
rect 16820 -23418 16878 -23373
rect 17838 -22863 17896 -22818
rect 17838 -22897 17850 -22863
rect 17884 -22897 17896 -22863
rect 17838 -22931 17896 -22897
rect 17838 -22965 17850 -22931
rect 17884 -22965 17896 -22931
rect 17838 -22999 17896 -22965
rect 17838 -23033 17850 -22999
rect 17884 -23033 17896 -22999
rect 17838 -23067 17896 -23033
rect 17838 -23101 17850 -23067
rect 17884 -23101 17896 -23067
rect 17838 -23135 17896 -23101
rect 17838 -23169 17850 -23135
rect 17884 -23169 17896 -23135
rect 17838 -23203 17896 -23169
rect 17838 -23237 17850 -23203
rect 17884 -23237 17896 -23203
rect 17838 -23271 17896 -23237
rect 17838 -23305 17850 -23271
rect 17884 -23305 17896 -23271
rect 17838 -23339 17896 -23305
rect 17838 -23373 17850 -23339
rect 17884 -23373 17896 -23339
rect 17838 -23418 17896 -23373
rect 18856 -22863 18914 -22818
rect 18856 -22897 18868 -22863
rect 18902 -22897 18914 -22863
rect 18856 -22931 18914 -22897
rect 18856 -22965 18868 -22931
rect 18902 -22965 18914 -22931
rect 18856 -22999 18914 -22965
rect 18856 -23033 18868 -22999
rect 18902 -23033 18914 -22999
rect 18856 -23067 18914 -23033
rect 18856 -23101 18868 -23067
rect 18902 -23101 18914 -23067
rect 18856 -23135 18914 -23101
rect 18856 -23169 18868 -23135
rect 18902 -23169 18914 -23135
rect 18856 -23203 18914 -23169
rect 18856 -23237 18868 -23203
rect 18902 -23237 18914 -23203
rect 18856 -23271 18914 -23237
rect 18856 -23305 18868 -23271
rect 18902 -23305 18914 -23271
rect 18856 -23339 18914 -23305
rect 18856 -23373 18868 -23339
rect 18902 -23373 18914 -23339
rect 18856 -23418 18914 -23373
rect 19874 -22863 19932 -22818
rect 19874 -22897 19886 -22863
rect 19920 -22897 19932 -22863
rect 19874 -22931 19932 -22897
rect 19874 -22965 19886 -22931
rect 19920 -22965 19932 -22931
rect 19874 -22999 19932 -22965
rect 19874 -23033 19886 -22999
rect 19920 -23033 19932 -22999
rect 19874 -23067 19932 -23033
rect 19874 -23101 19886 -23067
rect 19920 -23101 19932 -23067
rect 19874 -23135 19932 -23101
rect 19874 -23169 19886 -23135
rect 19920 -23169 19932 -23135
rect 19874 -23203 19932 -23169
rect 19874 -23237 19886 -23203
rect 19920 -23237 19932 -23203
rect 19874 -23271 19932 -23237
rect 19874 -23305 19886 -23271
rect 19920 -23305 19932 -23271
rect 19874 -23339 19932 -23305
rect 19874 -23373 19886 -23339
rect 19920 -23373 19932 -23339
rect 19874 -23418 19932 -23373
rect 20892 -22863 20950 -22818
rect 20892 -22897 20904 -22863
rect 20938 -22897 20950 -22863
rect 20892 -22931 20950 -22897
rect 20892 -22965 20904 -22931
rect 20938 -22965 20950 -22931
rect 20892 -22999 20950 -22965
rect 20892 -23033 20904 -22999
rect 20938 -23033 20950 -22999
rect 20892 -23067 20950 -23033
rect 20892 -23101 20904 -23067
rect 20938 -23101 20950 -23067
rect 20892 -23135 20950 -23101
rect 20892 -23169 20904 -23135
rect 20938 -23169 20950 -23135
rect 20892 -23203 20950 -23169
rect 20892 -23237 20904 -23203
rect 20938 -23237 20950 -23203
rect 20892 -23271 20950 -23237
rect 20892 -23305 20904 -23271
rect 20938 -23305 20950 -23271
rect 20892 -23339 20950 -23305
rect 20892 -23373 20904 -23339
rect 20938 -23373 20950 -23339
rect 20892 -23418 20950 -23373
rect 21910 -22863 21968 -22818
rect 21910 -22897 21922 -22863
rect 21956 -22897 21968 -22863
rect 21910 -22931 21968 -22897
rect 21910 -22965 21922 -22931
rect 21956 -22965 21968 -22931
rect 21910 -22999 21968 -22965
rect 21910 -23033 21922 -22999
rect 21956 -23033 21968 -22999
rect 21910 -23067 21968 -23033
rect 21910 -23101 21922 -23067
rect 21956 -23101 21968 -23067
rect 21910 -23135 21968 -23101
rect 21910 -23169 21922 -23135
rect 21956 -23169 21968 -23135
rect 21910 -23203 21968 -23169
rect 21910 -23237 21922 -23203
rect 21956 -23237 21968 -23203
rect 21910 -23271 21968 -23237
rect 21910 -23305 21922 -23271
rect 21956 -23305 21968 -23271
rect 21910 -23339 21968 -23305
rect 21910 -23373 21922 -23339
rect 21956 -23373 21968 -23339
rect 21910 -23418 21968 -23373
rect 22928 -22863 22986 -22818
rect 22928 -22897 22940 -22863
rect 22974 -22897 22986 -22863
rect 22928 -22931 22986 -22897
rect 22928 -22965 22940 -22931
rect 22974 -22965 22986 -22931
rect 22928 -22999 22986 -22965
rect 22928 -23033 22940 -22999
rect 22974 -23033 22986 -22999
rect 22928 -23067 22986 -23033
rect 22928 -23101 22940 -23067
rect 22974 -23101 22986 -23067
rect 22928 -23135 22986 -23101
rect 22928 -23169 22940 -23135
rect 22974 -23169 22986 -23135
rect 22928 -23203 22986 -23169
rect 22928 -23237 22940 -23203
rect 22974 -23237 22986 -23203
rect 22928 -23271 22986 -23237
rect 22928 -23305 22940 -23271
rect 22974 -23305 22986 -23271
rect 22928 -23339 22986 -23305
rect 22928 -23373 22940 -23339
rect 22974 -23373 22986 -23339
rect 22928 -23418 22986 -23373
rect 856 -23492 914 -23447
rect -9417 -24050 -9359 -24005
rect -9417 -24084 -9405 -24050
rect -9371 -24084 -9359 -24050
rect -9417 -24118 -9359 -24084
rect -9417 -24152 -9405 -24118
rect -9371 -24152 -9359 -24118
rect -9417 -24186 -9359 -24152
rect -9417 -24220 -9405 -24186
rect -9371 -24220 -9359 -24186
rect -9417 -24254 -9359 -24220
rect -9417 -24288 -9405 -24254
rect -9371 -24288 -9359 -24254
rect -9417 -24322 -9359 -24288
rect -9417 -24356 -9405 -24322
rect -9371 -24356 -9359 -24322
rect -9417 -24390 -9359 -24356
rect -9417 -24424 -9405 -24390
rect -9371 -24424 -9359 -24390
rect -9417 -24458 -9359 -24424
rect -9417 -24492 -9405 -24458
rect -9371 -24492 -9359 -24458
rect -9417 -24526 -9359 -24492
rect -9417 -24560 -9405 -24526
rect -9371 -24560 -9359 -24526
rect -9417 -24605 -9359 -24560
rect -8399 -24050 -8341 -24005
rect -8399 -24084 -8387 -24050
rect -8353 -24084 -8341 -24050
rect -8399 -24118 -8341 -24084
rect -8399 -24152 -8387 -24118
rect -8353 -24152 -8341 -24118
rect -8399 -24186 -8341 -24152
rect -8399 -24220 -8387 -24186
rect -8353 -24220 -8341 -24186
rect -8399 -24254 -8341 -24220
rect -8399 -24288 -8387 -24254
rect -8353 -24288 -8341 -24254
rect -8399 -24322 -8341 -24288
rect -8399 -24356 -8387 -24322
rect -8353 -24356 -8341 -24322
rect -8399 -24390 -8341 -24356
rect -8399 -24424 -8387 -24390
rect -8353 -24424 -8341 -24390
rect -8399 -24458 -8341 -24424
rect -8399 -24492 -8387 -24458
rect -8353 -24492 -8341 -24458
rect -8399 -24526 -8341 -24492
rect -8399 -24560 -8387 -24526
rect -8353 -24560 -8341 -24526
rect -8399 -24605 -8341 -24560
rect -7381 -24050 -7323 -24005
rect -7381 -24084 -7369 -24050
rect -7335 -24084 -7323 -24050
rect -7381 -24118 -7323 -24084
rect -7381 -24152 -7369 -24118
rect -7335 -24152 -7323 -24118
rect -7381 -24186 -7323 -24152
rect -7381 -24220 -7369 -24186
rect -7335 -24220 -7323 -24186
rect -7381 -24254 -7323 -24220
rect -7381 -24288 -7369 -24254
rect -7335 -24288 -7323 -24254
rect -7381 -24322 -7323 -24288
rect -7381 -24356 -7369 -24322
rect -7335 -24356 -7323 -24322
rect -7381 -24390 -7323 -24356
rect -7381 -24424 -7369 -24390
rect -7335 -24424 -7323 -24390
rect -7381 -24458 -7323 -24424
rect -7381 -24492 -7369 -24458
rect -7335 -24492 -7323 -24458
rect -7381 -24526 -7323 -24492
rect -7381 -24560 -7369 -24526
rect -7335 -24560 -7323 -24526
rect -7381 -24605 -7323 -24560
rect -6363 -24050 -6305 -24005
rect -6363 -24084 -6351 -24050
rect -6317 -24084 -6305 -24050
rect -6363 -24118 -6305 -24084
rect -6363 -24152 -6351 -24118
rect -6317 -24152 -6305 -24118
rect -6363 -24186 -6305 -24152
rect -6363 -24220 -6351 -24186
rect -6317 -24220 -6305 -24186
rect -6363 -24254 -6305 -24220
rect -6363 -24288 -6351 -24254
rect -6317 -24288 -6305 -24254
rect -6363 -24322 -6305 -24288
rect -6363 -24356 -6351 -24322
rect -6317 -24356 -6305 -24322
rect -6363 -24390 -6305 -24356
rect -6363 -24424 -6351 -24390
rect -6317 -24424 -6305 -24390
rect -6363 -24458 -6305 -24424
rect -6363 -24492 -6351 -24458
rect -6317 -24492 -6305 -24458
rect -6363 -24526 -6305 -24492
rect -6363 -24560 -6351 -24526
rect -6317 -24560 -6305 -24526
rect -6363 -24605 -6305 -24560
rect -5345 -24050 -5287 -24005
rect -5345 -24084 -5333 -24050
rect -5299 -24084 -5287 -24050
rect -5345 -24118 -5287 -24084
rect -5345 -24152 -5333 -24118
rect -5299 -24152 -5287 -24118
rect -5345 -24186 -5287 -24152
rect -5345 -24220 -5333 -24186
rect -5299 -24220 -5287 -24186
rect -5345 -24254 -5287 -24220
rect -5345 -24288 -5333 -24254
rect -5299 -24288 -5287 -24254
rect -5345 -24322 -5287 -24288
rect -5345 -24356 -5333 -24322
rect -5299 -24356 -5287 -24322
rect -5345 -24390 -5287 -24356
rect -5345 -24424 -5333 -24390
rect -5299 -24424 -5287 -24390
rect -5345 -24458 -5287 -24424
rect -5345 -24492 -5333 -24458
rect -5299 -24492 -5287 -24458
rect -5345 -24526 -5287 -24492
rect -5345 -24560 -5333 -24526
rect -5299 -24560 -5287 -24526
rect -5345 -24605 -5287 -24560
rect -4327 -24050 -4269 -24005
rect -4327 -24084 -4315 -24050
rect -4281 -24084 -4269 -24050
rect -4327 -24118 -4269 -24084
rect -4327 -24152 -4315 -24118
rect -4281 -24152 -4269 -24118
rect -4327 -24186 -4269 -24152
rect -4327 -24220 -4315 -24186
rect -4281 -24220 -4269 -24186
rect -4327 -24254 -4269 -24220
rect -4327 -24288 -4315 -24254
rect -4281 -24288 -4269 -24254
rect -4327 -24322 -4269 -24288
rect -4327 -24356 -4315 -24322
rect -4281 -24356 -4269 -24322
rect -4327 -24390 -4269 -24356
rect -4327 -24424 -4315 -24390
rect -4281 -24424 -4269 -24390
rect -4327 -24458 -4269 -24424
rect -4327 -24492 -4315 -24458
rect -4281 -24492 -4269 -24458
rect -4327 -24526 -4269 -24492
rect -4327 -24560 -4315 -24526
rect -4281 -24560 -4269 -24526
rect -4327 -24605 -4269 -24560
rect -3309 -24050 -3251 -24005
rect -3309 -24084 -3297 -24050
rect -3263 -24084 -3251 -24050
rect -3309 -24118 -3251 -24084
rect -3309 -24152 -3297 -24118
rect -3263 -24152 -3251 -24118
rect -3309 -24186 -3251 -24152
rect -3309 -24220 -3297 -24186
rect -3263 -24220 -3251 -24186
rect -3309 -24254 -3251 -24220
rect -3309 -24288 -3297 -24254
rect -3263 -24288 -3251 -24254
rect -3309 -24322 -3251 -24288
rect -3309 -24356 -3297 -24322
rect -3263 -24356 -3251 -24322
rect -3309 -24390 -3251 -24356
rect -3309 -24424 -3297 -24390
rect -3263 -24424 -3251 -24390
rect -3309 -24458 -3251 -24424
rect -3309 -24492 -3297 -24458
rect -3263 -24492 -3251 -24458
rect -3309 -24526 -3251 -24492
rect -3309 -24560 -3297 -24526
rect -3263 -24560 -3251 -24526
rect -3309 -24605 -3251 -24560
rect -2424 -24049 -2366 -24004
rect -2424 -24083 -2412 -24049
rect -2378 -24083 -2366 -24049
rect -2424 -24117 -2366 -24083
rect -2424 -24151 -2412 -24117
rect -2378 -24151 -2366 -24117
rect -2424 -24185 -2366 -24151
rect -2424 -24219 -2412 -24185
rect -2378 -24219 -2366 -24185
rect -2424 -24253 -2366 -24219
rect -2424 -24287 -2412 -24253
rect -2378 -24287 -2366 -24253
rect -2424 -24321 -2366 -24287
rect -2424 -24355 -2412 -24321
rect -2378 -24355 -2366 -24321
rect -2424 -24389 -2366 -24355
rect -2424 -24423 -2412 -24389
rect -2378 -24423 -2366 -24389
rect -2424 -24457 -2366 -24423
rect -2424 -24491 -2412 -24457
rect -2378 -24491 -2366 -24457
rect -2424 -24525 -2366 -24491
rect -2424 -24559 -2412 -24525
rect -2378 -24559 -2366 -24525
rect -2424 -24604 -2366 -24559
rect -2126 -24049 -2068 -24004
rect -2126 -24083 -2114 -24049
rect -2080 -24083 -2068 -24049
rect -2126 -24117 -2068 -24083
rect -2126 -24151 -2114 -24117
rect -2080 -24151 -2068 -24117
rect -2126 -24185 -2068 -24151
rect -2126 -24219 -2114 -24185
rect -2080 -24219 -2068 -24185
rect -2126 -24253 -2068 -24219
rect -2126 -24287 -2114 -24253
rect -2080 -24287 -2068 -24253
rect -2126 -24321 -2068 -24287
rect -2126 -24355 -2114 -24321
rect -2080 -24355 -2068 -24321
rect -2126 -24389 -2068 -24355
rect -2126 -24423 -2114 -24389
rect -2080 -24423 -2068 -24389
rect -2126 -24457 -2068 -24423
rect -2126 -24491 -2114 -24457
rect -2080 -24491 -2068 -24457
rect -2126 -24525 -2068 -24491
rect -2126 -24559 -2114 -24525
rect -2080 -24559 -2068 -24525
rect -2126 -24604 -2068 -24559
rect -1828 -24049 -1770 -24004
rect -1828 -24083 -1816 -24049
rect -1782 -24083 -1770 -24049
rect -1828 -24117 -1770 -24083
rect -1828 -24151 -1816 -24117
rect -1782 -24151 -1770 -24117
rect -1828 -24185 -1770 -24151
rect -1828 -24219 -1816 -24185
rect -1782 -24219 -1770 -24185
rect -1828 -24253 -1770 -24219
rect -1828 -24287 -1816 -24253
rect -1782 -24287 -1770 -24253
rect -1828 -24321 -1770 -24287
rect -1828 -24355 -1816 -24321
rect -1782 -24355 -1770 -24321
rect -1828 -24389 -1770 -24355
rect -1828 -24423 -1816 -24389
rect -1782 -24423 -1770 -24389
rect -1828 -24457 -1770 -24423
rect -1828 -24491 -1816 -24457
rect -1782 -24491 -1770 -24457
rect -1828 -24525 -1770 -24491
rect -1828 -24559 -1816 -24525
rect -1782 -24559 -1770 -24525
rect -1828 -24604 -1770 -24559
rect -1530 -24049 -1472 -24004
rect -1530 -24083 -1518 -24049
rect -1484 -24083 -1472 -24049
rect -1530 -24117 -1472 -24083
rect -1530 -24151 -1518 -24117
rect -1484 -24151 -1472 -24117
rect -1530 -24185 -1472 -24151
rect -1530 -24219 -1518 -24185
rect -1484 -24219 -1472 -24185
rect -1530 -24253 -1472 -24219
rect -1530 -24287 -1518 -24253
rect -1484 -24287 -1472 -24253
rect -1530 -24321 -1472 -24287
rect -1530 -24355 -1518 -24321
rect -1484 -24355 -1472 -24321
rect -1530 -24389 -1472 -24355
rect -1530 -24423 -1518 -24389
rect -1484 -24423 -1472 -24389
rect -1530 -24457 -1472 -24423
rect -1530 -24491 -1518 -24457
rect -1484 -24491 -1472 -24457
rect -1530 -24525 -1472 -24491
rect -1530 -24559 -1518 -24525
rect -1484 -24559 -1472 -24525
rect -1530 -24604 -1472 -24559
rect -1232 -24049 -1174 -24004
rect -1232 -24083 -1220 -24049
rect -1186 -24083 -1174 -24049
rect -1232 -24117 -1174 -24083
rect -1232 -24151 -1220 -24117
rect -1186 -24151 -1174 -24117
rect -1232 -24185 -1174 -24151
rect -1232 -24219 -1220 -24185
rect -1186 -24219 -1174 -24185
rect -1232 -24253 -1174 -24219
rect -1232 -24287 -1220 -24253
rect -1186 -24287 -1174 -24253
rect -1232 -24321 -1174 -24287
rect -1232 -24355 -1220 -24321
rect -1186 -24355 -1174 -24321
rect -1232 -24389 -1174 -24355
rect -1232 -24423 -1220 -24389
rect -1186 -24423 -1174 -24389
rect -1232 -24457 -1174 -24423
rect -1232 -24491 -1220 -24457
rect -1186 -24491 -1174 -24457
rect -1232 -24525 -1174 -24491
rect -1232 -24559 -1220 -24525
rect -1186 -24559 -1174 -24525
rect -1232 -24604 -1174 -24559
rect -934 -24049 -876 -24004
rect -934 -24083 -922 -24049
rect -888 -24083 -876 -24049
rect -934 -24117 -876 -24083
rect -934 -24151 -922 -24117
rect -888 -24151 -876 -24117
rect -934 -24185 -876 -24151
rect -934 -24219 -922 -24185
rect -888 -24219 -876 -24185
rect -934 -24253 -876 -24219
rect -934 -24287 -922 -24253
rect -888 -24287 -876 -24253
rect -934 -24321 -876 -24287
rect -934 -24355 -922 -24321
rect -888 -24355 -876 -24321
rect -934 -24389 -876 -24355
rect -934 -24423 -922 -24389
rect -888 -24423 -876 -24389
rect -934 -24457 -876 -24423
rect -934 -24491 -922 -24457
rect -888 -24491 -876 -24457
rect -934 -24525 -876 -24491
rect -934 -24559 -922 -24525
rect -888 -24559 -876 -24525
rect -934 -24604 -876 -24559
rect -636 -24049 -578 -24004
rect -636 -24083 -624 -24049
rect -590 -24083 -578 -24049
rect -636 -24117 -578 -24083
rect -636 -24151 -624 -24117
rect -590 -24151 -578 -24117
rect -636 -24185 -578 -24151
rect -636 -24219 -624 -24185
rect -590 -24219 -578 -24185
rect -636 -24253 -578 -24219
rect -636 -24287 -624 -24253
rect -590 -24287 -578 -24253
rect -636 -24321 -578 -24287
rect -636 -24355 -624 -24321
rect -590 -24355 -578 -24321
rect -636 -24389 -578 -24355
rect -636 -24423 -624 -24389
rect -590 -24423 -578 -24389
rect -636 -24457 -578 -24423
rect -636 -24491 -624 -24457
rect -590 -24491 -578 -24457
rect -636 -24525 -578 -24491
rect -636 -24559 -624 -24525
rect -590 -24559 -578 -24525
rect -636 -24604 -578 -24559
rect -338 -24049 -280 -24004
rect -338 -24083 -326 -24049
rect -292 -24083 -280 -24049
rect -338 -24117 -280 -24083
rect -338 -24151 -326 -24117
rect -292 -24151 -280 -24117
rect -338 -24185 -280 -24151
rect -338 -24219 -326 -24185
rect -292 -24219 -280 -24185
rect -338 -24253 -280 -24219
rect -338 -24287 -326 -24253
rect -292 -24287 -280 -24253
rect -338 -24321 -280 -24287
rect -338 -24355 -326 -24321
rect -292 -24355 -280 -24321
rect -338 -24389 -280 -24355
rect -338 -24423 -326 -24389
rect -292 -24423 -280 -24389
rect -338 -24457 -280 -24423
rect -338 -24491 -326 -24457
rect -292 -24491 -280 -24457
rect -338 -24525 -280 -24491
rect -338 -24559 -326 -24525
rect -292 -24559 -280 -24525
rect -338 -24604 -280 -24559
rect -40 -24049 18 -24004
rect -40 -24083 -28 -24049
rect 6 -24083 18 -24049
rect -40 -24117 18 -24083
rect -40 -24151 -28 -24117
rect 6 -24151 18 -24117
rect -40 -24185 18 -24151
rect -40 -24219 -28 -24185
rect 6 -24219 18 -24185
rect -40 -24253 18 -24219
rect -40 -24287 -28 -24253
rect 6 -24287 18 -24253
rect -40 -24321 18 -24287
rect -40 -24355 -28 -24321
rect 6 -24355 18 -24321
rect -40 -24389 18 -24355
rect -40 -24423 -28 -24389
rect 6 -24423 18 -24389
rect -40 -24457 18 -24423
rect -40 -24491 -28 -24457
rect 6 -24491 18 -24457
rect -40 -24525 18 -24491
rect -40 -24559 -28 -24525
rect 6 -24559 18 -24525
rect -40 -24604 18 -24559
rect 258 -24049 316 -24004
rect 258 -24083 270 -24049
rect 304 -24083 316 -24049
rect 258 -24117 316 -24083
rect 258 -24151 270 -24117
rect 304 -24151 316 -24117
rect 258 -24185 316 -24151
rect 258 -24219 270 -24185
rect 304 -24219 316 -24185
rect 258 -24253 316 -24219
rect 258 -24287 270 -24253
rect 304 -24287 316 -24253
rect 258 -24321 316 -24287
rect 258 -24355 270 -24321
rect 304 -24355 316 -24321
rect 258 -24389 316 -24355
rect 258 -24423 270 -24389
rect 304 -24423 316 -24389
rect 258 -24457 316 -24423
rect 258 -24491 270 -24457
rect 304 -24491 316 -24457
rect 258 -24525 316 -24491
rect 258 -24559 270 -24525
rect 304 -24559 316 -24525
rect 258 -24604 316 -24559
rect 556 -24049 614 -24004
rect 556 -24083 568 -24049
rect 602 -24083 614 -24049
rect 556 -24117 614 -24083
rect 556 -24151 568 -24117
rect 602 -24151 614 -24117
rect 556 -24185 614 -24151
rect 556 -24219 568 -24185
rect 602 -24219 614 -24185
rect 556 -24253 614 -24219
rect 556 -24287 568 -24253
rect 602 -24287 614 -24253
rect 556 -24321 614 -24287
rect 556 -24355 568 -24321
rect 602 -24355 614 -24321
rect 556 -24389 614 -24355
rect 556 -24423 568 -24389
rect 602 -24423 614 -24389
rect 556 -24457 614 -24423
rect 556 -24491 568 -24457
rect 602 -24491 614 -24457
rect 556 -24525 614 -24491
rect 556 -24559 568 -24525
rect 602 -24559 614 -24525
rect 556 -24604 614 -24559
rect 854 -24049 912 -24004
rect 854 -24083 866 -24049
rect 900 -24083 912 -24049
rect 854 -24117 912 -24083
rect 854 -24151 866 -24117
rect 900 -24151 912 -24117
rect 854 -24185 912 -24151
rect 854 -24219 866 -24185
rect 900 -24219 912 -24185
rect 854 -24253 912 -24219
rect 854 -24287 866 -24253
rect 900 -24287 912 -24253
rect 854 -24321 912 -24287
rect 854 -24355 866 -24321
rect 900 -24355 912 -24321
rect 854 -24389 912 -24355
rect 854 -24423 866 -24389
rect 900 -24423 912 -24389
rect 854 -24457 912 -24423
rect 854 -24491 866 -24457
rect 900 -24491 912 -24457
rect 854 -24525 912 -24491
rect 854 -24559 866 -24525
rect 900 -24559 912 -24525
rect 854 -24604 912 -24559
rect 2568 -24097 2626 -24052
rect 2568 -24131 2580 -24097
rect 2614 -24131 2626 -24097
rect 2568 -24165 2626 -24131
rect 2568 -24199 2580 -24165
rect 2614 -24199 2626 -24165
rect 2568 -24233 2626 -24199
rect 2568 -24267 2580 -24233
rect 2614 -24267 2626 -24233
rect 2568 -24301 2626 -24267
rect 2568 -24335 2580 -24301
rect 2614 -24335 2626 -24301
rect 2568 -24369 2626 -24335
rect 2568 -24403 2580 -24369
rect 2614 -24403 2626 -24369
rect 2568 -24437 2626 -24403
rect 2568 -24471 2580 -24437
rect 2614 -24471 2626 -24437
rect 2568 -24505 2626 -24471
rect 2568 -24539 2580 -24505
rect 2614 -24539 2626 -24505
rect 2568 -24573 2626 -24539
rect 2568 -24607 2580 -24573
rect 2614 -24607 2626 -24573
rect 2568 -24652 2626 -24607
rect 3586 -24097 3644 -24052
rect 3586 -24131 3598 -24097
rect 3632 -24131 3644 -24097
rect 3586 -24165 3644 -24131
rect 3586 -24199 3598 -24165
rect 3632 -24199 3644 -24165
rect 3586 -24233 3644 -24199
rect 3586 -24267 3598 -24233
rect 3632 -24267 3644 -24233
rect 3586 -24301 3644 -24267
rect 3586 -24335 3598 -24301
rect 3632 -24335 3644 -24301
rect 3586 -24369 3644 -24335
rect 3586 -24403 3598 -24369
rect 3632 -24403 3644 -24369
rect 3586 -24437 3644 -24403
rect 3586 -24471 3598 -24437
rect 3632 -24471 3644 -24437
rect 3586 -24505 3644 -24471
rect 3586 -24539 3598 -24505
rect 3632 -24539 3644 -24505
rect 3586 -24573 3644 -24539
rect 3586 -24607 3598 -24573
rect 3632 -24607 3644 -24573
rect 3586 -24652 3644 -24607
rect 4604 -24097 4662 -24052
rect 4604 -24131 4616 -24097
rect 4650 -24131 4662 -24097
rect 4604 -24165 4662 -24131
rect 4604 -24199 4616 -24165
rect 4650 -24199 4662 -24165
rect 4604 -24233 4662 -24199
rect 4604 -24267 4616 -24233
rect 4650 -24267 4662 -24233
rect 4604 -24301 4662 -24267
rect 4604 -24335 4616 -24301
rect 4650 -24335 4662 -24301
rect 4604 -24369 4662 -24335
rect 4604 -24403 4616 -24369
rect 4650 -24403 4662 -24369
rect 4604 -24437 4662 -24403
rect 4604 -24471 4616 -24437
rect 4650 -24471 4662 -24437
rect 4604 -24505 4662 -24471
rect 4604 -24539 4616 -24505
rect 4650 -24539 4662 -24505
rect 4604 -24573 4662 -24539
rect 4604 -24607 4616 -24573
rect 4650 -24607 4662 -24573
rect 4604 -24652 4662 -24607
rect 5622 -24097 5680 -24052
rect 5622 -24131 5634 -24097
rect 5668 -24131 5680 -24097
rect 5622 -24165 5680 -24131
rect 5622 -24199 5634 -24165
rect 5668 -24199 5680 -24165
rect 5622 -24233 5680 -24199
rect 5622 -24267 5634 -24233
rect 5668 -24267 5680 -24233
rect 5622 -24301 5680 -24267
rect 5622 -24335 5634 -24301
rect 5668 -24335 5680 -24301
rect 5622 -24369 5680 -24335
rect 5622 -24403 5634 -24369
rect 5668 -24403 5680 -24369
rect 5622 -24437 5680 -24403
rect 5622 -24471 5634 -24437
rect 5668 -24471 5680 -24437
rect 5622 -24505 5680 -24471
rect 5622 -24539 5634 -24505
rect 5668 -24539 5680 -24505
rect 5622 -24573 5680 -24539
rect 5622 -24607 5634 -24573
rect 5668 -24607 5680 -24573
rect 5622 -24652 5680 -24607
rect 6640 -24097 6698 -24052
rect 6640 -24131 6652 -24097
rect 6686 -24131 6698 -24097
rect 6640 -24165 6698 -24131
rect 6640 -24199 6652 -24165
rect 6686 -24199 6698 -24165
rect 6640 -24233 6698 -24199
rect 6640 -24267 6652 -24233
rect 6686 -24267 6698 -24233
rect 6640 -24301 6698 -24267
rect 6640 -24335 6652 -24301
rect 6686 -24335 6698 -24301
rect 6640 -24369 6698 -24335
rect 6640 -24403 6652 -24369
rect 6686 -24403 6698 -24369
rect 6640 -24437 6698 -24403
rect 6640 -24471 6652 -24437
rect 6686 -24471 6698 -24437
rect 6640 -24505 6698 -24471
rect 6640 -24539 6652 -24505
rect 6686 -24539 6698 -24505
rect 6640 -24573 6698 -24539
rect 6640 -24607 6652 -24573
rect 6686 -24607 6698 -24573
rect 6640 -24652 6698 -24607
rect 7658 -24097 7716 -24052
rect 7658 -24131 7670 -24097
rect 7704 -24131 7716 -24097
rect 7658 -24165 7716 -24131
rect 7658 -24199 7670 -24165
rect 7704 -24199 7716 -24165
rect 7658 -24233 7716 -24199
rect 7658 -24267 7670 -24233
rect 7704 -24267 7716 -24233
rect 7658 -24301 7716 -24267
rect 7658 -24335 7670 -24301
rect 7704 -24335 7716 -24301
rect 7658 -24369 7716 -24335
rect 7658 -24403 7670 -24369
rect 7704 -24403 7716 -24369
rect 7658 -24437 7716 -24403
rect 7658 -24471 7670 -24437
rect 7704 -24471 7716 -24437
rect 7658 -24505 7716 -24471
rect 7658 -24539 7670 -24505
rect 7704 -24539 7716 -24505
rect 7658 -24573 7716 -24539
rect 7658 -24607 7670 -24573
rect 7704 -24607 7716 -24573
rect 7658 -24652 7716 -24607
rect 8676 -24097 8734 -24052
rect 8676 -24131 8688 -24097
rect 8722 -24131 8734 -24097
rect 8676 -24165 8734 -24131
rect 8676 -24199 8688 -24165
rect 8722 -24199 8734 -24165
rect 8676 -24233 8734 -24199
rect 8676 -24267 8688 -24233
rect 8722 -24267 8734 -24233
rect 8676 -24301 8734 -24267
rect 8676 -24335 8688 -24301
rect 8722 -24335 8734 -24301
rect 8676 -24369 8734 -24335
rect 8676 -24403 8688 -24369
rect 8722 -24403 8734 -24369
rect 8676 -24437 8734 -24403
rect 8676 -24471 8688 -24437
rect 8722 -24471 8734 -24437
rect 8676 -24505 8734 -24471
rect 8676 -24539 8688 -24505
rect 8722 -24539 8734 -24505
rect 8676 -24573 8734 -24539
rect 8676 -24607 8688 -24573
rect 8722 -24607 8734 -24573
rect 8676 -24652 8734 -24607
rect 9694 -24097 9752 -24052
rect 9694 -24131 9706 -24097
rect 9740 -24131 9752 -24097
rect 9694 -24165 9752 -24131
rect 9694 -24199 9706 -24165
rect 9740 -24199 9752 -24165
rect 9694 -24233 9752 -24199
rect 9694 -24267 9706 -24233
rect 9740 -24267 9752 -24233
rect 9694 -24301 9752 -24267
rect 9694 -24335 9706 -24301
rect 9740 -24335 9752 -24301
rect 9694 -24369 9752 -24335
rect 9694 -24403 9706 -24369
rect 9740 -24403 9752 -24369
rect 9694 -24437 9752 -24403
rect 9694 -24471 9706 -24437
rect 9740 -24471 9752 -24437
rect 9694 -24505 9752 -24471
rect 9694 -24539 9706 -24505
rect 9740 -24539 9752 -24505
rect 9694 -24573 9752 -24539
rect 9694 -24607 9706 -24573
rect 9740 -24607 9752 -24573
rect 9694 -24652 9752 -24607
rect 10712 -24097 10770 -24052
rect 10712 -24131 10724 -24097
rect 10758 -24131 10770 -24097
rect 10712 -24165 10770 -24131
rect 10712 -24199 10724 -24165
rect 10758 -24199 10770 -24165
rect 10712 -24233 10770 -24199
rect 10712 -24267 10724 -24233
rect 10758 -24267 10770 -24233
rect 10712 -24301 10770 -24267
rect 10712 -24335 10724 -24301
rect 10758 -24335 10770 -24301
rect 10712 -24369 10770 -24335
rect 10712 -24403 10724 -24369
rect 10758 -24403 10770 -24369
rect 10712 -24437 10770 -24403
rect 10712 -24471 10724 -24437
rect 10758 -24471 10770 -24437
rect 10712 -24505 10770 -24471
rect 10712 -24539 10724 -24505
rect 10758 -24539 10770 -24505
rect 10712 -24573 10770 -24539
rect 10712 -24607 10724 -24573
rect 10758 -24607 10770 -24573
rect 10712 -24652 10770 -24607
rect 11730 -24097 11788 -24052
rect 11730 -24131 11742 -24097
rect 11776 -24131 11788 -24097
rect 11730 -24165 11788 -24131
rect 11730 -24199 11742 -24165
rect 11776 -24199 11788 -24165
rect 11730 -24233 11788 -24199
rect 11730 -24267 11742 -24233
rect 11776 -24267 11788 -24233
rect 11730 -24301 11788 -24267
rect 11730 -24335 11742 -24301
rect 11776 -24335 11788 -24301
rect 11730 -24369 11788 -24335
rect 11730 -24403 11742 -24369
rect 11776 -24403 11788 -24369
rect 11730 -24437 11788 -24403
rect 11730 -24471 11742 -24437
rect 11776 -24471 11788 -24437
rect 11730 -24505 11788 -24471
rect 11730 -24539 11742 -24505
rect 11776 -24539 11788 -24505
rect 11730 -24573 11788 -24539
rect 11730 -24607 11742 -24573
rect 11776 -24607 11788 -24573
rect 11730 -24652 11788 -24607
rect 12748 -24097 12806 -24052
rect 12748 -24131 12760 -24097
rect 12794 -24131 12806 -24097
rect 12748 -24165 12806 -24131
rect 12748 -24199 12760 -24165
rect 12794 -24199 12806 -24165
rect 12748 -24233 12806 -24199
rect 12748 -24267 12760 -24233
rect 12794 -24267 12806 -24233
rect 12748 -24301 12806 -24267
rect 12748 -24335 12760 -24301
rect 12794 -24335 12806 -24301
rect 12748 -24369 12806 -24335
rect 12748 -24403 12760 -24369
rect 12794 -24403 12806 -24369
rect 12748 -24437 12806 -24403
rect 12748 -24471 12760 -24437
rect 12794 -24471 12806 -24437
rect 12748 -24505 12806 -24471
rect 12748 -24539 12760 -24505
rect 12794 -24539 12806 -24505
rect 12748 -24573 12806 -24539
rect 12748 -24607 12760 -24573
rect 12794 -24607 12806 -24573
rect 12748 -24652 12806 -24607
rect 13766 -24097 13824 -24052
rect 13766 -24131 13778 -24097
rect 13812 -24131 13824 -24097
rect 13766 -24165 13824 -24131
rect 13766 -24199 13778 -24165
rect 13812 -24199 13824 -24165
rect 13766 -24233 13824 -24199
rect 13766 -24267 13778 -24233
rect 13812 -24267 13824 -24233
rect 13766 -24301 13824 -24267
rect 13766 -24335 13778 -24301
rect 13812 -24335 13824 -24301
rect 13766 -24369 13824 -24335
rect 13766 -24403 13778 -24369
rect 13812 -24403 13824 -24369
rect 13766 -24437 13824 -24403
rect 13766 -24471 13778 -24437
rect 13812 -24471 13824 -24437
rect 13766 -24505 13824 -24471
rect 13766 -24539 13778 -24505
rect 13812 -24539 13824 -24505
rect 13766 -24573 13824 -24539
rect 13766 -24607 13778 -24573
rect 13812 -24607 13824 -24573
rect 13766 -24652 13824 -24607
rect 14784 -24097 14842 -24052
rect 14784 -24131 14796 -24097
rect 14830 -24131 14842 -24097
rect 14784 -24165 14842 -24131
rect 14784 -24199 14796 -24165
rect 14830 -24199 14842 -24165
rect 14784 -24233 14842 -24199
rect 14784 -24267 14796 -24233
rect 14830 -24267 14842 -24233
rect 14784 -24301 14842 -24267
rect 14784 -24335 14796 -24301
rect 14830 -24335 14842 -24301
rect 14784 -24369 14842 -24335
rect 14784 -24403 14796 -24369
rect 14830 -24403 14842 -24369
rect 14784 -24437 14842 -24403
rect 14784 -24471 14796 -24437
rect 14830 -24471 14842 -24437
rect 14784 -24505 14842 -24471
rect 14784 -24539 14796 -24505
rect 14830 -24539 14842 -24505
rect 14784 -24573 14842 -24539
rect 14784 -24607 14796 -24573
rect 14830 -24607 14842 -24573
rect 14784 -24652 14842 -24607
rect 15802 -24097 15860 -24052
rect 15802 -24131 15814 -24097
rect 15848 -24131 15860 -24097
rect 15802 -24165 15860 -24131
rect 15802 -24199 15814 -24165
rect 15848 -24199 15860 -24165
rect 15802 -24233 15860 -24199
rect 15802 -24267 15814 -24233
rect 15848 -24267 15860 -24233
rect 15802 -24301 15860 -24267
rect 15802 -24335 15814 -24301
rect 15848 -24335 15860 -24301
rect 15802 -24369 15860 -24335
rect 15802 -24403 15814 -24369
rect 15848 -24403 15860 -24369
rect 15802 -24437 15860 -24403
rect 15802 -24471 15814 -24437
rect 15848 -24471 15860 -24437
rect 15802 -24505 15860 -24471
rect 15802 -24539 15814 -24505
rect 15848 -24539 15860 -24505
rect 15802 -24573 15860 -24539
rect 15802 -24607 15814 -24573
rect 15848 -24607 15860 -24573
rect 15802 -24652 15860 -24607
rect 16820 -24097 16878 -24052
rect 16820 -24131 16832 -24097
rect 16866 -24131 16878 -24097
rect 16820 -24165 16878 -24131
rect 16820 -24199 16832 -24165
rect 16866 -24199 16878 -24165
rect 16820 -24233 16878 -24199
rect 16820 -24267 16832 -24233
rect 16866 -24267 16878 -24233
rect 16820 -24301 16878 -24267
rect 16820 -24335 16832 -24301
rect 16866 -24335 16878 -24301
rect 16820 -24369 16878 -24335
rect 16820 -24403 16832 -24369
rect 16866 -24403 16878 -24369
rect 16820 -24437 16878 -24403
rect 16820 -24471 16832 -24437
rect 16866 -24471 16878 -24437
rect 16820 -24505 16878 -24471
rect 16820 -24539 16832 -24505
rect 16866 -24539 16878 -24505
rect 16820 -24573 16878 -24539
rect 16820 -24607 16832 -24573
rect 16866 -24607 16878 -24573
rect 16820 -24652 16878 -24607
rect 17838 -24097 17896 -24052
rect 17838 -24131 17850 -24097
rect 17884 -24131 17896 -24097
rect 17838 -24165 17896 -24131
rect 17838 -24199 17850 -24165
rect 17884 -24199 17896 -24165
rect 17838 -24233 17896 -24199
rect 17838 -24267 17850 -24233
rect 17884 -24267 17896 -24233
rect 17838 -24301 17896 -24267
rect 17838 -24335 17850 -24301
rect 17884 -24335 17896 -24301
rect 17838 -24369 17896 -24335
rect 17838 -24403 17850 -24369
rect 17884 -24403 17896 -24369
rect 17838 -24437 17896 -24403
rect 17838 -24471 17850 -24437
rect 17884 -24471 17896 -24437
rect 17838 -24505 17896 -24471
rect 17838 -24539 17850 -24505
rect 17884 -24539 17896 -24505
rect 17838 -24573 17896 -24539
rect 17838 -24607 17850 -24573
rect 17884 -24607 17896 -24573
rect 17838 -24652 17896 -24607
rect 18856 -24097 18914 -24052
rect 18856 -24131 18868 -24097
rect 18902 -24131 18914 -24097
rect 18856 -24165 18914 -24131
rect 18856 -24199 18868 -24165
rect 18902 -24199 18914 -24165
rect 18856 -24233 18914 -24199
rect 18856 -24267 18868 -24233
rect 18902 -24267 18914 -24233
rect 18856 -24301 18914 -24267
rect 18856 -24335 18868 -24301
rect 18902 -24335 18914 -24301
rect 18856 -24369 18914 -24335
rect 18856 -24403 18868 -24369
rect 18902 -24403 18914 -24369
rect 18856 -24437 18914 -24403
rect 18856 -24471 18868 -24437
rect 18902 -24471 18914 -24437
rect 18856 -24505 18914 -24471
rect 18856 -24539 18868 -24505
rect 18902 -24539 18914 -24505
rect 18856 -24573 18914 -24539
rect 18856 -24607 18868 -24573
rect 18902 -24607 18914 -24573
rect 18856 -24652 18914 -24607
rect 19874 -24097 19932 -24052
rect 19874 -24131 19886 -24097
rect 19920 -24131 19932 -24097
rect 19874 -24165 19932 -24131
rect 19874 -24199 19886 -24165
rect 19920 -24199 19932 -24165
rect 19874 -24233 19932 -24199
rect 19874 -24267 19886 -24233
rect 19920 -24267 19932 -24233
rect 19874 -24301 19932 -24267
rect 19874 -24335 19886 -24301
rect 19920 -24335 19932 -24301
rect 19874 -24369 19932 -24335
rect 19874 -24403 19886 -24369
rect 19920 -24403 19932 -24369
rect 19874 -24437 19932 -24403
rect 19874 -24471 19886 -24437
rect 19920 -24471 19932 -24437
rect 19874 -24505 19932 -24471
rect 19874 -24539 19886 -24505
rect 19920 -24539 19932 -24505
rect 19874 -24573 19932 -24539
rect 19874 -24607 19886 -24573
rect 19920 -24607 19932 -24573
rect 19874 -24652 19932 -24607
rect 20892 -24097 20950 -24052
rect 20892 -24131 20904 -24097
rect 20938 -24131 20950 -24097
rect 20892 -24165 20950 -24131
rect 20892 -24199 20904 -24165
rect 20938 -24199 20950 -24165
rect 20892 -24233 20950 -24199
rect 20892 -24267 20904 -24233
rect 20938 -24267 20950 -24233
rect 20892 -24301 20950 -24267
rect 20892 -24335 20904 -24301
rect 20938 -24335 20950 -24301
rect 20892 -24369 20950 -24335
rect 20892 -24403 20904 -24369
rect 20938 -24403 20950 -24369
rect 20892 -24437 20950 -24403
rect 20892 -24471 20904 -24437
rect 20938 -24471 20950 -24437
rect 20892 -24505 20950 -24471
rect 20892 -24539 20904 -24505
rect 20938 -24539 20950 -24505
rect 20892 -24573 20950 -24539
rect 20892 -24607 20904 -24573
rect 20938 -24607 20950 -24573
rect 20892 -24652 20950 -24607
rect 21910 -24097 21968 -24052
rect 21910 -24131 21922 -24097
rect 21956 -24131 21968 -24097
rect 21910 -24165 21968 -24131
rect 21910 -24199 21922 -24165
rect 21956 -24199 21968 -24165
rect 21910 -24233 21968 -24199
rect 21910 -24267 21922 -24233
rect 21956 -24267 21968 -24233
rect 21910 -24301 21968 -24267
rect 21910 -24335 21922 -24301
rect 21956 -24335 21968 -24301
rect 21910 -24369 21968 -24335
rect 21910 -24403 21922 -24369
rect 21956 -24403 21968 -24369
rect 21910 -24437 21968 -24403
rect 21910 -24471 21922 -24437
rect 21956 -24471 21968 -24437
rect 21910 -24505 21968 -24471
rect 21910 -24539 21922 -24505
rect 21956 -24539 21968 -24505
rect 21910 -24573 21968 -24539
rect 21910 -24607 21922 -24573
rect 21956 -24607 21968 -24573
rect 21910 -24652 21968 -24607
rect 22928 -24097 22986 -24052
rect 22928 -24131 22940 -24097
rect 22974 -24131 22986 -24097
rect 22928 -24165 22986 -24131
rect 22928 -24199 22940 -24165
rect 22974 -24199 22986 -24165
rect 22928 -24233 22986 -24199
rect 22928 -24267 22940 -24233
rect 22974 -24267 22986 -24233
rect 22928 -24301 22986 -24267
rect 22928 -24335 22940 -24301
rect 22974 -24335 22986 -24301
rect 22928 -24369 22986 -24335
rect 22928 -24403 22940 -24369
rect 22974 -24403 22986 -24369
rect 22928 -24437 22986 -24403
rect 22928 -24471 22940 -24437
rect 22974 -24471 22986 -24437
rect 22928 -24505 22986 -24471
rect 22928 -24539 22940 -24505
rect 22974 -24539 22986 -24505
rect 22928 -24573 22986 -24539
rect 22928 -24607 22940 -24573
rect 22974 -24607 22986 -24573
rect 22928 -24652 22986 -24607
rect -9418 -25163 -9360 -25118
rect -9418 -25197 -9406 -25163
rect -9372 -25197 -9360 -25163
rect -9418 -25231 -9360 -25197
rect -9418 -25265 -9406 -25231
rect -9372 -25265 -9360 -25231
rect -9418 -25299 -9360 -25265
rect -9418 -25333 -9406 -25299
rect -9372 -25333 -9360 -25299
rect -9418 -25367 -9360 -25333
rect -9418 -25401 -9406 -25367
rect -9372 -25401 -9360 -25367
rect -9418 -25435 -9360 -25401
rect -9418 -25469 -9406 -25435
rect -9372 -25469 -9360 -25435
rect -9418 -25503 -9360 -25469
rect -9418 -25537 -9406 -25503
rect -9372 -25537 -9360 -25503
rect -9418 -25571 -9360 -25537
rect -9418 -25605 -9406 -25571
rect -9372 -25605 -9360 -25571
rect -9418 -25639 -9360 -25605
rect -9418 -25673 -9406 -25639
rect -9372 -25673 -9360 -25639
rect -9418 -25718 -9360 -25673
rect -8400 -25163 -8342 -25118
rect -8400 -25197 -8388 -25163
rect -8354 -25197 -8342 -25163
rect -8400 -25231 -8342 -25197
rect -8400 -25265 -8388 -25231
rect -8354 -25265 -8342 -25231
rect -8400 -25299 -8342 -25265
rect -8400 -25333 -8388 -25299
rect -8354 -25333 -8342 -25299
rect -8400 -25367 -8342 -25333
rect -8400 -25401 -8388 -25367
rect -8354 -25401 -8342 -25367
rect -8400 -25435 -8342 -25401
rect -8400 -25469 -8388 -25435
rect -8354 -25469 -8342 -25435
rect -8400 -25503 -8342 -25469
rect -8400 -25537 -8388 -25503
rect -8354 -25537 -8342 -25503
rect -8400 -25571 -8342 -25537
rect -8400 -25605 -8388 -25571
rect -8354 -25605 -8342 -25571
rect -8400 -25639 -8342 -25605
rect -8400 -25673 -8388 -25639
rect -8354 -25673 -8342 -25639
rect -8400 -25718 -8342 -25673
rect -7382 -25163 -7324 -25118
rect -7382 -25197 -7370 -25163
rect -7336 -25197 -7324 -25163
rect -7382 -25231 -7324 -25197
rect -7382 -25265 -7370 -25231
rect -7336 -25265 -7324 -25231
rect -7382 -25299 -7324 -25265
rect -7382 -25333 -7370 -25299
rect -7336 -25333 -7324 -25299
rect -7382 -25367 -7324 -25333
rect -7382 -25401 -7370 -25367
rect -7336 -25401 -7324 -25367
rect -7382 -25435 -7324 -25401
rect -7382 -25469 -7370 -25435
rect -7336 -25469 -7324 -25435
rect -7382 -25503 -7324 -25469
rect -7382 -25537 -7370 -25503
rect -7336 -25537 -7324 -25503
rect -7382 -25571 -7324 -25537
rect -7382 -25605 -7370 -25571
rect -7336 -25605 -7324 -25571
rect -7382 -25639 -7324 -25605
rect -7382 -25673 -7370 -25639
rect -7336 -25673 -7324 -25639
rect -7382 -25718 -7324 -25673
rect -6364 -25163 -6306 -25118
rect -6364 -25197 -6352 -25163
rect -6318 -25197 -6306 -25163
rect -6364 -25231 -6306 -25197
rect -6364 -25265 -6352 -25231
rect -6318 -25265 -6306 -25231
rect -6364 -25299 -6306 -25265
rect -6364 -25333 -6352 -25299
rect -6318 -25333 -6306 -25299
rect -6364 -25367 -6306 -25333
rect -6364 -25401 -6352 -25367
rect -6318 -25401 -6306 -25367
rect -6364 -25435 -6306 -25401
rect -6364 -25469 -6352 -25435
rect -6318 -25469 -6306 -25435
rect -6364 -25503 -6306 -25469
rect -6364 -25537 -6352 -25503
rect -6318 -25537 -6306 -25503
rect -6364 -25571 -6306 -25537
rect -6364 -25605 -6352 -25571
rect -6318 -25605 -6306 -25571
rect -6364 -25639 -6306 -25605
rect -6364 -25673 -6352 -25639
rect -6318 -25673 -6306 -25639
rect -6364 -25718 -6306 -25673
rect -5346 -25163 -5288 -25118
rect -5346 -25197 -5334 -25163
rect -5300 -25197 -5288 -25163
rect -5346 -25231 -5288 -25197
rect -5346 -25265 -5334 -25231
rect -5300 -25265 -5288 -25231
rect -5346 -25299 -5288 -25265
rect -5346 -25333 -5334 -25299
rect -5300 -25333 -5288 -25299
rect -5346 -25367 -5288 -25333
rect -5346 -25401 -5334 -25367
rect -5300 -25401 -5288 -25367
rect -5346 -25435 -5288 -25401
rect -5346 -25469 -5334 -25435
rect -5300 -25469 -5288 -25435
rect -5346 -25503 -5288 -25469
rect -5346 -25537 -5334 -25503
rect -5300 -25537 -5288 -25503
rect -5346 -25571 -5288 -25537
rect -5346 -25605 -5334 -25571
rect -5300 -25605 -5288 -25571
rect -5346 -25639 -5288 -25605
rect -5346 -25673 -5334 -25639
rect -5300 -25673 -5288 -25639
rect -5346 -25718 -5288 -25673
rect -4328 -25163 -4270 -25118
rect -4328 -25197 -4316 -25163
rect -4282 -25197 -4270 -25163
rect -4328 -25231 -4270 -25197
rect -4328 -25265 -4316 -25231
rect -4282 -25265 -4270 -25231
rect -4328 -25299 -4270 -25265
rect -4328 -25333 -4316 -25299
rect -4282 -25333 -4270 -25299
rect -4328 -25367 -4270 -25333
rect -4328 -25401 -4316 -25367
rect -4282 -25401 -4270 -25367
rect -4328 -25435 -4270 -25401
rect -4328 -25469 -4316 -25435
rect -4282 -25469 -4270 -25435
rect -4328 -25503 -4270 -25469
rect -4328 -25537 -4316 -25503
rect -4282 -25537 -4270 -25503
rect -4328 -25571 -4270 -25537
rect -4328 -25605 -4316 -25571
rect -4282 -25605 -4270 -25571
rect -4328 -25639 -4270 -25605
rect -4328 -25673 -4316 -25639
rect -4282 -25673 -4270 -25639
rect -4328 -25718 -4270 -25673
rect -3310 -25163 -3252 -25118
rect -3310 -25197 -3298 -25163
rect -3264 -25197 -3252 -25163
rect -3310 -25231 -3252 -25197
rect -3310 -25265 -3298 -25231
rect -3264 -25265 -3252 -25231
rect -3310 -25299 -3252 -25265
rect -3310 -25333 -3298 -25299
rect -3264 -25333 -3252 -25299
rect -3310 -25367 -3252 -25333
rect -3310 -25401 -3298 -25367
rect -3264 -25401 -3252 -25367
rect -3310 -25435 -3252 -25401
rect -3310 -25469 -3298 -25435
rect -3264 -25469 -3252 -25435
rect -3310 -25503 -3252 -25469
rect -3310 -25537 -3298 -25503
rect -3264 -25537 -3252 -25503
rect -3310 -25571 -3252 -25537
rect -3310 -25605 -3298 -25571
rect -3264 -25605 -3252 -25571
rect -3310 -25639 -3252 -25605
rect -3310 -25673 -3298 -25639
rect -3264 -25673 -3252 -25639
rect -3310 -25718 -3252 -25673
rect -2424 -25159 -2366 -25114
rect -2424 -25193 -2412 -25159
rect -2378 -25193 -2366 -25159
rect -2424 -25227 -2366 -25193
rect -2424 -25261 -2412 -25227
rect -2378 -25261 -2366 -25227
rect -2424 -25295 -2366 -25261
rect -2424 -25329 -2412 -25295
rect -2378 -25329 -2366 -25295
rect -2424 -25363 -2366 -25329
rect -2424 -25397 -2412 -25363
rect -2378 -25397 -2366 -25363
rect -2424 -25431 -2366 -25397
rect -2424 -25465 -2412 -25431
rect -2378 -25465 -2366 -25431
rect -2424 -25499 -2366 -25465
rect -2424 -25533 -2412 -25499
rect -2378 -25533 -2366 -25499
rect -2424 -25567 -2366 -25533
rect -2424 -25601 -2412 -25567
rect -2378 -25601 -2366 -25567
rect -2424 -25635 -2366 -25601
rect -2424 -25669 -2412 -25635
rect -2378 -25669 -2366 -25635
rect -2424 -25714 -2366 -25669
rect -2126 -25159 -2068 -25114
rect -2126 -25193 -2114 -25159
rect -2080 -25193 -2068 -25159
rect -2126 -25227 -2068 -25193
rect -2126 -25261 -2114 -25227
rect -2080 -25261 -2068 -25227
rect -2126 -25295 -2068 -25261
rect -2126 -25329 -2114 -25295
rect -2080 -25329 -2068 -25295
rect -2126 -25363 -2068 -25329
rect -2126 -25397 -2114 -25363
rect -2080 -25397 -2068 -25363
rect -2126 -25431 -2068 -25397
rect -2126 -25465 -2114 -25431
rect -2080 -25465 -2068 -25431
rect -2126 -25499 -2068 -25465
rect -2126 -25533 -2114 -25499
rect -2080 -25533 -2068 -25499
rect -2126 -25567 -2068 -25533
rect -2126 -25601 -2114 -25567
rect -2080 -25601 -2068 -25567
rect -2126 -25635 -2068 -25601
rect -2126 -25669 -2114 -25635
rect -2080 -25669 -2068 -25635
rect -2126 -25714 -2068 -25669
rect -1828 -25159 -1770 -25114
rect -1828 -25193 -1816 -25159
rect -1782 -25193 -1770 -25159
rect -1828 -25227 -1770 -25193
rect -1828 -25261 -1816 -25227
rect -1782 -25261 -1770 -25227
rect -1828 -25295 -1770 -25261
rect -1828 -25329 -1816 -25295
rect -1782 -25329 -1770 -25295
rect -1828 -25363 -1770 -25329
rect -1828 -25397 -1816 -25363
rect -1782 -25397 -1770 -25363
rect -1828 -25431 -1770 -25397
rect -1828 -25465 -1816 -25431
rect -1782 -25465 -1770 -25431
rect -1828 -25499 -1770 -25465
rect -1828 -25533 -1816 -25499
rect -1782 -25533 -1770 -25499
rect -1828 -25567 -1770 -25533
rect -1828 -25601 -1816 -25567
rect -1782 -25601 -1770 -25567
rect -1828 -25635 -1770 -25601
rect -1828 -25669 -1816 -25635
rect -1782 -25669 -1770 -25635
rect -1828 -25714 -1770 -25669
rect -1530 -25159 -1472 -25114
rect -1530 -25193 -1518 -25159
rect -1484 -25193 -1472 -25159
rect -1530 -25227 -1472 -25193
rect -1530 -25261 -1518 -25227
rect -1484 -25261 -1472 -25227
rect -1530 -25295 -1472 -25261
rect -1530 -25329 -1518 -25295
rect -1484 -25329 -1472 -25295
rect -1530 -25363 -1472 -25329
rect -1530 -25397 -1518 -25363
rect -1484 -25397 -1472 -25363
rect -1530 -25431 -1472 -25397
rect -1530 -25465 -1518 -25431
rect -1484 -25465 -1472 -25431
rect -1530 -25499 -1472 -25465
rect -1530 -25533 -1518 -25499
rect -1484 -25533 -1472 -25499
rect -1530 -25567 -1472 -25533
rect -1530 -25601 -1518 -25567
rect -1484 -25601 -1472 -25567
rect -1530 -25635 -1472 -25601
rect -1530 -25669 -1518 -25635
rect -1484 -25669 -1472 -25635
rect -1530 -25714 -1472 -25669
rect -1232 -25159 -1174 -25114
rect -1232 -25193 -1220 -25159
rect -1186 -25193 -1174 -25159
rect -1232 -25227 -1174 -25193
rect -1232 -25261 -1220 -25227
rect -1186 -25261 -1174 -25227
rect -1232 -25295 -1174 -25261
rect -1232 -25329 -1220 -25295
rect -1186 -25329 -1174 -25295
rect -1232 -25363 -1174 -25329
rect -1232 -25397 -1220 -25363
rect -1186 -25397 -1174 -25363
rect -1232 -25431 -1174 -25397
rect -1232 -25465 -1220 -25431
rect -1186 -25465 -1174 -25431
rect -1232 -25499 -1174 -25465
rect -1232 -25533 -1220 -25499
rect -1186 -25533 -1174 -25499
rect -1232 -25567 -1174 -25533
rect -1232 -25601 -1220 -25567
rect -1186 -25601 -1174 -25567
rect -1232 -25635 -1174 -25601
rect -1232 -25669 -1220 -25635
rect -1186 -25669 -1174 -25635
rect -1232 -25714 -1174 -25669
rect -934 -25159 -876 -25114
rect -934 -25193 -922 -25159
rect -888 -25193 -876 -25159
rect -934 -25227 -876 -25193
rect -934 -25261 -922 -25227
rect -888 -25261 -876 -25227
rect -934 -25295 -876 -25261
rect -934 -25329 -922 -25295
rect -888 -25329 -876 -25295
rect -934 -25363 -876 -25329
rect -934 -25397 -922 -25363
rect -888 -25397 -876 -25363
rect -934 -25431 -876 -25397
rect -934 -25465 -922 -25431
rect -888 -25465 -876 -25431
rect -934 -25499 -876 -25465
rect -934 -25533 -922 -25499
rect -888 -25533 -876 -25499
rect -934 -25567 -876 -25533
rect -934 -25601 -922 -25567
rect -888 -25601 -876 -25567
rect -934 -25635 -876 -25601
rect -934 -25669 -922 -25635
rect -888 -25669 -876 -25635
rect -934 -25714 -876 -25669
rect -636 -25159 -578 -25114
rect -636 -25193 -624 -25159
rect -590 -25193 -578 -25159
rect -636 -25227 -578 -25193
rect -636 -25261 -624 -25227
rect -590 -25261 -578 -25227
rect -636 -25295 -578 -25261
rect -636 -25329 -624 -25295
rect -590 -25329 -578 -25295
rect -636 -25363 -578 -25329
rect -636 -25397 -624 -25363
rect -590 -25397 -578 -25363
rect -636 -25431 -578 -25397
rect -636 -25465 -624 -25431
rect -590 -25465 -578 -25431
rect -636 -25499 -578 -25465
rect -636 -25533 -624 -25499
rect -590 -25533 -578 -25499
rect -636 -25567 -578 -25533
rect -636 -25601 -624 -25567
rect -590 -25601 -578 -25567
rect -636 -25635 -578 -25601
rect -636 -25669 -624 -25635
rect -590 -25669 -578 -25635
rect -636 -25714 -578 -25669
rect -338 -25159 -280 -25114
rect -338 -25193 -326 -25159
rect -292 -25193 -280 -25159
rect -338 -25227 -280 -25193
rect -338 -25261 -326 -25227
rect -292 -25261 -280 -25227
rect -338 -25295 -280 -25261
rect -338 -25329 -326 -25295
rect -292 -25329 -280 -25295
rect -338 -25363 -280 -25329
rect -338 -25397 -326 -25363
rect -292 -25397 -280 -25363
rect -338 -25431 -280 -25397
rect -338 -25465 -326 -25431
rect -292 -25465 -280 -25431
rect -338 -25499 -280 -25465
rect -338 -25533 -326 -25499
rect -292 -25533 -280 -25499
rect -338 -25567 -280 -25533
rect -338 -25601 -326 -25567
rect -292 -25601 -280 -25567
rect -338 -25635 -280 -25601
rect -338 -25669 -326 -25635
rect -292 -25669 -280 -25635
rect -338 -25714 -280 -25669
rect -40 -25159 18 -25114
rect -40 -25193 -28 -25159
rect 6 -25193 18 -25159
rect -40 -25227 18 -25193
rect -40 -25261 -28 -25227
rect 6 -25261 18 -25227
rect -40 -25295 18 -25261
rect -40 -25329 -28 -25295
rect 6 -25329 18 -25295
rect -40 -25363 18 -25329
rect -40 -25397 -28 -25363
rect 6 -25397 18 -25363
rect -40 -25431 18 -25397
rect -40 -25465 -28 -25431
rect 6 -25465 18 -25431
rect -40 -25499 18 -25465
rect -40 -25533 -28 -25499
rect 6 -25533 18 -25499
rect -40 -25567 18 -25533
rect -40 -25601 -28 -25567
rect 6 -25601 18 -25567
rect -40 -25635 18 -25601
rect -40 -25669 -28 -25635
rect 6 -25669 18 -25635
rect -40 -25714 18 -25669
rect 258 -25159 316 -25114
rect 258 -25193 270 -25159
rect 304 -25193 316 -25159
rect 258 -25227 316 -25193
rect 258 -25261 270 -25227
rect 304 -25261 316 -25227
rect 258 -25295 316 -25261
rect 258 -25329 270 -25295
rect 304 -25329 316 -25295
rect 258 -25363 316 -25329
rect 258 -25397 270 -25363
rect 304 -25397 316 -25363
rect 258 -25431 316 -25397
rect 258 -25465 270 -25431
rect 304 -25465 316 -25431
rect 258 -25499 316 -25465
rect 258 -25533 270 -25499
rect 304 -25533 316 -25499
rect 258 -25567 316 -25533
rect 258 -25601 270 -25567
rect 304 -25601 316 -25567
rect 258 -25635 316 -25601
rect 258 -25669 270 -25635
rect 304 -25669 316 -25635
rect 258 -25714 316 -25669
rect 556 -25159 614 -25114
rect 556 -25193 568 -25159
rect 602 -25193 614 -25159
rect 556 -25227 614 -25193
rect 556 -25261 568 -25227
rect 602 -25261 614 -25227
rect 556 -25295 614 -25261
rect 556 -25329 568 -25295
rect 602 -25329 614 -25295
rect 556 -25363 614 -25329
rect 556 -25397 568 -25363
rect 602 -25397 614 -25363
rect 556 -25431 614 -25397
rect 556 -25465 568 -25431
rect 602 -25465 614 -25431
rect 556 -25499 614 -25465
rect 556 -25533 568 -25499
rect 602 -25533 614 -25499
rect 556 -25567 614 -25533
rect 556 -25601 568 -25567
rect 602 -25601 614 -25567
rect 556 -25635 614 -25601
rect 556 -25669 568 -25635
rect 602 -25669 614 -25635
rect 556 -25714 614 -25669
rect 854 -25159 912 -25114
rect 854 -25193 866 -25159
rect 900 -25193 912 -25159
rect 854 -25227 912 -25193
rect 854 -25261 866 -25227
rect 900 -25261 912 -25227
rect 854 -25295 912 -25261
rect 854 -25329 866 -25295
rect 900 -25329 912 -25295
rect 854 -25363 912 -25329
rect 854 -25397 866 -25363
rect 900 -25397 912 -25363
rect 854 -25431 912 -25397
rect 854 -25465 866 -25431
rect 900 -25465 912 -25431
rect 854 -25499 912 -25465
rect 854 -25533 866 -25499
rect 900 -25533 912 -25499
rect 854 -25567 912 -25533
rect 854 -25601 866 -25567
rect 900 -25601 912 -25567
rect 854 -25635 912 -25601
rect 854 -25669 866 -25635
rect 900 -25669 912 -25635
rect 854 -25714 912 -25669
rect 2568 -25329 2626 -25284
rect 2568 -25363 2580 -25329
rect 2614 -25363 2626 -25329
rect 2568 -25397 2626 -25363
rect 2568 -25431 2580 -25397
rect 2614 -25431 2626 -25397
rect 2568 -25465 2626 -25431
rect 2568 -25499 2580 -25465
rect 2614 -25499 2626 -25465
rect 2568 -25533 2626 -25499
rect 2568 -25567 2580 -25533
rect 2614 -25567 2626 -25533
rect 2568 -25601 2626 -25567
rect 2568 -25635 2580 -25601
rect 2614 -25635 2626 -25601
rect 2568 -25669 2626 -25635
rect 2568 -25703 2580 -25669
rect 2614 -25703 2626 -25669
rect 2568 -25737 2626 -25703
rect 2568 -25771 2580 -25737
rect 2614 -25771 2626 -25737
rect 2568 -25805 2626 -25771
rect 2568 -25839 2580 -25805
rect 2614 -25839 2626 -25805
rect 2568 -25884 2626 -25839
rect 3586 -25329 3644 -25284
rect 3586 -25363 3598 -25329
rect 3632 -25363 3644 -25329
rect 3586 -25397 3644 -25363
rect 3586 -25431 3598 -25397
rect 3632 -25431 3644 -25397
rect 3586 -25465 3644 -25431
rect 3586 -25499 3598 -25465
rect 3632 -25499 3644 -25465
rect 3586 -25533 3644 -25499
rect 3586 -25567 3598 -25533
rect 3632 -25567 3644 -25533
rect 3586 -25601 3644 -25567
rect 3586 -25635 3598 -25601
rect 3632 -25635 3644 -25601
rect 3586 -25669 3644 -25635
rect 3586 -25703 3598 -25669
rect 3632 -25703 3644 -25669
rect 3586 -25737 3644 -25703
rect 3586 -25771 3598 -25737
rect 3632 -25771 3644 -25737
rect 3586 -25805 3644 -25771
rect 3586 -25839 3598 -25805
rect 3632 -25839 3644 -25805
rect 3586 -25884 3644 -25839
rect 4604 -25329 4662 -25284
rect 4604 -25363 4616 -25329
rect 4650 -25363 4662 -25329
rect 4604 -25397 4662 -25363
rect 4604 -25431 4616 -25397
rect 4650 -25431 4662 -25397
rect 4604 -25465 4662 -25431
rect 4604 -25499 4616 -25465
rect 4650 -25499 4662 -25465
rect 4604 -25533 4662 -25499
rect 4604 -25567 4616 -25533
rect 4650 -25567 4662 -25533
rect 4604 -25601 4662 -25567
rect 4604 -25635 4616 -25601
rect 4650 -25635 4662 -25601
rect 4604 -25669 4662 -25635
rect 4604 -25703 4616 -25669
rect 4650 -25703 4662 -25669
rect 4604 -25737 4662 -25703
rect 4604 -25771 4616 -25737
rect 4650 -25771 4662 -25737
rect 4604 -25805 4662 -25771
rect 4604 -25839 4616 -25805
rect 4650 -25839 4662 -25805
rect 4604 -25884 4662 -25839
rect 5622 -25329 5680 -25284
rect 5622 -25363 5634 -25329
rect 5668 -25363 5680 -25329
rect 5622 -25397 5680 -25363
rect 5622 -25431 5634 -25397
rect 5668 -25431 5680 -25397
rect 5622 -25465 5680 -25431
rect 5622 -25499 5634 -25465
rect 5668 -25499 5680 -25465
rect 5622 -25533 5680 -25499
rect 5622 -25567 5634 -25533
rect 5668 -25567 5680 -25533
rect 5622 -25601 5680 -25567
rect 5622 -25635 5634 -25601
rect 5668 -25635 5680 -25601
rect 5622 -25669 5680 -25635
rect 5622 -25703 5634 -25669
rect 5668 -25703 5680 -25669
rect 5622 -25737 5680 -25703
rect 5622 -25771 5634 -25737
rect 5668 -25771 5680 -25737
rect 5622 -25805 5680 -25771
rect 5622 -25839 5634 -25805
rect 5668 -25839 5680 -25805
rect 5622 -25884 5680 -25839
rect 6640 -25329 6698 -25284
rect 6640 -25363 6652 -25329
rect 6686 -25363 6698 -25329
rect 6640 -25397 6698 -25363
rect 6640 -25431 6652 -25397
rect 6686 -25431 6698 -25397
rect 6640 -25465 6698 -25431
rect 6640 -25499 6652 -25465
rect 6686 -25499 6698 -25465
rect 6640 -25533 6698 -25499
rect 6640 -25567 6652 -25533
rect 6686 -25567 6698 -25533
rect 6640 -25601 6698 -25567
rect 6640 -25635 6652 -25601
rect 6686 -25635 6698 -25601
rect 6640 -25669 6698 -25635
rect 6640 -25703 6652 -25669
rect 6686 -25703 6698 -25669
rect 6640 -25737 6698 -25703
rect 6640 -25771 6652 -25737
rect 6686 -25771 6698 -25737
rect 6640 -25805 6698 -25771
rect 6640 -25839 6652 -25805
rect 6686 -25839 6698 -25805
rect 6640 -25884 6698 -25839
rect 7658 -25329 7716 -25284
rect 7658 -25363 7670 -25329
rect 7704 -25363 7716 -25329
rect 7658 -25397 7716 -25363
rect 7658 -25431 7670 -25397
rect 7704 -25431 7716 -25397
rect 7658 -25465 7716 -25431
rect 7658 -25499 7670 -25465
rect 7704 -25499 7716 -25465
rect 7658 -25533 7716 -25499
rect 7658 -25567 7670 -25533
rect 7704 -25567 7716 -25533
rect 7658 -25601 7716 -25567
rect 7658 -25635 7670 -25601
rect 7704 -25635 7716 -25601
rect 7658 -25669 7716 -25635
rect 7658 -25703 7670 -25669
rect 7704 -25703 7716 -25669
rect 7658 -25737 7716 -25703
rect 7658 -25771 7670 -25737
rect 7704 -25771 7716 -25737
rect 7658 -25805 7716 -25771
rect 7658 -25839 7670 -25805
rect 7704 -25839 7716 -25805
rect 7658 -25884 7716 -25839
rect 8676 -25329 8734 -25284
rect 8676 -25363 8688 -25329
rect 8722 -25363 8734 -25329
rect 8676 -25397 8734 -25363
rect 8676 -25431 8688 -25397
rect 8722 -25431 8734 -25397
rect 8676 -25465 8734 -25431
rect 8676 -25499 8688 -25465
rect 8722 -25499 8734 -25465
rect 8676 -25533 8734 -25499
rect 8676 -25567 8688 -25533
rect 8722 -25567 8734 -25533
rect 8676 -25601 8734 -25567
rect 8676 -25635 8688 -25601
rect 8722 -25635 8734 -25601
rect 8676 -25669 8734 -25635
rect 8676 -25703 8688 -25669
rect 8722 -25703 8734 -25669
rect 8676 -25737 8734 -25703
rect 8676 -25771 8688 -25737
rect 8722 -25771 8734 -25737
rect 8676 -25805 8734 -25771
rect 8676 -25839 8688 -25805
rect 8722 -25839 8734 -25805
rect 8676 -25884 8734 -25839
rect 9694 -25329 9752 -25284
rect 9694 -25363 9706 -25329
rect 9740 -25363 9752 -25329
rect 9694 -25397 9752 -25363
rect 9694 -25431 9706 -25397
rect 9740 -25431 9752 -25397
rect 9694 -25465 9752 -25431
rect 9694 -25499 9706 -25465
rect 9740 -25499 9752 -25465
rect 9694 -25533 9752 -25499
rect 9694 -25567 9706 -25533
rect 9740 -25567 9752 -25533
rect 9694 -25601 9752 -25567
rect 9694 -25635 9706 -25601
rect 9740 -25635 9752 -25601
rect 9694 -25669 9752 -25635
rect 9694 -25703 9706 -25669
rect 9740 -25703 9752 -25669
rect 9694 -25737 9752 -25703
rect 9694 -25771 9706 -25737
rect 9740 -25771 9752 -25737
rect 9694 -25805 9752 -25771
rect 9694 -25839 9706 -25805
rect 9740 -25839 9752 -25805
rect 9694 -25884 9752 -25839
rect 10712 -25329 10770 -25284
rect 10712 -25363 10724 -25329
rect 10758 -25363 10770 -25329
rect 10712 -25397 10770 -25363
rect 10712 -25431 10724 -25397
rect 10758 -25431 10770 -25397
rect 10712 -25465 10770 -25431
rect 10712 -25499 10724 -25465
rect 10758 -25499 10770 -25465
rect 10712 -25533 10770 -25499
rect 10712 -25567 10724 -25533
rect 10758 -25567 10770 -25533
rect 10712 -25601 10770 -25567
rect 10712 -25635 10724 -25601
rect 10758 -25635 10770 -25601
rect 10712 -25669 10770 -25635
rect 10712 -25703 10724 -25669
rect 10758 -25703 10770 -25669
rect 10712 -25737 10770 -25703
rect 10712 -25771 10724 -25737
rect 10758 -25771 10770 -25737
rect 10712 -25805 10770 -25771
rect 10712 -25839 10724 -25805
rect 10758 -25839 10770 -25805
rect 10712 -25884 10770 -25839
rect 11730 -25329 11788 -25284
rect 11730 -25363 11742 -25329
rect 11776 -25363 11788 -25329
rect 11730 -25397 11788 -25363
rect 11730 -25431 11742 -25397
rect 11776 -25431 11788 -25397
rect 11730 -25465 11788 -25431
rect 11730 -25499 11742 -25465
rect 11776 -25499 11788 -25465
rect 11730 -25533 11788 -25499
rect 11730 -25567 11742 -25533
rect 11776 -25567 11788 -25533
rect 11730 -25601 11788 -25567
rect 11730 -25635 11742 -25601
rect 11776 -25635 11788 -25601
rect 11730 -25669 11788 -25635
rect 11730 -25703 11742 -25669
rect 11776 -25703 11788 -25669
rect 11730 -25737 11788 -25703
rect 11730 -25771 11742 -25737
rect 11776 -25771 11788 -25737
rect 11730 -25805 11788 -25771
rect 11730 -25839 11742 -25805
rect 11776 -25839 11788 -25805
rect 11730 -25884 11788 -25839
rect 12748 -25329 12806 -25284
rect 12748 -25363 12760 -25329
rect 12794 -25363 12806 -25329
rect 12748 -25397 12806 -25363
rect 12748 -25431 12760 -25397
rect 12794 -25431 12806 -25397
rect 12748 -25465 12806 -25431
rect 12748 -25499 12760 -25465
rect 12794 -25499 12806 -25465
rect 12748 -25533 12806 -25499
rect 12748 -25567 12760 -25533
rect 12794 -25567 12806 -25533
rect 12748 -25601 12806 -25567
rect 12748 -25635 12760 -25601
rect 12794 -25635 12806 -25601
rect 12748 -25669 12806 -25635
rect 12748 -25703 12760 -25669
rect 12794 -25703 12806 -25669
rect 12748 -25737 12806 -25703
rect 12748 -25771 12760 -25737
rect 12794 -25771 12806 -25737
rect 12748 -25805 12806 -25771
rect 12748 -25839 12760 -25805
rect 12794 -25839 12806 -25805
rect 12748 -25884 12806 -25839
rect 13766 -25329 13824 -25284
rect 13766 -25363 13778 -25329
rect 13812 -25363 13824 -25329
rect 13766 -25397 13824 -25363
rect 13766 -25431 13778 -25397
rect 13812 -25431 13824 -25397
rect 13766 -25465 13824 -25431
rect 13766 -25499 13778 -25465
rect 13812 -25499 13824 -25465
rect 13766 -25533 13824 -25499
rect 13766 -25567 13778 -25533
rect 13812 -25567 13824 -25533
rect 13766 -25601 13824 -25567
rect 13766 -25635 13778 -25601
rect 13812 -25635 13824 -25601
rect 13766 -25669 13824 -25635
rect 13766 -25703 13778 -25669
rect 13812 -25703 13824 -25669
rect 13766 -25737 13824 -25703
rect 13766 -25771 13778 -25737
rect 13812 -25771 13824 -25737
rect 13766 -25805 13824 -25771
rect 13766 -25839 13778 -25805
rect 13812 -25839 13824 -25805
rect 13766 -25884 13824 -25839
rect 14784 -25329 14842 -25284
rect 14784 -25363 14796 -25329
rect 14830 -25363 14842 -25329
rect 14784 -25397 14842 -25363
rect 14784 -25431 14796 -25397
rect 14830 -25431 14842 -25397
rect 14784 -25465 14842 -25431
rect 14784 -25499 14796 -25465
rect 14830 -25499 14842 -25465
rect 14784 -25533 14842 -25499
rect 14784 -25567 14796 -25533
rect 14830 -25567 14842 -25533
rect 14784 -25601 14842 -25567
rect 14784 -25635 14796 -25601
rect 14830 -25635 14842 -25601
rect 14784 -25669 14842 -25635
rect 14784 -25703 14796 -25669
rect 14830 -25703 14842 -25669
rect 14784 -25737 14842 -25703
rect 14784 -25771 14796 -25737
rect 14830 -25771 14842 -25737
rect 14784 -25805 14842 -25771
rect 14784 -25839 14796 -25805
rect 14830 -25839 14842 -25805
rect 14784 -25884 14842 -25839
rect 15802 -25329 15860 -25284
rect 15802 -25363 15814 -25329
rect 15848 -25363 15860 -25329
rect 15802 -25397 15860 -25363
rect 15802 -25431 15814 -25397
rect 15848 -25431 15860 -25397
rect 15802 -25465 15860 -25431
rect 15802 -25499 15814 -25465
rect 15848 -25499 15860 -25465
rect 15802 -25533 15860 -25499
rect 15802 -25567 15814 -25533
rect 15848 -25567 15860 -25533
rect 15802 -25601 15860 -25567
rect 15802 -25635 15814 -25601
rect 15848 -25635 15860 -25601
rect 15802 -25669 15860 -25635
rect 15802 -25703 15814 -25669
rect 15848 -25703 15860 -25669
rect 15802 -25737 15860 -25703
rect 15802 -25771 15814 -25737
rect 15848 -25771 15860 -25737
rect 15802 -25805 15860 -25771
rect 15802 -25839 15814 -25805
rect 15848 -25839 15860 -25805
rect 15802 -25884 15860 -25839
rect 16820 -25329 16878 -25284
rect 16820 -25363 16832 -25329
rect 16866 -25363 16878 -25329
rect 16820 -25397 16878 -25363
rect 16820 -25431 16832 -25397
rect 16866 -25431 16878 -25397
rect 16820 -25465 16878 -25431
rect 16820 -25499 16832 -25465
rect 16866 -25499 16878 -25465
rect 16820 -25533 16878 -25499
rect 16820 -25567 16832 -25533
rect 16866 -25567 16878 -25533
rect 16820 -25601 16878 -25567
rect 16820 -25635 16832 -25601
rect 16866 -25635 16878 -25601
rect 16820 -25669 16878 -25635
rect 16820 -25703 16832 -25669
rect 16866 -25703 16878 -25669
rect 16820 -25737 16878 -25703
rect 16820 -25771 16832 -25737
rect 16866 -25771 16878 -25737
rect 16820 -25805 16878 -25771
rect 16820 -25839 16832 -25805
rect 16866 -25839 16878 -25805
rect 16820 -25884 16878 -25839
rect 17838 -25329 17896 -25284
rect 17838 -25363 17850 -25329
rect 17884 -25363 17896 -25329
rect 17838 -25397 17896 -25363
rect 17838 -25431 17850 -25397
rect 17884 -25431 17896 -25397
rect 17838 -25465 17896 -25431
rect 17838 -25499 17850 -25465
rect 17884 -25499 17896 -25465
rect 17838 -25533 17896 -25499
rect 17838 -25567 17850 -25533
rect 17884 -25567 17896 -25533
rect 17838 -25601 17896 -25567
rect 17838 -25635 17850 -25601
rect 17884 -25635 17896 -25601
rect 17838 -25669 17896 -25635
rect 17838 -25703 17850 -25669
rect 17884 -25703 17896 -25669
rect 17838 -25737 17896 -25703
rect 17838 -25771 17850 -25737
rect 17884 -25771 17896 -25737
rect 17838 -25805 17896 -25771
rect 17838 -25839 17850 -25805
rect 17884 -25839 17896 -25805
rect 17838 -25884 17896 -25839
rect 18856 -25329 18914 -25284
rect 18856 -25363 18868 -25329
rect 18902 -25363 18914 -25329
rect 18856 -25397 18914 -25363
rect 18856 -25431 18868 -25397
rect 18902 -25431 18914 -25397
rect 18856 -25465 18914 -25431
rect 18856 -25499 18868 -25465
rect 18902 -25499 18914 -25465
rect 18856 -25533 18914 -25499
rect 18856 -25567 18868 -25533
rect 18902 -25567 18914 -25533
rect 18856 -25601 18914 -25567
rect 18856 -25635 18868 -25601
rect 18902 -25635 18914 -25601
rect 18856 -25669 18914 -25635
rect 18856 -25703 18868 -25669
rect 18902 -25703 18914 -25669
rect 18856 -25737 18914 -25703
rect 18856 -25771 18868 -25737
rect 18902 -25771 18914 -25737
rect 18856 -25805 18914 -25771
rect 18856 -25839 18868 -25805
rect 18902 -25839 18914 -25805
rect 18856 -25884 18914 -25839
rect 19874 -25329 19932 -25284
rect 19874 -25363 19886 -25329
rect 19920 -25363 19932 -25329
rect 19874 -25397 19932 -25363
rect 19874 -25431 19886 -25397
rect 19920 -25431 19932 -25397
rect 19874 -25465 19932 -25431
rect 19874 -25499 19886 -25465
rect 19920 -25499 19932 -25465
rect 19874 -25533 19932 -25499
rect 19874 -25567 19886 -25533
rect 19920 -25567 19932 -25533
rect 19874 -25601 19932 -25567
rect 19874 -25635 19886 -25601
rect 19920 -25635 19932 -25601
rect 19874 -25669 19932 -25635
rect 19874 -25703 19886 -25669
rect 19920 -25703 19932 -25669
rect 19874 -25737 19932 -25703
rect 19874 -25771 19886 -25737
rect 19920 -25771 19932 -25737
rect 19874 -25805 19932 -25771
rect 19874 -25839 19886 -25805
rect 19920 -25839 19932 -25805
rect 19874 -25884 19932 -25839
rect 20892 -25329 20950 -25284
rect 20892 -25363 20904 -25329
rect 20938 -25363 20950 -25329
rect 20892 -25397 20950 -25363
rect 20892 -25431 20904 -25397
rect 20938 -25431 20950 -25397
rect 20892 -25465 20950 -25431
rect 20892 -25499 20904 -25465
rect 20938 -25499 20950 -25465
rect 20892 -25533 20950 -25499
rect 20892 -25567 20904 -25533
rect 20938 -25567 20950 -25533
rect 20892 -25601 20950 -25567
rect 20892 -25635 20904 -25601
rect 20938 -25635 20950 -25601
rect 20892 -25669 20950 -25635
rect 20892 -25703 20904 -25669
rect 20938 -25703 20950 -25669
rect 20892 -25737 20950 -25703
rect 20892 -25771 20904 -25737
rect 20938 -25771 20950 -25737
rect 20892 -25805 20950 -25771
rect 20892 -25839 20904 -25805
rect 20938 -25839 20950 -25805
rect 20892 -25884 20950 -25839
rect 21910 -25329 21968 -25284
rect 21910 -25363 21922 -25329
rect 21956 -25363 21968 -25329
rect 21910 -25397 21968 -25363
rect 21910 -25431 21922 -25397
rect 21956 -25431 21968 -25397
rect 21910 -25465 21968 -25431
rect 21910 -25499 21922 -25465
rect 21956 -25499 21968 -25465
rect 21910 -25533 21968 -25499
rect 21910 -25567 21922 -25533
rect 21956 -25567 21968 -25533
rect 21910 -25601 21968 -25567
rect 21910 -25635 21922 -25601
rect 21956 -25635 21968 -25601
rect 21910 -25669 21968 -25635
rect 21910 -25703 21922 -25669
rect 21956 -25703 21968 -25669
rect 21910 -25737 21968 -25703
rect 21910 -25771 21922 -25737
rect 21956 -25771 21968 -25737
rect 21910 -25805 21968 -25771
rect 21910 -25839 21922 -25805
rect 21956 -25839 21968 -25805
rect 21910 -25884 21968 -25839
rect 22928 -25329 22986 -25284
rect 22928 -25363 22940 -25329
rect 22974 -25363 22986 -25329
rect 22928 -25397 22986 -25363
rect 22928 -25431 22940 -25397
rect 22974 -25431 22986 -25397
rect 22928 -25465 22986 -25431
rect 22928 -25499 22940 -25465
rect 22974 -25499 22986 -25465
rect 22928 -25533 22986 -25499
rect 22928 -25567 22940 -25533
rect 22974 -25567 22986 -25533
rect 22928 -25601 22986 -25567
rect 22928 -25635 22940 -25601
rect 22974 -25635 22986 -25601
rect 22928 -25669 22986 -25635
rect 22928 -25703 22940 -25669
rect 22974 -25703 22986 -25669
rect 22928 -25737 22986 -25703
rect 22928 -25771 22940 -25737
rect 22974 -25771 22986 -25737
rect 22928 -25805 22986 -25771
rect 22928 -25839 22940 -25805
rect 22974 -25839 22986 -25805
rect 22928 -25884 22986 -25839
<< pdiff >>
rect 3614 -4703 3672 -4690
rect 3614 -4737 3626 -4703
rect 3660 -4737 3672 -4703
rect 3614 -4771 3672 -4737
rect 3614 -4805 3626 -4771
rect 3660 -4805 3672 -4771
rect 3614 -4839 3672 -4805
rect 3614 -4873 3626 -4839
rect 3660 -4873 3672 -4839
rect 3614 -4907 3672 -4873
rect 3614 -4941 3626 -4907
rect 3660 -4941 3672 -4907
rect 3614 -4975 3672 -4941
rect 3614 -5009 3626 -4975
rect 3660 -5009 3672 -4975
rect 3614 -5043 3672 -5009
rect 3614 -5077 3626 -5043
rect 3660 -5077 3672 -5043
rect 3614 -5090 3672 -5077
rect 3832 -4703 3890 -4690
rect 3832 -4737 3844 -4703
rect 3878 -4737 3890 -4703
rect 3832 -4771 3890 -4737
rect 3832 -4805 3844 -4771
rect 3878 -4805 3890 -4771
rect 3832 -4839 3890 -4805
rect 3832 -4873 3844 -4839
rect 3878 -4873 3890 -4839
rect 3832 -4907 3890 -4873
rect 3832 -4941 3844 -4907
rect 3878 -4941 3890 -4907
rect 3832 -4975 3890 -4941
rect 3832 -5009 3844 -4975
rect 3878 -5009 3890 -4975
rect 3832 -5043 3890 -5009
rect 3832 -5077 3844 -5043
rect 3878 -5077 3890 -5043
rect 3832 -5090 3890 -5077
rect 4050 -4703 4108 -4690
rect 4050 -4737 4062 -4703
rect 4096 -4737 4108 -4703
rect 4050 -4771 4108 -4737
rect 4050 -4805 4062 -4771
rect 4096 -4805 4108 -4771
rect 4050 -4839 4108 -4805
rect 4050 -4873 4062 -4839
rect 4096 -4873 4108 -4839
rect 4050 -4907 4108 -4873
rect 4050 -4941 4062 -4907
rect 4096 -4941 4108 -4907
rect 4050 -4975 4108 -4941
rect 4050 -5009 4062 -4975
rect 4096 -5009 4108 -4975
rect 4050 -5043 4108 -5009
rect 4050 -5077 4062 -5043
rect 4096 -5077 4108 -5043
rect 4050 -5090 4108 -5077
rect 4268 -4703 4326 -4690
rect 4268 -4737 4280 -4703
rect 4314 -4737 4326 -4703
rect 4268 -4771 4326 -4737
rect 4268 -4805 4280 -4771
rect 4314 -4805 4326 -4771
rect 4268 -4839 4326 -4805
rect 4268 -4873 4280 -4839
rect 4314 -4873 4326 -4839
rect 4268 -4907 4326 -4873
rect 4268 -4941 4280 -4907
rect 4314 -4941 4326 -4907
rect 4268 -4975 4326 -4941
rect 4268 -5009 4280 -4975
rect 4314 -5009 4326 -4975
rect 4268 -5043 4326 -5009
rect 4268 -5077 4280 -5043
rect 4314 -5077 4326 -5043
rect 4268 -5090 4326 -5077
rect 4486 -4703 4544 -4690
rect 4486 -4737 4498 -4703
rect 4532 -4737 4544 -4703
rect 4486 -4771 4544 -4737
rect 4486 -4805 4498 -4771
rect 4532 -4805 4544 -4771
rect 4486 -4839 4544 -4805
rect 4486 -4873 4498 -4839
rect 4532 -4873 4544 -4839
rect 4486 -4907 4544 -4873
rect 4486 -4941 4498 -4907
rect 4532 -4941 4544 -4907
rect 4486 -4975 4544 -4941
rect 4486 -5009 4498 -4975
rect 4532 -5009 4544 -4975
rect 4486 -5043 4544 -5009
rect 4486 -5077 4498 -5043
rect 4532 -5077 4544 -5043
rect 4486 -5090 4544 -5077
rect 4704 -4703 4762 -4690
rect 4704 -4737 4716 -4703
rect 4750 -4737 4762 -4703
rect 4704 -4771 4762 -4737
rect 4704 -4805 4716 -4771
rect 4750 -4805 4762 -4771
rect 4704 -4839 4762 -4805
rect 4704 -4873 4716 -4839
rect 4750 -4873 4762 -4839
rect 4704 -4907 4762 -4873
rect 4704 -4941 4716 -4907
rect 4750 -4941 4762 -4907
rect 4704 -4975 4762 -4941
rect 4704 -5009 4716 -4975
rect 4750 -5009 4762 -4975
rect 4704 -5043 4762 -5009
rect 4704 -5077 4716 -5043
rect 4750 -5077 4762 -5043
rect 4704 -5090 4762 -5077
rect 4922 -4703 4980 -4690
rect 4922 -4737 4934 -4703
rect 4968 -4737 4980 -4703
rect 4922 -4771 4980 -4737
rect 4922 -4805 4934 -4771
rect 4968 -4805 4980 -4771
rect 4922 -4839 4980 -4805
rect 4922 -4873 4934 -4839
rect 4968 -4873 4980 -4839
rect 4922 -4907 4980 -4873
rect 4922 -4941 4934 -4907
rect 4968 -4941 4980 -4907
rect 4922 -4975 4980 -4941
rect 4922 -5009 4934 -4975
rect 4968 -5009 4980 -4975
rect 4922 -5043 4980 -5009
rect 4922 -5077 4934 -5043
rect 4968 -5077 4980 -5043
rect 4922 -5090 4980 -5077
rect 5140 -4703 5198 -4690
rect 5140 -4737 5152 -4703
rect 5186 -4737 5198 -4703
rect 5140 -4771 5198 -4737
rect 5140 -4805 5152 -4771
rect 5186 -4805 5198 -4771
rect 5140 -4839 5198 -4805
rect 5140 -4873 5152 -4839
rect 5186 -4873 5198 -4839
rect 5140 -4907 5198 -4873
rect 5140 -4941 5152 -4907
rect 5186 -4941 5198 -4907
rect 5140 -4975 5198 -4941
rect 5140 -5009 5152 -4975
rect 5186 -5009 5198 -4975
rect 5140 -5043 5198 -5009
rect 5140 -5077 5152 -5043
rect 5186 -5077 5198 -5043
rect 5140 -5090 5198 -5077
rect 5358 -4703 5416 -4690
rect 5358 -4737 5370 -4703
rect 5404 -4737 5416 -4703
rect 5358 -4771 5416 -4737
rect 5358 -4805 5370 -4771
rect 5404 -4805 5416 -4771
rect 5358 -4839 5416 -4805
rect 5358 -4873 5370 -4839
rect 5404 -4873 5416 -4839
rect 5358 -4907 5416 -4873
rect 5358 -4941 5370 -4907
rect 5404 -4941 5416 -4907
rect 5358 -4975 5416 -4941
rect 5358 -5009 5370 -4975
rect 5404 -5009 5416 -4975
rect 5358 -5043 5416 -5009
rect 5358 -5077 5370 -5043
rect 5404 -5077 5416 -5043
rect 5358 -5090 5416 -5077
rect 5576 -4703 5634 -4690
rect 5576 -4737 5588 -4703
rect 5622 -4737 5634 -4703
rect 5576 -4771 5634 -4737
rect 5576 -4805 5588 -4771
rect 5622 -4805 5634 -4771
rect 5576 -4839 5634 -4805
rect 5576 -4873 5588 -4839
rect 5622 -4873 5634 -4839
rect 5576 -4907 5634 -4873
rect 5576 -4941 5588 -4907
rect 5622 -4941 5634 -4907
rect 5576 -4975 5634 -4941
rect 5576 -5009 5588 -4975
rect 5622 -5009 5634 -4975
rect 5576 -5043 5634 -5009
rect 5576 -5077 5588 -5043
rect 5622 -5077 5634 -5043
rect 5576 -5090 5634 -5077
rect 5794 -4703 5852 -4690
rect 5794 -4737 5806 -4703
rect 5840 -4737 5852 -4703
rect 5794 -4771 5852 -4737
rect 5794 -4805 5806 -4771
rect 5840 -4805 5852 -4771
rect 5794 -4839 5852 -4805
rect 5794 -4873 5806 -4839
rect 5840 -4873 5852 -4839
rect 5794 -4907 5852 -4873
rect 5794 -4941 5806 -4907
rect 5840 -4941 5852 -4907
rect 5794 -4975 5852 -4941
rect 5794 -5009 5806 -4975
rect 5840 -5009 5852 -4975
rect 5794 -5043 5852 -5009
rect 5794 -5077 5806 -5043
rect 5840 -5077 5852 -5043
rect 5794 -5090 5852 -5077
rect 3614 -5641 3672 -5628
rect 3614 -5675 3626 -5641
rect 3660 -5675 3672 -5641
rect 3614 -5709 3672 -5675
rect 3614 -5743 3626 -5709
rect 3660 -5743 3672 -5709
rect 3614 -5777 3672 -5743
rect 3614 -5811 3626 -5777
rect 3660 -5811 3672 -5777
rect 3614 -5845 3672 -5811
rect 3614 -5879 3626 -5845
rect 3660 -5879 3672 -5845
rect 3614 -5913 3672 -5879
rect 3614 -5947 3626 -5913
rect 3660 -5947 3672 -5913
rect 3614 -5981 3672 -5947
rect 3614 -6015 3626 -5981
rect 3660 -6015 3672 -5981
rect 3614 -6028 3672 -6015
rect 3832 -5641 3890 -5628
rect 3832 -5675 3844 -5641
rect 3878 -5675 3890 -5641
rect 3832 -5709 3890 -5675
rect 3832 -5743 3844 -5709
rect 3878 -5743 3890 -5709
rect 3832 -5777 3890 -5743
rect 3832 -5811 3844 -5777
rect 3878 -5811 3890 -5777
rect 3832 -5845 3890 -5811
rect 3832 -5879 3844 -5845
rect 3878 -5879 3890 -5845
rect 3832 -5913 3890 -5879
rect 3832 -5947 3844 -5913
rect 3878 -5947 3890 -5913
rect 3832 -5981 3890 -5947
rect 3832 -6015 3844 -5981
rect 3878 -6015 3890 -5981
rect 3832 -6028 3890 -6015
rect 4050 -5641 4108 -5628
rect 4050 -5675 4062 -5641
rect 4096 -5675 4108 -5641
rect 4050 -5709 4108 -5675
rect 4050 -5743 4062 -5709
rect 4096 -5743 4108 -5709
rect 4050 -5777 4108 -5743
rect 4050 -5811 4062 -5777
rect 4096 -5811 4108 -5777
rect 4050 -5845 4108 -5811
rect 4050 -5879 4062 -5845
rect 4096 -5879 4108 -5845
rect 4050 -5913 4108 -5879
rect 4050 -5947 4062 -5913
rect 4096 -5947 4108 -5913
rect 4050 -5981 4108 -5947
rect 4050 -6015 4062 -5981
rect 4096 -6015 4108 -5981
rect 4050 -6028 4108 -6015
rect 4268 -5641 4326 -5628
rect 4268 -5675 4280 -5641
rect 4314 -5675 4326 -5641
rect 4268 -5709 4326 -5675
rect 4268 -5743 4280 -5709
rect 4314 -5743 4326 -5709
rect 4268 -5777 4326 -5743
rect 4268 -5811 4280 -5777
rect 4314 -5811 4326 -5777
rect 4268 -5845 4326 -5811
rect 4268 -5879 4280 -5845
rect 4314 -5879 4326 -5845
rect 4268 -5913 4326 -5879
rect 4268 -5947 4280 -5913
rect 4314 -5947 4326 -5913
rect 4268 -5981 4326 -5947
rect 4268 -6015 4280 -5981
rect 4314 -6015 4326 -5981
rect 4268 -6028 4326 -6015
rect 4486 -5641 4544 -5628
rect 4486 -5675 4498 -5641
rect 4532 -5675 4544 -5641
rect 4486 -5709 4544 -5675
rect 4486 -5743 4498 -5709
rect 4532 -5743 4544 -5709
rect 4486 -5777 4544 -5743
rect 4486 -5811 4498 -5777
rect 4532 -5811 4544 -5777
rect 4486 -5845 4544 -5811
rect 4486 -5879 4498 -5845
rect 4532 -5879 4544 -5845
rect 4486 -5913 4544 -5879
rect 4486 -5947 4498 -5913
rect 4532 -5947 4544 -5913
rect 4486 -5981 4544 -5947
rect 4486 -6015 4498 -5981
rect 4532 -6015 4544 -5981
rect 4486 -6028 4544 -6015
rect 4704 -5641 4762 -5628
rect 4704 -5675 4716 -5641
rect 4750 -5675 4762 -5641
rect 4704 -5709 4762 -5675
rect 4704 -5743 4716 -5709
rect 4750 -5743 4762 -5709
rect 4704 -5777 4762 -5743
rect 4704 -5811 4716 -5777
rect 4750 -5811 4762 -5777
rect 4704 -5845 4762 -5811
rect 4704 -5879 4716 -5845
rect 4750 -5879 4762 -5845
rect 4704 -5913 4762 -5879
rect 4704 -5947 4716 -5913
rect 4750 -5947 4762 -5913
rect 4704 -5981 4762 -5947
rect 4704 -6015 4716 -5981
rect 4750 -6015 4762 -5981
rect 4704 -6028 4762 -6015
rect 4922 -5641 4980 -5628
rect 4922 -5675 4934 -5641
rect 4968 -5675 4980 -5641
rect 4922 -5709 4980 -5675
rect 4922 -5743 4934 -5709
rect 4968 -5743 4980 -5709
rect 4922 -5777 4980 -5743
rect 4922 -5811 4934 -5777
rect 4968 -5811 4980 -5777
rect 4922 -5845 4980 -5811
rect 4922 -5879 4934 -5845
rect 4968 -5879 4980 -5845
rect 4922 -5913 4980 -5879
rect 4922 -5947 4934 -5913
rect 4968 -5947 4980 -5913
rect 4922 -5981 4980 -5947
rect 4922 -6015 4934 -5981
rect 4968 -6015 4980 -5981
rect 4922 -6028 4980 -6015
rect 5140 -5641 5198 -5628
rect 5140 -5675 5152 -5641
rect 5186 -5675 5198 -5641
rect 5140 -5709 5198 -5675
rect 5140 -5743 5152 -5709
rect 5186 -5743 5198 -5709
rect 5140 -5777 5198 -5743
rect 5140 -5811 5152 -5777
rect 5186 -5811 5198 -5777
rect 5140 -5845 5198 -5811
rect 5140 -5879 5152 -5845
rect 5186 -5879 5198 -5845
rect 5140 -5913 5198 -5879
rect 5140 -5947 5152 -5913
rect 5186 -5947 5198 -5913
rect 5140 -5981 5198 -5947
rect 5140 -6015 5152 -5981
rect 5186 -6015 5198 -5981
rect 5140 -6028 5198 -6015
rect 5358 -5641 5416 -5628
rect 5358 -5675 5370 -5641
rect 5404 -5675 5416 -5641
rect 5358 -5709 5416 -5675
rect 5358 -5743 5370 -5709
rect 5404 -5743 5416 -5709
rect 5358 -5777 5416 -5743
rect 5358 -5811 5370 -5777
rect 5404 -5811 5416 -5777
rect 5358 -5845 5416 -5811
rect 5358 -5879 5370 -5845
rect 5404 -5879 5416 -5845
rect 5358 -5913 5416 -5879
rect 5358 -5947 5370 -5913
rect 5404 -5947 5416 -5913
rect 5358 -5981 5416 -5947
rect 5358 -6015 5370 -5981
rect 5404 -6015 5416 -5981
rect 5358 -6028 5416 -6015
rect 5576 -5641 5634 -5628
rect 5576 -5675 5588 -5641
rect 5622 -5675 5634 -5641
rect 5576 -5709 5634 -5675
rect 5576 -5743 5588 -5709
rect 5622 -5743 5634 -5709
rect 5576 -5777 5634 -5743
rect 5576 -5811 5588 -5777
rect 5622 -5811 5634 -5777
rect 5576 -5845 5634 -5811
rect 5576 -5879 5588 -5845
rect 5622 -5879 5634 -5845
rect 5576 -5913 5634 -5879
rect 5576 -5947 5588 -5913
rect 5622 -5947 5634 -5913
rect 5576 -5981 5634 -5947
rect 5576 -6015 5588 -5981
rect 5622 -6015 5634 -5981
rect 5576 -6028 5634 -6015
rect 5794 -5641 5852 -5628
rect 5794 -5675 5806 -5641
rect 5840 -5675 5852 -5641
rect 5794 -5709 5852 -5675
rect 5794 -5743 5806 -5709
rect 5840 -5743 5852 -5709
rect 5794 -5777 5852 -5743
rect 5794 -5811 5806 -5777
rect 5840 -5811 5852 -5777
rect 5794 -5845 5852 -5811
rect 5794 -5879 5806 -5845
rect 5840 -5879 5852 -5845
rect 5794 -5913 5852 -5879
rect 5794 -5947 5806 -5913
rect 5840 -5947 5852 -5913
rect 5794 -5981 5852 -5947
rect 5794 -6015 5806 -5981
rect 5840 -6015 5852 -5981
rect 5794 -6028 5852 -6015
rect 3614 -6579 3672 -6566
rect 3614 -6613 3626 -6579
rect 3660 -6613 3672 -6579
rect 3614 -6647 3672 -6613
rect 3614 -6681 3626 -6647
rect 3660 -6681 3672 -6647
rect 3614 -6715 3672 -6681
rect 3614 -6749 3626 -6715
rect 3660 -6749 3672 -6715
rect 3614 -6783 3672 -6749
rect 3614 -6817 3626 -6783
rect 3660 -6817 3672 -6783
rect 3614 -6851 3672 -6817
rect 3614 -6885 3626 -6851
rect 3660 -6885 3672 -6851
rect 3614 -6919 3672 -6885
rect 3614 -6953 3626 -6919
rect 3660 -6953 3672 -6919
rect 3614 -6966 3672 -6953
rect 3832 -6579 3890 -6566
rect 3832 -6613 3844 -6579
rect 3878 -6613 3890 -6579
rect 3832 -6647 3890 -6613
rect 3832 -6681 3844 -6647
rect 3878 -6681 3890 -6647
rect 3832 -6715 3890 -6681
rect 3832 -6749 3844 -6715
rect 3878 -6749 3890 -6715
rect 3832 -6783 3890 -6749
rect 3832 -6817 3844 -6783
rect 3878 -6817 3890 -6783
rect 3832 -6851 3890 -6817
rect 3832 -6885 3844 -6851
rect 3878 -6885 3890 -6851
rect 3832 -6919 3890 -6885
rect 3832 -6953 3844 -6919
rect 3878 -6953 3890 -6919
rect 3832 -6966 3890 -6953
rect 4050 -6579 4108 -6566
rect 4050 -6613 4062 -6579
rect 4096 -6613 4108 -6579
rect 4050 -6647 4108 -6613
rect 4050 -6681 4062 -6647
rect 4096 -6681 4108 -6647
rect 4050 -6715 4108 -6681
rect 4050 -6749 4062 -6715
rect 4096 -6749 4108 -6715
rect 4050 -6783 4108 -6749
rect 4050 -6817 4062 -6783
rect 4096 -6817 4108 -6783
rect 4050 -6851 4108 -6817
rect 4050 -6885 4062 -6851
rect 4096 -6885 4108 -6851
rect 4050 -6919 4108 -6885
rect 4050 -6953 4062 -6919
rect 4096 -6953 4108 -6919
rect 4050 -6966 4108 -6953
rect 4268 -6579 4326 -6566
rect 4268 -6613 4280 -6579
rect 4314 -6613 4326 -6579
rect 4268 -6647 4326 -6613
rect 4268 -6681 4280 -6647
rect 4314 -6681 4326 -6647
rect 4268 -6715 4326 -6681
rect 4268 -6749 4280 -6715
rect 4314 -6749 4326 -6715
rect 4268 -6783 4326 -6749
rect 4268 -6817 4280 -6783
rect 4314 -6817 4326 -6783
rect 4268 -6851 4326 -6817
rect 4268 -6885 4280 -6851
rect 4314 -6885 4326 -6851
rect 4268 -6919 4326 -6885
rect 4268 -6953 4280 -6919
rect 4314 -6953 4326 -6919
rect 4268 -6966 4326 -6953
rect 4486 -6579 4544 -6566
rect 4486 -6613 4498 -6579
rect 4532 -6613 4544 -6579
rect 4486 -6647 4544 -6613
rect 4486 -6681 4498 -6647
rect 4532 -6681 4544 -6647
rect 4486 -6715 4544 -6681
rect 4486 -6749 4498 -6715
rect 4532 -6749 4544 -6715
rect 4486 -6783 4544 -6749
rect 4486 -6817 4498 -6783
rect 4532 -6817 4544 -6783
rect 4486 -6851 4544 -6817
rect 4486 -6885 4498 -6851
rect 4532 -6885 4544 -6851
rect 4486 -6919 4544 -6885
rect 4486 -6953 4498 -6919
rect 4532 -6953 4544 -6919
rect 4486 -6966 4544 -6953
rect 4704 -6579 4762 -6566
rect 4704 -6613 4716 -6579
rect 4750 -6613 4762 -6579
rect 4704 -6647 4762 -6613
rect 4704 -6681 4716 -6647
rect 4750 -6681 4762 -6647
rect 4704 -6715 4762 -6681
rect 4704 -6749 4716 -6715
rect 4750 -6749 4762 -6715
rect 4704 -6783 4762 -6749
rect 4704 -6817 4716 -6783
rect 4750 -6817 4762 -6783
rect 4704 -6851 4762 -6817
rect 4704 -6885 4716 -6851
rect 4750 -6885 4762 -6851
rect 4704 -6919 4762 -6885
rect 4704 -6953 4716 -6919
rect 4750 -6953 4762 -6919
rect 4704 -6966 4762 -6953
rect 4922 -6579 4980 -6566
rect 4922 -6613 4934 -6579
rect 4968 -6613 4980 -6579
rect 4922 -6647 4980 -6613
rect 4922 -6681 4934 -6647
rect 4968 -6681 4980 -6647
rect 4922 -6715 4980 -6681
rect 4922 -6749 4934 -6715
rect 4968 -6749 4980 -6715
rect 4922 -6783 4980 -6749
rect 4922 -6817 4934 -6783
rect 4968 -6817 4980 -6783
rect 4922 -6851 4980 -6817
rect 4922 -6885 4934 -6851
rect 4968 -6885 4980 -6851
rect 4922 -6919 4980 -6885
rect 4922 -6953 4934 -6919
rect 4968 -6953 4980 -6919
rect 4922 -6966 4980 -6953
rect 5140 -6579 5198 -6566
rect 5140 -6613 5152 -6579
rect 5186 -6613 5198 -6579
rect 5140 -6647 5198 -6613
rect 5140 -6681 5152 -6647
rect 5186 -6681 5198 -6647
rect 5140 -6715 5198 -6681
rect 5140 -6749 5152 -6715
rect 5186 -6749 5198 -6715
rect 5140 -6783 5198 -6749
rect 5140 -6817 5152 -6783
rect 5186 -6817 5198 -6783
rect 5140 -6851 5198 -6817
rect 5140 -6885 5152 -6851
rect 5186 -6885 5198 -6851
rect 5140 -6919 5198 -6885
rect 5140 -6953 5152 -6919
rect 5186 -6953 5198 -6919
rect 5140 -6966 5198 -6953
rect 5358 -6579 5416 -6566
rect 5358 -6613 5370 -6579
rect 5404 -6613 5416 -6579
rect 5358 -6647 5416 -6613
rect 5358 -6681 5370 -6647
rect 5404 -6681 5416 -6647
rect 5358 -6715 5416 -6681
rect 5358 -6749 5370 -6715
rect 5404 -6749 5416 -6715
rect 5358 -6783 5416 -6749
rect 5358 -6817 5370 -6783
rect 5404 -6817 5416 -6783
rect 5358 -6851 5416 -6817
rect 5358 -6885 5370 -6851
rect 5404 -6885 5416 -6851
rect 5358 -6919 5416 -6885
rect 5358 -6953 5370 -6919
rect 5404 -6953 5416 -6919
rect 5358 -6966 5416 -6953
rect 5576 -6579 5634 -6566
rect 5576 -6613 5588 -6579
rect 5622 -6613 5634 -6579
rect 5576 -6647 5634 -6613
rect 5576 -6681 5588 -6647
rect 5622 -6681 5634 -6647
rect 5576 -6715 5634 -6681
rect 5576 -6749 5588 -6715
rect 5622 -6749 5634 -6715
rect 5576 -6783 5634 -6749
rect 5576 -6817 5588 -6783
rect 5622 -6817 5634 -6783
rect 5576 -6851 5634 -6817
rect 5576 -6885 5588 -6851
rect 5622 -6885 5634 -6851
rect 5576 -6919 5634 -6885
rect 5576 -6953 5588 -6919
rect 5622 -6953 5634 -6919
rect 5576 -6966 5634 -6953
rect 5794 -6579 5852 -6566
rect 5794 -6613 5806 -6579
rect 5840 -6613 5852 -6579
rect 5794 -6647 5852 -6613
rect 5794 -6681 5806 -6647
rect 5840 -6681 5852 -6647
rect 5794 -6715 5852 -6681
rect 5794 -6749 5806 -6715
rect 5840 -6749 5852 -6715
rect 5794 -6783 5852 -6749
rect 5794 -6817 5806 -6783
rect 5840 -6817 5852 -6783
rect 5794 -6851 5852 -6817
rect 5794 -6885 5806 -6851
rect 5840 -6885 5852 -6851
rect 5794 -6919 5852 -6885
rect 5794 -6953 5806 -6919
rect 5840 -6953 5852 -6919
rect 5794 -6966 5852 -6953
rect 3614 -7517 3672 -7504
rect 3614 -7551 3626 -7517
rect 3660 -7551 3672 -7517
rect 3614 -7585 3672 -7551
rect 3614 -7619 3626 -7585
rect 3660 -7619 3672 -7585
rect 3614 -7653 3672 -7619
rect 3614 -7687 3626 -7653
rect 3660 -7687 3672 -7653
rect 3614 -7721 3672 -7687
rect 3614 -7755 3626 -7721
rect 3660 -7755 3672 -7721
rect 3614 -7789 3672 -7755
rect 3614 -7823 3626 -7789
rect 3660 -7823 3672 -7789
rect 3614 -7857 3672 -7823
rect 3614 -7891 3626 -7857
rect 3660 -7891 3672 -7857
rect 3614 -7904 3672 -7891
rect 3832 -7517 3890 -7504
rect 3832 -7551 3844 -7517
rect 3878 -7551 3890 -7517
rect 3832 -7585 3890 -7551
rect 3832 -7619 3844 -7585
rect 3878 -7619 3890 -7585
rect 3832 -7653 3890 -7619
rect 3832 -7687 3844 -7653
rect 3878 -7687 3890 -7653
rect 3832 -7721 3890 -7687
rect 3832 -7755 3844 -7721
rect 3878 -7755 3890 -7721
rect 3832 -7789 3890 -7755
rect 3832 -7823 3844 -7789
rect 3878 -7823 3890 -7789
rect 3832 -7857 3890 -7823
rect 3832 -7891 3844 -7857
rect 3878 -7891 3890 -7857
rect 3832 -7904 3890 -7891
rect 4050 -7517 4108 -7504
rect 4050 -7551 4062 -7517
rect 4096 -7551 4108 -7517
rect 4050 -7585 4108 -7551
rect 4050 -7619 4062 -7585
rect 4096 -7619 4108 -7585
rect 4050 -7653 4108 -7619
rect 4050 -7687 4062 -7653
rect 4096 -7687 4108 -7653
rect 4050 -7721 4108 -7687
rect 4050 -7755 4062 -7721
rect 4096 -7755 4108 -7721
rect 4050 -7789 4108 -7755
rect 4050 -7823 4062 -7789
rect 4096 -7823 4108 -7789
rect 4050 -7857 4108 -7823
rect 4050 -7891 4062 -7857
rect 4096 -7891 4108 -7857
rect 4050 -7904 4108 -7891
rect 4268 -7517 4326 -7504
rect 4268 -7551 4280 -7517
rect 4314 -7551 4326 -7517
rect 4268 -7585 4326 -7551
rect 4268 -7619 4280 -7585
rect 4314 -7619 4326 -7585
rect 4268 -7653 4326 -7619
rect 4268 -7687 4280 -7653
rect 4314 -7687 4326 -7653
rect 4268 -7721 4326 -7687
rect 4268 -7755 4280 -7721
rect 4314 -7755 4326 -7721
rect 4268 -7789 4326 -7755
rect 4268 -7823 4280 -7789
rect 4314 -7823 4326 -7789
rect 4268 -7857 4326 -7823
rect 4268 -7891 4280 -7857
rect 4314 -7891 4326 -7857
rect 4268 -7904 4326 -7891
rect 4486 -7517 4544 -7504
rect 4486 -7551 4498 -7517
rect 4532 -7551 4544 -7517
rect 4486 -7585 4544 -7551
rect 4486 -7619 4498 -7585
rect 4532 -7619 4544 -7585
rect 4486 -7653 4544 -7619
rect 4486 -7687 4498 -7653
rect 4532 -7687 4544 -7653
rect 4486 -7721 4544 -7687
rect 4486 -7755 4498 -7721
rect 4532 -7755 4544 -7721
rect 4486 -7789 4544 -7755
rect 4486 -7823 4498 -7789
rect 4532 -7823 4544 -7789
rect 4486 -7857 4544 -7823
rect 4486 -7891 4498 -7857
rect 4532 -7891 4544 -7857
rect 4486 -7904 4544 -7891
rect 4704 -7517 4762 -7504
rect 4704 -7551 4716 -7517
rect 4750 -7551 4762 -7517
rect 4704 -7585 4762 -7551
rect 4704 -7619 4716 -7585
rect 4750 -7619 4762 -7585
rect 4704 -7653 4762 -7619
rect 4704 -7687 4716 -7653
rect 4750 -7687 4762 -7653
rect 4704 -7721 4762 -7687
rect 4704 -7755 4716 -7721
rect 4750 -7755 4762 -7721
rect 4704 -7789 4762 -7755
rect 4704 -7823 4716 -7789
rect 4750 -7823 4762 -7789
rect 4704 -7857 4762 -7823
rect 4704 -7891 4716 -7857
rect 4750 -7891 4762 -7857
rect 4704 -7904 4762 -7891
rect 4922 -7517 4980 -7504
rect 4922 -7551 4934 -7517
rect 4968 -7551 4980 -7517
rect 4922 -7585 4980 -7551
rect 4922 -7619 4934 -7585
rect 4968 -7619 4980 -7585
rect 4922 -7653 4980 -7619
rect 4922 -7687 4934 -7653
rect 4968 -7687 4980 -7653
rect 4922 -7721 4980 -7687
rect 4922 -7755 4934 -7721
rect 4968 -7755 4980 -7721
rect 4922 -7789 4980 -7755
rect 4922 -7823 4934 -7789
rect 4968 -7823 4980 -7789
rect 4922 -7857 4980 -7823
rect 4922 -7891 4934 -7857
rect 4968 -7891 4980 -7857
rect 4922 -7904 4980 -7891
rect 5140 -7517 5198 -7504
rect 5140 -7551 5152 -7517
rect 5186 -7551 5198 -7517
rect 5140 -7585 5198 -7551
rect 5140 -7619 5152 -7585
rect 5186 -7619 5198 -7585
rect 5140 -7653 5198 -7619
rect 5140 -7687 5152 -7653
rect 5186 -7687 5198 -7653
rect 5140 -7721 5198 -7687
rect 5140 -7755 5152 -7721
rect 5186 -7755 5198 -7721
rect 5140 -7789 5198 -7755
rect 5140 -7823 5152 -7789
rect 5186 -7823 5198 -7789
rect 5140 -7857 5198 -7823
rect 5140 -7891 5152 -7857
rect 5186 -7891 5198 -7857
rect 5140 -7904 5198 -7891
rect 5358 -7517 5416 -7504
rect 5358 -7551 5370 -7517
rect 5404 -7551 5416 -7517
rect 5358 -7585 5416 -7551
rect 5358 -7619 5370 -7585
rect 5404 -7619 5416 -7585
rect 5358 -7653 5416 -7619
rect 5358 -7687 5370 -7653
rect 5404 -7687 5416 -7653
rect 5358 -7721 5416 -7687
rect 5358 -7755 5370 -7721
rect 5404 -7755 5416 -7721
rect 5358 -7789 5416 -7755
rect 5358 -7823 5370 -7789
rect 5404 -7823 5416 -7789
rect 5358 -7857 5416 -7823
rect 5358 -7891 5370 -7857
rect 5404 -7891 5416 -7857
rect 5358 -7904 5416 -7891
rect 5576 -7517 5634 -7504
rect 5576 -7551 5588 -7517
rect 5622 -7551 5634 -7517
rect 5576 -7585 5634 -7551
rect 5576 -7619 5588 -7585
rect 5622 -7619 5634 -7585
rect 5576 -7653 5634 -7619
rect 5576 -7687 5588 -7653
rect 5622 -7687 5634 -7653
rect 5576 -7721 5634 -7687
rect 5576 -7755 5588 -7721
rect 5622 -7755 5634 -7721
rect 5576 -7789 5634 -7755
rect 5576 -7823 5588 -7789
rect 5622 -7823 5634 -7789
rect 5576 -7857 5634 -7823
rect 5576 -7891 5588 -7857
rect 5622 -7891 5634 -7857
rect 5576 -7904 5634 -7891
rect 5794 -7517 5852 -7504
rect 5794 -7551 5806 -7517
rect 5840 -7551 5852 -7517
rect 5794 -7585 5852 -7551
rect 5794 -7619 5806 -7585
rect 5840 -7619 5852 -7585
rect 5794 -7653 5852 -7619
rect 5794 -7687 5806 -7653
rect 5840 -7687 5852 -7653
rect 5794 -7721 5852 -7687
rect 5794 -7755 5806 -7721
rect 5840 -7755 5852 -7721
rect 5794 -7789 5852 -7755
rect 5794 -7823 5806 -7789
rect 5840 -7823 5852 -7789
rect 5794 -7857 5852 -7823
rect 5794 -7891 5806 -7857
rect 5840 -7891 5852 -7857
rect 5794 -7904 5852 -7891
<< ndiffc >>
rect 2582 -11797 2616 -11763
rect 2582 -11865 2616 -11831
rect 2582 -11933 2616 -11899
rect 2582 -12001 2616 -11967
rect 2582 -12069 2616 -12035
rect 2582 -12137 2616 -12103
rect 2582 -12205 2616 -12171
rect 2582 -12273 2616 -12239
rect 3600 -11797 3634 -11763
rect 3600 -11865 3634 -11831
rect 3600 -11933 3634 -11899
rect 3600 -12001 3634 -11967
rect 3600 -12069 3634 -12035
rect 3600 -12137 3634 -12103
rect 3600 -12205 3634 -12171
rect 3600 -12273 3634 -12239
rect 4618 -11797 4652 -11763
rect 4618 -11865 4652 -11831
rect 4618 -11933 4652 -11899
rect 4618 -12001 4652 -11967
rect 4618 -12069 4652 -12035
rect 4618 -12137 4652 -12103
rect 4618 -12205 4652 -12171
rect 4618 -12273 4652 -12239
rect 5636 -11797 5670 -11763
rect 5636 -11865 5670 -11831
rect 5636 -11933 5670 -11899
rect 5636 -12001 5670 -11967
rect 5636 -12069 5670 -12035
rect 5636 -12137 5670 -12103
rect 5636 -12205 5670 -12171
rect 5636 -12273 5670 -12239
rect 6654 -11797 6688 -11763
rect 6654 -11865 6688 -11831
rect 6654 -11933 6688 -11899
rect 6654 -12001 6688 -11967
rect 6654 -12069 6688 -12035
rect 6654 -12137 6688 -12103
rect 6654 -12205 6688 -12171
rect 6654 -12273 6688 -12239
rect 7672 -11797 7706 -11763
rect 7672 -11865 7706 -11831
rect 7672 -11933 7706 -11899
rect 7672 -12001 7706 -11967
rect 7672 -12069 7706 -12035
rect 7672 -12137 7706 -12103
rect 7672 -12205 7706 -12171
rect 7672 -12273 7706 -12239
rect 8690 -11797 8724 -11763
rect 8690 -11865 8724 -11831
rect 8690 -11933 8724 -11899
rect 8690 -12001 8724 -11967
rect 8690 -12069 8724 -12035
rect 8690 -12137 8724 -12103
rect 8690 -12205 8724 -12171
rect 8690 -12273 8724 -12239
rect 9708 -11797 9742 -11763
rect 9708 -11865 9742 -11831
rect 9708 -11933 9742 -11899
rect 9708 -12001 9742 -11967
rect 9708 -12069 9742 -12035
rect 9708 -12137 9742 -12103
rect 9708 -12205 9742 -12171
rect 9708 -12273 9742 -12239
rect 10726 -11797 10760 -11763
rect 10726 -11865 10760 -11831
rect 10726 -11933 10760 -11899
rect 10726 -12001 10760 -11967
rect 10726 -12069 10760 -12035
rect 10726 -12137 10760 -12103
rect 10726 -12205 10760 -12171
rect 10726 -12273 10760 -12239
rect 11744 -11797 11778 -11763
rect 11744 -11865 11778 -11831
rect 11744 -11933 11778 -11899
rect 11744 -12001 11778 -11967
rect 11744 -12069 11778 -12035
rect 11744 -12137 11778 -12103
rect 11744 -12205 11778 -12171
rect 11744 -12273 11778 -12239
rect 12762 -11797 12796 -11763
rect 12762 -11865 12796 -11831
rect 12762 -11933 12796 -11899
rect 12762 -12001 12796 -11967
rect 12762 -12069 12796 -12035
rect 12762 -12137 12796 -12103
rect 12762 -12205 12796 -12171
rect 12762 -12273 12796 -12239
rect 13780 -11797 13814 -11763
rect 13780 -11865 13814 -11831
rect 13780 -11933 13814 -11899
rect 13780 -12001 13814 -11967
rect 13780 -12069 13814 -12035
rect 13780 -12137 13814 -12103
rect 13780 -12205 13814 -12171
rect 13780 -12273 13814 -12239
rect 14798 -11797 14832 -11763
rect 14798 -11865 14832 -11831
rect 14798 -11933 14832 -11899
rect 14798 -12001 14832 -11967
rect 14798 -12069 14832 -12035
rect 14798 -12137 14832 -12103
rect 14798 -12205 14832 -12171
rect 14798 -12273 14832 -12239
rect 15816 -11797 15850 -11763
rect 15816 -11865 15850 -11831
rect 15816 -11933 15850 -11899
rect 15816 -12001 15850 -11967
rect 15816 -12069 15850 -12035
rect 15816 -12137 15850 -12103
rect 15816 -12205 15850 -12171
rect 15816 -12273 15850 -12239
rect 16834 -11797 16868 -11763
rect 16834 -11865 16868 -11831
rect 16834 -11933 16868 -11899
rect 16834 -12001 16868 -11967
rect 16834 -12069 16868 -12035
rect 16834 -12137 16868 -12103
rect 16834 -12205 16868 -12171
rect 16834 -12273 16868 -12239
rect 17852 -11797 17886 -11763
rect 17852 -11865 17886 -11831
rect 17852 -11933 17886 -11899
rect 17852 -12001 17886 -11967
rect 17852 -12069 17886 -12035
rect 17852 -12137 17886 -12103
rect 17852 -12205 17886 -12171
rect 17852 -12273 17886 -12239
rect 18870 -11797 18904 -11763
rect 18870 -11865 18904 -11831
rect 18870 -11933 18904 -11899
rect 18870 -12001 18904 -11967
rect 18870 -12069 18904 -12035
rect 18870 -12137 18904 -12103
rect 18870 -12205 18904 -12171
rect 18870 -12273 18904 -12239
rect 19888 -11797 19922 -11763
rect 19888 -11865 19922 -11831
rect 19888 -11933 19922 -11899
rect 19888 -12001 19922 -11967
rect 19888 -12069 19922 -12035
rect 19888 -12137 19922 -12103
rect 19888 -12205 19922 -12171
rect 19888 -12273 19922 -12239
rect 20906 -11797 20940 -11763
rect 20906 -11865 20940 -11831
rect 20906 -11933 20940 -11899
rect 20906 -12001 20940 -11967
rect 20906 -12069 20940 -12035
rect 20906 -12137 20940 -12103
rect 20906 -12205 20940 -12171
rect 20906 -12273 20940 -12239
rect 21924 -11797 21958 -11763
rect 21924 -11865 21958 -11831
rect 21924 -11933 21958 -11899
rect 21924 -12001 21958 -11967
rect 21924 -12069 21958 -12035
rect 21924 -12137 21958 -12103
rect 21924 -12205 21958 -12171
rect 21924 -12273 21958 -12239
rect 22942 -11797 22976 -11763
rect 22942 -11865 22976 -11831
rect 22942 -11933 22976 -11899
rect 22942 -12001 22976 -11967
rect 22942 -12069 22976 -12035
rect 22942 -12137 22976 -12103
rect 22942 -12205 22976 -12171
rect 22942 -12273 22976 -12239
rect -9184 -12591 -9150 -12557
rect -9184 -12659 -9150 -12625
rect -9184 -12727 -9150 -12693
rect -9184 -12795 -9150 -12761
rect -9184 -12863 -9150 -12829
rect -9184 -12931 -9150 -12897
rect -9184 -12999 -9150 -12965
rect -9184 -13067 -9150 -13033
rect -8166 -12591 -8132 -12557
rect -8166 -12659 -8132 -12625
rect -8166 -12727 -8132 -12693
rect -8166 -12795 -8132 -12761
rect -8166 -12863 -8132 -12829
rect -8166 -12931 -8132 -12897
rect -8166 -12999 -8132 -12965
rect -8166 -13067 -8132 -13033
rect -7148 -12591 -7114 -12557
rect -7148 -12659 -7114 -12625
rect -7148 -12727 -7114 -12693
rect -7148 -12795 -7114 -12761
rect -7148 -12863 -7114 -12829
rect -7148 -12931 -7114 -12897
rect -7148 -12999 -7114 -12965
rect -7148 -13067 -7114 -13033
rect -6130 -12591 -6096 -12557
rect -6130 -12659 -6096 -12625
rect -6130 -12727 -6096 -12693
rect -6130 -12795 -6096 -12761
rect -6130 -12863 -6096 -12829
rect -6130 -12931 -6096 -12897
rect -6130 -12999 -6096 -12965
rect -6130 -13067 -6096 -13033
rect -5112 -12591 -5078 -12557
rect -5112 -12659 -5078 -12625
rect -5112 -12727 -5078 -12693
rect -5112 -12795 -5078 -12761
rect -5112 -12863 -5078 -12829
rect -5112 -12931 -5078 -12897
rect -5112 -12999 -5078 -12965
rect -5112 -13067 -5078 -13033
rect -4094 -12591 -4060 -12557
rect -4094 -12659 -4060 -12625
rect -4094 -12727 -4060 -12693
rect -4094 -12795 -4060 -12761
rect -4094 -12863 -4060 -12829
rect -4094 -12931 -4060 -12897
rect -4094 -12999 -4060 -12965
rect -4094 -13067 -4060 -13033
rect -3076 -12591 -3042 -12557
rect -3076 -12659 -3042 -12625
rect -3076 -12727 -3042 -12693
rect -3076 -12795 -3042 -12761
rect -3076 -12863 -3042 -12829
rect -3076 -12931 -3042 -12897
rect -3076 -12999 -3042 -12965
rect -3076 -13067 -3042 -13033
rect -2058 -12591 -2024 -12557
rect -2058 -12659 -2024 -12625
rect -2058 -12727 -2024 -12693
rect -2058 -12795 -2024 -12761
rect -2058 -12863 -2024 -12829
rect -2058 -12931 -2024 -12897
rect -2058 -12999 -2024 -12965
rect -2058 -13067 -2024 -13033
rect -1040 -12591 -1006 -12557
rect -1040 -12659 -1006 -12625
rect -1040 -12727 -1006 -12693
rect -1040 -12795 -1006 -12761
rect -1040 -12863 -1006 -12829
rect -1040 -12931 -1006 -12897
rect -1040 -12999 -1006 -12965
rect -1040 -13067 -1006 -13033
rect -22 -12591 12 -12557
rect -22 -12659 12 -12625
rect -22 -12727 12 -12693
rect -22 -12795 12 -12761
rect -22 -12863 12 -12829
rect -22 -12931 12 -12897
rect -22 -12999 12 -12965
rect -22 -13067 12 -13033
rect 2582 -13031 2616 -12997
rect 2582 -13099 2616 -13065
rect 2582 -13167 2616 -13133
rect 2582 -13235 2616 -13201
rect 2582 -13303 2616 -13269
rect -9184 -13409 -9150 -13375
rect -9184 -13477 -9150 -13443
rect -9184 -13545 -9150 -13511
rect -9184 -13613 -9150 -13579
rect -9184 -13681 -9150 -13647
rect -9184 -13749 -9150 -13715
rect -9184 -13817 -9150 -13783
rect -9184 -13885 -9150 -13851
rect -8166 -13409 -8132 -13375
rect -8166 -13477 -8132 -13443
rect -8166 -13545 -8132 -13511
rect -8166 -13613 -8132 -13579
rect -8166 -13681 -8132 -13647
rect -8166 -13749 -8132 -13715
rect -8166 -13817 -8132 -13783
rect -8166 -13885 -8132 -13851
rect -7148 -13409 -7114 -13375
rect -7148 -13477 -7114 -13443
rect -7148 -13545 -7114 -13511
rect -7148 -13613 -7114 -13579
rect -7148 -13681 -7114 -13647
rect -7148 -13749 -7114 -13715
rect -7148 -13817 -7114 -13783
rect -7148 -13885 -7114 -13851
rect -6130 -13409 -6096 -13375
rect -6130 -13477 -6096 -13443
rect -6130 -13545 -6096 -13511
rect -6130 -13613 -6096 -13579
rect -6130 -13681 -6096 -13647
rect -6130 -13749 -6096 -13715
rect -6130 -13817 -6096 -13783
rect -6130 -13885 -6096 -13851
rect -5112 -13409 -5078 -13375
rect -5112 -13477 -5078 -13443
rect -5112 -13545 -5078 -13511
rect -5112 -13613 -5078 -13579
rect -5112 -13681 -5078 -13647
rect -5112 -13749 -5078 -13715
rect -5112 -13817 -5078 -13783
rect -5112 -13885 -5078 -13851
rect -4094 -13409 -4060 -13375
rect -4094 -13477 -4060 -13443
rect -4094 -13545 -4060 -13511
rect -4094 -13613 -4060 -13579
rect -4094 -13681 -4060 -13647
rect -4094 -13749 -4060 -13715
rect -4094 -13817 -4060 -13783
rect -4094 -13885 -4060 -13851
rect -3076 -13409 -3042 -13375
rect -3076 -13477 -3042 -13443
rect -3076 -13545 -3042 -13511
rect -3076 -13613 -3042 -13579
rect -3076 -13681 -3042 -13647
rect -3076 -13749 -3042 -13715
rect -3076 -13817 -3042 -13783
rect -3076 -13885 -3042 -13851
rect -2058 -13409 -2024 -13375
rect -2058 -13477 -2024 -13443
rect -2058 -13545 -2024 -13511
rect -2058 -13613 -2024 -13579
rect -2058 -13681 -2024 -13647
rect -2058 -13749 -2024 -13715
rect -2058 -13817 -2024 -13783
rect -2058 -13885 -2024 -13851
rect -1040 -13409 -1006 -13375
rect -1040 -13477 -1006 -13443
rect -1040 -13545 -1006 -13511
rect -1040 -13613 -1006 -13579
rect -1040 -13681 -1006 -13647
rect -1040 -13749 -1006 -13715
rect -1040 -13817 -1006 -13783
rect -1040 -13885 -1006 -13851
rect -22 -13409 12 -13375
rect -22 -13477 12 -13443
rect -22 -13545 12 -13511
rect 2582 -13371 2616 -13337
rect 2582 -13439 2616 -13405
rect 2582 -13507 2616 -13473
rect 3600 -13031 3634 -12997
rect 3600 -13099 3634 -13065
rect 3600 -13167 3634 -13133
rect 3600 -13235 3634 -13201
rect 3600 -13303 3634 -13269
rect 3600 -13371 3634 -13337
rect 3600 -13439 3634 -13405
rect 3600 -13507 3634 -13473
rect 4618 -13031 4652 -12997
rect 4618 -13099 4652 -13065
rect 4618 -13167 4652 -13133
rect 4618 -13235 4652 -13201
rect 4618 -13303 4652 -13269
rect 4618 -13371 4652 -13337
rect 4618 -13439 4652 -13405
rect 4618 -13507 4652 -13473
rect 5636 -13031 5670 -12997
rect 5636 -13099 5670 -13065
rect 5636 -13167 5670 -13133
rect 5636 -13235 5670 -13201
rect 5636 -13303 5670 -13269
rect 5636 -13371 5670 -13337
rect 5636 -13439 5670 -13405
rect 5636 -13507 5670 -13473
rect 6654 -13031 6688 -12997
rect 6654 -13099 6688 -13065
rect 6654 -13167 6688 -13133
rect 6654 -13235 6688 -13201
rect 6654 -13303 6688 -13269
rect 6654 -13371 6688 -13337
rect 6654 -13439 6688 -13405
rect 6654 -13507 6688 -13473
rect 7672 -13031 7706 -12997
rect 7672 -13099 7706 -13065
rect 7672 -13167 7706 -13133
rect 7672 -13235 7706 -13201
rect 7672 -13303 7706 -13269
rect 7672 -13371 7706 -13337
rect 7672 -13439 7706 -13405
rect 7672 -13507 7706 -13473
rect 8690 -13031 8724 -12997
rect 8690 -13099 8724 -13065
rect 8690 -13167 8724 -13133
rect 8690 -13235 8724 -13201
rect 8690 -13303 8724 -13269
rect 8690 -13371 8724 -13337
rect 8690 -13439 8724 -13405
rect 8690 -13507 8724 -13473
rect 9708 -13031 9742 -12997
rect 9708 -13099 9742 -13065
rect 9708 -13167 9742 -13133
rect 9708 -13235 9742 -13201
rect 9708 -13303 9742 -13269
rect 9708 -13371 9742 -13337
rect 9708 -13439 9742 -13405
rect 9708 -13507 9742 -13473
rect 10726 -13031 10760 -12997
rect 10726 -13099 10760 -13065
rect 10726 -13167 10760 -13133
rect 10726 -13235 10760 -13201
rect 10726 -13303 10760 -13269
rect 10726 -13371 10760 -13337
rect 10726 -13439 10760 -13405
rect 10726 -13507 10760 -13473
rect 11744 -13031 11778 -12997
rect 11744 -13099 11778 -13065
rect 11744 -13167 11778 -13133
rect 11744 -13235 11778 -13201
rect 11744 -13303 11778 -13269
rect 11744 -13371 11778 -13337
rect 11744 -13439 11778 -13405
rect 11744 -13507 11778 -13473
rect 12762 -13031 12796 -12997
rect 12762 -13099 12796 -13065
rect 12762 -13167 12796 -13133
rect 12762 -13235 12796 -13201
rect 12762 -13303 12796 -13269
rect 12762 -13371 12796 -13337
rect 12762 -13439 12796 -13405
rect 12762 -13507 12796 -13473
rect 13780 -13031 13814 -12997
rect 13780 -13099 13814 -13065
rect 13780 -13167 13814 -13133
rect 13780 -13235 13814 -13201
rect 13780 -13303 13814 -13269
rect 13780 -13371 13814 -13337
rect 13780 -13439 13814 -13405
rect 13780 -13507 13814 -13473
rect 14798 -13031 14832 -12997
rect 14798 -13099 14832 -13065
rect 14798 -13167 14832 -13133
rect 14798 -13235 14832 -13201
rect 14798 -13303 14832 -13269
rect 14798 -13371 14832 -13337
rect 14798 -13439 14832 -13405
rect 14798 -13507 14832 -13473
rect 15816 -13031 15850 -12997
rect 15816 -13099 15850 -13065
rect 15816 -13167 15850 -13133
rect 15816 -13235 15850 -13201
rect 15816 -13303 15850 -13269
rect 15816 -13371 15850 -13337
rect 15816 -13439 15850 -13405
rect 15816 -13507 15850 -13473
rect 16834 -13031 16868 -12997
rect 16834 -13099 16868 -13065
rect 16834 -13167 16868 -13133
rect 16834 -13235 16868 -13201
rect 16834 -13303 16868 -13269
rect 16834 -13371 16868 -13337
rect 16834 -13439 16868 -13405
rect 16834 -13507 16868 -13473
rect 17852 -13031 17886 -12997
rect 17852 -13099 17886 -13065
rect 17852 -13167 17886 -13133
rect 17852 -13235 17886 -13201
rect 17852 -13303 17886 -13269
rect 17852 -13371 17886 -13337
rect 17852 -13439 17886 -13405
rect 17852 -13507 17886 -13473
rect 18870 -13031 18904 -12997
rect 18870 -13099 18904 -13065
rect 18870 -13167 18904 -13133
rect 18870 -13235 18904 -13201
rect 18870 -13303 18904 -13269
rect 18870 -13371 18904 -13337
rect 18870 -13439 18904 -13405
rect 18870 -13507 18904 -13473
rect 19888 -13031 19922 -12997
rect 19888 -13099 19922 -13065
rect 19888 -13167 19922 -13133
rect 19888 -13235 19922 -13201
rect 19888 -13303 19922 -13269
rect 19888 -13371 19922 -13337
rect 19888 -13439 19922 -13405
rect 19888 -13507 19922 -13473
rect 20906 -13031 20940 -12997
rect 20906 -13099 20940 -13065
rect 20906 -13167 20940 -13133
rect 20906 -13235 20940 -13201
rect 20906 -13303 20940 -13269
rect 20906 -13371 20940 -13337
rect 20906 -13439 20940 -13405
rect 20906 -13507 20940 -13473
rect 21924 -13031 21958 -12997
rect 21924 -13099 21958 -13065
rect 21924 -13167 21958 -13133
rect 21924 -13235 21958 -13201
rect 21924 -13303 21958 -13269
rect 21924 -13371 21958 -13337
rect 21924 -13439 21958 -13405
rect 21924 -13507 21958 -13473
rect 22942 -13031 22976 -12997
rect 22942 -13099 22976 -13065
rect 22942 -13167 22976 -13133
rect 22942 -13235 22976 -13201
rect 22942 -13303 22976 -13269
rect 22942 -13371 22976 -13337
rect 22942 -13439 22976 -13405
rect 22942 -13507 22976 -13473
rect -22 -13613 12 -13579
rect -22 -13681 12 -13647
rect -22 -13749 12 -13715
rect -22 -13817 12 -13783
rect -22 -13885 12 -13851
rect -9184 -14227 -9150 -14193
rect -9184 -14295 -9150 -14261
rect -9184 -14363 -9150 -14329
rect -9184 -14431 -9150 -14397
rect -9184 -14499 -9150 -14465
rect -9184 -14567 -9150 -14533
rect -9184 -14635 -9150 -14601
rect -9184 -14703 -9150 -14669
rect -8166 -14227 -8132 -14193
rect -8166 -14295 -8132 -14261
rect -8166 -14363 -8132 -14329
rect -8166 -14431 -8132 -14397
rect -8166 -14499 -8132 -14465
rect -8166 -14567 -8132 -14533
rect -8166 -14635 -8132 -14601
rect -8166 -14703 -8132 -14669
rect -7148 -14227 -7114 -14193
rect -7148 -14295 -7114 -14261
rect -7148 -14363 -7114 -14329
rect -7148 -14431 -7114 -14397
rect -7148 -14499 -7114 -14465
rect -7148 -14567 -7114 -14533
rect -7148 -14635 -7114 -14601
rect -7148 -14703 -7114 -14669
rect -6130 -14227 -6096 -14193
rect -6130 -14295 -6096 -14261
rect -6130 -14363 -6096 -14329
rect -6130 -14431 -6096 -14397
rect -6130 -14499 -6096 -14465
rect -6130 -14567 -6096 -14533
rect -6130 -14635 -6096 -14601
rect -6130 -14703 -6096 -14669
rect -5112 -14227 -5078 -14193
rect -5112 -14295 -5078 -14261
rect -5112 -14363 -5078 -14329
rect -5112 -14431 -5078 -14397
rect -5112 -14499 -5078 -14465
rect -5112 -14567 -5078 -14533
rect -5112 -14635 -5078 -14601
rect -5112 -14703 -5078 -14669
rect -4094 -14227 -4060 -14193
rect -4094 -14295 -4060 -14261
rect -4094 -14363 -4060 -14329
rect -4094 -14431 -4060 -14397
rect -4094 -14499 -4060 -14465
rect -4094 -14567 -4060 -14533
rect -4094 -14635 -4060 -14601
rect -4094 -14703 -4060 -14669
rect -3076 -14227 -3042 -14193
rect -3076 -14295 -3042 -14261
rect -3076 -14363 -3042 -14329
rect -3076 -14431 -3042 -14397
rect -3076 -14499 -3042 -14465
rect -3076 -14567 -3042 -14533
rect -3076 -14635 -3042 -14601
rect -3076 -14703 -3042 -14669
rect -2058 -14227 -2024 -14193
rect -2058 -14295 -2024 -14261
rect -2058 -14363 -2024 -14329
rect -2058 -14431 -2024 -14397
rect -2058 -14499 -2024 -14465
rect -2058 -14567 -2024 -14533
rect -2058 -14635 -2024 -14601
rect -2058 -14703 -2024 -14669
rect -1040 -14227 -1006 -14193
rect -1040 -14295 -1006 -14261
rect -1040 -14363 -1006 -14329
rect -1040 -14431 -1006 -14397
rect -1040 -14499 -1006 -14465
rect -1040 -14567 -1006 -14533
rect -1040 -14635 -1006 -14601
rect -1040 -14703 -1006 -14669
rect -22 -14227 12 -14193
rect -22 -14295 12 -14261
rect -22 -14363 12 -14329
rect -22 -14431 12 -14397
rect -22 -14499 12 -14465
rect -22 -14567 12 -14533
rect -22 -14635 12 -14601
rect -22 -14703 12 -14669
rect 2582 -14263 2616 -14229
rect 2582 -14331 2616 -14297
rect 2582 -14399 2616 -14365
rect 2582 -14467 2616 -14433
rect 2582 -14535 2616 -14501
rect 2582 -14603 2616 -14569
rect 2582 -14671 2616 -14637
rect 2582 -14739 2616 -14705
rect 3600 -14263 3634 -14229
rect 3600 -14331 3634 -14297
rect 3600 -14399 3634 -14365
rect 3600 -14467 3634 -14433
rect 3600 -14535 3634 -14501
rect 3600 -14603 3634 -14569
rect 3600 -14671 3634 -14637
rect 3600 -14739 3634 -14705
rect 4618 -14263 4652 -14229
rect 4618 -14331 4652 -14297
rect 4618 -14399 4652 -14365
rect 4618 -14467 4652 -14433
rect 4618 -14535 4652 -14501
rect 4618 -14603 4652 -14569
rect 4618 -14671 4652 -14637
rect 4618 -14739 4652 -14705
rect 5636 -14263 5670 -14229
rect 5636 -14331 5670 -14297
rect 5636 -14399 5670 -14365
rect 5636 -14467 5670 -14433
rect 5636 -14535 5670 -14501
rect 5636 -14603 5670 -14569
rect 5636 -14671 5670 -14637
rect 5636 -14739 5670 -14705
rect 6654 -14263 6688 -14229
rect 6654 -14331 6688 -14297
rect 6654 -14399 6688 -14365
rect 6654 -14467 6688 -14433
rect 6654 -14535 6688 -14501
rect 6654 -14603 6688 -14569
rect 6654 -14671 6688 -14637
rect 6654 -14739 6688 -14705
rect 7672 -14263 7706 -14229
rect 7672 -14331 7706 -14297
rect 7672 -14399 7706 -14365
rect 7672 -14467 7706 -14433
rect 7672 -14535 7706 -14501
rect 7672 -14603 7706 -14569
rect 7672 -14671 7706 -14637
rect 7672 -14739 7706 -14705
rect 8690 -14263 8724 -14229
rect 8690 -14331 8724 -14297
rect 8690 -14399 8724 -14365
rect 8690 -14467 8724 -14433
rect 8690 -14535 8724 -14501
rect 8690 -14603 8724 -14569
rect 8690 -14671 8724 -14637
rect 8690 -14739 8724 -14705
rect 9708 -14263 9742 -14229
rect 9708 -14331 9742 -14297
rect 9708 -14399 9742 -14365
rect 9708 -14467 9742 -14433
rect 9708 -14535 9742 -14501
rect 9708 -14603 9742 -14569
rect 9708 -14671 9742 -14637
rect 9708 -14739 9742 -14705
rect 10726 -14263 10760 -14229
rect 10726 -14331 10760 -14297
rect 10726 -14399 10760 -14365
rect 10726 -14467 10760 -14433
rect 10726 -14535 10760 -14501
rect 10726 -14603 10760 -14569
rect 10726 -14671 10760 -14637
rect 10726 -14739 10760 -14705
rect 11744 -14263 11778 -14229
rect 11744 -14331 11778 -14297
rect 11744 -14399 11778 -14365
rect 11744 -14467 11778 -14433
rect 11744 -14535 11778 -14501
rect 11744 -14603 11778 -14569
rect 11744 -14671 11778 -14637
rect 11744 -14739 11778 -14705
rect 12762 -14263 12796 -14229
rect 12762 -14331 12796 -14297
rect 12762 -14399 12796 -14365
rect 12762 -14467 12796 -14433
rect 12762 -14535 12796 -14501
rect 12762 -14603 12796 -14569
rect 12762 -14671 12796 -14637
rect 12762 -14739 12796 -14705
rect 13780 -14263 13814 -14229
rect 13780 -14331 13814 -14297
rect 13780 -14399 13814 -14365
rect 13780 -14467 13814 -14433
rect 13780 -14535 13814 -14501
rect 13780 -14603 13814 -14569
rect 13780 -14671 13814 -14637
rect 13780 -14739 13814 -14705
rect 14798 -14263 14832 -14229
rect 14798 -14331 14832 -14297
rect 14798 -14399 14832 -14365
rect 14798 -14467 14832 -14433
rect 14798 -14535 14832 -14501
rect 14798 -14603 14832 -14569
rect 14798 -14671 14832 -14637
rect 14798 -14739 14832 -14705
rect 15816 -14263 15850 -14229
rect 15816 -14331 15850 -14297
rect 15816 -14399 15850 -14365
rect 15816 -14467 15850 -14433
rect 15816 -14535 15850 -14501
rect 15816 -14603 15850 -14569
rect 15816 -14671 15850 -14637
rect 15816 -14739 15850 -14705
rect 16834 -14263 16868 -14229
rect 16834 -14331 16868 -14297
rect 16834 -14399 16868 -14365
rect 16834 -14467 16868 -14433
rect 16834 -14535 16868 -14501
rect 16834 -14603 16868 -14569
rect 16834 -14671 16868 -14637
rect 16834 -14739 16868 -14705
rect 17852 -14263 17886 -14229
rect 17852 -14331 17886 -14297
rect 17852 -14399 17886 -14365
rect 17852 -14467 17886 -14433
rect 17852 -14535 17886 -14501
rect 17852 -14603 17886 -14569
rect 17852 -14671 17886 -14637
rect 17852 -14739 17886 -14705
rect 18870 -14263 18904 -14229
rect 18870 -14331 18904 -14297
rect 18870 -14399 18904 -14365
rect 18870 -14467 18904 -14433
rect 18870 -14535 18904 -14501
rect 18870 -14603 18904 -14569
rect 18870 -14671 18904 -14637
rect 18870 -14739 18904 -14705
rect 19888 -14263 19922 -14229
rect 19888 -14331 19922 -14297
rect 19888 -14399 19922 -14365
rect 19888 -14467 19922 -14433
rect 19888 -14535 19922 -14501
rect 19888 -14603 19922 -14569
rect 19888 -14671 19922 -14637
rect 19888 -14739 19922 -14705
rect 20906 -14263 20940 -14229
rect 20906 -14331 20940 -14297
rect 20906 -14399 20940 -14365
rect 20906 -14467 20940 -14433
rect 20906 -14535 20940 -14501
rect 20906 -14603 20940 -14569
rect 20906 -14671 20940 -14637
rect 20906 -14739 20940 -14705
rect 21924 -14263 21958 -14229
rect 21924 -14331 21958 -14297
rect 21924 -14399 21958 -14365
rect 21924 -14467 21958 -14433
rect 21924 -14535 21958 -14501
rect 21924 -14603 21958 -14569
rect 21924 -14671 21958 -14637
rect 21924 -14739 21958 -14705
rect 22942 -14263 22976 -14229
rect 22942 -14331 22976 -14297
rect 22942 -14399 22976 -14365
rect 22942 -14467 22976 -14433
rect 22942 -14535 22976 -14501
rect 22942 -14603 22976 -14569
rect 22942 -14671 22976 -14637
rect 22942 -14739 22976 -14705
rect -9184 -15045 -9150 -15011
rect -9184 -15113 -9150 -15079
rect -9184 -15181 -9150 -15147
rect -9184 -15249 -9150 -15215
rect -9184 -15317 -9150 -15283
rect -9184 -15385 -9150 -15351
rect -9184 -15453 -9150 -15419
rect -9184 -15521 -9150 -15487
rect -8166 -15045 -8132 -15011
rect -8166 -15113 -8132 -15079
rect -8166 -15181 -8132 -15147
rect -8166 -15249 -8132 -15215
rect -8166 -15317 -8132 -15283
rect -8166 -15385 -8132 -15351
rect -8166 -15453 -8132 -15419
rect -8166 -15521 -8132 -15487
rect -7148 -15045 -7114 -15011
rect -7148 -15113 -7114 -15079
rect -7148 -15181 -7114 -15147
rect -7148 -15249 -7114 -15215
rect -7148 -15317 -7114 -15283
rect -7148 -15385 -7114 -15351
rect -7148 -15453 -7114 -15419
rect -7148 -15521 -7114 -15487
rect -6130 -15045 -6096 -15011
rect -6130 -15113 -6096 -15079
rect -6130 -15181 -6096 -15147
rect -6130 -15249 -6096 -15215
rect -6130 -15317 -6096 -15283
rect -6130 -15385 -6096 -15351
rect -6130 -15453 -6096 -15419
rect -6130 -15521 -6096 -15487
rect -5112 -15045 -5078 -15011
rect -5112 -15113 -5078 -15079
rect -5112 -15181 -5078 -15147
rect -5112 -15249 -5078 -15215
rect -5112 -15317 -5078 -15283
rect -5112 -15385 -5078 -15351
rect -5112 -15453 -5078 -15419
rect -5112 -15521 -5078 -15487
rect -4094 -15045 -4060 -15011
rect -4094 -15113 -4060 -15079
rect -4094 -15181 -4060 -15147
rect -4094 -15249 -4060 -15215
rect -4094 -15317 -4060 -15283
rect -4094 -15385 -4060 -15351
rect -4094 -15453 -4060 -15419
rect -4094 -15521 -4060 -15487
rect -3076 -15045 -3042 -15011
rect -3076 -15113 -3042 -15079
rect -3076 -15181 -3042 -15147
rect -3076 -15249 -3042 -15215
rect -3076 -15317 -3042 -15283
rect -3076 -15385 -3042 -15351
rect -3076 -15453 -3042 -15419
rect -3076 -15521 -3042 -15487
rect -2058 -15045 -2024 -15011
rect -2058 -15113 -2024 -15079
rect -2058 -15181 -2024 -15147
rect -2058 -15249 -2024 -15215
rect -2058 -15317 -2024 -15283
rect -2058 -15385 -2024 -15351
rect -2058 -15453 -2024 -15419
rect -2058 -15521 -2024 -15487
rect -1040 -15045 -1006 -15011
rect -1040 -15113 -1006 -15079
rect -1040 -15181 -1006 -15147
rect -1040 -15249 -1006 -15215
rect -1040 -15317 -1006 -15283
rect -1040 -15385 -1006 -15351
rect -1040 -15453 -1006 -15419
rect -1040 -15521 -1006 -15487
rect -22 -15045 12 -15011
rect -22 -15113 12 -15079
rect -22 -15181 12 -15147
rect -22 -15249 12 -15215
rect -22 -15317 12 -15283
rect -22 -15385 12 -15351
rect -22 -15453 12 -15419
rect -22 -15521 12 -15487
rect 2580 -15497 2614 -15463
rect 2580 -15565 2614 -15531
rect 2580 -15633 2614 -15599
rect 2580 -15701 2614 -15667
rect 2580 -15769 2614 -15735
rect -9184 -15863 -9150 -15829
rect -9184 -15931 -9150 -15897
rect -9184 -15999 -9150 -15965
rect -9184 -16067 -9150 -16033
rect -9184 -16135 -9150 -16101
rect -9184 -16203 -9150 -16169
rect -9184 -16271 -9150 -16237
rect -9184 -16339 -9150 -16305
rect -8166 -15863 -8132 -15829
rect -8166 -15931 -8132 -15897
rect -8166 -15999 -8132 -15965
rect -8166 -16067 -8132 -16033
rect -8166 -16135 -8132 -16101
rect -8166 -16203 -8132 -16169
rect -8166 -16271 -8132 -16237
rect -8166 -16339 -8132 -16305
rect -7148 -15863 -7114 -15829
rect -7148 -15931 -7114 -15897
rect -7148 -15999 -7114 -15965
rect -7148 -16067 -7114 -16033
rect -7148 -16135 -7114 -16101
rect -7148 -16203 -7114 -16169
rect -7148 -16271 -7114 -16237
rect -7148 -16339 -7114 -16305
rect -6130 -15863 -6096 -15829
rect -6130 -15931 -6096 -15897
rect -6130 -15999 -6096 -15965
rect -6130 -16067 -6096 -16033
rect -6130 -16135 -6096 -16101
rect -6130 -16203 -6096 -16169
rect -6130 -16271 -6096 -16237
rect -6130 -16339 -6096 -16305
rect -5112 -15863 -5078 -15829
rect -5112 -15931 -5078 -15897
rect -5112 -15999 -5078 -15965
rect -5112 -16067 -5078 -16033
rect -5112 -16135 -5078 -16101
rect -5112 -16203 -5078 -16169
rect -5112 -16271 -5078 -16237
rect -5112 -16339 -5078 -16305
rect -4094 -15863 -4060 -15829
rect -4094 -15931 -4060 -15897
rect -4094 -15999 -4060 -15965
rect -4094 -16067 -4060 -16033
rect -4094 -16135 -4060 -16101
rect -4094 -16203 -4060 -16169
rect -4094 -16271 -4060 -16237
rect -4094 -16339 -4060 -16305
rect -3076 -15863 -3042 -15829
rect -3076 -15931 -3042 -15897
rect -3076 -15999 -3042 -15965
rect -3076 -16067 -3042 -16033
rect -3076 -16135 -3042 -16101
rect -3076 -16203 -3042 -16169
rect -3076 -16271 -3042 -16237
rect -3076 -16339 -3042 -16305
rect -2058 -15863 -2024 -15829
rect -2058 -15931 -2024 -15897
rect -2058 -15999 -2024 -15965
rect -2058 -16067 -2024 -16033
rect -2058 -16135 -2024 -16101
rect -2058 -16203 -2024 -16169
rect -2058 -16271 -2024 -16237
rect -2058 -16339 -2024 -16305
rect -1040 -15863 -1006 -15829
rect -1040 -15931 -1006 -15897
rect -1040 -15999 -1006 -15965
rect -1040 -16067 -1006 -16033
rect -1040 -16135 -1006 -16101
rect -1040 -16203 -1006 -16169
rect -1040 -16271 -1006 -16237
rect -1040 -16339 -1006 -16305
rect -22 -15863 12 -15829
rect -22 -15931 12 -15897
rect -22 -15999 12 -15965
rect 2580 -15837 2614 -15803
rect 2580 -15905 2614 -15871
rect 2580 -15973 2614 -15939
rect 3598 -15497 3632 -15463
rect 3598 -15565 3632 -15531
rect 3598 -15633 3632 -15599
rect 3598 -15701 3632 -15667
rect 3598 -15769 3632 -15735
rect 3598 -15837 3632 -15803
rect 3598 -15905 3632 -15871
rect 3598 -15973 3632 -15939
rect 4616 -15497 4650 -15463
rect 4616 -15565 4650 -15531
rect 4616 -15633 4650 -15599
rect 4616 -15701 4650 -15667
rect 4616 -15769 4650 -15735
rect 4616 -15837 4650 -15803
rect 4616 -15905 4650 -15871
rect 4616 -15973 4650 -15939
rect 5634 -15497 5668 -15463
rect 5634 -15565 5668 -15531
rect 5634 -15633 5668 -15599
rect 5634 -15701 5668 -15667
rect 5634 -15769 5668 -15735
rect 5634 -15837 5668 -15803
rect 5634 -15905 5668 -15871
rect 5634 -15973 5668 -15939
rect 6652 -15497 6686 -15463
rect 6652 -15565 6686 -15531
rect 6652 -15633 6686 -15599
rect 6652 -15701 6686 -15667
rect 6652 -15769 6686 -15735
rect 6652 -15837 6686 -15803
rect 6652 -15905 6686 -15871
rect 6652 -15973 6686 -15939
rect 7670 -15497 7704 -15463
rect 7670 -15565 7704 -15531
rect 7670 -15633 7704 -15599
rect 7670 -15701 7704 -15667
rect 7670 -15769 7704 -15735
rect 7670 -15837 7704 -15803
rect 7670 -15905 7704 -15871
rect 7670 -15973 7704 -15939
rect 8688 -15497 8722 -15463
rect 8688 -15565 8722 -15531
rect 8688 -15633 8722 -15599
rect 8688 -15701 8722 -15667
rect 8688 -15769 8722 -15735
rect 8688 -15837 8722 -15803
rect 8688 -15905 8722 -15871
rect 8688 -15973 8722 -15939
rect 9706 -15497 9740 -15463
rect 9706 -15565 9740 -15531
rect 9706 -15633 9740 -15599
rect 9706 -15701 9740 -15667
rect 9706 -15769 9740 -15735
rect 9706 -15837 9740 -15803
rect 9706 -15905 9740 -15871
rect 9706 -15973 9740 -15939
rect 10724 -15497 10758 -15463
rect 10724 -15565 10758 -15531
rect 10724 -15633 10758 -15599
rect 10724 -15701 10758 -15667
rect 10724 -15769 10758 -15735
rect 10724 -15837 10758 -15803
rect 10724 -15905 10758 -15871
rect 10724 -15973 10758 -15939
rect 11742 -15497 11776 -15463
rect 11742 -15565 11776 -15531
rect 11742 -15633 11776 -15599
rect 11742 -15701 11776 -15667
rect 11742 -15769 11776 -15735
rect 11742 -15837 11776 -15803
rect 11742 -15905 11776 -15871
rect 11742 -15973 11776 -15939
rect 12760 -15497 12794 -15463
rect 12760 -15565 12794 -15531
rect 12760 -15633 12794 -15599
rect 12760 -15701 12794 -15667
rect 12760 -15769 12794 -15735
rect 12760 -15837 12794 -15803
rect 12760 -15905 12794 -15871
rect 12760 -15973 12794 -15939
rect 13778 -15497 13812 -15463
rect 13778 -15565 13812 -15531
rect 13778 -15633 13812 -15599
rect 13778 -15701 13812 -15667
rect 13778 -15769 13812 -15735
rect 13778 -15837 13812 -15803
rect 13778 -15905 13812 -15871
rect 13778 -15973 13812 -15939
rect 14796 -15497 14830 -15463
rect 14796 -15565 14830 -15531
rect 14796 -15633 14830 -15599
rect 14796 -15701 14830 -15667
rect 14796 -15769 14830 -15735
rect 14796 -15837 14830 -15803
rect 14796 -15905 14830 -15871
rect 14796 -15973 14830 -15939
rect 15814 -15497 15848 -15463
rect 15814 -15565 15848 -15531
rect 15814 -15633 15848 -15599
rect 15814 -15701 15848 -15667
rect 15814 -15769 15848 -15735
rect 15814 -15837 15848 -15803
rect 15814 -15905 15848 -15871
rect 15814 -15973 15848 -15939
rect 16832 -15497 16866 -15463
rect 16832 -15565 16866 -15531
rect 16832 -15633 16866 -15599
rect 16832 -15701 16866 -15667
rect 16832 -15769 16866 -15735
rect 16832 -15837 16866 -15803
rect 16832 -15905 16866 -15871
rect 16832 -15973 16866 -15939
rect 17850 -15497 17884 -15463
rect 17850 -15565 17884 -15531
rect 17850 -15633 17884 -15599
rect 17850 -15701 17884 -15667
rect 17850 -15769 17884 -15735
rect 17850 -15837 17884 -15803
rect 17850 -15905 17884 -15871
rect 17850 -15973 17884 -15939
rect 18868 -15497 18902 -15463
rect 18868 -15565 18902 -15531
rect 18868 -15633 18902 -15599
rect 18868 -15701 18902 -15667
rect 18868 -15769 18902 -15735
rect 18868 -15837 18902 -15803
rect 18868 -15905 18902 -15871
rect 18868 -15973 18902 -15939
rect 19886 -15497 19920 -15463
rect 19886 -15565 19920 -15531
rect 19886 -15633 19920 -15599
rect 19886 -15701 19920 -15667
rect 19886 -15769 19920 -15735
rect 19886 -15837 19920 -15803
rect 19886 -15905 19920 -15871
rect 19886 -15973 19920 -15939
rect 20904 -15497 20938 -15463
rect 20904 -15565 20938 -15531
rect 20904 -15633 20938 -15599
rect 20904 -15701 20938 -15667
rect 20904 -15769 20938 -15735
rect 20904 -15837 20938 -15803
rect 20904 -15905 20938 -15871
rect 20904 -15973 20938 -15939
rect 21922 -15497 21956 -15463
rect 21922 -15565 21956 -15531
rect 21922 -15633 21956 -15599
rect 21922 -15701 21956 -15667
rect 21922 -15769 21956 -15735
rect 21922 -15837 21956 -15803
rect 21922 -15905 21956 -15871
rect 21922 -15973 21956 -15939
rect 22940 -15497 22974 -15463
rect 22940 -15565 22974 -15531
rect 22940 -15633 22974 -15599
rect 22940 -15701 22974 -15667
rect 22940 -15769 22974 -15735
rect 22940 -15837 22974 -15803
rect 22940 -15905 22974 -15871
rect 22940 -15973 22974 -15939
rect -22 -16067 12 -16033
rect -22 -16135 12 -16101
rect -22 -16203 12 -16169
rect -22 -16271 12 -16237
rect -22 -16339 12 -16305
rect -9184 -16681 -9150 -16647
rect -9184 -16749 -9150 -16715
rect -9184 -16817 -9150 -16783
rect -9184 -16885 -9150 -16851
rect -9184 -16953 -9150 -16919
rect -9184 -17021 -9150 -16987
rect -9184 -17089 -9150 -17055
rect -9184 -17157 -9150 -17123
rect -8166 -16681 -8132 -16647
rect -8166 -16749 -8132 -16715
rect -8166 -16817 -8132 -16783
rect -8166 -16885 -8132 -16851
rect -8166 -16953 -8132 -16919
rect -8166 -17021 -8132 -16987
rect -8166 -17089 -8132 -17055
rect -8166 -17157 -8132 -17123
rect -7148 -16681 -7114 -16647
rect -7148 -16749 -7114 -16715
rect -7148 -16817 -7114 -16783
rect -7148 -16885 -7114 -16851
rect -7148 -16953 -7114 -16919
rect -7148 -17021 -7114 -16987
rect -7148 -17089 -7114 -17055
rect -7148 -17157 -7114 -17123
rect -6130 -16681 -6096 -16647
rect -6130 -16749 -6096 -16715
rect -6130 -16817 -6096 -16783
rect -6130 -16885 -6096 -16851
rect -6130 -16953 -6096 -16919
rect -6130 -17021 -6096 -16987
rect -6130 -17089 -6096 -17055
rect -6130 -17157 -6096 -17123
rect -5112 -16681 -5078 -16647
rect -5112 -16749 -5078 -16715
rect -5112 -16817 -5078 -16783
rect -5112 -16885 -5078 -16851
rect -5112 -16953 -5078 -16919
rect -5112 -17021 -5078 -16987
rect -5112 -17089 -5078 -17055
rect -5112 -17157 -5078 -17123
rect -4094 -16681 -4060 -16647
rect -4094 -16749 -4060 -16715
rect -4094 -16817 -4060 -16783
rect -4094 -16885 -4060 -16851
rect -4094 -16953 -4060 -16919
rect -4094 -17021 -4060 -16987
rect -4094 -17089 -4060 -17055
rect -4094 -17157 -4060 -17123
rect -3076 -16681 -3042 -16647
rect -3076 -16749 -3042 -16715
rect -3076 -16817 -3042 -16783
rect -3076 -16885 -3042 -16851
rect -3076 -16953 -3042 -16919
rect -3076 -17021 -3042 -16987
rect -3076 -17089 -3042 -17055
rect -3076 -17157 -3042 -17123
rect -2058 -16681 -2024 -16647
rect -2058 -16749 -2024 -16715
rect -2058 -16817 -2024 -16783
rect -2058 -16885 -2024 -16851
rect -2058 -16953 -2024 -16919
rect -2058 -17021 -2024 -16987
rect -2058 -17089 -2024 -17055
rect -2058 -17157 -2024 -17123
rect -1040 -16681 -1006 -16647
rect -1040 -16749 -1006 -16715
rect -1040 -16817 -1006 -16783
rect -1040 -16885 -1006 -16851
rect -1040 -16953 -1006 -16919
rect -1040 -17021 -1006 -16987
rect -1040 -17089 -1006 -17055
rect -1040 -17157 -1006 -17123
rect -22 -16681 12 -16647
rect -22 -16749 12 -16715
rect -22 -16817 12 -16783
rect -22 -16885 12 -16851
rect -22 -16953 12 -16919
rect -22 -17021 12 -16987
rect -22 -17089 12 -17055
rect -22 -17157 12 -17123
rect 2580 -16731 2614 -16697
rect 2580 -16799 2614 -16765
rect 2580 -16867 2614 -16833
rect 2580 -16935 2614 -16901
rect 2580 -17003 2614 -16969
rect 2580 -17071 2614 -17037
rect 2580 -17139 2614 -17105
rect 2580 -17207 2614 -17173
rect 3598 -16731 3632 -16697
rect 3598 -16799 3632 -16765
rect 3598 -16867 3632 -16833
rect 3598 -16935 3632 -16901
rect 3598 -17003 3632 -16969
rect 3598 -17071 3632 -17037
rect 3598 -17139 3632 -17105
rect 3598 -17207 3632 -17173
rect 4616 -16731 4650 -16697
rect 4616 -16799 4650 -16765
rect 4616 -16867 4650 -16833
rect 4616 -16935 4650 -16901
rect 4616 -17003 4650 -16969
rect 4616 -17071 4650 -17037
rect 4616 -17139 4650 -17105
rect 4616 -17207 4650 -17173
rect 5634 -16731 5668 -16697
rect 5634 -16799 5668 -16765
rect 5634 -16867 5668 -16833
rect 5634 -16935 5668 -16901
rect 5634 -17003 5668 -16969
rect 5634 -17071 5668 -17037
rect 5634 -17139 5668 -17105
rect 5634 -17207 5668 -17173
rect 6652 -16731 6686 -16697
rect 6652 -16799 6686 -16765
rect 6652 -16867 6686 -16833
rect 6652 -16935 6686 -16901
rect 6652 -17003 6686 -16969
rect 6652 -17071 6686 -17037
rect 6652 -17139 6686 -17105
rect 6652 -17207 6686 -17173
rect 7670 -16731 7704 -16697
rect 7670 -16799 7704 -16765
rect 7670 -16867 7704 -16833
rect 7670 -16935 7704 -16901
rect 7670 -17003 7704 -16969
rect 7670 -17071 7704 -17037
rect 7670 -17139 7704 -17105
rect 7670 -17207 7704 -17173
rect 8688 -16731 8722 -16697
rect 8688 -16799 8722 -16765
rect 8688 -16867 8722 -16833
rect 8688 -16935 8722 -16901
rect 8688 -17003 8722 -16969
rect 8688 -17071 8722 -17037
rect 8688 -17139 8722 -17105
rect 8688 -17207 8722 -17173
rect 9706 -16731 9740 -16697
rect 9706 -16799 9740 -16765
rect 9706 -16867 9740 -16833
rect 9706 -16935 9740 -16901
rect 9706 -17003 9740 -16969
rect 9706 -17071 9740 -17037
rect 9706 -17139 9740 -17105
rect 9706 -17207 9740 -17173
rect 10724 -16731 10758 -16697
rect 10724 -16799 10758 -16765
rect 10724 -16867 10758 -16833
rect 10724 -16935 10758 -16901
rect 10724 -17003 10758 -16969
rect 10724 -17071 10758 -17037
rect 10724 -17139 10758 -17105
rect 10724 -17207 10758 -17173
rect 11742 -16731 11776 -16697
rect 11742 -16799 11776 -16765
rect 11742 -16867 11776 -16833
rect 11742 -16935 11776 -16901
rect 11742 -17003 11776 -16969
rect 11742 -17071 11776 -17037
rect 11742 -17139 11776 -17105
rect 11742 -17207 11776 -17173
rect 12760 -16731 12794 -16697
rect 12760 -16799 12794 -16765
rect 12760 -16867 12794 -16833
rect 12760 -16935 12794 -16901
rect 12760 -17003 12794 -16969
rect 12760 -17071 12794 -17037
rect 12760 -17139 12794 -17105
rect 12760 -17207 12794 -17173
rect 13778 -16731 13812 -16697
rect 13778 -16799 13812 -16765
rect 13778 -16867 13812 -16833
rect 13778 -16935 13812 -16901
rect 13778 -17003 13812 -16969
rect 13778 -17071 13812 -17037
rect 13778 -17139 13812 -17105
rect 13778 -17207 13812 -17173
rect 14796 -16731 14830 -16697
rect 14796 -16799 14830 -16765
rect 14796 -16867 14830 -16833
rect 14796 -16935 14830 -16901
rect 14796 -17003 14830 -16969
rect 14796 -17071 14830 -17037
rect 14796 -17139 14830 -17105
rect 14796 -17207 14830 -17173
rect 15814 -16731 15848 -16697
rect 15814 -16799 15848 -16765
rect 15814 -16867 15848 -16833
rect 15814 -16935 15848 -16901
rect 15814 -17003 15848 -16969
rect 15814 -17071 15848 -17037
rect 15814 -17139 15848 -17105
rect 15814 -17207 15848 -17173
rect 16832 -16731 16866 -16697
rect 16832 -16799 16866 -16765
rect 16832 -16867 16866 -16833
rect 16832 -16935 16866 -16901
rect 16832 -17003 16866 -16969
rect 16832 -17071 16866 -17037
rect 16832 -17139 16866 -17105
rect 16832 -17207 16866 -17173
rect 17850 -16731 17884 -16697
rect 17850 -16799 17884 -16765
rect 17850 -16867 17884 -16833
rect 17850 -16935 17884 -16901
rect 17850 -17003 17884 -16969
rect 17850 -17071 17884 -17037
rect 17850 -17139 17884 -17105
rect 17850 -17207 17884 -17173
rect 18868 -16731 18902 -16697
rect 18868 -16799 18902 -16765
rect 18868 -16867 18902 -16833
rect 18868 -16935 18902 -16901
rect 18868 -17003 18902 -16969
rect 18868 -17071 18902 -17037
rect 18868 -17139 18902 -17105
rect 18868 -17207 18902 -17173
rect 19886 -16731 19920 -16697
rect 19886 -16799 19920 -16765
rect 19886 -16867 19920 -16833
rect 19886 -16935 19920 -16901
rect 19886 -17003 19920 -16969
rect 19886 -17071 19920 -17037
rect 19886 -17139 19920 -17105
rect 19886 -17207 19920 -17173
rect 20904 -16731 20938 -16697
rect 20904 -16799 20938 -16765
rect 20904 -16867 20938 -16833
rect 20904 -16935 20938 -16901
rect 20904 -17003 20938 -16969
rect 20904 -17071 20938 -17037
rect 20904 -17139 20938 -17105
rect 20904 -17207 20938 -17173
rect 21922 -16731 21956 -16697
rect 21922 -16799 21956 -16765
rect 21922 -16867 21956 -16833
rect 21922 -16935 21956 -16901
rect 21922 -17003 21956 -16969
rect 21922 -17071 21956 -17037
rect 21922 -17139 21956 -17105
rect 21922 -17207 21956 -17173
rect 22940 -16731 22974 -16697
rect 22940 -16799 22974 -16765
rect 22940 -16867 22974 -16833
rect 22940 -16935 22974 -16901
rect 22940 -17003 22974 -16969
rect 22940 -17071 22974 -17037
rect 22940 -17139 22974 -17105
rect 22940 -17207 22974 -17173
rect -9184 -17499 -9150 -17465
rect -9184 -17567 -9150 -17533
rect -9184 -17635 -9150 -17601
rect -9184 -17703 -9150 -17669
rect -9184 -17771 -9150 -17737
rect -9184 -17839 -9150 -17805
rect -9184 -17907 -9150 -17873
rect -9184 -17975 -9150 -17941
rect -8166 -17499 -8132 -17465
rect -8166 -17567 -8132 -17533
rect -8166 -17635 -8132 -17601
rect -8166 -17703 -8132 -17669
rect -8166 -17771 -8132 -17737
rect -8166 -17839 -8132 -17805
rect -8166 -17907 -8132 -17873
rect -8166 -17975 -8132 -17941
rect -7148 -17499 -7114 -17465
rect -7148 -17567 -7114 -17533
rect -7148 -17635 -7114 -17601
rect -7148 -17703 -7114 -17669
rect -7148 -17771 -7114 -17737
rect -7148 -17839 -7114 -17805
rect -7148 -17907 -7114 -17873
rect -7148 -17975 -7114 -17941
rect -6130 -17499 -6096 -17465
rect -6130 -17567 -6096 -17533
rect -6130 -17635 -6096 -17601
rect -6130 -17703 -6096 -17669
rect -6130 -17771 -6096 -17737
rect -6130 -17839 -6096 -17805
rect -6130 -17907 -6096 -17873
rect -6130 -17975 -6096 -17941
rect -5112 -17499 -5078 -17465
rect -5112 -17567 -5078 -17533
rect -5112 -17635 -5078 -17601
rect -5112 -17703 -5078 -17669
rect -5112 -17771 -5078 -17737
rect -5112 -17839 -5078 -17805
rect -5112 -17907 -5078 -17873
rect -5112 -17975 -5078 -17941
rect -4094 -17499 -4060 -17465
rect -4094 -17567 -4060 -17533
rect -4094 -17635 -4060 -17601
rect -4094 -17703 -4060 -17669
rect -4094 -17771 -4060 -17737
rect -4094 -17839 -4060 -17805
rect -4094 -17907 -4060 -17873
rect -4094 -17975 -4060 -17941
rect -3076 -17499 -3042 -17465
rect -3076 -17567 -3042 -17533
rect -3076 -17635 -3042 -17601
rect -3076 -17703 -3042 -17669
rect -3076 -17771 -3042 -17737
rect -3076 -17839 -3042 -17805
rect -3076 -17907 -3042 -17873
rect -3076 -17975 -3042 -17941
rect -2058 -17499 -2024 -17465
rect -2058 -17567 -2024 -17533
rect -2058 -17635 -2024 -17601
rect -2058 -17703 -2024 -17669
rect -2058 -17771 -2024 -17737
rect -2058 -17839 -2024 -17805
rect -2058 -17907 -2024 -17873
rect -2058 -17975 -2024 -17941
rect -1040 -17499 -1006 -17465
rect -1040 -17567 -1006 -17533
rect -1040 -17635 -1006 -17601
rect -1040 -17703 -1006 -17669
rect -1040 -17771 -1006 -17737
rect -1040 -17839 -1006 -17805
rect -1040 -17907 -1006 -17873
rect -1040 -17975 -1006 -17941
rect -22 -17499 12 -17465
rect -22 -17567 12 -17533
rect -22 -17635 12 -17601
rect -22 -17703 12 -17669
rect -22 -17771 12 -17737
rect -22 -17839 12 -17805
rect -22 -17907 12 -17873
rect -22 -17975 12 -17941
rect 2580 -17963 2614 -17929
rect 2580 -18031 2614 -17997
rect 2580 -18099 2614 -18065
rect 2580 -18167 2614 -18133
rect 2580 -18235 2614 -18201
rect -9184 -18317 -9150 -18283
rect -9184 -18385 -9150 -18351
rect -9184 -18453 -9150 -18419
rect -9184 -18521 -9150 -18487
rect -9184 -18589 -9150 -18555
rect -9184 -18657 -9150 -18623
rect -9184 -18725 -9150 -18691
rect -9184 -18793 -9150 -18759
rect -8166 -18317 -8132 -18283
rect -8166 -18385 -8132 -18351
rect -8166 -18453 -8132 -18419
rect -8166 -18521 -8132 -18487
rect -8166 -18589 -8132 -18555
rect -8166 -18657 -8132 -18623
rect -8166 -18725 -8132 -18691
rect -8166 -18793 -8132 -18759
rect -7148 -18317 -7114 -18283
rect -7148 -18385 -7114 -18351
rect -7148 -18453 -7114 -18419
rect -7148 -18521 -7114 -18487
rect -7148 -18589 -7114 -18555
rect -7148 -18657 -7114 -18623
rect -7148 -18725 -7114 -18691
rect -7148 -18793 -7114 -18759
rect -6130 -18317 -6096 -18283
rect -6130 -18385 -6096 -18351
rect -6130 -18453 -6096 -18419
rect -6130 -18521 -6096 -18487
rect -6130 -18589 -6096 -18555
rect -6130 -18657 -6096 -18623
rect -6130 -18725 -6096 -18691
rect -6130 -18793 -6096 -18759
rect -5112 -18317 -5078 -18283
rect -5112 -18385 -5078 -18351
rect -5112 -18453 -5078 -18419
rect -5112 -18521 -5078 -18487
rect -5112 -18589 -5078 -18555
rect -5112 -18657 -5078 -18623
rect -5112 -18725 -5078 -18691
rect -5112 -18793 -5078 -18759
rect -4094 -18317 -4060 -18283
rect -4094 -18385 -4060 -18351
rect -4094 -18453 -4060 -18419
rect -4094 -18521 -4060 -18487
rect -4094 -18589 -4060 -18555
rect -4094 -18657 -4060 -18623
rect -4094 -18725 -4060 -18691
rect -4094 -18793 -4060 -18759
rect -3076 -18317 -3042 -18283
rect -3076 -18385 -3042 -18351
rect -3076 -18453 -3042 -18419
rect -3076 -18521 -3042 -18487
rect -3076 -18589 -3042 -18555
rect -3076 -18657 -3042 -18623
rect -3076 -18725 -3042 -18691
rect -3076 -18793 -3042 -18759
rect -2058 -18317 -2024 -18283
rect -2058 -18385 -2024 -18351
rect -2058 -18453 -2024 -18419
rect -2058 -18521 -2024 -18487
rect -2058 -18589 -2024 -18555
rect -2058 -18657 -2024 -18623
rect -2058 -18725 -2024 -18691
rect -2058 -18793 -2024 -18759
rect -1040 -18317 -1006 -18283
rect -1040 -18385 -1006 -18351
rect -1040 -18453 -1006 -18419
rect -1040 -18521 -1006 -18487
rect -1040 -18589 -1006 -18555
rect -1040 -18657 -1006 -18623
rect -1040 -18725 -1006 -18691
rect -1040 -18793 -1006 -18759
rect -22 -18317 12 -18283
rect -22 -18385 12 -18351
rect -22 -18453 12 -18419
rect 2580 -18303 2614 -18269
rect 2580 -18371 2614 -18337
rect 2580 -18439 2614 -18405
rect 3598 -17963 3632 -17929
rect 3598 -18031 3632 -17997
rect 3598 -18099 3632 -18065
rect 3598 -18167 3632 -18133
rect 3598 -18235 3632 -18201
rect 3598 -18303 3632 -18269
rect 3598 -18371 3632 -18337
rect 3598 -18439 3632 -18405
rect 4616 -17963 4650 -17929
rect 4616 -18031 4650 -17997
rect 4616 -18099 4650 -18065
rect 4616 -18167 4650 -18133
rect 4616 -18235 4650 -18201
rect 4616 -18303 4650 -18269
rect 4616 -18371 4650 -18337
rect 4616 -18439 4650 -18405
rect 5634 -17963 5668 -17929
rect 5634 -18031 5668 -17997
rect 5634 -18099 5668 -18065
rect 5634 -18167 5668 -18133
rect 5634 -18235 5668 -18201
rect 5634 -18303 5668 -18269
rect 5634 -18371 5668 -18337
rect 5634 -18439 5668 -18405
rect 6652 -17963 6686 -17929
rect 6652 -18031 6686 -17997
rect 6652 -18099 6686 -18065
rect 6652 -18167 6686 -18133
rect 6652 -18235 6686 -18201
rect 6652 -18303 6686 -18269
rect 6652 -18371 6686 -18337
rect 6652 -18439 6686 -18405
rect 7670 -17963 7704 -17929
rect 7670 -18031 7704 -17997
rect 7670 -18099 7704 -18065
rect 7670 -18167 7704 -18133
rect 7670 -18235 7704 -18201
rect 7670 -18303 7704 -18269
rect 7670 -18371 7704 -18337
rect 7670 -18439 7704 -18405
rect 8688 -17963 8722 -17929
rect 8688 -18031 8722 -17997
rect 8688 -18099 8722 -18065
rect 8688 -18167 8722 -18133
rect 8688 -18235 8722 -18201
rect 8688 -18303 8722 -18269
rect 8688 -18371 8722 -18337
rect 8688 -18439 8722 -18405
rect 9706 -17963 9740 -17929
rect 9706 -18031 9740 -17997
rect 9706 -18099 9740 -18065
rect 9706 -18167 9740 -18133
rect 9706 -18235 9740 -18201
rect 9706 -18303 9740 -18269
rect 9706 -18371 9740 -18337
rect 9706 -18439 9740 -18405
rect 10724 -17963 10758 -17929
rect 10724 -18031 10758 -17997
rect 10724 -18099 10758 -18065
rect 10724 -18167 10758 -18133
rect 10724 -18235 10758 -18201
rect 10724 -18303 10758 -18269
rect 10724 -18371 10758 -18337
rect 10724 -18439 10758 -18405
rect 11742 -17963 11776 -17929
rect 11742 -18031 11776 -17997
rect 11742 -18099 11776 -18065
rect 11742 -18167 11776 -18133
rect 11742 -18235 11776 -18201
rect 11742 -18303 11776 -18269
rect 11742 -18371 11776 -18337
rect 11742 -18439 11776 -18405
rect 12760 -17963 12794 -17929
rect 12760 -18031 12794 -17997
rect 12760 -18099 12794 -18065
rect 12760 -18167 12794 -18133
rect 12760 -18235 12794 -18201
rect 12760 -18303 12794 -18269
rect 12760 -18371 12794 -18337
rect 12760 -18439 12794 -18405
rect 13778 -17963 13812 -17929
rect 13778 -18031 13812 -17997
rect 13778 -18099 13812 -18065
rect 13778 -18167 13812 -18133
rect 13778 -18235 13812 -18201
rect 13778 -18303 13812 -18269
rect 13778 -18371 13812 -18337
rect 13778 -18439 13812 -18405
rect 14796 -17963 14830 -17929
rect 14796 -18031 14830 -17997
rect 14796 -18099 14830 -18065
rect 14796 -18167 14830 -18133
rect 14796 -18235 14830 -18201
rect 14796 -18303 14830 -18269
rect 14796 -18371 14830 -18337
rect 14796 -18439 14830 -18405
rect 15814 -17963 15848 -17929
rect 15814 -18031 15848 -17997
rect 15814 -18099 15848 -18065
rect 15814 -18167 15848 -18133
rect 15814 -18235 15848 -18201
rect 15814 -18303 15848 -18269
rect 15814 -18371 15848 -18337
rect 15814 -18439 15848 -18405
rect 16832 -17963 16866 -17929
rect 16832 -18031 16866 -17997
rect 16832 -18099 16866 -18065
rect 16832 -18167 16866 -18133
rect 16832 -18235 16866 -18201
rect 16832 -18303 16866 -18269
rect 16832 -18371 16866 -18337
rect 16832 -18439 16866 -18405
rect 17850 -17963 17884 -17929
rect 17850 -18031 17884 -17997
rect 17850 -18099 17884 -18065
rect 17850 -18167 17884 -18133
rect 17850 -18235 17884 -18201
rect 17850 -18303 17884 -18269
rect 17850 -18371 17884 -18337
rect 17850 -18439 17884 -18405
rect 18868 -17963 18902 -17929
rect 18868 -18031 18902 -17997
rect 18868 -18099 18902 -18065
rect 18868 -18167 18902 -18133
rect 18868 -18235 18902 -18201
rect 18868 -18303 18902 -18269
rect 18868 -18371 18902 -18337
rect 18868 -18439 18902 -18405
rect 19886 -17963 19920 -17929
rect 19886 -18031 19920 -17997
rect 19886 -18099 19920 -18065
rect 19886 -18167 19920 -18133
rect 19886 -18235 19920 -18201
rect 19886 -18303 19920 -18269
rect 19886 -18371 19920 -18337
rect 19886 -18439 19920 -18405
rect 20904 -17963 20938 -17929
rect 20904 -18031 20938 -17997
rect 20904 -18099 20938 -18065
rect 20904 -18167 20938 -18133
rect 20904 -18235 20938 -18201
rect 20904 -18303 20938 -18269
rect 20904 -18371 20938 -18337
rect 20904 -18439 20938 -18405
rect 21922 -17963 21956 -17929
rect 21922 -18031 21956 -17997
rect 21922 -18099 21956 -18065
rect 21922 -18167 21956 -18133
rect 21922 -18235 21956 -18201
rect 21922 -18303 21956 -18269
rect 21922 -18371 21956 -18337
rect 21922 -18439 21956 -18405
rect 22940 -17963 22974 -17929
rect 22940 -18031 22974 -17997
rect 22940 -18099 22974 -18065
rect 22940 -18167 22974 -18133
rect 22940 -18235 22974 -18201
rect 22940 -18303 22974 -18269
rect 22940 -18371 22974 -18337
rect 22940 -18439 22974 -18405
rect -22 -18521 12 -18487
rect -22 -18589 12 -18555
rect -22 -18657 12 -18623
rect -22 -18725 12 -18691
rect -22 -18793 12 -18759
rect 2580 -19197 2614 -19163
rect 2580 -19265 2614 -19231
rect 2580 -19333 2614 -19299
rect 2580 -19401 2614 -19367
rect 2580 -19469 2614 -19435
rect 2580 -19537 2614 -19503
rect 2580 -19605 2614 -19571
rect -2324 -19671 -2290 -19637
rect -2324 -19739 -2290 -19705
rect -2324 -19807 -2290 -19773
rect -2106 -19671 -2072 -19637
rect -2106 -19739 -2072 -19705
rect -2106 -19807 -2072 -19773
rect -1888 -19671 -1854 -19637
rect -1888 -19739 -1854 -19705
rect -1888 -19807 -1854 -19773
rect -1670 -19671 -1636 -19637
rect -1670 -19739 -1636 -19705
rect -1670 -19807 -1636 -19773
rect -1452 -19671 -1418 -19637
rect -1452 -19739 -1418 -19705
rect -1452 -19807 -1418 -19773
rect -1234 -19671 -1200 -19637
rect -1234 -19739 -1200 -19705
rect -1234 -19807 -1200 -19773
rect -1016 -19671 -982 -19637
rect -1016 -19739 -982 -19705
rect -1016 -19807 -982 -19773
rect -798 -19671 -764 -19637
rect -798 -19739 -764 -19705
rect -798 -19807 -764 -19773
rect -580 -19671 -546 -19637
rect -580 -19739 -546 -19705
rect -580 -19807 -546 -19773
rect -362 -19671 -328 -19637
rect -362 -19739 -328 -19705
rect -362 -19807 -328 -19773
rect -144 -19671 -110 -19637
rect -144 -19739 -110 -19705
rect 2580 -19673 2614 -19639
rect 3598 -19197 3632 -19163
rect 3598 -19265 3632 -19231
rect 3598 -19333 3632 -19299
rect 3598 -19401 3632 -19367
rect 3598 -19469 3632 -19435
rect 3598 -19537 3632 -19503
rect 3598 -19605 3632 -19571
rect 3598 -19673 3632 -19639
rect 4616 -19197 4650 -19163
rect 4616 -19265 4650 -19231
rect 4616 -19333 4650 -19299
rect 4616 -19401 4650 -19367
rect 4616 -19469 4650 -19435
rect 4616 -19537 4650 -19503
rect 4616 -19605 4650 -19571
rect 4616 -19673 4650 -19639
rect 5634 -19197 5668 -19163
rect 5634 -19265 5668 -19231
rect 5634 -19333 5668 -19299
rect 5634 -19401 5668 -19367
rect 5634 -19469 5668 -19435
rect 5634 -19537 5668 -19503
rect 5634 -19605 5668 -19571
rect 5634 -19673 5668 -19639
rect 6652 -19197 6686 -19163
rect 6652 -19265 6686 -19231
rect 6652 -19333 6686 -19299
rect 6652 -19401 6686 -19367
rect 6652 -19469 6686 -19435
rect 6652 -19537 6686 -19503
rect 6652 -19605 6686 -19571
rect 6652 -19673 6686 -19639
rect 7670 -19197 7704 -19163
rect 7670 -19265 7704 -19231
rect 7670 -19333 7704 -19299
rect 7670 -19401 7704 -19367
rect 7670 -19469 7704 -19435
rect 7670 -19537 7704 -19503
rect 7670 -19605 7704 -19571
rect 7670 -19673 7704 -19639
rect 8688 -19197 8722 -19163
rect 8688 -19265 8722 -19231
rect 8688 -19333 8722 -19299
rect 8688 -19401 8722 -19367
rect 8688 -19469 8722 -19435
rect 8688 -19537 8722 -19503
rect 8688 -19605 8722 -19571
rect 8688 -19673 8722 -19639
rect 9706 -19197 9740 -19163
rect 9706 -19265 9740 -19231
rect 9706 -19333 9740 -19299
rect 9706 -19401 9740 -19367
rect 9706 -19469 9740 -19435
rect 9706 -19537 9740 -19503
rect 9706 -19605 9740 -19571
rect 9706 -19673 9740 -19639
rect 10724 -19197 10758 -19163
rect 10724 -19265 10758 -19231
rect 10724 -19333 10758 -19299
rect 10724 -19401 10758 -19367
rect 10724 -19469 10758 -19435
rect 10724 -19537 10758 -19503
rect 10724 -19605 10758 -19571
rect 10724 -19673 10758 -19639
rect 11742 -19197 11776 -19163
rect 11742 -19265 11776 -19231
rect 11742 -19333 11776 -19299
rect 11742 -19401 11776 -19367
rect 11742 -19469 11776 -19435
rect 11742 -19537 11776 -19503
rect 11742 -19605 11776 -19571
rect 11742 -19673 11776 -19639
rect 12760 -19197 12794 -19163
rect 12760 -19265 12794 -19231
rect 12760 -19333 12794 -19299
rect 12760 -19401 12794 -19367
rect 12760 -19469 12794 -19435
rect 12760 -19537 12794 -19503
rect 12760 -19605 12794 -19571
rect 12760 -19673 12794 -19639
rect 13778 -19197 13812 -19163
rect 13778 -19265 13812 -19231
rect 13778 -19333 13812 -19299
rect 13778 -19401 13812 -19367
rect 13778 -19469 13812 -19435
rect 13778 -19537 13812 -19503
rect 13778 -19605 13812 -19571
rect 13778 -19673 13812 -19639
rect 14796 -19197 14830 -19163
rect 14796 -19265 14830 -19231
rect 14796 -19333 14830 -19299
rect 14796 -19401 14830 -19367
rect 14796 -19469 14830 -19435
rect 14796 -19537 14830 -19503
rect 14796 -19605 14830 -19571
rect 14796 -19673 14830 -19639
rect 15814 -19197 15848 -19163
rect 15814 -19265 15848 -19231
rect 15814 -19333 15848 -19299
rect 15814 -19401 15848 -19367
rect 15814 -19469 15848 -19435
rect 15814 -19537 15848 -19503
rect 15814 -19605 15848 -19571
rect 15814 -19673 15848 -19639
rect 16832 -19197 16866 -19163
rect 16832 -19265 16866 -19231
rect 16832 -19333 16866 -19299
rect 16832 -19401 16866 -19367
rect 16832 -19469 16866 -19435
rect 16832 -19537 16866 -19503
rect 16832 -19605 16866 -19571
rect 16832 -19673 16866 -19639
rect 17850 -19197 17884 -19163
rect 17850 -19265 17884 -19231
rect 17850 -19333 17884 -19299
rect 17850 -19401 17884 -19367
rect 17850 -19469 17884 -19435
rect 17850 -19537 17884 -19503
rect 17850 -19605 17884 -19571
rect 17850 -19673 17884 -19639
rect 18868 -19197 18902 -19163
rect 18868 -19265 18902 -19231
rect 18868 -19333 18902 -19299
rect 18868 -19401 18902 -19367
rect 18868 -19469 18902 -19435
rect 18868 -19537 18902 -19503
rect 18868 -19605 18902 -19571
rect 18868 -19673 18902 -19639
rect 19886 -19197 19920 -19163
rect 19886 -19265 19920 -19231
rect 19886 -19333 19920 -19299
rect 19886 -19401 19920 -19367
rect 19886 -19469 19920 -19435
rect 19886 -19537 19920 -19503
rect 19886 -19605 19920 -19571
rect 19886 -19673 19920 -19639
rect 20904 -19197 20938 -19163
rect 20904 -19265 20938 -19231
rect 20904 -19333 20938 -19299
rect 20904 -19401 20938 -19367
rect 20904 -19469 20938 -19435
rect 20904 -19537 20938 -19503
rect 20904 -19605 20938 -19571
rect 20904 -19673 20938 -19639
rect 21922 -19197 21956 -19163
rect 21922 -19265 21956 -19231
rect 21922 -19333 21956 -19299
rect 21922 -19401 21956 -19367
rect 21922 -19469 21956 -19435
rect 21922 -19537 21956 -19503
rect 21922 -19605 21956 -19571
rect 21922 -19673 21956 -19639
rect 22940 -19197 22974 -19163
rect 22940 -19265 22974 -19231
rect 22940 -19333 22974 -19299
rect 22940 -19401 22974 -19367
rect 22940 -19469 22974 -19435
rect 22940 -19537 22974 -19503
rect 22940 -19605 22974 -19571
rect 22940 -19673 22974 -19639
rect -144 -19807 -110 -19773
rect 2580 -20431 2614 -20397
rect -2324 -20503 -2290 -20469
rect -2324 -20571 -2290 -20537
rect -2324 -20639 -2290 -20605
rect -2106 -20503 -2072 -20469
rect -2106 -20571 -2072 -20537
rect -2106 -20639 -2072 -20605
rect -1888 -20503 -1854 -20469
rect -1888 -20571 -1854 -20537
rect -1888 -20639 -1854 -20605
rect -1670 -20503 -1636 -20469
rect -1670 -20571 -1636 -20537
rect -1670 -20639 -1636 -20605
rect -1452 -20503 -1418 -20469
rect -1452 -20571 -1418 -20537
rect -1452 -20639 -1418 -20605
rect -1234 -20503 -1200 -20469
rect -1234 -20571 -1200 -20537
rect -1234 -20639 -1200 -20605
rect -1016 -20503 -982 -20469
rect -1016 -20571 -982 -20537
rect -1016 -20639 -982 -20605
rect -798 -20503 -764 -20469
rect -798 -20571 -764 -20537
rect -798 -20639 -764 -20605
rect -580 -20503 -546 -20469
rect -580 -20571 -546 -20537
rect -580 -20639 -546 -20605
rect -362 -20503 -328 -20469
rect -362 -20571 -328 -20537
rect -362 -20639 -328 -20605
rect -144 -20503 -110 -20469
rect -144 -20571 -110 -20537
rect -144 -20639 -110 -20605
rect 2580 -20499 2614 -20465
rect 2580 -20567 2614 -20533
rect 2580 -20635 2614 -20601
rect 2580 -20703 2614 -20669
rect 2580 -20771 2614 -20737
rect 2580 -20839 2614 -20805
rect 2580 -20907 2614 -20873
rect 3598 -20431 3632 -20397
rect 3598 -20499 3632 -20465
rect 3598 -20567 3632 -20533
rect 3598 -20635 3632 -20601
rect 3598 -20703 3632 -20669
rect 3598 -20771 3632 -20737
rect 3598 -20839 3632 -20805
rect 3598 -20907 3632 -20873
rect 4616 -20431 4650 -20397
rect 4616 -20499 4650 -20465
rect 4616 -20567 4650 -20533
rect 4616 -20635 4650 -20601
rect 4616 -20703 4650 -20669
rect 4616 -20771 4650 -20737
rect 4616 -20839 4650 -20805
rect 4616 -20907 4650 -20873
rect 5634 -20431 5668 -20397
rect 5634 -20499 5668 -20465
rect 5634 -20567 5668 -20533
rect 5634 -20635 5668 -20601
rect 5634 -20703 5668 -20669
rect 5634 -20771 5668 -20737
rect 5634 -20839 5668 -20805
rect 5634 -20907 5668 -20873
rect 6652 -20431 6686 -20397
rect 6652 -20499 6686 -20465
rect 6652 -20567 6686 -20533
rect 6652 -20635 6686 -20601
rect 6652 -20703 6686 -20669
rect 6652 -20771 6686 -20737
rect 6652 -20839 6686 -20805
rect 6652 -20907 6686 -20873
rect 7670 -20431 7704 -20397
rect 7670 -20499 7704 -20465
rect 7670 -20567 7704 -20533
rect 7670 -20635 7704 -20601
rect 7670 -20703 7704 -20669
rect 7670 -20771 7704 -20737
rect 7670 -20839 7704 -20805
rect 7670 -20907 7704 -20873
rect 8688 -20431 8722 -20397
rect 8688 -20499 8722 -20465
rect 8688 -20567 8722 -20533
rect 8688 -20635 8722 -20601
rect 8688 -20703 8722 -20669
rect 8688 -20771 8722 -20737
rect 8688 -20839 8722 -20805
rect 8688 -20907 8722 -20873
rect 9706 -20431 9740 -20397
rect 9706 -20499 9740 -20465
rect 9706 -20567 9740 -20533
rect 9706 -20635 9740 -20601
rect 9706 -20703 9740 -20669
rect 9706 -20771 9740 -20737
rect 9706 -20839 9740 -20805
rect 9706 -20907 9740 -20873
rect 10724 -20431 10758 -20397
rect 10724 -20499 10758 -20465
rect 10724 -20567 10758 -20533
rect 10724 -20635 10758 -20601
rect 10724 -20703 10758 -20669
rect 10724 -20771 10758 -20737
rect 10724 -20839 10758 -20805
rect 10724 -20907 10758 -20873
rect 11742 -20431 11776 -20397
rect 11742 -20499 11776 -20465
rect 11742 -20567 11776 -20533
rect 11742 -20635 11776 -20601
rect 11742 -20703 11776 -20669
rect 11742 -20771 11776 -20737
rect 11742 -20839 11776 -20805
rect 11742 -20907 11776 -20873
rect 12760 -20431 12794 -20397
rect 12760 -20499 12794 -20465
rect 12760 -20567 12794 -20533
rect 12760 -20635 12794 -20601
rect 12760 -20703 12794 -20669
rect 12760 -20771 12794 -20737
rect 12760 -20839 12794 -20805
rect 12760 -20907 12794 -20873
rect 13778 -20431 13812 -20397
rect 13778 -20499 13812 -20465
rect 13778 -20567 13812 -20533
rect 13778 -20635 13812 -20601
rect 13778 -20703 13812 -20669
rect 13778 -20771 13812 -20737
rect 13778 -20839 13812 -20805
rect 13778 -20907 13812 -20873
rect 14796 -20431 14830 -20397
rect 14796 -20499 14830 -20465
rect 14796 -20567 14830 -20533
rect 14796 -20635 14830 -20601
rect 14796 -20703 14830 -20669
rect 14796 -20771 14830 -20737
rect 14796 -20839 14830 -20805
rect 14796 -20907 14830 -20873
rect 15814 -20431 15848 -20397
rect 15814 -20499 15848 -20465
rect 15814 -20567 15848 -20533
rect 15814 -20635 15848 -20601
rect 15814 -20703 15848 -20669
rect 15814 -20771 15848 -20737
rect 15814 -20839 15848 -20805
rect 15814 -20907 15848 -20873
rect 16832 -20431 16866 -20397
rect 16832 -20499 16866 -20465
rect 16832 -20567 16866 -20533
rect 16832 -20635 16866 -20601
rect 16832 -20703 16866 -20669
rect 16832 -20771 16866 -20737
rect 16832 -20839 16866 -20805
rect 16832 -20907 16866 -20873
rect 17850 -20431 17884 -20397
rect 17850 -20499 17884 -20465
rect 17850 -20567 17884 -20533
rect 17850 -20635 17884 -20601
rect 17850 -20703 17884 -20669
rect 17850 -20771 17884 -20737
rect 17850 -20839 17884 -20805
rect 17850 -20907 17884 -20873
rect 18868 -20431 18902 -20397
rect 18868 -20499 18902 -20465
rect 18868 -20567 18902 -20533
rect 18868 -20635 18902 -20601
rect 18868 -20703 18902 -20669
rect 18868 -20771 18902 -20737
rect 18868 -20839 18902 -20805
rect 18868 -20907 18902 -20873
rect 19886 -20431 19920 -20397
rect 19886 -20499 19920 -20465
rect 19886 -20567 19920 -20533
rect 19886 -20635 19920 -20601
rect 19886 -20703 19920 -20669
rect 19886 -20771 19920 -20737
rect 19886 -20839 19920 -20805
rect 19886 -20907 19920 -20873
rect 20904 -20431 20938 -20397
rect 20904 -20499 20938 -20465
rect 20904 -20567 20938 -20533
rect 20904 -20635 20938 -20601
rect 20904 -20703 20938 -20669
rect 20904 -20771 20938 -20737
rect 20904 -20839 20938 -20805
rect 20904 -20907 20938 -20873
rect 21922 -20431 21956 -20397
rect 21922 -20499 21956 -20465
rect 21922 -20567 21956 -20533
rect 21922 -20635 21956 -20601
rect 21922 -20703 21956 -20669
rect 21922 -20771 21956 -20737
rect 21922 -20839 21956 -20805
rect 21922 -20907 21956 -20873
rect 22940 -20431 22974 -20397
rect 22940 -20499 22974 -20465
rect 22940 -20567 22974 -20533
rect 22940 -20635 22974 -20601
rect 22940 -20703 22974 -20669
rect 22940 -20771 22974 -20737
rect 22940 -20839 22974 -20805
rect 22940 -20907 22974 -20873
rect 2580 -21663 2614 -21629
rect 2580 -21731 2614 -21697
rect -9405 -21860 -9371 -21826
rect -9405 -21928 -9371 -21894
rect -9405 -21996 -9371 -21962
rect -9405 -22064 -9371 -22030
rect -9405 -22132 -9371 -22098
rect -9405 -22200 -9371 -22166
rect -9405 -22268 -9371 -22234
rect -9405 -22336 -9371 -22302
rect -8387 -21860 -8353 -21826
rect -8387 -21928 -8353 -21894
rect -8387 -21996 -8353 -21962
rect -8387 -22064 -8353 -22030
rect -8387 -22132 -8353 -22098
rect -8387 -22200 -8353 -22166
rect -8387 -22268 -8353 -22234
rect -8387 -22336 -8353 -22302
rect -7369 -21860 -7335 -21826
rect -7369 -21928 -7335 -21894
rect -7369 -21996 -7335 -21962
rect -7369 -22064 -7335 -22030
rect -7369 -22132 -7335 -22098
rect -7369 -22200 -7335 -22166
rect -7369 -22268 -7335 -22234
rect -7369 -22336 -7335 -22302
rect -6351 -21860 -6317 -21826
rect -6351 -21928 -6317 -21894
rect -6351 -21996 -6317 -21962
rect -6351 -22064 -6317 -22030
rect -6351 -22132 -6317 -22098
rect -6351 -22200 -6317 -22166
rect -6351 -22268 -6317 -22234
rect -6351 -22336 -6317 -22302
rect -5333 -21860 -5299 -21826
rect -5333 -21928 -5299 -21894
rect -5333 -21996 -5299 -21962
rect -5333 -22064 -5299 -22030
rect -5333 -22132 -5299 -22098
rect -5333 -22200 -5299 -22166
rect -5333 -22268 -5299 -22234
rect -5333 -22336 -5299 -22302
rect -4315 -21860 -4281 -21826
rect -4315 -21928 -4281 -21894
rect -4315 -21996 -4281 -21962
rect -4315 -22064 -4281 -22030
rect -4315 -22132 -4281 -22098
rect -4315 -22200 -4281 -22166
rect -4315 -22268 -4281 -22234
rect -4315 -22336 -4281 -22302
rect -3297 -21860 -3263 -21826
rect -3297 -21928 -3263 -21894
rect -3297 -21996 -3263 -21962
rect -3297 -22064 -3263 -22030
rect -3297 -22132 -3263 -22098
rect -3297 -22200 -3263 -22166
rect -3297 -22268 -3263 -22234
rect -3297 -22336 -3263 -22302
rect -2410 -21859 -2376 -21825
rect -2410 -21927 -2376 -21893
rect -2410 -21995 -2376 -21961
rect -2410 -22063 -2376 -22029
rect -2410 -22131 -2376 -22097
rect -2410 -22199 -2376 -22165
rect -2410 -22267 -2376 -22233
rect -2410 -22335 -2376 -22301
rect -2112 -21859 -2078 -21825
rect -2112 -21927 -2078 -21893
rect -2112 -21995 -2078 -21961
rect -2112 -22063 -2078 -22029
rect -2112 -22131 -2078 -22097
rect -2112 -22199 -2078 -22165
rect -2112 -22267 -2078 -22233
rect -2112 -22335 -2078 -22301
rect -1814 -21859 -1780 -21825
rect -1814 -21927 -1780 -21893
rect -1814 -21995 -1780 -21961
rect -1814 -22063 -1780 -22029
rect -1814 -22131 -1780 -22097
rect -1814 -22199 -1780 -22165
rect -1814 -22267 -1780 -22233
rect -1814 -22335 -1780 -22301
rect -1516 -21859 -1482 -21825
rect -1516 -21927 -1482 -21893
rect -1516 -21995 -1482 -21961
rect -1516 -22063 -1482 -22029
rect -1516 -22131 -1482 -22097
rect -1516 -22199 -1482 -22165
rect -1516 -22267 -1482 -22233
rect -1516 -22335 -1482 -22301
rect -1218 -21859 -1184 -21825
rect -1218 -21927 -1184 -21893
rect -1218 -21995 -1184 -21961
rect -1218 -22063 -1184 -22029
rect -1218 -22131 -1184 -22097
rect -1218 -22199 -1184 -22165
rect -1218 -22267 -1184 -22233
rect -1218 -22335 -1184 -22301
rect -920 -21859 -886 -21825
rect -920 -21927 -886 -21893
rect -920 -21995 -886 -21961
rect -920 -22063 -886 -22029
rect -920 -22131 -886 -22097
rect -920 -22199 -886 -22165
rect -920 -22267 -886 -22233
rect -920 -22335 -886 -22301
rect -622 -21859 -588 -21825
rect -622 -21927 -588 -21893
rect -622 -21995 -588 -21961
rect -622 -22063 -588 -22029
rect -622 -22131 -588 -22097
rect -622 -22199 -588 -22165
rect -622 -22267 -588 -22233
rect -622 -22335 -588 -22301
rect -324 -21859 -290 -21825
rect -324 -21927 -290 -21893
rect -324 -21995 -290 -21961
rect -324 -22063 -290 -22029
rect -324 -22131 -290 -22097
rect -324 -22199 -290 -22165
rect -324 -22267 -290 -22233
rect -324 -22335 -290 -22301
rect -26 -21859 8 -21825
rect -26 -21927 8 -21893
rect -26 -21995 8 -21961
rect -26 -22063 8 -22029
rect -26 -22131 8 -22097
rect -26 -22199 8 -22165
rect -26 -22267 8 -22233
rect -26 -22335 8 -22301
rect 272 -21859 306 -21825
rect 272 -21927 306 -21893
rect 272 -21995 306 -21961
rect 272 -22063 306 -22029
rect 272 -22131 306 -22097
rect 272 -22199 306 -22165
rect 272 -22267 306 -22233
rect 272 -22335 306 -22301
rect 570 -21859 604 -21825
rect 570 -21927 604 -21893
rect 570 -21995 604 -21961
rect 570 -22063 604 -22029
rect 570 -22131 604 -22097
rect 570 -22199 604 -22165
rect 570 -22267 604 -22233
rect 570 -22335 604 -22301
rect 868 -21859 902 -21825
rect 868 -21927 902 -21893
rect 868 -21995 902 -21961
rect 868 -22063 902 -22029
rect 868 -22131 902 -22097
rect 868 -22199 902 -22165
rect 2580 -21799 2614 -21765
rect 2580 -21867 2614 -21833
rect 2580 -21935 2614 -21901
rect 2580 -22003 2614 -21969
rect 2580 -22071 2614 -22037
rect 2580 -22139 2614 -22105
rect 3598 -21663 3632 -21629
rect 3598 -21731 3632 -21697
rect 3598 -21799 3632 -21765
rect 3598 -21867 3632 -21833
rect 3598 -21935 3632 -21901
rect 3598 -22003 3632 -21969
rect 3598 -22071 3632 -22037
rect 3598 -22139 3632 -22105
rect 4616 -21663 4650 -21629
rect 4616 -21731 4650 -21697
rect 4616 -21799 4650 -21765
rect 4616 -21867 4650 -21833
rect 4616 -21935 4650 -21901
rect 4616 -22003 4650 -21969
rect 4616 -22071 4650 -22037
rect 4616 -22139 4650 -22105
rect 5634 -21663 5668 -21629
rect 5634 -21731 5668 -21697
rect 5634 -21799 5668 -21765
rect 5634 -21867 5668 -21833
rect 5634 -21935 5668 -21901
rect 5634 -22003 5668 -21969
rect 5634 -22071 5668 -22037
rect 5634 -22139 5668 -22105
rect 6652 -21663 6686 -21629
rect 6652 -21731 6686 -21697
rect 6652 -21799 6686 -21765
rect 6652 -21867 6686 -21833
rect 6652 -21935 6686 -21901
rect 6652 -22003 6686 -21969
rect 6652 -22071 6686 -22037
rect 6652 -22139 6686 -22105
rect 7670 -21663 7704 -21629
rect 7670 -21731 7704 -21697
rect 7670 -21799 7704 -21765
rect 7670 -21867 7704 -21833
rect 7670 -21935 7704 -21901
rect 7670 -22003 7704 -21969
rect 7670 -22071 7704 -22037
rect 7670 -22139 7704 -22105
rect 8688 -21663 8722 -21629
rect 8688 -21731 8722 -21697
rect 8688 -21799 8722 -21765
rect 8688 -21867 8722 -21833
rect 8688 -21935 8722 -21901
rect 8688 -22003 8722 -21969
rect 8688 -22071 8722 -22037
rect 8688 -22139 8722 -22105
rect 9706 -21663 9740 -21629
rect 9706 -21731 9740 -21697
rect 9706 -21799 9740 -21765
rect 9706 -21867 9740 -21833
rect 9706 -21935 9740 -21901
rect 9706 -22003 9740 -21969
rect 9706 -22071 9740 -22037
rect 9706 -22139 9740 -22105
rect 10724 -21663 10758 -21629
rect 10724 -21731 10758 -21697
rect 10724 -21799 10758 -21765
rect 10724 -21867 10758 -21833
rect 10724 -21935 10758 -21901
rect 10724 -22003 10758 -21969
rect 10724 -22071 10758 -22037
rect 10724 -22139 10758 -22105
rect 11742 -21663 11776 -21629
rect 11742 -21731 11776 -21697
rect 11742 -21799 11776 -21765
rect 11742 -21867 11776 -21833
rect 11742 -21935 11776 -21901
rect 11742 -22003 11776 -21969
rect 11742 -22071 11776 -22037
rect 11742 -22139 11776 -22105
rect 12760 -21663 12794 -21629
rect 12760 -21731 12794 -21697
rect 12760 -21799 12794 -21765
rect 12760 -21867 12794 -21833
rect 12760 -21935 12794 -21901
rect 12760 -22003 12794 -21969
rect 12760 -22071 12794 -22037
rect 12760 -22139 12794 -22105
rect 13778 -21663 13812 -21629
rect 13778 -21731 13812 -21697
rect 13778 -21799 13812 -21765
rect 13778 -21867 13812 -21833
rect 13778 -21935 13812 -21901
rect 13778 -22003 13812 -21969
rect 13778 -22071 13812 -22037
rect 13778 -22139 13812 -22105
rect 14796 -21663 14830 -21629
rect 14796 -21731 14830 -21697
rect 14796 -21799 14830 -21765
rect 14796 -21867 14830 -21833
rect 14796 -21935 14830 -21901
rect 14796 -22003 14830 -21969
rect 14796 -22071 14830 -22037
rect 14796 -22139 14830 -22105
rect 15814 -21663 15848 -21629
rect 15814 -21731 15848 -21697
rect 15814 -21799 15848 -21765
rect 15814 -21867 15848 -21833
rect 15814 -21935 15848 -21901
rect 15814 -22003 15848 -21969
rect 15814 -22071 15848 -22037
rect 15814 -22139 15848 -22105
rect 16832 -21663 16866 -21629
rect 16832 -21731 16866 -21697
rect 16832 -21799 16866 -21765
rect 16832 -21867 16866 -21833
rect 16832 -21935 16866 -21901
rect 16832 -22003 16866 -21969
rect 16832 -22071 16866 -22037
rect 16832 -22139 16866 -22105
rect 17850 -21663 17884 -21629
rect 17850 -21731 17884 -21697
rect 17850 -21799 17884 -21765
rect 17850 -21867 17884 -21833
rect 17850 -21935 17884 -21901
rect 17850 -22003 17884 -21969
rect 17850 -22071 17884 -22037
rect 17850 -22139 17884 -22105
rect 18868 -21663 18902 -21629
rect 18868 -21731 18902 -21697
rect 18868 -21799 18902 -21765
rect 18868 -21867 18902 -21833
rect 18868 -21935 18902 -21901
rect 18868 -22003 18902 -21969
rect 18868 -22071 18902 -22037
rect 18868 -22139 18902 -22105
rect 19886 -21663 19920 -21629
rect 19886 -21731 19920 -21697
rect 19886 -21799 19920 -21765
rect 19886 -21867 19920 -21833
rect 19886 -21935 19920 -21901
rect 19886 -22003 19920 -21969
rect 19886 -22071 19920 -22037
rect 19886 -22139 19920 -22105
rect 20904 -21663 20938 -21629
rect 20904 -21731 20938 -21697
rect 20904 -21799 20938 -21765
rect 20904 -21867 20938 -21833
rect 20904 -21935 20938 -21901
rect 20904 -22003 20938 -21969
rect 20904 -22071 20938 -22037
rect 20904 -22139 20938 -22105
rect 21922 -21663 21956 -21629
rect 21922 -21731 21956 -21697
rect 21922 -21799 21956 -21765
rect 21922 -21867 21956 -21833
rect 21922 -21935 21956 -21901
rect 21922 -22003 21956 -21969
rect 21922 -22071 21956 -22037
rect 21922 -22139 21956 -22105
rect 22940 -21663 22974 -21629
rect 22940 -21731 22974 -21697
rect 22940 -21799 22974 -21765
rect 22940 -21867 22974 -21833
rect 22940 -21935 22974 -21901
rect 22940 -22003 22974 -21969
rect 22940 -22071 22974 -22037
rect 22940 -22139 22974 -22105
rect 868 -22267 902 -22233
rect 868 -22335 902 -22301
rect -9406 -22973 -9372 -22939
rect -9406 -23041 -9372 -23007
rect -9406 -23109 -9372 -23075
rect -9406 -23177 -9372 -23143
rect -9406 -23245 -9372 -23211
rect -9406 -23313 -9372 -23279
rect -9406 -23381 -9372 -23347
rect -9406 -23449 -9372 -23415
rect -8388 -22973 -8354 -22939
rect -8388 -23041 -8354 -23007
rect -8388 -23109 -8354 -23075
rect -8388 -23177 -8354 -23143
rect -8388 -23245 -8354 -23211
rect -8388 -23313 -8354 -23279
rect -8388 -23381 -8354 -23347
rect -8388 -23449 -8354 -23415
rect -7370 -22973 -7336 -22939
rect -7370 -23041 -7336 -23007
rect -7370 -23109 -7336 -23075
rect -7370 -23177 -7336 -23143
rect -7370 -23245 -7336 -23211
rect -7370 -23313 -7336 -23279
rect -7370 -23381 -7336 -23347
rect -7370 -23449 -7336 -23415
rect -6352 -22973 -6318 -22939
rect -6352 -23041 -6318 -23007
rect -6352 -23109 -6318 -23075
rect -6352 -23177 -6318 -23143
rect -6352 -23245 -6318 -23211
rect -6352 -23313 -6318 -23279
rect -6352 -23381 -6318 -23347
rect -6352 -23449 -6318 -23415
rect -5334 -22973 -5300 -22939
rect -5334 -23041 -5300 -23007
rect -5334 -23109 -5300 -23075
rect -5334 -23177 -5300 -23143
rect -5334 -23245 -5300 -23211
rect -5334 -23313 -5300 -23279
rect -5334 -23381 -5300 -23347
rect -5334 -23449 -5300 -23415
rect -4316 -22973 -4282 -22939
rect -4316 -23041 -4282 -23007
rect -4316 -23109 -4282 -23075
rect -4316 -23177 -4282 -23143
rect -4316 -23245 -4282 -23211
rect -4316 -23313 -4282 -23279
rect -4316 -23381 -4282 -23347
rect -4316 -23449 -4282 -23415
rect -3298 -22973 -3264 -22939
rect -3298 -23041 -3264 -23007
rect -3298 -23109 -3264 -23075
rect -3298 -23177 -3264 -23143
rect -3298 -23245 -3264 -23211
rect -3298 -23313 -3264 -23279
rect -3298 -23381 -3264 -23347
rect -3298 -23449 -3264 -23415
rect -2410 -22971 -2376 -22937
rect -2410 -23039 -2376 -23005
rect -2410 -23107 -2376 -23073
rect -2410 -23175 -2376 -23141
rect -2410 -23243 -2376 -23209
rect -2410 -23311 -2376 -23277
rect -2410 -23379 -2376 -23345
rect -2410 -23447 -2376 -23413
rect -2112 -22971 -2078 -22937
rect -2112 -23039 -2078 -23005
rect -2112 -23107 -2078 -23073
rect -2112 -23175 -2078 -23141
rect -2112 -23243 -2078 -23209
rect -2112 -23311 -2078 -23277
rect -2112 -23379 -2078 -23345
rect -2112 -23447 -2078 -23413
rect -1814 -22971 -1780 -22937
rect -1814 -23039 -1780 -23005
rect -1814 -23107 -1780 -23073
rect -1814 -23175 -1780 -23141
rect -1814 -23243 -1780 -23209
rect -1814 -23311 -1780 -23277
rect -1814 -23379 -1780 -23345
rect -1814 -23447 -1780 -23413
rect -1516 -22971 -1482 -22937
rect -1516 -23039 -1482 -23005
rect -1516 -23107 -1482 -23073
rect -1516 -23175 -1482 -23141
rect -1516 -23243 -1482 -23209
rect -1516 -23311 -1482 -23277
rect -1516 -23379 -1482 -23345
rect -1516 -23447 -1482 -23413
rect -1218 -22971 -1184 -22937
rect -1218 -23039 -1184 -23005
rect -1218 -23107 -1184 -23073
rect -1218 -23175 -1184 -23141
rect -1218 -23243 -1184 -23209
rect -1218 -23311 -1184 -23277
rect -1218 -23379 -1184 -23345
rect -1218 -23447 -1184 -23413
rect -920 -22971 -886 -22937
rect -920 -23039 -886 -23005
rect -920 -23107 -886 -23073
rect -920 -23175 -886 -23141
rect -920 -23243 -886 -23209
rect -920 -23311 -886 -23277
rect -920 -23379 -886 -23345
rect -920 -23447 -886 -23413
rect -622 -22971 -588 -22937
rect -622 -23039 -588 -23005
rect -622 -23107 -588 -23073
rect -622 -23175 -588 -23141
rect -622 -23243 -588 -23209
rect -622 -23311 -588 -23277
rect -622 -23379 -588 -23345
rect -622 -23447 -588 -23413
rect -324 -22971 -290 -22937
rect -324 -23039 -290 -23005
rect -324 -23107 -290 -23073
rect -324 -23175 -290 -23141
rect -324 -23243 -290 -23209
rect -324 -23311 -290 -23277
rect -324 -23379 -290 -23345
rect -324 -23447 -290 -23413
rect -26 -22971 8 -22937
rect -26 -23039 8 -23005
rect -26 -23107 8 -23073
rect -26 -23175 8 -23141
rect -26 -23243 8 -23209
rect -26 -23311 8 -23277
rect -26 -23379 8 -23345
rect -26 -23447 8 -23413
rect 272 -22971 306 -22937
rect 272 -23039 306 -23005
rect 272 -23107 306 -23073
rect 272 -23175 306 -23141
rect 272 -23243 306 -23209
rect 272 -23311 306 -23277
rect 272 -23379 306 -23345
rect 272 -23447 306 -23413
rect 570 -22971 604 -22937
rect 570 -23039 604 -23005
rect 570 -23107 604 -23073
rect 570 -23175 604 -23141
rect 570 -23243 604 -23209
rect 570 -23311 604 -23277
rect 570 -23379 604 -23345
rect 570 -23447 604 -23413
rect 868 -22971 902 -22937
rect 868 -23039 902 -23005
rect 868 -23107 902 -23073
rect 868 -23175 902 -23141
rect 868 -23243 902 -23209
rect 868 -23311 902 -23277
rect 868 -23379 902 -23345
rect 868 -23447 902 -23413
rect 2580 -22897 2614 -22863
rect 2580 -22965 2614 -22931
rect 2580 -23033 2614 -22999
rect 2580 -23101 2614 -23067
rect 2580 -23169 2614 -23135
rect 2580 -23237 2614 -23203
rect 2580 -23305 2614 -23271
rect 2580 -23373 2614 -23339
rect 3598 -22897 3632 -22863
rect 3598 -22965 3632 -22931
rect 3598 -23033 3632 -22999
rect 3598 -23101 3632 -23067
rect 3598 -23169 3632 -23135
rect 3598 -23237 3632 -23203
rect 3598 -23305 3632 -23271
rect 3598 -23373 3632 -23339
rect 4616 -22897 4650 -22863
rect 4616 -22965 4650 -22931
rect 4616 -23033 4650 -22999
rect 4616 -23101 4650 -23067
rect 4616 -23169 4650 -23135
rect 4616 -23237 4650 -23203
rect 4616 -23305 4650 -23271
rect 4616 -23373 4650 -23339
rect 5634 -22897 5668 -22863
rect 5634 -22965 5668 -22931
rect 5634 -23033 5668 -22999
rect 5634 -23101 5668 -23067
rect 5634 -23169 5668 -23135
rect 5634 -23237 5668 -23203
rect 5634 -23305 5668 -23271
rect 5634 -23373 5668 -23339
rect 6652 -22897 6686 -22863
rect 6652 -22965 6686 -22931
rect 6652 -23033 6686 -22999
rect 6652 -23101 6686 -23067
rect 6652 -23169 6686 -23135
rect 6652 -23237 6686 -23203
rect 6652 -23305 6686 -23271
rect 6652 -23373 6686 -23339
rect 7670 -22897 7704 -22863
rect 7670 -22965 7704 -22931
rect 7670 -23033 7704 -22999
rect 7670 -23101 7704 -23067
rect 7670 -23169 7704 -23135
rect 7670 -23237 7704 -23203
rect 7670 -23305 7704 -23271
rect 7670 -23373 7704 -23339
rect 8688 -22897 8722 -22863
rect 8688 -22965 8722 -22931
rect 8688 -23033 8722 -22999
rect 8688 -23101 8722 -23067
rect 8688 -23169 8722 -23135
rect 8688 -23237 8722 -23203
rect 8688 -23305 8722 -23271
rect 8688 -23373 8722 -23339
rect 9706 -22897 9740 -22863
rect 9706 -22965 9740 -22931
rect 9706 -23033 9740 -22999
rect 9706 -23101 9740 -23067
rect 9706 -23169 9740 -23135
rect 9706 -23237 9740 -23203
rect 9706 -23305 9740 -23271
rect 9706 -23373 9740 -23339
rect 10724 -22897 10758 -22863
rect 10724 -22965 10758 -22931
rect 10724 -23033 10758 -22999
rect 10724 -23101 10758 -23067
rect 10724 -23169 10758 -23135
rect 10724 -23237 10758 -23203
rect 10724 -23305 10758 -23271
rect 10724 -23373 10758 -23339
rect 11742 -22897 11776 -22863
rect 11742 -22965 11776 -22931
rect 11742 -23033 11776 -22999
rect 11742 -23101 11776 -23067
rect 11742 -23169 11776 -23135
rect 11742 -23237 11776 -23203
rect 11742 -23305 11776 -23271
rect 11742 -23373 11776 -23339
rect 12760 -22897 12794 -22863
rect 12760 -22965 12794 -22931
rect 12760 -23033 12794 -22999
rect 12760 -23101 12794 -23067
rect 12760 -23169 12794 -23135
rect 12760 -23237 12794 -23203
rect 12760 -23305 12794 -23271
rect 12760 -23373 12794 -23339
rect 13778 -22897 13812 -22863
rect 13778 -22965 13812 -22931
rect 13778 -23033 13812 -22999
rect 13778 -23101 13812 -23067
rect 13778 -23169 13812 -23135
rect 13778 -23237 13812 -23203
rect 13778 -23305 13812 -23271
rect 13778 -23373 13812 -23339
rect 14796 -22897 14830 -22863
rect 14796 -22965 14830 -22931
rect 14796 -23033 14830 -22999
rect 14796 -23101 14830 -23067
rect 14796 -23169 14830 -23135
rect 14796 -23237 14830 -23203
rect 14796 -23305 14830 -23271
rect 14796 -23373 14830 -23339
rect 15814 -22897 15848 -22863
rect 15814 -22965 15848 -22931
rect 15814 -23033 15848 -22999
rect 15814 -23101 15848 -23067
rect 15814 -23169 15848 -23135
rect 15814 -23237 15848 -23203
rect 15814 -23305 15848 -23271
rect 15814 -23373 15848 -23339
rect 16832 -22897 16866 -22863
rect 16832 -22965 16866 -22931
rect 16832 -23033 16866 -22999
rect 16832 -23101 16866 -23067
rect 16832 -23169 16866 -23135
rect 16832 -23237 16866 -23203
rect 16832 -23305 16866 -23271
rect 16832 -23373 16866 -23339
rect 17850 -22897 17884 -22863
rect 17850 -22965 17884 -22931
rect 17850 -23033 17884 -22999
rect 17850 -23101 17884 -23067
rect 17850 -23169 17884 -23135
rect 17850 -23237 17884 -23203
rect 17850 -23305 17884 -23271
rect 17850 -23373 17884 -23339
rect 18868 -22897 18902 -22863
rect 18868 -22965 18902 -22931
rect 18868 -23033 18902 -22999
rect 18868 -23101 18902 -23067
rect 18868 -23169 18902 -23135
rect 18868 -23237 18902 -23203
rect 18868 -23305 18902 -23271
rect 18868 -23373 18902 -23339
rect 19886 -22897 19920 -22863
rect 19886 -22965 19920 -22931
rect 19886 -23033 19920 -22999
rect 19886 -23101 19920 -23067
rect 19886 -23169 19920 -23135
rect 19886 -23237 19920 -23203
rect 19886 -23305 19920 -23271
rect 19886 -23373 19920 -23339
rect 20904 -22897 20938 -22863
rect 20904 -22965 20938 -22931
rect 20904 -23033 20938 -22999
rect 20904 -23101 20938 -23067
rect 20904 -23169 20938 -23135
rect 20904 -23237 20938 -23203
rect 20904 -23305 20938 -23271
rect 20904 -23373 20938 -23339
rect 21922 -22897 21956 -22863
rect 21922 -22965 21956 -22931
rect 21922 -23033 21956 -22999
rect 21922 -23101 21956 -23067
rect 21922 -23169 21956 -23135
rect 21922 -23237 21956 -23203
rect 21922 -23305 21956 -23271
rect 21922 -23373 21956 -23339
rect 22940 -22897 22974 -22863
rect 22940 -22965 22974 -22931
rect 22940 -23033 22974 -22999
rect 22940 -23101 22974 -23067
rect 22940 -23169 22974 -23135
rect 22940 -23237 22974 -23203
rect 22940 -23305 22974 -23271
rect 22940 -23373 22974 -23339
rect -9405 -24084 -9371 -24050
rect -9405 -24152 -9371 -24118
rect -9405 -24220 -9371 -24186
rect -9405 -24288 -9371 -24254
rect -9405 -24356 -9371 -24322
rect -9405 -24424 -9371 -24390
rect -9405 -24492 -9371 -24458
rect -9405 -24560 -9371 -24526
rect -8387 -24084 -8353 -24050
rect -8387 -24152 -8353 -24118
rect -8387 -24220 -8353 -24186
rect -8387 -24288 -8353 -24254
rect -8387 -24356 -8353 -24322
rect -8387 -24424 -8353 -24390
rect -8387 -24492 -8353 -24458
rect -8387 -24560 -8353 -24526
rect -7369 -24084 -7335 -24050
rect -7369 -24152 -7335 -24118
rect -7369 -24220 -7335 -24186
rect -7369 -24288 -7335 -24254
rect -7369 -24356 -7335 -24322
rect -7369 -24424 -7335 -24390
rect -7369 -24492 -7335 -24458
rect -7369 -24560 -7335 -24526
rect -6351 -24084 -6317 -24050
rect -6351 -24152 -6317 -24118
rect -6351 -24220 -6317 -24186
rect -6351 -24288 -6317 -24254
rect -6351 -24356 -6317 -24322
rect -6351 -24424 -6317 -24390
rect -6351 -24492 -6317 -24458
rect -6351 -24560 -6317 -24526
rect -5333 -24084 -5299 -24050
rect -5333 -24152 -5299 -24118
rect -5333 -24220 -5299 -24186
rect -5333 -24288 -5299 -24254
rect -5333 -24356 -5299 -24322
rect -5333 -24424 -5299 -24390
rect -5333 -24492 -5299 -24458
rect -5333 -24560 -5299 -24526
rect -4315 -24084 -4281 -24050
rect -4315 -24152 -4281 -24118
rect -4315 -24220 -4281 -24186
rect -4315 -24288 -4281 -24254
rect -4315 -24356 -4281 -24322
rect -4315 -24424 -4281 -24390
rect -4315 -24492 -4281 -24458
rect -4315 -24560 -4281 -24526
rect -3297 -24084 -3263 -24050
rect -3297 -24152 -3263 -24118
rect -3297 -24220 -3263 -24186
rect -3297 -24288 -3263 -24254
rect -3297 -24356 -3263 -24322
rect -3297 -24424 -3263 -24390
rect -3297 -24492 -3263 -24458
rect -3297 -24560 -3263 -24526
rect -2412 -24083 -2378 -24049
rect -2412 -24151 -2378 -24117
rect -2412 -24219 -2378 -24185
rect -2412 -24287 -2378 -24253
rect -2412 -24355 -2378 -24321
rect -2412 -24423 -2378 -24389
rect -2412 -24491 -2378 -24457
rect -2412 -24559 -2378 -24525
rect -2114 -24083 -2080 -24049
rect -2114 -24151 -2080 -24117
rect -2114 -24219 -2080 -24185
rect -2114 -24287 -2080 -24253
rect -2114 -24355 -2080 -24321
rect -2114 -24423 -2080 -24389
rect -2114 -24491 -2080 -24457
rect -2114 -24559 -2080 -24525
rect -1816 -24083 -1782 -24049
rect -1816 -24151 -1782 -24117
rect -1816 -24219 -1782 -24185
rect -1816 -24287 -1782 -24253
rect -1816 -24355 -1782 -24321
rect -1816 -24423 -1782 -24389
rect -1816 -24491 -1782 -24457
rect -1816 -24559 -1782 -24525
rect -1518 -24083 -1484 -24049
rect -1518 -24151 -1484 -24117
rect -1518 -24219 -1484 -24185
rect -1518 -24287 -1484 -24253
rect -1518 -24355 -1484 -24321
rect -1518 -24423 -1484 -24389
rect -1518 -24491 -1484 -24457
rect -1518 -24559 -1484 -24525
rect -1220 -24083 -1186 -24049
rect -1220 -24151 -1186 -24117
rect -1220 -24219 -1186 -24185
rect -1220 -24287 -1186 -24253
rect -1220 -24355 -1186 -24321
rect -1220 -24423 -1186 -24389
rect -1220 -24491 -1186 -24457
rect -1220 -24559 -1186 -24525
rect -922 -24083 -888 -24049
rect -922 -24151 -888 -24117
rect -922 -24219 -888 -24185
rect -922 -24287 -888 -24253
rect -922 -24355 -888 -24321
rect -922 -24423 -888 -24389
rect -922 -24491 -888 -24457
rect -922 -24559 -888 -24525
rect -624 -24083 -590 -24049
rect -624 -24151 -590 -24117
rect -624 -24219 -590 -24185
rect -624 -24287 -590 -24253
rect -624 -24355 -590 -24321
rect -624 -24423 -590 -24389
rect -624 -24491 -590 -24457
rect -624 -24559 -590 -24525
rect -326 -24083 -292 -24049
rect -326 -24151 -292 -24117
rect -326 -24219 -292 -24185
rect -326 -24287 -292 -24253
rect -326 -24355 -292 -24321
rect -326 -24423 -292 -24389
rect -326 -24491 -292 -24457
rect -326 -24559 -292 -24525
rect -28 -24083 6 -24049
rect -28 -24151 6 -24117
rect -28 -24219 6 -24185
rect -28 -24287 6 -24253
rect -28 -24355 6 -24321
rect -28 -24423 6 -24389
rect -28 -24491 6 -24457
rect -28 -24559 6 -24525
rect 270 -24083 304 -24049
rect 270 -24151 304 -24117
rect 270 -24219 304 -24185
rect 270 -24287 304 -24253
rect 270 -24355 304 -24321
rect 270 -24423 304 -24389
rect 270 -24491 304 -24457
rect 270 -24559 304 -24525
rect 568 -24083 602 -24049
rect 568 -24151 602 -24117
rect 568 -24219 602 -24185
rect 568 -24287 602 -24253
rect 568 -24355 602 -24321
rect 568 -24423 602 -24389
rect 568 -24491 602 -24457
rect 568 -24559 602 -24525
rect 866 -24083 900 -24049
rect 866 -24151 900 -24117
rect 866 -24219 900 -24185
rect 866 -24287 900 -24253
rect 866 -24355 900 -24321
rect 866 -24423 900 -24389
rect 866 -24491 900 -24457
rect 866 -24559 900 -24525
rect 2580 -24131 2614 -24097
rect 2580 -24199 2614 -24165
rect 2580 -24267 2614 -24233
rect 2580 -24335 2614 -24301
rect 2580 -24403 2614 -24369
rect 2580 -24471 2614 -24437
rect 2580 -24539 2614 -24505
rect 2580 -24607 2614 -24573
rect 3598 -24131 3632 -24097
rect 3598 -24199 3632 -24165
rect 3598 -24267 3632 -24233
rect 3598 -24335 3632 -24301
rect 3598 -24403 3632 -24369
rect 3598 -24471 3632 -24437
rect 3598 -24539 3632 -24505
rect 3598 -24607 3632 -24573
rect 4616 -24131 4650 -24097
rect 4616 -24199 4650 -24165
rect 4616 -24267 4650 -24233
rect 4616 -24335 4650 -24301
rect 4616 -24403 4650 -24369
rect 4616 -24471 4650 -24437
rect 4616 -24539 4650 -24505
rect 4616 -24607 4650 -24573
rect 5634 -24131 5668 -24097
rect 5634 -24199 5668 -24165
rect 5634 -24267 5668 -24233
rect 5634 -24335 5668 -24301
rect 5634 -24403 5668 -24369
rect 5634 -24471 5668 -24437
rect 5634 -24539 5668 -24505
rect 5634 -24607 5668 -24573
rect 6652 -24131 6686 -24097
rect 6652 -24199 6686 -24165
rect 6652 -24267 6686 -24233
rect 6652 -24335 6686 -24301
rect 6652 -24403 6686 -24369
rect 6652 -24471 6686 -24437
rect 6652 -24539 6686 -24505
rect 6652 -24607 6686 -24573
rect 7670 -24131 7704 -24097
rect 7670 -24199 7704 -24165
rect 7670 -24267 7704 -24233
rect 7670 -24335 7704 -24301
rect 7670 -24403 7704 -24369
rect 7670 -24471 7704 -24437
rect 7670 -24539 7704 -24505
rect 7670 -24607 7704 -24573
rect 8688 -24131 8722 -24097
rect 8688 -24199 8722 -24165
rect 8688 -24267 8722 -24233
rect 8688 -24335 8722 -24301
rect 8688 -24403 8722 -24369
rect 8688 -24471 8722 -24437
rect 8688 -24539 8722 -24505
rect 8688 -24607 8722 -24573
rect 9706 -24131 9740 -24097
rect 9706 -24199 9740 -24165
rect 9706 -24267 9740 -24233
rect 9706 -24335 9740 -24301
rect 9706 -24403 9740 -24369
rect 9706 -24471 9740 -24437
rect 9706 -24539 9740 -24505
rect 9706 -24607 9740 -24573
rect 10724 -24131 10758 -24097
rect 10724 -24199 10758 -24165
rect 10724 -24267 10758 -24233
rect 10724 -24335 10758 -24301
rect 10724 -24403 10758 -24369
rect 10724 -24471 10758 -24437
rect 10724 -24539 10758 -24505
rect 10724 -24607 10758 -24573
rect 11742 -24131 11776 -24097
rect 11742 -24199 11776 -24165
rect 11742 -24267 11776 -24233
rect 11742 -24335 11776 -24301
rect 11742 -24403 11776 -24369
rect 11742 -24471 11776 -24437
rect 11742 -24539 11776 -24505
rect 11742 -24607 11776 -24573
rect 12760 -24131 12794 -24097
rect 12760 -24199 12794 -24165
rect 12760 -24267 12794 -24233
rect 12760 -24335 12794 -24301
rect 12760 -24403 12794 -24369
rect 12760 -24471 12794 -24437
rect 12760 -24539 12794 -24505
rect 12760 -24607 12794 -24573
rect 13778 -24131 13812 -24097
rect 13778 -24199 13812 -24165
rect 13778 -24267 13812 -24233
rect 13778 -24335 13812 -24301
rect 13778 -24403 13812 -24369
rect 13778 -24471 13812 -24437
rect 13778 -24539 13812 -24505
rect 13778 -24607 13812 -24573
rect 14796 -24131 14830 -24097
rect 14796 -24199 14830 -24165
rect 14796 -24267 14830 -24233
rect 14796 -24335 14830 -24301
rect 14796 -24403 14830 -24369
rect 14796 -24471 14830 -24437
rect 14796 -24539 14830 -24505
rect 14796 -24607 14830 -24573
rect 15814 -24131 15848 -24097
rect 15814 -24199 15848 -24165
rect 15814 -24267 15848 -24233
rect 15814 -24335 15848 -24301
rect 15814 -24403 15848 -24369
rect 15814 -24471 15848 -24437
rect 15814 -24539 15848 -24505
rect 15814 -24607 15848 -24573
rect 16832 -24131 16866 -24097
rect 16832 -24199 16866 -24165
rect 16832 -24267 16866 -24233
rect 16832 -24335 16866 -24301
rect 16832 -24403 16866 -24369
rect 16832 -24471 16866 -24437
rect 16832 -24539 16866 -24505
rect 16832 -24607 16866 -24573
rect 17850 -24131 17884 -24097
rect 17850 -24199 17884 -24165
rect 17850 -24267 17884 -24233
rect 17850 -24335 17884 -24301
rect 17850 -24403 17884 -24369
rect 17850 -24471 17884 -24437
rect 17850 -24539 17884 -24505
rect 17850 -24607 17884 -24573
rect 18868 -24131 18902 -24097
rect 18868 -24199 18902 -24165
rect 18868 -24267 18902 -24233
rect 18868 -24335 18902 -24301
rect 18868 -24403 18902 -24369
rect 18868 -24471 18902 -24437
rect 18868 -24539 18902 -24505
rect 18868 -24607 18902 -24573
rect 19886 -24131 19920 -24097
rect 19886 -24199 19920 -24165
rect 19886 -24267 19920 -24233
rect 19886 -24335 19920 -24301
rect 19886 -24403 19920 -24369
rect 19886 -24471 19920 -24437
rect 19886 -24539 19920 -24505
rect 19886 -24607 19920 -24573
rect 20904 -24131 20938 -24097
rect 20904 -24199 20938 -24165
rect 20904 -24267 20938 -24233
rect 20904 -24335 20938 -24301
rect 20904 -24403 20938 -24369
rect 20904 -24471 20938 -24437
rect 20904 -24539 20938 -24505
rect 20904 -24607 20938 -24573
rect 21922 -24131 21956 -24097
rect 21922 -24199 21956 -24165
rect 21922 -24267 21956 -24233
rect 21922 -24335 21956 -24301
rect 21922 -24403 21956 -24369
rect 21922 -24471 21956 -24437
rect 21922 -24539 21956 -24505
rect 21922 -24607 21956 -24573
rect 22940 -24131 22974 -24097
rect 22940 -24199 22974 -24165
rect 22940 -24267 22974 -24233
rect 22940 -24335 22974 -24301
rect 22940 -24403 22974 -24369
rect 22940 -24471 22974 -24437
rect 22940 -24539 22974 -24505
rect 22940 -24607 22974 -24573
rect -9406 -25197 -9372 -25163
rect -9406 -25265 -9372 -25231
rect -9406 -25333 -9372 -25299
rect -9406 -25401 -9372 -25367
rect -9406 -25469 -9372 -25435
rect -9406 -25537 -9372 -25503
rect -9406 -25605 -9372 -25571
rect -9406 -25673 -9372 -25639
rect -8388 -25197 -8354 -25163
rect -8388 -25265 -8354 -25231
rect -8388 -25333 -8354 -25299
rect -8388 -25401 -8354 -25367
rect -8388 -25469 -8354 -25435
rect -8388 -25537 -8354 -25503
rect -8388 -25605 -8354 -25571
rect -8388 -25673 -8354 -25639
rect -7370 -25197 -7336 -25163
rect -7370 -25265 -7336 -25231
rect -7370 -25333 -7336 -25299
rect -7370 -25401 -7336 -25367
rect -7370 -25469 -7336 -25435
rect -7370 -25537 -7336 -25503
rect -7370 -25605 -7336 -25571
rect -7370 -25673 -7336 -25639
rect -6352 -25197 -6318 -25163
rect -6352 -25265 -6318 -25231
rect -6352 -25333 -6318 -25299
rect -6352 -25401 -6318 -25367
rect -6352 -25469 -6318 -25435
rect -6352 -25537 -6318 -25503
rect -6352 -25605 -6318 -25571
rect -6352 -25673 -6318 -25639
rect -5334 -25197 -5300 -25163
rect -5334 -25265 -5300 -25231
rect -5334 -25333 -5300 -25299
rect -5334 -25401 -5300 -25367
rect -5334 -25469 -5300 -25435
rect -5334 -25537 -5300 -25503
rect -5334 -25605 -5300 -25571
rect -5334 -25673 -5300 -25639
rect -4316 -25197 -4282 -25163
rect -4316 -25265 -4282 -25231
rect -4316 -25333 -4282 -25299
rect -4316 -25401 -4282 -25367
rect -4316 -25469 -4282 -25435
rect -4316 -25537 -4282 -25503
rect -4316 -25605 -4282 -25571
rect -4316 -25673 -4282 -25639
rect -3298 -25197 -3264 -25163
rect -3298 -25265 -3264 -25231
rect -3298 -25333 -3264 -25299
rect -3298 -25401 -3264 -25367
rect -3298 -25469 -3264 -25435
rect -3298 -25537 -3264 -25503
rect -3298 -25605 -3264 -25571
rect -3298 -25673 -3264 -25639
rect -2412 -25193 -2378 -25159
rect -2412 -25261 -2378 -25227
rect -2412 -25329 -2378 -25295
rect -2412 -25397 -2378 -25363
rect -2412 -25465 -2378 -25431
rect -2412 -25533 -2378 -25499
rect -2412 -25601 -2378 -25567
rect -2412 -25669 -2378 -25635
rect -2114 -25193 -2080 -25159
rect -2114 -25261 -2080 -25227
rect -2114 -25329 -2080 -25295
rect -2114 -25397 -2080 -25363
rect -2114 -25465 -2080 -25431
rect -2114 -25533 -2080 -25499
rect -2114 -25601 -2080 -25567
rect -2114 -25669 -2080 -25635
rect -1816 -25193 -1782 -25159
rect -1816 -25261 -1782 -25227
rect -1816 -25329 -1782 -25295
rect -1816 -25397 -1782 -25363
rect -1816 -25465 -1782 -25431
rect -1816 -25533 -1782 -25499
rect -1816 -25601 -1782 -25567
rect -1816 -25669 -1782 -25635
rect -1518 -25193 -1484 -25159
rect -1518 -25261 -1484 -25227
rect -1518 -25329 -1484 -25295
rect -1518 -25397 -1484 -25363
rect -1518 -25465 -1484 -25431
rect -1518 -25533 -1484 -25499
rect -1518 -25601 -1484 -25567
rect -1518 -25669 -1484 -25635
rect -1220 -25193 -1186 -25159
rect -1220 -25261 -1186 -25227
rect -1220 -25329 -1186 -25295
rect -1220 -25397 -1186 -25363
rect -1220 -25465 -1186 -25431
rect -1220 -25533 -1186 -25499
rect -1220 -25601 -1186 -25567
rect -1220 -25669 -1186 -25635
rect -922 -25193 -888 -25159
rect -922 -25261 -888 -25227
rect -922 -25329 -888 -25295
rect -922 -25397 -888 -25363
rect -922 -25465 -888 -25431
rect -922 -25533 -888 -25499
rect -922 -25601 -888 -25567
rect -922 -25669 -888 -25635
rect -624 -25193 -590 -25159
rect -624 -25261 -590 -25227
rect -624 -25329 -590 -25295
rect -624 -25397 -590 -25363
rect -624 -25465 -590 -25431
rect -624 -25533 -590 -25499
rect -624 -25601 -590 -25567
rect -624 -25669 -590 -25635
rect -326 -25193 -292 -25159
rect -326 -25261 -292 -25227
rect -326 -25329 -292 -25295
rect -326 -25397 -292 -25363
rect -326 -25465 -292 -25431
rect -326 -25533 -292 -25499
rect -326 -25601 -292 -25567
rect -326 -25669 -292 -25635
rect -28 -25193 6 -25159
rect -28 -25261 6 -25227
rect -28 -25329 6 -25295
rect -28 -25397 6 -25363
rect -28 -25465 6 -25431
rect -28 -25533 6 -25499
rect -28 -25601 6 -25567
rect -28 -25669 6 -25635
rect 270 -25193 304 -25159
rect 270 -25261 304 -25227
rect 270 -25329 304 -25295
rect 270 -25397 304 -25363
rect 270 -25465 304 -25431
rect 270 -25533 304 -25499
rect 270 -25601 304 -25567
rect 270 -25669 304 -25635
rect 568 -25193 602 -25159
rect 568 -25261 602 -25227
rect 568 -25329 602 -25295
rect 568 -25397 602 -25363
rect 568 -25465 602 -25431
rect 568 -25533 602 -25499
rect 568 -25601 602 -25567
rect 568 -25669 602 -25635
rect 866 -25193 900 -25159
rect 866 -25261 900 -25227
rect 866 -25329 900 -25295
rect 866 -25397 900 -25363
rect 866 -25465 900 -25431
rect 866 -25533 900 -25499
rect 866 -25601 900 -25567
rect 866 -25669 900 -25635
rect 2580 -25363 2614 -25329
rect 2580 -25431 2614 -25397
rect 2580 -25499 2614 -25465
rect 2580 -25567 2614 -25533
rect 2580 -25635 2614 -25601
rect 2580 -25703 2614 -25669
rect 2580 -25771 2614 -25737
rect 2580 -25839 2614 -25805
rect 3598 -25363 3632 -25329
rect 3598 -25431 3632 -25397
rect 3598 -25499 3632 -25465
rect 3598 -25567 3632 -25533
rect 3598 -25635 3632 -25601
rect 3598 -25703 3632 -25669
rect 3598 -25771 3632 -25737
rect 3598 -25839 3632 -25805
rect 4616 -25363 4650 -25329
rect 4616 -25431 4650 -25397
rect 4616 -25499 4650 -25465
rect 4616 -25567 4650 -25533
rect 4616 -25635 4650 -25601
rect 4616 -25703 4650 -25669
rect 4616 -25771 4650 -25737
rect 4616 -25839 4650 -25805
rect 5634 -25363 5668 -25329
rect 5634 -25431 5668 -25397
rect 5634 -25499 5668 -25465
rect 5634 -25567 5668 -25533
rect 5634 -25635 5668 -25601
rect 5634 -25703 5668 -25669
rect 5634 -25771 5668 -25737
rect 5634 -25839 5668 -25805
rect 6652 -25363 6686 -25329
rect 6652 -25431 6686 -25397
rect 6652 -25499 6686 -25465
rect 6652 -25567 6686 -25533
rect 6652 -25635 6686 -25601
rect 6652 -25703 6686 -25669
rect 6652 -25771 6686 -25737
rect 6652 -25839 6686 -25805
rect 7670 -25363 7704 -25329
rect 7670 -25431 7704 -25397
rect 7670 -25499 7704 -25465
rect 7670 -25567 7704 -25533
rect 7670 -25635 7704 -25601
rect 7670 -25703 7704 -25669
rect 7670 -25771 7704 -25737
rect 7670 -25839 7704 -25805
rect 8688 -25363 8722 -25329
rect 8688 -25431 8722 -25397
rect 8688 -25499 8722 -25465
rect 8688 -25567 8722 -25533
rect 8688 -25635 8722 -25601
rect 8688 -25703 8722 -25669
rect 8688 -25771 8722 -25737
rect 8688 -25839 8722 -25805
rect 9706 -25363 9740 -25329
rect 9706 -25431 9740 -25397
rect 9706 -25499 9740 -25465
rect 9706 -25567 9740 -25533
rect 9706 -25635 9740 -25601
rect 9706 -25703 9740 -25669
rect 9706 -25771 9740 -25737
rect 9706 -25839 9740 -25805
rect 10724 -25363 10758 -25329
rect 10724 -25431 10758 -25397
rect 10724 -25499 10758 -25465
rect 10724 -25567 10758 -25533
rect 10724 -25635 10758 -25601
rect 10724 -25703 10758 -25669
rect 10724 -25771 10758 -25737
rect 10724 -25839 10758 -25805
rect 11742 -25363 11776 -25329
rect 11742 -25431 11776 -25397
rect 11742 -25499 11776 -25465
rect 11742 -25567 11776 -25533
rect 11742 -25635 11776 -25601
rect 11742 -25703 11776 -25669
rect 11742 -25771 11776 -25737
rect 11742 -25839 11776 -25805
rect 12760 -25363 12794 -25329
rect 12760 -25431 12794 -25397
rect 12760 -25499 12794 -25465
rect 12760 -25567 12794 -25533
rect 12760 -25635 12794 -25601
rect 12760 -25703 12794 -25669
rect 12760 -25771 12794 -25737
rect 12760 -25839 12794 -25805
rect 13778 -25363 13812 -25329
rect 13778 -25431 13812 -25397
rect 13778 -25499 13812 -25465
rect 13778 -25567 13812 -25533
rect 13778 -25635 13812 -25601
rect 13778 -25703 13812 -25669
rect 13778 -25771 13812 -25737
rect 13778 -25839 13812 -25805
rect 14796 -25363 14830 -25329
rect 14796 -25431 14830 -25397
rect 14796 -25499 14830 -25465
rect 14796 -25567 14830 -25533
rect 14796 -25635 14830 -25601
rect 14796 -25703 14830 -25669
rect 14796 -25771 14830 -25737
rect 14796 -25839 14830 -25805
rect 15814 -25363 15848 -25329
rect 15814 -25431 15848 -25397
rect 15814 -25499 15848 -25465
rect 15814 -25567 15848 -25533
rect 15814 -25635 15848 -25601
rect 15814 -25703 15848 -25669
rect 15814 -25771 15848 -25737
rect 15814 -25839 15848 -25805
rect 16832 -25363 16866 -25329
rect 16832 -25431 16866 -25397
rect 16832 -25499 16866 -25465
rect 16832 -25567 16866 -25533
rect 16832 -25635 16866 -25601
rect 16832 -25703 16866 -25669
rect 16832 -25771 16866 -25737
rect 16832 -25839 16866 -25805
rect 17850 -25363 17884 -25329
rect 17850 -25431 17884 -25397
rect 17850 -25499 17884 -25465
rect 17850 -25567 17884 -25533
rect 17850 -25635 17884 -25601
rect 17850 -25703 17884 -25669
rect 17850 -25771 17884 -25737
rect 17850 -25839 17884 -25805
rect 18868 -25363 18902 -25329
rect 18868 -25431 18902 -25397
rect 18868 -25499 18902 -25465
rect 18868 -25567 18902 -25533
rect 18868 -25635 18902 -25601
rect 18868 -25703 18902 -25669
rect 18868 -25771 18902 -25737
rect 18868 -25839 18902 -25805
rect 19886 -25363 19920 -25329
rect 19886 -25431 19920 -25397
rect 19886 -25499 19920 -25465
rect 19886 -25567 19920 -25533
rect 19886 -25635 19920 -25601
rect 19886 -25703 19920 -25669
rect 19886 -25771 19920 -25737
rect 19886 -25839 19920 -25805
rect 20904 -25363 20938 -25329
rect 20904 -25431 20938 -25397
rect 20904 -25499 20938 -25465
rect 20904 -25567 20938 -25533
rect 20904 -25635 20938 -25601
rect 20904 -25703 20938 -25669
rect 20904 -25771 20938 -25737
rect 20904 -25839 20938 -25805
rect 21922 -25363 21956 -25329
rect 21922 -25431 21956 -25397
rect 21922 -25499 21956 -25465
rect 21922 -25567 21956 -25533
rect 21922 -25635 21956 -25601
rect 21922 -25703 21956 -25669
rect 21922 -25771 21956 -25737
rect 21922 -25839 21956 -25805
rect 22940 -25363 22974 -25329
rect 22940 -25431 22974 -25397
rect 22940 -25499 22974 -25465
rect 22940 -25567 22974 -25533
rect 22940 -25635 22974 -25601
rect 22940 -25703 22974 -25669
rect 22940 -25771 22974 -25737
rect 22940 -25839 22974 -25805
<< pdiffc >>
rect 3626 -4737 3660 -4703
rect 3626 -4805 3660 -4771
rect 3626 -4873 3660 -4839
rect 3626 -4941 3660 -4907
rect 3626 -5009 3660 -4975
rect 3626 -5077 3660 -5043
rect 3844 -4737 3878 -4703
rect 3844 -4805 3878 -4771
rect 3844 -4873 3878 -4839
rect 3844 -4941 3878 -4907
rect 3844 -5009 3878 -4975
rect 3844 -5077 3878 -5043
rect 4062 -4737 4096 -4703
rect 4062 -4805 4096 -4771
rect 4062 -4873 4096 -4839
rect 4062 -4941 4096 -4907
rect 4062 -5009 4096 -4975
rect 4062 -5077 4096 -5043
rect 4280 -4737 4314 -4703
rect 4280 -4805 4314 -4771
rect 4280 -4873 4314 -4839
rect 4280 -4941 4314 -4907
rect 4280 -5009 4314 -4975
rect 4280 -5077 4314 -5043
rect 4498 -4737 4532 -4703
rect 4498 -4805 4532 -4771
rect 4498 -4873 4532 -4839
rect 4498 -4941 4532 -4907
rect 4498 -5009 4532 -4975
rect 4498 -5077 4532 -5043
rect 4716 -4737 4750 -4703
rect 4716 -4805 4750 -4771
rect 4716 -4873 4750 -4839
rect 4716 -4941 4750 -4907
rect 4716 -5009 4750 -4975
rect 4716 -5077 4750 -5043
rect 4934 -4737 4968 -4703
rect 4934 -4805 4968 -4771
rect 4934 -4873 4968 -4839
rect 4934 -4941 4968 -4907
rect 4934 -5009 4968 -4975
rect 4934 -5077 4968 -5043
rect 5152 -4737 5186 -4703
rect 5152 -4805 5186 -4771
rect 5152 -4873 5186 -4839
rect 5152 -4941 5186 -4907
rect 5152 -5009 5186 -4975
rect 5152 -5077 5186 -5043
rect 5370 -4737 5404 -4703
rect 5370 -4805 5404 -4771
rect 5370 -4873 5404 -4839
rect 5370 -4941 5404 -4907
rect 5370 -5009 5404 -4975
rect 5370 -5077 5404 -5043
rect 5588 -4737 5622 -4703
rect 5588 -4805 5622 -4771
rect 5588 -4873 5622 -4839
rect 5588 -4941 5622 -4907
rect 5588 -5009 5622 -4975
rect 5588 -5077 5622 -5043
rect 5806 -4737 5840 -4703
rect 5806 -4805 5840 -4771
rect 5806 -4873 5840 -4839
rect 5806 -4941 5840 -4907
rect 5806 -5009 5840 -4975
rect 5806 -5077 5840 -5043
rect 3626 -5675 3660 -5641
rect 3626 -5743 3660 -5709
rect 3626 -5811 3660 -5777
rect 3626 -5879 3660 -5845
rect 3626 -5947 3660 -5913
rect 3626 -6015 3660 -5981
rect 3844 -5675 3878 -5641
rect 3844 -5743 3878 -5709
rect 3844 -5811 3878 -5777
rect 3844 -5879 3878 -5845
rect 3844 -5947 3878 -5913
rect 3844 -6015 3878 -5981
rect 4062 -5675 4096 -5641
rect 4062 -5743 4096 -5709
rect 4062 -5811 4096 -5777
rect 4062 -5879 4096 -5845
rect 4062 -5947 4096 -5913
rect 4062 -6015 4096 -5981
rect 4280 -5675 4314 -5641
rect 4280 -5743 4314 -5709
rect 4280 -5811 4314 -5777
rect 4280 -5879 4314 -5845
rect 4280 -5947 4314 -5913
rect 4280 -6015 4314 -5981
rect 4498 -5675 4532 -5641
rect 4498 -5743 4532 -5709
rect 4498 -5811 4532 -5777
rect 4498 -5879 4532 -5845
rect 4498 -5947 4532 -5913
rect 4498 -6015 4532 -5981
rect 4716 -5675 4750 -5641
rect 4716 -5743 4750 -5709
rect 4716 -5811 4750 -5777
rect 4716 -5879 4750 -5845
rect 4716 -5947 4750 -5913
rect 4716 -6015 4750 -5981
rect 4934 -5675 4968 -5641
rect 4934 -5743 4968 -5709
rect 4934 -5811 4968 -5777
rect 4934 -5879 4968 -5845
rect 4934 -5947 4968 -5913
rect 4934 -6015 4968 -5981
rect 5152 -5675 5186 -5641
rect 5152 -5743 5186 -5709
rect 5152 -5811 5186 -5777
rect 5152 -5879 5186 -5845
rect 5152 -5947 5186 -5913
rect 5152 -6015 5186 -5981
rect 5370 -5675 5404 -5641
rect 5370 -5743 5404 -5709
rect 5370 -5811 5404 -5777
rect 5370 -5879 5404 -5845
rect 5370 -5947 5404 -5913
rect 5370 -6015 5404 -5981
rect 5588 -5675 5622 -5641
rect 5588 -5743 5622 -5709
rect 5588 -5811 5622 -5777
rect 5588 -5879 5622 -5845
rect 5588 -5947 5622 -5913
rect 5588 -6015 5622 -5981
rect 5806 -5675 5840 -5641
rect 5806 -5743 5840 -5709
rect 5806 -5811 5840 -5777
rect 5806 -5879 5840 -5845
rect 5806 -5947 5840 -5913
rect 5806 -6015 5840 -5981
rect 3626 -6613 3660 -6579
rect 3626 -6681 3660 -6647
rect 3626 -6749 3660 -6715
rect 3626 -6817 3660 -6783
rect 3626 -6885 3660 -6851
rect 3626 -6953 3660 -6919
rect 3844 -6613 3878 -6579
rect 3844 -6681 3878 -6647
rect 3844 -6749 3878 -6715
rect 3844 -6817 3878 -6783
rect 3844 -6885 3878 -6851
rect 3844 -6953 3878 -6919
rect 4062 -6613 4096 -6579
rect 4062 -6681 4096 -6647
rect 4062 -6749 4096 -6715
rect 4062 -6817 4096 -6783
rect 4062 -6885 4096 -6851
rect 4062 -6953 4096 -6919
rect 4280 -6613 4314 -6579
rect 4280 -6681 4314 -6647
rect 4280 -6749 4314 -6715
rect 4280 -6817 4314 -6783
rect 4280 -6885 4314 -6851
rect 4280 -6953 4314 -6919
rect 4498 -6613 4532 -6579
rect 4498 -6681 4532 -6647
rect 4498 -6749 4532 -6715
rect 4498 -6817 4532 -6783
rect 4498 -6885 4532 -6851
rect 4498 -6953 4532 -6919
rect 4716 -6613 4750 -6579
rect 4716 -6681 4750 -6647
rect 4716 -6749 4750 -6715
rect 4716 -6817 4750 -6783
rect 4716 -6885 4750 -6851
rect 4716 -6953 4750 -6919
rect 4934 -6613 4968 -6579
rect 4934 -6681 4968 -6647
rect 4934 -6749 4968 -6715
rect 4934 -6817 4968 -6783
rect 4934 -6885 4968 -6851
rect 4934 -6953 4968 -6919
rect 5152 -6613 5186 -6579
rect 5152 -6681 5186 -6647
rect 5152 -6749 5186 -6715
rect 5152 -6817 5186 -6783
rect 5152 -6885 5186 -6851
rect 5152 -6953 5186 -6919
rect 5370 -6613 5404 -6579
rect 5370 -6681 5404 -6647
rect 5370 -6749 5404 -6715
rect 5370 -6817 5404 -6783
rect 5370 -6885 5404 -6851
rect 5370 -6953 5404 -6919
rect 5588 -6613 5622 -6579
rect 5588 -6681 5622 -6647
rect 5588 -6749 5622 -6715
rect 5588 -6817 5622 -6783
rect 5588 -6885 5622 -6851
rect 5588 -6953 5622 -6919
rect 5806 -6613 5840 -6579
rect 5806 -6681 5840 -6647
rect 5806 -6749 5840 -6715
rect 5806 -6817 5840 -6783
rect 5806 -6885 5840 -6851
rect 5806 -6953 5840 -6919
rect 3626 -7551 3660 -7517
rect 3626 -7619 3660 -7585
rect 3626 -7687 3660 -7653
rect 3626 -7755 3660 -7721
rect 3626 -7823 3660 -7789
rect 3626 -7891 3660 -7857
rect 3844 -7551 3878 -7517
rect 3844 -7619 3878 -7585
rect 3844 -7687 3878 -7653
rect 3844 -7755 3878 -7721
rect 3844 -7823 3878 -7789
rect 3844 -7891 3878 -7857
rect 4062 -7551 4096 -7517
rect 4062 -7619 4096 -7585
rect 4062 -7687 4096 -7653
rect 4062 -7755 4096 -7721
rect 4062 -7823 4096 -7789
rect 4062 -7891 4096 -7857
rect 4280 -7551 4314 -7517
rect 4280 -7619 4314 -7585
rect 4280 -7687 4314 -7653
rect 4280 -7755 4314 -7721
rect 4280 -7823 4314 -7789
rect 4280 -7891 4314 -7857
rect 4498 -7551 4532 -7517
rect 4498 -7619 4532 -7585
rect 4498 -7687 4532 -7653
rect 4498 -7755 4532 -7721
rect 4498 -7823 4532 -7789
rect 4498 -7891 4532 -7857
rect 4716 -7551 4750 -7517
rect 4716 -7619 4750 -7585
rect 4716 -7687 4750 -7653
rect 4716 -7755 4750 -7721
rect 4716 -7823 4750 -7789
rect 4716 -7891 4750 -7857
rect 4934 -7551 4968 -7517
rect 4934 -7619 4968 -7585
rect 4934 -7687 4968 -7653
rect 4934 -7755 4968 -7721
rect 4934 -7823 4968 -7789
rect 4934 -7891 4968 -7857
rect 5152 -7551 5186 -7517
rect 5152 -7619 5186 -7585
rect 5152 -7687 5186 -7653
rect 5152 -7755 5186 -7721
rect 5152 -7823 5186 -7789
rect 5152 -7891 5186 -7857
rect 5370 -7551 5404 -7517
rect 5370 -7619 5404 -7585
rect 5370 -7687 5404 -7653
rect 5370 -7755 5404 -7721
rect 5370 -7823 5404 -7789
rect 5370 -7891 5404 -7857
rect 5588 -7551 5622 -7517
rect 5588 -7619 5622 -7585
rect 5588 -7687 5622 -7653
rect 5588 -7755 5622 -7721
rect 5588 -7823 5622 -7789
rect 5588 -7891 5622 -7857
rect 5806 -7551 5840 -7517
rect 5806 -7619 5840 -7585
rect 5806 -7687 5840 -7653
rect 5806 -7755 5840 -7721
rect 5806 -7823 5840 -7789
rect 5806 -7891 5840 -7857
<< psubdiff >>
rect -12322 -11211 24922 -11178
rect -12322 -11245 -12145 -11211
rect -12111 -11245 -12077 -11211
rect -12043 -11245 -12009 -11211
rect -11975 -11245 -11941 -11211
rect -11907 -11245 -11873 -11211
rect -11839 -11245 -11805 -11211
rect -11771 -11245 -11737 -11211
rect -11703 -11245 -11669 -11211
rect -11635 -11245 -11601 -11211
rect -11567 -11245 -11533 -11211
rect -11499 -11245 -11465 -11211
rect -11431 -11245 -11397 -11211
rect -11363 -11245 -11329 -11211
rect -11295 -11245 -11261 -11211
rect -11227 -11245 -11193 -11211
rect -11159 -11245 -11125 -11211
rect -11091 -11245 -11057 -11211
rect -11023 -11245 -10989 -11211
rect -10955 -11245 -10921 -11211
rect -10887 -11245 -10853 -11211
rect -10819 -11245 -10785 -11211
rect -10751 -11245 -10717 -11211
rect -10683 -11245 -10649 -11211
rect -10615 -11245 -10581 -11211
rect -10547 -11245 -10513 -11211
rect -10479 -11245 -10445 -11211
rect -10411 -11245 -10377 -11211
rect -10343 -11245 -10309 -11211
rect -10275 -11245 -10241 -11211
rect -10207 -11245 -10173 -11211
rect -10139 -11245 -10105 -11211
rect -10071 -11245 -10037 -11211
rect -10003 -11245 -9969 -11211
rect -9935 -11245 -9901 -11211
rect -9867 -11245 -9833 -11211
rect -9799 -11245 -9765 -11211
rect -9731 -11245 -9697 -11211
rect -9663 -11245 -9629 -11211
rect -9595 -11245 -9561 -11211
rect -9527 -11245 -9493 -11211
rect -9459 -11245 -9425 -11211
rect -9391 -11245 -9357 -11211
rect -9323 -11245 -9289 -11211
rect -9255 -11245 -9221 -11211
rect -9187 -11245 -9153 -11211
rect -9119 -11245 -9085 -11211
rect -9051 -11245 -9017 -11211
rect -8983 -11245 -8949 -11211
rect -8915 -11245 -8881 -11211
rect -8847 -11245 -8813 -11211
rect -8779 -11245 -8745 -11211
rect -8711 -11245 -8677 -11211
rect -8643 -11245 -8609 -11211
rect -8575 -11245 -8541 -11211
rect -8507 -11245 -8473 -11211
rect -8439 -11245 -8405 -11211
rect -8371 -11245 -8337 -11211
rect -8303 -11245 -8269 -11211
rect -8235 -11245 -8201 -11211
rect -8167 -11245 -8133 -11211
rect -8099 -11245 -8065 -11211
rect -8031 -11245 -7997 -11211
rect -7963 -11245 -7929 -11211
rect -7895 -11245 -7861 -11211
rect -7827 -11245 -7793 -11211
rect -7759 -11245 -7725 -11211
rect -7691 -11245 -7657 -11211
rect -7623 -11245 -7589 -11211
rect -7555 -11245 -7521 -11211
rect -7487 -11245 -7453 -11211
rect -7419 -11245 -7385 -11211
rect -7351 -11245 -7317 -11211
rect -7283 -11245 -7249 -11211
rect -7215 -11245 -7181 -11211
rect -7147 -11245 -7113 -11211
rect -7079 -11245 -7045 -11211
rect -7011 -11245 -6977 -11211
rect -6943 -11245 -6909 -11211
rect -6875 -11245 -6841 -11211
rect -6807 -11245 -6773 -11211
rect -6739 -11245 -6705 -11211
rect -6671 -11245 -6637 -11211
rect -6603 -11245 -6569 -11211
rect -6535 -11245 -6501 -11211
rect -6467 -11245 -6433 -11211
rect -6399 -11245 -6365 -11211
rect -6331 -11245 -6297 -11211
rect -6263 -11245 -6229 -11211
rect -6195 -11245 -6161 -11211
rect -6127 -11245 -6093 -11211
rect -6059 -11245 -6025 -11211
rect -5991 -11245 -5957 -11211
rect -5923 -11245 -5889 -11211
rect -5855 -11245 -5821 -11211
rect -5787 -11245 -5753 -11211
rect -5719 -11245 -5685 -11211
rect -5651 -11245 -5617 -11211
rect -5583 -11245 -5549 -11211
rect -5515 -11245 -5481 -11211
rect -5447 -11245 -5413 -11211
rect -5379 -11245 -5345 -11211
rect -5311 -11245 -5277 -11211
rect -5243 -11245 -5209 -11211
rect -5175 -11245 -5141 -11211
rect -5107 -11245 -5073 -11211
rect -5039 -11245 -5005 -11211
rect -4971 -11245 -4937 -11211
rect -4903 -11245 -4869 -11211
rect -4835 -11245 -4801 -11211
rect -4767 -11245 -4733 -11211
rect -4699 -11245 -4665 -11211
rect -4631 -11245 -4597 -11211
rect -4563 -11245 -4529 -11211
rect -4495 -11245 -4461 -11211
rect -4427 -11245 -4393 -11211
rect -4359 -11245 -4325 -11211
rect -4291 -11245 -4257 -11211
rect -4223 -11245 -4189 -11211
rect -4155 -11245 -4121 -11211
rect -4087 -11245 -4053 -11211
rect -4019 -11245 -3985 -11211
rect -3951 -11245 -3917 -11211
rect -3883 -11245 -3849 -11211
rect -3815 -11245 -3781 -11211
rect -3747 -11245 -3713 -11211
rect -3679 -11245 -3645 -11211
rect -3611 -11245 -3577 -11211
rect -3543 -11245 -3509 -11211
rect -3475 -11245 -3441 -11211
rect -3407 -11245 -3373 -11211
rect -3339 -11245 -3305 -11211
rect -3271 -11245 -3237 -11211
rect -3203 -11245 -3169 -11211
rect -3135 -11245 -3101 -11211
rect -3067 -11245 -3033 -11211
rect -2999 -11245 -2965 -11211
rect -2931 -11245 -2897 -11211
rect -2863 -11245 -2829 -11211
rect -2795 -11245 -2761 -11211
rect -2727 -11245 -2693 -11211
rect -2659 -11245 -2625 -11211
rect -2591 -11245 -2557 -11211
rect -2523 -11245 -2489 -11211
rect -2455 -11245 -2421 -11211
rect -2387 -11245 -2353 -11211
rect -2319 -11245 -2285 -11211
rect -2251 -11245 -2217 -11211
rect -2183 -11245 -2149 -11211
rect -2115 -11245 -2081 -11211
rect -2047 -11245 -2013 -11211
rect -1979 -11245 -1945 -11211
rect -1911 -11245 -1877 -11211
rect -1843 -11245 -1809 -11211
rect -1775 -11245 -1741 -11211
rect -1707 -11245 -1673 -11211
rect -1639 -11245 -1605 -11211
rect -1571 -11245 -1537 -11211
rect -1503 -11245 -1469 -11211
rect -1435 -11245 -1401 -11211
rect -1367 -11245 -1333 -11211
rect -1299 -11245 -1265 -11211
rect -1231 -11245 -1197 -11211
rect -1163 -11245 -1129 -11211
rect -1095 -11245 -1061 -11211
rect -1027 -11245 -993 -11211
rect -959 -11245 -925 -11211
rect -891 -11245 -857 -11211
rect -823 -11245 -789 -11211
rect -755 -11245 -721 -11211
rect -687 -11245 -653 -11211
rect -619 -11245 -585 -11211
rect -551 -11245 -517 -11211
rect -483 -11245 -449 -11211
rect -415 -11245 -381 -11211
rect -347 -11245 -313 -11211
rect -279 -11245 -245 -11211
rect -211 -11245 -177 -11211
rect -143 -11245 -109 -11211
rect -75 -11245 -41 -11211
rect -7 -11245 27 -11211
rect 61 -11245 95 -11211
rect 129 -11245 163 -11211
rect 197 -11245 231 -11211
rect 265 -11245 299 -11211
rect 333 -11245 367 -11211
rect 401 -11245 435 -11211
rect 469 -11245 503 -11211
rect 537 -11245 571 -11211
rect 605 -11245 639 -11211
rect 673 -11245 707 -11211
rect 741 -11245 775 -11211
rect 809 -11245 843 -11211
rect 877 -11245 911 -11211
rect 945 -11245 979 -11211
rect 1013 -11245 1047 -11211
rect 1081 -11245 1115 -11211
rect 1149 -11245 1183 -11211
rect 1217 -11245 1251 -11211
rect 1285 -11245 1319 -11211
rect 1353 -11245 1387 -11211
rect 1421 -11245 1455 -11211
rect 1489 -11245 1523 -11211
rect 1557 -11245 1591 -11211
rect 1625 -11245 1659 -11211
rect 1693 -11245 1727 -11211
rect 1761 -11245 1795 -11211
rect 1829 -11245 1863 -11211
rect 1897 -11245 1931 -11211
rect 1965 -11245 1999 -11211
rect 2033 -11245 2067 -11211
rect 2101 -11245 2135 -11211
rect 2169 -11245 2203 -11211
rect 2237 -11245 2271 -11211
rect 2305 -11245 2339 -11211
rect 2373 -11245 2407 -11211
rect 2441 -11245 2475 -11211
rect 2509 -11245 2543 -11211
rect 2577 -11245 2611 -11211
rect 2645 -11245 2679 -11211
rect 2713 -11245 2747 -11211
rect 2781 -11245 2815 -11211
rect 2849 -11245 2883 -11211
rect 2917 -11245 2951 -11211
rect 2985 -11245 3019 -11211
rect 3053 -11245 3087 -11211
rect 3121 -11245 3155 -11211
rect 3189 -11245 3223 -11211
rect 3257 -11245 3291 -11211
rect 3325 -11245 3359 -11211
rect 3393 -11245 3427 -11211
rect 3461 -11245 3495 -11211
rect 3529 -11245 3563 -11211
rect 3597 -11245 3631 -11211
rect 3665 -11245 3699 -11211
rect 3733 -11245 3767 -11211
rect 3801 -11245 3835 -11211
rect 3869 -11245 3903 -11211
rect 3937 -11245 3971 -11211
rect 4005 -11245 4039 -11211
rect 4073 -11245 4107 -11211
rect 4141 -11245 4175 -11211
rect 4209 -11245 4243 -11211
rect 4277 -11245 4311 -11211
rect 4345 -11245 4379 -11211
rect 4413 -11245 4447 -11211
rect 4481 -11245 4515 -11211
rect 4549 -11245 4583 -11211
rect 4617 -11245 4651 -11211
rect 4685 -11245 4719 -11211
rect 4753 -11245 4787 -11211
rect 4821 -11245 4855 -11211
rect 4889 -11245 4923 -11211
rect 4957 -11245 4991 -11211
rect 5025 -11245 5059 -11211
rect 5093 -11245 5127 -11211
rect 5161 -11245 5195 -11211
rect 5229 -11245 5263 -11211
rect 5297 -11245 5331 -11211
rect 5365 -11245 5399 -11211
rect 5433 -11245 5467 -11211
rect 5501 -11245 5535 -11211
rect 5569 -11245 5603 -11211
rect 5637 -11245 5671 -11211
rect 5705 -11245 5739 -11211
rect 5773 -11245 5807 -11211
rect 5841 -11245 5875 -11211
rect 5909 -11245 5943 -11211
rect 5977 -11245 6011 -11211
rect 6045 -11245 6079 -11211
rect 6113 -11245 6147 -11211
rect 6181 -11245 6215 -11211
rect 6249 -11245 6283 -11211
rect 6317 -11245 6351 -11211
rect 6385 -11245 6419 -11211
rect 6453 -11245 6487 -11211
rect 6521 -11245 6555 -11211
rect 6589 -11245 6623 -11211
rect 6657 -11245 6691 -11211
rect 6725 -11245 6759 -11211
rect 6793 -11245 6827 -11211
rect 6861 -11245 6895 -11211
rect 6929 -11245 6963 -11211
rect 6997 -11245 7031 -11211
rect 7065 -11245 7099 -11211
rect 7133 -11245 7167 -11211
rect 7201 -11245 7235 -11211
rect 7269 -11245 7303 -11211
rect 7337 -11245 7371 -11211
rect 7405 -11245 7439 -11211
rect 7473 -11245 7507 -11211
rect 7541 -11245 7575 -11211
rect 7609 -11245 7643 -11211
rect 7677 -11245 7711 -11211
rect 7745 -11245 7779 -11211
rect 7813 -11245 7847 -11211
rect 7881 -11245 7915 -11211
rect 7949 -11245 7983 -11211
rect 8017 -11245 8051 -11211
rect 8085 -11245 8119 -11211
rect 8153 -11245 8187 -11211
rect 8221 -11245 8255 -11211
rect 8289 -11245 8323 -11211
rect 8357 -11245 8391 -11211
rect 8425 -11245 8459 -11211
rect 8493 -11245 8527 -11211
rect 8561 -11245 8595 -11211
rect 8629 -11245 8663 -11211
rect 8697 -11245 8731 -11211
rect 8765 -11245 8799 -11211
rect 8833 -11245 8867 -11211
rect 8901 -11245 8935 -11211
rect 8969 -11245 9003 -11211
rect 9037 -11245 9071 -11211
rect 9105 -11245 9139 -11211
rect 9173 -11245 9207 -11211
rect 9241 -11245 9275 -11211
rect 9309 -11245 9343 -11211
rect 9377 -11245 9411 -11211
rect 9445 -11245 9479 -11211
rect 9513 -11245 9547 -11211
rect 9581 -11245 9615 -11211
rect 9649 -11245 9683 -11211
rect 9717 -11245 9751 -11211
rect 9785 -11245 9819 -11211
rect 9853 -11245 9887 -11211
rect 9921 -11245 9955 -11211
rect 9989 -11245 10023 -11211
rect 10057 -11245 10091 -11211
rect 10125 -11245 10159 -11211
rect 10193 -11245 10227 -11211
rect 10261 -11245 10295 -11211
rect 10329 -11245 10363 -11211
rect 10397 -11245 10431 -11211
rect 10465 -11245 10499 -11211
rect 10533 -11245 10567 -11211
rect 10601 -11245 10635 -11211
rect 10669 -11245 10703 -11211
rect 10737 -11245 10771 -11211
rect 10805 -11245 10839 -11211
rect 10873 -11245 10907 -11211
rect 10941 -11245 10975 -11211
rect 11009 -11245 11043 -11211
rect 11077 -11245 11111 -11211
rect 11145 -11245 11179 -11211
rect 11213 -11245 11247 -11211
rect 11281 -11245 11315 -11211
rect 11349 -11245 11383 -11211
rect 11417 -11245 11451 -11211
rect 11485 -11245 11519 -11211
rect 11553 -11245 11587 -11211
rect 11621 -11245 11655 -11211
rect 11689 -11245 11723 -11211
rect 11757 -11245 11791 -11211
rect 11825 -11245 11859 -11211
rect 11893 -11245 11927 -11211
rect 11961 -11245 11995 -11211
rect 12029 -11245 12063 -11211
rect 12097 -11245 12131 -11211
rect 12165 -11245 12199 -11211
rect 12233 -11245 12267 -11211
rect 12301 -11245 12335 -11211
rect 12369 -11245 12403 -11211
rect 12437 -11245 12471 -11211
rect 12505 -11245 12539 -11211
rect 12573 -11245 12607 -11211
rect 12641 -11245 12675 -11211
rect 12709 -11245 12743 -11211
rect 12777 -11245 12811 -11211
rect 12845 -11245 12879 -11211
rect 12913 -11245 12947 -11211
rect 12981 -11245 13015 -11211
rect 13049 -11245 13083 -11211
rect 13117 -11245 13151 -11211
rect 13185 -11245 13219 -11211
rect 13253 -11245 13287 -11211
rect 13321 -11245 13355 -11211
rect 13389 -11245 13423 -11211
rect 13457 -11245 13491 -11211
rect 13525 -11245 13559 -11211
rect 13593 -11245 13627 -11211
rect 13661 -11245 13695 -11211
rect 13729 -11245 13763 -11211
rect 13797 -11245 13831 -11211
rect 13865 -11245 13899 -11211
rect 13933 -11245 13967 -11211
rect 14001 -11245 14035 -11211
rect 14069 -11245 14103 -11211
rect 14137 -11245 14171 -11211
rect 14205 -11245 14239 -11211
rect 14273 -11245 14307 -11211
rect 14341 -11245 14375 -11211
rect 14409 -11245 14443 -11211
rect 14477 -11245 14511 -11211
rect 14545 -11245 14579 -11211
rect 14613 -11245 14647 -11211
rect 14681 -11245 14715 -11211
rect 14749 -11245 14783 -11211
rect 14817 -11245 14851 -11211
rect 14885 -11245 14919 -11211
rect 14953 -11245 14987 -11211
rect 15021 -11245 15055 -11211
rect 15089 -11245 15123 -11211
rect 15157 -11245 15191 -11211
rect 15225 -11245 15259 -11211
rect 15293 -11245 15327 -11211
rect 15361 -11245 15395 -11211
rect 15429 -11245 15463 -11211
rect 15497 -11245 15531 -11211
rect 15565 -11245 15599 -11211
rect 15633 -11245 15667 -11211
rect 15701 -11245 15735 -11211
rect 15769 -11245 15803 -11211
rect 15837 -11245 15871 -11211
rect 15905 -11245 15939 -11211
rect 15973 -11245 16007 -11211
rect 16041 -11245 16075 -11211
rect 16109 -11245 16143 -11211
rect 16177 -11245 16211 -11211
rect 16245 -11245 16279 -11211
rect 16313 -11245 16347 -11211
rect 16381 -11245 16415 -11211
rect 16449 -11245 16483 -11211
rect 16517 -11245 16551 -11211
rect 16585 -11245 16619 -11211
rect 16653 -11245 16687 -11211
rect 16721 -11245 16755 -11211
rect 16789 -11245 16823 -11211
rect 16857 -11245 16891 -11211
rect 16925 -11245 16959 -11211
rect 16993 -11245 17027 -11211
rect 17061 -11245 17095 -11211
rect 17129 -11245 17163 -11211
rect 17197 -11245 17231 -11211
rect 17265 -11245 17299 -11211
rect 17333 -11245 17367 -11211
rect 17401 -11245 17435 -11211
rect 17469 -11245 17503 -11211
rect 17537 -11245 17571 -11211
rect 17605 -11245 17639 -11211
rect 17673 -11245 17707 -11211
rect 17741 -11245 17775 -11211
rect 17809 -11245 17843 -11211
rect 17877 -11245 17911 -11211
rect 17945 -11245 17979 -11211
rect 18013 -11245 18047 -11211
rect 18081 -11245 18115 -11211
rect 18149 -11245 18183 -11211
rect 18217 -11245 18251 -11211
rect 18285 -11245 18319 -11211
rect 18353 -11245 18387 -11211
rect 18421 -11245 18455 -11211
rect 18489 -11245 18523 -11211
rect 18557 -11245 18591 -11211
rect 18625 -11245 18659 -11211
rect 18693 -11245 18727 -11211
rect 18761 -11245 18795 -11211
rect 18829 -11245 18863 -11211
rect 18897 -11245 18931 -11211
rect 18965 -11245 18999 -11211
rect 19033 -11245 19067 -11211
rect 19101 -11245 19135 -11211
rect 19169 -11245 19203 -11211
rect 19237 -11245 19271 -11211
rect 19305 -11245 19339 -11211
rect 19373 -11245 19407 -11211
rect 19441 -11245 19475 -11211
rect 19509 -11245 19543 -11211
rect 19577 -11245 19611 -11211
rect 19645 -11245 19679 -11211
rect 19713 -11245 19747 -11211
rect 19781 -11245 19815 -11211
rect 19849 -11245 19883 -11211
rect 19917 -11245 19951 -11211
rect 19985 -11245 20019 -11211
rect 20053 -11245 20087 -11211
rect 20121 -11245 20155 -11211
rect 20189 -11245 20223 -11211
rect 20257 -11245 20291 -11211
rect 20325 -11245 20359 -11211
rect 20393 -11245 20427 -11211
rect 20461 -11245 20495 -11211
rect 20529 -11245 20563 -11211
rect 20597 -11245 20631 -11211
rect 20665 -11245 20699 -11211
rect 20733 -11245 20767 -11211
rect 20801 -11245 20835 -11211
rect 20869 -11245 20903 -11211
rect 20937 -11245 20971 -11211
rect 21005 -11245 21039 -11211
rect 21073 -11245 21107 -11211
rect 21141 -11245 21175 -11211
rect 21209 -11245 21243 -11211
rect 21277 -11245 21311 -11211
rect 21345 -11245 21379 -11211
rect 21413 -11245 21447 -11211
rect 21481 -11245 21515 -11211
rect 21549 -11245 21583 -11211
rect 21617 -11245 21651 -11211
rect 21685 -11245 21719 -11211
rect 21753 -11245 21787 -11211
rect 21821 -11245 21855 -11211
rect 21889 -11245 21923 -11211
rect 21957 -11245 21991 -11211
rect 22025 -11245 22059 -11211
rect 22093 -11245 22127 -11211
rect 22161 -11245 22195 -11211
rect 22229 -11245 22263 -11211
rect 22297 -11245 22331 -11211
rect 22365 -11245 22399 -11211
rect 22433 -11245 22467 -11211
rect 22501 -11245 22535 -11211
rect 22569 -11245 22603 -11211
rect 22637 -11245 22671 -11211
rect 22705 -11245 22739 -11211
rect 22773 -11245 22807 -11211
rect 22841 -11245 22875 -11211
rect 22909 -11245 22943 -11211
rect 22977 -11245 23011 -11211
rect 23045 -11245 23079 -11211
rect 23113 -11245 23147 -11211
rect 23181 -11245 23215 -11211
rect 23249 -11245 23283 -11211
rect 23317 -11245 23351 -11211
rect 23385 -11245 23419 -11211
rect 23453 -11245 23487 -11211
rect 23521 -11245 23555 -11211
rect 23589 -11245 23623 -11211
rect 23657 -11245 23691 -11211
rect 23725 -11245 23759 -11211
rect 23793 -11245 23827 -11211
rect 23861 -11245 23895 -11211
rect 23929 -11245 23963 -11211
rect 23997 -11245 24031 -11211
rect 24065 -11245 24099 -11211
rect 24133 -11245 24167 -11211
rect 24201 -11245 24235 -11211
rect 24269 -11245 24303 -11211
rect 24337 -11245 24371 -11211
rect 24405 -11245 24439 -11211
rect 24473 -11245 24507 -11211
rect 24541 -11245 24575 -11211
rect 24609 -11245 24643 -11211
rect 24677 -11245 24711 -11211
rect 24745 -11245 24922 -11211
rect -12322 -11278 24922 -11245
rect -12322 -11363 -12222 -11278
rect -12322 -11397 -12289 -11363
rect -12255 -11397 -12222 -11363
rect -12322 -11431 -12222 -11397
rect -12322 -11465 -12289 -11431
rect -12255 -11465 -12222 -11431
rect -12322 -11499 -12222 -11465
rect -12322 -11533 -12289 -11499
rect -12255 -11533 -12222 -11499
rect -12322 -11567 -12222 -11533
rect -12322 -11601 -12289 -11567
rect -12255 -11601 -12222 -11567
rect -12322 -11635 -12222 -11601
rect 24822 -11363 24922 -11278
rect 24822 -11397 24855 -11363
rect 24889 -11397 24922 -11363
rect 24822 -11431 24922 -11397
rect 24822 -11465 24855 -11431
rect 24889 -11465 24922 -11431
rect 24822 -11499 24922 -11465
rect 24822 -11533 24855 -11499
rect 24889 -11533 24922 -11499
rect 24822 -11567 24922 -11533
rect 24822 -11601 24855 -11567
rect 24889 -11601 24922 -11567
rect -12322 -11669 -12289 -11635
rect -12255 -11669 -12222 -11635
rect -12322 -11703 -12222 -11669
rect -12322 -11737 -12289 -11703
rect -12255 -11737 -12222 -11703
rect 24822 -11635 24922 -11601
rect 24822 -11669 24855 -11635
rect 24889 -11669 24922 -11635
rect 24822 -11703 24922 -11669
rect -12322 -11771 -12222 -11737
rect -12322 -11805 -12289 -11771
rect -12255 -11805 -12222 -11771
rect -12322 -11839 -12222 -11805
rect -12322 -11873 -12289 -11839
rect -12255 -11873 -12222 -11839
rect -12322 -11907 -12222 -11873
rect -12322 -11941 -12289 -11907
rect -12255 -11941 -12222 -11907
rect -12322 -11975 -12222 -11941
rect -12322 -12009 -12289 -11975
rect -12255 -12009 -12222 -11975
rect -12322 -12043 -12222 -12009
rect -12322 -12077 -12289 -12043
rect -12255 -12077 -12222 -12043
rect -12322 -12111 -12222 -12077
rect -12322 -12145 -12289 -12111
rect -12255 -12145 -12222 -12111
rect -12322 -12179 -12222 -12145
rect -12322 -12213 -12289 -12179
rect -12255 -12213 -12222 -12179
rect -12322 -12247 -12222 -12213
rect -12322 -12281 -12289 -12247
rect -12255 -12281 -12222 -12247
rect -12322 -12315 -12222 -12281
rect -12322 -12349 -12289 -12315
rect -12255 -12349 -12222 -12315
rect 24822 -11737 24855 -11703
rect 24889 -11737 24922 -11703
rect 24822 -11771 24922 -11737
rect 24822 -11805 24855 -11771
rect 24889 -11805 24922 -11771
rect 24822 -11839 24922 -11805
rect 24822 -11873 24855 -11839
rect 24889 -11873 24922 -11839
rect 24822 -11907 24922 -11873
rect 24822 -11941 24855 -11907
rect 24889 -11941 24922 -11907
rect 24822 -11975 24922 -11941
rect 24822 -12009 24855 -11975
rect 24889 -12009 24922 -11975
rect 24822 -12043 24922 -12009
rect 24822 -12077 24855 -12043
rect 24889 -12077 24922 -12043
rect 24822 -12111 24922 -12077
rect 24822 -12145 24855 -12111
rect 24889 -12145 24922 -12111
rect 24822 -12179 24922 -12145
rect 24822 -12213 24855 -12179
rect 24889 -12213 24922 -12179
rect 24822 -12247 24922 -12213
rect 24822 -12281 24855 -12247
rect 24889 -12281 24922 -12247
rect 24822 -12315 24922 -12281
rect -12322 -12383 -12222 -12349
rect -12322 -12417 -12289 -12383
rect -12255 -12417 -12222 -12383
rect 24822 -12349 24855 -12315
rect 24889 -12349 24922 -12315
rect 24822 -12383 24922 -12349
rect -12322 -12451 -12222 -12417
rect 24822 -12417 24855 -12383
rect 24889 -12417 24922 -12383
rect -12322 -12485 -12289 -12451
rect -12255 -12485 -12222 -12451
rect -12322 -12519 -12222 -12485
rect 24822 -12451 24922 -12417
rect 24822 -12485 24855 -12451
rect 24889 -12485 24922 -12451
rect -12322 -12553 -12289 -12519
rect -12255 -12553 -12222 -12519
rect -12322 -12587 -12222 -12553
rect -12322 -12621 -12289 -12587
rect -12255 -12621 -12222 -12587
rect -12322 -12655 -12222 -12621
rect -12322 -12689 -12289 -12655
rect -12255 -12689 -12222 -12655
rect -12322 -12723 -12222 -12689
rect -12322 -12757 -12289 -12723
rect -12255 -12757 -12222 -12723
rect -12322 -12791 -12222 -12757
rect -12322 -12825 -12289 -12791
rect -12255 -12825 -12222 -12791
rect -12322 -12859 -12222 -12825
rect -12322 -12893 -12289 -12859
rect -12255 -12893 -12222 -12859
rect -12322 -12927 -12222 -12893
rect -12322 -12961 -12289 -12927
rect -12255 -12961 -12222 -12927
rect -12322 -12995 -12222 -12961
rect -12322 -13029 -12289 -12995
rect -12255 -13029 -12222 -12995
rect -12322 -13063 -12222 -13029
rect -12322 -13097 -12289 -13063
rect -12255 -13097 -12222 -13063
rect -12322 -13131 -12222 -13097
rect 24822 -12519 24922 -12485
rect 24822 -12553 24855 -12519
rect 24889 -12553 24922 -12519
rect 24822 -12587 24922 -12553
rect 24822 -12621 24855 -12587
rect 24889 -12621 24922 -12587
rect 24822 -12655 24922 -12621
rect 24822 -12689 24855 -12655
rect 24889 -12689 24922 -12655
rect 24822 -12723 24922 -12689
rect 24822 -12757 24855 -12723
rect 24889 -12757 24922 -12723
rect 24822 -12791 24922 -12757
rect 24822 -12825 24855 -12791
rect 24889 -12825 24922 -12791
rect 24822 -12859 24922 -12825
rect 24822 -12893 24855 -12859
rect 24889 -12893 24922 -12859
rect 24822 -12927 24922 -12893
rect -12322 -13165 -12289 -13131
rect -12255 -13165 -12222 -13131
rect -12322 -13199 -12222 -13165
rect -12322 -13233 -12289 -13199
rect -12255 -13233 -12222 -13199
rect -12322 -13267 -12222 -13233
rect -12322 -13301 -12289 -13267
rect -12255 -13301 -12222 -13267
rect -12322 -13335 -12222 -13301
rect -12322 -13369 -12289 -13335
rect -12255 -13369 -12222 -13335
rect -12322 -13403 -12222 -13369
rect -12322 -13437 -12289 -13403
rect -12255 -13437 -12222 -13403
rect -12322 -13471 -12222 -13437
rect -12322 -13505 -12289 -13471
rect -12255 -13505 -12222 -13471
rect -12322 -13539 -12222 -13505
rect -12322 -13573 -12289 -13539
rect -12255 -13573 -12222 -13539
rect -12322 -13607 -12222 -13573
rect -12322 -13641 -12289 -13607
rect -12255 -13641 -12222 -13607
rect -12322 -13675 -12222 -13641
rect -12322 -13709 -12289 -13675
rect -12255 -13709 -12222 -13675
rect -12322 -13743 -12222 -13709
rect -12322 -13777 -12289 -13743
rect -12255 -13777 -12222 -13743
rect -12322 -13811 -12222 -13777
rect -12322 -13845 -12289 -13811
rect -12255 -13845 -12222 -13811
rect -12322 -13879 -12222 -13845
rect -12322 -13913 -12289 -13879
rect -12255 -13913 -12222 -13879
rect -12322 -13947 -12222 -13913
rect 24822 -12961 24855 -12927
rect 24889 -12961 24922 -12927
rect 24822 -12995 24922 -12961
rect 24822 -13029 24855 -12995
rect 24889 -13029 24922 -12995
rect 24822 -13063 24922 -13029
rect 24822 -13097 24855 -13063
rect 24889 -13097 24922 -13063
rect 24822 -13131 24922 -13097
rect 24822 -13165 24855 -13131
rect 24889 -13165 24922 -13131
rect 24822 -13199 24922 -13165
rect 24822 -13233 24855 -13199
rect 24889 -13233 24922 -13199
rect 24822 -13267 24922 -13233
rect 24822 -13301 24855 -13267
rect 24889 -13301 24922 -13267
rect 24822 -13335 24922 -13301
rect 24822 -13369 24855 -13335
rect 24889 -13369 24922 -13335
rect 24822 -13403 24922 -13369
rect 24822 -13437 24855 -13403
rect 24889 -13437 24922 -13403
rect 24822 -13471 24922 -13437
rect 24822 -13505 24855 -13471
rect 24889 -13505 24922 -13471
rect 24822 -13539 24922 -13505
rect 24822 -13573 24855 -13539
rect 24889 -13573 24922 -13539
rect 24822 -13607 24922 -13573
rect 24822 -13641 24855 -13607
rect 24889 -13641 24922 -13607
rect 24822 -13675 24922 -13641
rect 24822 -13709 24855 -13675
rect 24889 -13709 24922 -13675
rect 24822 -13743 24922 -13709
rect 24822 -13777 24855 -13743
rect 24889 -13777 24922 -13743
rect 24822 -13811 24922 -13777
rect 24822 -13845 24855 -13811
rect 24889 -13845 24922 -13811
rect 24822 -13879 24922 -13845
rect 24822 -13913 24855 -13879
rect 24889 -13913 24922 -13879
rect -12322 -13981 -12289 -13947
rect -12255 -13981 -12222 -13947
rect -12322 -14015 -12222 -13981
rect -12322 -14049 -12289 -14015
rect -12255 -14049 -12222 -14015
rect 24822 -13947 24922 -13913
rect 24822 -13981 24855 -13947
rect 24889 -13981 24922 -13947
rect 24822 -14015 24922 -13981
rect -12322 -14083 -12222 -14049
rect 24822 -14049 24855 -14015
rect 24889 -14049 24922 -14015
rect -12322 -14117 -12289 -14083
rect -12255 -14117 -12222 -14083
rect -12322 -14151 -12222 -14117
rect 24822 -14083 24922 -14049
rect -12322 -14185 -12289 -14151
rect -12255 -14185 -12222 -14151
rect -12322 -14219 -12222 -14185
rect -12322 -14253 -12289 -14219
rect -12255 -14253 -12222 -14219
rect -12322 -14287 -12222 -14253
rect -12322 -14321 -12289 -14287
rect -12255 -14321 -12222 -14287
rect -12322 -14355 -12222 -14321
rect -12322 -14389 -12289 -14355
rect -12255 -14389 -12222 -14355
rect -12322 -14423 -12222 -14389
rect -12322 -14457 -12289 -14423
rect -12255 -14457 -12222 -14423
rect -12322 -14491 -12222 -14457
rect -12322 -14525 -12289 -14491
rect -12255 -14525 -12222 -14491
rect -12322 -14559 -12222 -14525
rect -12322 -14593 -12289 -14559
rect -12255 -14593 -12222 -14559
rect -12322 -14627 -12222 -14593
rect -12322 -14661 -12289 -14627
rect -12255 -14661 -12222 -14627
rect -12322 -14695 -12222 -14661
rect -12322 -14729 -12289 -14695
rect -12255 -14729 -12222 -14695
rect -12322 -14763 -12222 -14729
rect 24822 -14117 24855 -14083
rect 24889 -14117 24922 -14083
rect 24822 -14151 24922 -14117
rect -12322 -14797 -12289 -14763
rect -12255 -14797 -12222 -14763
rect -12322 -14831 -12222 -14797
rect -12322 -14865 -12289 -14831
rect -12255 -14865 -12222 -14831
rect 24822 -14185 24855 -14151
rect 24889 -14185 24922 -14151
rect 24822 -14219 24922 -14185
rect 24822 -14253 24855 -14219
rect 24889 -14253 24922 -14219
rect 24822 -14287 24922 -14253
rect 24822 -14321 24855 -14287
rect 24889 -14321 24922 -14287
rect 24822 -14355 24922 -14321
rect 24822 -14389 24855 -14355
rect 24889 -14389 24922 -14355
rect 24822 -14423 24922 -14389
rect 24822 -14457 24855 -14423
rect 24889 -14457 24922 -14423
rect 24822 -14491 24922 -14457
rect 24822 -14525 24855 -14491
rect 24889 -14525 24922 -14491
rect 24822 -14559 24922 -14525
rect 24822 -14593 24855 -14559
rect 24889 -14593 24922 -14559
rect 24822 -14627 24922 -14593
rect 24822 -14661 24855 -14627
rect 24889 -14661 24922 -14627
rect 24822 -14695 24922 -14661
rect 24822 -14729 24855 -14695
rect 24889 -14729 24922 -14695
rect 24822 -14763 24922 -14729
rect -12322 -14899 -12222 -14865
rect 24822 -14797 24855 -14763
rect 24889 -14797 24922 -14763
rect 24822 -14831 24922 -14797
rect 24822 -14865 24855 -14831
rect 24889 -14865 24922 -14831
rect -12322 -14933 -12289 -14899
rect -12255 -14933 -12222 -14899
rect -12322 -14967 -12222 -14933
rect 24822 -14899 24922 -14865
rect 24822 -14933 24855 -14899
rect 24889 -14933 24922 -14899
rect -12322 -15001 -12289 -14967
rect -12255 -15001 -12222 -14967
rect -12322 -15035 -12222 -15001
rect -12322 -15069 -12289 -15035
rect -12255 -15069 -12222 -15035
rect -12322 -15103 -12222 -15069
rect -12322 -15137 -12289 -15103
rect -12255 -15137 -12222 -15103
rect -12322 -15171 -12222 -15137
rect -12322 -15205 -12289 -15171
rect -12255 -15205 -12222 -15171
rect -12322 -15239 -12222 -15205
rect -12322 -15273 -12289 -15239
rect -12255 -15273 -12222 -15239
rect -12322 -15307 -12222 -15273
rect -12322 -15341 -12289 -15307
rect -12255 -15341 -12222 -15307
rect -12322 -15375 -12222 -15341
rect -12322 -15409 -12289 -15375
rect -12255 -15409 -12222 -15375
rect -12322 -15443 -12222 -15409
rect -12322 -15477 -12289 -15443
rect -12255 -15477 -12222 -15443
rect -12322 -15511 -12222 -15477
rect -12322 -15545 -12289 -15511
rect -12255 -15545 -12222 -15511
rect -12322 -15579 -12222 -15545
rect 24822 -14967 24922 -14933
rect 24822 -15001 24855 -14967
rect 24889 -15001 24922 -14967
rect 24822 -15035 24922 -15001
rect 24822 -15069 24855 -15035
rect 24889 -15069 24922 -15035
rect 24822 -15103 24922 -15069
rect 24822 -15137 24855 -15103
rect 24889 -15137 24922 -15103
rect 24822 -15171 24922 -15137
rect 24822 -15205 24855 -15171
rect 24889 -15205 24922 -15171
rect 24822 -15239 24922 -15205
rect 24822 -15273 24855 -15239
rect 24889 -15273 24922 -15239
rect 24822 -15307 24922 -15273
rect 24822 -15341 24855 -15307
rect 24889 -15341 24922 -15307
rect 24822 -15375 24922 -15341
rect 24822 -15409 24855 -15375
rect 24889 -15409 24922 -15375
rect -12322 -15613 -12289 -15579
rect -12255 -15613 -12222 -15579
rect -12322 -15647 -12222 -15613
rect -12322 -15681 -12289 -15647
rect -12255 -15681 -12222 -15647
rect -12322 -15715 -12222 -15681
rect -12322 -15749 -12289 -15715
rect -12255 -15749 -12222 -15715
rect -12322 -15783 -12222 -15749
rect -12322 -15817 -12289 -15783
rect -12255 -15817 -12222 -15783
rect -12322 -15851 -12222 -15817
rect -12322 -15885 -12289 -15851
rect -12255 -15885 -12222 -15851
rect -12322 -15919 -12222 -15885
rect -12322 -15953 -12289 -15919
rect -12255 -15953 -12222 -15919
rect -12322 -15987 -12222 -15953
rect -12322 -16021 -12289 -15987
rect -12255 -16021 -12222 -15987
rect -12322 -16055 -12222 -16021
rect -12322 -16089 -12289 -16055
rect -12255 -16089 -12222 -16055
rect -12322 -16123 -12222 -16089
rect -12322 -16157 -12289 -16123
rect -12255 -16157 -12222 -16123
rect -12322 -16191 -12222 -16157
rect -12322 -16225 -12289 -16191
rect -12255 -16225 -12222 -16191
rect -12322 -16259 -12222 -16225
rect -12322 -16293 -12289 -16259
rect -12255 -16293 -12222 -16259
rect -12322 -16327 -12222 -16293
rect -12322 -16361 -12289 -16327
rect -12255 -16361 -12222 -16327
rect -12322 -16395 -12222 -16361
rect 24822 -15443 24922 -15409
rect 24822 -15477 24855 -15443
rect 24889 -15477 24922 -15443
rect 24822 -15511 24922 -15477
rect 24822 -15545 24855 -15511
rect 24889 -15545 24922 -15511
rect 24822 -15579 24922 -15545
rect 24822 -15613 24855 -15579
rect 24889 -15613 24922 -15579
rect 24822 -15647 24922 -15613
rect 24822 -15681 24855 -15647
rect 24889 -15681 24922 -15647
rect 24822 -15715 24922 -15681
rect 24822 -15749 24855 -15715
rect 24889 -15749 24922 -15715
rect 24822 -15783 24922 -15749
rect 24822 -15817 24855 -15783
rect 24889 -15817 24922 -15783
rect 24822 -15851 24922 -15817
rect 24822 -15885 24855 -15851
rect 24889 -15885 24922 -15851
rect 24822 -15919 24922 -15885
rect 24822 -15953 24855 -15919
rect 24889 -15953 24922 -15919
rect 24822 -15987 24922 -15953
rect 24822 -16021 24855 -15987
rect 24889 -16021 24922 -15987
rect 24822 -16055 24922 -16021
rect 24822 -16089 24855 -16055
rect 24889 -16089 24922 -16055
rect 24822 -16123 24922 -16089
rect 24822 -16157 24855 -16123
rect 24889 -16157 24922 -16123
rect 24822 -16191 24922 -16157
rect 24822 -16225 24855 -16191
rect 24889 -16225 24922 -16191
rect 24822 -16259 24922 -16225
rect 24822 -16293 24855 -16259
rect 24889 -16293 24922 -16259
rect 24822 -16327 24922 -16293
rect 24822 -16361 24855 -16327
rect 24889 -16361 24922 -16327
rect -12322 -16429 -12289 -16395
rect -12255 -16429 -12222 -16395
rect -12322 -16463 -12222 -16429
rect -12322 -16497 -12289 -16463
rect -12255 -16497 -12222 -16463
rect 24822 -16395 24922 -16361
rect 24822 -16429 24855 -16395
rect 24889 -16429 24922 -16395
rect 24822 -16463 24922 -16429
rect -12322 -16531 -12222 -16497
rect 24822 -16497 24855 -16463
rect 24889 -16497 24922 -16463
rect -12322 -16565 -12289 -16531
rect -12255 -16565 -12222 -16531
rect -12322 -16599 -12222 -16565
rect -12322 -16633 -12289 -16599
rect -12255 -16633 -12222 -16599
rect 24822 -16531 24922 -16497
rect -12322 -16667 -12222 -16633
rect -12322 -16701 -12289 -16667
rect -12255 -16701 -12222 -16667
rect -12322 -16735 -12222 -16701
rect -12322 -16769 -12289 -16735
rect -12255 -16769 -12222 -16735
rect -12322 -16803 -12222 -16769
rect -12322 -16837 -12289 -16803
rect -12255 -16837 -12222 -16803
rect -12322 -16871 -12222 -16837
rect -12322 -16905 -12289 -16871
rect -12255 -16905 -12222 -16871
rect -12322 -16939 -12222 -16905
rect -12322 -16973 -12289 -16939
rect -12255 -16973 -12222 -16939
rect -12322 -17007 -12222 -16973
rect -12322 -17041 -12289 -17007
rect -12255 -17041 -12222 -17007
rect -12322 -17075 -12222 -17041
rect -12322 -17109 -12289 -17075
rect -12255 -17109 -12222 -17075
rect -12322 -17143 -12222 -17109
rect -12322 -17177 -12289 -17143
rect -12255 -17177 -12222 -17143
rect -12322 -17211 -12222 -17177
rect 24822 -16565 24855 -16531
rect 24889 -16565 24922 -16531
rect 24822 -16599 24922 -16565
rect 24822 -16633 24855 -16599
rect 24889 -16633 24922 -16599
rect -12322 -17245 -12289 -17211
rect -12255 -17245 -12222 -17211
rect -12322 -17279 -12222 -17245
rect -12322 -17313 -12289 -17279
rect -12255 -17313 -12222 -17279
rect 24822 -16667 24922 -16633
rect 24822 -16701 24855 -16667
rect 24889 -16701 24922 -16667
rect 24822 -16735 24922 -16701
rect 24822 -16769 24855 -16735
rect 24889 -16769 24922 -16735
rect 24822 -16803 24922 -16769
rect 24822 -16837 24855 -16803
rect 24889 -16837 24922 -16803
rect 24822 -16871 24922 -16837
rect 24822 -16905 24855 -16871
rect 24889 -16905 24922 -16871
rect 24822 -16939 24922 -16905
rect 24822 -16973 24855 -16939
rect 24889 -16973 24922 -16939
rect 24822 -17007 24922 -16973
rect 24822 -17041 24855 -17007
rect 24889 -17041 24922 -17007
rect 24822 -17075 24922 -17041
rect 24822 -17109 24855 -17075
rect 24889 -17109 24922 -17075
rect 24822 -17143 24922 -17109
rect 24822 -17177 24855 -17143
rect 24889 -17177 24922 -17143
rect 24822 -17211 24922 -17177
rect 24822 -17245 24855 -17211
rect 24889 -17245 24922 -17211
rect -12322 -17347 -12222 -17313
rect -12322 -17381 -12289 -17347
rect -12255 -17381 -12222 -17347
rect -12322 -17415 -12222 -17381
rect -12322 -17449 -12289 -17415
rect -12255 -17449 -12222 -17415
rect 24822 -17279 24922 -17245
rect 24822 -17313 24855 -17279
rect 24889 -17313 24922 -17279
rect 24822 -17347 24922 -17313
rect 24822 -17381 24855 -17347
rect 24889 -17381 24922 -17347
rect 24822 -17415 24922 -17381
rect -12322 -17483 -12222 -17449
rect -12322 -17517 -12289 -17483
rect -12255 -17517 -12222 -17483
rect -12322 -17551 -12222 -17517
rect -12322 -17585 -12289 -17551
rect -12255 -17585 -12222 -17551
rect -12322 -17619 -12222 -17585
rect -12322 -17653 -12289 -17619
rect -12255 -17653 -12222 -17619
rect -12322 -17687 -12222 -17653
rect -12322 -17721 -12289 -17687
rect -12255 -17721 -12222 -17687
rect -12322 -17755 -12222 -17721
rect -12322 -17789 -12289 -17755
rect -12255 -17789 -12222 -17755
rect -12322 -17823 -12222 -17789
rect -12322 -17857 -12289 -17823
rect -12255 -17857 -12222 -17823
rect -12322 -17891 -12222 -17857
rect -12322 -17925 -12289 -17891
rect -12255 -17925 -12222 -17891
rect -12322 -17959 -12222 -17925
rect -12322 -17993 -12289 -17959
rect -12255 -17993 -12222 -17959
rect -12322 -18027 -12222 -17993
rect 24822 -17449 24855 -17415
rect 24889 -17449 24922 -17415
rect 24822 -17483 24922 -17449
rect 24822 -17517 24855 -17483
rect 24889 -17517 24922 -17483
rect 24822 -17551 24922 -17517
rect 24822 -17585 24855 -17551
rect 24889 -17585 24922 -17551
rect 24822 -17619 24922 -17585
rect 24822 -17653 24855 -17619
rect 24889 -17653 24922 -17619
rect 24822 -17687 24922 -17653
rect 24822 -17721 24855 -17687
rect 24889 -17721 24922 -17687
rect 24822 -17755 24922 -17721
rect 24822 -17789 24855 -17755
rect 24889 -17789 24922 -17755
rect 24822 -17823 24922 -17789
rect 24822 -17857 24855 -17823
rect 24889 -17857 24922 -17823
rect -12322 -18061 -12289 -18027
rect -12255 -18061 -12222 -18027
rect -12322 -18095 -12222 -18061
rect -12322 -18129 -12289 -18095
rect -12255 -18129 -12222 -18095
rect -12322 -18163 -12222 -18129
rect -12322 -18197 -12289 -18163
rect -12255 -18197 -12222 -18163
rect -12322 -18231 -12222 -18197
rect -12322 -18265 -12289 -18231
rect -12255 -18265 -12222 -18231
rect -12322 -18299 -12222 -18265
rect -12322 -18333 -12289 -18299
rect -12255 -18333 -12222 -18299
rect -12322 -18367 -12222 -18333
rect -12322 -18401 -12289 -18367
rect -12255 -18401 -12222 -18367
rect -12322 -18435 -12222 -18401
rect -12322 -18469 -12289 -18435
rect -12255 -18469 -12222 -18435
rect -12322 -18503 -12222 -18469
rect -12322 -18537 -12289 -18503
rect -12255 -18537 -12222 -18503
rect -12322 -18571 -12222 -18537
rect -12322 -18605 -12289 -18571
rect -12255 -18605 -12222 -18571
rect -12322 -18639 -12222 -18605
rect -12322 -18673 -12289 -18639
rect -12255 -18673 -12222 -18639
rect -12322 -18707 -12222 -18673
rect -12322 -18741 -12289 -18707
rect -12255 -18741 -12222 -18707
rect -12322 -18775 -12222 -18741
rect -12322 -18809 -12289 -18775
rect -12255 -18809 -12222 -18775
rect -12322 -18843 -12222 -18809
rect 24822 -17891 24922 -17857
rect 24822 -17925 24855 -17891
rect 24889 -17925 24922 -17891
rect 24822 -17959 24922 -17925
rect 24822 -17993 24855 -17959
rect 24889 -17993 24922 -17959
rect 24822 -18027 24922 -17993
rect 24822 -18061 24855 -18027
rect 24889 -18061 24922 -18027
rect 24822 -18095 24922 -18061
rect 24822 -18129 24855 -18095
rect 24889 -18129 24922 -18095
rect 24822 -18163 24922 -18129
rect 24822 -18197 24855 -18163
rect 24889 -18197 24922 -18163
rect 24822 -18231 24922 -18197
rect 24822 -18265 24855 -18231
rect 24889 -18265 24922 -18231
rect 24822 -18299 24922 -18265
rect 24822 -18333 24855 -18299
rect 24889 -18333 24922 -18299
rect 24822 -18367 24922 -18333
rect 24822 -18401 24855 -18367
rect 24889 -18401 24922 -18367
rect 24822 -18435 24922 -18401
rect 24822 -18469 24855 -18435
rect 24889 -18469 24922 -18435
rect 24822 -18503 24922 -18469
rect 24822 -18537 24855 -18503
rect 24889 -18537 24922 -18503
rect 24822 -18571 24922 -18537
rect 24822 -18605 24855 -18571
rect 24889 -18605 24922 -18571
rect 24822 -18639 24922 -18605
rect 24822 -18673 24855 -18639
rect 24889 -18673 24922 -18639
rect 24822 -18707 24922 -18673
rect 24822 -18741 24855 -18707
rect 24889 -18741 24922 -18707
rect 24822 -18775 24922 -18741
rect 24822 -18809 24855 -18775
rect 24889 -18809 24922 -18775
rect -12322 -18877 -12289 -18843
rect -12255 -18877 -12222 -18843
rect -12322 -18911 -12222 -18877
rect -12322 -18945 -12289 -18911
rect -12255 -18945 -12222 -18911
rect 24822 -18843 24922 -18809
rect 24822 -18877 24855 -18843
rect 24889 -18877 24922 -18843
rect 24822 -18911 24922 -18877
rect -12322 -18979 -12222 -18945
rect -12322 -19013 -12289 -18979
rect -12255 -19013 -12222 -18979
rect -12322 -19047 -12222 -19013
rect 24822 -18945 24855 -18911
rect 24889 -18945 24922 -18911
rect 24822 -18979 24922 -18945
rect 24822 -19013 24855 -18979
rect 24889 -19013 24922 -18979
rect -12322 -19081 -12289 -19047
rect -12255 -19081 -12222 -19047
rect -12322 -19115 -12222 -19081
rect -12322 -19149 -12289 -19115
rect -12255 -19149 -12222 -19115
rect 24822 -19047 24922 -19013
rect 24822 -19081 24855 -19047
rect 24889 -19081 24922 -19047
rect 24822 -19115 24922 -19081
rect -12322 -19183 -12222 -19149
rect -12322 -19217 -12289 -19183
rect -12255 -19217 -12222 -19183
rect -12322 -19251 -12222 -19217
rect -12322 -19285 -12289 -19251
rect -12255 -19285 -12222 -19251
rect -12322 -19319 -12222 -19285
rect -12322 -19353 -12289 -19319
rect -12255 -19353 -12222 -19319
rect -12322 -19387 -12222 -19353
rect -12322 -19421 -12289 -19387
rect -12255 -19421 -12222 -19387
rect -12322 -19455 -12222 -19421
rect -12322 -19489 -12289 -19455
rect -12255 -19489 -12222 -19455
rect -12322 -19523 -12222 -19489
rect -12322 -19557 -12289 -19523
rect -12255 -19557 -12222 -19523
rect -12322 -19591 -12222 -19557
rect -12322 -19625 -12289 -19591
rect -12255 -19625 -12222 -19591
rect -12322 -19659 -12222 -19625
rect -12322 -19693 -12289 -19659
rect -12255 -19693 -12222 -19659
rect -12322 -19727 -12222 -19693
rect -12322 -19761 -12289 -19727
rect -12255 -19761 -12222 -19727
rect -12322 -19795 -12222 -19761
rect -12322 -19829 -12289 -19795
rect -12255 -19829 -12222 -19795
rect 24822 -19149 24855 -19115
rect 24889 -19149 24922 -19115
rect 24822 -19183 24922 -19149
rect 24822 -19217 24855 -19183
rect 24889 -19217 24922 -19183
rect 24822 -19251 24922 -19217
rect 24822 -19285 24855 -19251
rect 24889 -19285 24922 -19251
rect 24822 -19319 24922 -19285
rect 24822 -19353 24855 -19319
rect 24889 -19353 24922 -19319
rect 24822 -19387 24922 -19353
rect 24822 -19421 24855 -19387
rect 24889 -19421 24922 -19387
rect 24822 -19455 24922 -19421
rect 24822 -19489 24855 -19455
rect 24889 -19489 24922 -19455
rect 24822 -19523 24922 -19489
rect 24822 -19557 24855 -19523
rect 24889 -19557 24922 -19523
rect 24822 -19591 24922 -19557
rect 24822 -19625 24855 -19591
rect 24889 -19625 24922 -19591
rect 24822 -19659 24922 -19625
rect 24822 -19693 24855 -19659
rect 24889 -19693 24922 -19659
rect 24822 -19727 24922 -19693
rect 24822 -19761 24855 -19727
rect 24889 -19761 24922 -19727
rect 24822 -19795 24922 -19761
rect -12322 -19863 -12222 -19829
rect -12322 -19897 -12289 -19863
rect -12255 -19897 -12222 -19863
rect -12322 -19931 -12222 -19897
rect 24822 -19829 24855 -19795
rect 24889 -19829 24922 -19795
rect 24822 -19863 24922 -19829
rect 24822 -19897 24855 -19863
rect 24889 -19897 24922 -19863
rect -12322 -19965 -12289 -19931
rect -12255 -19965 -12222 -19931
rect -12322 -19999 -12222 -19965
rect -12322 -20033 -12289 -19999
rect -12255 -20033 -12222 -19999
rect -12322 -20067 -12222 -20033
rect -12322 -20101 -12289 -20067
rect -12255 -20101 -12222 -20067
rect -12322 -20135 -12222 -20101
rect -12322 -20169 -12289 -20135
rect -12255 -20169 -12222 -20135
rect -12322 -20203 -12222 -20169
rect -12322 -20237 -12289 -20203
rect -12255 -20237 -12222 -20203
rect -12322 -20271 -12222 -20237
rect 24822 -19931 24922 -19897
rect 24822 -19965 24855 -19931
rect 24889 -19965 24922 -19931
rect 24822 -19999 24922 -19965
rect 24822 -20033 24855 -19999
rect 24889 -20033 24922 -19999
rect 24822 -20067 24922 -20033
rect 24822 -20101 24855 -20067
rect 24889 -20101 24922 -20067
rect 24822 -20135 24922 -20101
rect 24822 -20169 24855 -20135
rect 24889 -20169 24922 -20135
rect 24822 -20203 24922 -20169
rect 24822 -20237 24855 -20203
rect 24889 -20237 24922 -20203
rect -12322 -20305 -12289 -20271
rect -12255 -20305 -12222 -20271
rect -12322 -20339 -12222 -20305
rect -12322 -20373 -12289 -20339
rect -12255 -20373 -12222 -20339
rect 24822 -20271 24922 -20237
rect 24822 -20305 24855 -20271
rect 24889 -20305 24922 -20271
rect 24822 -20339 24922 -20305
rect -12322 -20407 -12222 -20373
rect -12322 -20441 -12289 -20407
rect -12255 -20441 -12222 -20407
rect -12322 -20475 -12222 -20441
rect -12322 -20509 -12289 -20475
rect -12255 -20509 -12222 -20475
rect -12322 -20543 -12222 -20509
rect -12322 -20577 -12289 -20543
rect -12255 -20577 -12222 -20543
rect -12322 -20611 -12222 -20577
rect -12322 -20645 -12289 -20611
rect -12255 -20645 -12222 -20611
rect -12322 -20679 -12222 -20645
rect -12322 -20713 -12289 -20679
rect -12255 -20713 -12222 -20679
rect -12322 -20747 -12222 -20713
rect -12322 -20781 -12289 -20747
rect -12255 -20781 -12222 -20747
rect -12322 -20815 -12222 -20781
rect -12322 -20849 -12289 -20815
rect -12255 -20849 -12222 -20815
rect -12322 -20883 -12222 -20849
rect -12322 -20917 -12289 -20883
rect -12255 -20917 -12222 -20883
rect -12322 -20951 -12222 -20917
rect -12322 -20985 -12289 -20951
rect -12255 -20985 -12222 -20951
rect 24822 -20373 24855 -20339
rect 24889 -20373 24922 -20339
rect 24822 -20407 24922 -20373
rect 24822 -20441 24855 -20407
rect 24889 -20441 24922 -20407
rect 24822 -20475 24922 -20441
rect 24822 -20509 24855 -20475
rect 24889 -20509 24922 -20475
rect 24822 -20543 24922 -20509
rect 24822 -20577 24855 -20543
rect 24889 -20577 24922 -20543
rect 24822 -20611 24922 -20577
rect 24822 -20645 24855 -20611
rect 24889 -20645 24922 -20611
rect 24822 -20679 24922 -20645
rect 24822 -20713 24855 -20679
rect 24889 -20713 24922 -20679
rect 24822 -20747 24922 -20713
rect 24822 -20781 24855 -20747
rect 24889 -20781 24922 -20747
rect 24822 -20815 24922 -20781
rect 24822 -20849 24855 -20815
rect 24889 -20849 24922 -20815
rect 24822 -20883 24922 -20849
rect 24822 -20917 24855 -20883
rect 24889 -20917 24922 -20883
rect 24822 -20951 24922 -20917
rect -12322 -21019 -12222 -20985
rect -12322 -21053 -12289 -21019
rect -12255 -21053 -12222 -21019
rect 24822 -20985 24855 -20951
rect 24889 -20985 24922 -20951
rect 24822 -21019 24922 -20985
rect -12322 -21087 -12222 -21053
rect -12322 -21121 -12289 -21087
rect -12255 -21121 -12222 -21087
rect -12322 -21155 -12222 -21121
rect -12322 -21189 -12289 -21155
rect -12255 -21189 -12222 -21155
rect -12322 -21223 -12222 -21189
rect -12322 -21257 -12289 -21223
rect -12255 -21257 -12222 -21223
rect -12322 -21291 -12222 -21257
rect -12322 -21325 -12289 -21291
rect -12255 -21325 -12222 -21291
rect -12322 -21359 -12222 -21325
rect -12322 -21393 -12289 -21359
rect -12255 -21393 -12222 -21359
rect -12322 -21427 -12222 -21393
rect -12322 -21461 -12289 -21427
rect -12255 -21461 -12222 -21427
rect -12322 -21495 -12222 -21461
rect -12322 -21529 -12289 -21495
rect -12255 -21529 -12222 -21495
rect 24822 -21053 24855 -21019
rect 24889 -21053 24922 -21019
rect 24822 -21087 24922 -21053
rect 24822 -21121 24855 -21087
rect 24889 -21121 24922 -21087
rect 24822 -21155 24922 -21121
rect 24822 -21189 24855 -21155
rect 24889 -21189 24922 -21155
rect 24822 -21223 24922 -21189
rect 24822 -21257 24855 -21223
rect 24889 -21257 24922 -21223
rect 24822 -21291 24922 -21257
rect 24822 -21325 24855 -21291
rect 24889 -21325 24922 -21291
rect 24822 -21359 24922 -21325
rect 24822 -21393 24855 -21359
rect 24889 -21393 24922 -21359
rect 24822 -21427 24922 -21393
rect 24822 -21461 24855 -21427
rect 24889 -21461 24922 -21427
rect 24822 -21495 24922 -21461
rect -12322 -21563 -12222 -21529
rect -12322 -21597 -12289 -21563
rect -12255 -21597 -12222 -21563
rect 24822 -21529 24855 -21495
rect 24889 -21529 24922 -21495
rect 24822 -21563 24922 -21529
rect -12322 -21631 -12222 -21597
rect -12322 -21665 -12289 -21631
rect -12255 -21665 -12222 -21631
rect -12322 -21699 -12222 -21665
rect -12322 -21733 -12289 -21699
rect -12255 -21733 -12222 -21699
rect -12322 -21767 -12222 -21733
rect -12322 -21801 -12289 -21767
rect -12255 -21801 -12222 -21767
rect -12322 -21835 -12222 -21801
rect -12322 -21869 -12289 -21835
rect -12255 -21869 -12222 -21835
rect -12322 -21903 -12222 -21869
rect -12322 -21937 -12289 -21903
rect -12255 -21937 -12222 -21903
rect -12322 -21971 -12222 -21937
rect -12322 -22005 -12289 -21971
rect -12255 -22005 -12222 -21971
rect -12322 -22039 -12222 -22005
rect -12322 -22073 -12289 -22039
rect -12255 -22073 -12222 -22039
rect -12322 -22107 -12222 -22073
rect -12322 -22141 -12289 -22107
rect -12255 -22141 -12222 -22107
rect -12322 -22175 -12222 -22141
rect -12322 -22209 -12289 -22175
rect -12255 -22209 -12222 -22175
rect -12322 -22243 -12222 -22209
rect -12322 -22277 -12289 -22243
rect -12255 -22277 -12222 -22243
rect -12322 -22311 -12222 -22277
rect -12322 -22345 -12289 -22311
rect -12255 -22345 -12222 -22311
rect -12322 -22379 -12222 -22345
rect -12322 -22413 -12289 -22379
rect -12255 -22413 -12222 -22379
rect 24822 -21597 24855 -21563
rect 24889 -21597 24922 -21563
rect 24822 -21631 24922 -21597
rect 24822 -21665 24855 -21631
rect 24889 -21665 24922 -21631
rect 24822 -21699 24922 -21665
rect 24822 -21733 24855 -21699
rect 24889 -21733 24922 -21699
rect 24822 -21767 24922 -21733
rect 24822 -21801 24855 -21767
rect 24889 -21801 24922 -21767
rect 24822 -21835 24922 -21801
rect 24822 -21869 24855 -21835
rect 24889 -21869 24922 -21835
rect 24822 -21903 24922 -21869
rect 24822 -21937 24855 -21903
rect 24889 -21937 24922 -21903
rect 24822 -21971 24922 -21937
rect 24822 -22005 24855 -21971
rect 24889 -22005 24922 -21971
rect 24822 -22039 24922 -22005
rect 24822 -22073 24855 -22039
rect 24889 -22073 24922 -22039
rect 24822 -22107 24922 -22073
rect 24822 -22141 24855 -22107
rect 24889 -22141 24922 -22107
rect 24822 -22175 24922 -22141
rect 24822 -22209 24855 -22175
rect 24889 -22209 24922 -22175
rect 24822 -22243 24922 -22209
rect 24822 -22277 24855 -22243
rect 24889 -22277 24922 -22243
rect 24822 -22311 24922 -22277
rect 24822 -22345 24855 -22311
rect 24889 -22345 24922 -22311
rect 24822 -22379 24922 -22345
rect -12322 -22447 -12222 -22413
rect -12322 -22481 -12289 -22447
rect -12255 -22481 -12222 -22447
rect 24822 -22413 24855 -22379
rect 24889 -22413 24922 -22379
rect 24822 -22447 24922 -22413
rect -12322 -22515 -12222 -22481
rect -12322 -22549 -12289 -22515
rect -12255 -22549 -12222 -22515
rect -12322 -22583 -12222 -22549
rect -12322 -22617 -12289 -22583
rect -12255 -22617 -12222 -22583
rect -12322 -22651 -12222 -22617
rect -12322 -22685 -12289 -22651
rect -12255 -22685 -12222 -22651
rect -12322 -22719 -12222 -22685
rect -12322 -22753 -12289 -22719
rect -12255 -22753 -12222 -22719
rect 24822 -22481 24855 -22447
rect 24889 -22481 24922 -22447
rect 24822 -22515 24922 -22481
rect 24822 -22549 24855 -22515
rect 24889 -22549 24922 -22515
rect 24822 -22583 24922 -22549
rect 24822 -22617 24855 -22583
rect 24889 -22617 24922 -22583
rect 24822 -22651 24922 -22617
rect 24822 -22685 24855 -22651
rect 24889 -22685 24922 -22651
rect 24822 -22719 24922 -22685
rect -12322 -22787 -12222 -22753
rect -12322 -22821 -12289 -22787
rect -12255 -22821 -12222 -22787
rect -12322 -22855 -12222 -22821
rect -12322 -22889 -12289 -22855
rect -12255 -22889 -12222 -22855
rect -12322 -22923 -12222 -22889
rect 24822 -22753 24855 -22719
rect 24889 -22753 24922 -22719
rect 24822 -22787 24922 -22753
rect -12322 -22957 -12289 -22923
rect -12255 -22957 -12222 -22923
rect -12322 -22991 -12222 -22957
rect -12322 -23025 -12289 -22991
rect -12255 -23025 -12222 -22991
rect -12322 -23059 -12222 -23025
rect -12322 -23093 -12289 -23059
rect -12255 -23093 -12222 -23059
rect -12322 -23127 -12222 -23093
rect -12322 -23161 -12289 -23127
rect -12255 -23161 -12222 -23127
rect -12322 -23195 -12222 -23161
rect -12322 -23229 -12289 -23195
rect -12255 -23229 -12222 -23195
rect -12322 -23263 -12222 -23229
rect -12322 -23297 -12289 -23263
rect -12255 -23297 -12222 -23263
rect -12322 -23331 -12222 -23297
rect -12322 -23365 -12289 -23331
rect -12255 -23365 -12222 -23331
rect -12322 -23399 -12222 -23365
rect -12322 -23433 -12289 -23399
rect -12255 -23433 -12222 -23399
rect -12322 -23467 -12222 -23433
rect -12322 -23501 -12289 -23467
rect -12255 -23501 -12222 -23467
rect 24822 -22821 24855 -22787
rect 24889 -22821 24922 -22787
rect 24822 -22855 24922 -22821
rect 24822 -22889 24855 -22855
rect 24889 -22889 24922 -22855
rect 24822 -22923 24922 -22889
rect 24822 -22957 24855 -22923
rect 24889 -22957 24922 -22923
rect 24822 -22991 24922 -22957
rect 24822 -23025 24855 -22991
rect 24889 -23025 24922 -22991
rect 24822 -23059 24922 -23025
rect 24822 -23093 24855 -23059
rect 24889 -23093 24922 -23059
rect 24822 -23127 24922 -23093
rect 24822 -23161 24855 -23127
rect 24889 -23161 24922 -23127
rect 24822 -23195 24922 -23161
rect 24822 -23229 24855 -23195
rect 24889 -23229 24922 -23195
rect 24822 -23263 24922 -23229
rect 24822 -23297 24855 -23263
rect 24889 -23297 24922 -23263
rect 24822 -23331 24922 -23297
rect 24822 -23365 24855 -23331
rect 24889 -23365 24922 -23331
rect 24822 -23399 24922 -23365
rect -12322 -23535 -12222 -23501
rect -12322 -23569 -12289 -23535
rect -12255 -23569 -12222 -23535
rect -12322 -23603 -12222 -23569
rect 24822 -23433 24855 -23399
rect 24889 -23433 24922 -23399
rect 24822 -23467 24922 -23433
rect 24822 -23501 24855 -23467
rect 24889 -23501 24922 -23467
rect 24822 -23535 24922 -23501
rect 24822 -23569 24855 -23535
rect 24889 -23569 24922 -23535
rect -12322 -23637 -12289 -23603
rect -12255 -23637 -12222 -23603
rect -12322 -23671 -12222 -23637
rect -12322 -23705 -12289 -23671
rect -12255 -23705 -12222 -23671
rect -12322 -23739 -12222 -23705
rect -12322 -23773 -12289 -23739
rect -12255 -23773 -12222 -23739
rect -12322 -23807 -12222 -23773
rect -12322 -23841 -12289 -23807
rect -12255 -23841 -12222 -23807
rect -12322 -23875 -12222 -23841
rect -12322 -23909 -12289 -23875
rect -12255 -23909 -12222 -23875
rect -12322 -23943 -12222 -23909
rect 24822 -23603 24922 -23569
rect 24822 -23637 24855 -23603
rect 24889 -23637 24922 -23603
rect 24822 -23671 24922 -23637
rect 24822 -23705 24855 -23671
rect 24889 -23705 24922 -23671
rect 24822 -23739 24922 -23705
rect 24822 -23773 24855 -23739
rect 24889 -23773 24922 -23739
rect 24822 -23807 24922 -23773
rect 24822 -23841 24855 -23807
rect 24889 -23841 24922 -23807
rect 24822 -23875 24922 -23841
rect 24822 -23909 24855 -23875
rect 24889 -23909 24922 -23875
rect -12322 -23977 -12289 -23943
rect -12255 -23977 -12222 -23943
rect -12322 -24011 -12222 -23977
rect 24822 -23943 24922 -23909
rect -12322 -24045 -12289 -24011
rect -12255 -24045 -12222 -24011
rect -12322 -24079 -12222 -24045
rect -12322 -24113 -12289 -24079
rect -12255 -24113 -12222 -24079
rect -12322 -24147 -12222 -24113
rect -12322 -24181 -12289 -24147
rect -12255 -24181 -12222 -24147
rect -12322 -24215 -12222 -24181
rect -12322 -24249 -12289 -24215
rect -12255 -24249 -12222 -24215
rect -12322 -24283 -12222 -24249
rect -12322 -24317 -12289 -24283
rect -12255 -24317 -12222 -24283
rect -12322 -24351 -12222 -24317
rect -12322 -24385 -12289 -24351
rect -12255 -24385 -12222 -24351
rect -12322 -24419 -12222 -24385
rect -12322 -24453 -12289 -24419
rect -12255 -24453 -12222 -24419
rect -12322 -24487 -12222 -24453
rect -12322 -24521 -12289 -24487
rect -12255 -24521 -12222 -24487
rect -12322 -24555 -12222 -24521
rect -12322 -24589 -12289 -24555
rect -12255 -24589 -12222 -24555
rect -12322 -24623 -12222 -24589
rect 24822 -23977 24855 -23943
rect 24889 -23977 24922 -23943
rect 24822 -24011 24922 -23977
rect 24822 -24045 24855 -24011
rect 24889 -24045 24922 -24011
rect -12322 -24657 -12289 -24623
rect -12255 -24657 -12222 -24623
rect -12322 -24691 -12222 -24657
rect -12322 -24725 -12289 -24691
rect -12255 -24725 -12222 -24691
rect 24822 -24079 24922 -24045
rect 24822 -24113 24855 -24079
rect 24889 -24113 24922 -24079
rect 24822 -24147 24922 -24113
rect 24822 -24181 24855 -24147
rect 24889 -24181 24922 -24147
rect 24822 -24215 24922 -24181
rect 24822 -24249 24855 -24215
rect 24889 -24249 24922 -24215
rect 24822 -24283 24922 -24249
rect 24822 -24317 24855 -24283
rect 24889 -24317 24922 -24283
rect 24822 -24351 24922 -24317
rect 24822 -24385 24855 -24351
rect 24889 -24385 24922 -24351
rect 24822 -24419 24922 -24385
rect 24822 -24453 24855 -24419
rect 24889 -24453 24922 -24419
rect 24822 -24487 24922 -24453
rect 24822 -24521 24855 -24487
rect 24889 -24521 24922 -24487
rect 24822 -24555 24922 -24521
rect 24822 -24589 24855 -24555
rect 24889 -24589 24922 -24555
rect 24822 -24623 24922 -24589
rect -12322 -24759 -12222 -24725
rect 24822 -24657 24855 -24623
rect 24889 -24657 24922 -24623
rect 24822 -24691 24922 -24657
rect 24822 -24725 24855 -24691
rect 24889 -24725 24922 -24691
rect -12322 -24793 -12289 -24759
rect -12255 -24793 -12222 -24759
rect -12322 -24827 -12222 -24793
rect -12322 -24861 -12289 -24827
rect -12255 -24861 -12222 -24827
rect -12322 -24895 -12222 -24861
rect -12322 -24929 -12289 -24895
rect -12255 -24929 -12222 -24895
rect -12322 -24963 -12222 -24929
rect -12322 -24997 -12289 -24963
rect -12255 -24997 -12222 -24963
rect -12322 -25031 -12222 -24997
rect 24822 -24759 24922 -24725
rect 24822 -24793 24855 -24759
rect 24889 -24793 24922 -24759
rect 24822 -24827 24922 -24793
rect 24822 -24861 24855 -24827
rect 24889 -24861 24922 -24827
rect 24822 -24895 24922 -24861
rect 24822 -24929 24855 -24895
rect 24889 -24929 24922 -24895
rect 24822 -24963 24922 -24929
rect 24822 -24997 24855 -24963
rect 24889 -24997 24922 -24963
rect -12322 -25065 -12289 -25031
rect -12255 -25065 -12222 -25031
rect -12322 -25099 -12222 -25065
rect -12322 -25133 -12289 -25099
rect -12255 -25133 -12222 -25099
rect 24822 -25031 24922 -24997
rect 24822 -25065 24855 -25031
rect 24889 -25065 24922 -25031
rect 24822 -25099 24922 -25065
rect -12322 -25167 -12222 -25133
rect -12322 -25201 -12289 -25167
rect -12255 -25201 -12222 -25167
rect -12322 -25235 -12222 -25201
rect -12322 -25269 -12289 -25235
rect -12255 -25269 -12222 -25235
rect -12322 -25303 -12222 -25269
rect -12322 -25337 -12289 -25303
rect -12255 -25337 -12222 -25303
rect -12322 -25371 -12222 -25337
rect -12322 -25405 -12289 -25371
rect -12255 -25405 -12222 -25371
rect -12322 -25439 -12222 -25405
rect -12322 -25473 -12289 -25439
rect -12255 -25473 -12222 -25439
rect -12322 -25507 -12222 -25473
rect -12322 -25541 -12289 -25507
rect -12255 -25541 -12222 -25507
rect -12322 -25575 -12222 -25541
rect -12322 -25609 -12289 -25575
rect -12255 -25609 -12222 -25575
rect -12322 -25643 -12222 -25609
rect -12322 -25677 -12289 -25643
rect -12255 -25677 -12222 -25643
rect -12322 -25711 -12222 -25677
rect -12322 -25745 -12289 -25711
rect -12255 -25745 -12222 -25711
rect 24822 -25133 24855 -25099
rect 24889 -25133 24922 -25099
rect 24822 -25167 24922 -25133
rect 24822 -25201 24855 -25167
rect 24889 -25201 24922 -25167
rect 24822 -25235 24922 -25201
rect 24822 -25269 24855 -25235
rect 24889 -25269 24922 -25235
rect -12322 -25779 -12222 -25745
rect -12322 -25813 -12289 -25779
rect -12255 -25813 -12222 -25779
rect -12322 -25847 -12222 -25813
rect -12322 -25881 -12289 -25847
rect -12255 -25881 -12222 -25847
rect -12322 -25915 -12222 -25881
rect 24822 -25303 24922 -25269
rect 24822 -25337 24855 -25303
rect 24889 -25337 24922 -25303
rect 24822 -25371 24922 -25337
rect 24822 -25405 24855 -25371
rect 24889 -25405 24922 -25371
rect 24822 -25439 24922 -25405
rect 24822 -25473 24855 -25439
rect 24889 -25473 24922 -25439
rect 24822 -25507 24922 -25473
rect 24822 -25541 24855 -25507
rect 24889 -25541 24922 -25507
rect 24822 -25575 24922 -25541
rect 24822 -25609 24855 -25575
rect 24889 -25609 24922 -25575
rect 24822 -25643 24922 -25609
rect 24822 -25677 24855 -25643
rect 24889 -25677 24922 -25643
rect 24822 -25711 24922 -25677
rect 24822 -25745 24855 -25711
rect 24889 -25745 24922 -25711
rect 24822 -25779 24922 -25745
rect 24822 -25813 24855 -25779
rect 24889 -25813 24922 -25779
rect 24822 -25847 24922 -25813
rect 24822 -25881 24855 -25847
rect 24889 -25881 24922 -25847
rect -12322 -25949 -12289 -25915
rect -12255 -25949 -12222 -25915
rect -12322 -25983 -12222 -25949
rect 24822 -25915 24922 -25881
rect 24822 -25949 24855 -25915
rect 24889 -25949 24922 -25915
rect -12322 -26017 -12289 -25983
rect -12255 -26017 -12222 -25983
rect -12322 -26051 -12222 -26017
rect -12322 -26085 -12289 -26051
rect -12255 -26085 -12222 -26051
rect -12322 -26119 -12222 -26085
rect -12322 -26153 -12289 -26119
rect -12255 -26153 -12222 -26119
rect -12322 -26187 -12222 -26153
rect -12322 -26221 -12289 -26187
rect -12255 -26221 -12222 -26187
rect -12322 -26255 -12222 -26221
rect -12322 -26289 -12289 -26255
rect -12255 -26289 -12222 -26255
rect -12322 -26323 -12222 -26289
rect -12322 -26357 -12289 -26323
rect -12255 -26357 -12222 -26323
rect -12322 -26391 -12222 -26357
rect -12322 -26425 -12289 -26391
rect -12255 -26425 -12222 -26391
rect -12322 -26459 -12222 -26425
rect -12322 -26493 -12289 -26459
rect -12255 -26493 -12222 -26459
rect -12322 -26527 -12222 -26493
rect -12322 -26561 -12289 -26527
rect -12255 -26561 -12222 -26527
rect -12322 -26595 -12222 -26561
rect -12322 -26629 -12289 -26595
rect -12255 -26629 -12222 -26595
rect -12322 -26663 -12222 -26629
rect -12322 -26697 -12289 -26663
rect -12255 -26697 -12222 -26663
rect -12322 -26731 -12222 -26697
rect -12322 -26765 -12289 -26731
rect -12255 -26765 -12222 -26731
rect -12322 -26799 -12222 -26765
rect -12322 -26833 -12289 -26799
rect -12255 -26833 -12222 -26799
rect -12322 -26867 -12222 -26833
rect -12322 -26901 -12289 -26867
rect -12255 -26901 -12222 -26867
rect -12322 -26935 -12222 -26901
rect -12322 -26969 -12289 -26935
rect -12255 -26969 -12222 -26935
rect -12322 -27003 -12222 -26969
rect -12322 -27037 -12289 -27003
rect -12255 -27037 -12222 -27003
rect -12322 -27122 -12222 -27037
rect 24822 -25983 24922 -25949
rect 24822 -26017 24855 -25983
rect 24889 -26017 24922 -25983
rect 24822 -26051 24922 -26017
rect 24822 -26085 24855 -26051
rect 24889 -26085 24922 -26051
rect 24822 -26119 24922 -26085
rect 24822 -26153 24855 -26119
rect 24889 -26153 24922 -26119
rect 24822 -26187 24922 -26153
rect 24822 -26221 24855 -26187
rect 24889 -26221 24922 -26187
rect 24822 -26255 24922 -26221
rect 24822 -26289 24855 -26255
rect 24889 -26289 24922 -26255
rect 24822 -26323 24922 -26289
rect 24822 -26357 24855 -26323
rect 24889 -26357 24922 -26323
rect 24822 -26391 24922 -26357
rect 24822 -26425 24855 -26391
rect 24889 -26425 24922 -26391
rect 24822 -26459 24922 -26425
rect 24822 -26493 24855 -26459
rect 24889 -26493 24922 -26459
rect 24822 -26527 24922 -26493
rect 24822 -26561 24855 -26527
rect 24889 -26561 24922 -26527
rect 24822 -26595 24922 -26561
rect 24822 -26629 24855 -26595
rect 24889 -26629 24922 -26595
rect 24822 -26663 24922 -26629
rect 24822 -26697 24855 -26663
rect 24889 -26697 24922 -26663
rect 24822 -26731 24922 -26697
rect 24822 -26765 24855 -26731
rect 24889 -26765 24922 -26731
rect 24822 -26799 24922 -26765
rect 24822 -26833 24855 -26799
rect 24889 -26833 24922 -26799
rect 24822 -26867 24922 -26833
rect 24822 -26901 24855 -26867
rect 24889 -26901 24922 -26867
rect 24822 -26935 24922 -26901
rect 24822 -26969 24855 -26935
rect 24889 -26969 24922 -26935
rect 24822 -27003 24922 -26969
rect 24822 -27037 24855 -27003
rect 24889 -27037 24922 -27003
rect 24822 -27122 24922 -27037
rect -12322 -27155 24922 -27122
rect -12322 -27189 -12145 -27155
rect -12111 -27189 -12077 -27155
rect -12043 -27189 -12009 -27155
rect -11975 -27189 -11941 -27155
rect -11907 -27189 -11873 -27155
rect -11839 -27189 -11805 -27155
rect -11771 -27189 -11737 -27155
rect -11703 -27189 -11669 -27155
rect -11635 -27189 -11601 -27155
rect -11567 -27189 -11533 -27155
rect -11499 -27189 -11465 -27155
rect -11431 -27189 -11397 -27155
rect -11363 -27189 -11329 -27155
rect -11295 -27189 -11261 -27155
rect -11227 -27189 -11193 -27155
rect -11159 -27189 -11125 -27155
rect -11091 -27189 -11057 -27155
rect -11023 -27189 -10989 -27155
rect -10955 -27189 -10921 -27155
rect -10887 -27189 -10853 -27155
rect -10819 -27189 -10785 -27155
rect -10751 -27189 -10717 -27155
rect -10683 -27189 -10649 -27155
rect -10615 -27189 -10581 -27155
rect -10547 -27189 -10513 -27155
rect -10479 -27189 -10445 -27155
rect -10411 -27189 -10377 -27155
rect -10343 -27189 -10309 -27155
rect -10275 -27189 -10241 -27155
rect -10207 -27189 -10173 -27155
rect -10139 -27189 -10105 -27155
rect -10071 -27189 -10037 -27155
rect -10003 -27189 -9969 -27155
rect -9935 -27189 -9901 -27155
rect -9867 -27189 -9833 -27155
rect -9799 -27189 -9765 -27155
rect -9731 -27189 -9697 -27155
rect -9663 -27189 -9629 -27155
rect -9595 -27189 -9561 -27155
rect -9527 -27189 -9493 -27155
rect -9459 -27189 -9425 -27155
rect -9391 -27189 -9357 -27155
rect -9323 -27189 -9289 -27155
rect -9255 -27189 -9221 -27155
rect -9187 -27189 -9153 -27155
rect -9119 -27189 -9085 -27155
rect -9051 -27189 -9017 -27155
rect -8983 -27189 -8949 -27155
rect -8915 -27189 -8881 -27155
rect -8847 -27189 -8813 -27155
rect -8779 -27189 -8745 -27155
rect -8711 -27189 -8677 -27155
rect -8643 -27189 -8609 -27155
rect -8575 -27189 -8541 -27155
rect -8507 -27189 -8473 -27155
rect -8439 -27189 -8405 -27155
rect -8371 -27189 -8337 -27155
rect -8303 -27189 -8269 -27155
rect -8235 -27189 -8201 -27155
rect -8167 -27189 -8133 -27155
rect -8099 -27189 -8065 -27155
rect -8031 -27189 -7997 -27155
rect -7963 -27189 -7929 -27155
rect -7895 -27189 -7861 -27155
rect -7827 -27189 -7793 -27155
rect -7759 -27189 -7725 -27155
rect -7691 -27189 -7657 -27155
rect -7623 -27189 -7589 -27155
rect -7555 -27189 -7521 -27155
rect -7487 -27189 -7453 -27155
rect -7419 -27189 -7385 -27155
rect -7351 -27189 -7317 -27155
rect -7283 -27189 -7249 -27155
rect -7215 -27189 -7181 -27155
rect -7147 -27189 -7113 -27155
rect -7079 -27189 -7045 -27155
rect -7011 -27189 -6977 -27155
rect -6943 -27189 -6909 -27155
rect -6875 -27189 -6841 -27155
rect -6807 -27189 -6773 -27155
rect -6739 -27189 -6705 -27155
rect -6671 -27189 -6637 -27155
rect -6603 -27189 -6569 -27155
rect -6535 -27189 -6501 -27155
rect -6467 -27189 -6433 -27155
rect -6399 -27189 -6365 -27155
rect -6331 -27189 -6297 -27155
rect -6263 -27189 -6229 -27155
rect -6195 -27189 -6161 -27155
rect -6127 -27189 -6093 -27155
rect -6059 -27189 -6025 -27155
rect -5991 -27189 -5957 -27155
rect -5923 -27189 -5889 -27155
rect -5855 -27189 -5821 -27155
rect -5787 -27189 -5753 -27155
rect -5719 -27189 -5685 -27155
rect -5651 -27189 -5617 -27155
rect -5583 -27189 -5549 -27155
rect -5515 -27189 -5481 -27155
rect -5447 -27189 -5413 -27155
rect -5379 -27189 -5345 -27155
rect -5311 -27189 -5277 -27155
rect -5243 -27189 -5209 -27155
rect -5175 -27189 -5141 -27155
rect -5107 -27189 -5073 -27155
rect -5039 -27189 -5005 -27155
rect -4971 -27189 -4937 -27155
rect -4903 -27189 -4869 -27155
rect -4835 -27189 -4801 -27155
rect -4767 -27189 -4733 -27155
rect -4699 -27189 -4665 -27155
rect -4631 -27189 -4597 -27155
rect -4563 -27189 -4529 -27155
rect -4495 -27189 -4461 -27155
rect -4427 -27189 -4393 -27155
rect -4359 -27189 -4325 -27155
rect -4291 -27189 -4257 -27155
rect -4223 -27189 -4189 -27155
rect -4155 -27189 -4121 -27155
rect -4087 -27189 -4053 -27155
rect -4019 -27189 -3985 -27155
rect -3951 -27189 -3917 -27155
rect -3883 -27189 -3849 -27155
rect -3815 -27189 -3781 -27155
rect -3747 -27189 -3713 -27155
rect -3679 -27189 -3645 -27155
rect -3611 -27189 -3577 -27155
rect -3543 -27189 -3509 -27155
rect -3475 -27189 -3441 -27155
rect -3407 -27189 -3373 -27155
rect -3339 -27189 -3305 -27155
rect -3271 -27189 -3237 -27155
rect -3203 -27189 -3169 -27155
rect -3135 -27189 -3101 -27155
rect -3067 -27189 -3033 -27155
rect -2999 -27189 -2965 -27155
rect -2931 -27189 -2897 -27155
rect -2863 -27189 -2829 -27155
rect -2795 -27189 -2761 -27155
rect -2727 -27189 -2693 -27155
rect -2659 -27189 -2625 -27155
rect -2591 -27189 -2557 -27155
rect -2523 -27189 -2489 -27155
rect -2455 -27189 -2421 -27155
rect -2387 -27189 -2353 -27155
rect -2319 -27189 -2285 -27155
rect -2251 -27189 -2217 -27155
rect -2183 -27189 -2149 -27155
rect -2115 -27189 -2081 -27155
rect -2047 -27189 -2013 -27155
rect -1979 -27189 -1945 -27155
rect -1911 -27189 -1877 -27155
rect -1843 -27189 -1809 -27155
rect -1775 -27189 -1741 -27155
rect -1707 -27189 -1673 -27155
rect -1639 -27189 -1605 -27155
rect -1571 -27189 -1537 -27155
rect -1503 -27189 -1469 -27155
rect -1435 -27189 -1401 -27155
rect -1367 -27189 -1333 -27155
rect -1299 -27189 -1265 -27155
rect -1231 -27189 -1197 -27155
rect -1163 -27189 -1129 -27155
rect -1095 -27189 -1061 -27155
rect -1027 -27189 -993 -27155
rect -959 -27189 -925 -27155
rect -891 -27189 -857 -27155
rect -823 -27189 -789 -27155
rect -755 -27189 -721 -27155
rect -687 -27189 -653 -27155
rect -619 -27189 -585 -27155
rect -551 -27189 -517 -27155
rect -483 -27189 -449 -27155
rect -415 -27189 -381 -27155
rect -347 -27189 -313 -27155
rect -279 -27189 -245 -27155
rect -211 -27189 -177 -27155
rect -143 -27189 -109 -27155
rect -75 -27189 -41 -27155
rect -7 -27189 27 -27155
rect 61 -27189 95 -27155
rect 129 -27189 163 -27155
rect 197 -27189 231 -27155
rect 265 -27189 299 -27155
rect 333 -27189 367 -27155
rect 401 -27189 435 -27155
rect 469 -27189 503 -27155
rect 537 -27189 571 -27155
rect 605 -27189 639 -27155
rect 673 -27189 707 -27155
rect 741 -27189 775 -27155
rect 809 -27189 843 -27155
rect 877 -27189 911 -27155
rect 945 -27189 979 -27155
rect 1013 -27189 1047 -27155
rect 1081 -27189 1115 -27155
rect 1149 -27189 1183 -27155
rect 1217 -27189 1251 -27155
rect 1285 -27189 1319 -27155
rect 1353 -27189 1387 -27155
rect 1421 -27189 1455 -27155
rect 1489 -27189 1523 -27155
rect 1557 -27189 1591 -27155
rect 1625 -27189 1659 -27155
rect 1693 -27189 1727 -27155
rect 1761 -27189 1795 -27155
rect 1829 -27189 1863 -27155
rect 1897 -27189 1931 -27155
rect 1965 -27189 1999 -27155
rect 2033 -27189 2067 -27155
rect 2101 -27189 2135 -27155
rect 2169 -27189 2203 -27155
rect 2237 -27189 2271 -27155
rect 2305 -27189 2339 -27155
rect 2373 -27189 2407 -27155
rect 2441 -27189 2475 -27155
rect 2509 -27189 2543 -27155
rect 2577 -27189 2611 -27155
rect 2645 -27189 2679 -27155
rect 2713 -27189 2747 -27155
rect 2781 -27189 2815 -27155
rect 2849 -27189 2883 -27155
rect 2917 -27189 2951 -27155
rect 2985 -27189 3019 -27155
rect 3053 -27189 3087 -27155
rect 3121 -27189 3155 -27155
rect 3189 -27189 3223 -27155
rect 3257 -27189 3291 -27155
rect 3325 -27189 3359 -27155
rect 3393 -27189 3427 -27155
rect 3461 -27189 3495 -27155
rect 3529 -27189 3563 -27155
rect 3597 -27189 3631 -27155
rect 3665 -27189 3699 -27155
rect 3733 -27189 3767 -27155
rect 3801 -27189 3835 -27155
rect 3869 -27189 3903 -27155
rect 3937 -27189 3971 -27155
rect 4005 -27189 4039 -27155
rect 4073 -27189 4107 -27155
rect 4141 -27189 4175 -27155
rect 4209 -27189 4243 -27155
rect 4277 -27189 4311 -27155
rect 4345 -27189 4379 -27155
rect 4413 -27189 4447 -27155
rect 4481 -27189 4515 -27155
rect 4549 -27189 4583 -27155
rect 4617 -27189 4651 -27155
rect 4685 -27189 4719 -27155
rect 4753 -27189 4787 -27155
rect 4821 -27189 4855 -27155
rect 4889 -27189 4923 -27155
rect 4957 -27189 4991 -27155
rect 5025 -27189 5059 -27155
rect 5093 -27189 5127 -27155
rect 5161 -27189 5195 -27155
rect 5229 -27189 5263 -27155
rect 5297 -27189 5331 -27155
rect 5365 -27189 5399 -27155
rect 5433 -27189 5467 -27155
rect 5501 -27189 5535 -27155
rect 5569 -27189 5603 -27155
rect 5637 -27189 5671 -27155
rect 5705 -27189 5739 -27155
rect 5773 -27189 5807 -27155
rect 5841 -27189 5875 -27155
rect 5909 -27189 5943 -27155
rect 5977 -27189 6011 -27155
rect 6045 -27189 6079 -27155
rect 6113 -27189 6147 -27155
rect 6181 -27189 6215 -27155
rect 6249 -27189 6283 -27155
rect 6317 -27189 6351 -27155
rect 6385 -27189 6419 -27155
rect 6453 -27189 6487 -27155
rect 6521 -27189 6555 -27155
rect 6589 -27189 6623 -27155
rect 6657 -27189 6691 -27155
rect 6725 -27189 6759 -27155
rect 6793 -27189 6827 -27155
rect 6861 -27189 6895 -27155
rect 6929 -27189 6963 -27155
rect 6997 -27189 7031 -27155
rect 7065 -27189 7099 -27155
rect 7133 -27189 7167 -27155
rect 7201 -27189 7235 -27155
rect 7269 -27189 7303 -27155
rect 7337 -27189 7371 -27155
rect 7405 -27189 7439 -27155
rect 7473 -27189 7507 -27155
rect 7541 -27189 7575 -27155
rect 7609 -27189 7643 -27155
rect 7677 -27189 7711 -27155
rect 7745 -27189 7779 -27155
rect 7813 -27189 7847 -27155
rect 7881 -27189 7915 -27155
rect 7949 -27189 7983 -27155
rect 8017 -27189 8051 -27155
rect 8085 -27189 8119 -27155
rect 8153 -27189 8187 -27155
rect 8221 -27189 8255 -27155
rect 8289 -27189 8323 -27155
rect 8357 -27189 8391 -27155
rect 8425 -27189 8459 -27155
rect 8493 -27189 8527 -27155
rect 8561 -27189 8595 -27155
rect 8629 -27189 8663 -27155
rect 8697 -27189 8731 -27155
rect 8765 -27189 8799 -27155
rect 8833 -27189 8867 -27155
rect 8901 -27189 8935 -27155
rect 8969 -27189 9003 -27155
rect 9037 -27189 9071 -27155
rect 9105 -27189 9139 -27155
rect 9173 -27189 9207 -27155
rect 9241 -27189 9275 -27155
rect 9309 -27189 9343 -27155
rect 9377 -27189 9411 -27155
rect 9445 -27189 9479 -27155
rect 9513 -27189 9547 -27155
rect 9581 -27189 9615 -27155
rect 9649 -27189 9683 -27155
rect 9717 -27189 9751 -27155
rect 9785 -27189 9819 -27155
rect 9853 -27189 9887 -27155
rect 9921 -27189 9955 -27155
rect 9989 -27189 10023 -27155
rect 10057 -27189 10091 -27155
rect 10125 -27189 10159 -27155
rect 10193 -27189 10227 -27155
rect 10261 -27189 10295 -27155
rect 10329 -27189 10363 -27155
rect 10397 -27189 10431 -27155
rect 10465 -27189 10499 -27155
rect 10533 -27189 10567 -27155
rect 10601 -27189 10635 -27155
rect 10669 -27189 10703 -27155
rect 10737 -27189 10771 -27155
rect 10805 -27189 10839 -27155
rect 10873 -27189 10907 -27155
rect 10941 -27189 10975 -27155
rect 11009 -27189 11043 -27155
rect 11077 -27189 11111 -27155
rect 11145 -27189 11179 -27155
rect 11213 -27189 11247 -27155
rect 11281 -27189 11315 -27155
rect 11349 -27189 11383 -27155
rect 11417 -27189 11451 -27155
rect 11485 -27189 11519 -27155
rect 11553 -27189 11587 -27155
rect 11621 -27189 11655 -27155
rect 11689 -27189 11723 -27155
rect 11757 -27189 11791 -27155
rect 11825 -27189 11859 -27155
rect 11893 -27189 11927 -27155
rect 11961 -27189 11995 -27155
rect 12029 -27189 12063 -27155
rect 12097 -27189 12131 -27155
rect 12165 -27189 12199 -27155
rect 12233 -27189 12267 -27155
rect 12301 -27189 12335 -27155
rect 12369 -27189 12403 -27155
rect 12437 -27189 12471 -27155
rect 12505 -27189 12539 -27155
rect 12573 -27189 12607 -27155
rect 12641 -27189 12675 -27155
rect 12709 -27189 12743 -27155
rect 12777 -27189 12811 -27155
rect 12845 -27189 12879 -27155
rect 12913 -27189 12947 -27155
rect 12981 -27189 13015 -27155
rect 13049 -27189 13083 -27155
rect 13117 -27189 13151 -27155
rect 13185 -27189 13219 -27155
rect 13253 -27189 13287 -27155
rect 13321 -27189 13355 -27155
rect 13389 -27189 13423 -27155
rect 13457 -27189 13491 -27155
rect 13525 -27189 13559 -27155
rect 13593 -27189 13627 -27155
rect 13661 -27189 13695 -27155
rect 13729 -27189 13763 -27155
rect 13797 -27189 13831 -27155
rect 13865 -27189 13899 -27155
rect 13933 -27189 13967 -27155
rect 14001 -27189 14035 -27155
rect 14069 -27189 14103 -27155
rect 14137 -27189 14171 -27155
rect 14205 -27189 14239 -27155
rect 14273 -27189 14307 -27155
rect 14341 -27189 14375 -27155
rect 14409 -27189 14443 -27155
rect 14477 -27189 14511 -27155
rect 14545 -27189 14579 -27155
rect 14613 -27189 14647 -27155
rect 14681 -27189 14715 -27155
rect 14749 -27189 14783 -27155
rect 14817 -27189 14851 -27155
rect 14885 -27189 14919 -27155
rect 14953 -27189 14987 -27155
rect 15021 -27189 15055 -27155
rect 15089 -27189 15123 -27155
rect 15157 -27189 15191 -27155
rect 15225 -27189 15259 -27155
rect 15293 -27189 15327 -27155
rect 15361 -27189 15395 -27155
rect 15429 -27189 15463 -27155
rect 15497 -27189 15531 -27155
rect 15565 -27189 15599 -27155
rect 15633 -27189 15667 -27155
rect 15701 -27189 15735 -27155
rect 15769 -27189 15803 -27155
rect 15837 -27189 15871 -27155
rect 15905 -27189 15939 -27155
rect 15973 -27189 16007 -27155
rect 16041 -27189 16075 -27155
rect 16109 -27189 16143 -27155
rect 16177 -27189 16211 -27155
rect 16245 -27189 16279 -27155
rect 16313 -27189 16347 -27155
rect 16381 -27189 16415 -27155
rect 16449 -27189 16483 -27155
rect 16517 -27189 16551 -27155
rect 16585 -27189 16619 -27155
rect 16653 -27189 16687 -27155
rect 16721 -27189 16755 -27155
rect 16789 -27189 16823 -27155
rect 16857 -27189 16891 -27155
rect 16925 -27189 16959 -27155
rect 16993 -27189 17027 -27155
rect 17061 -27189 17095 -27155
rect 17129 -27189 17163 -27155
rect 17197 -27189 17231 -27155
rect 17265 -27189 17299 -27155
rect 17333 -27189 17367 -27155
rect 17401 -27189 17435 -27155
rect 17469 -27189 17503 -27155
rect 17537 -27189 17571 -27155
rect 17605 -27189 17639 -27155
rect 17673 -27189 17707 -27155
rect 17741 -27189 17775 -27155
rect 17809 -27189 17843 -27155
rect 17877 -27189 17911 -27155
rect 17945 -27189 17979 -27155
rect 18013 -27189 18047 -27155
rect 18081 -27189 18115 -27155
rect 18149 -27189 18183 -27155
rect 18217 -27189 18251 -27155
rect 18285 -27189 18319 -27155
rect 18353 -27189 18387 -27155
rect 18421 -27189 18455 -27155
rect 18489 -27189 18523 -27155
rect 18557 -27189 18591 -27155
rect 18625 -27189 18659 -27155
rect 18693 -27189 18727 -27155
rect 18761 -27189 18795 -27155
rect 18829 -27189 18863 -27155
rect 18897 -27189 18931 -27155
rect 18965 -27189 18999 -27155
rect 19033 -27189 19067 -27155
rect 19101 -27189 19135 -27155
rect 19169 -27189 19203 -27155
rect 19237 -27189 19271 -27155
rect 19305 -27189 19339 -27155
rect 19373 -27189 19407 -27155
rect 19441 -27189 19475 -27155
rect 19509 -27189 19543 -27155
rect 19577 -27189 19611 -27155
rect 19645 -27189 19679 -27155
rect 19713 -27189 19747 -27155
rect 19781 -27189 19815 -27155
rect 19849 -27189 19883 -27155
rect 19917 -27189 19951 -27155
rect 19985 -27189 20019 -27155
rect 20053 -27189 20087 -27155
rect 20121 -27189 20155 -27155
rect 20189 -27189 20223 -27155
rect 20257 -27189 20291 -27155
rect 20325 -27189 20359 -27155
rect 20393 -27189 20427 -27155
rect 20461 -27189 20495 -27155
rect 20529 -27189 20563 -27155
rect 20597 -27189 20631 -27155
rect 20665 -27189 20699 -27155
rect 20733 -27189 20767 -27155
rect 20801 -27189 20835 -27155
rect 20869 -27189 20903 -27155
rect 20937 -27189 20971 -27155
rect 21005 -27189 21039 -27155
rect 21073 -27189 21107 -27155
rect 21141 -27189 21175 -27155
rect 21209 -27189 21243 -27155
rect 21277 -27189 21311 -27155
rect 21345 -27189 21379 -27155
rect 21413 -27189 21447 -27155
rect 21481 -27189 21515 -27155
rect 21549 -27189 21583 -27155
rect 21617 -27189 21651 -27155
rect 21685 -27189 21719 -27155
rect 21753 -27189 21787 -27155
rect 21821 -27189 21855 -27155
rect 21889 -27189 21923 -27155
rect 21957 -27189 21991 -27155
rect 22025 -27189 22059 -27155
rect 22093 -27189 22127 -27155
rect 22161 -27189 22195 -27155
rect 22229 -27189 22263 -27155
rect 22297 -27189 22331 -27155
rect 22365 -27189 22399 -27155
rect 22433 -27189 22467 -27155
rect 22501 -27189 22535 -27155
rect 22569 -27189 22603 -27155
rect 22637 -27189 22671 -27155
rect 22705 -27189 22739 -27155
rect 22773 -27189 22807 -27155
rect 22841 -27189 22875 -27155
rect 22909 -27189 22943 -27155
rect 22977 -27189 23011 -27155
rect 23045 -27189 23079 -27155
rect 23113 -27189 23147 -27155
rect 23181 -27189 23215 -27155
rect 23249 -27189 23283 -27155
rect 23317 -27189 23351 -27155
rect 23385 -27189 23419 -27155
rect 23453 -27189 23487 -27155
rect 23521 -27189 23555 -27155
rect 23589 -27189 23623 -27155
rect 23657 -27189 23691 -27155
rect 23725 -27189 23759 -27155
rect 23793 -27189 23827 -27155
rect 23861 -27189 23895 -27155
rect 23929 -27189 23963 -27155
rect 23997 -27189 24031 -27155
rect 24065 -27189 24099 -27155
rect 24133 -27189 24167 -27155
rect 24201 -27189 24235 -27155
rect 24269 -27189 24303 -27155
rect 24337 -27189 24371 -27155
rect 24405 -27189 24439 -27155
rect 24473 -27189 24507 -27155
rect 24541 -27189 24575 -27155
rect 24609 -27189 24643 -27155
rect 24677 -27189 24711 -27155
rect 24745 -27189 24922 -27155
rect -12322 -27222 24922 -27189
<< nsubdiff >>
rect 378 1689 24822 1722
rect 378 1655 547 1689
rect 581 1655 615 1689
rect 649 1655 683 1689
rect 717 1655 751 1689
rect 785 1655 819 1689
rect 853 1655 887 1689
rect 921 1655 955 1689
rect 989 1655 1023 1689
rect 1057 1655 1091 1689
rect 1125 1655 1159 1689
rect 1193 1655 1227 1689
rect 1261 1655 1295 1689
rect 1329 1655 1363 1689
rect 1397 1655 1431 1689
rect 1465 1655 1499 1689
rect 1533 1655 1567 1689
rect 1601 1655 1635 1689
rect 1669 1655 1703 1689
rect 1737 1655 1771 1689
rect 1805 1655 1839 1689
rect 1873 1655 1907 1689
rect 1941 1655 1975 1689
rect 2009 1655 2043 1689
rect 2077 1655 2111 1689
rect 2145 1655 2179 1689
rect 2213 1655 2247 1689
rect 2281 1655 2315 1689
rect 2349 1655 2383 1689
rect 2417 1655 2451 1689
rect 2485 1655 2519 1689
rect 2553 1655 2587 1689
rect 2621 1655 2655 1689
rect 2689 1655 2723 1689
rect 2757 1655 2791 1689
rect 2825 1655 2859 1689
rect 2893 1655 2927 1689
rect 2961 1655 2995 1689
rect 3029 1655 3063 1689
rect 3097 1655 3131 1689
rect 3165 1655 3199 1689
rect 3233 1655 3267 1689
rect 3301 1655 3335 1689
rect 3369 1655 3403 1689
rect 3437 1655 3471 1689
rect 3505 1655 3539 1689
rect 3573 1655 3607 1689
rect 3641 1655 3675 1689
rect 3709 1655 3743 1689
rect 3777 1655 3811 1689
rect 3845 1655 3879 1689
rect 3913 1655 3947 1689
rect 3981 1655 4015 1689
rect 4049 1655 4083 1689
rect 4117 1655 4151 1689
rect 4185 1655 4219 1689
rect 4253 1655 4287 1689
rect 4321 1655 4355 1689
rect 4389 1655 4423 1689
rect 4457 1655 4491 1689
rect 4525 1655 4559 1689
rect 4593 1655 4627 1689
rect 4661 1655 4695 1689
rect 4729 1655 4763 1689
rect 4797 1655 4831 1689
rect 4865 1655 4899 1689
rect 4933 1655 4967 1689
rect 5001 1655 5035 1689
rect 5069 1655 5103 1689
rect 5137 1655 5171 1689
rect 5205 1655 5239 1689
rect 5273 1655 5307 1689
rect 5341 1655 5375 1689
rect 5409 1655 5443 1689
rect 5477 1655 5511 1689
rect 5545 1655 5579 1689
rect 5613 1655 5647 1689
rect 5681 1655 5715 1689
rect 5749 1655 5783 1689
rect 5817 1655 5851 1689
rect 5885 1655 5919 1689
rect 5953 1655 5987 1689
rect 6021 1655 6055 1689
rect 6089 1655 6123 1689
rect 6157 1655 6191 1689
rect 6225 1655 6259 1689
rect 6293 1655 6327 1689
rect 6361 1655 6395 1689
rect 6429 1655 6463 1689
rect 6497 1655 6531 1689
rect 6565 1655 6599 1689
rect 6633 1655 6667 1689
rect 6701 1655 6735 1689
rect 6769 1655 6803 1689
rect 6837 1655 6871 1689
rect 6905 1655 6939 1689
rect 6973 1655 7007 1689
rect 7041 1655 7075 1689
rect 7109 1655 7143 1689
rect 7177 1655 7211 1689
rect 7245 1655 7279 1689
rect 7313 1655 7347 1689
rect 7381 1655 7415 1689
rect 7449 1655 7483 1689
rect 7517 1655 7551 1689
rect 7585 1655 7619 1689
rect 7653 1655 7687 1689
rect 7721 1655 7755 1689
rect 7789 1655 7823 1689
rect 7857 1655 7891 1689
rect 7925 1655 7959 1689
rect 7993 1655 8027 1689
rect 8061 1655 8095 1689
rect 8129 1655 8163 1689
rect 8197 1655 8231 1689
rect 8265 1655 8299 1689
rect 8333 1655 8367 1689
rect 8401 1655 8435 1689
rect 8469 1655 8503 1689
rect 8537 1655 8571 1689
rect 8605 1655 8639 1689
rect 8673 1655 8707 1689
rect 8741 1655 8775 1689
rect 8809 1655 8843 1689
rect 8877 1655 8911 1689
rect 8945 1655 8979 1689
rect 9013 1655 9047 1689
rect 9081 1655 9115 1689
rect 9149 1655 9183 1689
rect 9217 1655 9251 1689
rect 9285 1655 9319 1689
rect 9353 1655 9387 1689
rect 9421 1655 9455 1689
rect 9489 1655 9523 1689
rect 9557 1655 9591 1689
rect 9625 1655 9659 1689
rect 9693 1655 9727 1689
rect 9761 1655 9795 1689
rect 9829 1655 9863 1689
rect 9897 1655 9931 1689
rect 9965 1655 9999 1689
rect 10033 1655 10067 1689
rect 10101 1655 10135 1689
rect 10169 1655 10203 1689
rect 10237 1655 10271 1689
rect 10305 1655 10339 1689
rect 10373 1655 10407 1689
rect 10441 1655 10475 1689
rect 10509 1655 10543 1689
rect 10577 1655 10611 1689
rect 10645 1655 10679 1689
rect 10713 1655 10747 1689
rect 10781 1655 10815 1689
rect 10849 1655 10883 1689
rect 10917 1655 10951 1689
rect 10985 1655 11019 1689
rect 11053 1655 11087 1689
rect 11121 1655 11155 1689
rect 11189 1655 11223 1689
rect 11257 1655 11291 1689
rect 11325 1655 11359 1689
rect 11393 1655 11427 1689
rect 11461 1655 11495 1689
rect 11529 1655 11563 1689
rect 11597 1655 11631 1689
rect 11665 1655 11699 1689
rect 11733 1655 11767 1689
rect 11801 1655 11835 1689
rect 11869 1655 11903 1689
rect 11937 1655 11971 1689
rect 12005 1655 12039 1689
rect 12073 1655 12107 1689
rect 12141 1655 12175 1689
rect 12209 1655 12243 1689
rect 12277 1655 12311 1689
rect 12345 1655 12379 1689
rect 12413 1655 12447 1689
rect 12481 1655 12515 1689
rect 12549 1655 12583 1689
rect 12617 1655 12651 1689
rect 12685 1655 12719 1689
rect 12753 1655 12787 1689
rect 12821 1655 12855 1689
rect 12889 1655 12923 1689
rect 12957 1655 12991 1689
rect 13025 1655 13059 1689
rect 13093 1655 13127 1689
rect 13161 1655 13195 1689
rect 13229 1655 13263 1689
rect 13297 1655 13331 1689
rect 13365 1655 13399 1689
rect 13433 1655 13467 1689
rect 13501 1655 13535 1689
rect 13569 1655 13603 1689
rect 13637 1655 13671 1689
rect 13705 1655 13739 1689
rect 13773 1655 13807 1689
rect 13841 1655 13875 1689
rect 13909 1655 13943 1689
rect 13977 1655 14011 1689
rect 14045 1655 14079 1689
rect 14113 1655 14147 1689
rect 14181 1655 14215 1689
rect 14249 1655 14283 1689
rect 14317 1655 14351 1689
rect 14385 1655 14419 1689
rect 14453 1655 14487 1689
rect 14521 1655 14555 1689
rect 14589 1655 14623 1689
rect 14657 1655 14691 1689
rect 14725 1655 14759 1689
rect 14793 1655 14827 1689
rect 14861 1655 14895 1689
rect 14929 1655 14963 1689
rect 14997 1655 15031 1689
rect 15065 1655 15099 1689
rect 15133 1655 15167 1689
rect 15201 1655 15235 1689
rect 15269 1655 15303 1689
rect 15337 1655 15371 1689
rect 15405 1655 15439 1689
rect 15473 1655 15507 1689
rect 15541 1655 15575 1689
rect 15609 1655 15643 1689
rect 15677 1655 15711 1689
rect 15745 1655 15779 1689
rect 15813 1655 15847 1689
rect 15881 1655 15915 1689
rect 15949 1655 15983 1689
rect 16017 1655 16051 1689
rect 16085 1655 16119 1689
rect 16153 1655 16187 1689
rect 16221 1655 16255 1689
rect 16289 1655 16323 1689
rect 16357 1655 16391 1689
rect 16425 1655 16459 1689
rect 16493 1655 16527 1689
rect 16561 1655 16595 1689
rect 16629 1655 16663 1689
rect 16697 1655 16731 1689
rect 16765 1655 16799 1689
rect 16833 1655 16867 1689
rect 16901 1655 16935 1689
rect 16969 1655 17003 1689
rect 17037 1655 17071 1689
rect 17105 1655 17139 1689
rect 17173 1655 17207 1689
rect 17241 1655 17275 1689
rect 17309 1655 17343 1689
rect 17377 1655 17411 1689
rect 17445 1655 17479 1689
rect 17513 1655 17547 1689
rect 17581 1655 17615 1689
rect 17649 1655 17683 1689
rect 17717 1655 17751 1689
rect 17785 1655 17819 1689
rect 17853 1655 17887 1689
rect 17921 1655 17955 1689
rect 17989 1655 18023 1689
rect 18057 1655 18091 1689
rect 18125 1655 18159 1689
rect 18193 1655 18227 1689
rect 18261 1655 18295 1689
rect 18329 1655 18363 1689
rect 18397 1655 18431 1689
rect 18465 1655 18499 1689
rect 18533 1655 18567 1689
rect 18601 1655 18635 1689
rect 18669 1655 18703 1689
rect 18737 1655 18771 1689
rect 18805 1655 18839 1689
rect 18873 1655 18907 1689
rect 18941 1655 18975 1689
rect 19009 1655 19043 1689
rect 19077 1655 19111 1689
rect 19145 1655 19179 1689
rect 19213 1655 19247 1689
rect 19281 1655 19315 1689
rect 19349 1655 19383 1689
rect 19417 1655 19451 1689
rect 19485 1655 19519 1689
rect 19553 1655 19587 1689
rect 19621 1655 19655 1689
rect 19689 1655 19723 1689
rect 19757 1655 19791 1689
rect 19825 1655 19859 1689
rect 19893 1655 19927 1689
rect 19961 1655 19995 1689
rect 20029 1655 20063 1689
rect 20097 1655 20131 1689
rect 20165 1655 20199 1689
rect 20233 1655 20267 1689
rect 20301 1655 20335 1689
rect 20369 1655 20403 1689
rect 20437 1655 20471 1689
rect 20505 1655 20539 1689
rect 20573 1655 20607 1689
rect 20641 1655 20675 1689
rect 20709 1655 20743 1689
rect 20777 1655 20811 1689
rect 20845 1655 20879 1689
rect 20913 1655 20947 1689
rect 20981 1655 21015 1689
rect 21049 1655 21083 1689
rect 21117 1655 21151 1689
rect 21185 1655 21219 1689
rect 21253 1655 21287 1689
rect 21321 1655 21355 1689
rect 21389 1655 21423 1689
rect 21457 1655 21491 1689
rect 21525 1655 21559 1689
rect 21593 1655 21627 1689
rect 21661 1655 21695 1689
rect 21729 1655 21763 1689
rect 21797 1655 21831 1689
rect 21865 1655 21899 1689
rect 21933 1655 21967 1689
rect 22001 1655 22035 1689
rect 22069 1655 22103 1689
rect 22137 1655 22171 1689
rect 22205 1655 22239 1689
rect 22273 1655 22307 1689
rect 22341 1655 22375 1689
rect 22409 1655 22443 1689
rect 22477 1655 22511 1689
rect 22545 1655 22579 1689
rect 22613 1655 22647 1689
rect 22681 1655 22715 1689
rect 22749 1655 22783 1689
rect 22817 1655 22851 1689
rect 22885 1655 22919 1689
rect 22953 1655 22987 1689
rect 23021 1655 23055 1689
rect 23089 1655 23123 1689
rect 23157 1655 23191 1689
rect 23225 1655 23259 1689
rect 23293 1655 23327 1689
rect 23361 1655 23395 1689
rect 23429 1655 23463 1689
rect 23497 1655 23531 1689
rect 23565 1655 23599 1689
rect 23633 1655 23667 1689
rect 23701 1655 23735 1689
rect 23769 1655 23803 1689
rect 23837 1655 23871 1689
rect 23905 1655 23939 1689
rect 23973 1655 24007 1689
rect 24041 1655 24075 1689
rect 24109 1655 24143 1689
rect 24177 1655 24211 1689
rect 24245 1655 24279 1689
rect 24313 1655 24347 1689
rect 24381 1655 24415 1689
rect 24449 1655 24483 1689
rect 24517 1655 24551 1689
rect 24585 1655 24619 1689
rect 24653 1655 24822 1689
rect 378 1622 24822 1655
rect 378 1537 478 1622
rect 378 1503 411 1537
rect 445 1503 478 1537
rect 378 1469 478 1503
rect 378 1435 411 1469
rect 445 1435 478 1469
rect 378 1401 478 1435
rect 378 1367 411 1401
rect 445 1367 478 1401
rect 378 1333 478 1367
rect 378 1299 411 1333
rect 445 1299 478 1333
rect 378 1265 478 1299
rect 378 1231 411 1265
rect 445 1231 478 1265
rect 378 1197 478 1231
rect 378 1163 411 1197
rect 445 1163 478 1197
rect 378 1129 478 1163
rect 378 1095 411 1129
rect 445 1095 478 1129
rect 378 1061 478 1095
rect 378 1027 411 1061
rect 445 1027 478 1061
rect 378 993 478 1027
rect 378 959 411 993
rect 445 959 478 993
rect 378 925 478 959
rect 378 891 411 925
rect 445 891 478 925
rect 378 857 478 891
rect 378 823 411 857
rect 445 823 478 857
rect 378 789 478 823
rect 378 755 411 789
rect 445 755 478 789
rect 378 721 478 755
rect 378 687 411 721
rect 445 687 478 721
rect 378 653 478 687
rect 378 619 411 653
rect 445 619 478 653
rect 378 585 478 619
rect 378 551 411 585
rect 445 551 478 585
rect 378 517 478 551
rect 378 483 411 517
rect 445 483 478 517
rect 378 449 478 483
rect 378 415 411 449
rect 445 415 478 449
rect 378 381 478 415
rect 378 347 411 381
rect 445 347 478 381
rect 378 313 478 347
rect 378 279 411 313
rect 445 279 478 313
rect 378 245 478 279
rect 378 211 411 245
rect 445 211 478 245
rect 378 177 478 211
rect 378 143 411 177
rect 445 143 478 177
rect 378 109 478 143
rect 378 75 411 109
rect 445 75 478 109
rect 378 41 478 75
rect 378 7 411 41
rect 445 7 478 41
rect 378 -27 478 7
rect 378 -61 411 -27
rect 445 -61 478 -27
rect 378 -95 478 -61
rect 378 -129 411 -95
rect 445 -129 478 -95
rect 378 -163 478 -129
rect 378 -197 411 -163
rect 445 -197 478 -163
rect 378 -231 478 -197
rect 378 -265 411 -231
rect 445 -265 478 -231
rect 378 -299 478 -265
rect 378 -333 411 -299
rect 445 -333 478 -299
rect 378 -367 478 -333
rect 378 -401 411 -367
rect 445 -401 478 -367
rect 378 -435 478 -401
rect 378 -469 411 -435
rect 445 -469 478 -435
rect 378 -503 478 -469
rect 378 -537 411 -503
rect 445 -537 478 -503
rect 378 -571 478 -537
rect 378 -605 411 -571
rect 445 -605 478 -571
rect 378 -639 478 -605
rect 378 -673 411 -639
rect 445 -673 478 -639
rect 378 -707 478 -673
rect 378 -741 411 -707
rect 445 -741 478 -707
rect 378 -775 478 -741
rect 378 -809 411 -775
rect 445 -809 478 -775
rect 378 -843 478 -809
rect 378 -877 411 -843
rect 445 -877 478 -843
rect 378 -911 478 -877
rect 378 -945 411 -911
rect 445 -945 478 -911
rect 378 -979 478 -945
rect 378 -1013 411 -979
rect 445 -1013 478 -979
rect 378 -1047 478 -1013
rect 378 -1081 411 -1047
rect 445 -1081 478 -1047
rect 378 -1115 478 -1081
rect 378 -1149 411 -1115
rect 445 -1149 478 -1115
rect 378 -1183 478 -1149
rect 378 -1217 411 -1183
rect 445 -1217 478 -1183
rect 378 -1251 478 -1217
rect 378 -1285 411 -1251
rect 445 -1285 478 -1251
rect 378 -1319 478 -1285
rect 378 -1353 411 -1319
rect 445 -1353 478 -1319
rect 378 -1387 478 -1353
rect 378 -1421 411 -1387
rect 445 -1421 478 -1387
rect 378 -1455 478 -1421
rect 378 -1489 411 -1455
rect 445 -1489 478 -1455
rect 378 -1523 478 -1489
rect 378 -1557 411 -1523
rect 445 -1557 478 -1523
rect 378 -1591 478 -1557
rect 378 -1625 411 -1591
rect 445 -1625 478 -1591
rect 378 -1659 478 -1625
rect 378 -1693 411 -1659
rect 445 -1693 478 -1659
rect 378 -1727 478 -1693
rect 378 -1761 411 -1727
rect 445 -1761 478 -1727
rect 378 -1795 478 -1761
rect 378 -1829 411 -1795
rect 445 -1829 478 -1795
rect 378 -1863 478 -1829
rect 378 -1897 411 -1863
rect 445 -1897 478 -1863
rect 378 -1931 478 -1897
rect 378 -1965 411 -1931
rect 445 -1965 478 -1931
rect 378 -1999 478 -1965
rect 378 -2033 411 -1999
rect 445 -2033 478 -1999
rect 378 -2067 478 -2033
rect 378 -2101 411 -2067
rect 445 -2101 478 -2067
rect 378 -2135 478 -2101
rect 378 -2169 411 -2135
rect 445 -2169 478 -2135
rect 378 -2203 478 -2169
rect 378 -2237 411 -2203
rect 445 -2237 478 -2203
rect 378 -2271 478 -2237
rect 378 -2305 411 -2271
rect 445 -2305 478 -2271
rect 378 -2339 478 -2305
rect 378 -2373 411 -2339
rect 445 -2373 478 -2339
rect 378 -2407 478 -2373
rect 378 -2441 411 -2407
rect 445 -2441 478 -2407
rect 378 -2475 478 -2441
rect 378 -2509 411 -2475
rect 445 -2509 478 -2475
rect 378 -2543 478 -2509
rect 378 -2577 411 -2543
rect 445 -2577 478 -2543
rect 378 -2611 478 -2577
rect 378 -2645 411 -2611
rect 445 -2645 478 -2611
rect 378 -2679 478 -2645
rect 378 -2713 411 -2679
rect 445 -2713 478 -2679
rect 378 -2747 478 -2713
rect 378 -2781 411 -2747
rect 445 -2781 478 -2747
rect 378 -2815 478 -2781
rect 378 -2849 411 -2815
rect 445 -2849 478 -2815
rect 378 -2883 478 -2849
rect 378 -2917 411 -2883
rect 445 -2917 478 -2883
rect 378 -2951 478 -2917
rect 378 -2985 411 -2951
rect 445 -2985 478 -2951
rect 378 -3019 478 -2985
rect 378 -3053 411 -3019
rect 445 -3053 478 -3019
rect 378 -3087 478 -3053
rect 378 -3121 411 -3087
rect 445 -3121 478 -3087
rect 378 -3155 478 -3121
rect 378 -3189 411 -3155
rect 445 -3189 478 -3155
rect 378 -3223 478 -3189
rect 378 -3257 411 -3223
rect 445 -3257 478 -3223
rect 378 -3291 478 -3257
rect 378 -3325 411 -3291
rect 445 -3325 478 -3291
rect 378 -3359 478 -3325
rect 378 -3393 411 -3359
rect 445 -3393 478 -3359
rect 378 -3427 478 -3393
rect 378 -3461 411 -3427
rect 445 -3461 478 -3427
rect 378 -3495 478 -3461
rect 378 -3529 411 -3495
rect 445 -3529 478 -3495
rect 378 -3563 478 -3529
rect 378 -3597 411 -3563
rect 445 -3597 478 -3563
rect 378 -3631 478 -3597
rect 378 -3665 411 -3631
rect 445 -3665 478 -3631
rect 378 -3699 478 -3665
rect 378 -3733 411 -3699
rect 445 -3733 478 -3699
rect 378 -3767 478 -3733
rect 378 -3801 411 -3767
rect 445 -3801 478 -3767
rect 378 -3835 478 -3801
rect 378 -3869 411 -3835
rect 445 -3869 478 -3835
rect 378 -3903 478 -3869
rect 378 -3937 411 -3903
rect 445 -3937 478 -3903
rect 378 -3971 478 -3937
rect 378 -4005 411 -3971
rect 445 -4005 478 -3971
rect 378 -4039 478 -4005
rect 378 -4073 411 -4039
rect 445 -4073 478 -4039
rect 378 -4107 478 -4073
rect 378 -4141 411 -4107
rect 445 -4141 478 -4107
rect 378 -4175 478 -4141
rect 378 -4209 411 -4175
rect 445 -4209 478 -4175
rect 378 -4243 478 -4209
rect 378 -4277 411 -4243
rect 445 -4277 478 -4243
rect 378 -4311 478 -4277
rect 378 -4345 411 -4311
rect 445 -4345 478 -4311
rect 378 -4379 478 -4345
rect 378 -4413 411 -4379
rect 445 -4413 478 -4379
rect 378 -4447 478 -4413
rect 378 -4481 411 -4447
rect 445 -4481 478 -4447
rect 378 -4515 478 -4481
rect 378 -4549 411 -4515
rect 445 -4549 478 -4515
rect 378 -4583 478 -4549
rect 378 -4617 411 -4583
rect 445 -4617 478 -4583
rect 24722 1537 24822 1622
rect 24722 1503 24755 1537
rect 24789 1503 24822 1537
rect 24722 1469 24822 1503
rect 24722 1435 24755 1469
rect 24789 1435 24822 1469
rect 24722 1401 24822 1435
rect 24722 1367 24755 1401
rect 24789 1367 24822 1401
rect 24722 1333 24822 1367
rect 24722 1299 24755 1333
rect 24789 1299 24822 1333
rect 24722 1265 24822 1299
rect 24722 1231 24755 1265
rect 24789 1231 24822 1265
rect 24722 1197 24822 1231
rect 24722 1163 24755 1197
rect 24789 1163 24822 1197
rect 24722 1129 24822 1163
rect 24722 1095 24755 1129
rect 24789 1095 24822 1129
rect 24722 1061 24822 1095
rect 24722 1027 24755 1061
rect 24789 1027 24822 1061
rect 24722 993 24822 1027
rect 24722 959 24755 993
rect 24789 959 24822 993
rect 24722 925 24822 959
rect 24722 891 24755 925
rect 24789 891 24822 925
rect 24722 857 24822 891
rect 24722 823 24755 857
rect 24789 823 24822 857
rect 24722 789 24822 823
rect 24722 755 24755 789
rect 24789 755 24822 789
rect 24722 721 24822 755
rect 24722 687 24755 721
rect 24789 687 24822 721
rect 24722 653 24822 687
rect 24722 619 24755 653
rect 24789 619 24822 653
rect 24722 585 24822 619
rect 24722 551 24755 585
rect 24789 551 24822 585
rect 24722 517 24822 551
rect 24722 483 24755 517
rect 24789 483 24822 517
rect 24722 449 24822 483
rect 24722 415 24755 449
rect 24789 415 24822 449
rect 24722 381 24822 415
rect 24722 347 24755 381
rect 24789 347 24822 381
rect 24722 313 24822 347
rect 24722 279 24755 313
rect 24789 279 24822 313
rect 24722 245 24822 279
rect 24722 211 24755 245
rect 24789 211 24822 245
rect 24722 177 24822 211
rect 24722 143 24755 177
rect 24789 143 24822 177
rect 24722 109 24822 143
rect 24722 75 24755 109
rect 24789 75 24822 109
rect 24722 41 24822 75
rect 24722 7 24755 41
rect 24789 7 24822 41
rect 24722 -27 24822 7
rect 24722 -61 24755 -27
rect 24789 -61 24822 -27
rect 24722 -95 24822 -61
rect 24722 -129 24755 -95
rect 24789 -129 24822 -95
rect 24722 -163 24822 -129
rect 24722 -197 24755 -163
rect 24789 -197 24822 -163
rect 24722 -231 24822 -197
rect 24722 -265 24755 -231
rect 24789 -265 24822 -231
rect 24722 -299 24822 -265
rect 24722 -333 24755 -299
rect 24789 -333 24822 -299
rect 24722 -367 24822 -333
rect 24722 -401 24755 -367
rect 24789 -401 24822 -367
rect 24722 -435 24822 -401
rect 24722 -469 24755 -435
rect 24789 -469 24822 -435
rect 24722 -503 24822 -469
rect 24722 -537 24755 -503
rect 24789 -537 24822 -503
rect 24722 -571 24822 -537
rect 24722 -605 24755 -571
rect 24789 -605 24822 -571
rect 24722 -639 24822 -605
rect 24722 -673 24755 -639
rect 24789 -673 24822 -639
rect 24722 -707 24822 -673
rect 24722 -741 24755 -707
rect 24789 -741 24822 -707
rect 24722 -775 24822 -741
rect 24722 -809 24755 -775
rect 24789 -809 24822 -775
rect 24722 -843 24822 -809
rect 24722 -877 24755 -843
rect 24789 -877 24822 -843
rect 24722 -911 24822 -877
rect 24722 -945 24755 -911
rect 24789 -945 24822 -911
rect 24722 -979 24822 -945
rect 24722 -1013 24755 -979
rect 24789 -1013 24822 -979
rect 24722 -1047 24822 -1013
rect 24722 -1081 24755 -1047
rect 24789 -1081 24822 -1047
rect 24722 -1115 24822 -1081
rect 24722 -1149 24755 -1115
rect 24789 -1149 24822 -1115
rect 24722 -1183 24822 -1149
rect 24722 -1217 24755 -1183
rect 24789 -1217 24822 -1183
rect 24722 -1251 24822 -1217
rect 24722 -1285 24755 -1251
rect 24789 -1285 24822 -1251
rect 24722 -1319 24822 -1285
rect 24722 -1353 24755 -1319
rect 24789 -1353 24822 -1319
rect 24722 -1387 24822 -1353
rect 24722 -1421 24755 -1387
rect 24789 -1421 24822 -1387
rect 24722 -1455 24822 -1421
rect 24722 -1489 24755 -1455
rect 24789 -1489 24822 -1455
rect 24722 -1523 24822 -1489
rect 24722 -1557 24755 -1523
rect 24789 -1557 24822 -1523
rect 24722 -1591 24822 -1557
rect 24722 -1625 24755 -1591
rect 24789 -1625 24822 -1591
rect 24722 -1659 24822 -1625
rect 24722 -1693 24755 -1659
rect 24789 -1693 24822 -1659
rect 24722 -1727 24822 -1693
rect 24722 -1761 24755 -1727
rect 24789 -1761 24822 -1727
rect 24722 -1795 24822 -1761
rect 24722 -1829 24755 -1795
rect 24789 -1829 24822 -1795
rect 24722 -1863 24822 -1829
rect 24722 -1897 24755 -1863
rect 24789 -1897 24822 -1863
rect 24722 -1931 24822 -1897
rect 24722 -1965 24755 -1931
rect 24789 -1965 24822 -1931
rect 24722 -1999 24822 -1965
rect 24722 -2033 24755 -1999
rect 24789 -2033 24822 -1999
rect 24722 -2067 24822 -2033
rect 24722 -2101 24755 -2067
rect 24789 -2101 24822 -2067
rect 24722 -2135 24822 -2101
rect 24722 -2169 24755 -2135
rect 24789 -2169 24822 -2135
rect 24722 -2203 24822 -2169
rect 24722 -2237 24755 -2203
rect 24789 -2237 24822 -2203
rect 24722 -2271 24822 -2237
rect 24722 -2305 24755 -2271
rect 24789 -2305 24822 -2271
rect 24722 -2339 24822 -2305
rect 24722 -2373 24755 -2339
rect 24789 -2373 24822 -2339
rect 24722 -2407 24822 -2373
rect 24722 -2441 24755 -2407
rect 24789 -2441 24822 -2407
rect 24722 -2475 24822 -2441
rect 24722 -2509 24755 -2475
rect 24789 -2509 24822 -2475
rect 24722 -2543 24822 -2509
rect 24722 -2577 24755 -2543
rect 24789 -2577 24822 -2543
rect 24722 -2611 24822 -2577
rect 24722 -2645 24755 -2611
rect 24789 -2645 24822 -2611
rect 24722 -2679 24822 -2645
rect 24722 -2713 24755 -2679
rect 24789 -2713 24822 -2679
rect 24722 -2747 24822 -2713
rect 24722 -2781 24755 -2747
rect 24789 -2781 24822 -2747
rect 24722 -2815 24822 -2781
rect 24722 -2849 24755 -2815
rect 24789 -2849 24822 -2815
rect 24722 -2883 24822 -2849
rect 24722 -2917 24755 -2883
rect 24789 -2917 24822 -2883
rect 24722 -2951 24822 -2917
rect 24722 -2985 24755 -2951
rect 24789 -2985 24822 -2951
rect 24722 -3019 24822 -2985
rect 24722 -3053 24755 -3019
rect 24789 -3053 24822 -3019
rect 24722 -3087 24822 -3053
rect 24722 -3121 24755 -3087
rect 24789 -3121 24822 -3087
rect 24722 -3155 24822 -3121
rect 24722 -3189 24755 -3155
rect 24789 -3189 24822 -3155
rect 24722 -3223 24822 -3189
rect 24722 -3257 24755 -3223
rect 24789 -3257 24822 -3223
rect 24722 -3291 24822 -3257
rect 24722 -3325 24755 -3291
rect 24789 -3325 24822 -3291
rect 24722 -3359 24822 -3325
rect 24722 -3393 24755 -3359
rect 24789 -3393 24822 -3359
rect 24722 -3427 24822 -3393
rect 24722 -3461 24755 -3427
rect 24789 -3461 24822 -3427
rect 24722 -3495 24822 -3461
rect 24722 -3529 24755 -3495
rect 24789 -3529 24822 -3495
rect 24722 -3563 24822 -3529
rect 24722 -3597 24755 -3563
rect 24789 -3597 24822 -3563
rect 24722 -3631 24822 -3597
rect 24722 -3665 24755 -3631
rect 24789 -3665 24822 -3631
rect 24722 -3699 24822 -3665
rect 24722 -3733 24755 -3699
rect 24789 -3733 24822 -3699
rect 24722 -3767 24822 -3733
rect 24722 -3801 24755 -3767
rect 24789 -3801 24822 -3767
rect 24722 -3835 24822 -3801
rect 24722 -3869 24755 -3835
rect 24789 -3869 24822 -3835
rect 24722 -3903 24822 -3869
rect 24722 -3937 24755 -3903
rect 24789 -3937 24822 -3903
rect 24722 -3971 24822 -3937
rect 24722 -4005 24755 -3971
rect 24789 -4005 24822 -3971
rect 24722 -4039 24822 -4005
rect 24722 -4073 24755 -4039
rect 24789 -4073 24822 -4039
rect 24722 -4107 24822 -4073
rect 24722 -4141 24755 -4107
rect 24789 -4141 24822 -4107
rect 24722 -4175 24822 -4141
rect 24722 -4209 24755 -4175
rect 24789 -4209 24822 -4175
rect 24722 -4243 24822 -4209
rect 24722 -4277 24755 -4243
rect 24789 -4277 24822 -4243
rect 24722 -4311 24822 -4277
rect 24722 -4345 24755 -4311
rect 24789 -4345 24822 -4311
rect 24722 -4379 24822 -4345
rect 24722 -4413 24755 -4379
rect 24789 -4413 24822 -4379
rect 24722 -4447 24822 -4413
rect 24722 -4481 24755 -4447
rect 24789 -4481 24822 -4447
rect 24722 -4515 24822 -4481
rect 24722 -4549 24755 -4515
rect 24789 -4549 24822 -4515
rect 24722 -4583 24822 -4549
rect 378 -4651 478 -4617
rect 378 -4685 411 -4651
rect 445 -4685 478 -4651
rect 378 -4719 478 -4685
rect 24722 -4617 24755 -4583
rect 24789 -4617 24822 -4583
rect 24722 -4651 24822 -4617
rect 24722 -4685 24755 -4651
rect 24789 -4685 24822 -4651
rect 378 -4753 411 -4719
rect 445 -4753 478 -4719
rect 378 -4787 478 -4753
rect 378 -4821 411 -4787
rect 445 -4821 478 -4787
rect 378 -4855 478 -4821
rect 378 -4889 411 -4855
rect 445 -4889 478 -4855
rect 378 -4923 478 -4889
rect 378 -4957 411 -4923
rect 445 -4957 478 -4923
rect 378 -4991 478 -4957
rect 378 -5025 411 -4991
rect 445 -5025 478 -4991
rect 378 -5059 478 -5025
rect 378 -5093 411 -5059
rect 445 -5093 478 -5059
rect 24722 -4719 24822 -4685
rect 24722 -4753 24755 -4719
rect 24789 -4753 24822 -4719
rect 24722 -4787 24822 -4753
rect 24722 -4821 24755 -4787
rect 24789 -4821 24822 -4787
rect 24722 -4855 24822 -4821
rect 24722 -4889 24755 -4855
rect 24789 -4889 24822 -4855
rect 24722 -4923 24822 -4889
rect 24722 -4957 24755 -4923
rect 24789 -4957 24822 -4923
rect 24722 -4991 24822 -4957
rect 24722 -5025 24755 -4991
rect 24789 -5025 24822 -4991
rect 24722 -5059 24822 -5025
rect 378 -5127 478 -5093
rect 378 -5161 411 -5127
rect 445 -5161 478 -5127
rect 378 -5195 478 -5161
rect 24722 -5093 24755 -5059
rect 24789 -5093 24822 -5059
rect 24722 -5127 24822 -5093
rect 24722 -5161 24755 -5127
rect 24789 -5161 24822 -5127
rect 378 -5229 411 -5195
rect 445 -5229 478 -5195
rect 378 -5263 478 -5229
rect 378 -5297 411 -5263
rect 445 -5297 478 -5263
rect 378 -5331 478 -5297
rect 378 -5365 411 -5331
rect 445 -5365 478 -5331
rect 378 -5399 478 -5365
rect 378 -5433 411 -5399
rect 445 -5433 478 -5399
rect 378 -5467 478 -5433
rect 378 -5501 411 -5467
rect 445 -5501 478 -5467
rect 378 -5535 478 -5501
rect 24722 -5195 24822 -5161
rect 24722 -5229 24755 -5195
rect 24789 -5229 24822 -5195
rect 24722 -5263 24822 -5229
rect 24722 -5297 24755 -5263
rect 24789 -5297 24822 -5263
rect 24722 -5331 24822 -5297
rect 24722 -5365 24755 -5331
rect 24789 -5365 24822 -5331
rect 24722 -5399 24822 -5365
rect 24722 -5433 24755 -5399
rect 24789 -5433 24822 -5399
rect 24722 -5467 24822 -5433
rect 24722 -5501 24755 -5467
rect 24789 -5501 24822 -5467
rect 378 -5569 411 -5535
rect 445 -5569 478 -5535
rect 378 -5603 478 -5569
rect 378 -5637 411 -5603
rect 445 -5637 478 -5603
rect 24722 -5535 24822 -5501
rect 24722 -5569 24755 -5535
rect 24789 -5569 24822 -5535
rect 24722 -5603 24822 -5569
rect 378 -5671 478 -5637
rect 378 -5705 411 -5671
rect 445 -5705 478 -5671
rect 378 -5739 478 -5705
rect 378 -5773 411 -5739
rect 445 -5773 478 -5739
rect 378 -5807 478 -5773
rect 378 -5841 411 -5807
rect 445 -5841 478 -5807
rect 378 -5875 478 -5841
rect 378 -5909 411 -5875
rect 445 -5909 478 -5875
rect 378 -5943 478 -5909
rect 378 -5977 411 -5943
rect 445 -5977 478 -5943
rect 378 -6011 478 -5977
rect 378 -6045 411 -6011
rect 445 -6045 478 -6011
rect 24722 -5637 24755 -5603
rect 24789 -5637 24822 -5603
rect 24722 -5671 24822 -5637
rect 24722 -5705 24755 -5671
rect 24789 -5705 24822 -5671
rect 24722 -5739 24822 -5705
rect 24722 -5773 24755 -5739
rect 24789 -5773 24822 -5739
rect 24722 -5807 24822 -5773
rect 24722 -5841 24755 -5807
rect 24789 -5841 24822 -5807
rect 24722 -5875 24822 -5841
rect 24722 -5909 24755 -5875
rect 24789 -5909 24822 -5875
rect 24722 -5943 24822 -5909
rect 24722 -5977 24755 -5943
rect 24789 -5977 24822 -5943
rect 24722 -6011 24822 -5977
rect 378 -6079 478 -6045
rect 378 -6113 411 -6079
rect 445 -6113 478 -6079
rect 378 -6147 478 -6113
rect 24722 -6045 24755 -6011
rect 24789 -6045 24822 -6011
rect 24722 -6079 24822 -6045
rect 24722 -6113 24755 -6079
rect 24789 -6113 24822 -6079
rect 378 -6181 411 -6147
rect 445 -6181 478 -6147
rect 378 -6215 478 -6181
rect 378 -6249 411 -6215
rect 445 -6249 478 -6215
rect 378 -6283 478 -6249
rect 378 -6317 411 -6283
rect 445 -6317 478 -6283
rect 378 -6351 478 -6317
rect 378 -6385 411 -6351
rect 445 -6385 478 -6351
rect 378 -6419 478 -6385
rect 378 -6453 411 -6419
rect 445 -6453 478 -6419
rect 378 -6487 478 -6453
rect 24722 -6147 24822 -6113
rect 24722 -6181 24755 -6147
rect 24789 -6181 24822 -6147
rect 24722 -6215 24822 -6181
rect 24722 -6249 24755 -6215
rect 24789 -6249 24822 -6215
rect 24722 -6283 24822 -6249
rect 24722 -6317 24755 -6283
rect 24789 -6317 24822 -6283
rect 24722 -6351 24822 -6317
rect 24722 -6385 24755 -6351
rect 24789 -6385 24822 -6351
rect 24722 -6419 24822 -6385
rect 24722 -6453 24755 -6419
rect 24789 -6453 24822 -6419
rect 378 -6521 411 -6487
rect 445 -6521 478 -6487
rect 378 -6555 478 -6521
rect 378 -6589 411 -6555
rect 445 -6589 478 -6555
rect 24722 -6487 24822 -6453
rect 24722 -6521 24755 -6487
rect 24789 -6521 24822 -6487
rect 24722 -6555 24822 -6521
rect 378 -6623 478 -6589
rect 378 -6657 411 -6623
rect 445 -6657 478 -6623
rect 378 -6691 478 -6657
rect 378 -6725 411 -6691
rect 445 -6725 478 -6691
rect 378 -6759 478 -6725
rect 378 -6793 411 -6759
rect 445 -6793 478 -6759
rect 378 -6827 478 -6793
rect 378 -6861 411 -6827
rect 445 -6861 478 -6827
rect 378 -6895 478 -6861
rect 378 -6929 411 -6895
rect 445 -6929 478 -6895
rect 378 -6963 478 -6929
rect 378 -6997 411 -6963
rect 445 -6997 478 -6963
rect 24722 -6589 24755 -6555
rect 24789 -6589 24822 -6555
rect 24722 -6623 24822 -6589
rect 24722 -6657 24755 -6623
rect 24789 -6657 24822 -6623
rect 24722 -6691 24822 -6657
rect 24722 -6725 24755 -6691
rect 24789 -6725 24822 -6691
rect 24722 -6759 24822 -6725
rect 24722 -6793 24755 -6759
rect 24789 -6793 24822 -6759
rect 24722 -6827 24822 -6793
rect 24722 -6861 24755 -6827
rect 24789 -6861 24822 -6827
rect 24722 -6895 24822 -6861
rect 24722 -6929 24755 -6895
rect 24789 -6929 24822 -6895
rect 24722 -6963 24822 -6929
rect 378 -7031 478 -6997
rect 378 -7065 411 -7031
rect 445 -7065 478 -7031
rect 24722 -6997 24755 -6963
rect 24789 -6997 24822 -6963
rect 24722 -7031 24822 -6997
rect 378 -7099 478 -7065
rect 378 -7133 411 -7099
rect 445 -7133 478 -7099
rect 378 -7167 478 -7133
rect 378 -7201 411 -7167
rect 445 -7201 478 -7167
rect 378 -7235 478 -7201
rect 378 -7269 411 -7235
rect 445 -7269 478 -7235
rect 378 -7303 478 -7269
rect 378 -7337 411 -7303
rect 445 -7337 478 -7303
rect 378 -7371 478 -7337
rect 378 -7405 411 -7371
rect 445 -7405 478 -7371
rect 378 -7439 478 -7405
rect 24722 -7065 24755 -7031
rect 24789 -7065 24822 -7031
rect 24722 -7099 24822 -7065
rect 24722 -7133 24755 -7099
rect 24789 -7133 24822 -7099
rect 24722 -7167 24822 -7133
rect 24722 -7201 24755 -7167
rect 24789 -7201 24822 -7167
rect 24722 -7235 24822 -7201
rect 24722 -7269 24755 -7235
rect 24789 -7269 24822 -7235
rect 24722 -7303 24822 -7269
rect 24722 -7337 24755 -7303
rect 24789 -7337 24822 -7303
rect 24722 -7371 24822 -7337
rect 24722 -7405 24755 -7371
rect 24789 -7405 24822 -7371
rect 378 -7473 411 -7439
rect 445 -7473 478 -7439
rect 378 -7507 478 -7473
rect 24722 -7439 24822 -7405
rect 24722 -7473 24755 -7439
rect 24789 -7473 24822 -7439
rect 378 -7541 411 -7507
rect 445 -7541 478 -7507
rect 378 -7575 478 -7541
rect 378 -7609 411 -7575
rect 445 -7609 478 -7575
rect 378 -7643 478 -7609
rect 378 -7677 411 -7643
rect 445 -7677 478 -7643
rect 378 -7711 478 -7677
rect 378 -7745 411 -7711
rect 445 -7745 478 -7711
rect 378 -7779 478 -7745
rect 378 -7813 411 -7779
rect 445 -7813 478 -7779
rect 378 -7847 478 -7813
rect 378 -7881 411 -7847
rect 445 -7881 478 -7847
rect 378 -7915 478 -7881
rect 24722 -7507 24822 -7473
rect 24722 -7541 24755 -7507
rect 24789 -7541 24822 -7507
rect 24722 -7575 24822 -7541
rect 24722 -7609 24755 -7575
rect 24789 -7609 24822 -7575
rect 24722 -7643 24822 -7609
rect 24722 -7677 24755 -7643
rect 24789 -7677 24822 -7643
rect 24722 -7711 24822 -7677
rect 24722 -7745 24755 -7711
rect 24789 -7745 24822 -7711
rect 24722 -7779 24822 -7745
rect 24722 -7813 24755 -7779
rect 24789 -7813 24822 -7779
rect 24722 -7847 24822 -7813
rect 24722 -7881 24755 -7847
rect 24789 -7881 24822 -7847
rect 378 -7949 411 -7915
rect 445 -7949 478 -7915
rect 378 -7983 478 -7949
rect 378 -8017 411 -7983
rect 445 -8017 478 -7983
rect 24722 -7915 24822 -7881
rect 24722 -7949 24755 -7915
rect 24789 -7949 24822 -7915
rect 24722 -7983 24822 -7949
rect 378 -8051 478 -8017
rect 378 -8085 411 -8051
rect 445 -8085 478 -8051
rect 378 -8119 478 -8085
rect 378 -8153 411 -8119
rect 445 -8153 478 -8119
rect 378 -8187 478 -8153
rect 378 -8221 411 -8187
rect 445 -8221 478 -8187
rect 378 -8255 478 -8221
rect 378 -8289 411 -8255
rect 445 -8289 478 -8255
rect 378 -8323 478 -8289
rect 378 -8357 411 -8323
rect 445 -8357 478 -8323
rect 378 -8391 478 -8357
rect 378 -8425 411 -8391
rect 445 -8425 478 -8391
rect 378 -8459 478 -8425
rect 378 -8493 411 -8459
rect 445 -8493 478 -8459
rect 378 -8527 478 -8493
rect 378 -8561 411 -8527
rect 445 -8561 478 -8527
rect 378 -8595 478 -8561
rect 378 -8629 411 -8595
rect 445 -8629 478 -8595
rect 378 -8663 478 -8629
rect 378 -8697 411 -8663
rect 445 -8697 478 -8663
rect 378 -8782 478 -8697
rect 24722 -8017 24755 -7983
rect 24789 -8017 24822 -7983
rect 24722 -8051 24822 -8017
rect 24722 -8085 24755 -8051
rect 24789 -8085 24822 -8051
rect 24722 -8119 24822 -8085
rect 24722 -8153 24755 -8119
rect 24789 -8153 24822 -8119
rect 24722 -8187 24822 -8153
rect 24722 -8221 24755 -8187
rect 24789 -8221 24822 -8187
rect 24722 -8255 24822 -8221
rect 24722 -8289 24755 -8255
rect 24789 -8289 24822 -8255
rect 24722 -8323 24822 -8289
rect 24722 -8357 24755 -8323
rect 24789 -8357 24822 -8323
rect 24722 -8391 24822 -8357
rect 24722 -8425 24755 -8391
rect 24789 -8425 24822 -8391
rect 24722 -8459 24822 -8425
rect 24722 -8493 24755 -8459
rect 24789 -8493 24822 -8459
rect 24722 -8527 24822 -8493
rect 24722 -8561 24755 -8527
rect 24789 -8561 24822 -8527
rect 24722 -8595 24822 -8561
rect 24722 -8629 24755 -8595
rect 24789 -8629 24822 -8595
rect 24722 -8663 24822 -8629
rect 24722 -8697 24755 -8663
rect 24789 -8697 24822 -8663
rect 24722 -8782 24822 -8697
rect 378 -8815 24822 -8782
rect 378 -8849 547 -8815
rect 581 -8849 615 -8815
rect 649 -8849 683 -8815
rect 717 -8849 751 -8815
rect 785 -8849 819 -8815
rect 853 -8849 887 -8815
rect 921 -8849 955 -8815
rect 989 -8849 1023 -8815
rect 1057 -8849 1091 -8815
rect 1125 -8849 1159 -8815
rect 1193 -8849 1227 -8815
rect 1261 -8849 1295 -8815
rect 1329 -8849 1363 -8815
rect 1397 -8849 1431 -8815
rect 1465 -8849 1499 -8815
rect 1533 -8849 1567 -8815
rect 1601 -8849 1635 -8815
rect 1669 -8849 1703 -8815
rect 1737 -8849 1771 -8815
rect 1805 -8849 1839 -8815
rect 1873 -8849 1907 -8815
rect 1941 -8849 1975 -8815
rect 2009 -8849 2043 -8815
rect 2077 -8849 2111 -8815
rect 2145 -8849 2179 -8815
rect 2213 -8849 2247 -8815
rect 2281 -8849 2315 -8815
rect 2349 -8849 2383 -8815
rect 2417 -8849 2451 -8815
rect 2485 -8849 2519 -8815
rect 2553 -8849 2587 -8815
rect 2621 -8849 2655 -8815
rect 2689 -8849 2723 -8815
rect 2757 -8849 2791 -8815
rect 2825 -8849 2859 -8815
rect 2893 -8849 2927 -8815
rect 2961 -8849 2995 -8815
rect 3029 -8849 3063 -8815
rect 3097 -8849 3131 -8815
rect 3165 -8849 3199 -8815
rect 3233 -8849 3267 -8815
rect 3301 -8849 3335 -8815
rect 3369 -8849 3403 -8815
rect 3437 -8849 3471 -8815
rect 3505 -8849 3539 -8815
rect 3573 -8849 3607 -8815
rect 3641 -8849 3675 -8815
rect 3709 -8849 3743 -8815
rect 3777 -8849 3811 -8815
rect 3845 -8849 3879 -8815
rect 3913 -8849 3947 -8815
rect 3981 -8849 4015 -8815
rect 4049 -8849 4083 -8815
rect 4117 -8849 4151 -8815
rect 4185 -8849 4219 -8815
rect 4253 -8849 4287 -8815
rect 4321 -8849 4355 -8815
rect 4389 -8849 4423 -8815
rect 4457 -8849 4491 -8815
rect 4525 -8849 4559 -8815
rect 4593 -8849 4627 -8815
rect 4661 -8849 4695 -8815
rect 4729 -8849 4763 -8815
rect 4797 -8849 4831 -8815
rect 4865 -8849 4899 -8815
rect 4933 -8849 4967 -8815
rect 5001 -8849 5035 -8815
rect 5069 -8849 5103 -8815
rect 5137 -8849 5171 -8815
rect 5205 -8849 5239 -8815
rect 5273 -8849 5307 -8815
rect 5341 -8849 5375 -8815
rect 5409 -8849 5443 -8815
rect 5477 -8849 5511 -8815
rect 5545 -8849 5579 -8815
rect 5613 -8849 5647 -8815
rect 5681 -8849 5715 -8815
rect 5749 -8849 5783 -8815
rect 5817 -8849 5851 -8815
rect 5885 -8849 5919 -8815
rect 5953 -8849 5987 -8815
rect 6021 -8849 6055 -8815
rect 6089 -8849 6123 -8815
rect 6157 -8849 6191 -8815
rect 6225 -8849 6259 -8815
rect 6293 -8849 6327 -8815
rect 6361 -8849 6395 -8815
rect 6429 -8849 6463 -8815
rect 6497 -8849 6531 -8815
rect 6565 -8849 6599 -8815
rect 6633 -8849 6667 -8815
rect 6701 -8849 6735 -8815
rect 6769 -8849 6803 -8815
rect 6837 -8849 6871 -8815
rect 6905 -8849 6939 -8815
rect 6973 -8849 7007 -8815
rect 7041 -8849 7075 -8815
rect 7109 -8849 7143 -8815
rect 7177 -8849 7211 -8815
rect 7245 -8849 7279 -8815
rect 7313 -8849 7347 -8815
rect 7381 -8849 7415 -8815
rect 7449 -8849 7483 -8815
rect 7517 -8849 7551 -8815
rect 7585 -8849 7619 -8815
rect 7653 -8849 7687 -8815
rect 7721 -8849 7755 -8815
rect 7789 -8849 7823 -8815
rect 7857 -8849 7891 -8815
rect 7925 -8849 7959 -8815
rect 7993 -8849 8027 -8815
rect 8061 -8849 8095 -8815
rect 8129 -8849 8163 -8815
rect 8197 -8849 8231 -8815
rect 8265 -8849 8299 -8815
rect 8333 -8849 8367 -8815
rect 8401 -8849 8435 -8815
rect 8469 -8849 8503 -8815
rect 8537 -8849 8571 -8815
rect 8605 -8849 8639 -8815
rect 8673 -8849 8707 -8815
rect 8741 -8849 8775 -8815
rect 8809 -8849 8843 -8815
rect 8877 -8849 8911 -8815
rect 8945 -8849 8979 -8815
rect 9013 -8849 9047 -8815
rect 9081 -8849 9115 -8815
rect 9149 -8849 9183 -8815
rect 9217 -8849 9251 -8815
rect 9285 -8849 9319 -8815
rect 9353 -8849 9387 -8815
rect 9421 -8849 9455 -8815
rect 9489 -8849 9523 -8815
rect 9557 -8849 9591 -8815
rect 9625 -8849 9659 -8815
rect 9693 -8849 9727 -8815
rect 9761 -8849 9795 -8815
rect 9829 -8849 9863 -8815
rect 9897 -8849 9931 -8815
rect 9965 -8849 9999 -8815
rect 10033 -8849 10067 -8815
rect 10101 -8849 10135 -8815
rect 10169 -8849 10203 -8815
rect 10237 -8849 10271 -8815
rect 10305 -8849 10339 -8815
rect 10373 -8849 10407 -8815
rect 10441 -8849 10475 -8815
rect 10509 -8849 10543 -8815
rect 10577 -8849 10611 -8815
rect 10645 -8849 10679 -8815
rect 10713 -8849 10747 -8815
rect 10781 -8849 10815 -8815
rect 10849 -8849 10883 -8815
rect 10917 -8849 10951 -8815
rect 10985 -8849 11019 -8815
rect 11053 -8849 11087 -8815
rect 11121 -8849 11155 -8815
rect 11189 -8849 11223 -8815
rect 11257 -8849 11291 -8815
rect 11325 -8849 11359 -8815
rect 11393 -8849 11427 -8815
rect 11461 -8849 11495 -8815
rect 11529 -8849 11563 -8815
rect 11597 -8849 11631 -8815
rect 11665 -8849 11699 -8815
rect 11733 -8849 11767 -8815
rect 11801 -8849 11835 -8815
rect 11869 -8849 11903 -8815
rect 11937 -8849 11971 -8815
rect 12005 -8849 12039 -8815
rect 12073 -8849 12107 -8815
rect 12141 -8849 12175 -8815
rect 12209 -8849 12243 -8815
rect 12277 -8849 12311 -8815
rect 12345 -8849 12379 -8815
rect 12413 -8849 12447 -8815
rect 12481 -8849 12515 -8815
rect 12549 -8849 12583 -8815
rect 12617 -8849 12651 -8815
rect 12685 -8849 12719 -8815
rect 12753 -8849 12787 -8815
rect 12821 -8849 12855 -8815
rect 12889 -8849 12923 -8815
rect 12957 -8849 12991 -8815
rect 13025 -8849 13059 -8815
rect 13093 -8849 13127 -8815
rect 13161 -8849 13195 -8815
rect 13229 -8849 13263 -8815
rect 13297 -8849 13331 -8815
rect 13365 -8849 13399 -8815
rect 13433 -8849 13467 -8815
rect 13501 -8849 13535 -8815
rect 13569 -8849 13603 -8815
rect 13637 -8849 13671 -8815
rect 13705 -8849 13739 -8815
rect 13773 -8849 13807 -8815
rect 13841 -8849 13875 -8815
rect 13909 -8849 13943 -8815
rect 13977 -8849 14011 -8815
rect 14045 -8849 14079 -8815
rect 14113 -8849 14147 -8815
rect 14181 -8849 14215 -8815
rect 14249 -8849 14283 -8815
rect 14317 -8849 14351 -8815
rect 14385 -8849 14419 -8815
rect 14453 -8849 14487 -8815
rect 14521 -8849 14555 -8815
rect 14589 -8849 14623 -8815
rect 14657 -8849 14691 -8815
rect 14725 -8849 14759 -8815
rect 14793 -8849 14827 -8815
rect 14861 -8849 14895 -8815
rect 14929 -8849 14963 -8815
rect 14997 -8849 15031 -8815
rect 15065 -8849 15099 -8815
rect 15133 -8849 15167 -8815
rect 15201 -8849 15235 -8815
rect 15269 -8849 15303 -8815
rect 15337 -8849 15371 -8815
rect 15405 -8849 15439 -8815
rect 15473 -8849 15507 -8815
rect 15541 -8849 15575 -8815
rect 15609 -8849 15643 -8815
rect 15677 -8849 15711 -8815
rect 15745 -8849 15779 -8815
rect 15813 -8849 15847 -8815
rect 15881 -8849 15915 -8815
rect 15949 -8849 15983 -8815
rect 16017 -8849 16051 -8815
rect 16085 -8849 16119 -8815
rect 16153 -8849 16187 -8815
rect 16221 -8849 16255 -8815
rect 16289 -8849 16323 -8815
rect 16357 -8849 16391 -8815
rect 16425 -8849 16459 -8815
rect 16493 -8849 16527 -8815
rect 16561 -8849 16595 -8815
rect 16629 -8849 16663 -8815
rect 16697 -8849 16731 -8815
rect 16765 -8849 16799 -8815
rect 16833 -8849 16867 -8815
rect 16901 -8849 16935 -8815
rect 16969 -8849 17003 -8815
rect 17037 -8849 17071 -8815
rect 17105 -8849 17139 -8815
rect 17173 -8849 17207 -8815
rect 17241 -8849 17275 -8815
rect 17309 -8849 17343 -8815
rect 17377 -8849 17411 -8815
rect 17445 -8849 17479 -8815
rect 17513 -8849 17547 -8815
rect 17581 -8849 17615 -8815
rect 17649 -8849 17683 -8815
rect 17717 -8849 17751 -8815
rect 17785 -8849 17819 -8815
rect 17853 -8849 17887 -8815
rect 17921 -8849 17955 -8815
rect 17989 -8849 18023 -8815
rect 18057 -8849 18091 -8815
rect 18125 -8849 18159 -8815
rect 18193 -8849 18227 -8815
rect 18261 -8849 18295 -8815
rect 18329 -8849 18363 -8815
rect 18397 -8849 18431 -8815
rect 18465 -8849 18499 -8815
rect 18533 -8849 18567 -8815
rect 18601 -8849 18635 -8815
rect 18669 -8849 18703 -8815
rect 18737 -8849 18771 -8815
rect 18805 -8849 18839 -8815
rect 18873 -8849 18907 -8815
rect 18941 -8849 18975 -8815
rect 19009 -8849 19043 -8815
rect 19077 -8849 19111 -8815
rect 19145 -8849 19179 -8815
rect 19213 -8849 19247 -8815
rect 19281 -8849 19315 -8815
rect 19349 -8849 19383 -8815
rect 19417 -8849 19451 -8815
rect 19485 -8849 19519 -8815
rect 19553 -8849 19587 -8815
rect 19621 -8849 19655 -8815
rect 19689 -8849 19723 -8815
rect 19757 -8849 19791 -8815
rect 19825 -8849 19859 -8815
rect 19893 -8849 19927 -8815
rect 19961 -8849 19995 -8815
rect 20029 -8849 20063 -8815
rect 20097 -8849 20131 -8815
rect 20165 -8849 20199 -8815
rect 20233 -8849 20267 -8815
rect 20301 -8849 20335 -8815
rect 20369 -8849 20403 -8815
rect 20437 -8849 20471 -8815
rect 20505 -8849 20539 -8815
rect 20573 -8849 20607 -8815
rect 20641 -8849 20675 -8815
rect 20709 -8849 20743 -8815
rect 20777 -8849 20811 -8815
rect 20845 -8849 20879 -8815
rect 20913 -8849 20947 -8815
rect 20981 -8849 21015 -8815
rect 21049 -8849 21083 -8815
rect 21117 -8849 21151 -8815
rect 21185 -8849 21219 -8815
rect 21253 -8849 21287 -8815
rect 21321 -8849 21355 -8815
rect 21389 -8849 21423 -8815
rect 21457 -8849 21491 -8815
rect 21525 -8849 21559 -8815
rect 21593 -8849 21627 -8815
rect 21661 -8849 21695 -8815
rect 21729 -8849 21763 -8815
rect 21797 -8849 21831 -8815
rect 21865 -8849 21899 -8815
rect 21933 -8849 21967 -8815
rect 22001 -8849 22035 -8815
rect 22069 -8849 22103 -8815
rect 22137 -8849 22171 -8815
rect 22205 -8849 22239 -8815
rect 22273 -8849 22307 -8815
rect 22341 -8849 22375 -8815
rect 22409 -8849 22443 -8815
rect 22477 -8849 22511 -8815
rect 22545 -8849 22579 -8815
rect 22613 -8849 22647 -8815
rect 22681 -8849 22715 -8815
rect 22749 -8849 22783 -8815
rect 22817 -8849 22851 -8815
rect 22885 -8849 22919 -8815
rect 22953 -8849 22987 -8815
rect 23021 -8849 23055 -8815
rect 23089 -8849 23123 -8815
rect 23157 -8849 23191 -8815
rect 23225 -8849 23259 -8815
rect 23293 -8849 23327 -8815
rect 23361 -8849 23395 -8815
rect 23429 -8849 23463 -8815
rect 23497 -8849 23531 -8815
rect 23565 -8849 23599 -8815
rect 23633 -8849 23667 -8815
rect 23701 -8849 23735 -8815
rect 23769 -8849 23803 -8815
rect 23837 -8849 23871 -8815
rect 23905 -8849 23939 -8815
rect 23973 -8849 24007 -8815
rect 24041 -8849 24075 -8815
rect 24109 -8849 24143 -8815
rect 24177 -8849 24211 -8815
rect 24245 -8849 24279 -8815
rect 24313 -8849 24347 -8815
rect 24381 -8849 24415 -8815
rect 24449 -8849 24483 -8815
rect 24517 -8849 24551 -8815
rect 24585 -8849 24619 -8815
rect 24653 -8849 24822 -8815
rect 378 -8882 24822 -8849
<< psubdiffcont >>
rect -12145 -11245 -12111 -11211
rect -12077 -11245 -12043 -11211
rect -12009 -11245 -11975 -11211
rect -11941 -11245 -11907 -11211
rect -11873 -11245 -11839 -11211
rect -11805 -11245 -11771 -11211
rect -11737 -11245 -11703 -11211
rect -11669 -11245 -11635 -11211
rect -11601 -11245 -11567 -11211
rect -11533 -11245 -11499 -11211
rect -11465 -11245 -11431 -11211
rect -11397 -11245 -11363 -11211
rect -11329 -11245 -11295 -11211
rect -11261 -11245 -11227 -11211
rect -11193 -11245 -11159 -11211
rect -11125 -11245 -11091 -11211
rect -11057 -11245 -11023 -11211
rect -10989 -11245 -10955 -11211
rect -10921 -11245 -10887 -11211
rect -10853 -11245 -10819 -11211
rect -10785 -11245 -10751 -11211
rect -10717 -11245 -10683 -11211
rect -10649 -11245 -10615 -11211
rect -10581 -11245 -10547 -11211
rect -10513 -11245 -10479 -11211
rect -10445 -11245 -10411 -11211
rect -10377 -11245 -10343 -11211
rect -10309 -11245 -10275 -11211
rect -10241 -11245 -10207 -11211
rect -10173 -11245 -10139 -11211
rect -10105 -11245 -10071 -11211
rect -10037 -11245 -10003 -11211
rect -9969 -11245 -9935 -11211
rect -9901 -11245 -9867 -11211
rect -9833 -11245 -9799 -11211
rect -9765 -11245 -9731 -11211
rect -9697 -11245 -9663 -11211
rect -9629 -11245 -9595 -11211
rect -9561 -11245 -9527 -11211
rect -9493 -11245 -9459 -11211
rect -9425 -11245 -9391 -11211
rect -9357 -11245 -9323 -11211
rect -9289 -11245 -9255 -11211
rect -9221 -11245 -9187 -11211
rect -9153 -11245 -9119 -11211
rect -9085 -11245 -9051 -11211
rect -9017 -11245 -8983 -11211
rect -8949 -11245 -8915 -11211
rect -8881 -11245 -8847 -11211
rect -8813 -11245 -8779 -11211
rect -8745 -11245 -8711 -11211
rect -8677 -11245 -8643 -11211
rect -8609 -11245 -8575 -11211
rect -8541 -11245 -8507 -11211
rect -8473 -11245 -8439 -11211
rect -8405 -11245 -8371 -11211
rect -8337 -11245 -8303 -11211
rect -8269 -11245 -8235 -11211
rect -8201 -11245 -8167 -11211
rect -8133 -11245 -8099 -11211
rect -8065 -11245 -8031 -11211
rect -7997 -11245 -7963 -11211
rect -7929 -11245 -7895 -11211
rect -7861 -11245 -7827 -11211
rect -7793 -11245 -7759 -11211
rect -7725 -11245 -7691 -11211
rect -7657 -11245 -7623 -11211
rect -7589 -11245 -7555 -11211
rect -7521 -11245 -7487 -11211
rect -7453 -11245 -7419 -11211
rect -7385 -11245 -7351 -11211
rect -7317 -11245 -7283 -11211
rect -7249 -11245 -7215 -11211
rect -7181 -11245 -7147 -11211
rect -7113 -11245 -7079 -11211
rect -7045 -11245 -7011 -11211
rect -6977 -11245 -6943 -11211
rect -6909 -11245 -6875 -11211
rect -6841 -11245 -6807 -11211
rect -6773 -11245 -6739 -11211
rect -6705 -11245 -6671 -11211
rect -6637 -11245 -6603 -11211
rect -6569 -11245 -6535 -11211
rect -6501 -11245 -6467 -11211
rect -6433 -11245 -6399 -11211
rect -6365 -11245 -6331 -11211
rect -6297 -11245 -6263 -11211
rect -6229 -11245 -6195 -11211
rect -6161 -11245 -6127 -11211
rect -6093 -11245 -6059 -11211
rect -6025 -11245 -5991 -11211
rect -5957 -11245 -5923 -11211
rect -5889 -11245 -5855 -11211
rect -5821 -11245 -5787 -11211
rect -5753 -11245 -5719 -11211
rect -5685 -11245 -5651 -11211
rect -5617 -11245 -5583 -11211
rect -5549 -11245 -5515 -11211
rect -5481 -11245 -5447 -11211
rect -5413 -11245 -5379 -11211
rect -5345 -11245 -5311 -11211
rect -5277 -11245 -5243 -11211
rect -5209 -11245 -5175 -11211
rect -5141 -11245 -5107 -11211
rect -5073 -11245 -5039 -11211
rect -5005 -11245 -4971 -11211
rect -4937 -11245 -4903 -11211
rect -4869 -11245 -4835 -11211
rect -4801 -11245 -4767 -11211
rect -4733 -11245 -4699 -11211
rect -4665 -11245 -4631 -11211
rect -4597 -11245 -4563 -11211
rect -4529 -11245 -4495 -11211
rect -4461 -11245 -4427 -11211
rect -4393 -11245 -4359 -11211
rect -4325 -11245 -4291 -11211
rect -4257 -11245 -4223 -11211
rect -4189 -11245 -4155 -11211
rect -4121 -11245 -4087 -11211
rect -4053 -11245 -4019 -11211
rect -3985 -11245 -3951 -11211
rect -3917 -11245 -3883 -11211
rect -3849 -11245 -3815 -11211
rect -3781 -11245 -3747 -11211
rect -3713 -11245 -3679 -11211
rect -3645 -11245 -3611 -11211
rect -3577 -11245 -3543 -11211
rect -3509 -11245 -3475 -11211
rect -3441 -11245 -3407 -11211
rect -3373 -11245 -3339 -11211
rect -3305 -11245 -3271 -11211
rect -3237 -11245 -3203 -11211
rect -3169 -11245 -3135 -11211
rect -3101 -11245 -3067 -11211
rect -3033 -11245 -2999 -11211
rect -2965 -11245 -2931 -11211
rect -2897 -11245 -2863 -11211
rect -2829 -11245 -2795 -11211
rect -2761 -11245 -2727 -11211
rect -2693 -11245 -2659 -11211
rect -2625 -11245 -2591 -11211
rect -2557 -11245 -2523 -11211
rect -2489 -11245 -2455 -11211
rect -2421 -11245 -2387 -11211
rect -2353 -11245 -2319 -11211
rect -2285 -11245 -2251 -11211
rect -2217 -11245 -2183 -11211
rect -2149 -11245 -2115 -11211
rect -2081 -11245 -2047 -11211
rect -2013 -11245 -1979 -11211
rect -1945 -11245 -1911 -11211
rect -1877 -11245 -1843 -11211
rect -1809 -11245 -1775 -11211
rect -1741 -11245 -1707 -11211
rect -1673 -11245 -1639 -11211
rect -1605 -11245 -1571 -11211
rect -1537 -11245 -1503 -11211
rect -1469 -11245 -1435 -11211
rect -1401 -11245 -1367 -11211
rect -1333 -11245 -1299 -11211
rect -1265 -11245 -1231 -11211
rect -1197 -11245 -1163 -11211
rect -1129 -11245 -1095 -11211
rect -1061 -11245 -1027 -11211
rect -993 -11245 -959 -11211
rect -925 -11245 -891 -11211
rect -857 -11245 -823 -11211
rect -789 -11245 -755 -11211
rect -721 -11245 -687 -11211
rect -653 -11245 -619 -11211
rect -585 -11245 -551 -11211
rect -517 -11245 -483 -11211
rect -449 -11245 -415 -11211
rect -381 -11245 -347 -11211
rect -313 -11245 -279 -11211
rect -245 -11245 -211 -11211
rect -177 -11245 -143 -11211
rect -109 -11245 -75 -11211
rect -41 -11245 -7 -11211
rect 27 -11245 61 -11211
rect 95 -11245 129 -11211
rect 163 -11245 197 -11211
rect 231 -11245 265 -11211
rect 299 -11245 333 -11211
rect 367 -11245 401 -11211
rect 435 -11245 469 -11211
rect 503 -11245 537 -11211
rect 571 -11245 605 -11211
rect 639 -11245 673 -11211
rect 707 -11245 741 -11211
rect 775 -11245 809 -11211
rect 843 -11245 877 -11211
rect 911 -11245 945 -11211
rect 979 -11245 1013 -11211
rect 1047 -11245 1081 -11211
rect 1115 -11245 1149 -11211
rect 1183 -11245 1217 -11211
rect 1251 -11245 1285 -11211
rect 1319 -11245 1353 -11211
rect 1387 -11245 1421 -11211
rect 1455 -11245 1489 -11211
rect 1523 -11245 1557 -11211
rect 1591 -11245 1625 -11211
rect 1659 -11245 1693 -11211
rect 1727 -11245 1761 -11211
rect 1795 -11245 1829 -11211
rect 1863 -11245 1897 -11211
rect 1931 -11245 1965 -11211
rect 1999 -11245 2033 -11211
rect 2067 -11245 2101 -11211
rect 2135 -11245 2169 -11211
rect 2203 -11245 2237 -11211
rect 2271 -11245 2305 -11211
rect 2339 -11245 2373 -11211
rect 2407 -11245 2441 -11211
rect 2475 -11245 2509 -11211
rect 2543 -11245 2577 -11211
rect 2611 -11245 2645 -11211
rect 2679 -11245 2713 -11211
rect 2747 -11245 2781 -11211
rect 2815 -11245 2849 -11211
rect 2883 -11245 2917 -11211
rect 2951 -11245 2985 -11211
rect 3019 -11245 3053 -11211
rect 3087 -11245 3121 -11211
rect 3155 -11245 3189 -11211
rect 3223 -11245 3257 -11211
rect 3291 -11245 3325 -11211
rect 3359 -11245 3393 -11211
rect 3427 -11245 3461 -11211
rect 3495 -11245 3529 -11211
rect 3563 -11245 3597 -11211
rect 3631 -11245 3665 -11211
rect 3699 -11245 3733 -11211
rect 3767 -11245 3801 -11211
rect 3835 -11245 3869 -11211
rect 3903 -11245 3937 -11211
rect 3971 -11245 4005 -11211
rect 4039 -11245 4073 -11211
rect 4107 -11245 4141 -11211
rect 4175 -11245 4209 -11211
rect 4243 -11245 4277 -11211
rect 4311 -11245 4345 -11211
rect 4379 -11245 4413 -11211
rect 4447 -11245 4481 -11211
rect 4515 -11245 4549 -11211
rect 4583 -11245 4617 -11211
rect 4651 -11245 4685 -11211
rect 4719 -11245 4753 -11211
rect 4787 -11245 4821 -11211
rect 4855 -11245 4889 -11211
rect 4923 -11245 4957 -11211
rect 4991 -11245 5025 -11211
rect 5059 -11245 5093 -11211
rect 5127 -11245 5161 -11211
rect 5195 -11245 5229 -11211
rect 5263 -11245 5297 -11211
rect 5331 -11245 5365 -11211
rect 5399 -11245 5433 -11211
rect 5467 -11245 5501 -11211
rect 5535 -11245 5569 -11211
rect 5603 -11245 5637 -11211
rect 5671 -11245 5705 -11211
rect 5739 -11245 5773 -11211
rect 5807 -11245 5841 -11211
rect 5875 -11245 5909 -11211
rect 5943 -11245 5977 -11211
rect 6011 -11245 6045 -11211
rect 6079 -11245 6113 -11211
rect 6147 -11245 6181 -11211
rect 6215 -11245 6249 -11211
rect 6283 -11245 6317 -11211
rect 6351 -11245 6385 -11211
rect 6419 -11245 6453 -11211
rect 6487 -11245 6521 -11211
rect 6555 -11245 6589 -11211
rect 6623 -11245 6657 -11211
rect 6691 -11245 6725 -11211
rect 6759 -11245 6793 -11211
rect 6827 -11245 6861 -11211
rect 6895 -11245 6929 -11211
rect 6963 -11245 6997 -11211
rect 7031 -11245 7065 -11211
rect 7099 -11245 7133 -11211
rect 7167 -11245 7201 -11211
rect 7235 -11245 7269 -11211
rect 7303 -11245 7337 -11211
rect 7371 -11245 7405 -11211
rect 7439 -11245 7473 -11211
rect 7507 -11245 7541 -11211
rect 7575 -11245 7609 -11211
rect 7643 -11245 7677 -11211
rect 7711 -11245 7745 -11211
rect 7779 -11245 7813 -11211
rect 7847 -11245 7881 -11211
rect 7915 -11245 7949 -11211
rect 7983 -11245 8017 -11211
rect 8051 -11245 8085 -11211
rect 8119 -11245 8153 -11211
rect 8187 -11245 8221 -11211
rect 8255 -11245 8289 -11211
rect 8323 -11245 8357 -11211
rect 8391 -11245 8425 -11211
rect 8459 -11245 8493 -11211
rect 8527 -11245 8561 -11211
rect 8595 -11245 8629 -11211
rect 8663 -11245 8697 -11211
rect 8731 -11245 8765 -11211
rect 8799 -11245 8833 -11211
rect 8867 -11245 8901 -11211
rect 8935 -11245 8969 -11211
rect 9003 -11245 9037 -11211
rect 9071 -11245 9105 -11211
rect 9139 -11245 9173 -11211
rect 9207 -11245 9241 -11211
rect 9275 -11245 9309 -11211
rect 9343 -11245 9377 -11211
rect 9411 -11245 9445 -11211
rect 9479 -11245 9513 -11211
rect 9547 -11245 9581 -11211
rect 9615 -11245 9649 -11211
rect 9683 -11245 9717 -11211
rect 9751 -11245 9785 -11211
rect 9819 -11245 9853 -11211
rect 9887 -11245 9921 -11211
rect 9955 -11245 9989 -11211
rect 10023 -11245 10057 -11211
rect 10091 -11245 10125 -11211
rect 10159 -11245 10193 -11211
rect 10227 -11245 10261 -11211
rect 10295 -11245 10329 -11211
rect 10363 -11245 10397 -11211
rect 10431 -11245 10465 -11211
rect 10499 -11245 10533 -11211
rect 10567 -11245 10601 -11211
rect 10635 -11245 10669 -11211
rect 10703 -11245 10737 -11211
rect 10771 -11245 10805 -11211
rect 10839 -11245 10873 -11211
rect 10907 -11245 10941 -11211
rect 10975 -11245 11009 -11211
rect 11043 -11245 11077 -11211
rect 11111 -11245 11145 -11211
rect 11179 -11245 11213 -11211
rect 11247 -11245 11281 -11211
rect 11315 -11245 11349 -11211
rect 11383 -11245 11417 -11211
rect 11451 -11245 11485 -11211
rect 11519 -11245 11553 -11211
rect 11587 -11245 11621 -11211
rect 11655 -11245 11689 -11211
rect 11723 -11245 11757 -11211
rect 11791 -11245 11825 -11211
rect 11859 -11245 11893 -11211
rect 11927 -11245 11961 -11211
rect 11995 -11245 12029 -11211
rect 12063 -11245 12097 -11211
rect 12131 -11245 12165 -11211
rect 12199 -11245 12233 -11211
rect 12267 -11245 12301 -11211
rect 12335 -11245 12369 -11211
rect 12403 -11245 12437 -11211
rect 12471 -11245 12505 -11211
rect 12539 -11245 12573 -11211
rect 12607 -11245 12641 -11211
rect 12675 -11245 12709 -11211
rect 12743 -11245 12777 -11211
rect 12811 -11245 12845 -11211
rect 12879 -11245 12913 -11211
rect 12947 -11245 12981 -11211
rect 13015 -11245 13049 -11211
rect 13083 -11245 13117 -11211
rect 13151 -11245 13185 -11211
rect 13219 -11245 13253 -11211
rect 13287 -11245 13321 -11211
rect 13355 -11245 13389 -11211
rect 13423 -11245 13457 -11211
rect 13491 -11245 13525 -11211
rect 13559 -11245 13593 -11211
rect 13627 -11245 13661 -11211
rect 13695 -11245 13729 -11211
rect 13763 -11245 13797 -11211
rect 13831 -11245 13865 -11211
rect 13899 -11245 13933 -11211
rect 13967 -11245 14001 -11211
rect 14035 -11245 14069 -11211
rect 14103 -11245 14137 -11211
rect 14171 -11245 14205 -11211
rect 14239 -11245 14273 -11211
rect 14307 -11245 14341 -11211
rect 14375 -11245 14409 -11211
rect 14443 -11245 14477 -11211
rect 14511 -11245 14545 -11211
rect 14579 -11245 14613 -11211
rect 14647 -11245 14681 -11211
rect 14715 -11245 14749 -11211
rect 14783 -11245 14817 -11211
rect 14851 -11245 14885 -11211
rect 14919 -11245 14953 -11211
rect 14987 -11245 15021 -11211
rect 15055 -11245 15089 -11211
rect 15123 -11245 15157 -11211
rect 15191 -11245 15225 -11211
rect 15259 -11245 15293 -11211
rect 15327 -11245 15361 -11211
rect 15395 -11245 15429 -11211
rect 15463 -11245 15497 -11211
rect 15531 -11245 15565 -11211
rect 15599 -11245 15633 -11211
rect 15667 -11245 15701 -11211
rect 15735 -11245 15769 -11211
rect 15803 -11245 15837 -11211
rect 15871 -11245 15905 -11211
rect 15939 -11245 15973 -11211
rect 16007 -11245 16041 -11211
rect 16075 -11245 16109 -11211
rect 16143 -11245 16177 -11211
rect 16211 -11245 16245 -11211
rect 16279 -11245 16313 -11211
rect 16347 -11245 16381 -11211
rect 16415 -11245 16449 -11211
rect 16483 -11245 16517 -11211
rect 16551 -11245 16585 -11211
rect 16619 -11245 16653 -11211
rect 16687 -11245 16721 -11211
rect 16755 -11245 16789 -11211
rect 16823 -11245 16857 -11211
rect 16891 -11245 16925 -11211
rect 16959 -11245 16993 -11211
rect 17027 -11245 17061 -11211
rect 17095 -11245 17129 -11211
rect 17163 -11245 17197 -11211
rect 17231 -11245 17265 -11211
rect 17299 -11245 17333 -11211
rect 17367 -11245 17401 -11211
rect 17435 -11245 17469 -11211
rect 17503 -11245 17537 -11211
rect 17571 -11245 17605 -11211
rect 17639 -11245 17673 -11211
rect 17707 -11245 17741 -11211
rect 17775 -11245 17809 -11211
rect 17843 -11245 17877 -11211
rect 17911 -11245 17945 -11211
rect 17979 -11245 18013 -11211
rect 18047 -11245 18081 -11211
rect 18115 -11245 18149 -11211
rect 18183 -11245 18217 -11211
rect 18251 -11245 18285 -11211
rect 18319 -11245 18353 -11211
rect 18387 -11245 18421 -11211
rect 18455 -11245 18489 -11211
rect 18523 -11245 18557 -11211
rect 18591 -11245 18625 -11211
rect 18659 -11245 18693 -11211
rect 18727 -11245 18761 -11211
rect 18795 -11245 18829 -11211
rect 18863 -11245 18897 -11211
rect 18931 -11245 18965 -11211
rect 18999 -11245 19033 -11211
rect 19067 -11245 19101 -11211
rect 19135 -11245 19169 -11211
rect 19203 -11245 19237 -11211
rect 19271 -11245 19305 -11211
rect 19339 -11245 19373 -11211
rect 19407 -11245 19441 -11211
rect 19475 -11245 19509 -11211
rect 19543 -11245 19577 -11211
rect 19611 -11245 19645 -11211
rect 19679 -11245 19713 -11211
rect 19747 -11245 19781 -11211
rect 19815 -11245 19849 -11211
rect 19883 -11245 19917 -11211
rect 19951 -11245 19985 -11211
rect 20019 -11245 20053 -11211
rect 20087 -11245 20121 -11211
rect 20155 -11245 20189 -11211
rect 20223 -11245 20257 -11211
rect 20291 -11245 20325 -11211
rect 20359 -11245 20393 -11211
rect 20427 -11245 20461 -11211
rect 20495 -11245 20529 -11211
rect 20563 -11245 20597 -11211
rect 20631 -11245 20665 -11211
rect 20699 -11245 20733 -11211
rect 20767 -11245 20801 -11211
rect 20835 -11245 20869 -11211
rect 20903 -11245 20937 -11211
rect 20971 -11245 21005 -11211
rect 21039 -11245 21073 -11211
rect 21107 -11245 21141 -11211
rect 21175 -11245 21209 -11211
rect 21243 -11245 21277 -11211
rect 21311 -11245 21345 -11211
rect 21379 -11245 21413 -11211
rect 21447 -11245 21481 -11211
rect 21515 -11245 21549 -11211
rect 21583 -11245 21617 -11211
rect 21651 -11245 21685 -11211
rect 21719 -11245 21753 -11211
rect 21787 -11245 21821 -11211
rect 21855 -11245 21889 -11211
rect 21923 -11245 21957 -11211
rect 21991 -11245 22025 -11211
rect 22059 -11245 22093 -11211
rect 22127 -11245 22161 -11211
rect 22195 -11245 22229 -11211
rect 22263 -11245 22297 -11211
rect 22331 -11245 22365 -11211
rect 22399 -11245 22433 -11211
rect 22467 -11245 22501 -11211
rect 22535 -11245 22569 -11211
rect 22603 -11245 22637 -11211
rect 22671 -11245 22705 -11211
rect 22739 -11245 22773 -11211
rect 22807 -11245 22841 -11211
rect 22875 -11245 22909 -11211
rect 22943 -11245 22977 -11211
rect 23011 -11245 23045 -11211
rect 23079 -11245 23113 -11211
rect 23147 -11245 23181 -11211
rect 23215 -11245 23249 -11211
rect 23283 -11245 23317 -11211
rect 23351 -11245 23385 -11211
rect 23419 -11245 23453 -11211
rect 23487 -11245 23521 -11211
rect 23555 -11245 23589 -11211
rect 23623 -11245 23657 -11211
rect 23691 -11245 23725 -11211
rect 23759 -11245 23793 -11211
rect 23827 -11245 23861 -11211
rect 23895 -11245 23929 -11211
rect 23963 -11245 23997 -11211
rect 24031 -11245 24065 -11211
rect 24099 -11245 24133 -11211
rect 24167 -11245 24201 -11211
rect 24235 -11245 24269 -11211
rect 24303 -11245 24337 -11211
rect 24371 -11245 24405 -11211
rect 24439 -11245 24473 -11211
rect 24507 -11245 24541 -11211
rect 24575 -11245 24609 -11211
rect 24643 -11245 24677 -11211
rect 24711 -11245 24745 -11211
rect -12289 -11397 -12255 -11363
rect -12289 -11465 -12255 -11431
rect -12289 -11533 -12255 -11499
rect -12289 -11601 -12255 -11567
rect 24855 -11397 24889 -11363
rect 24855 -11465 24889 -11431
rect 24855 -11533 24889 -11499
rect 24855 -11601 24889 -11567
rect -12289 -11669 -12255 -11635
rect -12289 -11737 -12255 -11703
rect 24855 -11669 24889 -11635
rect -12289 -11805 -12255 -11771
rect -12289 -11873 -12255 -11839
rect -12289 -11941 -12255 -11907
rect -12289 -12009 -12255 -11975
rect -12289 -12077 -12255 -12043
rect -12289 -12145 -12255 -12111
rect -12289 -12213 -12255 -12179
rect -12289 -12281 -12255 -12247
rect -12289 -12349 -12255 -12315
rect 24855 -11737 24889 -11703
rect 24855 -11805 24889 -11771
rect 24855 -11873 24889 -11839
rect 24855 -11941 24889 -11907
rect 24855 -12009 24889 -11975
rect 24855 -12077 24889 -12043
rect 24855 -12145 24889 -12111
rect 24855 -12213 24889 -12179
rect 24855 -12281 24889 -12247
rect -12289 -12417 -12255 -12383
rect 24855 -12349 24889 -12315
rect 24855 -12417 24889 -12383
rect -12289 -12485 -12255 -12451
rect 24855 -12485 24889 -12451
rect -12289 -12553 -12255 -12519
rect -12289 -12621 -12255 -12587
rect -12289 -12689 -12255 -12655
rect -12289 -12757 -12255 -12723
rect -12289 -12825 -12255 -12791
rect -12289 -12893 -12255 -12859
rect -12289 -12961 -12255 -12927
rect -12289 -13029 -12255 -12995
rect -12289 -13097 -12255 -13063
rect 24855 -12553 24889 -12519
rect 24855 -12621 24889 -12587
rect 24855 -12689 24889 -12655
rect 24855 -12757 24889 -12723
rect 24855 -12825 24889 -12791
rect 24855 -12893 24889 -12859
rect -12289 -13165 -12255 -13131
rect -12289 -13233 -12255 -13199
rect -12289 -13301 -12255 -13267
rect -12289 -13369 -12255 -13335
rect -12289 -13437 -12255 -13403
rect -12289 -13505 -12255 -13471
rect -12289 -13573 -12255 -13539
rect -12289 -13641 -12255 -13607
rect -12289 -13709 -12255 -13675
rect -12289 -13777 -12255 -13743
rect -12289 -13845 -12255 -13811
rect -12289 -13913 -12255 -13879
rect 24855 -12961 24889 -12927
rect 24855 -13029 24889 -12995
rect 24855 -13097 24889 -13063
rect 24855 -13165 24889 -13131
rect 24855 -13233 24889 -13199
rect 24855 -13301 24889 -13267
rect 24855 -13369 24889 -13335
rect 24855 -13437 24889 -13403
rect 24855 -13505 24889 -13471
rect 24855 -13573 24889 -13539
rect 24855 -13641 24889 -13607
rect 24855 -13709 24889 -13675
rect 24855 -13777 24889 -13743
rect 24855 -13845 24889 -13811
rect 24855 -13913 24889 -13879
rect -12289 -13981 -12255 -13947
rect -12289 -14049 -12255 -14015
rect 24855 -13981 24889 -13947
rect 24855 -14049 24889 -14015
rect -12289 -14117 -12255 -14083
rect -12289 -14185 -12255 -14151
rect -12289 -14253 -12255 -14219
rect -12289 -14321 -12255 -14287
rect -12289 -14389 -12255 -14355
rect -12289 -14457 -12255 -14423
rect -12289 -14525 -12255 -14491
rect -12289 -14593 -12255 -14559
rect -12289 -14661 -12255 -14627
rect -12289 -14729 -12255 -14695
rect 24855 -14117 24889 -14083
rect -12289 -14797 -12255 -14763
rect -12289 -14865 -12255 -14831
rect 24855 -14185 24889 -14151
rect 24855 -14253 24889 -14219
rect 24855 -14321 24889 -14287
rect 24855 -14389 24889 -14355
rect 24855 -14457 24889 -14423
rect 24855 -14525 24889 -14491
rect 24855 -14593 24889 -14559
rect 24855 -14661 24889 -14627
rect 24855 -14729 24889 -14695
rect 24855 -14797 24889 -14763
rect 24855 -14865 24889 -14831
rect -12289 -14933 -12255 -14899
rect 24855 -14933 24889 -14899
rect -12289 -15001 -12255 -14967
rect -12289 -15069 -12255 -15035
rect -12289 -15137 -12255 -15103
rect -12289 -15205 -12255 -15171
rect -12289 -15273 -12255 -15239
rect -12289 -15341 -12255 -15307
rect -12289 -15409 -12255 -15375
rect -12289 -15477 -12255 -15443
rect -12289 -15545 -12255 -15511
rect 24855 -15001 24889 -14967
rect 24855 -15069 24889 -15035
rect 24855 -15137 24889 -15103
rect 24855 -15205 24889 -15171
rect 24855 -15273 24889 -15239
rect 24855 -15341 24889 -15307
rect 24855 -15409 24889 -15375
rect -12289 -15613 -12255 -15579
rect -12289 -15681 -12255 -15647
rect -12289 -15749 -12255 -15715
rect -12289 -15817 -12255 -15783
rect -12289 -15885 -12255 -15851
rect -12289 -15953 -12255 -15919
rect -12289 -16021 -12255 -15987
rect -12289 -16089 -12255 -16055
rect -12289 -16157 -12255 -16123
rect -12289 -16225 -12255 -16191
rect -12289 -16293 -12255 -16259
rect -12289 -16361 -12255 -16327
rect 24855 -15477 24889 -15443
rect 24855 -15545 24889 -15511
rect 24855 -15613 24889 -15579
rect 24855 -15681 24889 -15647
rect 24855 -15749 24889 -15715
rect 24855 -15817 24889 -15783
rect 24855 -15885 24889 -15851
rect 24855 -15953 24889 -15919
rect 24855 -16021 24889 -15987
rect 24855 -16089 24889 -16055
rect 24855 -16157 24889 -16123
rect 24855 -16225 24889 -16191
rect 24855 -16293 24889 -16259
rect 24855 -16361 24889 -16327
rect -12289 -16429 -12255 -16395
rect -12289 -16497 -12255 -16463
rect 24855 -16429 24889 -16395
rect 24855 -16497 24889 -16463
rect -12289 -16565 -12255 -16531
rect -12289 -16633 -12255 -16599
rect -12289 -16701 -12255 -16667
rect -12289 -16769 -12255 -16735
rect -12289 -16837 -12255 -16803
rect -12289 -16905 -12255 -16871
rect -12289 -16973 -12255 -16939
rect -12289 -17041 -12255 -17007
rect -12289 -17109 -12255 -17075
rect -12289 -17177 -12255 -17143
rect 24855 -16565 24889 -16531
rect 24855 -16633 24889 -16599
rect -12289 -17245 -12255 -17211
rect -12289 -17313 -12255 -17279
rect 24855 -16701 24889 -16667
rect 24855 -16769 24889 -16735
rect 24855 -16837 24889 -16803
rect 24855 -16905 24889 -16871
rect 24855 -16973 24889 -16939
rect 24855 -17041 24889 -17007
rect 24855 -17109 24889 -17075
rect 24855 -17177 24889 -17143
rect 24855 -17245 24889 -17211
rect -12289 -17381 -12255 -17347
rect -12289 -17449 -12255 -17415
rect 24855 -17313 24889 -17279
rect 24855 -17381 24889 -17347
rect -12289 -17517 -12255 -17483
rect -12289 -17585 -12255 -17551
rect -12289 -17653 -12255 -17619
rect -12289 -17721 -12255 -17687
rect -12289 -17789 -12255 -17755
rect -12289 -17857 -12255 -17823
rect -12289 -17925 -12255 -17891
rect -12289 -17993 -12255 -17959
rect 24855 -17449 24889 -17415
rect 24855 -17517 24889 -17483
rect 24855 -17585 24889 -17551
rect 24855 -17653 24889 -17619
rect 24855 -17721 24889 -17687
rect 24855 -17789 24889 -17755
rect 24855 -17857 24889 -17823
rect -12289 -18061 -12255 -18027
rect -12289 -18129 -12255 -18095
rect -12289 -18197 -12255 -18163
rect -12289 -18265 -12255 -18231
rect -12289 -18333 -12255 -18299
rect -12289 -18401 -12255 -18367
rect -12289 -18469 -12255 -18435
rect -12289 -18537 -12255 -18503
rect -12289 -18605 -12255 -18571
rect -12289 -18673 -12255 -18639
rect -12289 -18741 -12255 -18707
rect -12289 -18809 -12255 -18775
rect 24855 -17925 24889 -17891
rect 24855 -17993 24889 -17959
rect 24855 -18061 24889 -18027
rect 24855 -18129 24889 -18095
rect 24855 -18197 24889 -18163
rect 24855 -18265 24889 -18231
rect 24855 -18333 24889 -18299
rect 24855 -18401 24889 -18367
rect 24855 -18469 24889 -18435
rect 24855 -18537 24889 -18503
rect 24855 -18605 24889 -18571
rect 24855 -18673 24889 -18639
rect 24855 -18741 24889 -18707
rect 24855 -18809 24889 -18775
rect -12289 -18877 -12255 -18843
rect -12289 -18945 -12255 -18911
rect 24855 -18877 24889 -18843
rect -12289 -19013 -12255 -18979
rect 24855 -18945 24889 -18911
rect 24855 -19013 24889 -18979
rect -12289 -19081 -12255 -19047
rect -12289 -19149 -12255 -19115
rect 24855 -19081 24889 -19047
rect -12289 -19217 -12255 -19183
rect -12289 -19285 -12255 -19251
rect -12289 -19353 -12255 -19319
rect -12289 -19421 -12255 -19387
rect -12289 -19489 -12255 -19455
rect -12289 -19557 -12255 -19523
rect -12289 -19625 -12255 -19591
rect -12289 -19693 -12255 -19659
rect -12289 -19761 -12255 -19727
rect -12289 -19829 -12255 -19795
rect 24855 -19149 24889 -19115
rect 24855 -19217 24889 -19183
rect 24855 -19285 24889 -19251
rect 24855 -19353 24889 -19319
rect 24855 -19421 24889 -19387
rect 24855 -19489 24889 -19455
rect 24855 -19557 24889 -19523
rect 24855 -19625 24889 -19591
rect 24855 -19693 24889 -19659
rect 24855 -19761 24889 -19727
rect -12289 -19897 -12255 -19863
rect 24855 -19829 24889 -19795
rect 24855 -19897 24889 -19863
rect -12289 -19965 -12255 -19931
rect -12289 -20033 -12255 -19999
rect -12289 -20101 -12255 -20067
rect -12289 -20169 -12255 -20135
rect -12289 -20237 -12255 -20203
rect 24855 -19965 24889 -19931
rect 24855 -20033 24889 -19999
rect 24855 -20101 24889 -20067
rect 24855 -20169 24889 -20135
rect 24855 -20237 24889 -20203
rect -12289 -20305 -12255 -20271
rect -12289 -20373 -12255 -20339
rect 24855 -20305 24889 -20271
rect -12289 -20441 -12255 -20407
rect -12289 -20509 -12255 -20475
rect -12289 -20577 -12255 -20543
rect -12289 -20645 -12255 -20611
rect -12289 -20713 -12255 -20679
rect -12289 -20781 -12255 -20747
rect -12289 -20849 -12255 -20815
rect -12289 -20917 -12255 -20883
rect -12289 -20985 -12255 -20951
rect 24855 -20373 24889 -20339
rect 24855 -20441 24889 -20407
rect 24855 -20509 24889 -20475
rect 24855 -20577 24889 -20543
rect 24855 -20645 24889 -20611
rect 24855 -20713 24889 -20679
rect 24855 -20781 24889 -20747
rect 24855 -20849 24889 -20815
rect 24855 -20917 24889 -20883
rect -12289 -21053 -12255 -21019
rect 24855 -20985 24889 -20951
rect -12289 -21121 -12255 -21087
rect -12289 -21189 -12255 -21155
rect -12289 -21257 -12255 -21223
rect -12289 -21325 -12255 -21291
rect -12289 -21393 -12255 -21359
rect -12289 -21461 -12255 -21427
rect -12289 -21529 -12255 -21495
rect 24855 -21053 24889 -21019
rect 24855 -21121 24889 -21087
rect 24855 -21189 24889 -21155
rect 24855 -21257 24889 -21223
rect 24855 -21325 24889 -21291
rect 24855 -21393 24889 -21359
rect 24855 -21461 24889 -21427
rect -12289 -21597 -12255 -21563
rect 24855 -21529 24889 -21495
rect -12289 -21665 -12255 -21631
rect -12289 -21733 -12255 -21699
rect -12289 -21801 -12255 -21767
rect -12289 -21869 -12255 -21835
rect -12289 -21937 -12255 -21903
rect -12289 -22005 -12255 -21971
rect -12289 -22073 -12255 -22039
rect -12289 -22141 -12255 -22107
rect -12289 -22209 -12255 -22175
rect -12289 -22277 -12255 -22243
rect -12289 -22345 -12255 -22311
rect -12289 -22413 -12255 -22379
rect 24855 -21597 24889 -21563
rect 24855 -21665 24889 -21631
rect 24855 -21733 24889 -21699
rect 24855 -21801 24889 -21767
rect 24855 -21869 24889 -21835
rect 24855 -21937 24889 -21903
rect 24855 -22005 24889 -21971
rect 24855 -22073 24889 -22039
rect 24855 -22141 24889 -22107
rect 24855 -22209 24889 -22175
rect 24855 -22277 24889 -22243
rect 24855 -22345 24889 -22311
rect -12289 -22481 -12255 -22447
rect 24855 -22413 24889 -22379
rect -12289 -22549 -12255 -22515
rect -12289 -22617 -12255 -22583
rect -12289 -22685 -12255 -22651
rect -12289 -22753 -12255 -22719
rect 24855 -22481 24889 -22447
rect 24855 -22549 24889 -22515
rect 24855 -22617 24889 -22583
rect 24855 -22685 24889 -22651
rect -12289 -22821 -12255 -22787
rect -12289 -22889 -12255 -22855
rect 24855 -22753 24889 -22719
rect -12289 -22957 -12255 -22923
rect -12289 -23025 -12255 -22991
rect -12289 -23093 -12255 -23059
rect -12289 -23161 -12255 -23127
rect -12289 -23229 -12255 -23195
rect -12289 -23297 -12255 -23263
rect -12289 -23365 -12255 -23331
rect -12289 -23433 -12255 -23399
rect -12289 -23501 -12255 -23467
rect 24855 -22821 24889 -22787
rect 24855 -22889 24889 -22855
rect 24855 -22957 24889 -22923
rect 24855 -23025 24889 -22991
rect 24855 -23093 24889 -23059
rect 24855 -23161 24889 -23127
rect 24855 -23229 24889 -23195
rect 24855 -23297 24889 -23263
rect 24855 -23365 24889 -23331
rect -12289 -23569 -12255 -23535
rect 24855 -23433 24889 -23399
rect 24855 -23501 24889 -23467
rect 24855 -23569 24889 -23535
rect -12289 -23637 -12255 -23603
rect -12289 -23705 -12255 -23671
rect -12289 -23773 -12255 -23739
rect -12289 -23841 -12255 -23807
rect -12289 -23909 -12255 -23875
rect 24855 -23637 24889 -23603
rect 24855 -23705 24889 -23671
rect 24855 -23773 24889 -23739
rect 24855 -23841 24889 -23807
rect 24855 -23909 24889 -23875
rect -12289 -23977 -12255 -23943
rect -12289 -24045 -12255 -24011
rect -12289 -24113 -12255 -24079
rect -12289 -24181 -12255 -24147
rect -12289 -24249 -12255 -24215
rect -12289 -24317 -12255 -24283
rect -12289 -24385 -12255 -24351
rect -12289 -24453 -12255 -24419
rect -12289 -24521 -12255 -24487
rect -12289 -24589 -12255 -24555
rect 24855 -23977 24889 -23943
rect 24855 -24045 24889 -24011
rect -12289 -24657 -12255 -24623
rect -12289 -24725 -12255 -24691
rect 24855 -24113 24889 -24079
rect 24855 -24181 24889 -24147
rect 24855 -24249 24889 -24215
rect 24855 -24317 24889 -24283
rect 24855 -24385 24889 -24351
rect 24855 -24453 24889 -24419
rect 24855 -24521 24889 -24487
rect 24855 -24589 24889 -24555
rect 24855 -24657 24889 -24623
rect 24855 -24725 24889 -24691
rect -12289 -24793 -12255 -24759
rect -12289 -24861 -12255 -24827
rect -12289 -24929 -12255 -24895
rect -12289 -24997 -12255 -24963
rect 24855 -24793 24889 -24759
rect 24855 -24861 24889 -24827
rect 24855 -24929 24889 -24895
rect 24855 -24997 24889 -24963
rect -12289 -25065 -12255 -25031
rect -12289 -25133 -12255 -25099
rect 24855 -25065 24889 -25031
rect -12289 -25201 -12255 -25167
rect -12289 -25269 -12255 -25235
rect -12289 -25337 -12255 -25303
rect -12289 -25405 -12255 -25371
rect -12289 -25473 -12255 -25439
rect -12289 -25541 -12255 -25507
rect -12289 -25609 -12255 -25575
rect -12289 -25677 -12255 -25643
rect -12289 -25745 -12255 -25711
rect 24855 -25133 24889 -25099
rect 24855 -25201 24889 -25167
rect 24855 -25269 24889 -25235
rect -12289 -25813 -12255 -25779
rect -12289 -25881 -12255 -25847
rect 24855 -25337 24889 -25303
rect 24855 -25405 24889 -25371
rect 24855 -25473 24889 -25439
rect 24855 -25541 24889 -25507
rect 24855 -25609 24889 -25575
rect 24855 -25677 24889 -25643
rect 24855 -25745 24889 -25711
rect 24855 -25813 24889 -25779
rect 24855 -25881 24889 -25847
rect -12289 -25949 -12255 -25915
rect 24855 -25949 24889 -25915
rect -12289 -26017 -12255 -25983
rect -12289 -26085 -12255 -26051
rect -12289 -26153 -12255 -26119
rect -12289 -26221 -12255 -26187
rect -12289 -26289 -12255 -26255
rect -12289 -26357 -12255 -26323
rect -12289 -26425 -12255 -26391
rect -12289 -26493 -12255 -26459
rect -12289 -26561 -12255 -26527
rect -12289 -26629 -12255 -26595
rect -12289 -26697 -12255 -26663
rect -12289 -26765 -12255 -26731
rect -12289 -26833 -12255 -26799
rect -12289 -26901 -12255 -26867
rect -12289 -26969 -12255 -26935
rect -12289 -27037 -12255 -27003
rect 24855 -26017 24889 -25983
rect 24855 -26085 24889 -26051
rect 24855 -26153 24889 -26119
rect 24855 -26221 24889 -26187
rect 24855 -26289 24889 -26255
rect 24855 -26357 24889 -26323
rect 24855 -26425 24889 -26391
rect 24855 -26493 24889 -26459
rect 24855 -26561 24889 -26527
rect 24855 -26629 24889 -26595
rect 24855 -26697 24889 -26663
rect 24855 -26765 24889 -26731
rect 24855 -26833 24889 -26799
rect 24855 -26901 24889 -26867
rect 24855 -26969 24889 -26935
rect 24855 -27037 24889 -27003
rect -12145 -27189 -12111 -27155
rect -12077 -27189 -12043 -27155
rect -12009 -27189 -11975 -27155
rect -11941 -27189 -11907 -27155
rect -11873 -27189 -11839 -27155
rect -11805 -27189 -11771 -27155
rect -11737 -27189 -11703 -27155
rect -11669 -27189 -11635 -27155
rect -11601 -27189 -11567 -27155
rect -11533 -27189 -11499 -27155
rect -11465 -27189 -11431 -27155
rect -11397 -27189 -11363 -27155
rect -11329 -27189 -11295 -27155
rect -11261 -27189 -11227 -27155
rect -11193 -27189 -11159 -27155
rect -11125 -27189 -11091 -27155
rect -11057 -27189 -11023 -27155
rect -10989 -27189 -10955 -27155
rect -10921 -27189 -10887 -27155
rect -10853 -27189 -10819 -27155
rect -10785 -27189 -10751 -27155
rect -10717 -27189 -10683 -27155
rect -10649 -27189 -10615 -27155
rect -10581 -27189 -10547 -27155
rect -10513 -27189 -10479 -27155
rect -10445 -27189 -10411 -27155
rect -10377 -27189 -10343 -27155
rect -10309 -27189 -10275 -27155
rect -10241 -27189 -10207 -27155
rect -10173 -27189 -10139 -27155
rect -10105 -27189 -10071 -27155
rect -10037 -27189 -10003 -27155
rect -9969 -27189 -9935 -27155
rect -9901 -27189 -9867 -27155
rect -9833 -27189 -9799 -27155
rect -9765 -27189 -9731 -27155
rect -9697 -27189 -9663 -27155
rect -9629 -27189 -9595 -27155
rect -9561 -27189 -9527 -27155
rect -9493 -27189 -9459 -27155
rect -9425 -27189 -9391 -27155
rect -9357 -27189 -9323 -27155
rect -9289 -27189 -9255 -27155
rect -9221 -27189 -9187 -27155
rect -9153 -27189 -9119 -27155
rect -9085 -27189 -9051 -27155
rect -9017 -27189 -8983 -27155
rect -8949 -27189 -8915 -27155
rect -8881 -27189 -8847 -27155
rect -8813 -27189 -8779 -27155
rect -8745 -27189 -8711 -27155
rect -8677 -27189 -8643 -27155
rect -8609 -27189 -8575 -27155
rect -8541 -27189 -8507 -27155
rect -8473 -27189 -8439 -27155
rect -8405 -27189 -8371 -27155
rect -8337 -27189 -8303 -27155
rect -8269 -27189 -8235 -27155
rect -8201 -27189 -8167 -27155
rect -8133 -27189 -8099 -27155
rect -8065 -27189 -8031 -27155
rect -7997 -27189 -7963 -27155
rect -7929 -27189 -7895 -27155
rect -7861 -27189 -7827 -27155
rect -7793 -27189 -7759 -27155
rect -7725 -27189 -7691 -27155
rect -7657 -27189 -7623 -27155
rect -7589 -27189 -7555 -27155
rect -7521 -27189 -7487 -27155
rect -7453 -27189 -7419 -27155
rect -7385 -27189 -7351 -27155
rect -7317 -27189 -7283 -27155
rect -7249 -27189 -7215 -27155
rect -7181 -27189 -7147 -27155
rect -7113 -27189 -7079 -27155
rect -7045 -27189 -7011 -27155
rect -6977 -27189 -6943 -27155
rect -6909 -27189 -6875 -27155
rect -6841 -27189 -6807 -27155
rect -6773 -27189 -6739 -27155
rect -6705 -27189 -6671 -27155
rect -6637 -27189 -6603 -27155
rect -6569 -27189 -6535 -27155
rect -6501 -27189 -6467 -27155
rect -6433 -27189 -6399 -27155
rect -6365 -27189 -6331 -27155
rect -6297 -27189 -6263 -27155
rect -6229 -27189 -6195 -27155
rect -6161 -27189 -6127 -27155
rect -6093 -27189 -6059 -27155
rect -6025 -27189 -5991 -27155
rect -5957 -27189 -5923 -27155
rect -5889 -27189 -5855 -27155
rect -5821 -27189 -5787 -27155
rect -5753 -27189 -5719 -27155
rect -5685 -27189 -5651 -27155
rect -5617 -27189 -5583 -27155
rect -5549 -27189 -5515 -27155
rect -5481 -27189 -5447 -27155
rect -5413 -27189 -5379 -27155
rect -5345 -27189 -5311 -27155
rect -5277 -27189 -5243 -27155
rect -5209 -27189 -5175 -27155
rect -5141 -27189 -5107 -27155
rect -5073 -27189 -5039 -27155
rect -5005 -27189 -4971 -27155
rect -4937 -27189 -4903 -27155
rect -4869 -27189 -4835 -27155
rect -4801 -27189 -4767 -27155
rect -4733 -27189 -4699 -27155
rect -4665 -27189 -4631 -27155
rect -4597 -27189 -4563 -27155
rect -4529 -27189 -4495 -27155
rect -4461 -27189 -4427 -27155
rect -4393 -27189 -4359 -27155
rect -4325 -27189 -4291 -27155
rect -4257 -27189 -4223 -27155
rect -4189 -27189 -4155 -27155
rect -4121 -27189 -4087 -27155
rect -4053 -27189 -4019 -27155
rect -3985 -27189 -3951 -27155
rect -3917 -27189 -3883 -27155
rect -3849 -27189 -3815 -27155
rect -3781 -27189 -3747 -27155
rect -3713 -27189 -3679 -27155
rect -3645 -27189 -3611 -27155
rect -3577 -27189 -3543 -27155
rect -3509 -27189 -3475 -27155
rect -3441 -27189 -3407 -27155
rect -3373 -27189 -3339 -27155
rect -3305 -27189 -3271 -27155
rect -3237 -27189 -3203 -27155
rect -3169 -27189 -3135 -27155
rect -3101 -27189 -3067 -27155
rect -3033 -27189 -2999 -27155
rect -2965 -27189 -2931 -27155
rect -2897 -27189 -2863 -27155
rect -2829 -27189 -2795 -27155
rect -2761 -27189 -2727 -27155
rect -2693 -27189 -2659 -27155
rect -2625 -27189 -2591 -27155
rect -2557 -27189 -2523 -27155
rect -2489 -27189 -2455 -27155
rect -2421 -27189 -2387 -27155
rect -2353 -27189 -2319 -27155
rect -2285 -27189 -2251 -27155
rect -2217 -27189 -2183 -27155
rect -2149 -27189 -2115 -27155
rect -2081 -27189 -2047 -27155
rect -2013 -27189 -1979 -27155
rect -1945 -27189 -1911 -27155
rect -1877 -27189 -1843 -27155
rect -1809 -27189 -1775 -27155
rect -1741 -27189 -1707 -27155
rect -1673 -27189 -1639 -27155
rect -1605 -27189 -1571 -27155
rect -1537 -27189 -1503 -27155
rect -1469 -27189 -1435 -27155
rect -1401 -27189 -1367 -27155
rect -1333 -27189 -1299 -27155
rect -1265 -27189 -1231 -27155
rect -1197 -27189 -1163 -27155
rect -1129 -27189 -1095 -27155
rect -1061 -27189 -1027 -27155
rect -993 -27189 -959 -27155
rect -925 -27189 -891 -27155
rect -857 -27189 -823 -27155
rect -789 -27189 -755 -27155
rect -721 -27189 -687 -27155
rect -653 -27189 -619 -27155
rect -585 -27189 -551 -27155
rect -517 -27189 -483 -27155
rect -449 -27189 -415 -27155
rect -381 -27189 -347 -27155
rect -313 -27189 -279 -27155
rect -245 -27189 -211 -27155
rect -177 -27189 -143 -27155
rect -109 -27189 -75 -27155
rect -41 -27189 -7 -27155
rect 27 -27189 61 -27155
rect 95 -27189 129 -27155
rect 163 -27189 197 -27155
rect 231 -27189 265 -27155
rect 299 -27189 333 -27155
rect 367 -27189 401 -27155
rect 435 -27189 469 -27155
rect 503 -27189 537 -27155
rect 571 -27189 605 -27155
rect 639 -27189 673 -27155
rect 707 -27189 741 -27155
rect 775 -27189 809 -27155
rect 843 -27189 877 -27155
rect 911 -27189 945 -27155
rect 979 -27189 1013 -27155
rect 1047 -27189 1081 -27155
rect 1115 -27189 1149 -27155
rect 1183 -27189 1217 -27155
rect 1251 -27189 1285 -27155
rect 1319 -27189 1353 -27155
rect 1387 -27189 1421 -27155
rect 1455 -27189 1489 -27155
rect 1523 -27189 1557 -27155
rect 1591 -27189 1625 -27155
rect 1659 -27189 1693 -27155
rect 1727 -27189 1761 -27155
rect 1795 -27189 1829 -27155
rect 1863 -27189 1897 -27155
rect 1931 -27189 1965 -27155
rect 1999 -27189 2033 -27155
rect 2067 -27189 2101 -27155
rect 2135 -27189 2169 -27155
rect 2203 -27189 2237 -27155
rect 2271 -27189 2305 -27155
rect 2339 -27189 2373 -27155
rect 2407 -27189 2441 -27155
rect 2475 -27189 2509 -27155
rect 2543 -27189 2577 -27155
rect 2611 -27189 2645 -27155
rect 2679 -27189 2713 -27155
rect 2747 -27189 2781 -27155
rect 2815 -27189 2849 -27155
rect 2883 -27189 2917 -27155
rect 2951 -27189 2985 -27155
rect 3019 -27189 3053 -27155
rect 3087 -27189 3121 -27155
rect 3155 -27189 3189 -27155
rect 3223 -27189 3257 -27155
rect 3291 -27189 3325 -27155
rect 3359 -27189 3393 -27155
rect 3427 -27189 3461 -27155
rect 3495 -27189 3529 -27155
rect 3563 -27189 3597 -27155
rect 3631 -27189 3665 -27155
rect 3699 -27189 3733 -27155
rect 3767 -27189 3801 -27155
rect 3835 -27189 3869 -27155
rect 3903 -27189 3937 -27155
rect 3971 -27189 4005 -27155
rect 4039 -27189 4073 -27155
rect 4107 -27189 4141 -27155
rect 4175 -27189 4209 -27155
rect 4243 -27189 4277 -27155
rect 4311 -27189 4345 -27155
rect 4379 -27189 4413 -27155
rect 4447 -27189 4481 -27155
rect 4515 -27189 4549 -27155
rect 4583 -27189 4617 -27155
rect 4651 -27189 4685 -27155
rect 4719 -27189 4753 -27155
rect 4787 -27189 4821 -27155
rect 4855 -27189 4889 -27155
rect 4923 -27189 4957 -27155
rect 4991 -27189 5025 -27155
rect 5059 -27189 5093 -27155
rect 5127 -27189 5161 -27155
rect 5195 -27189 5229 -27155
rect 5263 -27189 5297 -27155
rect 5331 -27189 5365 -27155
rect 5399 -27189 5433 -27155
rect 5467 -27189 5501 -27155
rect 5535 -27189 5569 -27155
rect 5603 -27189 5637 -27155
rect 5671 -27189 5705 -27155
rect 5739 -27189 5773 -27155
rect 5807 -27189 5841 -27155
rect 5875 -27189 5909 -27155
rect 5943 -27189 5977 -27155
rect 6011 -27189 6045 -27155
rect 6079 -27189 6113 -27155
rect 6147 -27189 6181 -27155
rect 6215 -27189 6249 -27155
rect 6283 -27189 6317 -27155
rect 6351 -27189 6385 -27155
rect 6419 -27189 6453 -27155
rect 6487 -27189 6521 -27155
rect 6555 -27189 6589 -27155
rect 6623 -27189 6657 -27155
rect 6691 -27189 6725 -27155
rect 6759 -27189 6793 -27155
rect 6827 -27189 6861 -27155
rect 6895 -27189 6929 -27155
rect 6963 -27189 6997 -27155
rect 7031 -27189 7065 -27155
rect 7099 -27189 7133 -27155
rect 7167 -27189 7201 -27155
rect 7235 -27189 7269 -27155
rect 7303 -27189 7337 -27155
rect 7371 -27189 7405 -27155
rect 7439 -27189 7473 -27155
rect 7507 -27189 7541 -27155
rect 7575 -27189 7609 -27155
rect 7643 -27189 7677 -27155
rect 7711 -27189 7745 -27155
rect 7779 -27189 7813 -27155
rect 7847 -27189 7881 -27155
rect 7915 -27189 7949 -27155
rect 7983 -27189 8017 -27155
rect 8051 -27189 8085 -27155
rect 8119 -27189 8153 -27155
rect 8187 -27189 8221 -27155
rect 8255 -27189 8289 -27155
rect 8323 -27189 8357 -27155
rect 8391 -27189 8425 -27155
rect 8459 -27189 8493 -27155
rect 8527 -27189 8561 -27155
rect 8595 -27189 8629 -27155
rect 8663 -27189 8697 -27155
rect 8731 -27189 8765 -27155
rect 8799 -27189 8833 -27155
rect 8867 -27189 8901 -27155
rect 8935 -27189 8969 -27155
rect 9003 -27189 9037 -27155
rect 9071 -27189 9105 -27155
rect 9139 -27189 9173 -27155
rect 9207 -27189 9241 -27155
rect 9275 -27189 9309 -27155
rect 9343 -27189 9377 -27155
rect 9411 -27189 9445 -27155
rect 9479 -27189 9513 -27155
rect 9547 -27189 9581 -27155
rect 9615 -27189 9649 -27155
rect 9683 -27189 9717 -27155
rect 9751 -27189 9785 -27155
rect 9819 -27189 9853 -27155
rect 9887 -27189 9921 -27155
rect 9955 -27189 9989 -27155
rect 10023 -27189 10057 -27155
rect 10091 -27189 10125 -27155
rect 10159 -27189 10193 -27155
rect 10227 -27189 10261 -27155
rect 10295 -27189 10329 -27155
rect 10363 -27189 10397 -27155
rect 10431 -27189 10465 -27155
rect 10499 -27189 10533 -27155
rect 10567 -27189 10601 -27155
rect 10635 -27189 10669 -27155
rect 10703 -27189 10737 -27155
rect 10771 -27189 10805 -27155
rect 10839 -27189 10873 -27155
rect 10907 -27189 10941 -27155
rect 10975 -27189 11009 -27155
rect 11043 -27189 11077 -27155
rect 11111 -27189 11145 -27155
rect 11179 -27189 11213 -27155
rect 11247 -27189 11281 -27155
rect 11315 -27189 11349 -27155
rect 11383 -27189 11417 -27155
rect 11451 -27189 11485 -27155
rect 11519 -27189 11553 -27155
rect 11587 -27189 11621 -27155
rect 11655 -27189 11689 -27155
rect 11723 -27189 11757 -27155
rect 11791 -27189 11825 -27155
rect 11859 -27189 11893 -27155
rect 11927 -27189 11961 -27155
rect 11995 -27189 12029 -27155
rect 12063 -27189 12097 -27155
rect 12131 -27189 12165 -27155
rect 12199 -27189 12233 -27155
rect 12267 -27189 12301 -27155
rect 12335 -27189 12369 -27155
rect 12403 -27189 12437 -27155
rect 12471 -27189 12505 -27155
rect 12539 -27189 12573 -27155
rect 12607 -27189 12641 -27155
rect 12675 -27189 12709 -27155
rect 12743 -27189 12777 -27155
rect 12811 -27189 12845 -27155
rect 12879 -27189 12913 -27155
rect 12947 -27189 12981 -27155
rect 13015 -27189 13049 -27155
rect 13083 -27189 13117 -27155
rect 13151 -27189 13185 -27155
rect 13219 -27189 13253 -27155
rect 13287 -27189 13321 -27155
rect 13355 -27189 13389 -27155
rect 13423 -27189 13457 -27155
rect 13491 -27189 13525 -27155
rect 13559 -27189 13593 -27155
rect 13627 -27189 13661 -27155
rect 13695 -27189 13729 -27155
rect 13763 -27189 13797 -27155
rect 13831 -27189 13865 -27155
rect 13899 -27189 13933 -27155
rect 13967 -27189 14001 -27155
rect 14035 -27189 14069 -27155
rect 14103 -27189 14137 -27155
rect 14171 -27189 14205 -27155
rect 14239 -27189 14273 -27155
rect 14307 -27189 14341 -27155
rect 14375 -27189 14409 -27155
rect 14443 -27189 14477 -27155
rect 14511 -27189 14545 -27155
rect 14579 -27189 14613 -27155
rect 14647 -27189 14681 -27155
rect 14715 -27189 14749 -27155
rect 14783 -27189 14817 -27155
rect 14851 -27189 14885 -27155
rect 14919 -27189 14953 -27155
rect 14987 -27189 15021 -27155
rect 15055 -27189 15089 -27155
rect 15123 -27189 15157 -27155
rect 15191 -27189 15225 -27155
rect 15259 -27189 15293 -27155
rect 15327 -27189 15361 -27155
rect 15395 -27189 15429 -27155
rect 15463 -27189 15497 -27155
rect 15531 -27189 15565 -27155
rect 15599 -27189 15633 -27155
rect 15667 -27189 15701 -27155
rect 15735 -27189 15769 -27155
rect 15803 -27189 15837 -27155
rect 15871 -27189 15905 -27155
rect 15939 -27189 15973 -27155
rect 16007 -27189 16041 -27155
rect 16075 -27189 16109 -27155
rect 16143 -27189 16177 -27155
rect 16211 -27189 16245 -27155
rect 16279 -27189 16313 -27155
rect 16347 -27189 16381 -27155
rect 16415 -27189 16449 -27155
rect 16483 -27189 16517 -27155
rect 16551 -27189 16585 -27155
rect 16619 -27189 16653 -27155
rect 16687 -27189 16721 -27155
rect 16755 -27189 16789 -27155
rect 16823 -27189 16857 -27155
rect 16891 -27189 16925 -27155
rect 16959 -27189 16993 -27155
rect 17027 -27189 17061 -27155
rect 17095 -27189 17129 -27155
rect 17163 -27189 17197 -27155
rect 17231 -27189 17265 -27155
rect 17299 -27189 17333 -27155
rect 17367 -27189 17401 -27155
rect 17435 -27189 17469 -27155
rect 17503 -27189 17537 -27155
rect 17571 -27189 17605 -27155
rect 17639 -27189 17673 -27155
rect 17707 -27189 17741 -27155
rect 17775 -27189 17809 -27155
rect 17843 -27189 17877 -27155
rect 17911 -27189 17945 -27155
rect 17979 -27189 18013 -27155
rect 18047 -27189 18081 -27155
rect 18115 -27189 18149 -27155
rect 18183 -27189 18217 -27155
rect 18251 -27189 18285 -27155
rect 18319 -27189 18353 -27155
rect 18387 -27189 18421 -27155
rect 18455 -27189 18489 -27155
rect 18523 -27189 18557 -27155
rect 18591 -27189 18625 -27155
rect 18659 -27189 18693 -27155
rect 18727 -27189 18761 -27155
rect 18795 -27189 18829 -27155
rect 18863 -27189 18897 -27155
rect 18931 -27189 18965 -27155
rect 18999 -27189 19033 -27155
rect 19067 -27189 19101 -27155
rect 19135 -27189 19169 -27155
rect 19203 -27189 19237 -27155
rect 19271 -27189 19305 -27155
rect 19339 -27189 19373 -27155
rect 19407 -27189 19441 -27155
rect 19475 -27189 19509 -27155
rect 19543 -27189 19577 -27155
rect 19611 -27189 19645 -27155
rect 19679 -27189 19713 -27155
rect 19747 -27189 19781 -27155
rect 19815 -27189 19849 -27155
rect 19883 -27189 19917 -27155
rect 19951 -27189 19985 -27155
rect 20019 -27189 20053 -27155
rect 20087 -27189 20121 -27155
rect 20155 -27189 20189 -27155
rect 20223 -27189 20257 -27155
rect 20291 -27189 20325 -27155
rect 20359 -27189 20393 -27155
rect 20427 -27189 20461 -27155
rect 20495 -27189 20529 -27155
rect 20563 -27189 20597 -27155
rect 20631 -27189 20665 -27155
rect 20699 -27189 20733 -27155
rect 20767 -27189 20801 -27155
rect 20835 -27189 20869 -27155
rect 20903 -27189 20937 -27155
rect 20971 -27189 21005 -27155
rect 21039 -27189 21073 -27155
rect 21107 -27189 21141 -27155
rect 21175 -27189 21209 -27155
rect 21243 -27189 21277 -27155
rect 21311 -27189 21345 -27155
rect 21379 -27189 21413 -27155
rect 21447 -27189 21481 -27155
rect 21515 -27189 21549 -27155
rect 21583 -27189 21617 -27155
rect 21651 -27189 21685 -27155
rect 21719 -27189 21753 -27155
rect 21787 -27189 21821 -27155
rect 21855 -27189 21889 -27155
rect 21923 -27189 21957 -27155
rect 21991 -27189 22025 -27155
rect 22059 -27189 22093 -27155
rect 22127 -27189 22161 -27155
rect 22195 -27189 22229 -27155
rect 22263 -27189 22297 -27155
rect 22331 -27189 22365 -27155
rect 22399 -27189 22433 -27155
rect 22467 -27189 22501 -27155
rect 22535 -27189 22569 -27155
rect 22603 -27189 22637 -27155
rect 22671 -27189 22705 -27155
rect 22739 -27189 22773 -27155
rect 22807 -27189 22841 -27155
rect 22875 -27189 22909 -27155
rect 22943 -27189 22977 -27155
rect 23011 -27189 23045 -27155
rect 23079 -27189 23113 -27155
rect 23147 -27189 23181 -27155
rect 23215 -27189 23249 -27155
rect 23283 -27189 23317 -27155
rect 23351 -27189 23385 -27155
rect 23419 -27189 23453 -27155
rect 23487 -27189 23521 -27155
rect 23555 -27189 23589 -27155
rect 23623 -27189 23657 -27155
rect 23691 -27189 23725 -27155
rect 23759 -27189 23793 -27155
rect 23827 -27189 23861 -27155
rect 23895 -27189 23929 -27155
rect 23963 -27189 23997 -27155
rect 24031 -27189 24065 -27155
rect 24099 -27189 24133 -27155
rect 24167 -27189 24201 -27155
rect 24235 -27189 24269 -27155
rect 24303 -27189 24337 -27155
rect 24371 -27189 24405 -27155
rect 24439 -27189 24473 -27155
rect 24507 -27189 24541 -27155
rect 24575 -27189 24609 -27155
rect 24643 -27189 24677 -27155
rect 24711 -27189 24745 -27155
<< nsubdiffcont >>
rect 547 1655 581 1689
rect 615 1655 649 1689
rect 683 1655 717 1689
rect 751 1655 785 1689
rect 819 1655 853 1689
rect 887 1655 921 1689
rect 955 1655 989 1689
rect 1023 1655 1057 1689
rect 1091 1655 1125 1689
rect 1159 1655 1193 1689
rect 1227 1655 1261 1689
rect 1295 1655 1329 1689
rect 1363 1655 1397 1689
rect 1431 1655 1465 1689
rect 1499 1655 1533 1689
rect 1567 1655 1601 1689
rect 1635 1655 1669 1689
rect 1703 1655 1737 1689
rect 1771 1655 1805 1689
rect 1839 1655 1873 1689
rect 1907 1655 1941 1689
rect 1975 1655 2009 1689
rect 2043 1655 2077 1689
rect 2111 1655 2145 1689
rect 2179 1655 2213 1689
rect 2247 1655 2281 1689
rect 2315 1655 2349 1689
rect 2383 1655 2417 1689
rect 2451 1655 2485 1689
rect 2519 1655 2553 1689
rect 2587 1655 2621 1689
rect 2655 1655 2689 1689
rect 2723 1655 2757 1689
rect 2791 1655 2825 1689
rect 2859 1655 2893 1689
rect 2927 1655 2961 1689
rect 2995 1655 3029 1689
rect 3063 1655 3097 1689
rect 3131 1655 3165 1689
rect 3199 1655 3233 1689
rect 3267 1655 3301 1689
rect 3335 1655 3369 1689
rect 3403 1655 3437 1689
rect 3471 1655 3505 1689
rect 3539 1655 3573 1689
rect 3607 1655 3641 1689
rect 3675 1655 3709 1689
rect 3743 1655 3777 1689
rect 3811 1655 3845 1689
rect 3879 1655 3913 1689
rect 3947 1655 3981 1689
rect 4015 1655 4049 1689
rect 4083 1655 4117 1689
rect 4151 1655 4185 1689
rect 4219 1655 4253 1689
rect 4287 1655 4321 1689
rect 4355 1655 4389 1689
rect 4423 1655 4457 1689
rect 4491 1655 4525 1689
rect 4559 1655 4593 1689
rect 4627 1655 4661 1689
rect 4695 1655 4729 1689
rect 4763 1655 4797 1689
rect 4831 1655 4865 1689
rect 4899 1655 4933 1689
rect 4967 1655 5001 1689
rect 5035 1655 5069 1689
rect 5103 1655 5137 1689
rect 5171 1655 5205 1689
rect 5239 1655 5273 1689
rect 5307 1655 5341 1689
rect 5375 1655 5409 1689
rect 5443 1655 5477 1689
rect 5511 1655 5545 1689
rect 5579 1655 5613 1689
rect 5647 1655 5681 1689
rect 5715 1655 5749 1689
rect 5783 1655 5817 1689
rect 5851 1655 5885 1689
rect 5919 1655 5953 1689
rect 5987 1655 6021 1689
rect 6055 1655 6089 1689
rect 6123 1655 6157 1689
rect 6191 1655 6225 1689
rect 6259 1655 6293 1689
rect 6327 1655 6361 1689
rect 6395 1655 6429 1689
rect 6463 1655 6497 1689
rect 6531 1655 6565 1689
rect 6599 1655 6633 1689
rect 6667 1655 6701 1689
rect 6735 1655 6769 1689
rect 6803 1655 6837 1689
rect 6871 1655 6905 1689
rect 6939 1655 6973 1689
rect 7007 1655 7041 1689
rect 7075 1655 7109 1689
rect 7143 1655 7177 1689
rect 7211 1655 7245 1689
rect 7279 1655 7313 1689
rect 7347 1655 7381 1689
rect 7415 1655 7449 1689
rect 7483 1655 7517 1689
rect 7551 1655 7585 1689
rect 7619 1655 7653 1689
rect 7687 1655 7721 1689
rect 7755 1655 7789 1689
rect 7823 1655 7857 1689
rect 7891 1655 7925 1689
rect 7959 1655 7993 1689
rect 8027 1655 8061 1689
rect 8095 1655 8129 1689
rect 8163 1655 8197 1689
rect 8231 1655 8265 1689
rect 8299 1655 8333 1689
rect 8367 1655 8401 1689
rect 8435 1655 8469 1689
rect 8503 1655 8537 1689
rect 8571 1655 8605 1689
rect 8639 1655 8673 1689
rect 8707 1655 8741 1689
rect 8775 1655 8809 1689
rect 8843 1655 8877 1689
rect 8911 1655 8945 1689
rect 8979 1655 9013 1689
rect 9047 1655 9081 1689
rect 9115 1655 9149 1689
rect 9183 1655 9217 1689
rect 9251 1655 9285 1689
rect 9319 1655 9353 1689
rect 9387 1655 9421 1689
rect 9455 1655 9489 1689
rect 9523 1655 9557 1689
rect 9591 1655 9625 1689
rect 9659 1655 9693 1689
rect 9727 1655 9761 1689
rect 9795 1655 9829 1689
rect 9863 1655 9897 1689
rect 9931 1655 9965 1689
rect 9999 1655 10033 1689
rect 10067 1655 10101 1689
rect 10135 1655 10169 1689
rect 10203 1655 10237 1689
rect 10271 1655 10305 1689
rect 10339 1655 10373 1689
rect 10407 1655 10441 1689
rect 10475 1655 10509 1689
rect 10543 1655 10577 1689
rect 10611 1655 10645 1689
rect 10679 1655 10713 1689
rect 10747 1655 10781 1689
rect 10815 1655 10849 1689
rect 10883 1655 10917 1689
rect 10951 1655 10985 1689
rect 11019 1655 11053 1689
rect 11087 1655 11121 1689
rect 11155 1655 11189 1689
rect 11223 1655 11257 1689
rect 11291 1655 11325 1689
rect 11359 1655 11393 1689
rect 11427 1655 11461 1689
rect 11495 1655 11529 1689
rect 11563 1655 11597 1689
rect 11631 1655 11665 1689
rect 11699 1655 11733 1689
rect 11767 1655 11801 1689
rect 11835 1655 11869 1689
rect 11903 1655 11937 1689
rect 11971 1655 12005 1689
rect 12039 1655 12073 1689
rect 12107 1655 12141 1689
rect 12175 1655 12209 1689
rect 12243 1655 12277 1689
rect 12311 1655 12345 1689
rect 12379 1655 12413 1689
rect 12447 1655 12481 1689
rect 12515 1655 12549 1689
rect 12583 1655 12617 1689
rect 12651 1655 12685 1689
rect 12719 1655 12753 1689
rect 12787 1655 12821 1689
rect 12855 1655 12889 1689
rect 12923 1655 12957 1689
rect 12991 1655 13025 1689
rect 13059 1655 13093 1689
rect 13127 1655 13161 1689
rect 13195 1655 13229 1689
rect 13263 1655 13297 1689
rect 13331 1655 13365 1689
rect 13399 1655 13433 1689
rect 13467 1655 13501 1689
rect 13535 1655 13569 1689
rect 13603 1655 13637 1689
rect 13671 1655 13705 1689
rect 13739 1655 13773 1689
rect 13807 1655 13841 1689
rect 13875 1655 13909 1689
rect 13943 1655 13977 1689
rect 14011 1655 14045 1689
rect 14079 1655 14113 1689
rect 14147 1655 14181 1689
rect 14215 1655 14249 1689
rect 14283 1655 14317 1689
rect 14351 1655 14385 1689
rect 14419 1655 14453 1689
rect 14487 1655 14521 1689
rect 14555 1655 14589 1689
rect 14623 1655 14657 1689
rect 14691 1655 14725 1689
rect 14759 1655 14793 1689
rect 14827 1655 14861 1689
rect 14895 1655 14929 1689
rect 14963 1655 14997 1689
rect 15031 1655 15065 1689
rect 15099 1655 15133 1689
rect 15167 1655 15201 1689
rect 15235 1655 15269 1689
rect 15303 1655 15337 1689
rect 15371 1655 15405 1689
rect 15439 1655 15473 1689
rect 15507 1655 15541 1689
rect 15575 1655 15609 1689
rect 15643 1655 15677 1689
rect 15711 1655 15745 1689
rect 15779 1655 15813 1689
rect 15847 1655 15881 1689
rect 15915 1655 15949 1689
rect 15983 1655 16017 1689
rect 16051 1655 16085 1689
rect 16119 1655 16153 1689
rect 16187 1655 16221 1689
rect 16255 1655 16289 1689
rect 16323 1655 16357 1689
rect 16391 1655 16425 1689
rect 16459 1655 16493 1689
rect 16527 1655 16561 1689
rect 16595 1655 16629 1689
rect 16663 1655 16697 1689
rect 16731 1655 16765 1689
rect 16799 1655 16833 1689
rect 16867 1655 16901 1689
rect 16935 1655 16969 1689
rect 17003 1655 17037 1689
rect 17071 1655 17105 1689
rect 17139 1655 17173 1689
rect 17207 1655 17241 1689
rect 17275 1655 17309 1689
rect 17343 1655 17377 1689
rect 17411 1655 17445 1689
rect 17479 1655 17513 1689
rect 17547 1655 17581 1689
rect 17615 1655 17649 1689
rect 17683 1655 17717 1689
rect 17751 1655 17785 1689
rect 17819 1655 17853 1689
rect 17887 1655 17921 1689
rect 17955 1655 17989 1689
rect 18023 1655 18057 1689
rect 18091 1655 18125 1689
rect 18159 1655 18193 1689
rect 18227 1655 18261 1689
rect 18295 1655 18329 1689
rect 18363 1655 18397 1689
rect 18431 1655 18465 1689
rect 18499 1655 18533 1689
rect 18567 1655 18601 1689
rect 18635 1655 18669 1689
rect 18703 1655 18737 1689
rect 18771 1655 18805 1689
rect 18839 1655 18873 1689
rect 18907 1655 18941 1689
rect 18975 1655 19009 1689
rect 19043 1655 19077 1689
rect 19111 1655 19145 1689
rect 19179 1655 19213 1689
rect 19247 1655 19281 1689
rect 19315 1655 19349 1689
rect 19383 1655 19417 1689
rect 19451 1655 19485 1689
rect 19519 1655 19553 1689
rect 19587 1655 19621 1689
rect 19655 1655 19689 1689
rect 19723 1655 19757 1689
rect 19791 1655 19825 1689
rect 19859 1655 19893 1689
rect 19927 1655 19961 1689
rect 19995 1655 20029 1689
rect 20063 1655 20097 1689
rect 20131 1655 20165 1689
rect 20199 1655 20233 1689
rect 20267 1655 20301 1689
rect 20335 1655 20369 1689
rect 20403 1655 20437 1689
rect 20471 1655 20505 1689
rect 20539 1655 20573 1689
rect 20607 1655 20641 1689
rect 20675 1655 20709 1689
rect 20743 1655 20777 1689
rect 20811 1655 20845 1689
rect 20879 1655 20913 1689
rect 20947 1655 20981 1689
rect 21015 1655 21049 1689
rect 21083 1655 21117 1689
rect 21151 1655 21185 1689
rect 21219 1655 21253 1689
rect 21287 1655 21321 1689
rect 21355 1655 21389 1689
rect 21423 1655 21457 1689
rect 21491 1655 21525 1689
rect 21559 1655 21593 1689
rect 21627 1655 21661 1689
rect 21695 1655 21729 1689
rect 21763 1655 21797 1689
rect 21831 1655 21865 1689
rect 21899 1655 21933 1689
rect 21967 1655 22001 1689
rect 22035 1655 22069 1689
rect 22103 1655 22137 1689
rect 22171 1655 22205 1689
rect 22239 1655 22273 1689
rect 22307 1655 22341 1689
rect 22375 1655 22409 1689
rect 22443 1655 22477 1689
rect 22511 1655 22545 1689
rect 22579 1655 22613 1689
rect 22647 1655 22681 1689
rect 22715 1655 22749 1689
rect 22783 1655 22817 1689
rect 22851 1655 22885 1689
rect 22919 1655 22953 1689
rect 22987 1655 23021 1689
rect 23055 1655 23089 1689
rect 23123 1655 23157 1689
rect 23191 1655 23225 1689
rect 23259 1655 23293 1689
rect 23327 1655 23361 1689
rect 23395 1655 23429 1689
rect 23463 1655 23497 1689
rect 23531 1655 23565 1689
rect 23599 1655 23633 1689
rect 23667 1655 23701 1689
rect 23735 1655 23769 1689
rect 23803 1655 23837 1689
rect 23871 1655 23905 1689
rect 23939 1655 23973 1689
rect 24007 1655 24041 1689
rect 24075 1655 24109 1689
rect 24143 1655 24177 1689
rect 24211 1655 24245 1689
rect 24279 1655 24313 1689
rect 24347 1655 24381 1689
rect 24415 1655 24449 1689
rect 24483 1655 24517 1689
rect 24551 1655 24585 1689
rect 24619 1655 24653 1689
rect 411 1503 445 1537
rect 411 1435 445 1469
rect 411 1367 445 1401
rect 411 1299 445 1333
rect 411 1231 445 1265
rect 411 1163 445 1197
rect 411 1095 445 1129
rect 411 1027 445 1061
rect 411 959 445 993
rect 411 891 445 925
rect 411 823 445 857
rect 411 755 445 789
rect 411 687 445 721
rect 411 619 445 653
rect 411 551 445 585
rect 411 483 445 517
rect 411 415 445 449
rect 411 347 445 381
rect 411 279 445 313
rect 411 211 445 245
rect 411 143 445 177
rect 411 75 445 109
rect 411 7 445 41
rect 411 -61 445 -27
rect 411 -129 445 -95
rect 411 -197 445 -163
rect 411 -265 445 -231
rect 411 -333 445 -299
rect 411 -401 445 -367
rect 411 -469 445 -435
rect 411 -537 445 -503
rect 411 -605 445 -571
rect 411 -673 445 -639
rect 411 -741 445 -707
rect 411 -809 445 -775
rect 411 -877 445 -843
rect 411 -945 445 -911
rect 411 -1013 445 -979
rect 411 -1081 445 -1047
rect 411 -1149 445 -1115
rect 411 -1217 445 -1183
rect 411 -1285 445 -1251
rect 411 -1353 445 -1319
rect 411 -1421 445 -1387
rect 411 -1489 445 -1455
rect 411 -1557 445 -1523
rect 411 -1625 445 -1591
rect 411 -1693 445 -1659
rect 411 -1761 445 -1727
rect 411 -1829 445 -1795
rect 411 -1897 445 -1863
rect 411 -1965 445 -1931
rect 411 -2033 445 -1999
rect 411 -2101 445 -2067
rect 411 -2169 445 -2135
rect 411 -2237 445 -2203
rect 411 -2305 445 -2271
rect 411 -2373 445 -2339
rect 411 -2441 445 -2407
rect 411 -2509 445 -2475
rect 411 -2577 445 -2543
rect 411 -2645 445 -2611
rect 411 -2713 445 -2679
rect 411 -2781 445 -2747
rect 411 -2849 445 -2815
rect 411 -2917 445 -2883
rect 411 -2985 445 -2951
rect 411 -3053 445 -3019
rect 411 -3121 445 -3087
rect 411 -3189 445 -3155
rect 411 -3257 445 -3223
rect 411 -3325 445 -3291
rect 411 -3393 445 -3359
rect 411 -3461 445 -3427
rect 411 -3529 445 -3495
rect 411 -3597 445 -3563
rect 411 -3665 445 -3631
rect 411 -3733 445 -3699
rect 411 -3801 445 -3767
rect 411 -3869 445 -3835
rect 411 -3937 445 -3903
rect 411 -4005 445 -3971
rect 411 -4073 445 -4039
rect 411 -4141 445 -4107
rect 411 -4209 445 -4175
rect 411 -4277 445 -4243
rect 411 -4345 445 -4311
rect 411 -4413 445 -4379
rect 411 -4481 445 -4447
rect 411 -4549 445 -4515
rect 411 -4617 445 -4583
rect 24755 1503 24789 1537
rect 24755 1435 24789 1469
rect 24755 1367 24789 1401
rect 24755 1299 24789 1333
rect 24755 1231 24789 1265
rect 24755 1163 24789 1197
rect 24755 1095 24789 1129
rect 24755 1027 24789 1061
rect 24755 959 24789 993
rect 24755 891 24789 925
rect 24755 823 24789 857
rect 24755 755 24789 789
rect 24755 687 24789 721
rect 24755 619 24789 653
rect 24755 551 24789 585
rect 24755 483 24789 517
rect 24755 415 24789 449
rect 24755 347 24789 381
rect 24755 279 24789 313
rect 24755 211 24789 245
rect 24755 143 24789 177
rect 24755 75 24789 109
rect 24755 7 24789 41
rect 24755 -61 24789 -27
rect 24755 -129 24789 -95
rect 24755 -197 24789 -163
rect 24755 -265 24789 -231
rect 24755 -333 24789 -299
rect 24755 -401 24789 -367
rect 24755 -469 24789 -435
rect 24755 -537 24789 -503
rect 24755 -605 24789 -571
rect 24755 -673 24789 -639
rect 24755 -741 24789 -707
rect 24755 -809 24789 -775
rect 24755 -877 24789 -843
rect 24755 -945 24789 -911
rect 24755 -1013 24789 -979
rect 24755 -1081 24789 -1047
rect 24755 -1149 24789 -1115
rect 24755 -1217 24789 -1183
rect 24755 -1285 24789 -1251
rect 24755 -1353 24789 -1319
rect 24755 -1421 24789 -1387
rect 24755 -1489 24789 -1455
rect 24755 -1557 24789 -1523
rect 24755 -1625 24789 -1591
rect 24755 -1693 24789 -1659
rect 24755 -1761 24789 -1727
rect 24755 -1829 24789 -1795
rect 24755 -1897 24789 -1863
rect 24755 -1965 24789 -1931
rect 24755 -2033 24789 -1999
rect 24755 -2101 24789 -2067
rect 24755 -2169 24789 -2135
rect 24755 -2237 24789 -2203
rect 24755 -2305 24789 -2271
rect 24755 -2373 24789 -2339
rect 24755 -2441 24789 -2407
rect 24755 -2509 24789 -2475
rect 24755 -2577 24789 -2543
rect 24755 -2645 24789 -2611
rect 24755 -2713 24789 -2679
rect 24755 -2781 24789 -2747
rect 24755 -2849 24789 -2815
rect 24755 -2917 24789 -2883
rect 24755 -2985 24789 -2951
rect 24755 -3053 24789 -3019
rect 24755 -3121 24789 -3087
rect 24755 -3189 24789 -3155
rect 24755 -3257 24789 -3223
rect 24755 -3325 24789 -3291
rect 24755 -3393 24789 -3359
rect 24755 -3461 24789 -3427
rect 24755 -3529 24789 -3495
rect 24755 -3597 24789 -3563
rect 24755 -3665 24789 -3631
rect 24755 -3733 24789 -3699
rect 24755 -3801 24789 -3767
rect 24755 -3869 24789 -3835
rect 24755 -3937 24789 -3903
rect 24755 -4005 24789 -3971
rect 24755 -4073 24789 -4039
rect 24755 -4141 24789 -4107
rect 24755 -4209 24789 -4175
rect 24755 -4277 24789 -4243
rect 24755 -4345 24789 -4311
rect 24755 -4413 24789 -4379
rect 24755 -4481 24789 -4447
rect 24755 -4549 24789 -4515
rect 411 -4685 445 -4651
rect 24755 -4617 24789 -4583
rect 24755 -4685 24789 -4651
rect 411 -4753 445 -4719
rect 411 -4821 445 -4787
rect 411 -4889 445 -4855
rect 411 -4957 445 -4923
rect 411 -5025 445 -4991
rect 411 -5093 445 -5059
rect 24755 -4753 24789 -4719
rect 24755 -4821 24789 -4787
rect 24755 -4889 24789 -4855
rect 24755 -4957 24789 -4923
rect 24755 -5025 24789 -4991
rect 411 -5161 445 -5127
rect 24755 -5093 24789 -5059
rect 24755 -5161 24789 -5127
rect 411 -5229 445 -5195
rect 411 -5297 445 -5263
rect 411 -5365 445 -5331
rect 411 -5433 445 -5399
rect 411 -5501 445 -5467
rect 24755 -5229 24789 -5195
rect 24755 -5297 24789 -5263
rect 24755 -5365 24789 -5331
rect 24755 -5433 24789 -5399
rect 24755 -5501 24789 -5467
rect 411 -5569 445 -5535
rect 411 -5637 445 -5603
rect 24755 -5569 24789 -5535
rect 411 -5705 445 -5671
rect 411 -5773 445 -5739
rect 411 -5841 445 -5807
rect 411 -5909 445 -5875
rect 411 -5977 445 -5943
rect 411 -6045 445 -6011
rect 24755 -5637 24789 -5603
rect 24755 -5705 24789 -5671
rect 24755 -5773 24789 -5739
rect 24755 -5841 24789 -5807
rect 24755 -5909 24789 -5875
rect 24755 -5977 24789 -5943
rect 411 -6113 445 -6079
rect 24755 -6045 24789 -6011
rect 24755 -6113 24789 -6079
rect 411 -6181 445 -6147
rect 411 -6249 445 -6215
rect 411 -6317 445 -6283
rect 411 -6385 445 -6351
rect 411 -6453 445 -6419
rect 24755 -6181 24789 -6147
rect 24755 -6249 24789 -6215
rect 24755 -6317 24789 -6283
rect 24755 -6385 24789 -6351
rect 24755 -6453 24789 -6419
rect 411 -6521 445 -6487
rect 411 -6589 445 -6555
rect 24755 -6521 24789 -6487
rect 411 -6657 445 -6623
rect 411 -6725 445 -6691
rect 411 -6793 445 -6759
rect 411 -6861 445 -6827
rect 411 -6929 445 -6895
rect 411 -6997 445 -6963
rect 24755 -6589 24789 -6555
rect 24755 -6657 24789 -6623
rect 24755 -6725 24789 -6691
rect 24755 -6793 24789 -6759
rect 24755 -6861 24789 -6827
rect 24755 -6929 24789 -6895
rect 411 -7065 445 -7031
rect 24755 -6997 24789 -6963
rect 411 -7133 445 -7099
rect 411 -7201 445 -7167
rect 411 -7269 445 -7235
rect 411 -7337 445 -7303
rect 411 -7405 445 -7371
rect 24755 -7065 24789 -7031
rect 24755 -7133 24789 -7099
rect 24755 -7201 24789 -7167
rect 24755 -7269 24789 -7235
rect 24755 -7337 24789 -7303
rect 24755 -7405 24789 -7371
rect 411 -7473 445 -7439
rect 24755 -7473 24789 -7439
rect 411 -7541 445 -7507
rect 411 -7609 445 -7575
rect 411 -7677 445 -7643
rect 411 -7745 445 -7711
rect 411 -7813 445 -7779
rect 411 -7881 445 -7847
rect 24755 -7541 24789 -7507
rect 24755 -7609 24789 -7575
rect 24755 -7677 24789 -7643
rect 24755 -7745 24789 -7711
rect 24755 -7813 24789 -7779
rect 24755 -7881 24789 -7847
rect 411 -7949 445 -7915
rect 411 -8017 445 -7983
rect 24755 -7949 24789 -7915
rect 411 -8085 445 -8051
rect 411 -8153 445 -8119
rect 411 -8221 445 -8187
rect 411 -8289 445 -8255
rect 411 -8357 445 -8323
rect 411 -8425 445 -8391
rect 411 -8493 445 -8459
rect 411 -8561 445 -8527
rect 411 -8629 445 -8595
rect 411 -8697 445 -8663
rect 24755 -8017 24789 -7983
rect 24755 -8085 24789 -8051
rect 24755 -8153 24789 -8119
rect 24755 -8221 24789 -8187
rect 24755 -8289 24789 -8255
rect 24755 -8357 24789 -8323
rect 24755 -8425 24789 -8391
rect 24755 -8493 24789 -8459
rect 24755 -8561 24789 -8527
rect 24755 -8629 24789 -8595
rect 24755 -8697 24789 -8663
rect 547 -8849 581 -8815
rect 615 -8849 649 -8815
rect 683 -8849 717 -8815
rect 751 -8849 785 -8815
rect 819 -8849 853 -8815
rect 887 -8849 921 -8815
rect 955 -8849 989 -8815
rect 1023 -8849 1057 -8815
rect 1091 -8849 1125 -8815
rect 1159 -8849 1193 -8815
rect 1227 -8849 1261 -8815
rect 1295 -8849 1329 -8815
rect 1363 -8849 1397 -8815
rect 1431 -8849 1465 -8815
rect 1499 -8849 1533 -8815
rect 1567 -8849 1601 -8815
rect 1635 -8849 1669 -8815
rect 1703 -8849 1737 -8815
rect 1771 -8849 1805 -8815
rect 1839 -8849 1873 -8815
rect 1907 -8849 1941 -8815
rect 1975 -8849 2009 -8815
rect 2043 -8849 2077 -8815
rect 2111 -8849 2145 -8815
rect 2179 -8849 2213 -8815
rect 2247 -8849 2281 -8815
rect 2315 -8849 2349 -8815
rect 2383 -8849 2417 -8815
rect 2451 -8849 2485 -8815
rect 2519 -8849 2553 -8815
rect 2587 -8849 2621 -8815
rect 2655 -8849 2689 -8815
rect 2723 -8849 2757 -8815
rect 2791 -8849 2825 -8815
rect 2859 -8849 2893 -8815
rect 2927 -8849 2961 -8815
rect 2995 -8849 3029 -8815
rect 3063 -8849 3097 -8815
rect 3131 -8849 3165 -8815
rect 3199 -8849 3233 -8815
rect 3267 -8849 3301 -8815
rect 3335 -8849 3369 -8815
rect 3403 -8849 3437 -8815
rect 3471 -8849 3505 -8815
rect 3539 -8849 3573 -8815
rect 3607 -8849 3641 -8815
rect 3675 -8849 3709 -8815
rect 3743 -8849 3777 -8815
rect 3811 -8849 3845 -8815
rect 3879 -8849 3913 -8815
rect 3947 -8849 3981 -8815
rect 4015 -8849 4049 -8815
rect 4083 -8849 4117 -8815
rect 4151 -8849 4185 -8815
rect 4219 -8849 4253 -8815
rect 4287 -8849 4321 -8815
rect 4355 -8849 4389 -8815
rect 4423 -8849 4457 -8815
rect 4491 -8849 4525 -8815
rect 4559 -8849 4593 -8815
rect 4627 -8849 4661 -8815
rect 4695 -8849 4729 -8815
rect 4763 -8849 4797 -8815
rect 4831 -8849 4865 -8815
rect 4899 -8849 4933 -8815
rect 4967 -8849 5001 -8815
rect 5035 -8849 5069 -8815
rect 5103 -8849 5137 -8815
rect 5171 -8849 5205 -8815
rect 5239 -8849 5273 -8815
rect 5307 -8849 5341 -8815
rect 5375 -8849 5409 -8815
rect 5443 -8849 5477 -8815
rect 5511 -8849 5545 -8815
rect 5579 -8849 5613 -8815
rect 5647 -8849 5681 -8815
rect 5715 -8849 5749 -8815
rect 5783 -8849 5817 -8815
rect 5851 -8849 5885 -8815
rect 5919 -8849 5953 -8815
rect 5987 -8849 6021 -8815
rect 6055 -8849 6089 -8815
rect 6123 -8849 6157 -8815
rect 6191 -8849 6225 -8815
rect 6259 -8849 6293 -8815
rect 6327 -8849 6361 -8815
rect 6395 -8849 6429 -8815
rect 6463 -8849 6497 -8815
rect 6531 -8849 6565 -8815
rect 6599 -8849 6633 -8815
rect 6667 -8849 6701 -8815
rect 6735 -8849 6769 -8815
rect 6803 -8849 6837 -8815
rect 6871 -8849 6905 -8815
rect 6939 -8849 6973 -8815
rect 7007 -8849 7041 -8815
rect 7075 -8849 7109 -8815
rect 7143 -8849 7177 -8815
rect 7211 -8849 7245 -8815
rect 7279 -8849 7313 -8815
rect 7347 -8849 7381 -8815
rect 7415 -8849 7449 -8815
rect 7483 -8849 7517 -8815
rect 7551 -8849 7585 -8815
rect 7619 -8849 7653 -8815
rect 7687 -8849 7721 -8815
rect 7755 -8849 7789 -8815
rect 7823 -8849 7857 -8815
rect 7891 -8849 7925 -8815
rect 7959 -8849 7993 -8815
rect 8027 -8849 8061 -8815
rect 8095 -8849 8129 -8815
rect 8163 -8849 8197 -8815
rect 8231 -8849 8265 -8815
rect 8299 -8849 8333 -8815
rect 8367 -8849 8401 -8815
rect 8435 -8849 8469 -8815
rect 8503 -8849 8537 -8815
rect 8571 -8849 8605 -8815
rect 8639 -8849 8673 -8815
rect 8707 -8849 8741 -8815
rect 8775 -8849 8809 -8815
rect 8843 -8849 8877 -8815
rect 8911 -8849 8945 -8815
rect 8979 -8849 9013 -8815
rect 9047 -8849 9081 -8815
rect 9115 -8849 9149 -8815
rect 9183 -8849 9217 -8815
rect 9251 -8849 9285 -8815
rect 9319 -8849 9353 -8815
rect 9387 -8849 9421 -8815
rect 9455 -8849 9489 -8815
rect 9523 -8849 9557 -8815
rect 9591 -8849 9625 -8815
rect 9659 -8849 9693 -8815
rect 9727 -8849 9761 -8815
rect 9795 -8849 9829 -8815
rect 9863 -8849 9897 -8815
rect 9931 -8849 9965 -8815
rect 9999 -8849 10033 -8815
rect 10067 -8849 10101 -8815
rect 10135 -8849 10169 -8815
rect 10203 -8849 10237 -8815
rect 10271 -8849 10305 -8815
rect 10339 -8849 10373 -8815
rect 10407 -8849 10441 -8815
rect 10475 -8849 10509 -8815
rect 10543 -8849 10577 -8815
rect 10611 -8849 10645 -8815
rect 10679 -8849 10713 -8815
rect 10747 -8849 10781 -8815
rect 10815 -8849 10849 -8815
rect 10883 -8849 10917 -8815
rect 10951 -8849 10985 -8815
rect 11019 -8849 11053 -8815
rect 11087 -8849 11121 -8815
rect 11155 -8849 11189 -8815
rect 11223 -8849 11257 -8815
rect 11291 -8849 11325 -8815
rect 11359 -8849 11393 -8815
rect 11427 -8849 11461 -8815
rect 11495 -8849 11529 -8815
rect 11563 -8849 11597 -8815
rect 11631 -8849 11665 -8815
rect 11699 -8849 11733 -8815
rect 11767 -8849 11801 -8815
rect 11835 -8849 11869 -8815
rect 11903 -8849 11937 -8815
rect 11971 -8849 12005 -8815
rect 12039 -8849 12073 -8815
rect 12107 -8849 12141 -8815
rect 12175 -8849 12209 -8815
rect 12243 -8849 12277 -8815
rect 12311 -8849 12345 -8815
rect 12379 -8849 12413 -8815
rect 12447 -8849 12481 -8815
rect 12515 -8849 12549 -8815
rect 12583 -8849 12617 -8815
rect 12651 -8849 12685 -8815
rect 12719 -8849 12753 -8815
rect 12787 -8849 12821 -8815
rect 12855 -8849 12889 -8815
rect 12923 -8849 12957 -8815
rect 12991 -8849 13025 -8815
rect 13059 -8849 13093 -8815
rect 13127 -8849 13161 -8815
rect 13195 -8849 13229 -8815
rect 13263 -8849 13297 -8815
rect 13331 -8849 13365 -8815
rect 13399 -8849 13433 -8815
rect 13467 -8849 13501 -8815
rect 13535 -8849 13569 -8815
rect 13603 -8849 13637 -8815
rect 13671 -8849 13705 -8815
rect 13739 -8849 13773 -8815
rect 13807 -8849 13841 -8815
rect 13875 -8849 13909 -8815
rect 13943 -8849 13977 -8815
rect 14011 -8849 14045 -8815
rect 14079 -8849 14113 -8815
rect 14147 -8849 14181 -8815
rect 14215 -8849 14249 -8815
rect 14283 -8849 14317 -8815
rect 14351 -8849 14385 -8815
rect 14419 -8849 14453 -8815
rect 14487 -8849 14521 -8815
rect 14555 -8849 14589 -8815
rect 14623 -8849 14657 -8815
rect 14691 -8849 14725 -8815
rect 14759 -8849 14793 -8815
rect 14827 -8849 14861 -8815
rect 14895 -8849 14929 -8815
rect 14963 -8849 14997 -8815
rect 15031 -8849 15065 -8815
rect 15099 -8849 15133 -8815
rect 15167 -8849 15201 -8815
rect 15235 -8849 15269 -8815
rect 15303 -8849 15337 -8815
rect 15371 -8849 15405 -8815
rect 15439 -8849 15473 -8815
rect 15507 -8849 15541 -8815
rect 15575 -8849 15609 -8815
rect 15643 -8849 15677 -8815
rect 15711 -8849 15745 -8815
rect 15779 -8849 15813 -8815
rect 15847 -8849 15881 -8815
rect 15915 -8849 15949 -8815
rect 15983 -8849 16017 -8815
rect 16051 -8849 16085 -8815
rect 16119 -8849 16153 -8815
rect 16187 -8849 16221 -8815
rect 16255 -8849 16289 -8815
rect 16323 -8849 16357 -8815
rect 16391 -8849 16425 -8815
rect 16459 -8849 16493 -8815
rect 16527 -8849 16561 -8815
rect 16595 -8849 16629 -8815
rect 16663 -8849 16697 -8815
rect 16731 -8849 16765 -8815
rect 16799 -8849 16833 -8815
rect 16867 -8849 16901 -8815
rect 16935 -8849 16969 -8815
rect 17003 -8849 17037 -8815
rect 17071 -8849 17105 -8815
rect 17139 -8849 17173 -8815
rect 17207 -8849 17241 -8815
rect 17275 -8849 17309 -8815
rect 17343 -8849 17377 -8815
rect 17411 -8849 17445 -8815
rect 17479 -8849 17513 -8815
rect 17547 -8849 17581 -8815
rect 17615 -8849 17649 -8815
rect 17683 -8849 17717 -8815
rect 17751 -8849 17785 -8815
rect 17819 -8849 17853 -8815
rect 17887 -8849 17921 -8815
rect 17955 -8849 17989 -8815
rect 18023 -8849 18057 -8815
rect 18091 -8849 18125 -8815
rect 18159 -8849 18193 -8815
rect 18227 -8849 18261 -8815
rect 18295 -8849 18329 -8815
rect 18363 -8849 18397 -8815
rect 18431 -8849 18465 -8815
rect 18499 -8849 18533 -8815
rect 18567 -8849 18601 -8815
rect 18635 -8849 18669 -8815
rect 18703 -8849 18737 -8815
rect 18771 -8849 18805 -8815
rect 18839 -8849 18873 -8815
rect 18907 -8849 18941 -8815
rect 18975 -8849 19009 -8815
rect 19043 -8849 19077 -8815
rect 19111 -8849 19145 -8815
rect 19179 -8849 19213 -8815
rect 19247 -8849 19281 -8815
rect 19315 -8849 19349 -8815
rect 19383 -8849 19417 -8815
rect 19451 -8849 19485 -8815
rect 19519 -8849 19553 -8815
rect 19587 -8849 19621 -8815
rect 19655 -8849 19689 -8815
rect 19723 -8849 19757 -8815
rect 19791 -8849 19825 -8815
rect 19859 -8849 19893 -8815
rect 19927 -8849 19961 -8815
rect 19995 -8849 20029 -8815
rect 20063 -8849 20097 -8815
rect 20131 -8849 20165 -8815
rect 20199 -8849 20233 -8815
rect 20267 -8849 20301 -8815
rect 20335 -8849 20369 -8815
rect 20403 -8849 20437 -8815
rect 20471 -8849 20505 -8815
rect 20539 -8849 20573 -8815
rect 20607 -8849 20641 -8815
rect 20675 -8849 20709 -8815
rect 20743 -8849 20777 -8815
rect 20811 -8849 20845 -8815
rect 20879 -8849 20913 -8815
rect 20947 -8849 20981 -8815
rect 21015 -8849 21049 -8815
rect 21083 -8849 21117 -8815
rect 21151 -8849 21185 -8815
rect 21219 -8849 21253 -8815
rect 21287 -8849 21321 -8815
rect 21355 -8849 21389 -8815
rect 21423 -8849 21457 -8815
rect 21491 -8849 21525 -8815
rect 21559 -8849 21593 -8815
rect 21627 -8849 21661 -8815
rect 21695 -8849 21729 -8815
rect 21763 -8849 21797 -8815
rect 21831 -8849 21865 -8815
rect 21899 -8849 21933 -8815
rect 21967 -8849 22001 -8815
rect 22035 -8849 22069 -8815
rect 22103 -8849 22137 -8815
rect 22171 -8849 22205 -8815
rect 22239 -8849 22273 -8815
rect 22307 -8849 22341 -8815
rect 22375 -8849 22409 -8815
rect 22443 -8849 22477 -8815
rect 22511 -8849 22545 -8815
rect 22579 -8849 22613 -8815
rect 22647 -8849 22681 -8815
rect 22715 -8849 22749 -8815
rect 22783 -8849 22817 -8815
rect 22851 -8849 22885 -8815
rect 22919 -8849 22953 -8815
rect 22987 -8849 23021 -8815
rect 23055 -8849 23089 -8815
rect 23123 -8849 23157 -8815
rect 23191 -8849 23225 -8815
rect 23259 -8849 23293 -8815
rect 23327 -8849 23361 -8815
rect 23395 -8849 23429 -8815
rect 23463 -8849 23497 -8815
rect 23531 -8849 23565 -8815
rect 23599 -8849 23633 -8815
rect 23667 -8849 23701 -8815
rect 23735 -8849 23769 -8815
rect 23803 -8849 23837 -8815
rect 23871 -8849 23905 -8815
rect 23939 -8849 23973 -8815
rect 24007 -8849 24041 -8815
rect 24075 -8849 24109 -8815
rect 24143 -8849 24177 -8815
rect 24211 -8849 24245 -8815
rect 24279 -8849 24313 -8815
rect 24347 -8849 24381 -8815
rect 24415 -8849 24449 -8815
rect 24483 -8849 24517 -8815
rect 24551 -8849 24585 -8815
rect 24619 -8849 24653 -8815
<< poly >>
rect 3698 -4609 3806 -4593
rect 3698 -4626 3735 -4609
rect 3672 -4643 3735 -4626
rect 3769 -4626 3806 -4609
rect 3916 -4609 4024 -4593
rect 3916 -4626 3953 -4609
rect 3769 -4643 3832 -4626
rect 3672 -4690 3832 -4643
rect 3890 -4643 3953 -4626
rect 3987 -4626 4024 -4609
rect 4134 -4609 4242 -4593
rect 4134 -4626 4171 -4609
rect 3987 -4643 4050 -4626
rect 3890 -4690 4050 -4643
rect 4108 -4643 4171 -4626
rect 4205 -4626 4242 -4609
rect 4352 -4609 4460 -4593
rect 4352 -4626 4389 -4609
rect 4205 -4643 4268 -4626
rect 4108 -4690 4268 -4643
rect 4326 -4643 4389 -4626
rect 4423 -4626 4460 -4609
rect 4570 -4609 4678 -4593
rect 4570 -4626 4607 -4609
rect 4423 -4643 4486 -4626
rect 4326 -4690 4486 -4643
rect 4544 -4643 4607 -4626
rect 4641 -4626 4678 -4609
rect 4788 -4609 4896 -4593
rect 4788 -4626 4825 -4609
rect 4641 -4643 4704 -4626
rect 4544 -4690 4704 -4643
rect 4762 -4643 4825 -4626
rect 4859 -4626 4896 -4609
rect 5006 -4609 5114 -4593
rect 5006 -4626 5043 -4609
rect 4859 -4643 4922 -4626
rect 4762 -4690 4922 -4643
rect 4980 -4643 5043 -4626
rect 5077 -4626 5114 -4609
rect 5224 -4609 5332 -4593
rect 5224 -4626 5261 -4609
rect 5077 -4643 5140 -4626
rect 4980 -4690 5140 -4643
rect 5198 -4643 5261 -4626
rect 5295 -4626 5332 -4609
rect 5442 -4609 5550 -4593
rect 5442 -4626 5479 -4609
rect 5295 -4643 5358 -4626
rect 5198 -4690 5358 -4643
rect 5416 -4643 5479 -4626
rect 5513 -4626 5550 -4609
rect 5660 -4609 5768 -4593
rect 5660 -4626 5697 -4609
rect 5513 -4643 5576 -4626
rect 5416 -4690 5576 -4643
rect 5634 -4643 5697 -4626
rect 5731 -4626 5768 -4609
rect 5731 -4643 5794 -4626
rect 5634 -4690 5794 -4643
rect 3672 -5137 3832 -5090
rect 3672 -5154 3735 -5137
rect 3698 -5171 3735 -5154
rect 3769 -5154 3832 -5137
rect 3890 -5137 4050 -5090
rect 3890 -5154 3953 -5137
rect 3769 -5171 3806 -5154
rect 3698 -5187 3806 -5171
rect 3916 -5171 3953 -5154
rect 3987 -5154 4050 -5137
rect 4108 -5137 4268 -5090
rect 4108 -5154 4171 -5137
rect 3987 -5171 4024 -5154
rect 3916 -5187 4024 -5171
rect 4134 -5171 4171 -5154
rect 4205 -5154 4268 -5137
rect 4326 -5137 4486 -5090
rect 4326 -5154 4389 -5137
rect 4205 -5171 4242 -5154
rect 4134 -5187 4242 -5171
rect 4352 -5171 4389 -5154
rect 4423 -5154 4486 -5137
rect 4544 -5137 4704 -5090
rect 4544 -5154 4607 -5137
rect 4423 -5171 4460 -5154
rect 4352 -5187 4460 -5171
rect 4570 -5171 4607 -5154
rect 4641 -5154 4704 -5137
rect 4762 -5137 4922 -5090
rect 4762 -5154 4825 -5137
rect 4641 -5171 4678 -5154
rect 4570 -5187 4678 -5171
rect 4788 -5171 4825 -5154
rect 4859 -5154 4922 -5137
rect 4980 -5137 5140 -5090
rect 4980 -5154 5043 -5137
rect 4859 -5171 4896 -5154
rect 4788 -5187 4896 -5171
rect 5006 -5171 5043 -5154
rect 5077 -5154 5140 -5137
rect 5198 -5137 5358 -5090
rect 5198 -5154 5261 -5137
rect 5077 -5171 5114 -5154
rect 5006 -5187 5114 -5171
rect 5224 -5171 5261 -5154
rect 5295 -5154 5358 -5137
rect 5416 -5137 5576 -5090
rect 5416 -5154 5479 -5137
rect 5295 -5171 5332 -5154
rect 5224 -5187 5332 -5171
rect 5442 -5171 5479 -5154
rect 5513 -5154 5576 -5137
rect 5634 -5137 5794 -5090
rect 5634 -5154 5697 -5137
rect 5513 -5171 5550 -5154
rect 5442 -5187 5550 -5171
rect 5660 -5171 5697 -5154
rect 5731 -5154 5794 -5137
rect 5731 -5171 5768 -5154
rect 5660 -5187 5768 -5171
rect 3698 -5547 3806 -5531
rect 3698 -5564 3735 -5547
rect 3672 -5581 3735 -5564
rect 3769 -5564 3806 -5547
rect 3916 -5547 4024 -5531
rect 3916 -5564 3953 -5547
rect 3769 -5581 3832 -5564
rect 3672 -5628 3832 -5581
rect 3890 -5581 3953 -5564
rect 3987 -5564 4024 -5547
rect 4134 -5547 4242 -5531
rect 4134 -5564 4171 -5547
rect 3987 -5581 4050 -5564
rect 3890 -5628 4050 -5581
rect 4108 -5581 4171 -5564
rect 4205 -5564 4242 -5547
rect 4352 -5547 4460 -5531
rect 4352 -5564 4389 -5547
rect 4205 -5581 4268 -5564
rect 4108 -5628 4268 -5581
rect 4326 -5581 4389 -5564
rect 4423 -5564 4460 -5547
rect 4570 -5547 4678 -5531
rect 4570 -5564 4607 -5547
rect 4423 -5581 4486 -5564
rect 4326 -5628 4486 -5581
rect 4544 -5581 4607 -5564
rect 4641 -5564 4678 -5547
rect 4788 -5547 4896 -5531
rect 4788 -5564 4825 -5547
rect 4641 -5581 4704 -5564
rect 4544 -5628 4704 -5581
rect 4762 -5581 4825 -5564
rect 4859 -5564 4896 -5547
rect 5006 -5547 5114 -5531
rect 5006 -5564 5043 -5547
rect 4859 -5581 4922 -5564
rect 4762 -5628 4922 -5581
rect 4980 -5581 5043 -5564
rect 5077 -5564 5114 -5547
rect 5224 -5547 5332 -5531
rect 5224 -5564 5261 -5547
rect 5077 -5581 5140 -5564
rect 4980 -5628 5140 -5581
rect 5198 -5581 5261 -5564
rect 5295 -5564 5332 -5547
rect 5442 -5547 5550 -5531
rect 5442 -5564 5479 -5547
rect 5295 -5581 5358 -5564
rect 5198 -5628 5358 -5581
rect 5416 -5581 5479 -5564
rect 5513 -5564 5550 -5547
rect 5660 -5547 5768 -5531
rect 5660 -5564 5697 -5547
rect 5513 -5581 5576 -5564
rect 5416 -5628 5576 -5581
rect 5634 -5581 5697 -5564
rect 5731 -5564 5768 -5547
rect 5731 -5581 5794 -5564
rect 5634 -5628 5794 -5581
rect 3672 -6075 3832 -6028
rect 3672 -6092 3735 -6075
rect 3698 -6109 3735 -6092
rect 3769 -6092 3832 -6075
rect 3890 -6075 4050 -6028
rect 3890 -6092 3953 -6075
rect 3769 -6109 3806 -6092
rect 3698 -6125 3806 -6109
rect 3916 -6109 3953 -6092
rect 3987 -6092 4050 -6075
rect 4108 -6075 4268 -6028
rect 4108 -6092 4171 -6075
rect 3987 -6109 4024 -6092
rect 3916 -6125 4024 -6109
rect 4134 -6109 4171 -6092
rect 4205 -6092 4268 -6075
rect 4326 -6075 4486 -6028
rect 4326 -6092 4389 -6075
rect 4205 -6109 4242 -6092
rect 4134 -6125 4242 -6109
rect 4352 -6109 4389 -6092
rect 4423 -6092 4486 -6075
rect 4544 -6075 4704 -6028
rect 4544 -6092 4607 -6075
rect 4423 -6109 4460 -6092
rect 4352 -6125 4460 -6109
rect 4570 -6109 4607 -6092
rect 4641 -6092 4704 -6075
rect 4762 -6075 4922 -6028
rect 4762 -6092 4825 -6075
rect 4641 -6109 4678 -6092
rect 4570 -6125 4678 -6109
rect 4788 -6109 4825 -6092
rect 4859 -6092 4922 -6075
rect 4980 -6075 5140 -6028
rect 4980 -6092 5043 -6075
rect 4859 -6109 4896 -6092
rect 4788 -6125 4896 -6109
rect 5006 -6109 5043 -6092
rect 5077 -6092 5140 -6075
rect 5198 -6075 5358 -6028
rect 5198 -6092 5261 -6075
rect 5077 -6109 5114 -6092
rect 5006 -6125 5114 -6109
rect 5224 -6109 5261 -6092
rect 5295 -6092 5358 -6075
rect 5416 -6075 5576 -6028
rect 5416 -6092 5479 -6075
rect 5295 -6109 5332 -6092
rect 5224 -6125 5332 -6109
rect 5442 -6109 5479 -6092
rect 5513 -6092 5576 -6075
rect 5634 -6075 5794 -6028
rect 5634 -6092 5697 -6075
rect 5513 -6109 5550 -6092
rect 5442 -6125 5550 -6109
rect 5660 -6109 5697 -6092
rect 5731 -6092 5794 -6075
rect 5731 -6109 5768 -6092
rect 5660 -6125 5768 -6109
rect 3698 -6485 3806 -6469
rect 3698 -6502 3735 -6485
rect 3672 -6519 3735 -6502
rect 3769 -6502 3806 -6485
rect 3916 -6485 4024 -6469
rect 3916 -6502 3953 -6485
rect 3769 -6519 3832 -6502
rect 3672 -6566 3832 -6519
rect 3890 -6519 3953 -6502
rect 3987 -6502 4024 -6485
rect 4134 -6485 4242 -6469
rect 4134 -6502 4171 -6485
rect 3987 -6519 4050 -6502
rect 3890 -6566 4050 -6519
rect 4108 -6519 4171 -6502
rect 4205 -6502 4242 -6485
rect 4352 -6485 4460 -6469
rect 4352 -6502 4389 -6485
rect 4205 -6519 4268 -6502
rect 4108 -6566 4268 -6519
rect 4326 -6519 4389 -6502
rect 4423 -6502 4460 -6485
rect 4570 -6485 4678 -6469
rect 4570 -6502 4607 -6485
rect 4423 -6519 4486 -6502
rect 4326 -6566 4486 -6519
rect 4544 -6519 4607 -6502
rect 4641 -6502 4678 -6485
rect 4788 -6485 4896 -6469
rect 4788 -6502 4825 -6485
rect 4641 -6519 4704 -6502
rect 4544 -6566 4704 -6519
rect 4762 -6519 4825 -6502
rect 4859 -6502 4896 -6485
rect 5006 -6485 5114 -6469
rect 5006 -6502 5043 -6485
rect 4859 -6519 4922 -6502
rect 4762 -6566 4922 -6519
rect 4980 -6519 5043 -6502
rect 5077 -6502 5114 -6485
rect 5224 -6485 5332 -6469
rect 5224 -6502 5261 -6485
rect 5077 -6519 5140 -6502
rect 4980 -6566 5140 -6519
rect 5198 -6519 5261 -6502
rect 5295 -6502 5332 -6485
rect 5442 -6485 5550 -6469
rect 5442 -6502 5479 -6485
rect 5295 -6519 5358 -6502
rect 5198 -6566 5358 -6519
rect 5416 -6519 5479 -6502
rect 5513 -6502 5550 -6485
rect 5660 -6485 5768 -6469
rect 5660 -6502 5697 -6485
rect 5513 -6519 5576 -6502
rect 5416 -6566 5576 -6519
rect 5634 -6519 5697 -6502
rect 5731 -6502 5768 -6485
rect 5731 -6519 5794 -6502
rect 5634 -6566 5794 -6519
rect 3672 -7013 3832 -6966
rect 3672 -7030 3735 -7013
rect 3698 -7047 3735 -7030
rect 3769 -7030 3832 -7013
rect 3890 -7013 4050 -6966
rect 3890 -7030 3953 -7013
rect 3769 -7047 3806 -7030
rect 3698 -7063 3806 -7047
rect 3916 -7047 3953 -7030
rect 3987 -7030 4050 -7013
rect 4108 -7013 4268 -6966
rect 4108 -7030 4171 -7013
rect 3987 -7047 4024 -7030
rect 3916 -7063 4024 -7047
rect 4134 -7047 4171 -7030
rect 4205 -7030 4268 -7013
rect 4326 -7013 4486 -6966
rect 4326 -7030 4389 -7013
rect 4205 -7047 4242 -7030
rect 4134 -7063 4242 -7047
rect 4352 -7047 4389 -7030
rect 4423 -7030 4486 -7013
rect 4544 -7013 4704 -6966
rect 4544 -7030 4607 -7013
rect 4423 -7047 4460 -7030
rect 4352 -7063 4460 -7047
rect 4570 -7047 4607 -7030
rect 4641 -7030 4704 -7013
rect 4762 -7013 4922 -6966
rect 4762 -7030 4825 -7013
rect 4641 -7047 4678 -7030
rect 4570 -7063 4678 -7047
rect 4788 -7047 4825 -7030
rect 4859 -7030 4922 -7013
rect 4980 -7013 5140 -6966
rect 4980 -7030 5043 -7013
rect 4859 -7047 4896 -7030
rect 4788 -7063 4896 -7047
rect 5006 -7047 5043 -7030
rect 5077 -7030 5140 -7013
rect 5198 -7013 5358 -6966
rect 5198 -7030 5261 -7013
rect 5077 -7047 5114 -7030
rect 5006 -7063 5114 -7047
rect 5224 -7047 5261 -7030
rect 5295 -7030 5358 -7013
rect 5416 -7013 5576 -6966
rect 5416 -7030 5479 -7013
rect 5295 -7047 5332 -7030
rect 5224 -7063 5332 -7047
rect 5442 -7047 5479 -7030
rect 5513 -7030 5576 -7013
rect 5634 -7013 5794 -6966
rect 5634 -7030 5697 -7013
rect 5513 -7047 5550 -7030
rect 5442 -7063 5550 -7047
rect 5660 -7047 5697 -7030
rect 5731 -7030 5794 -7013
rect 5731 -7047 5768 -7030
rect 5660 -7063 5768 -7047
rect 3698 -7423 3806 -7407
rect 3698 -7440 3735 -7423
rect 3672 -7457 3735 -7440
rect 3769 -7440 3806 -7423
rect 3916 -7423 4024 -7407
rect 3916 -7440 3953 -7423
rect 3769 -7457 3832 -7440
rect 3672 -7504 3832 -7457
rect 3890 -7457 3953 -7440
rect 3987 -7440 4024 -7423
rect 4134 -7423 4242 -7407
rect 4134 -7440 4171 -7423
rect 3987 -7457 4050 -7440
rect 3890 -7504 4050 -7457
rect 4108 -7457 4171 -7440
rect 4205 -7440 4242 -7423
rect 4352 -7423 4460 -7407
rect 4352 -7440 4389 -7423
rect 4205 -7457 4268 -7440
rect 4108 -7504 4268 -7457
rect 4326 -7457 4389 -7440
rect 4423 -7440 4460 -7423
rect 4570 -7423 4678 -7407
rect 4570 -7440 4607 -7423
rect 4423 -7457 4486 -7440
rect 4326 -7504 4486 -7457
rect 4544 -7457 4607 -7440
rect 4641 -7440 4678 -7423
rect 4788 -7423 4896 -7407
rect 4788 -7440 4825 -7423
rect 4641 -7457 4704 -7440
rect 4544 -7504 4704 -7457
rect 4762 -7457 4825 -7440
rect 4859 -7440 4896 -7423
rect 5006 -7423 5114 -7407
rect 5006 -7440 5043 -7423
rect 4859 -7457 4922 -7440
rect 4762 -7504 4922 -7457
rect 4980 -7457 5043 -7440
rect 5077 -7440 5114 -7423
rect 5224 -7423 5332 -7407
rect 5224 -7440 5261 -7423
rect 5077 -7457 5140 -7440
rect 4980 -7504 5140 -7457
rect 5198 -7457 5261 -7440
rect 5295 -7440 5332 -7423
rect 5442 -7423 5550 -7407
rect 5442 -7440 5479 -7423
rect 5295 -7457 5358 -7440
rect 5198 -7504 5358 -7457
rect 5416 -7457 5479 -7440
rect 5513 -7440 5550 -7423
rect 5660 -7423 5768 -7407
rect 5660 -7440 5697 -7423
rect 5513 -7457 5576 -7440
rect 5416 -7504 5576 -7457
rect 5634 -7457 5697 -7440
rect 5731 -7440 5768 -7423
rect 5731 -7457 5794 -7440
rect 5634 -7504 5794 -7457
rect 3672 -7951 3832 -7904
rect 3672 -7968 3735 -7951
rect 3698 -7985 3735 -7968
rect 3769 -7968 3832 -7951
rect 3890 -7951 4050 -7904
rect 3890 -7968 3953 -7951
rect 3769 -7985 3806 -7968
rect 3698 -8001 3806 -7985
rect 3916 -7985 3953 -7968
rect 3987 -7968 4050 -7951
rect 4108 -7951 4268 -7904
rect 4108 -7968 4171 -7951
rect 3987 -7985 4024 -7968
rect 3916 -8001 4024 -7985
rect 4134 -7985 4171 -7968
rect 4205 -7968 4268 -7951
rect 4326 -7951 4486 -7904
rect 4326 -7968 4389 -7951
rect 4205 -7985 4242 -7968
rect 4134 -8001 4242 -7985
rect 4352 -7985 4389 -7968
rect 4423 -7968 4486 -7951
rect 4544 -7951 4704 -7904
rect 4544 -7968 4607 -7951
rect 4423 -7985 4460 -7968
rect 4352 -8001 4460 -7985
rect 4570 -7985 4607 -7968
rect 4641 -7968 4704 -7951
rect 4762 -7951 4922 -7904
rect 4762 -7968 4825 -7951
rect 4641 -7985 4678 -7968
rect 4570 -8001 4678 -7985
rect 4788 -7985 4825 -7968
rect 4859 -7968 4922 -7951
rect 4980 -7951 5140 -7904
rect 4980 -7968 5043 -7951
rect 4859 -7985 4896 -7968
rect 4788 -8001 4896 -7985
rect 5006 -7985 5043 -7968
rect 5077 -7968 5140 -7951
rect 5198 -7951 5358 -7904
rect 5198 -7968 5261 -7951
rect 5077 -7985 5114 -7968
rect 5006 -8001 5114 -7985
rect 5224 -7985 5261 -7968
rect 5295 -7968 5358 -7951
rect 5416 -7951 5576 -7904
rect 5416 -7968 5479 -7951
rect 5295 -7985 5332 -7968
rect 5224 -8001 5332 -7985
rect 5442 -7985 5479 -7968
rect 5513 -7968 5576 -7951
rect 5634 -7951 5794 -7904
rect 5634 -7968 5697 -7951
rect 5513 -7985 5550 -7968
rect 5442 -8001 5550 -7985
rect 5660 -7985 5697 -7968
rect 5731 -7968 5794 -7951
rect 5731 -7985 5768 -7968
rect 5660 -8001 5768 -7985
rect 2814 -11646 3402 -11630
rect 2814 -11663 2853 -11646
rect 2628 -11680 2853 -11663
rect 2887 -11680 2921 -11646
rect 2955 -11680 2989 -11646
rect 3023 -11680 3057 -11646
rect 3091 -11680 3125 -11646
rect 3159 -11680 3193 -11646
rect 3227 -11680 3261 -11646
rect 3295 -11680 3329 -11646
rect 3363 -11663 3402 -11646
rect 3832 -11646 4420 -11630
rect 3832 -11663 3871 -11646
rect 3363 -11680 3588 -11663
rect 2628 -11718 3588 -11680
rect 3646 -11680 3871 -11663
rect 3905 -11680 3939 -11646
rect 3973 -11680 4007 -11646
rect 4041 -11680 4075 -11646
rect 4109 -11680 4143 -11646
rect 4177 -11680 4211 -11646
rect 4245 -11680 4279 -11646
rect 4313 -11680 4347 -11646
rect 4381 -11663 4420 -11646
rect 4850 -11646 5438 -11630
rect 4850 -11663 4889 -11646
rect 4381 -11680 4606 -11663
rect 3646 -11718 4606 -11680
rect 4664 -11680 4889 -11663
rect 4923 -11680 4957 -11646
rect 4991 -11680 5025 -11646
rect 5059 -11680 5093 -11646
rect 5127 -11680 5161 -11646
rect 5195 -11680 5229 -11646
rect 5263 -11680 5297 -11646
rect 5331 -11680 5365 -11646
rect 5399 -11663 5438 -11646
rect 5868 -11646 6456 -11630
rect 5868 -11663 5907 -11646
rect 5399 -11680 5624 -11663
rect 4664 -11718 5624 -11680
rect 5682 -11680 5907 -11663
rect 5941 -11680 5975 -11646
rect 6009 -11680 6043 -11646
rect 6077 -11680 6111 -11646
rect 6145 -11680 6179 -11646
rect 6213 -11680 6247 -11646
rect 6281 -11680 6315 -11646
rect 6349 -11680 6383 -11646
rect 6417 -11663 6456 -11646
rect 6886 -11646 7474 -11630
rect 6886 -11663 6925 -11646
rect 6417 -11680 6642 -11663
rect 5682 -11718 6642 -11680
rect 6700 -11680 6925 -11663
rect 6959 -11680 6993 -11646
rect 7027 -11680 7061 -11646
rect 7095 -11680 7129 -11646
rect 7163 -11680 7197 -11646
rect 7231 -11680 7265 -11646
rect 7299 -11680 7333 -11646
rect 7367 -11680 7401 -11646
rect 7435 -11663 7474 -11646
rect 7904 -11646 8492 -11630
rect 7904 -11663 7943 -11646
rect 7435 -11680 7660 -11663
rect 6700 -11718 7660 -11680
rect 7718 -11680 7943 -11663
rect 7977 -11680 8011 -11646
rect 8045 -11680 8079 -11646
rect 8113 -11680 8147 -11646
rect 8181 -11680 8215 -11646
rect 8249 -11680 8283 -11646
rect 8317 -11680 8351 -11646
rect 8385 -11680 8419 -11646
rect 8453 -11663 8492 -11646
rect 8922 -11646 9510 -11630
rect 8922 -11663 8961 -11646
rect 8453 -11680 8678 -11663
rect 7718 -11718 8678 -11680
rect 8736 -11680 8961 -11663
rect 8995 -11680 9029 -11646
rect 9063 -11680 9097 -11646
rect 9131 -11680 9165 -11646
rect 9199 -11680 9233 -11646
rect 9267 -11680 9301 -11646
rect 9335 -11680 9369 -11646
rect 9403 -11680 9437 -11646
rect 9471 -11663 9510 -11646
rect 9940 -11646 10528 -11630
rect 9940 -11663 9979 -11646
rect 9471 -11680 9696 -11663
rect 8736 -11718 9696 -11680
rect 9754 -11680 9979 -11663
rect 10013 -11680 10047 -11646
rect 10081 -11680 10115 -11646
rect 10149 -11680 10183 -11646
rect 10217 -11680 10251 -11646
rect 10285 -11680 10319 -11646
rect 10353 -11680 10387 -11646
rect 10421 -11680 10455 -11646
rect 10489 -11663 10528 -11646
rect 10958 -11646 11546 -11630
rect 10958 -11663 10997 -11646
rect 10489 -11680 10714 -11663
rect 9754 -11718 10714 -11680
rect 10772 -11680 10997 -11663
rect 11031 -11680 11065 -11646
rect 11099 -11680 11133 -11646
rect 11167 -11680 11201 -11646
rect 11235 -11680 11269 -11646
rect 11303 -11680 11337 -11646
rect 11371 -11680 11405 -11646
rect 11439 -11680 11473 -11646
rect 11507 -11663 11546 -11646
rect 11976 -11646 12564 -11630
rect 11976 -11663 12015 -11646
rect 11507 -11680 11732 -11663
rect 10772 -11718 11732 -11680
rect 11790 -11680 12015 -11663
rect 12049 -11680 12083 -11646
rect 12117 -11680 12151 -11646
rect 12185 -11680 12219 -11646
rect 12253 -11680 12287 -11646
rect 12321 -11680 12355 -11646
rect 12389 -11680 12423 -11646
rect 12457 -11680 12491 -11646
rect 12525 -11663 12564 -11646
rect 12994 -11646 13582 -11630
rect 12994 -11663 13033 -11646
rect 12525 -11680 12750 -11663
rect 11790 -11718 12750 -11680
rect 12808 -11680 13033 -11663
rect 13067 -11680 13101 -11646
rect 13135 -11680 13169 -11646
rect 13203 -11680 13237 -11646
rect 13271 -11680 13305 -11646
rect 13339 -11680 13373 -11646
rect 13407 -11680 13441 -11646
rect 13475 -11680 13509 -11646
rect 13543 -11663 13582 -11646
rect 14012 -11646 14600 -11630
rect 14012 -11663 14051 -11646
rect 13543 -11680 13768 -11663
rect 12808 -11718 13768 -11680
rect 13826 -11680 14051 -11663
rect 14085 -11680 14119 -11646
rect 14153 -11680 14187 -11646
rect 14221 -11680 14255 -11646
rect 14289 -11680 14323 -11646
rect 14357 -11680 14391 -11646
rect 14425 -11680 14459 -11646
rect 14493 -11680 14527 -11646
rect 14561 -11663 14600 -11646
rect 15030 -11646 15618 -11630
rect 15030 -11663 15069 -11646
rect 14561 -11680 14786 -11663
rect 13826 -11718 14786 -11680
rect 14844 -11680 15069 -11663
rect 15103 -11680 15137 -11646
rect 15171 -11680 15205 -11646
rect 15239 -11680 15273 -11646
rect 15307 -11680 15341 -11646
rect 15375 -11680 15409 -11646
rect 15443 -11680 15477 -11646
rect 15511 -11680 15545 -11646
rect 15579 -11663 15618 -11646
rect 16048 -11646 16636 -11630
rect 16048 -11663 16087 -11646
rect 15579 -11680 15804 -11663
rect 14844 -11718 15804 -11680
rect 15862 -11680 16087 -11663
rect 16121 -11680 16155 -11646
rect 16189 -11680 16223 -11646
rect 16257 -11680 16291 -11646
rect 16325 -11680 16359 -11646
rect 16393 -11680 16427 -11646
rect 16461 -11680 16495 -11646
rect 16529 -11680 16563 -11646
rect 16597 -11663 16636 -11646
rect 17066 -11646 17654 -11630
rect 17066 -11663 17105 -11646
rect 16597 -11680 16822 -11663
rect 15862 -11718 16822 -11680
rect 16880 -11680 17105 -11663
rect 17139 -11680 17173 -11646
rect 17207 -11680 17241 -11646
rect 17275 -11680 17309 -11646
rect 17343 -11680 17377 -11646
rect 17411 -11680 17445 -11646
rect 17479 -11680 17513 -11646
rect 17547 -11680 17581 -11646
rect 17615 -11663 17654 -11646
rect 18084 -11646 18672 -11630
rect 18084 -11663 18123 -11646
rect 17615 -11680 17840 -11663
rect 16880 -11718 17840 -11680
rect 17898 -11680 18123 -11663
rect 18157 -11680 18191 -11646
rect 18225 -11680 18259 -11646
rect 18293 -11680 18327 -11646
rect 18361 -11680 18395 -11646
rect 18429 -11680 18463 -11646
rect 18497 -11680 18531 -11646
rect 18565 -11680 18599 -11646
rect 18633 -11663 18672 -11646
rect 19102 -11646 19690 -11630
rect 19102 -11663 19141 -11646
rect 18633 -11680 18858 -11663
rect 17898 -11718 18858 -11680
rect 18916 -11680 19141 -11663
rect 19175 -11680 19209 -11646
rect 19243 -11680 19277 -11646
rect 19311 -11680 19345 -11646
rect 19379 -11680 19413 -11646
rect 19447 -11680 19481 -11646
rect 19515 -11680 19549 -11646
rect 19583 -11680 19617 -11646
rect 19651 -11663 19690 -11646
rect 20120 -11646 20708 -11630
rect 20120 -11663 20159 -11646
rect 19651 -11680 19876 -11663
rect 18916 -11718 19876 -11680
rect 19934 -11680 20159 -11663
rect 20193 -11680 20227 -11646
rect 20261 -11680 20295 -11646
rect 20329 -11680 20363 -11646
rect 20397 -11680 20431 -11646
rect 20465 -11680 20499 -11646
rect 20533 -11680 20567 -11646
rect 20601 -11680 20635 -11646
rect 20669 -11663 20708 -11646
rect 21138 -11646 21726 -11630
rect 21138 -11663 21177 -11646
rect 20669 -11680 20894 -11663
rect 19934 -11718 20894 -11680
rect 20952 -11680 21177 -11663
rect 21211 -11680 21245 -11646
rect 21279 -11680 21313 -11646
rect 21347 -11680 21381 -11646
rect 21415 -11680 21449 -11646
rect 21483 -11680 21517 -11646
rect 21551 -11680 21585 -11646
rect 21619 -11680 21653 -11646
rect 21687 -11663 21726 -11646
rect 22156 -11646 22744 -11630
rect 22156 -11663 22195 -11646
rect 21687 -11680 21912 -11663
rect 20952 -11718 21912 -11680
rect 21970 -11680 22195 -11663
rect 22229 -11680 22263 -11646
rect 22297 -11680 22331 -11646
rect 22365 -11680 22399 -11646
rect 22433 -11680 22467 -11646
rect 22501 -11680 22535 -11646
rect 22569 -11680 22603 -11646
rect 22637 -11680 22671 -11646
rect 22705 -11663 22744 -11646
rect 22705 -11680 22930 -11663
rect 21970 -11718 22930 -11680
rect 2628 -12356 3588 -12318
rect 2628 -12373 2853 -12356
rect 2814 -12390 2853 -12373
rect 2887 -12390 2921 -12356
rect 2955 -12390 2989 -12356
rect 3023 -12390 3057 -12356
rect 3091 -12390 3125 -12356
rect 3159 -12390 3193 -12356
rect 3227 -12390 3261 -12356
rect 3295 -12390 3329 -12356
rect 3363 -12373 3588 -12356
rect 3646 -12356 4606 -12318
rect 3646 -12373 3871 -12356
rect 3363 -12390 3402 -12373
rect 2814 -12406 3402 -12390
rect 3832 -12390 3871 -12373
rect 3905 -12390 3939 -12356
rect 3973 -12390 4007 -12356
rect 4041 -12390 4075 -12356
rect 4109 -12390 4143 -12356
rect 4177 -12390 4211 -12356
rect 4245 -12390 4279 -12356
rect 4313 -12390 4347 -12356
rect 4381 -12373 4606 -12356
rect 4664 -12356 5624 -12318
rect 4664 -12373 4889 -12356
rect 4381 -12390 4420 -12373
rect 3832 -12406 4420 -12390
rect 4850 -12390 4889 -12373
rect 4923 -12390 4957 -12356
rect 4991 -12390 5025 -12356
rect 5059 -12390 5093 -12356
rect 5127 -12390 5161 -12356
rect 5195 -12390 5229 -12356
rect 5263 -12390 5297 -12356
rect 5331 -12390 5365 -12356
rect 5399 -12373 5624 -12356
rect 5682 -12356 6642 -12318
rect 5682 -12373 5907 -12356
rect 5399 -12390 5438 -12373
rect 4850 -12406 5438 -12390
rect 5868 -12390 5907 -12373
rect 5941 -12390 5975 -12356
rect 6009 -12390 6043 -12356
rect 6077 -12390 6111 -12356
rect 6145 -12390 6179 -12356
rect 6213 -12390 6247 -12356
rect 6281 -12390 6315 -12356
rect 6349 -12390 6383 -12356
rect 6417 -12373 6642 -12356
rect 6700 -12356 7660 -12318
rect 6700 -12373 6925 -12356
rect 6417 -12390 6456 -12373
rect 5868 -12406 6456 -12390
rect 6886 -12390 6925 -12373
rect 6959 -12390 6993 -12356
rect 7027 -12390 7061 -12356
rect 7095 -12390 7129 -12356
rect 7163 -12390 7197 -12356
rect 7231 -12390 7265 -12356
rect 7299 -12390 7333 -12356
rect 7367 -12390 7401 -12356
rect 7435 -12373 7660 -12356
rect 7718 -12356 8678 -12318
rect 7718 -12373 7943 -12356
rect 7435 -12390 7474 -12373
rect 6886 -12406 7474 -12390
rect 7904 -12390 7943 -12373
rect 7977 -12390 8011 -12356
rect 8045 -12390 8079 -12356
rect 8113 -12390 8147 -12356
rect 8181 -12390 8215 -12356
rect 8249 -12390 8283 -12356
rect 8317 -12390 8351 -12356
rect 8385 -12390 8419 -12356
rect 8453 -12373 8678 -12356
rect 8736 -12356 9696 -12318
rect 8736 -12373 8961 -12356
rect 8453 -12390 8492 -12373
rect 7904 -12406 8492 -12390
rect 8922 -12390 8961 -12373
rect 8995 -12390 9029 -12356
rect 9063 -12390 9097 -12356
rect 9131 -12390 9165 -12356
rect 9199 -12390 9233 -12356
rect 9267 -12390 9301 -12356
rect 9335 -12390 9369 -12356
rect 9403 -12390 9437 -12356
rect 9471 -12373 9696 -12356
rect 9754 -12356 10714 -12318
rect 9754 -12373 9979 -12356
rect 9471 -12390 9510 -12373
rect 8922 -12406 9510 -12390
rect 9940 -12390 9979 -12373
rect 10013 -12390 10047 -12356
rect 10081 -12390 10115 -12356
rect 10149 -12390 10183 -12356
rect 10217 -12390 10251 -12356
rect 10285 -12390 10319 -12356
rect 10353 -12390 10387 -12356
rect 10421 -12390 10455 -12356
rect 10489 -12373 10714 -12356
rect 10772 -12356 11732 -12318
rect 10772 -12373 10997 -12356
rect 10489 -12390 10528 -12373
rect 9940 -12406 10528 -12390
rect 10958 -12390 10997 -12373
rect 11031 -12390 11065 -12356
rect 11099 -12390 11133 -12356
rect 11167 -12390 11201 -12356
rect 11235 -12390 11269 -12356
rect 11303 -12390 11337 -12356
rect 11371 -12390 11405 -12356
rect 11439 -12390 11473 -12356
rect 11507 -12373 11732 -12356
rect 11790 -12356 12750 -12318
rect 11790 -12373 12015 -12356
rect 11507 -12390 11546 -12373
rect 10958 -12406 11546 -12390
rect 11976 -12390 12015 -12373
rect 12049 -12390 12083 -12356
rect 12117 -12390 12151 -12356
rect 12185 -12390 12219 -12356
rect 12253 -12390 12287 -12356
rect 12321 -12390 12355 -12356
rect 12389 -12390 12423 -12356
rect 12457 -12390 12491 -12356
rect 12525 -12373 12750 -12356
rect 12808 -12356 13768 -12318
rect 12808 -12373 13033 -12356
rect 12525 -12390 12564 -12373
rect 11976 -12406 12564 -12390
rect 12994 -12390 13033 -12373
rect 13067 -12390 13101 -12356
rect 13135 -12390 13169 -12356
rect 13203 -12390 13237 -12356
rect 13271 -12390 13305 -12356
rect 13339 -12390 13373 -12356
rect 13407 -12390 13441 -12356
rect 13475 -12390 13509 -12356
rect 13543 -12373 13768 -12356
rect 13826 -12356 14786 -12318
rect 13826 -12373 14051 -12356
rect 13543 -12390 13582 -12373
rect 12994 -12406 13582 -12390
rect 14012 -12390 14051 -12373
rect 14085 -12390 14119 -12356
rect 14153 -12390 14187 -12356
rect 14221 -12390 14255 -12356
rect 14289 -12390 14323 -12356
rect 14357 -12390 14391 -12356
rect 14425 -12390 14459 -12356
rect 14493 -12390 14527 -12356
rect 14561 -12373 14786 -12356
rect 14844 -12356 15804 -12318
rect 14844 -12373 15069 -12356
rect 14561 -12390 14600 -12373
rect 14012 -12406 14600 -12390
rect 15030 -12390 15069 -12373
rect 15103 -12390 15137 -12356
rect 15171 -12390 15205 -12356
rect 15239 -12390 15273 -12356
rect 15307 -12390 15341 -12356
rect 15375 -12390 15409 -12356
rect 15443 -12390 15477 -12356
rect 15511 -12390 15545 -12356
rect 15579 -12373 15804 -12356
rect 15862 -12356 16822 -12318
rect 15862 -12373 16087 -12356
rect 15579 -12390 15618 -12373
rect 15030 -12406 15618 -12390
rect 16048 -12390 16087 -12373
rect 16121 -12390 16155 -12356
rect 16189 -12390 16223 -12356
rect 16257 -12390 16291 -12356
rect 16325 -12390 16359 -12356
rect 16393 -12390 16427 -12356
rect 16461 -12390 16495 -12356
rect 16529 -12390 16563 -12356
rect 16597 -12373 16822 -12356
rect 16880 -12356 17840 -12318
rect 16880 -12373 17105 -12356
rect 16597 -12390 16636 -12373
rect 16048 -12406 16636 -12390
rect 17066 -12390 17105 -12373
rect 17139 -12390 17173 -12356
rect 17207 -12390 17241 -12356
rect 17275 -12390 17309 -12356
rect 17343 -12390 17377 -12356
rect 17411 -12390 17445 -12356
rect 17479 -12390 17513 -12356
rect 17547 -12390 17581 -12356
rect 17615 -12373 17840 -12356
rect 17898 -12356 18858 -12318
rect 17898 -12373 18123 -12356
rect 17615 -12390 17654 -12373
rect 17066 -12406 17654 -12390
rect 18084 -12390 18123 -12373
rect 18157 -12390 18191 -12356
rect 18225 -12390 18259 -12356
rect 18293 -12390 18327 -12356
rect 18361 -12390 18395 -12356
rect 18429 -12390 18463 -12356
rect 18497 -12390 18531 -12356
rect 18565 -12390 18599 -12356
rect 18633 -12373 18858 -12356
rect 18916 -12356 19876 -12318
rect 18916 -12373 19141 -12356
rect 18633 -12390 18672 -12373
rect 18084 -12406 18672 -12390
rect 19102 -12390 19141 -12373
rect 19175 -12390 19209 -12356
rect 19243 -12390 19277 -12356
rect 19311 -12390 19345 -12356
rect 19379 -12390 19413 -12356
rect 19447 -12390 19481 -12356
rect 19515 -12390 19549 -12356
rect 19583 -12390 19617 -12356
rect 19651 -12373 19876 -12356
rect 19934 -12356 20894 -12318
rect 19934 -12373 20159 -12356
rect 19651 -12390 19690 -12373
rect 19102 -12406 19690 -12390
rect 20120 -12390 20159 -12373
rect 20193 -12390 20227 -12356
rect 20261 -12390 20295 -12356
rect 20329 -12390 20363 -12356
rect 20397 -12390 20431 -12356
rect 20465 -12390 20499 -12356
rect 20533 -12390 20567 -12356
rect 20601 -12390 20635 -12356
rect 20669 -12373 20894 -12356
rect 20952 -12356 21912 -12318
rect 20952 -12373 21177 -12356
rect 20669 -12390 20708 -12373
rect 20120 -12406 20708 -12390
rect 21138 -12390 21177 -12373
rect 21211 -12390 21245 -12356
rect 21279 -12390 21313 -12356
rect 21347 -12390 21381 -12356
rect 21415 -12390 21449 -12356
rect 21483 -12390 21517 -12356
rect 21551 -12390 21585 -12356
rect 21619 -12390 21653 -12356
rect 21687 -12373 21912 -12356
rect 21970 -12356 22930 -12318
rect 21970 -12373 22195 -12356
rect 21687 -12390 21726 -12373
rect 21138 -12406 21726 -12390
rect 22156 -12390 22195 -12373
rect 22229 -12390 22263 -12356
rect 22297 -12390 22331 -12356
rect 22365 -12390 22399 -12356
rect 22433 -12390 22467 -12356
rect 22501 -12390 22535 -12356
rect 22569 -12390 22603 -12356
rect 22637 -12390 22671 -12356
rect 22705 -12373 22930 -12356
rect 22705 -12390 22744 -12373
rect 22156 -12406 22744 -12390
rect -8952 -12440 -8364 -12424
rect -8952 -12457 -8913 -12440
rect -9138 -12474 -8913 -12457
rect -8879 -12474 -8845 -12440
rect -8811 -12474 -8777 -12440
rect -8743 -12474 -8709 -12440
rect -8675 -12474 -8641 -12440
rect -8607 -12474 -8573 -12440
rect -8539 -12474 -8505 -12440
rect -8471 -12474 -8437 -12440
rect -8403 -12457 -8364 -12440
rect -7934 -12440 -7346 -12424
rect -7934 -12457 -7895 -12440
rect -8403 -12474 -8178 -12457
rect -9138 -12512 -8178 -12474
rect -8120 -12474 -7895 -12457
rect -7861 -12474 -7827 -12440
rect -7793 -12474 -7759 -12440
rect -7725 -12474 -7691 -12440
rect -7657 -12474 -7623 -12440
rect -7589 -12474 -7555 -12440
rect -7521 -12474 -7487 -12440
rect -7453 -12474 -7419 -12440
rect -7385 -12457 -7346 -12440
rect -6916 -12440 -6328 -12424
rect -6916 -12457 -6877 -12440
rect -7385 -12474 -7160 -12457
rect -8120 -12512 -7160 -12474
rect -7102 -12474 -6877 -12457
rect -6843 -12474 -6809 -12440
rect -6775 -12474 -6741 -12440
rect -6707 -12474 -6673 -12440
rect -6639 -12474 -6605 -12440
rect -6571 -12474 -6537 -12440
rect -6503 -12474 -6469 -12440
rect -6435 -12474 -6401 -12440
rect -6367 -12457 -6328 -12440
rect -5898 -12440 -5310 -12424
rect -5898 -12457 -5859 -12440
rect -6367 -12474 -6142 -12457
rect -7102 -12512 -6142 -12474
rect -6084 -12474 -5859 -12457
rect -5825 -12474 -5791 -12440
rect -5757 -12474 -5723 -12440
rect -5689 -12474 -5655 -12440
rect -5621 -12474 -5587 -12440
rect -5553 -12474 -5519 -12440
rect -5485 -12474 -5451 -12440
rect -5417 -12474 -5383 -12440
rect -5349 -12457 -5310 -12440
rect -4880 -12440 -4292 -12424
rect -4880 -12457 -4841 -12440
rect -5349 -12474 -5124 -12457
rect -6084 -12512 -5124 -12474
rect -5066 -12474 -4841 -12457
rect -4807 -12474 -4773 -12440
rect -4739 -12474 -4705 -12440
rect -4671 -12474 -4637 -12440
rect -4603 -12474 -4569 -12440
rect -4535 -12474 -4501 -12440
rect -4467 -12474 -4433 -12440
rect -4399 -12474 -4365 -12440
rect -4331 -12457 -4292 -12440
rect -3862 -12440 -3274 -12424
rect -3862 -12457 -3823 -12440
rect -4331 -12474 -4106 -12457
rect -5066 -12512 -4106 -12474
rect -4048 -12474 -3823 -12457
rect -3789 -12474 -3755 -12440
rect -3721 -12474 -3687 -12440
rect -3653 -12474 -3619 -12440
rect -3585 -12474 -3551 -12440
rect -3517 -12474 -3483 -12440
rect -3449 -12474 -3415 -12440
rect -3381 -12474 -3347 -12440
rect -3313 -12457 -3274 -12440
rect -2844 -12440 -2256 -12424
rect -2844 -12457 -2805 -12440
rect -3313 -12474 -3088 -12457
rect -4048 -12512 -3088 -12474
rect -3030 -12474 -2805 -12457
rect -2771 -12474 -2737 -12440
rect -2703 -12474 -2669 -12440
rect -2635 -12474 -2601 -12440
rect -2567 -12474 -2533 -12440
rect -2499 -12474 -2465 -12440
rect -2431 -12474 -2397 -12440
rect -2363 -12474 -2329 -12440
rect -2295 -12457 -2256 -12440
rect -1826 -12440 -1238 -12424
rect -1826 -12457 -1787 -12440
rect -2295 -12474 -2070 -12457
rect -3030 -12512 -2070 -12474
rect -2012 -12474 -1787 -12457
rect -1753 -12474 -1719 -12440
rect -1685 -12474 -1651 -12440
rect -1617 -12474 -1583 -12440
rect -1549 -12474 -1515 -12440
rect -1481 -12474 -1447 -12440
rect -1413 -12474 -1379 -12440
rect -1345 -12474 -1311 -12440
rect -1277 -12457 -1238 -12440
rect -808 -12440 -220 -12424
rect -808 -12457 -769 -12440
rect -1277 -12474 -1052 -12457
rect -2012 -12512 -1052 -12474
rect -994 -12474 -769 -12457
rect -735 -12474 -701 -12440
rect -667 -12474 -633 -12440
rect -599 -12474 -565 -12440
rect -531 -12474 -497 -12440
rect -463 -12474 -429 -12440
rect -395 -12474 -361 -12440
rect -327 -12474 -293 -12440
rect -259 -12457 -220 -12440
rect -259 -12474 -34 -12457
rect -994 -12512 -34 -12474
rect 2814 -12880 3402 -12864
rect 2814 -12897 2853 -12880
rect 2628 -12914 2853 -12897
rect 2887 -12914 2921 -12880
rect 2955 -12914 2989 -12880
rect 3023 -12914 3057 -12880
rect 3091 -12914 3125 -12880
rect 3159 -12914 3193 -12880
rect 3227 -12914 3261 -12880
rect 3295 -12914 3329 -12880
rect 3363 -12897 3402 -12880
rect 3832 -12880 4420 -12864
rect 3832 -12897 3871 -12880
rect 3363 -12914 3588 -12897
rect 2628 -12952 3588 -12914
rect 3646 -12914 3871 -12897
rect 3905 -12914 3939 -12880
rect 3973 -12914 4007 -12880
rect 4041 -12914 4075 -12880
rect 4109 -12914 4143 -12880
rect 4177 -12914 4211 -12880
rect 4245 -12914 4279 -12880
rect 4313 -12914 4347 -12880
rect 4381 -12897 4420 -12880
rect 4850 -12880 5438 -12864
rect 4850 -12897 4889 -12880
rect 4381 -12914 4606 -12897
rect 3646 -12952 4606 -12914
rect 4664 -12914 4889 -12897
rect 4923 -12914 4957 -12880
rect 4991 -12914 5025 -12880
rect 5059 -12914 5093 -12880
rect 5127 -12914 5161 -12880
rect 5195 -12914 5229 -12880
rect 5263 -12914 5297 -12880
rect 5331 -12914 5365 -12880
rect 5399 -12897 5438 -12880
rect 5868 -12880 6456 -12864
rect 5868 -12897 5907 -12880
rect 5399 -12914 5624 -12897
rect 4664 -12952 5624 -12914
rect 5682 -12914 5907 -12897
rect 5941 -12914 5975 -12880
rect 6009 -12914 6043 -12880
rect 6077 -12914 6111 -12880
rect 6145 -12914 6179 -12880
rect 6213 -12914 6247 -12880
rect 6281 -12914 6315 -12880
rect 6349 -12914 6383 -12880
rect 6417 -12897 6456 -12880
rect 6886 -12880 7474 -12864
rect 6886 -12897 6925 -12880
rect 6417 -12914 6642 -12897
rect 5682 -12952 6642 -12914
rect 6700 -12914 6925 -12897
rect 6959 -12914 6993 -12880
rect 7027 -12914 7061 -12880
rect 7095 -12914 7129 -12880
rect 7163 -12914 7197 -12880
rect 7231 -12914 7265 -12880
rect 7299 -12914 7333 -12880
rect 7367 -12914 7401 -12880
rect 7435 -12897 7474 -12880
rect 7904 -12880 8492 -12864
rect 7904 -12897 7943 -12880
rect 7435 -12914 7660 -12897
rect 6700 -12952 7660 -12914
rect 7718 -12914 7943 -12897
rect 7977 -12914 8011 -12880
rect 8045 -12914 8079 -12880
rect 8113 -12914 8147 -12880
rect 8181 -12914 8215 -12880
rect 8249 -12914 8283 -12880
rect 8317 -12914 8351 -12880
rect 8385 -12914 8419 -12880
rect 8453 -12897 8492 -12880
rect 8922 -12880 9510 -12864
rect 8922 -12897 8961 -12880
rect 8453 -12914 8678 -12897
rect 7718 -12952 8678 -12914
rect 8736 -12914 8961 -12897
rect 8995 -12914 9029 -12880
rect 9063 -12914 9097 -12880
rect 9131 -12914 9165 -12880
rect 9199 -12914 9233 -12880
rect 9267 -12914 9301 -12880
rect 9335 -12914 9369 -12880
rect 9403 -12914 9437 -12880
rect 9471 -12897 9510 -12880
rect 9940 -12880 10528 -12864
rect 9940 -12897 9979 -12880
rect 9471 -12914 9696 -12897
rect 8736 -12952 9696 -12914
rect 9754 -12914 9979 -12897
rect 10013 -12914 10047 -12880
rect 10081 -12914 10115 -12880
rect 10149 -12914 10183 -12880
rect 10217 -12914 10251 -12880
rect 10285 -12914 10319 -12880
rect 10353 -12914 10387 -12880
rect 10421 -12914 10455 -12880
rect 10489 -12897 10528 -12880
rect 10958 -12880 11546 -12864
rect 10958 -12897 10997 -12880
rect 10489 -12914 10714 -12897
rect 9754 -12952 10714 -12914
rect 10772 -12914 10997 -12897
rect 11031 -12914 11065 -12880
rect 11099 -12914 11133 -12880
rect 11167 -12914 11201 -12880
rect 11235 -12914 11269 -12880
rect 11303 -12914 11337 -12880
rect 11371 -12914 11405 -12880
rect 11439 -12914 11473 -12880
rect 11507 -12897 11546 -12880
rect 11976 -12880 12564 -12864
rect 11976 -12897 12015 -12880
rect 11507 -12914 11732 -12897
rect 10772 -12952 11732 -12914
rect 11790 -12914 12015 -12897
rect 12049 -12914 12083 -12880
rect 12117 -12914 12151 -12880
rect 12185 -12914 12219 -12880
rect 12253 -12914 12287 -12880
rect 12321 -12914 12355 -12880
rect 12389 -12914 12423 -12880
rect 12457 -12914 12491 -12880
rect 12525 -12897 12564 -12880
rect 12994 -12880 13582 -12864
rect 12994 -12897 13033 -12880
rect 12525 -12914 12750 -12897
rect 11790 -12952 12750 -12914
rect 12808 -12914 13033 -12897
rect 13067 -12914 13101 -12880
rect 13135 -12914 13169 -12880
rect 13203 -12914 13237 -12880
rect 13271 -12914 13305 -12880
rect 13339 -12914 13373 -12880
rect 13407 -12914 13441 -12880
rect 13475 -12914 13509 -12880
rect 13543 -12897 13582 -12880
rect 14012 -12880 14600 -12864
rect 14012 -12897 14051 -12880
rect 13543 -12914 13768 -12897
rect 12808 -12952 13768 -12914
rect 13826 -12914 14051 -12897
rect 14085 -12914 14119 -12880
rect 14153 -12914 14187 -12880
rect 14221 -12914 14255 -12880
rect 14289 -12914 14323 -12880
rect 14357 -12914 14391 -12880
rect 14425 -12914 14459 -12880
rect 14493 -12914 14527 -12880
rect 14561 -12897 14600 -12880
rect 15030 -12880 15618 -12864
rect 15030 -12897 15069 -12880
rect 14561 -12914 14786 -12897
rect 13826 -12952 14786 -12914
rect 14844 -12914 15069 -12897
rect 15103 -12914 15137 -12880
rect 15171 -12914 15205 -12880
rect 15239 -12914 15273 -12880
rect 15307 -12914 15341 -12880
rect 15375 -12914 15409 -12880
rect 15443 -12914 15477 -12880
rect 15511 -12914 15545 -12880
rect 15579 -12897 15618 -12880
rect 16048 -12880 16636 -12864
rect 16048 -12897 16087 -12880
rect 15579 -12914 15804 -12897
rect 14844 -12952 15804 -12914
rect 15862 -12914 16087 -12897
rect 16121 -12914 16155 -12880
rect 16189 -12914 16223 -12880
rect 16257 -12914 16291 -12880
rect 16325 -12914 16359 -12880
rect 16393 -12914 16427 -12880
rect 16461 -12914 16495 -12880
rect 16529 -12914 16563 -12880
rect 16597 -12897 16636 -12880
rect 17066 -12880 17654 -12864
rect 17066 -12897 17105 -12880
rect 16597 -12914 16822 -12897
rect 15862 -12952 16822 -12914
rect 16880 -12914 17105 -12897
rect 17139 -12914 17173 -12880
rect 17207 -12914 17241 -12880
rect 17275 -12914 17309 -12880
rect 17343 -12914 17377 -12880
rect 17411 -12914 17445 -12880
rect 17479 -12914 17513 -12880
rect 17547 -12914 17581 -12880
rect 17615 -12897 17654 -12880
rect 18084 -12880 18672 -12864
rect 18084 -12897 18123 -12880
rect 17615 -12914 17840 -12897
rect 16880 -12952 17840 -12914
rect 17898 -12914 18123 -12897
rect 18157 -12914 18191 -12880
rect 18225 -12914 18259 -12880
rect 18293 -12914 18327 -12880
rect 18361 -12914 18395 -12880
rect 18429 -12914 18463 -12880
rect 18497 -12914 18531 -12880
rect 18565 -12914 18599 -12880
rect 18633 -12897 18672 -12880
rect 19102 -12880 19690 -12864
rect 19102 -12897 19141 -12880
rect 18633 -12914 18858 -12897
rect 17898 -12952 18858 -12914
rect 18916 -12914 19141 -12897
rect 19175 -12914 19209 -12880
rect 19243 -12914 19277 -12880
rect 19311 -12914 19345 -12880
rect 19379 -12914 19413 -12880
rect 19447 -12914 19481 -12880
rect 19515 -12914 19549 -12880
rect 19583 -12914 19617 -12880
rect 19651 -12897 19690 -12880
rect 20120 -12880 20708 -12864
rect 20120 -12897 20159 -12880
rect 19651 -12914 19876 -12897
rect 18916 -12952 19876 -12914
rect 19934 -12914 20159 -12897
rect 20193 -12914 20227 -12880
rect 20261 -12914 20295 -12880
rect 20329 -12914 20363 -12880
rect 20397 -12914 20431 -12880
rect 20465 -12914 20499 -12880
rect 20533 -12914 20567 -12880
rect 20601 -12914 20635 -12880
rect 20669 -12897 20708 -12880
rect 21138 -12880 21726 -12864
rect 21138 -12897 21177 -12880
rect 20669 -12914 20894 -12897
rect 19934 -12952 20894 -12914
rect 20952 -12914 21177 -12897
rect 21211 -12914 21245 -12880
rect 21279 -12914 21313 -12880
rect 21347 -12914 21381 -12880
rect 21415 -12914 21449 -12880
rect 21483 -12914 21517 -12880
rect 21551 -12914 21585 -12880
rect 21619 -12914 21653 -12880
rect 21687 -12897 21726 -12880
rect 22156 -12880 22744 -12864
rect 22156 -12897 22195 -12880
rect 21687 -12914 21912 -12897
rect 20952 -12952 21912 -12914
rect 21970 -12914 22195 -12897
rect 22229 -12914 22263 -12880
rect 22297 -12914 22331 -12880
rect 22365 -12914 22399 -12880
rect 22433 -12914 22467 -12880
rect 22501 -12914 22535 -12880
rect 22569 -12914 22603 -12880
rect 22637 -12914 22671 -12880
rect 22705 -12897 22744 -12880
rect 22705 -12914 22930 -12897
rect 21970 -12952 22930 -12914
rect -9138 -13150 -8178 -13112
rect -9138 -13167 -8913 -13150
rect -8952 -13184 -8913 -13167
rect -8879 -13184 -8845 -13150
rect -8811 -13184 -8777 -13150
rect -8743 -13184 -8709 -13150
rect -8675 -13184 -8641 -13150
rect -8607 -13184 -8573 -13150
rect -8539 -13184 -8505 -13150
rect -8471 -13184 -8437 -13150
rect -8403 -13167 -8178 -13150
rect -8120 -13150 -7160 -13112
rect -8120 -13167 -7895 -13150
rect -8403 -13184 -8364 -13167
rect -8952 -13200 -8364 -13184
rect -7934 -13184 -7895 -13167
rect -7861 -13184 -7827 -13150
rect -7793 -13184 -7759 -13150
rect -7725 -13184 -7691 -13150
rect -7657 -13184 -7623 -13150
rect -7589 -13184 -7555 -13150
rect -7521 -13184 -7487 -13150
rect -7453 -13184 -7419 -13150
rect -7385 -13167 -7160 -13150
rect -7102 -13150 -6142 -13112
rect -7102 -13167 -6877 -13150
rect -7385 -13184 -7346 -13167
rect -7934 -13200 -7346 -13184
rect -6916 -13184 -6877 -13167
rect -6843 -13184 -6809 -13150
rect -6775 -13184 -6741 -13150
rect -6707 -13184 -6673 -13150
rect -6639 -13184 -6605 -13150
rect -6571 -13184 -6537 -13150
rect -6503 -13184 -6469 -13150
rect -6435 -13184 -6401 -13150
rect -6367 -13167 -6142 -13150
rect -6084 -13150 -5124 -13112
rect -6084 -13167 -5859 -13150
rect -6367 -13184 -6328 -13167
rect -6916 -13200 -6328 -13184
rect -5898 -13184 -5859 -13167
rect -5825 -13184 -5791 -13150
rect -5757 -13184 -5723 -13150
rect -5689 -13184 -5655 -13150
rect -5621 -13184 -5587 -13150
rect -5553 -13184 -5519 -13150
rect -5485 -13184 -5451 -13150
rect -5417 -13184 -5383 -13150
rect -5349 -13167 -5124 -13150
rect -5066 -13150 -4106 -13112
rect -5066 -13167 -4841 -13150
rect -5349 -13184 -5310 -13167
rect -5898 -13200 -5310 -13184
rect -4880 -13184 -4841 -13167
rect -4807 -13184 -4773 -13150
rect -4739 -13184 -4705 -13150
rect -4671 -13184 -4637 -13150
rect -4603 -13184 -4569 -13150
rect -4535 -13184 -4501 -13150
rect -4467 -13184 -4433 -13150
rect -4399 -13184 -4365 -13150
rect -4331 -13167 -4106 -13150
rect -4048 -13150 -3088 -13112
rect -4048 -13167 -3823 -13150
rect -4331 -13184 -4292 -13167
rect -4880 -13200 -4292 -13184
rect -3862 -13184 -3823 -13167
rect -3789 -13184 -3755 -13150
rect -3721 -13184 -3687 -13150
rect -3653 -13184 -3619 -13150
rect -3585 -13184 -3551 -13150
rect -3517 -13184 -3483 -13150
rect -3449 -13184 -3415 -13150
rect -3381 -13184 -3347 -13150
rect -3313 -13167 -3088 -13150
rect -3030 -13150 -2070 -13112
rect -3030 -13167 -2805 -13150
rect -3313 -13184 -3274 -13167
rect -3862 -13200 -3274 -13184
rect -2844 -13184 -2805 -13167
rect -2771 -13184 -2737 -13150
rect -2703 -13184 -2669 -13150
rect -2635 -13184 -2601 -13150
rect -2567 -13184 -2533 -13150
rect -2499 -13184 -2465 -13150
rect -2431 -13184 -2397 -13150
rect -2363 -13184 -2329 -13150
rect -2295 -13167 -2070 -13150
rect -2012 -13150 -1052 -13112
rect -2012 -13167 -1787 -13150
rect -2295 -13184 -2256 -13167
rect -2844 -13200 -2256 -13184
rect -1826 -13184 -1787 -13167
rect -1753 -13184 -1719 -13150
rect -1685 -13184 -1651 -13150
rect -1617 -13184 -1583 -13150
rect -1549 -13184 -1515 -13150
rect -1481 -13184 -1447 -13150
rect -1413 -13184 -1379 -13150
rect -1345 -13184 -1311 -13150
rect -1277 -13167 -1052 -13150
rect -994 -13150 -34 -13112
rect -994 -13167 -769 -13150
rect -1277 -13184 -1238 -13167
rect -1826 -13200 -1238 -13184
rect -808 -13184 -769 -13167
rect -735 -13184 -701 -13150
rect -667 -13184 -633 -13150
rect -599 -13184 -565 -13150
rect -531 -13184 -497 -13150
rect -463 -13184 -429 -13150
rect -395 -13184 -361 -13150
rect -327 -13184 -293 -13150
rect -259 -13167 -34 -13150
rect -259 -13184 -220 -13167
rect -808 -13200 -220 -13184
rect -8952 -13258 -8364 -13242
rect -8952 -13275 -8913 -13258
rect -9138 -13292 -8913 -13275
rect -8879 -13292 -8845 -13258
rect -8811 -13292 -8777 -13258
rect -8743 -13292 -8709 -13258
rect -8675 -13292 -8641 -13258
rect -8607 -13292 -8573 -13258
rect -8539 -13292 -8505 -13258
rect -8471 -13292 -8437 -13258
rect -8403 -13275 -8364 -13258
rect -7934 -13258 -7346 -13242
rect -7934 -13275 -7895 -13258
rect -8403 -13292 -8178 -13275
rect -9138 -13330 -8178 -13292
rect -8120 -13292 -7895 -13275
rect -7861 -13292 -7827 -13258
rect -7793 -13292 -7759 -13258
rect -7725 -13292 -7691 -13258
rect -7657 -13292 -7623 -13258
rect -7589 -13292 -7555 -13258
rect -7521 -13292 -7487 -13258
rect -7453 -13292 -7419 -13258
rect -7385 -13275 -7346 -13258
rect -6916 -13258 -6328 -13242
rect -6916 -13275 -6877 -13258
rect -7385 -13292 -7160 -13275
rect -8120 -13330 -7160 -13292
rect -7102 -13292 -6877 -13275
rect -6843 -13292 -6809 -13258
rect -6775 -13292 -6741 -13258
rect -6707 -13292 -6673 -13258
rect -6639 -13292 -6605 -13258
rect -6571 -13292 -6537 -13258
rect -6503 -13292 -6469 -13258
rect -6435 -13292 -6401 -13258
rect -6367 -13275 -6328 -13258
rect -5898 -13258 -5310 -13242
rect -5898 -13275 -5859 -13258
rect -6367 -13292 -6142 -13275
rect -7102 -13330 -6142 -13292
rect -6084 -13292 -5859 -13275
rect -5825 -13292 -5791 -13258
rect -5757 -13292 -5723 -13258
rect -5689 -13292 -5655 -13258
rect -5621 -13292 -5587 -13258
rect -5553 -13292 -5519 -13258
rect -5485 -13292 -5451 -13258
rect -5417 -13292 -5383 -13258
rect -5349 -13275 -5310 -13258
rect -4880 -13258 -4292 -13242
rect -4880 -13275 -4841 -13258
rect -5349 -13292 -5124 -13275
rect -6084 -13330 -5124 -13292
rect -5066 -13292 -4841 -13275
rect -4807 -13292 -4773 -13258
rect -4739 -13292 -4705 -13258
rect -4671 -13292 -4637 -13258
rect -4603 -13292 -4569 -13258
rect -4535 -13292 -4501 -13258
rect -4467 -13292 -4433 -13258
rect -4399 -13292 -4365 -13258
rect -4331 -13275 -4292 -13258
rect -3862 -13258 -3274 -13242
rect -3862 -13275 -3823 -13258
rect -4331 -13292 -4106 -13275
rect -5066 -13330 -4106 -13292
rect -4048 -13292 -3823 -13275
rect -3789 -13292 -3755 -13258
rect -3721 -13292 -3687 -13258
rect -3653 -13292 -3619 -13258
rect -3585 -13292 -3551 -13258
rect -3517 -13292 -3483 -13258
rect -3449 -13292 -3415 -13258
rect -3381 -13292 -3347 -13258
rect -3313 -13275 -3274 -13258
rect -2844 -13258 -2256 -13242
rect -2844 -13275 -2805 -13258
rect -3313 -13292 -3088 -13275
rect -4048 -13330 -3088 -13292
rect -3030 -13292 -2805 -13275
rect -2771 -13292 -2737 -13258
rect -2703 -13292 -2669 -13258
rect -2635 -13292 -2601 -13258
rect -2567 -13292 -2533 -13258
rect -2499 -13292 -2465 -13258
rect -2431 -13292 -2397 -13258
rect -2363 -13292 -2329 -13258
rect -2295 -13275 -2256 -13258
rect -1826 -13258 -1238 -13242
rect -1826 -13275 -1787 -13258
rect -2295 -13292 -2070 -13275
rect -3030 -13330 -2070 -13292
rect -2012 -13292 -1787 -13275
rect -1753 -13292 -1719 -13258
rect -1685 -13292 -1651 -13258
rect -1617 -13292 -1583 -13258
rect -1549 -13292 -1515 -13258
rect -1481 -13292 -1447 -13258
rect -1413 -13292 -1379 -13258
rect -1345 -13292 -1311 -13258
rect -1277 -13275 -1238 -13258
rect -808 -13258 -220 -13242
rect -808 -13275 -769 -13258
rect -1277 -13292 -1052 -13275
rect -2012 -13330 -1052 -13292
rect -994 -13292 -769 -13275
rect -735 -13292 -701 -13258
rect -667 -13292 -633 -13258
rect -599 -13292 -565 -13258
rect -531 -13292 -497 -13258
rect -463 -13292 -429 -13258
rect -395 -13292 -361 -13258
rect -327 -13292 -293 -13258
rect -259 -13275 -220 -13258
rect -259 -13292 -34 -13275
rect -994 -13330 -34 -13292
rect 2628 -13590 3588 -13552
rect 2628 -13607 2853 -13590
rect 2814 -13624 2853 -13607
rect 2887 -13624 2921 -13590
rect 2955 -13624 2989 -13590
rect 3023 -13624 3057 -13590
rect 3091 -13624 3125 -13590
rect 3159 -13624 3193 -13590
rect 3227 -13624 3261 -13590
rect 3295 -13624 3329 -13590
rect 3363 -13607 3588 -13590
rect 3646 -13590 4606 -13552
rect 3646 -13607 3871 -13590
rect 3363 -13624 3402 -13607
rect 2814 -13640 3402 -13624
rect 3832 -13624 3871 -13607
rect 3905 -13624 3939 -13590
rect 3973 -13624 4007 -13590
rect 4041 -13624 4075 -13590
rect 4109 -13624 4143 -13590
rect 4177 -13624 4211 -13590
rect 4245 -13624 4279 -13590
rect 4313 -13624 4347 -13590
rect 4381 -13607 4606 -13590
rect 4664 -13590 5624 -13552
rect 4664 -13607 4889 -13590
rect 4381 -13624 4420 -13607
rect 3832 -13640 4420 -13624
rect 4850 -13624 4889 -13607
rect 4923 -13624 4957 -13590
rect 4991 -13624 5025 -13590
rect 5059 -13624 5093 -13590
rect 5127 -13624 5161 -13590
rect 5195 -13624 5229 -13590
rect 5263 -13624 5297 -13590
rect 5331 -13624 5365 -13590
rect 5399 -13607 5624 -13590
rect 5682 -13590 6642 -13552
rect 5682 -13607 5907 -13590
rect 5399 -13624 5438 -13607
rect 4850 -13640 5438 -13624
rect 5868 -13624 5907 -13607
rect 5941 -13624 5975 -13590
rect 6009 -13624 6043 -13590
rect 6077 -13624 6111 -13590
rect 6145 -13624 6179 -13590
rect 6213 -13624 6247 -13590
rect 6281 -13624 6315 -13590
rect 6349 -13624 6383 -13590
rect 6417 -13607 6642 -13590
rect 6700 -13590 7660 -13552
rect 6700 -13607 6925 -13590
rect 6417 -13624 6456 -13607
rect 5868 -13640 6456 -13624
rect 6886 -13624 6925 -13607
rect 6959 -13624 6993 -13590
rect 7027 -13624 7061 -13590
rect 7095 -13624 7129 -13590
rect 7163 -13624 7197 -13590
rect 7231 -13624 7265 -13590
rect 7299 -13624 7333 -13590
rect 7367 -13624 7401 -13590
rect 7435 -13607 7660 -13590
rect 7718 -13590 8678 -13552
rect 7718 -13607 7943 -13590
rect 7435 -13624 7474 -13607
rect 6886 -13640 7474 -13624
rect 7904 -13624 7943 -13607
rect 7977 -13624 8011 -13590
rect 8045 -13624 8079 -13590
rect 8113 -13624 8147 -13590
rect 8181 -13624 8215 -13590
rect 8249 -13624 8283 -13590
rect 8317 -13624 8351 -13590
rect 8385 -13624 8419 -13590
rect 8453 -13607 8678 -13590
rect 8736 -13590 9696 -13552
rect 8736 -13607 8961 -13590
rect 8453 -13624 8492 -13607
rect 7904 -13640 8492 -13624
rect 8922 -13624 8961 -13607
rect 8995 -13624 9029 -13590
rect 9063 -13624 9097 -13590
rect 9131 -13624 9165 -13590
rect 9199 -13624 9233 -13590
rect 9267 -13624 9301 -13590
rect 9335 -13624 9369 -13590
rect 9403 -13624 9437 -13590
rect 9471 -13607 9696 -13590
rect 9754 -13590 10714 -13552
rect 9754 -13607 9979 -13590
rect 9471 -13624 9510 -13607
rect 8922 -13640 9510 -13624
rect 9940 -13624 9979 -13607
rect 10013 -13624 10047 -13590
rect 10081 -13624 10115 -13590
rect 10149 -13624 10183 -13590
rect 10217 -13624 10251 -13590
rect 10285 -13624 10319 -13590
rect 10353 -13624 10387 -13590
rect 10421 -13624 10455 -13590
rect 10489 -13607 10714 -13590
rect 10772 -13590 11732 -13552
rect 10772 -13607 10997 -13590
rect 10489 -13624 10528 -13607
rect 9940 -13640 10528 -13624
rect 10958 -13624 10997 -13607
rect 11031 -13624 11065 -13590
rect 11099 -13624 11133 -13590
rect 11167 -13624 11201 -13590
rect 11235 -13624 11269 -13590
rect 11303 -13624 11337 -13590
rect 11371 -13624 11405 -13590
rect 11439 -13624 11473 -13590
rect 11507 -13607 11732 -13590
rect 11790 -13590 12750 -13552
rect 11790 -13607 12015 -13590
rect 11507 -13624 11546 -13607
rect 10958 -13640 11546 -13624
rect 11976 -13624 12015 -13607
rect 12049 -13624 12083 -13590
rect 12117 -13624 12151 -13590
rect 12185 -13624 12219 -13590
rect 12253 -13624 12287 -13590
rect 12321 -13624 12355 -13590
rect 12389 -13624 12423 -13590
rect 12457 -13624 12491 -13590
rect 12525 -13607 12750 -13590
rect 12808 -13590 13768 -13552
rect 12808 -13607 13033 -13590
rect 12525 -13624 12564 -13607
rect 11976 -13640 12564 -13624
rect 12994 -13624 13033 -13607
rect 13067 -13624 13101 -13590
rect 13135 -13624 13169 -13590
rect 13203 -13624 13237 -13590
rect 13271 -13624 13305 -13590
rect 13339 -13624 13373 -13590
rect 13407 -13624 13441 -13590
rect 13475 -13624 13509 -13590
rect 13543 -13607 13768 -13590
rect 13826 -13590 14786 -13552
rect 13826 -13607 14051 -13590
rect 13543 -13624 13582 -13607
rect 12994 -13640 13582 -13624
rect 14012 -13624 14051 -13607
rect 14085 -13624 14119 -13590
rect 14153 -13624 14187 -13590
rect 14221 -13624 14255 -13590
rect 14289 -13624 14323 -13590
rect 14357 -13624 14391 -13590
rect 14425 -13624 14459 -13590
rect 14493 -13624 14527 -13590
rect 14561 -13607 14786 -13590
rect 14844 -13590 15804 -13552
rect 14844 -13607 15069 -13590
rect 14561 -13624 14600 -13607
rect 14012 -13640 14600 -13624
rect 15030 -13624 15069 -13607
rect 15103 -13624 15137 -13590
rect 15171 -13624 15205 -13590
rect 15239 -13624 15273 -13590
rect 15307 -13624 15341 -13590
rect 15375 -13624 15409 -13590
rect 15443 -13624 15477 -13590
rect 15511 -13624 15545 -13590
rect 15579 -13607 15804 -13590
rect 15862 -13590 16822 -13552
rect 15862 -13607 16087 -13590
rect 15579 -13624 15618 -13607
rect 15030 -13640 15618 -13624
rect 16048 -13624 16087 -13607
rect 16121 -13624 16155 -13590
rect 16189 -13624 16223 -13590
rect 16257 -13624 16291 -13590
rect 16325 -13624 16359 -13590
rect 16393 -13624 16427 -13590
rect 16461 -13624 16495 -13590
rect 16529 -13624 16563 -13590
rect 16597 -13607 16822 -13590
rect 16880 -13590 17840 -13552
rect 16880 -13607 17105 -13590
rect 16597 -13624 16636 -13607
rect 16048 -13640 16636 -13624
rect 17066 -13624 17105 -13607
rect 17139 -13624 17173 -13590
rect 17207 -13624 17241 -13590
rect 17275 -13624 17309 -13590
rect 17343 -13624 17377 -13590
rect 17411 -13624 17445 -13590
rect 17479 -13624 17513 -13590
rect 17547 -13624 17581 -13590
rect 17615 -13607 17840 -13590
rect 17898 -13590 18858 -13552
rect 17898 -13607 18123 -13590
rect 17615 -13624 17654 -13607
rect 17066 -13640 17654 -13624
rect 18084 -13624 18123 -13607
rect 18157 -13624 18191 -13590
rect 18225 -13624 18259 -13590
rect 18293 -13624 18327 -13590
rect 18361 -13624 18395 -13590
rect 18429 -13624 18463 -13590
rect 18497 -13624 18531 -13590
rect 18565 -13624 18599 -13590
rect 18633 -13607 18858 -13590
rect 18916 -13590 19876 -13552
rect 18916 -13607 19141 -13590
rect 18633 -13624 18672 -13607
rect 18084 -13640 18672 -13624
rect 19102 -13624 19141 -13607
rect 19175 -13624 19209 -13590
rect 19243 -13624 19277 -13590
rect 19311 -13624 19345 -13590
rect 19379 -13624 19413 -13590
rect 19447 -13624 19481 -13590
rect 19515 -13624 19549 -13590
rect 19583 -13624 19617 -13590
rect 19651 -13607 19876 -13590
rect 19934 -13590 20894 -13552
rect 19934 -13607 20159 -13590
rect 19651 -13624 19690 -13607
rect 19102 -13640 19690 -13624
rect 20120 -13624 20159 -13607
rect 20193 -13624 20227 -13590
rect 20261 -13624 20295 -13590
rect 20329 -13624 20363 -13590
rect 20397 -13624 20431 -13590
rect 20465 -13624 20499 -13590
rect 20533 -13624 20567 -13590
rect 20601 -13624 20635 -13590
rect 20669 -13607 20894 -13590
rect 20952 -13590 21912 -13552
rect 20952 -13607 21177 -13590
rect 20669 -13624 20708 -13607
rect 20120 -13640 20708 -13624
rect 21138 -13624 21177 -13607
rect 21211 -13624 21245 -13590
rect 21279 -13624 21313 -13590
rect 21347 -13624 21381 -13590
rect 21415 -13624 21449 -13590
rect 21483 -13624 21517 -13590
rect 21551 -13624 21585 -13590
rect 21619 -13624 21653 -13590
rect 21687 -13607 21912 -13590
rect 21970 -13590 22930 -13552
rect 21970 -13607 22195 -13590
rect 21687 -13624 21726 -13607
rect 21138 -13640 21726 -13624
rect 22156 -13624 22195 -13607
rect 22229 -13624 22263 -13590
rect 22297 -13624 22331 -13590
rect 22365 -13624 22399 -13590
rect 22433 -13624 22467 -13590
rect 22501 -13624 22535 -13590
rect 22569 -13624 22603 -13590
rect 22637 -13624 22671 -13590
rect 22705 -13607 22930 -13590
rect 22705 -13624 22744 -13607
rect 22156 -13640 22744 -13624
rect -9138 -13968 -8178 -13930
rect -9138 -13985 -8913 -13968
rect -8952 -14002 -8913 -13985
rect -8879 -14002 -8845 -13968
rect -8811 -14002 -8777 -13968
rect -8743 -14002 -8709 -13968
rect -8675 -14002 -8641 -13968
rect -8607 -14002 -8573 -13968
rect -8539 -14002 -8505 -13968
rect -8471 -14002 -8437 -13968
rect -8403 -13985 -8178 -13968
rect -8120 -13968 -7160 -13930
rect -8120 -13985 -7895 -13968
rect -8403 -14002 -8364 -13985
rect -8952 -14018 -8364 -14002
rect -7934 -14002 -7895 -13985
rect -7861 -14002 -7827 -13968
rect -7793 -14002 -7759 -13968
rect -7725 -14002 -7691 -13968
rect -7657 -14002 -7623 -13968
rect -7589 -14002 -7555 -13968
rect -7521 -14002 -7487 -13968
rect -7453 -14002 -7419 -13968
rect -7385 -13985 -7160 -13968
rect -7102 -13968 -6142 -13930
rect -7102 -13985 -6877 -13968
rect -7385 -14002 -7346 -13985
rect -7934 -14018 -7346 -14002
rect -6916 -14002 -6877 -13985
rect -6843 -14002 -6809 -13968
rect -6775 -14002 -6741 -13968
rect -6707 -14002 -6673 -13968
rect -6639 -14002 -6605 -13968
rect -6571 -14002 -6537 -13968
rect -6503 -14002 -6469 -13968
rect -6435 -14002 -6401 -13968
rect -6367 -13985 -6142 -13968
rect -6084 -13968 -5124 -13930
rect -6084 -13985 -5859 -13968
rect -6367 -14002 -6328 -13985
rect -6916 -14018 -6328 -14002
rect -5898 -14002 -5859 -13985
rect -5825 -14002 -5791 -13968
rect -5757 -14002 -5723 -13968
rect -5689 -14002 -5655 -13968
rect -5621 -14002 -5587 -13968
rect -5553 -14002 -5519 -13968
rect -5485 -14002 -5451 -13968
rect -5417 -14002 -5383 -13968
rect -5349 -13985 -5124 -13968
rect -5066 -13968 -4106 -13930
rect -5066 -13985 -4841 -13968
rect -5349 -14002 -5310 -13985
rect -5898 -14018 -5310 -14002
rect -4880 -14002 -4841 -13985
rect -4807 -14002 -4773 -13968
rect -4739 -14002 -4705 -13968
rect -4671 -14002 -4637 -13968
rect -4603 -14002 -4569 -13968
rect -4535 -14002 -4501 -13968
rect -4467 -14002 -4433 -13968
rect -4399 -14002 -4365 -13968
rect -4331 -13985 -4106 -13968
rect -4048 -13968 -3088 -13930
rect -4048 -13985 -3823 -13968
rect -4331 -14002 -4292 -13985
rect -4880 -14018 -4292 -14002
rect -3862 -14002 -3823 -13985
rect -3789 -14002 -3755 -13968
rect -3721 -14002 -3687 -13968
rect -3653 -14002 -3619 -13968
rect -3585 -14002 -3551 -13968
rect -3517 -14002 -3483 -13968
rect -3449 -14002 -3415 -13968
rect -3381 -14002 -3347 -13968
rect -3313 -13985 -3088 -13968
rect -3030 -13968 -2070 -13930
rect -3030 -13985 -2805 -13968
rect -3313 -14002 -3274 -13985
rect -3862 -14018 -3274 -14002
rect -2844 -14002 -2805 -13985
rect -2771 -14002 -2737 -13968
rect -2703 -14002 -2669 -13968
rect -2635 -14002 -2601 -13968
rect -2567 -14002 -2533 -13968
rect -2499 -14002 -2465 -13968
rect -2431 -14002 -2397 -13968
rect -2363 -14002 -2329 -13968
rect -2295 -13985 -2070 -13968
rect -2012 -13968 -1052 -13930
rect -2012 -13985 -1787 -13968
rect -2295 -14002 -2256 -13985
rect -2844 -14018 -2256 -14002
rect -1826 -14002 -1787 -13985
rect -1753 -14002 -1719 -13968
rect -1685 -14002 -1651 -13968
rect -1617 -14002 -1583 -13968
rect -1549 -14002 -1515 -13968
rect -1481 -14002 -1447 -13968
rect -1413 -14002 -1379 -13968
rect -1345 -14002 -1311 -13968
rect -1277 -13985 -1052 -13968
rect -994 -13968 -34 -13930
rect -994 -13985 -769 -13968
rect -1277 -14002 -1238 -13985
rect -1826 -14018 -1238 -14002
rect -808 -14002 -769 -13985
rect -735 -14002 -701 -13968
rect -667 -14002 -633 -13968
rect -599 -14002 -565 -13968
rect -531 -14002 -497 -13968
rect -463 -14002 -429 -13968
rect -395 -14002 -361 -13968
rect -327 -14002 -293 -13968
rect -259 -13985 -34 -13968
rect -259 -14002 -220 -13985
rect -808 -14018 -220 -14002
rect -8952 -14076 -8364 -14060
rect -8952 -14093 -8913 -14076
rect -9138 -14110 -8913 -14093
rect -8879 -14110 -8845 -14076
rect -8811 -14110 -8777 -14076
rect -8743 -14110 -8709 -14076
rect -8675 -14110 -8641 -14076
rect -8607 -14110 -8573 -14076
rect -8539 -14110 -8505 -14076
rect -8471 -14110 -8437 -14076
rect -8403 -14093 -8364 -14076
rect -7934 -14076 -7346 -14060
rect -7934 -14093 -7895 -14076
rect -8403 -14110 -8178 -14093
rect -9138 -14148 -8178 -14110
rect -8120 -14110 -7895 -14093
rect -7861 -14110 -7827 -14076
rect -7793 -14110 -7759 -14076
rect -7725 -14110 -7691 -14076
rect -7657 -14110 -7623 -14076
rect -7589 -14110 -7555 -14076
rect -7521 -14110 -7487 -14076
rect -7453 -14110 -7419 -14076
rect -7385 -14093 -7346 -14076
rect -6916 -14076 -6328 -14060
rect -6916 -14093 -6877 -14076
rect -7385 -14110 -7160 -14093
rect -8120 -14148 -7160 -14110
rect -7102 -14110 -6877 -14093
rect -6843 -14110 -6809 -14076
rect -6775 -14110 -6741 -14076
rect -6707 -14110 -6673 -14076
rect -6639 -14110 -6605 -14076
rect -6571 -14110 -6537 -14076
rect -6503 -14110 -6469 -14076
rect -6435 -14110 -6401 -14076
rect -6367 -14093 -6328 -14076
rect -5898 -14076 -5310 -14060
rect -5898 -14093 -5859 -14076
rect -6367 -14110 -6142 -14093
rect -7102 -14148 -6142 -14110
rect -6084 -14110 -5859 -14093
rect -5825 -14110 -5791 -14076
rect -5757 -14110 -5723 -14076
rect -5689 -14110 -5655 -14076
rect -5621 -14110 -5587 -14076
rect -5553 -14110 -5519 -14076
rect -5485 -14110 -5451 -14076
rect -5417 -14110 -5383 -14076
rect -5349 -14093 -5310 -14076
rect -4880 -14076 -4292 -14060
rect -4880 -14093 -4841 -14076
rect -5349 -14110 -5124 -14093
rect -6084 -14148 -5124 -14110
rect -5066 -14110 -4841 -14093
rect -4807 -14110 -4773 -14076
rect -4739 -14110 -4705 -14076
rect -4671 -14110 -4637 -14076
rect -4603 -14110 -4569 -14076
rect -4535 -14110 -4501 -14076
rect -4467 -14110 -4433 -14076
rect -4399 -14110 -4365 -14076
rect -4331 -14093 -4292 -14076
rect -3862 -14076 -3274 -14060
rect -3862 -14093 -3823 -14076
rect -4331 -14110 -4106 -14093
rect -5066 -14148 -4106 -14110
rect -4048 -14110 -3823 -14093
rect -3789 -14110 -3755 -14076
rect -3721 -14110 -3687 -14076
rect -3653 -14110 -3619 -14076
rect -3585 -14110 -3551 -14076
rect -3517 -14110 -3483 -14076
rect -3449 -14110 -3415 -14076
rect -3381 -14110 -3347 -14076
rect -3313 -14093 -3274 -14076
rect -2844 -14076 -2256 -14060
rect -2844 -14093 -2805 -14076
rect -3313 -14110 -3088 -14093
rect -4048 -14148 -3088 -14110
rect -3030 -14110 -2805 -14093
rect -2771 -14110 -2737 -14076
rect -2703 -14110 -2669 -14076
rect -2635 -14110 -2601 -14076
rect -2567 -14110 -2533 -14076
rect -2499 -14110 -2465 -14076
rect -2431 -14110 -2397 -14076
rect -2363 -14110 -2329 -14076
rect -2295 -14093 -2256 -14076
rect -1826 -14076 -1238 -14060
rect -1826 -14093 -1787 -14076
rect -2295 -14110 -2070 -14093
rect -3030 -14148 -2070 -14110
rect -2012 -14110 -1787 -14093
rect -1753 -14110 -1719 -14076
rect -1685 -14110 -1651 -14076
rect -1617 -14110 -1583 -14076
rect -1549 -14110 -1515 -14076
rect -1481 -14110 -1447 -14076
rect -1413 -14110 -1379 -14076
rect -1345 -14110 -1311 -14076
rect -1277 -14093 -1238 -14076
rect -808 -14076 -220 -14060
rect -808 -14093 -769 -14076
rect -1277 -14110 -1052 -14093
rect -2012 -14148 -1052 -14110
rect -994 -14110 -769 -14093
rect -735 -14110 -701 -14076
rect -667 -14110 -633 -14076
rect -599 -14110 -565 -14076
rect -531 -14110 -497 -14076
rect -463 -14110 -429 -14076
rect -395 -14110 -361 -14076
rect -327 -14110 -293 -14076
rect -259 -14093 -220 -14076
rect -259 -14110 -34 -14093
rect -994 -14148 -34 -14110
rect 2814 -14112 3402 -14096
rect 2814 -14129 2853 -14112
rect 2628 -14146 2853 -14129
rect 2887 -14146 2921 -14112
rect 2955 -14146 2989 -14112
rect 3023 -14146 3057 -14112
rect 3091 -14146 3125 -14112
rect 3159 -14146 3193 -14112
rect 3227 -14146 3261 -14112
rect 3295 -14146 3329 -14112
rect 3363 -14129 3402 -14112
rect 3832 -14112 4420 -14096
rect 3832 -14129 3871 -14112
rect 3363 -14146 3588 -14129
rect 2628 -14184 3588 -14146
rect 3646 -14146 3871 -14129
rect 3905 -14146 3939 -14112
rect 3973 -14146 4007 -14112
rect 4041 -14146 4075 -14112
rect 4109 -14146 4143 -14112
rect 4177 -14146 4211 -14112
rect 4245 -14146 4279 -14112
rect 4313 -14146 4347 -14112
rect 4381 -14129 4420 -14112
rect 4850 -14112 5438 -14096
rect 4850 -14129 4889 -14112
rect 4381 -14146 4606 -14129
rect 3646 -14184 4606 -14146
rect 4664 -14146 4889 -14129
rect 4923 -14146 4957 -14112
rect 4991 -14146 5025 -14112
rect 5059 -14146 5093 -14112
rect 5127 -14146 5161 -14112
rect 5195 -14146 5229 -14112
rect 5263 -14146 5297 -14112
rect 5331 -14146 5365 -14112
rect 5399 -14129 5438 -14112
rect 5868 -14112 6456 -14096
rect 5868 -14129 5907 -14112
rect 5399 -14146 5624 -14129
rect 4664 -14184 5624 -14146
rect 5682 -14146 5907 -14129
rect 5941 -14146 5975 -14112
rect 6009 -14146 6043 -14112
rect 6077 -14146 6111 -14112
rect 6145 -14146 6179 -14112
rect 6213 -14146 6247 -14112
rect 6281 -14146 6315 -14112
rect 6349 -14146 6383 -14112
rect 6417 -14129 6456 -14112
rect 6886 -14112 7474 -14096
rect 6886 -14129 6925 -14112
rect 6417 -14146 6642 -14129
rect 5682 -14184 6642 -14146
rect 6700 -14146 6925 -14129
rect 6959 -14146 6993 -14112
rect 7027 -14146 7061 -14112
rect 7095 -14146 7129 -14112
rect 7163 -14146 7197 -14112
rect 7231 -14146 7265 -14112
rect 7299 -14146 7333 -14112
rect 7367 -14146 7401 -14112
rect 7435 -14129 7474 -14112
rect 7904 -14112 8492 -14096
rect 7904 -14129 7943 -14112
rect 7435 -14146 7660 -14129
rect 6700 -14184 7660 -14146
rect 7718 -14146 7943 -14129
rect 7977 -14146 8011 -14112
rect 8045 -14146 8079 -14112
rect 8113 -14146 8147 -14112
rect 8181 -14146 8215 -14112
rect 8249 -14146 8283 -14112
rect 8317 -14146 8351 -14112
rect 8385 -14146 8419 -14112
rect 8453 -14129 8492 -14112
rect 8922 -14112 9510 -14096
rect 8922 -14129 8961 -14112
rect 8453 -14146 8678 -14129
rect 7718 -14184 8678 -14146
rect 8736 -14146 8961 -14129
rect 8995 -14146 9029 -14112
rect 9063 -14146 9097 -14112
rect 9131 -14146 9165 -14112
rect 9199 -14146 9233 -14112
rect 9267 -14146 9301 -14112
rect 9335 -14146 9369 -14112
rect 9403 -14146 9437 -14112
rect 9471 -14129 9510 -14112
rect 9940 -14112 10528 -14096
rect 9940 -14129 9979 -14112
rect 9471 -14146 9696 -14129
rect 8736 -14184 9696 -14146
rect 9754 -14146 9979 -14129
rect 10013 -14146 10047 -14112
rect 10081 -14146 10115 -14112
rect 10149 -14146 10183 -14112
rect 10217 -14146 10251 -14112
rect 10285 -14146 10319 -14112
rect 10353 -14146 10387 -14112
rect 10421 -14146 10455 -14112
rect 10489 -14129 10528 -14112
rect 10958 -14112 11546 -14096
rect 10958 -14129 10997 -14112
rect 10489 -14146 10714 -14129
rect 9754 -14184 10714 -14146
rect 10772 -14146 10997 -14129
rect 11031 -14146 11065 -14112
rect 11099 -14146 11133 -14112
rect 11167 -14146 11201 -14112
rect 11235 -14146 11269 -14112
rect 11303 -14146 11337 -14112
rect 11371 -14146 11405 -14112
rect 11439 -14146 11473 -14112
rect 11507 -14129 11546 -14112
rect 11976 -14112 12564 -14096
rect 11976 -14129 12015 -14112
rect 11507 -14146 11732 -14129
rect 10772 -14184 11732 -14146
rect 11790 -14146 12015 -14129
rect 12049 -14146 12083 -14112
rect 12117 -14146 12151 -14112
rect 12185 -14146 12219 -14112
rect 12253 -14146 12287 -14112
rect 12321 -14146 12355 -14112
rect 12389 -14146 12423 -14112
rect 12457 -14146 12491 -14112
rect 12525 -14129 12564 -14112
rect 12994 -14112 13582 -14096
rect 12994 -14129 13033 -14112
rect 12525 -14146 12750 -14129
rect 11790 -14184 12750 -14146
rect 12808 -14146 13033 -14129
rect 13067 -14146 13101 -14112
rect 13135 -14146 13169 -14112
rect 13203 -14146 13237 -14112
rect 13271 -14146 13305 -14112
rect 13339 -14146 13373 -14112
rect 13407 -14146 13441 -14112
rect 13475 -14146 13509 -14112
rect 13543 -14129 13582 -14112
rect 14012 -14112 14600 -14096
rect 14012 -14129 14051 -14112
rect 13543 -14146 13768 -14129
rect 12808 -14184 13768 -14146
rect 13826 -14146 14051 -14129
rect 14085 -14146 14119 -14112
rect 14153 -14146 14187 -14112
rect 14221 -14146 14255 -14112
rect 14289 -14146 14323 -14112
rect 14357 -14146 14391 -14112
rect 14425 -14146 14459 -14112
rect 14493 -14146 14527 -14112
rect 14561 -14129 14600 -14112
rect 15030 -14112 15618 -14096
rect 15030 -14129 15069 -14112
rect 14561 -14146 14786 -14129
rect 13826 -14184 14786 -14146
rect 14844 -14146 15069 -14129
rect 15103 -14146 15137 -14112
rect 15171 -14146 15205 -14112
rect 15239 -14146 15273 -14112
rect 15307 -14146 15341 -14112
rect 15375 -14146 15409 -14112
rect 15443 -14146 15477 -14112
rect 15511 -14146 15545 -14112
rect 15579 -14129 15618 -14112
rect 16048 -14112 16636 -14096
rect 16048 -14129 16087 -14112
rect 15579 -14146 15804 -14129
rect 14844 -14184 15804 -14146
rect 15862 -14146 16087 -14129
rect 16121 -14146 16155 -14112
rect 16189 -14146 16223 -14112
rect 16257 -14146 16291 -14112
rect 16325 -14146 16359 -14112
rect 16393 -14146 16427 -14112
rect 16461 -14146 16495 -14112
rect 16529 -14146 16563 -14112
rect 16597 -14129 16636 -14112
rect 17066 -14112 17654 -14096
rect 17066 -14129 17105 -14112
rect 16597 -14146 16822 -14129
rect 15862 -14184 16822 -14146
rect 16880 -14146 17105 -14129
rect 17139 -14146 17173 -14112
rect 17207 -14146 17241 -14112
rect 17275 -14146 17309 -14112
rect 17343 -14146 17377 -14112
rect 17411 -14146 17445 -14112
rect 17479 -14146 17513 -14112
rect 17547 -14146 17581 -14112
rect 17615 -14129 17654 -14112
rect 18084 -14112 18672 -14096
rect 18084 -14129 18123 -14112
rect 17615 -14146 17840 -14129
rect 16880 -14184 17840 -14146
rect 17898 -14146 18123 -14129
rect 18157 -14146 18191 -14112
rect 18225 -14146 18259 -14112
rect 18293 -14146 18327 -14112
rect 18361 -14146 18395 -14112
rect 18429 -14146 18463 -14112
rect 18497 -14146 18531 -14112
rect 18565 -14146 18599 -14112
rect 18633 -14129 18672 -14112
rect 19102 -14112 19690 -14096
rect 19102 -14129 19141 -14112
rect 18633 -14146 18858 -14129
rect 17898 -14184 18858 -14146
rect 18916 -14146 19141 -14129
rect 19175 -14146 19209 -14112
rect 19243 -14146 19277 -14112
rect 19311 -14146 19345 -14112
rect 19379 -14146 19413 -14112
rect 19447 -14146 19481 -14112
rect 19515 -14146 19549 -14112
rect 19583 -14146 19617 -14112
rect 19651 -14129 19690 -14112
rect 20120 -14112 20708 -14096
rect 20120 -14129 20159 -14112
rect 19651 -14146 19876 -14129
rect 18916 -14184 19876 -14146
rect 19934 -14146 20159 -14129
rect 20193 -14146 20227 -14112
rect 20261 -14146 20295 -14112
rect 20329 -14146 20363 -14112
rect 20397 -14146 20431 -14112
rect 20465 -14146 20499 -14112
rect 20533 -14146 20567 -14112
rect 20601 -14146 20635 -14112
rect 20669 -14129 20708 -14112
rect 21138 -14112 21726 -14096
rect 21138 -14129 21177 -14112
rect 20669 -14146 20894 -14129
rect 19934 -14184 20894 -14146
rect 20952 -14146 21177 -14129
rect 21211 -14146 21245 -14112
rect 21279 -14146 21313 -14112
rect 21347 -14146 21381 -14112
rect 21415 -14146 21449 -14112
rect 21483 -14146 21517 -14112
rect 21551 -14146 21585 -14112
rect 21619 -14146 21653 -14112
rect 21687 -14129 21726 -14112
rect 22156 -14112 22744 -14096
rect 22156 -14129 22195 -14112
rect 21687 -14146 21912 -14129
rect 20952 -14184 21912 -14146
rect 21970 -14146 22195 -14129
rect 22229 -14146 22263 -14112
rect 22297 -14146 22331 -14112
rect 22365 -14146 22399 -14112
rect 22433 -14146 22467 -14112
rect 22501 -14146 22535 -14112
rect 22569 -14146 22603 -14112
rect 22637 -14146 22671 -14112
rect 22705 -14129 22744 -14112
rect 22705 -14146 22930 -14129
rect 21970 -14184 22930 -14146
rect -9138 -14786 -8178 -14748
rect -9138 -14803 -8913 -14786
rect -8952 -14820 -8913 -14803
rect -8879 -14820 -8845 -14786
rect -8811 -14820 -8777 -14786
rect -8743 -14820 -8709 -14786
rect -8675 -14820 -8641 -14786
rect -8607 -14820 -8573 -14786
rect -8539 -14820 -8505 -14786
rect -8471 -14820 -8437 -14786
rect -8403 -14803 -8178 -14786
rect -8120 -14786 -7160 -14748
rect -8120 -14803 -7895 -14786
rect -8403 -14820 -8364 -14803
rect -8952 -14836 -8364 -14820
rect -7934 -14820 -7895 -14803
rect -7861 -14820 -7827 -14786
rect -7793 -14820 -7759 -14786
rect -7725 -14820 -7691 -14786
rect -7657 -14820 -7623 -14786
rect -7589 -14820 -7555 -14786
rect -7521 -14820 -7487 -14786
rect -7453 -14820 -7419 -14786
rect -7385 -14803 -7160 -14786
rect -7102 -14786 -6142 -14748
rect -7102 -14803 -6877 -14786
rect -7385 -14820 -7346 -14803
rect -7934 -14836 -7346 -14820
rect -6916 -14820 -6877 -14803
rect -6843 -14820 -6809 -14786
rect -6775 -14820 -6741 -14786
rect -6707 -14820 -6673 -14786
rect -6639 -14820 -6605 -14786
rect -6571 -14820 -6537 -14786
rect -6503 -14820 -6469 -14786
rect -6435 -14820 -6401 -14786
rect -6367 -14803 -6142 -14786
rect -6084 -14786 -5124 -14748
rect -6084 -14803 -5859 -14786
rect -6367 -14820 -6328 -14803
rect -6916 -14836 -6328 -14820
rect -5898 -14820 -5859 -14803
rect -5825 -14820 -5791 -14786
rect -5757 -14820 -5723 -14786
rect -5689 -14820 -5655 -14786
rect -5621 -14820 -5587 -14786
rect -5553 -14820 -5519 -14786
rect -5485 -14820 -5451 -14786
rect -5417 -14820 -5383 -14786
rect -5349 -14803 -5124 -14786
rect -5066 -14786 -4106 -14748
rect -5066 -14803 -4841 -14786
rect -5349 -14820 -5310 -14803
rect -5898 -14836 -5310 -14820
rect -4880 -14820 -4841 -14803
rect -4807 -14820 -4773 -14786
rect -4739 -14820 -4705 -14786
rect -4671 -14820 -4637 -14786
rect -4603 -14820 -4569 -14786
rect -4535 -14820 -4501 -14786
rect -4467 -14820 -4433 -14786
rect -4399 -14820 -4365 -14786
rect -4331 -14803 -4106 -14786
rect -4048 -14786 -3088 -14748
rect -4048 -14803 -3823 -14786
rect -4331 -14820 -4292 -14803
rect -4880 -14836 -4292 -14820
rect -3862 -14820 -3823 -14803
rect -3789 -14820 -3755 -14786
rect -3721 -14820 -3687 -14786
rect -3653 -14820 -3619 -14786
rect -3585 -14820 -3551 -14786
rect -3517 -14820 -3483 -14786
rect -3449 -14820 -3415 -14786
rect -3381 -14820 -3347 -14786
rect -3313 -14803 -3088 -14786
rect -3030 -14786 -2070 -14748
rect -3030 -14803 -2805 -14786
rect -3313 -14820 -3274 -14803
rect -3862 -14836 -3274 -14820
rect -2844 -14820 -2805 -14803
rect -2771 -14820 -2737 -14786
rect -2703 -14820 -2669 -14786
rect -2635 -14820 -2601 -14786
rect -2567 -14820 -2533 -14786
rect -2499 -14820 -2465 -14786
rect -2431 -14820 -2397 -14786
rect -2363 -14820 -2329 -14786
rect -2295 -14803 -2070 -14786
rect -2012 -14786 -1052 -14748
rect -2012 -14803 -1787 -14786
rect -2295 -14820 -2256 -14803
rect -2844 -14836 -2256 -14820
rect -1826 -14820 -1787 -14803
rect -1753 -14820 -1719 -14786
rect -1685 -14820 -1651 -14786
rect -1617 -14820 -1583 -14786
rect -1549 -14820 -1515 -14786
rect -1481 -14820 -1447 -14786
rect -1413 -14820 -1379 -14786
rect -1345 -14820 -1311 -14786
rect -1277 -14803 -1052 -14786
rect -994 -14786 -34 -14748
rect -994 -14803 -769 -14786
rect -1277 -14820 -1238 -14803
rect -1826 -14836 -1238 -14820
rect -808 -14820 -769 -14803
rect -735 -14820 -701 -14786
rect -667 -14820 -633 -14786
rect -599 -14820 -565 -14786
rect -531 -14820 -497 -14786
rect -463 -14820 -429 -14786
rect -395 -14820 -361 -14786
rect -327 -14820 -293 -14786
rect -259 -14803 -34 -14786
rect -259 -14820 -220 -14803
rect -808 -14836 -220 -14820
rect 2628 -14822 3588 -14784
rect 2628 -14839 2853 -14822
rect 2814 -14856 2853 -14839
rect 2887 -14856 2921 -14822
rect 2955 -14856 2989 -14822
rect 3023 -14856 3057 -14822
rect 3091 -14856 3125 -14822
rect 3159 -14856 3193 -14822
rect 3227 -14856 3261 -14822
rect 3295 -14856 3329 -14822
rect 3363 -14839 3588 -14822
rect 3646 -14822 4606 -14784
rect 3646 -14839 3871 -14822
rect 3363 -14856 3402 -14839
rect 2814 -14872 3402 -14856
rect 3832 -14856 3871 -14839
rect 3905 -14856 3939 -14822
rect 3973 -14856 4007 -14822
rect 4041 -14856 4075 -14822
rect 4109 -14856 4143 -14822
rect 4177 -14856 4211 -14822
rect 4245 -14856 4279 -14822
rect 4313 -14856 4347 -14822
rect 4381 -14839 4606 -14822
rect 4664 -14822 5624 -14784
rect 4664 -14839 4889 -14822
rect 4381 -14856 4420 -14839
rect 3832 -14872 4420 -14856
rect 4850 -14856 4889 -14839
rect 4923 -14856 4957 -14822
rect 4991 -14856 5025 -14822
rect 5059 -14856 5093 -14822
rect 5127 -14856 5161 -14822
rect 5195 -14856 5229 -14822
rect 5263 -14856 5297 -14822
rect 5331 -14856 5365 -14822
rect 5399 -14839 5624 -14822
rect 5682 -14822 6642 -14784
rect 5682 -14839 5907 -14822
rect 5399 -14856 5438 -14839
rect 4850 -14872 5438 -14856
rect 5868 -14856 5907 -14839
rect 5941 -14856 5975 -14822
rect 6009 -14856 6043 -14822
rect 6077 -14856 6111 -14822
rect 6145 -14856 6179 -14822
rect 6213 -14856 6247 -14822
rect 6281 -14856 6315 -14822
rect 6349 -14856 6383 -14822
rect 6417 -14839 6642 -14822
rect 6700 -14822 7660 -14784
rect 6700 -14839 6925 -14822
rect 6417 -14856 6456 -14839
rect 5868 -14872 6456 -14856
rect 6886 -14856 6925 -14839
rect 6959 -14856 6993 -14822
rect 7027 -14856 7061 -14822
rect 7095 -14856 7129 -14822
rect 7163 -14856 7197 -14822
rect 7231 -14856 7265 -14822
rect 7299 -14856 7333 -14822
rect 7367 -14856 7401 -14822
rect 7435 -14839 7660 -14822
rect 7718 -14822 8678 -14784
rect 7718 -14839 7943 -14822
rect 7435 -14856 7474 -14839
rect 6886 -14872 7474 -14856
rect 7904 -14856 7943 -14839
rect 7977 -14856 8011 -14822
rect 8045 -14856 8079 -14822
rect 8113 -14856 8147 -14822
rect 8181 -14856 8215 -14822
rect 8249 -14856 8283 -14822
rect 8317 -14856 8351 -14822
rect 8385 -14856 8419 -14822
rect 8453 -14839 8678 -14822
rect 8736 -14822 9696 -14784
rect 8736 -14839 8961 -14822
rect 8453 -14856 8492 -14839
rect 7904 -14872 8492 -14856
rect 8922 -14856 8961 -14839
rect 8995 -14856 9029 -14822
rect 9063 -14856 9097 -14822
rect 9131 -14856 9165 -14822
rect 9199 -14856 9233 -14822
rect 9267 -14856 9301 -14822
rect 9335 -14856 9369 -14822
rect 9403 -14856 9437 -14822
rect 9471 -14839 9696 -14822
rect 9754 -14822 10714 -14784
rect 9754 -14839 9979 -14822
rect 9471 -14856 9510 -14839
rect 8922 -14872 9510 -14856
rect 9940 -14856 9979 -14839
rect 10013 -14856 10047 -14822
rect 10081 -14856 10115 -14822
rect 10149 -14856 10183 -14822
rect 10217 -14856 10251 -14822
rect 10285 -14856 10319 -14822
rect 10353 -14856 10387 -14822
rect 10421 -14856 10455 -14822
rect 10489 -14839 10714 -14822
rect 10772 -14822 11732 -14784
rect 10772 -14839 10997 -14822
rect 10489 -14856 10528 -14839
rect 9940 -14872 10528 -14856
rect 10958 -14856 10997 -14839
rect 11031 -14856 11065 -14822
rect 11099 -14856 11133 -14822
rect 11167 -14856 11201 -14822
rect 11235 -14856 11269 -14822
rect 11303 -14856 11337 -14822
rect 11371 -14856 11405 -14822
rect 11439 -14856 11473 -14822
rect 11507 -14839 11732 -14822
rect 11790 -14822 12750 -14784
rect 11790 -14839 12015 -14822
rect 11507 -14856 11546 -14839
rect 10958 -14872 11546 -14856
rect 11976 -14856 12015 -14839
rect 12049 -14856 12083 -14822
rect 12117 -14856 12151 -14822
rect 12185 -14856 12219 -14822
rect 12253 -14856 12287 -14822
rect 12321 -14856 12355 -14822
rect 12389 -14856 12423 -14822
rect 12457 -14856 12491 -14822
rect 12525 -14839 12750 -14822
rect 12808 -14822 13768 -14784
rect 12808 -14839 13033 -14822
rect 12525 -14856 12564 -14839
rect 11976 -14872 12564 -14856
rect 12994 -14856 13033 -14839
rect 13067 -14856 13101 -14822
rect 13135 -14856 13169 -14822
rect 13203 -14856 13237 -14822
rect 13271 -14856 13305 -14822
rect 13339 -14856 13373 -14822
rect 13407 -14856 13441 -14822
rect 13475 -14856 13509 -14822
rect 13543 -14839 13768 -14822
rect 13826 -14822 14786 -14784
rect 13826 -14839 14051 -14822
rect 13543 -14856 13582 -14839
rect 12994 -14872 13582 -14856
rect 14012 -14856 14051 -14839
rect 14085 -14856 14119 -14822
rect 14153 -14856 14187 -14822
rect 14221 -14856 14255 -14822
rect 14289 -14856 14323 -14822
rect 14357 -14856 14391 -14822
rect 14425 -14856 14459 -14822
rect 14493 -14856 14527 -14822
rect 14561 -14839 14786 -14822
rect 14844 -14822 15804 -14784
rect 14844 -14839 15069 -14822
rect 14561 -14856 14600 -14839
rect 14012 -14872 14600 -14856
rect 15030 -14856 15069 -14839
rect 15103 -14856 15137 -14822
rect 15171 -14856 15205 -14822
rect 15239 -14856 15273 -14822
rect 15307 -14856 15341 -14822
rect 15375 -14856 15409 -14822
rect 15443 -14856 15477 -14822
rect 15511 -14856 15545 -14822
rect 15579 -14839 15804 -14822
rect 15862 -14822 16822 -14784
rect 15862 -14839 16087 -14822
rect 15579 -14856 15618 -14839
rect 15030 -14872 15618 -14856
rect 16048 -14856 16087 -14839
rect 16121 -14856 16155 -14822
rect 16189 -14856 16223 -14822
rect 16257 -14856 16291 -14822
rect 16325 -14856 16359 -14822
rect 16393 -14856 16427 -14822
rect 16461 -14856 16495 -14822
rect 16529 -14856 16563 -14822
rect 16597 -14839 16822 -14822
rect 16880 -14822 17840 -14784
rect 16880 -14839 17105 -14822
rect 16597 -14856 16636 -14839
rect 16048 -14872 16636 -14856
rect 17066 -14856 17105 -14839
rect 17139 -14856 17173 -14822
rect 17207 -14856 17241 -14822
rect 17275 -14856 17309 -14822
rect 17343 -14856 17377 -14822
rect 17411 -14856 17445 -14822
rect 17479 -14856 17513 -14822
rect 17547 -14856 17581 -14822
rect 17615 -14839 17840 -14822
rect 17898 -14822 18858 -14784
rect 17898 -14839 18123 -14822
rect 17615 -14856 17654 -14839
rect 17066 -14872 17654 -14856
rect 18084 -14856 18123 -14839
rect 18157 -14856 18191 -14822
rect 18225 -14856 18259 -14822
rect 18293 -14856 18327 -14822
rect 18361 -14856 18395 -14822
rect 18429 -14856 18463 -14822
rect 18497 -14856 18531 -14822
rect 18565 -14856 18599 -14822
rect 18633 -14839 18858 -14822
rect 18916 -14822 19876 -14784
rect 18916 -14839 19141 -14822
rect 18633 -14856 18672 -14839
rect 18084 -14872 18672 -14856
rect 19102 -14856 19141 -14839
rect 19175 -14856 19209 -14822
rect 19243 -14856 19277 -14822
rect 19311 -14856 19345 -14822
rect 19379 -14856 19413 -14822
rect 19447 -14856 19481 -14822
rect 19515 -14856 19549 -14822
rect 19583 -14856 19617 -14822
rect 19651 -14839 19876 -14822
rect 19934 -14822 20894 -14784
rect 19934 -14839 20159 -14822
rect 19651 -14856 19690 -14839
rect 19102 -14872 19690 -14856
rect 20120 -14856 20159 -14839
rect 20193 -14856 20227 -14822
rect 20261 -14856 20295 -14822
rect 20329 -14856 20363 -14822
rect 20397 -14856 20431 -14822
rect 20465 -14856 20499 -14822
rect 20533 -14856 20567 -14822
rect 20601 -14856 20635 -14822
rect 20669 -14839 20894 -14822
rect 20952 -14822 21912 -14784
rect 20952 -14839 21177 -14822
rect 20669 -14856 20708 -14839
rect 20120 -14872 20708 -14856
rect 21138 -14856 21177 -14839
rect 21211 -14856 21245 -14822
rect 21279 -14856 21313 -14822
rect 21347 -14856 21381 -14822
rect 21415 -14856 21449 -14822
rect 21483 -14856 21517 -14822
rect 21551 -14856 21585 -14822
rect 21619 -14856 21653 -14822
rect 21687 -14839 21912 -14822
rect 21970 -14822 22930 -14784
rect 21970 -14839 22195 -14822
rect 21687 -14856 21726 -14839
rect 21138 -14872 21726 -14856
rect 22156 -14856 22195 -14839
rect 22229 -14856 22263 -14822
rect 22297 -14856 22331 -14822
rect 22365 -14856 22399 -14822
rect 22433 -14856 22467 -14822
rect 22501 -14856 22535 -14822
rect 22569 -14856 22603 -14822
rect 22637 -14856 22671 -14822
rect 22705 -14839 22930 -14822
rect 22705 -14856 22744 -14839
rect 22156 -14872 22744 -14856
rect -8952 -14894 -8364 -14878
rect -8952 -14911 -8913 -14894
rect -9138 -14928 -8913 -14911
rect -8879 -14928 -8845 -14894
rect -8811 -14928 -8777 -14894
rect -8743 -14928 -8709 -14894
rect -8675 -14928 -8641 -14894
rect -8607 -14928 -8573 -14894
rect -8539 -14928 -8505 -14894
rect -8471 -14928 -8437 -14894
rect -8403 -14911 -8364 -14894
rect -7934 -14894 -7346 -14878
rect -7934 -14911 -7895 -14894
rect -8403 -14928 -8178 -14911
rect -9138 -14966 -8178 -14928
rect -8120 -14928 -7895 -14911
rect -7861 -14928 -7827 -14894
rect -7793 -14928 -7759 -14894
rect -7725 -14928 -7691 -14894
rect -7657 -14928 -7623 -14894
rect -7589 -14928 -7555 -14894
rect -7521 -14928 -7487 -14894
rect -7453 -14928 -7419 -14894
rect -7385 -14911 -7346 -14894
rect -6916 -14894 -6328 -14878
rect -6916 -14911 -6877 -14894
rect -7385 -14928 -7160 -14911
rect -8120 -14966 -7160 -14928
rect -7102 -14928 -6877 -14911
rect -6843 -14928 -6809 -14894
rect -6775 -14928 -6741 -14894
rect -6707 -14928 -6673 -14894
rect -6639 -14928 -6605 -14894
rect -6571 -14928 -6537 -14894
rect -6503 -14928 -6469 -14894
rect -6435 -14928 -6401 -14894
rect -6367 -14911 -6328 -14894
rect -5898 -14894 -5310 -14878
rect -5898 -14911 -5859 -14894
rect -6367 -14928 -6142 -14911
rect -7102 -14966 -6142 -14928
rect -6084 -14928 -5859 -14911
rect -5825 -14928 -5791 -14894
rect -5757 -14928 -5723 -14894
rect -5689 -14928 -5655 -14894
rect -5621 -14928 -5587 -14894
rect -5553 -14928 -5519 -14894
rect -5485 -14928 -5451 -14894
rect -5417 -14928 -5383 -14894
rect -5349 -14911 -5310 -14894
rect -4880 -14894 -4292 -14878
rect -4880 -14911 -4841 -14894
rect -5349 -14928 -5124 -14911
rect -6084 -14966 -5124 -14928
rect -5066 -14928 -4841 -14911
rect -4807 -14928 -4773 -14894
rect -4739 -14928 -4705 -14894
rect -4671 -14928 -4637 -14894
rect -4603 -14928 -4569 -14894
rect -4535 -14928 -4501 -14894
rect -4467 -14928 -4433 -14894
rect -4399 -14928 -4365 -14894
rect -4331 -14911 -4292 -14894
rect -3862 -14894 -3274 -14878
rect -3862 -14911 -3823 -14894
rect -4331 -14928 -4106 -14911
rect -5066 -14966 -4106 -14928
rect -4048 -14928 -3823 -14911
rect -3789 -14928 -3755 -14894
rect -3721 -14928 -3687 -14894
rect -3653 -14928 -3619 -14894
rect -3585 -14928 -3551 -14894
rect -3517 -14928 -3483 -14894
rect -3449 -14928 -3415 -14894
rect -3381 -14928 -3347 -14894
rect -3313 -14911 -3274 -14894
rect -2844 -14894 -2256 -14878
rect -2844 -14911 -2805 -14894
rect -3313 -14928 -3088 -14911
rect -4048 -14966 -3088 -14928
rect -3030 -14928 -2805 -14911
rect -2771 -14928 -2737 -14894
rect -2703 -14928 -2669 -14894
rect -2635 -14928 -2601 -14894
rect -2567 -14928 -2533 -14894
rect -2499 -14928 -2465 -14894
rect -2431 -14928 -2397 -14894
rect -2363 -14928 -2329 -14894
rect -2295 -14911 -2256 -14894
rect -1826 -14894 -1238 -14878
rect -1826 -14911 -1787 -14894
rect -2295 -14928 -2070 -14911
rect -3030 -14966 -2070 -14928
rect -2012 -14928 -1787 -14911
rect -1753 -14928 -1719 -14894
rect -1685 -14928 -1651 -14894
rect -1617 -14928 -1583 -14894
rect -1549 -14928 -1515 -14894
rect -1481 -14928 -1447 -14894
rect -1413 -14928 -1379 -14894
rect -1345 -14928 -1311 -14894
rect -1277 -14911 -1238 -14894
rect -808 -14894 -220 -14878
rect -808 -14911 -769 -14894
rect -1277 -14928 -1052 -14911
rect -2012 -14966 -1052 -14928
rect -994 -14928 -769 -14911
rect -735 -14928 -701 -14894
rect -667 -14928 -633 -14894
rect -599 -14928 -565 -14894
rect -531 -14928 -497 -14894
rect -463 -14928 -429 -14894
rect -395 -14928 -361 -14894
rect -327 -14928 -293 -14894
rect -259 -14911 -220 -14894
rect -259 -14928 -34 -14911
rect -994 -14966 -34 -14928
rect 2812 -15346 3400 -15330
rect 2812 -15363 2851 -15346
rect 2626 -15380 2851 -15363
rect 2885 -15380 2919 -15346
rect 2953 -15380 2987 -15346
rect 3021 -15380 3055 -15346
rect 3089 -15380 3123 -15346
rect 3157 -15380 3191 -15346
rect 3225 -15380 3259 -15346
rect 3293 -15380 3327 -15346
rect 3361 -15363 3400 -15346
rect 3830 -15346 4418 -15330
rect 3830 -15363 3869 -15346
rect 3361 -15380 3586 -15363
rect 2626 -15418 3586 -15380
rect 3644 -15380 3869 -15363
rect 3903 -15380 3937 -15346
rect 3971 -15380 4005 -15346
rect 4039 -15380 4073 -15346
rect 4107 -15380 4141 -15346
rect 4175 -15380 4209 -15346
rect 4243 -15380 4277 -15346
rect 4311 -15380 4345 -15346
rect 4379 -15363 4418 -15346
rect 4848 -15346 5436 -15330
rect 4848 -15363 4887 -15346
rect 4379 -15380 4604 -15363
rect 3644 -15418 4604 -15380
rect 4662 -15380 4887 -15363
rect 4921 -15380 4955 -15346
rect 4989 -15380 5023 -15346
rect 5057 -15380 5091 -15346
rect 5125 -15380 5159 -15346
rect 5193 -15380 5227 -15346
rect 5261 -15380 5295 -15346
rect 5329 -15380 5363 -15346
rect 5397 -15363 5436 -15346
rect 5866 -15346 6454 -15330
rect 5866 -15363 5905 -15346
rect 5397 -15380 5622 -15363
rect 4662 -15418 5622 -15380
rect 5680 -15380 5905 -15363
rect 5939 -15380 5973 -15346
rect 6007 -15380 6041 -15346
rect 6075 -15380 6109 -15346
rect 6143 -15380 6177 -15346
rect 6211 -15380 6245 -15346
rect 6279 -15380 6313 -15346
rect 6347 -15380 6381 -15346
rect 6415 -15363 6454 -15346
rect 6884 -15346 7472 -15330
rect 6884 -15363 6923 -15346
rect 6415 -15380 6640 -15363
rect 5680 -15418 6640 -15380
rect 6698 -15380 6923 -15363
rect 6957 -15380 6991 -15346
rect 7025 -15380 7059 -15346
rect 7093 -15380 7127 -15346
rect 7161 -15380 7195 -15346
rect 7229 -15380 7263 -15346
rect 7297 -15380 7331 -15346
rect 7365 -15380 7399 -15346
rect 7433 -15363 7472 -15346
rect 7902 -15346 8490 -15330
rect 7902 -15363 7941 -15346
rect 7433 -15380 7658 -15363
rect 6698 -15418 7658 -15380
rect 7716 -15380 7941 -15363
rect 7975 -15380 8009 -15346
rect 8043 -15380 8077 -15346
rect 8111 -15380 8145 -15346
rect 8179 -15380 8213 -15346
rect 8247 -15380 8281 -15346
rect 8315 -15380 8349 -15346
rect 8383 -15380 8417 -15346
rect 8451 -15363 8490 -15346
rect 8920 -15346 9508 -15330
rect 8920 -15363 8959 -15346
rect 8451 -15380 8676 -15363
rect 7716 -15418 8676 -15380
rect 8734 -15380 8959 -15363
rect 8993 -15380 9027 -15346
rect 9061 -15380 9095 -15346
rect 9129 -15380 9163 -15346
rect 9197 -15380 9231 -15346
rect 9265 -15380 9299 -15346
rect 9333 -15380 9367 -15346
rect 9401 -15380 9435 -15346
rect 9469 -15363 9508 -15346
rect 9938 -15346 10526 -15330
rect 9938 -15363 9977 -15346
rect 9469 -15380 9694 -15363
rect 8734 -15418 9694 -15380
rect 9752 -15380 9977 -15363
rect 10011 -15380 10045 -15346
rect 10079 -15380 10113 -15346
rect 10147 -15380 10181 -15346
rect 10215 -15380 10249 -15346
rect 10283 -15380 10317 -15346
rect 10351 -15380 10385 -15346
rect 10419 -15380 10453 -15346
rect 10487 -15363 10526 -15346
rect 10956 -15346 11544 -15330
rect 10956 -15363 10995 -15346
rect 10487 -15380 10712 -15363
rect 9752 -15418 10712 -15380
rect 10770 -15380 10995 -15363
rect 11029 -15380 11063 -15346
rect 11097 -15380 11131 -15346
rect 11165 -15380 11199 -15346
rect 11233 -15380 11267 -15346
rect 11301 -15380 11335 -15346
rect 11369 -15380 11403 -15346
rect 11437 -15380 11471 -15346
rect 11505 -15363 11544 -15346
rect 11974 -15346 12562 -15330
rect 11974 -15363 12013 -15346
rect 11505 -15380 11730 -15363
rect 10770 -15418 11730 -15380
rect 11788 -15380 12013 -15363
rect 12047 -15380 12081 -15346
rect 12115 -15380 12149 -15346
rect 12183 -15380 12217 -15346
rect 12251 -15380 12285 -15346
rect 12319 -15380 12353 -15346
rect 12387 -15380 12421 -15346
rect 12455 -15380 12489 -15346
rect 12523 -15363 12562 -15346
rect 12992 -15346 13580 -15330
rect 12992 -15363 13031 -15346
rect 12523 -15380 12748 -15363
rect 11788 -15418 12748 -15380
rect 12806 -15380 13031 -15363
rect 13065 -15380 13099 -15346
rect 13133 -15380 13167 -15346
rect 13201 -15380 13235 -15346
rect 13269 -15380 13303 -15346
rect 13337 -15380 13371 -15346
rect 13405 -15380 13439 -15346
rect 13473 -15380 13507 -15346
rect 13541 -15363 13580 -15346
rect 14010 -15346 14598 -15330
rect 14010 -15363 14049 -15346
rect 13541 -15380 13766 -15363
rect 12806 -15418 13766 -15380
rect 13824 -15380 14049 -15363
rect 14083 -15380 14117 -15346
rect 14151 -15380 14185 -15346
rect 14219 -15380 14253 -15346
rect 14287 -15380 14321 -15346
rect 14355 -15380 14389 -15346
rect 14423 -15380 14457 -15346
rect 14491 -15380 14525 -15346
rect 14559 -15363 14598 -15346
rect 15028 -15346 15616 -15330
rect 15028 -15363 15067 -15346
rect 14559 -15380 14784 -15363
rect 13824 -15418 14784 -15380
rect 14842 -15380 15067 -15363
rect 15101 -15380 15135 -15346
rect 15169 -15380 15203 -15346
rect 15237 -15380 15271 -15346
rect 15305 -15380 15339 -15346
rect 15373 -15380 15407 -15346
rect 15441 -15380 15475 -15346
rect 15509 -15380 15543 -15346
rect 15577 -15363 15616 -15346
rect 16046 -15346 16634 -15330
rect 16046 -15363 16085 -15346
rect 15577 -15380 15802 -15363
rect 14842 -15418 15802 -15380
rect 15860 -15380 16085 -15363
rect 16119 -15380 16153 -15346
rect 16187 -15380 16221 -15346
rect 16255 -15380 16289 -15346
rect 16323 -15380 16357 -15346
rect 16391 -15380 16425 -15346
rect 16459 -15380 16493 -15346
rect 16527 -15380 16561 -15346
rect 16595 -15363 16634 -15346
rect 17064 -15346 17652 -15330
rect 17064 -15363 17103 -15346
rect 16595 -15380 16820 -15363
rect 15860 -15418 16820 -15380
rect 16878 -15380 17103 -15363
rect 17137 -15380 17171 -15346
rect 17205 -15380 17239 -15346
rect 17273 -15380 17307 -15346
rect 17341 -15380 17375 -15346
rect 17409 -15380 17443 -15346
rect 17477 -15380 17511 -15346
rect 17545 -15380 17579 -15346
rect 17613 -15363 17652 -15346
rect 18082 -15346 18670 -15330
rect 18082 -15363 18121 -15346
rect 17613 -15380 17838 -15363
rect 16878 -15418 17838 -15380
rect 17896 -15380 18121 -15363
rect 18155 -15380 18189 -15346
rect 18223 -15380 18257 -15346
rect 18291 -15380 18325 -15346
rect 18359 -15380 18393 -15346
rect 18427 -15380 18461 -15346
rect 18495 -15380 18529 -15346
rect 18563 -15380 18597 -15346
rect 18631 -15363 18670 -15346
rect 19100 -15346 19688 -15330
rect 19100 -15363 19139 -15346
rect 18631 -15380 18856 -15363
rect 17896 -15418 18856 -15380
rect 18914 -15380 19139 -15363
rect 19173 -15380 19207 -15346
rect 19241 -15380 19275 -15346
rect 19309 -15380 19343 -15346
rect 19377 -15380 19411 -15346
rect 19445 -15380 19479 -15346
rect 19513 -15380 19547 -15346
rect 19581 -15380 19615 -15346
rect 19649 -15363 19688 -15346
rect 20118 -15346 20706 -15330
rect 20118 -15363 20157 -15346
rect 19649 -15380 19874 -15363
rect 18914 -15418 19874 -15380
rect 19932 -15380 20157 -15363
rect 20191 -15380 20225 -15346
rect 20259 -15380 20293 -15346
rect 20327 -15380 20361 -15346
rect 20395 -15380 20429 -15346
rect 20463 -15380 20497 -15346
rect 20531 -15380 20565 -15346
rect 20599 -15380 20633 -15346
rect 20667 -15363 20706 -15346
rect 21136 -15346 21724 -15330
rect 21136 -15363 21175 -15346
rect 20667 -15380 20892 -15363
rect 19932 -15418 20892 -15380
rect 20950 -15380 21175 -15363
rect 21209 -15380 21243 -15346
rect 21277 -15380 21311 -15346
rect 21345 -15380 21379 -15346
rect 21413 -15380 21447 -15346
rect 21481 -15380 21515 -15346
rect 21549 -15380 21583 -15346
rect 21617 -15380 21651 -15346
rect 21685 -15363 21724 -15346
rect 22154 -15346 22742 -15330
rect 22154 -15363 22193 -15346
rect 21685 -15380 21910 -15363
rect 20950 -15418 21910 -15380
rect 21968 -15380 22193 -15363
rect 22227 -15380 22261 -15346
rect 22295 -15380 22329 -15346
rect 22363 -15380 22397 -15346
rect 22431 -15380 22465 -15346
rect 22499 -15380 22533 -15346
rect 22567 -15380 22601 -15346
rect 22635 -15380 22669 -15346
rect 22703 -15363 22742 -15346
rect 22703 -15380 22928 -15363
rect 21968 -15418 22928 -15380
rect -9138 -15604 -8178 -15566
rect -9138 -15621 -8913 -15604
rect -8952 -15638 -8913 -15621
rect -8879 -15638 -8845 -15604
rect -8811 -15638 -8777 -15604
rect -8743 -15638 -8709 -15604
rect -8675 -15638 -8641 -15604
rect -8607 -15638 -8573 -15604
rect -8539 -15638 -8505 -15604
rect -8471 -15638 -8437 -15604
rect -8403 -15621 -8178 -15604
rect -8120 -15604 -7160 -15566
rect -8120 -15621 -7895 -15604
rect -8403 -15638 -8364 -15621
rect -8952 -15654 -8364 -15638
rect -7934 -15638 -7895 -15621
rect -7861 -15638 -7827 -15604
rect -7793 -15638 -7759 -15604
rect -7725 -15638 -7691 -15604
rect -7657 -15638 -7623 -15604
rect -7589 -15638 -7555 -15604
rect -7521 -15638 -7487 -15604
rect -7453 -15638 -7419 -15604
rect -7385 -15621 -7160 -15604
rect -7102 -15604 -6142 -15566
rect -7102 -15621 -6877 -15604
rect -7385 -15638 -7346 -15621
rect -7934 -15654 -7346 -15638
rect -6916 -15638 -6877 -15621
rect -6843 -15638 -6809 -15604
rect -6775 -15638 -6741 -15604
rect -6707 -15638 -6673 -15604
rect -6639 -15638 -6605 -15604
rect -6571 -15638 -6537 -15604
rect -6503 -15638 -6469 -15604
rect -6435 -15638 -6401 -15604
rect -6367 -15621 -6142 -15604
rect -6084 -15604 -5124 -15566
rect -6084 -15621 -5859 -15604
rect -6367 -15638 -6328 -15621
rect -6916 -15654 -6328 -15638
rect -5898 -15638 -5859 -15621
rect -5825 -15638 -5791 -15604
rect -5757 -15638 -5723 -15604
rect -5689 -15638 -5655 -15604
rect -5621 -15638 -5587 -15604
rect -5553 -15638 -5519 -15604
rect -5485 -15638 -5451 -15604
rect -5417 -15638 -5383 -15604
rect -5349 -15621 -5124 -15604
rect -5066 -15604 -4106 -15566
rect -5066 -15621 -4841 -15604
rect -5349 -15638 -5310 -15621
rect -5898 -15654 -5310 -15638
rect -4880 -15638 -4841 -15621
rect -4807 -15638 -4773 -15604
rect -4739 -15638 -4705 -15604
rect -4671 -15638 -4637 -15604
rect -4603 -15638 -4569 -15604
rect -4535 -15638 -4501 -15604
rect -4467 -15638 -4433 -15604
rect -4399 -15638 -4365 -15604
rect -4331 -15621 -4106 -15604
rect -4048 -15604 -3088 -15566
rect -4048 -15621 -3823 -15604
rect -4331 -15638 -4292 -15621
rect -4880 -15654 -4292 -15638
rect -3862 -15638 -3823 -15621
rect -3789 -15638 -3755 -15604
rect -3721 -15638 -3687 -15604
rect -3653 -15638 -3619 -15604
rect -3585 -15638 -3551 -15604
rect -3517 -15638 -3483 -15604
rect -3449 -15638 -3415 -15604
rect -3381 -15638 -3347 -15604
rect -3313 -15621 -3088 -15604
rect -3030 -15604 -2070 -15566
rect -3030 -15621 -2805 -15604
rect -3313 -15638 -3274 -15621
rect -3862 -15654 -3274 -15638
rect -2844 -15638 -2805 -15621
rect -2771 -15638 -2737 -15604
rect -2703 -15638 -2669 -15604
rect -2635 -15638 -2601 -15604
rect -2567 -15638 -2533 -15604
rect -2499 -15638 -2465 -15604
rect -2431 -15638 -2397 -15604
rect -2363 -15638 -2329 -15604
rect -2295 -15621 -2070 -15604
rect -2012 -15604 -1052 -15566
rect -2012 -15621 -1787 -15604
rect -2295 -15638 -2256 -15621
rect -2844 -15654 -2256 -15638
rect -1826 -15638 -1787 -15621
rect -1753 -15638 -1719 -15604
rect -1685 -15638 -1651 -15604
rect -1617 -15638 -1583 -15604
rect -1549 -15638 -1515 -15604
rect -1481 -15638 -1447 -15604
rect -1413 -15638 -1379 -15604
rect -1345 -15638 -1311 -15604
rect -1277 -15621 -1052 -15604
rect -994 -15604 -34 -15566
rect -994 -15621 -769 -15604
rect -1277 -15638 -1238 -15621
rect -1826 -15654 -1238 -15638
rect -808 -15638 -769 -15621
rect -735 -15638 -701 -15604
rect -667 -15638 -633 -15604
rect -599 -15638 -565 -15604
rect -531 -15638 -497 -15604
rect -463 -15638 -429 -15604
rect -395 -15638 -361 -15604
rect -327 -15638 -293 -15604
rect -259 -15621 -34 -15604
rect -259 -15638 -220 -15621
rect -808 -15654 -220 -15638
rect -8952 -15712 -8364 -15696
rect -8952 -15729 -8913 -15712
rect -9138 -15746 -8913 -15729
rect -8879 -15746 -8845 -15712
rect -8811 -15746 -8777 -15712
rect -8743 -15746 -8709 -15712
rect -8675 -15746 -8641 -15712
rect -8607 -15746 -8573 -15712
rect -8539 -15746 -8505 -15712
rect -8471 -15746 -8437 -15712
rect -8403 -15729 -8364 -15712
rect -7934 -15712 -7346 -15696
rect -7934 -15729 -7895 -15712
rect -8403 -15746 -8178 -15729
rect -9138 -15784 -8178 -15746
rect -8120 -15746 -7895 -15729
rect -7861 -15746 -7827 -15712
rect -7793 -15746 -7759 -15712
rect -7725 -15746 -7691 -15712
rect -7657 -15746 -7623 -15712
rect -7589 -15746 -7555 -15712
rect -7521 -15746 -7487 -15712
rect -7453 -15746 -7419 -15712
rect -7385 -15729 -7346 -15712
rect -6916 -15712 -6328 -15696
rect -6916 -15729 -6877 -15712
rect -7385 -15746 -7160 -15729
rect -8120 -15784 -7160 -15746
rect -7102 -15746 -6877 -15729
rect -6843 -15746 -6809 -15712
rect -6775 -15746 -6741 -15712
rect -6707 -15746 -6673 -15712
rect -6639 -15746 -6605 -15712
rect -6571 -15746 -6537 -15712
rect -6503 -15746 -6469 -15712
rect -6435 -15746 -6401 -15712
rect -6367 -15729 -6328 -15712
rect -5898 -15712 -5310 -15696
rect -5898 -15729 -5859 -15712
rect -6367 -15746 -6142 -15729
rect -7102 -15784 -6142 -15746
rect -6084 -15746 -5859 -15729
rect -5825 -15746 -5791 -15712
rect -5757 -15746 -5723 -15712
rect -5689 -15746 -5655 -15712
rect -5621 -15746 -5587 -15712
rect -5553 -15746 -5519 -15712
rect -5485 -15746 -5451 -15712
rect -5417 -15746 -5383 -15712
rect -5349 -15729 -5310 -15712
rect -4880 -15712 -4292 -15696
rect -4880 -15729 -4841 -15712
rect -5349 -15746 -5124 -15729
rect -6084 -15784 -5124 -15746
rect -5066 -15746 -4841 -15729
rect -4807 -15746 -4773 -15712
rect -4739 -15746 -4705 -15712
rect -4671 -15746 -4637 -15712
rect -4603 -15746 -4569 -15712
rect -4535 -15746 -4501 -15712
rect -4467 -15746 -4433 -15712
rect -4399 -15746 -4365 -15712
rect -4331 -15729 -4292 -15712
rect -3862 -15712 -3274 -15696
rect -3862 -15729 -3823 -15712
rect -4331 -15746 -4106 -15729
rect -5066 -15784 -4106 -15746
rect -4048 -15746 -3823 -15729
rect -3789 -15746 -3755 -15712
rect -3721 -15746 -3687 -15712
rect -3653 -15746 -3619 -15712
rect -3585 -15746 -3551 -15712
rect -3517 -15746 -3483 -15712
rect -3449 -15746 -3415 -15712
rect -3381 -15746 -3347 -15712
rect -3313 -15729 -3274 -15712
rect -2844 -15712 -2256 -15696
rect -2844 -15729 -2805 -15712
rect -3313 -15746 -3088 -15729
rect -4048 -15784 -3088 -15746
rect -3030 -15746 -2805 -15729
rect -2771 -15746 -2737 -15712
rect -2703 -15746 -2669 -15712
rect -2635 -15746 -2601 -15712
rect -2567 -15746 -2533 -15712
rect -2499 -15746 -2465 -15712
rect -2431 -15746 -2397 -15712
rect -2363 -15746 -2329 -15712
rect -2295 -15729 -2256 -15712
rect -1826 -15712 -1238 -15696
rect -1826 -15729 -1787 -15712
rect -2295 -15746 -2070 -15729
rect -3030 -15784 -2070 -15746
rect -2012 -15746 -1787 -15729
rect -1753 -15746 -1719 -15712
rect -1685 -15746 -1651 -15712
rect -1617 -15746 -1583 -15712
rect -1549 -15746 -1515 -15712
rect -1481 -15746 -1447 -15712
rect -1413 -15746 -1379 -15712
rect -1345 -15746 -1311 -15712
rect -1277 -15729 -1238 -15712
rect -808 -15712 -220 -15696
rect -808 -15729 -769 -15712
rect -1277 -15746 -1052 -15729
rect -2012 -15784 -1052 -15746
rect -994 -15746 -769 -15729
rect -735 -15746 -701 -15712
rect -667 -15746 -633 -15712
rect -599 -15746 -565 -15712
rect -531 -15746 -497 -15712
rect -463 -15746 -429 -15712
rect -395 -15746 -361 -15712
rect -327 -15746 -293 -15712
rect -259 -15729 -220 -15712
rect -259 -15746 -34 -15729
rect -994 -15784 -34 -15746
rect 2626 -16056 3586 -16018
rect 2626 -16073 2851 -16056
rect 2812 -16090 2851 -16073
rect 2885 -16090 2919 -16056
rect 2953 -16090 2987 -16056
rect 3021 -16090 3055 -16056
rect 3089 -16090 3123 -16056
rect 3157 -16090 3191 -16056
rect 3225 -16090 3259 -16056
rect 3293 -16090 3327 -16056
rect 3361 -16073 3586 -16056
rect 3644 -16056 4604 -16018
rect 3644 -16073 3869 -16056
rect 3361 -16090 3400 -16073
rect 2812 -16106 3400 -16090
rect 3830 -16090 3869 -16073
rect 3903 -16090 3937 -16056
rect 3971 -16090 4005 -16056
rect 4039 -16090 4073 -16056
rect 4107 -16090 4141 -16056
rect 4175 -16090 4209 -16056
rect 4243 -16090 4277 -16056
rect 4311 -16090 4345 -16056
rect 4379 -16073 4604 -16056
rect 4662 -16056 5622 -16018
rect 4662 -16073 4887 -16056
rect 4379 -16090 4418 -16073
rect 3830 -16106 4418 -16090
rect 4848 -16090 4887 -16073
rect 4921 -16090 4955 -16056
rect 4989 -16090 5023 -16056
rect 5057 -16090 5091 -16056
rect 5125 -16090 5159 -16056
rect 5193 -16090 5227 -16056
rect 5261 -16090 5295 -16056
rect 5329 -16090 5363 -16056
rect 5397 -16073 5622 -16056
rect 5680 -16056 6640 -16018
rect 5680 -16073 5905 -16056
rect 5397 -16090 5436 -16073
rect 4848 -16106 5436 -16090
rect 5866 -16090 5905 -16073
rect 5939 -16090 5973 -16056
rect 6007 -16090 6041 -16056
rect 6075 -16090 6109 -16056
rect 6143 -16090 6177 -16056
rect 6211 -16090 6245 -16056
rect 6279 -16090 6313 -16056
rect 6347 -16090 6381 -16056
rect 6415 -16073 6640 -16056
rect 6698 -16056 7658 -16018
rect 6698 -16073 6923 -16056
rect 6415 -16090 6454 -16073
rect 5866 -16106 6454 -16090
rect 6884 -16090 6923 -16073
rect 6957 -16090 6991 -16056
rect 7025 -16090 7059 -16056
rect 7093 -16090 7127 -16056
rect 7161 -16090 7195 -16056
rect 7229 -16090 7263 -16056
rect 7297 -16090 7331 -16056
rect 7365 -16090 7399 -16056
rect 7433 -16073 7658 -16056
rect 7716 -16056 8676 -16018
rect 7716 -16073 7941 -16056
rect 7433 -16090 7472 -16073
rect 6884 -16106 7472 -16090
rect 7902 -16090 7941 -16073
rect 7975 -16090 8009 -16056
rect 8043 -16090 8077 -16056
rect 8111 -16090 8145 -16056
rect 8179 -16090 8213 -16056
rect 8247 -16090 8281 -16056
rect 8315 -16090 8349 -16056
rect 8383 -16090 8417 -16056
rect 8451 -16073 8676 -16056
rect 8734 -16056 9694 -16018
rect 8734 -16073 8959 -16056
rect 8451 -16090 8490 -16073
rect 7902 -16106 8490 -16090
rect 8920 -16090 8959 -16073
rect 8993 -16090 9027 -16056
rect 9061 -16090 9095 -16056
rect 9129 -16090 9163 -16056
rect 9197 -16090 9231 -16056
rect 9265 -16090 9299 -16056
rect 9333 -16090 9367 -16056
rect 9401 -16090 9435 -16056
rect 9469 -16073 9694 -16056
rect 9752 -16056 10712 -16018
rect 9752 -16073 9977 -16056
rect 9469 -16090 9508 -16073
rect 8920 -16106 9508 -16090
rect 9938 -16090 9977 -16073
rect 10011 -16090 10045 -16056
rect 10079 -16090 10113 -16056
rect 10147 -16090 10181 -16056
rect 10215 -16090 10249 -16056
rect 10283 -16090 10317 -16056
rect 10351 -16090 10385 -16056
rect 10419 -16090 10453 -16056
rect 10487 -16073 10712 -16056
rect 10770 -16056 11730 -16018
rect 10770 -16073 10995 -16056
rect 10487 -16090 10526 -16073
rect 9938 -16106 10526 -16090
rect 10956 -16090 10995 -16073
rect 11029 -16090 11063 -16056
rect 11097 -16090 11131 -16056
rect 11165 -16090 11199 -16056
rect 11233 -16090 11267 -16056
rect 11301 -16090 11335 -16056
rect 11369 -16090 11403 -16056
rect 11437 -16090 11471 -16056
rect 11505 -16073 11730 -16056
rect 11788 -16056 12748 -16018
rect 11788 -16073 12013 -16056
rect 11505 -16090 11544 -16073
rect 10956 -16106 11544 -16090
rect 11974 -16090 12013 -16073
rect 12047 -16090 12081 -16056
rect 12115 -16090 12149 -16056
rect 12183 -16090 12217 -16056
rect 12251 -16090 12285 -16056
rect 12319 -16090 12353 -16056
rect 12387 -16090 12421 -16056
rect 12455 -16090 12489 -16056
rect 12523 -16073 12748 -16056
rect 12806 -16056 13766 -16018
rect 12806 -16073 13031 -16056
rect 12523 -16090 12562 -16073
rect 11974 -16106 12562 -16090
rect 12992 -16090 13031 -16073
rect 13065 -16090 13099 -16056
rect 13133 -16090 13167 -16056
rect 13201 -16090 13235 -16056
rect 13269 -16090 13303 -16056
rect 13337 -16090 13371 -16056
rect 13405 -16090 13439 -16056
rect 13473 -16090 13507 -16056
rect 13541 -16073 13766 -16056
rect 13824 -16056 14784 -16018
rect 13824 -16073 14049 -16056
rect 13541 -16090 13580 -16073
rect 12992 -16106 13580 -16090
rect 14010 -16090 14049 -16073
rect 14083 -16090 14117 -16056
rect 14151 -16090 14185 -16056
rect 14219 -16090 14253 -16056
rect 14287 -16090 14321 -16056
rect 14355 -16090 14389 -16056
rect 14423 -16090 14457 -16056
rect 14491 -16090 14525 -16056
rect 14559 -16073 14784 -16056
rect 14842 -16056 15802 -16018
rect 14842 -16073 15067 -16056
rect 14559 -16090 14598 -16073
rect 14010 -16106 14598 -16090
rect 15028 -16090 15067 -16073
rect 15101 -16090 15135 -16056
rect 15169 -16090 15203 -16056
rect 15237 -16090 15271 -16056
rect 15305 -16090 15339 -16056
rect 15373 -16090 15407 -16056
rect 15441 -16090 15475 -16056
rect 15509 -16090 15543 -16056
rect 15577 -16073 15802 -16056
rect 15860 -16056 16820 -16018
rect 15860 -16073 16085 -16056
rect 15577 -16090 15616 -16073
rect 15028 -16106 15616 -16090
rect 16046 -16090 16085 -16073
rect 16119 -16090 16153 -16056
rect 16187 -16090 16221 -16056
rect 16255 -16090 16289 -16056
rect 16323 -16090 16357 -16056
rect 16391 -16090 16425 -16056
rect 16459 -16090 16493 -16056
rect 16527 -16090 16561 -16056
rect 16595 -16073 16820 -16056
rect 16878 -16056 17838 -16018
rect 16878 -16073 17103 -16056
rect 16595 -16090 16634 -16073
rect 16046 -16106 16634 -16090
rect 17064 -16090 17103 -16073
rect 17137 -16090 17171 -16056
rect 17205 -16090 17239 -16056
rect 17273 -16090 17307 -16056
rect 17341 -16090 17375 -16056
rect 17409 -16090 17443 -16056
rect 17477 -16090 17511 -16056
rect 17545 -16090 17579 -16056
rect 17613 -16073 17838 -16056
rect 17896 -16056 18856 -16018
rect 17896 -16073 18121 -16056
rect 17613 -16090 17652 -16073
rect 17064 -16106 17652 -16090
rect 18082 -16090 18121 -16073
rect 18155 -16090 18189 -16056
rect 18223 -16090 18257 -16056
rect 18291 -16090 18325 -16056
rect 18359 -16090 18393 -16056
rect 18427 -16090 18461 -16056
rect 18495 -16090 18529 -16056
rect 18563 -16090 18597 -16056
rect 18631 -16073 18856 -16056
rect 18914 -16056 19874 -16018
rect 18914 -16073 19139 -16056
rect 18631 -16090 18670 -16073
rect 18082 -16106 18670 -16090
rect 19100 -16090 19139 -16073
rect 19173 -16090 19207 -16056
rect 19241 -16090 19275 -16056
rect 19309 -16090 19343 -16056
rect 19377 -16090 19411 -16056
rect 19445 -16090 19479 -16056
rect 19513 -16090 19547 -16056
rect 19581 -16090 19615 -16056
rect 19649 -16073 19874 -16056
rect 19932 -16056 20892 -16018
rect 19932 -16073 20157 -16056
rect 19649 -16090 19688 -16073
rect 19100 -16106 19688 -16090
rect 20118 -16090 20157 -16073
rect 20191 -16090 20225 -16056
rect 20259 -16090 20293 -16056
rect 20327 -16090 20361 -16056
rect 20395 -16090 20429 -16056
rect 20463 -16090 20497 -16056
rect 20531 -16090 20565 -16056
rect 20599 -16090 20633 -16056
rect 20667 -16073 20892 -16056
rect 20950 -16056 21910 -16018
rect 20950 -16073 21175 -16056
rect 20667 -16090 20706 -16073
rect 20118 -16106 20706 -16090
rect 21136 -16090 21175 -16073
rect 21209 -16090 21243 -16056
rect 21277 -16090 21311 -16056
rect 21345 -16090 21379 -16056
rect 21413 -16090 21447 -16056
rect 21481 -16090 21515 -16056
rect 21549 -16090 21583 -16056
rect 21617 -16090 21651 -16056
rect 21685 -16073 21910 -16056
rect 21968 -16056 22928 -16018
rect 21968 -16073 22193 -16056
rect 21685 -16090 21724 -16073
rect 21136 -16106 21724 -16090
rect 22154 -16090 22193 -16073
rect 22227 -16090 22261 -16056
rect 22295 -16090 22329 -16056
rect 22363 -16090 22397 -16056
rect 22431 -16090 22465 -16056
rect 22499 -16090 22533 -16056
rect 22567 -16090 22601 -16056
rect 22635 -16090 22669 -16056
rect 22703 -16073 22928 -16056
rect 22703 -16090 22742 -16073
rect 22154 -16106 22742 -16090
rect -9138 -16422 -8178 -16384
rect -9138 -16439 -8913 -16422
rect -8952 -16456 -8913 -16439
rect -8879 -16456 -8845 -16422
rect -8811 -16456 -8777 -16422
rect -8743 -16456 -8709 -16422
rect -8675 -16456 -8641 -16422
rect -8607 -16456 -8573 -16422
rect -8539 -16456 -8505 -16422
rect -8471 -16456 -8437 -16422
rect -8403 -16439 -8178 -16422
rect -8120 -16422 -7160 -16384
rect -8120 -16439 -7895 -16422
rect -8403 -16456 -8364 -16439
rect -8952 -16472 -8364 -16456
rect -7934 -16456 -7895 -16439
rect -7861 -16456 -7827 -16422
rect -7793 -16456 -7759 -16422
rect -7725 -16456 -7691 -16422
rect -7657 -16456 -7623 -16422
rect -7589 -16456 -7555 -16422
rect -7521 -16456 -7487 -16422
rect -7453 -16456 -7419 -16422
rect -7385 -16439 -7160 -16422
rect -7102 -16422 -6142 -16384
rect -7102 -16439 -6877 -16422
rect -7385 -16456 -7346 -16439
rect -7934 -16472 -7346 -16456
rect -6916 -16456 -6877 -16439
rect -6843 -16456 -6809 -16422
rect -6775 -16456 -6741 -16422
rect -6707 -16456 -6673 -16422
rect -6639 -16456 -6605 -16422
rect -6571 -16456 -6537 -16422
rect -6503 -16456 -6469 -16422
rect -6435 -16456 -6401 -16422
rect -6367 -16439 -6142 -16422
rect -6084 -16422 -5124 -16384
rect -6084 -16439 -5859 -16422
rect -6367 -16456 -6328 -16439
rect -6916 -16472 -6328 -16456
rect -5898 -16456 -5859 -16439
rect -5825 -16456 -5791 -16422
rect -5757 -16456 -5723 -16422
rect -5689 -16456 -5655 -16422
rect -5621 -16456 -5587 -16422
rect -5553 -16456 -5519 -16422
rect -5485 -16456 -5451 -16422
rect -5417 -16456 -5383 -16422
rect -5349 -16439 -5124 -16422
rect -5066 -16422 -4106 -16384
rect -5066 -16439 -4841 -16422
rect -5349 -16456 -5310 -16439
rect -5898 -16472 -5310 -16456
rect -4880 -16456 -4841 -16439
rect -4807 -16456 -4773 -16422
rect -4739 -16456 -4705 -16422
rect -4671 -16456 -4637 -16422
rect -4603 -16456 -4569 -16422
rect -4535 -16456 -4501 -16422
rect -4467 -16456 -4433 -16422
rect -4399 -16456 -4365 -16422
rect -4331 -16439 -4106 -16422
rect -4048 -16422 -3088 -16384
rect -4048 -16439 -3823 -16422
rect -4331 -16456 -4292 -16439
rect -4880 -16472 -4292 -16456
rect -3862 -16456 -3823 -16439
rect -3789 -16456 -3755 -16422
rect -3721 -16456 -3687 -16422
rect -3653 -16456 -3619 -16422
rect -3585 -16456 -3551 -16422
rect -3517 -16456 -3483 -16422
rect -3449 -16456 -3415 -16422
rect -3381 -16456 -3347 -16422
rect -3313 -16439 -3088 -16422
rect -3030 -16422 -2070 -16384
rect -3030 -16439 -2805 -16422
rect -3313 -16456 -3274 -16439
rect -3862 -16472 -3274 -16456
rect -2844 -16456 -2805 -16439
rect -2771 -16456 -2737 -16422
rect -2703 -16456 -2669 -16422
rect -2635 -16456 -2601 -16422
rect -2567 -16456 -2533 -16422
rect -2499 -16456 -2465 -16422
rect -2431 -16456 -2397 -16422
rect -2363 -16456 -2329 -16422
rect -2295 -16439 -2070 -16422
rect -2012 -16422 -1052 -16384
rect -2012 -16439 -1787 -16422
rect -2295 -16456 -2256 -16439
rect -2844 -16472 -2256 -16456
rect -1826 -16456 -1787 -16439
rect -1753 -16456 -1719 -16422
rect -1685 -16456 -1651 -16422
rect -1617 -16456 -1583 -16422
rect -1549 -16456 -1515 -16422
rect -1481 -16456 -1447 -16422
rect -1413 -16456 -1379 -16422
rect -1345 -16456 -1311 -16422
rect -1277 -16439 -1052 -16422
rect -994 -16422 -34 -16384
rect -994 -16439 -769 -16422
rect -1277 -16456 -1238 -16439
rect -1826 -16472 -1238 -16456
rect -808 -16456 -769 -16439
rect -735 -16456 -701 -16422
rect -667 -16456 -633 -16422
rect -599 -16456 -565 -16422
rect -531 -16456 -497 -16422
rect -463 -16456 -429 -16422
rect -395 -16456 -361 -16422
rect -327 -16456 -293 -16422
rect -259 -16439 -34 -16422
rect -259 -16456 -220 -16439
rect -808 -16472 -220 -16456
rect -8952 -16530 -8364 -16514
rect -8952 -16547 -8913 -16530
rect -9138 -16564 -8913 -16547
rect -8879 -16564 -8845 -16530
rect -8811 -16564 -8777 -16530
rect -8743 -16564 -8709 -16530
rect -8675 -16564 -8641 -16530
rect -8607 -16564 -8573 -16530
rect -8539 -16564 -8505 -16530
rect -8471 -16564 -8437 -16530
rect -8403 -16547 -8364 -16530
rect -7934 -16530 -7346 -16514
rect -7934 -16547 -7895 -16530
rect -8403 -16564 -8178 -16547
rect -9138 -16602 -8178 -16564
rect -8120 -16564 -7895 -16547
rect -7861 -16564 -7827 -16530
rect -7793 -16564 -7759 -16530
rect -7725 -16564 -7691 -16530
rect -7657 -16564 -7623 -16530
rect -7589 -16564 -7555 -16530
rect -7521 -16564 -7487 -16530
rect -7453 -16564 -7419 -16530
rect -7385 -16547 -7346 -16530
rect -6916 -16530 -6328 -16514
rect -6916 -16547 -6877 -16530
rect -7385 -16564 -7160 -16547
rect -8120 -16602 -7160 -16564
rect -7102 -16564 -6877 -16547
rect -6843 -16564 -6809 -16530
rect -6775 -16564 -6741 -16530
rect -6707 -16564 -6673 -16530
rect -6639 -16564 -6605 -16530
rect -6571 -16564 -6537 -16530
rect -6503 -16564 -6469 -16530
rect -6435 -16564 -6401 -16530
rect -6367 -16547 -6328 -16530
rect -5898 -16530 -5310 -16514
rect -5898 -16547 -5859 -16530
rect -6367 -16564 -6142 -16547
rect -7102 -16602 -6142 -16564
rect -6084 -16564 -5859 -16547
rect -5825 -16564 -5791 -16530
rect -5757 -16564 -5723 -16530
rect -5689 -16564 -5655 -16530
rect -5621 -16564 -5587 -16530
rect -5553 -16564 -5519 -16530
rect -5485 -16564 -5451 -16530
rect -5417 -16564 -5383 -16530
rect -5349 -16547 -5310 -16530
rect -4880 -16530 -4292 -16514
rect -4880 -16547 -4841 -16530
rect -5349 -16564 -5124 -16547
rect -6084 -16602 -5124 -16564
rect -5066 -16564 -4841 -16547
rect -4807 -16564 -4773 -16530
rect -4739 -16564 -4705 -16530
rect -4671 -16564 -4637 -16530
rect -4603 -16564 -4569 -16530
rect -4535 -16564 -4501 -16530
rect -4467 -16564 -4433 -16530
rect -4399 -16564 -4365 -16530
rect -4331 -16547 -4292 -16530
rect -3862 -16530 -3274 -16514
rect -3862 -16547 -3823 -16530
rect -4331 -16564 -4106 -16547
rect -5066 -16602 -4106 -16564
rect -4048 -16564 -3823 -16547
rect -3789 -16564 -3755 -16530
rect -3721 -16564 -3687 -16530
rect -3653 -16564 -3619 -16530
rect -3585 -16564 -3551 -16530
rect -3517 -16564 -3483 -16530
rect -3449 -16564 -3415 -16530
rect -3381 -16564 -3347 -16530
rect -3313 -16547 -3274 -16530
rect -2844 -16530 -2256 -16514
rect -2844 -16547 -2805 -16530
rect -3313 -16564 -3088 -16547
rect -4048 -16602 -3088 -16564
rect -3030 -16564 -2805 -16547
rect -2771 -16564 -2737 -16530
rect -2703 -16564 -2669 -16530
rect -2635 -16564 -2601 -16530
rect -2567 -16564 -2533 -16530
rect -2499 -16564 -2465 -16530
rect -2431 -16564 -2397 -16530
rect -2363 -16564 -2329 -16530
rect -2295 -16547 -2256 -16530
rect -1826 -16530 -1238 -16514
rect -1826 -16547 -1787 -16530
rect -2295 -16564 -2070 -16547
rect -3030 -16602 -2070 -16564
rect -2012 -16564 -1787 -16547
rect -1753 -16564 -1719 -16530
rect -1685 -16564 -1651 -16530
rect -1617 -16564 -1583 -16530
rect -1549 -16564 -1515 -16530
rect -1481 -16564 -1447 -16530
rect -1413 -16564 -1379 -16530
rect -1345 -16564 -1311 -16530
rect -1277 -16547 -1238 -16530
rect -808 -16530 -220 -16514
rect -808 -16547 -769 -16530
rect -1277 -16564 -1052 -16547
rect -2012 -16602 -1052 -16564
rect -994 -16564 -769 -16547
rect -735 -16564 -701 -16530
rect -667 -16564 -633 -16530
rect -599 -16564 -565 -16530
rect -531 -16564 -497 -16530
rect -463 -16564 -429 -16530
rect -395 -16564 -361 -16530
rect -327 -16564 -293 -16530
rect -259 -16547 -220 -16530
rect -259 -16564 -34 -16547
rect -994 -16602 -34 -16564
rect 2812 -16580 3400 -16564
rect 2812 -16597 2851 -16580
rect 2626 -16614 2851 -16597
rect 2885 -16614 2919 -16580
rect 2953 -16614 2987 -16580
rect 3021 -16614 3055 -16580
rect 3089 -16614 3123 -16580
rect 3157 -16614 3191 -16580
rect 3225 -16614 3259 -16580
rect 3293 -16614 3327 -16580
rect 3361 -16597 3400 -16580
rect 3830 -16580 4418 -16564
rect 3830 -16597 3869 -16580
rect 3361 -16614 3586 -16597
rect 2626 -16652 3586 -16614
rect 3644 -16614 3869 -16597
rect 3903 -16614 3937 -16580
rect 3971 -16614 4005 -16580
rect 4039 -16614 4073 -16580
rect 4107 -16614 4141 -16580
rect 4175 -16614 4209 -16580
rect 4243 -16614 4277 -16580
rect 4311 -16614 4345 -16580
rect 4379 -16597 4418 -16580
rect 4848 -16580 5436 -16564
rect 4848 -16597 4887 -16580
rect 4379 -16614 4604 -16597
rect 3644 -16652 4604 -16614
rect 4662 -16614 4887 -16597
rect 4921 -16614 4955 -16580
rect 4989 -16614 5023 -16580
rect 5057 -16614 5091 -16580
rect 5125 -16614 5159 -16580
rect 5193 -16614 5227 -16580
rect 5261 -16614 5295 -16580
rect 5329 -16614 5363 -16580
rect 5397 -16597 5436 -16580
rect 5866 -16580 6454 -16564
rect 5866 -16597 5905 -16580
rect 5397 -16614 5622 -16597
rect 4662 -16652 5622 -16614
rect 5680 -16614 5905 -16597
rect 5939 -16614 5973 -16580
rect 6007 -16614 6041 -16580
rect 6075 -16614 6109 -16580
rect 6143 -16614 6177 -16580
rect 6211 -16614 6245 -16580
rect 6279 -16614 6313 -16580
rect 6347 -16614 6381 -16580
rect 6415 -16597 6454 -16580
rect 6884 -16580 7472 -16564
rect 6884 -16597 6923 -16580
rect 6415 -16614 6640 -16597
rect 5680 -16652 6640 -16614
rect 6698 -16614 6923 -16597
rect 6957 -16614 6991 -16580
rect 7025 -16614 7059 -16580
rect 7093 -16614 7127 -16580
rect 7161 -16614 7195 -16580
rect 7229 -16614 7263 -16580
rect 7297 -16614 7331 -16580
rect 7365 -16614 7399 -16580
rect 7433 -16597 7472 -16580
rect 7902 -16580 8490 -16564
rect 7902 -16597 7941 -16580
rect 7433 -16614 7658 -16597
rect 6698 -16652 7658 -16614
rect 7716 -16614 7941 -16597
rect 7975 -16614 8009 -16580
rect 8043 -16614 8077 -16580
rect 8111 -16614 8145 -16580
rect 8179 -16614 8213 -16580
rect 8247 -16614 8281 -16580
rect 8315 -16614 8349 -16580
rect 8383 -16614 8417 -16580
rect 8451 -16597 8490 -16580
rect 8920 -16580 9508 -16564
rect 8920 -16597 8959 -16580
rect 8451 -16614 8676 -16597
rect 7716 -16652 8676 -16614
rect 8734 -16614 8959 -16597
rect 8993 -16614 9027 -16580
rect 9061 -16614 9095 -16580
rect 9129 -16614 9163 -16580
rect 9197 -16614 9231 -16580
rect 9265 -16614 9299 -16580
rect 9333 -16614 9367 -16580
rect 9401 -16614 9435 -16580
rect 9469 -16597 9508 -16580
rect 9938 -16580 10526 -16564
rect 9938 -16597 9977 -16580
rect 9469 -16614 9694 -16597
rect 8734 -16652 9694 -16614
rect 9752 -16614 9977 -16597
rect 10011 -16614 10045 -16580
rect 10079 -16614 10113 -16580
rect 10147 -16614 10181 -16580
rect 10215 -16614 10249 -16580
rect 10283 -16614 10317 -16580
rect 10351 -16614 10385 -16580
rect 10419 -16614 10453 -16580
rect 10487 -16597 10526 -16580
rect 10956 -16580 11544 -16564
rect 10956 -16597 10995 -16580
rect 10487 -16614 10712 -16597
rect 9752 -16652 10712 -16614
rect 10770 -16614 10995 -16597
rect 11029 -16614 11063 -16580
rect 11097 -16614 11131 -16580
rect 11165 -16614 11199 -16580
rect 11233 -16614 11267 -16580
rect 11301 -16614 11335 -16580
rect 11369 -16614 11403 -16580
rect 11437 -16614 11471 -16580
rect 11505 -16597 11544 -16580
rect 11974 -16580 12562 -16564
rect 11974 -16597 12013 -16580
rect 11505 -16614 11730 -16597
rect 10770 -16652 11730 -16614
rect 11788 -16614 12013 -16597
rect 12047 -16614 12081 -16580
rect 12115 -16614 12149 -16580
rect 12183 -16614 12217 -16580
rect 12251 -16614 12285 -16580
rect 12319 -16614 12353 -16580
rect 12387 -16614 12421 -16580
rect 12455 -16614 12489 -16580
rect 12523 -16597 12562 -16580
rect 12992 -16580 13580 -16564
rect 12992 -16597 13031 -16580
rect 12523 -16614 12748 -16597
rect 11788 -16652 12748 -16614
rect 12806 -16614 13031 -16597
rect 13065 -16614 13099 -16580
rect 13133 -16614 13167 -16580
rect 13201 -16614 13235 -16580
rect 13269 -16614 13303 -16580
rect 13337 -16614 13371 -16580
rect 13405 -16614 13439 -16580
rect 13473 -16614 13507 -16580
rect 13541 -16597 13580 -16580
rect 14010 -16580 14598 -16564
rect 14010 -16597 14049 -16580
rect 13541 -16614 13766 -16597
rect 12806 -16652 13766 -16614
rect 13824 -16614 14049 -16597
rect 14083 -16614 14117 -16580
rect 14151 -16614 14185 -16580
rect 14219 -16614 14253 -16580
rect 14287 -16614 14321 -16580
rect 14355 -16614 14389 -16580
rect 14423 -16614 14457 -16580
rect 14491 -16614 14525 -16580
rect 14559 -16597 14598 -16580
rect 15028 -16580 15616 -16564
rect 15028 -16597 15067 -16580
rect 14559 -16614 14784 -16597
rect 13824 -16652 14784 -16614
rect 14842 -16614 15067 -16597
rect 15101 -16614 15135 -16580
rect 15169 -16614 15203 -16580
rect 15237 -16614 15271 -16580
rect 15305 -16614 15339 -16580
rect 15373 -16614 15407 -16580
rect 15441 -16614 15475 -16580
rect 15509 -16614 15543 -16580
rect 15577 -16597 15616 -16580
rect 16046 -16580 16634 -16564
rect 16046 -16597 16085 -16580
rect 15577 -16614 15802 -16597
rect 14842 -16652 15802 -16614
rect 15860 -16614 16085 -16597
rect 16119 -16614 16153 -16580
rect 16187 -16614 16221 -16580
rect 16255 -16614 16289 -16580
rect 16323 -16614 16357 -16580
rect 16391 -16614 16425 -16580
rect 16459 -16614 16493 -16580
rect 16527 -16614 16561 -16580
rect 16595 -16597 16634 -16580
rect 17064 -16580 17652 -16564
rect 17064 -16597 17103 -16580
rect 16595 -16614 16820 -16597
rect 15860 -16652 16820 -16614
rect 16878 -16614 17103 -16597
rect 17137 -16614 17171 -16580
rect 17205 -16614 17239 -16580
rect 17273 -16614 17307 -16580
rect 17341 -16614 17375 -16580
rect 17409 -16614 17443 -16580
rect 17477 -16614 17511 -16580
rect 17545 -16614 17579 -16580
rect 17613 -16597 17652 -16580
rect 18082 -16580 18670 -16564
rect 18082 -16597 18121 -16580
rect 17613 -16614 17838 -16597
rect 16878 -16652 17838 -16614
rect 17896 -16614 18121 -16597
rect 18155 -16614 18189 -16580
rect 18223 -16614 18257 -16580
rect 18291 -16614 18325 -16580
rect 18359 -16614 18393 -16580
rect 18427 -16614 18461 -16580
rect 18495 -16614 18529 -16580
rect 18563 -16614 18597 -16580
rect 18631 -16597 18670 -16580
rect 19100 -16580 19688 -16564
rect 19100 -16597 19139 -16580
rect 18631 -16614 18856 -16597
rect 17896 -16652 18856 -16614
rect 18914 -16614 19139 -16597
rect 19173 -16614 19207 -16580
rect 19241 -16614 19275 -16580
rect 19309 -16614 19343 -16580
rect 19377 -16614 19411 -16580
rect 19445 -16614 19479 -16580
rect 19513 -16614 19547 -16580
rect 19581 -16614 19615 -16580
rect 19649 -16597 19688 -16580
rect 20118 -16580 20706 -16564
rect 20118 -16597 20157 -16580
rect 19649 -16614 19874 -16597
rect 18914 -16652 19874 -16614
rect 19932 -16614 20157 -16597
rect 20191 -16614 20225 -16580
rect 20259 -16614 20293 -16580
rect 20327 -16614 20361 -16580
rect 20395 -16614 20429 -16580
rect 20463 -16614 20497 -16580
rect 20531 -16614 20565 -16580
rect 20599 -16614 20633 -16580
rect 20667 -16597 20706 -16580
rect 21136 -16580 21724 -16564
rect 21136 -16597 21175 -16580
rect 20667 -16614 20892 -16597
rect 19932 -16652 20892 -16614
rect 20950 -16614 21175 -16597
rect 21209 -16614 21243 -16580
rect 21277 -16614 21311 -16580
rect 21345 -16614 21379 -16580
rect 21413 -16614 21447 -16580
rect 21481 -16614 21515 -16580
rect 21549 -16614 21583 -16580
rect 21617 -16614 21651 -16580
rect 21685 -16597 21724 -16580
rect 22154 -16580 22742 -16564
rect 22154 -16597 22193 -16580
rect 21685 -16614 21910 -16597
rect 20950 -16652 21910 -16614
rect 21968 -16614 22193 -16597
rect 22227 -16614 22261 -16580
rect 22295 -16614 22329 -16580
rect 22363 -16614 22397 -16580
rect 22431 -16614 22465 -16580
rect 22499 -16614 22533 -16580
rect 22567 -16614 22601 -16580
rect 22635 -16614 22669 -16580
rect 22703 -16597 22742 -16580
rect 22703 -16614 22928 -16597
rect 21968 -16652 22928 -16614
rect -9138 -17240 -8178 -17202
rect -9138 -17257 -8913 -17240
rect -8952 -17274 -8913 -17257
rect -8879 -17274 -8845 -17240
rect -8811 -17274 -8777 -17240
rect -8743 -17274 -8709 -17240
rect -8675 -17274 -8641 -17240
rect -8607 -17274 -8573 -17240
rect -8539 -17274 -8505 -17240
rect -8471 -17274 -8437 -17240
rect -8403 -17257 -8178 -17240
rect -8120 -17240 -7160 -17202
rect -8120 -17257 -7895 -17240
rect -8403 -17274 -8364 -17257
rect -8952 -17290 -8364 -17274
rect -7934 -17274 -7895 -17257
rect -7861 -17274 -7827 -17240
rect -7793 -17274 -7759 -17240
rect -7725 -17274 -7691 -17240
rect -7657 -17274 -7623 -17240
rect -7589 -17274 -7555 -17240
rect -7521 -17274 -7487 -17240
rect -7453 -17274 -7419 -17240
rect -7385 -17257 -7160 -17240
rect -7102 -17240 -6142 -17202
rect -7102 -17257 -6877 -17240
rect -7385 -17274 -7346 -17257
rect -7934 -17290 -7346 -17274
rect -6916 -17274 -6877 -17257
rect -6843 -17274 -6809 -17240
rect -6775 -17274 -6741 -17240
rect -6707 -17274 -6673 -17240
rect -6639 -17274 -6605 -17240
rect -6571 -17274 -6537 -17240
rect -6503 -17274 -6469 -17240
rect -6435 -17274 -6401 -17240
rect -6367 -17257 -6142 -17240
rect -6084 -17240 -5124 -17202
rect -6084 -17257 -5859 -17240
rect -6367 -17274 -6328 -17257
rect -6916 -17290 -6328 -17274
rect -5898 -17274 -5859 -17257
rect -5825 -17274 -5791 -17240
rect -5757 -17274 -5723 -17240
rect -5689 -17274 -5655 -17240
rect -5621 -17274 -5587 -17240
rect -5553 -17274 -5519 -17240
rect -5485 -17274 -5451 -17240
rect -5417 -17274 -5383 -17240
rect -5349 -17257 -5124 -17240
rect -5066 -17240 -4106 -17202
rect -5066 -17257 -4841 -17240
rect -5349 -17274 -5310 -17257
rect -5898 -17290 -5310 -17274
rect -4880 -17274 -4841 -17257
rect -4807 -17274 -4773 -17240
rect -4739 -17274 -4705 -17240
rect -4671 -17274 -4637 -17240
rect -4603 -17274 -4569 -17240
rect -4535 -17274 -4501 -17240
rect -4467 -17274 -4433 -17240
rect -4399 -17274 -4365 -17240
rect -4331 -17257 -4106 -17240
rect -4048 -17240 -3088 -17202
rect -4048 -17257 -3823 -17240
rect -4331 -17274 -4292 -17257
rect -4880 -17290 -4292 -17274
rect -3862 -17274 -3823 -17257
rect -3789 -17274 -3755 -17240
rect -3721 -17274 -3687 -17240
rect -3653 -17274 -3619 -17240
rect -3585 -17274 -3551 -17240
rect -3517 -17274 -3483 -17240
rect -3449 -17274 -3415 -17240
rect -3381 -17274 -3347 -17240
rect -3313 -17257 -3088 -17240
rect -3030 -17240 -2070 -17202
rect -3030 -17257 -2805 -17240
rect -3313 -17274 -3274 -17257
rect -3862 -17290 -3274 -17274
rect -2844 -17274 -2805 -17257
rect -2771 -17274 -2737 -17240
rect -2703 -17274 -2669 -17240
rect -2635 -17274 -2601 -17240
rect -2567 -17274 -2533 -17240
rect -2499 -17274 -2465 -17240
rect -2431 -17274 -2397 -17240
rect -2363 -17274 -2329 -17240
rect -2295 -17257 -2070 -17240
rect -2012 -17240 -1052 -17202
rect -2012 -17257 -1787 -17240
rect -2295 -17274 -2256 -17257
rect -2844 -17290 -2256 -17274
rect -1826 -17274 -1787 -17257
rect -1753 -17274 -1719 -17240
rect -1685 -17274 -1651 -17240
rect -1617 -17274 -1583 -17240
rect -1549 -17274 -1515 -17240
rect -1481 -17274 -1447 -17240
rect -1413 -17274 -1379 -17240
rect -1345 -17274 -1311 -17240
rect -1277 -17257 -1052 -17240
rect -994 -17240 -34 -17202
rect -994 -17257 -769 -17240
rect -1277 -17274 -1238 -17257
rect -1826 -17290 -1238 -17274
rect -808 -17274 -769 -17257
rect -735 -17274 -701 -17240
rect -667 -17274 -633 -17240
rect -599 -17274 -565 -17240
rect -531 -17274 -497 -17240
rect -463 -17274 -429 -17240
rect -395 -17274 -361 -17240
rect -327 -17274 -293 -17240
rect -259 -17257 -34 -17240
rect -259 -17274 -220 -17257
rect -808 -17290 -220 -17274
rect 2626 -17290 3586 -17252
rect 2626 -17307 2851 -17290
rect 2812 -17324 2851 -17307
rect 2885 -17324 2919 -17290
rect 2953 -17324 2987 -17290
rect 3021 -17324 3055 -17290
rect 3089 -17324 3123 -17290
rect 3157 -17324 3191 -17290
rect 3225 -17324 3259 -17290
rect 3293 -17324 3327 -17290
rect 3361 -17307 3586 -17290
rect 3644 -17290 4604 -17252
rect 3644 -17307 3869 -17290
rect 3361 -17324 3400 -17307
rect -8952 -17348 -8364 -17332
rect -8952 -17365 -8913 -17348
rect -9138 -17382 -8913 -17365
rect -8879 -17382 -8845 -17348
rect -8811 -17382 -8777 -17348
rect -8743 -17382 -8709 -17348
rect -8675 -17382 -8641 -17348
rect -8607 -17382 -8573 -17348
rect -8539 -17382 -8505 -17348
rect -8471 -17382 -8437 -17348
rect -8403 -17365 -8364 -17348
rect -7934 -17348 -7346 -17332
rect -7934 -17365 -7895 -17348
rect -8403 -17382 -8178 -17365
rect -9138 -17420 -8178 -17382
rect -8120 -17382 -7895 -17365
rect -7861 -17382 -7827 -17348
rect -7793 -17382 -7759 -17348
rect -7725 -17382 -7691 -17348
rect -7657 -17382 -7623 -17348
rect -7589 -17382 -7555 -17348
rect -7521 -17382 -7487 -17348
rect -7453 -17382 -7419 -17348
rect -7385 -17365 -7346 -17348
rect -6916 -17348 -6328 -17332
rect -6916 -17365 -6877 -17348
rect -7385 -17382 -7160 -17365
rect -8120 -17420 -7160 -17382
rect -7102 -17382 -6877 -17365
rect -6843 -17382 -6809 -17348
rect -6775 -17382 -6741 -17348
rect -6707 -17382 -6673 -17348
rect -6639 -17382 -6605 -17348
rect -6571 -17382 -6537 -17348
rect -6503 -17382 -6469 -17348
rect -6435 -17382 -6401 -17348
rect -6367 -17365 -6328 -17348
rect -5898 -17348 -5310 -17332
rect -5898 -17365 -5859 -17348
rect -6367 -17382 -6142 -17365
rect -7102 -17420 -6142 -17382
rect -6084 -17382 -5859 -17365
rect -5825 -17382 -5791 -17348
rect -5757 -17382 -5723 -17348
rect -5689 -17382 -5655 -17348
rect -5621 -17382 -5587 -17348
rect -5553 -17382 -5519 -17348
rect -5485 -17382 -5451 -17348
rect -5417 -17382 -5383 -17348
rect -5349 -17365 -5310 -17348
rect -4880 -17348 -4292 -17332
rect -4880 -17365 -4841 -17348
rect -5349 -17382 -5124 -17365
rect -6084 -17420 -5124 -17382
rect -5066 -17382 -4841 -17365
rect -4807 -17382 -4773 -17348
rect -4739 -17382 -4705 -17348
rect -4671 -17382 -4637 -17348
rect -4603 -17382 -4569 -17348
rect -4535 -17382 -4501 -17348
rect -4467 -17382 -4433 -17348
rect -4399 -17382 -4365 -17348
rect -4331 -17365 -4292 -17348
rect -3862 -17348 -3274 -17332
rect -3862 -17365 -3823 -17348
rect -4331 -17382 -4106 -17365
rect -5066 -17420 -4106 -17382
rect -4048 -17382 -3823 -17365
rect -3789 -17382 -3755 -17348
rect -3721 -17382 -3687 -17348
rect -3653 -17382 -3619 -17348
rect -3585 -17382 -3551 -17348
rect -3517 -17382 -3483 -17348
rect -3449 -17382 -3415 -17348
rect -3381 -17382 -3347 -17348
rect -3313 -17365 -3274 -17348
rect -2844 -17348 -2256 -17332
rect -2844 -17365 -2805 -17348
rect -3313 -17382 -3088 -17365
rect -4048 -17420 -3088 -17382
rect -3030 -17382 -2805 -17365
rect -2771 -17382 -2737 -17348
rect -2703 -17382 -2669 -17348
rect -2635 -17382 -2601 -17348
rect -2567 -17382 -2533 -17348
rect -2499 -17382 -2465 -17348
rect -2431 -17382 -2397 -17348
rect -2363 -17382 -2329 -17348
rect -2295 -17365 -2256 -17348
rect -1826 -17348 -1238 -17332
rect -1826 -17365 -1787 -17348
rect -2295 -17382 -2070 -17365
rect -3030 -17420 -2070 -17382
rect -2012 -17382 -1787 -17365
rect -1753 -17382 -1719 -17348
rect -1685 -17382 -1651 -17348
rect -1617 -17382 -1583 -17348
rect -1549 -17382 -1515 -17348
rect -1481 -17382 -1447 -17348
rect -1413 -17382 -1379 -17348
rect -1345 -17382 -1311 -17348
rect -1277 -17365 -1238 -17348
rect -808 -17348 -220 -17332
rect 2812 -17340 3400 -17324
rect 3830 -17324 3869 -17307
rect 3903 -17324 3937 -17290
rect 3971 -17324 4005 -17290
rect 4039 -17324 4073 -17290
rect 4107 -17324 4141 -17290
rect 4175 -17324 4209 -17290
rect 4243 -17324 4277 -17290
rect 4311 -17324 4345 -17290
rect 4379 -17307 4604 -17290
rect 4662 -17290 5622 -17252
rect 4662 -17307 4887 -17290
rect 4379 -17324 4418 -17307
rect 3830 -17340 4418 -17324
rect 4848 -17324 4887 -17307
rect 4921 -17324 4955 -17290
rect 4989 -17324 5023 -17290
rect 5057 -17324 5091 -17290
rect 5125 -17324 5159 -17290
rect 5193 -17324 5227 -17290
rect 5261 -17324 5295 -17290
rect 5329 -17324 5363 -17290
rect 5397 -17307 5622 -17290
rect 5680 -17290 6640 -17252
rect 5680 -17307 5905 -17290
rect 5397 -17324 5436 -17307
rect 4848 -17340 5436 -17324
rect 5866 -17324 5905 -17307
rect 5939 -17324 5973 -17290
rect 6007 -17324 6041 -17290
rect 6075 -17324 6109 -17290
rect 6143 -17324 6177 -17290
rect 6211 -17324 6245 -17290
rect 6279 -17324 6313 -17290
rect 6347 -17324 6381 -17290
rect 6415 -17307 6640 -17290
rect 6698 -17290 7658 -17252
rect 6698 -17307 6923 -17290
rect 6415 -17324 6454 -17307
rect 5866 -17340 6454 -17324
rect 6884 -17324 6923 -17307
rect 6957 -17324 6991 -17290
rect 7025 -17324 7059 -17290
rect 7093 -17324 7127 -17290
rect 7161 -17324 7195 -17290
rect 7229 -17324 7263 -17290
rect 7297 -17324 7331 -17290
rect 7365 -17324 7399 -17290
rect 7433 -17307 7658 -17290
rect 7716 -17290 8676 -17252
rect 7716 -17307 7941 -17290
rect 7433 -17324 7472 -17307
rect 6884 -17340 7472 -17324
rect 7902 -17324 7941 -17307
rect 7975 -17324 8009 -17290
rect 8043 -17324 8077 -17290
rect 8111 -17324 8145 -17290
rect 8179 -17324 8213 -17290
rect 8247 -17324 8281 -17290
rect 8315 -17324 8349 -17290
rect 8383 -17324 8417 -17290
rect 8451 -17307 8676 -17290
rect 8734 -17290 9694 -17252
rect 8734 -17307 8959 -17290
rect 8451 -17324 8490 -17307
rect 7902 -17340 8490 -17324
rect 8920 -17324 8959 -17307
rect 8993 -17324 9027 -17290
rect 9061 -17324 9095 -17290
rect 9129 -17324 9163 -17290
rect 9197 -17324 9231 -17290
rect 9265 -17324 9299 -17290
rect 9333 -17324 9367 -17290
rect 9401 -17324 9435 -17290
rect 9469 -17307 9694 -17290
rect 9752 -17290 10712 -17252
rect 9752 -17307 9977 -17290
rect 9469 -17324 9508 -17307
rect 8920 -17340 9508 -17324
rect 9938 -17324 9977 -17307
rect 10011 -17324 10045 -17290
rect 10079 -17324 10113 -17290
rect 10147 -17324 10181 -17290
rect 10215 -17324 10249 -17290
rect 10283 -17324 10317 -17290
rect 10351 -17324 10385 -17290
rect 10419 -17324 10453 -17290
rect 10487 -17307 10712 -17290
rect 10770 -17290 11730 -17252
rect 10770 -17307 10995 -17290
rect 10487 -17324 10526 -17307
rect 9938 -17340 10526 -17324
rect 10956 -17324 10995 -17307
rect 11029 -17324 11063 -17290
rect 11097 -17324 11131 -17290
rect 11165 -17324 11199 -17290
rect 11233 -17324 11267 -17290
rect 11301 -17324 11335 -17290
rect 11369 -17324 11403 -17290
rect 11437 -17324 11471 -17290
rect 11505 -17307 11730 -17290
rect 11788 -17290 12748 -17252
rect 11788 -17307 12013 -17290
rect 11505 -17324 11544 -17307
rect 10956 -17340 11544 -17324
rect 11974 -17324 12013 -17307
rect 12047 -17324 12081 -17290
rect 12115 -17324 12149 -17290
rect 12183 -17324 12217 -17290
rect 12251 -17324 12285 -17290
rect 12319 -17324 12353 -17290
rect 12387 -17324 12421 -17290
rect 12455 -17324 12489 -17290
rect 12523 -17307 12748 -17290
rect 12806 -17290 13766 -17252
rect 12806 -17307 13031 -17290
rect 12523 -17324 12562 -17307
rect 11974 -17340 12562 -17324
rect 12992 -17324 13031 -17307
rect 13065 -17324 13099 -17290
rect 13133 -17324 13167 -17290
rect 13201 -17324 13235 -17290
rect 13269 -17324 13303 -17290
rect 13337 -17324 13371 -17290
rect 13405 -17324 13439 -17290
rect 13473 -17324 13507 -17290
rect 13541 -17307 13766 -17290
rect 13824 -17290 14784 -17252
rect 13824 -17307 14049 -17290
rect 13541 -17324 13580 -17307
rect 12992 -17340 13580 -17324
rect 14010 -17324 14049 -17307
rect 14083 -17324 14117 -17290
rect 14151 -17324 14185 -17290
rect 14219 -17324 14253 -17290
rect 14287 -17324 14321 -17290
rect 14355 -17324 14389 -17290
rect 14423 -17324 14457 -17290
rect 14491 -17324 14525 -17290
rect 14559 -17307 14784 -17290
rect 14842 -17290 15802 -17252
rect 14842 -17307 15067 -17290
rect 14559 -17324 14598 -17307
rect 14010 -17340 14598 -17324
rect 15028 -17324 15067 -17307
rect 15101 -17324 15135 -17290
rect 15169 -17324 15203 -17290
rect 15237 -17324 15271 -17290
rect 15305 -17324 15339 -17290
rect 15373 -17324 15407 -17290
rect 15441 -17324 15475 -17290
rect 15509 -17324 15543 -17290
rect 15577 -17307 15802 -17290
rect 15860 -17290 16820 -17252
rect 15860 -17307 16085 -17290
rect 15577 -17324 15616 -17307
rect 15028 -17340 15616 -17324
rect 16046 -17324 16085 -17307
rect 16119 -17324 16153 -17290
rect 16187 -17324 16221 -17290
rect 16255 -17324 16289 -17290
rect 16323 -17324 16357 -17290
rect 16391 -17324 16425 -17290
rect 16459 -17324 16493 -17290
rect 16527 -17324 16561 -17290
rect 16595 -17307 16820 -17290
rect 16878 -17290 17838 -17252
rect 16878 -17307 17103 -17290
rect 16595 -17324 16634 -17307
rect 16046 -17340 16634 -17324
rect 17064 -17324 17103 -17307
rect 17137 -17324 17171 -17290
rect 17205 -17324 17239 -17290
rect 17273 -17324 17307 -17290
rect 17341 -17324 17375 -17290
rect 17409 -17324 17443 -17290
rect 17477 -17324 17511 -17290
rect 17545 -17324 17579 -17290
rect 17613 -17307 17838 -17290
rect 17896 -17290 18856 -17252
rect 17896 -17307 18121 -17290
rect 17613 -17324 17652 -17307
rect 17064 -17340 17652 -17324
rect 18082 -17324 18121 -17307
rect 18155 -17324 18189 -17290
rect 18223 -17324 18257 -17290
rect 18291 -17324 18325 -17290
rect 18359 -17324 18393 -17290
rect 18427 -17324 18461 -17290
rect 18495 -17324 18529 -17290
rect 18563 -17324 18597 -17290
rect 18631 -17307 18856 -17290
rect 18914 -17290 19874 -17252
rect 18914 -17307 19139 -17290
rect 18631 -17324 18670 -17307
rect 18082 -17340 18670 -17324
rect 19100 -17324 19139 -17307
rect 19173 -17324 19207 -17290
rect 19241 -17324 19275 -17290
rect 19309 -17324 19343 -17290
rect 19377 -17324 19411 -17290
rect 19445 -17324 19479 -17290
rect 19513 -17324 19547 -17290
rect 19581 -17324 19615 -17290
rect 19649 -17307 19874 -17290
rect 19932 -17290 20892 -17252
rect 19932 -17307 20157 -17290
rect 19649 -17324 19688 -17307
rect 19100 -17340 19688 -17324
rect 20118 -17324 20157 -17307
rect 20191 -17324 20225 -17290
rect 20259 -17324 20293 -17290
rect 20327 -17324 20361 -17290
rect 20395 -17324 20429 -17290
rect 20463 -17324 20497 -17290
rect 20531 -17324 20565 -17290
rect 20599 -17324 20633 -17290
rect 20667 -17307 20892 -17290
rect 20950 -17290 21910 -17252
rect 20950 -17307 21175 -17290
rect 20667 -17324 20706 -17307
rect 20118 -17340 20706 -17324
rect 21136 -17324 21175 -17307
rect 21209 -17324 21243 -17290
rect 21277 -17324 21311 -17290
rect 21345 -17324 21379 -17290
rect 21413 -17324 21447 -17290
rect 21481 -17324 21515 -17290
rect 21549 -17324 21583 -17290
rect 21617 -17324 21651 -17290
rect 21685 -17307 21910 -17290
rect 21968 -17290 22928 -17252
rect 21968 -17307 22193 -17290
rect 21685 -17324 21724 -17307
rect 21136 -17340 21724 -17324
rect 22154 -17324 22193 -17307
rect 22227 -17324 22261 -17290
rect 22295 -17324 22329 -17290
rect 22363 -17324 22397 -17290
rect 22431 -17324 22465 -17290
rect 22499 -17324 22533 -17290
rect 22567 -17324 22601 -17290
rect 22635 -17324 22669 -17290
rect 22703 -17307 22928 -17290
rect 22703 -17324 22742 -17307
rect 22154 -17340 22742 -17324
rect -808 -17365 -769 -17348
rect -1277 -17382 -1052 -17365
rect -2012 -17420 -1052 -17382
rect -994 -17382 -769 -17365
rect -735 -17382 -701 -17348
rect -667 -17382 -633 -17348
rect -599 -17382 -565 -17348
rect -531 -17382 -497 -17348
rect -463 -17382 -429 -17348
rect -395 -17382 -361 -17348
rect -327 -17382 -293 -17348
rect -259 -17365 -220 -17348
rect -259 -17382 -34 -17365
rect -994 -17420 -34 -17382
rect 2812 -17812 3400 -17796
rect 2812 -17829 2851 -17812
rect 2626 -17846 2851 -17829
rect 2885 -17846 2919 -17812
rect 2953 -17846 2987 -17812
rect 3021 -17846 3055 -17812
rect 3089 -17846 3123 -17812
rect 3157 -17846 3191 -17812
rect 3225 -17846 3259 -17812
rect 3293 -17846 3327 -17812
rect 3361 -17829 3400 -17812
rect 3830 -17812 4418 -17796
rect 3830 -17829 3869 -17812
rect 3361 -17846 3586 -17829
rect 2626 -17884 3586 -17846
rect 3644 -17846 3869 -17829
rect 3903 -17846 3937 -17812
rect 3971 -17846 4005 -17812
rect 4039 -17846 4073 -17812
rect 4107 -17846 4141 -17812
rect 4175 -17846 4209 -17812
rect 4243 -17846 4277 -17812
rect 4311 -17846 4345 -17812
rect 4379 -17829 4418 -17812
rect 4848 -17812 5436 -17796
rect 4848 -17829 4887 -17812
rect 4379 -17846 4604 -17829
rect 3644 -17884 4604 -17846
rect 4662 -17846 4887 -17829
rect 4921 -17846 4955 -17812
rect 4989 -17846 5023 -17812
rect 5057 -17846 5091 -17812
rect 5125 -17846 5159 -17812
rect 5193 -17846 5227 -17812
rect 5261 -17846 5295 -17812
rect 5329 -17846 5363 -17812
rect 5397 -17829 5436 -17812
rect 5866 -17812 6454 -17796
rect 5866 -17829 5905 -17812
rect 5397 -17846 5622 -17829
rect 4662 -17884 5622 -17846
rect 5680 -17846 5905 -17829
rect 5939 -17846 5973 -17812
rect 6007 -17846 6041 -17812
rect 6075 -17846 6109 -17812
rect 6143 -17846 6177 -17812
rect 6211 -17846 6245 -17812
rect 6279 -17846 6313 -17812
rect 6347 -17846 6381 -17812
rect 6415 -17829 6454 -17812
rect 6884 -17812 7472 -17796
rect 6884 -17829 6923 -17812
rect 6415 -17846 6640 -17829
rect 5680 -17884 6640 -17846
rect 6698 -17846 6923 -17829
rect 6957 -17846 6991 -17812
rect 7025 -17846 7059 -17812
rect 7093 -17846 7127 -17812
rect 7161 -17846 7195 -17812
rect 7229 -17846 7263 -17812
rect 7297 -17846 7331 -17812
rect 7365 -17846 7399 -17812
rect 7433 -17829 7472 -17812
rect 7902 -17812 8490 -17796
rect 7902 -17829 7941 -17812
rect 7433 -17846 7658 -17829
rect 6698 -17884 7658 -17846
rect 7716 -17846 7941 -17829
rect 7975 -17846 8009 -17812
rect 8043 -17846 8077 -17812
rect 8111 -17846 8145 -17812
rect 8179 -17846 8213 -17812
rect 8247 -17846 8281 -17812
rect 8315 -17846 8349 -17812
rect 8383 -17846 8417 -17812
rect 8451 -17829 8490 -17812
rect 8920 -17812 9508 -17796
rect 8920 -17829 8959 -17812
rect 8451 -17846 8676 -17829
rect 7716 -17884 8676 -17846
rect 8734 -17846 8959 -17829
rect 8993 -17846 9027 -17812
rect 9061 -17846 9095 -17812
rect 9129 -17846 9163 -17812
rect 9197 -17846 9231 -17812
rect 9265 -17846 9299 -17812
rect 9333 -17846 9367 -17812
rect 9401 -17846 9435 -17812
rect 9469 -17829 9508 -17812
rect 9938 -17812 10526 -17796
rect 9938 -17829 9977 -17812
rect 9469 -17846 9694 -17829
rect 8734 -17884 9694 -17846
rect 9752 -17846 9977 -17829
rect 10011 -17846 10045 -17812
rect 10079 -17846 10113 -17812
rect 10147 -17846 10181 -17812
rect 10215 -17846 10249 -17812
rect 10283 -17846 10317 -17812
rect 10351 -17846 10385 -17812
rect 10419 -17846 10453 -17812
rect 10487 -17829 10526 -17812
rect 10956 -17812 11544 -17796
rect 10956 -17829 10995 -17812
rect 10487 -17846 10712 -17829
rect 9752 -17884 10712 -17846
rect 10770 -17846 10995 -17829
rect 11029 -17846 11063 -17812
rect 11097 -17846 11131 -17812
rect 11165 -17846 11199 -17812
rect 11233 -17846 11267 -17812
rect 11301 -17846 11335 -17812
rect 11369 -17846 11403 -17812
rect 11437 -17846 11471 -17812
rect 11505 -17829 11544 -17812
rect 11974 -17812 12562 -17796
rect 11974 -17829 12013 -17812
rect 11505 -17846 11730 -17829
rect 10770 -17884 11730 -17846
rect 11788 -17846 12013 -17829
rect 12047 -17846 12081 -17812
rect 12115 -17846 12149 -17812
rect 12183 -17846 12217 -17812
rect 12251 -17846 12285 -17812
rect 12319 -17846 12353 -17812
rect 12387 -17846 12421 -17812
rect 12455 -17846 12489 -17812
rect 12523 -17829 12562 -17812
rect 12992 -17812 13580 -17796
rect 12992 -17829 13031 -17812
rect 12523 -17846 12748 -17829
rect 11788 -17884 12748 -17846
rect 12806 -17846 13031 -17829
rect 13065 -17846 13099 -17812
rect 13133 -17846 13167 -17812
rect 13201 -17846 13235 -17812
rect 13269 -17846 13303 -17812
rect 13337 -17846 13371 -17812
rect 13405 -17846 13439 -17812
rect 13473 -17846 13507 -17812
rect 13541 -17829 13580 -17812
rect 14010 -17812 14598 -17796
rect 14010 -17829 14049 -17812
rect 13541 -17846 13766 -17829
rect 12806 -17884 13766 -17846
rect 13824 -17846 14049 -17829
rect 14083 -17846 14117 -17812
rect 14151 -17846 14185 -17812
rect 14219 -17846 14253 -17812
rect 14287 -17846 14321 -17812
rect 14355 -17846 14389 -17812
rect 14423 -17846 14457 -17812
rect 14491 -17846 14525 -17812
rect 14559 -17829 14598 -17812
rect 15028 -17812 15616 -17796
rect 15028 -17829 15067 -17812
rect 14559 -17846 14784 -17829
rect 13824 -17884 14784 -17846
rect 14842 -17846 15067 -17829
rect 15101 -17846 15135 -17812
rect 15169 -17846 15203 -17812
rect 15237 -17846 15271 -17812
rect 15305 -17846 15339 -17812
rect 15373 -17846 15407 -17812
rect 15441 -17846 15475 -17812
rect 15509 -17846 15543 -17812
rect 15577 -17829 15616 -17812
rect 16046 -17812 16634 -17796
rect 16046 -17829 16085 -17812
rect 15577 -17846 15802 -17829
rect 14842 -17884 15802 -17846
rect 15860 -17846 16085 -17829
rect 16119 -17846 16153 -17812
rect 16187 -17846 16221 -17812
rect 16255 -17846 16289 -17812
rect 16323 -17846 16357 -17812
rect 16391 -17846 16425 -17812
rect 16459 -17846 16493 -17812
rect 16527 -17846 16561 -17812
rect 16595 -17829 16634 -17812
rect 17064 -17812 17652 -17796
rect 17064 -17829 17103 -17812
rect 16595 -17846 16820 -17829
rect 15860 -17884 16820 -17846
rect 16878 -17846 17103 -17829
rect 17137 -17846 17171 -17812
rect 17205 -17846 17239 -17812
rect 17273 -17846 17307 -17812
rect 17341 -17846 17375 -17812
rect 17409 -17846 17443 -17812
rect 17477 -17846 17511 -17812
rect 17545 -17846 17579 -17812
rect 17613 -17829 17652 -17812
rect 18082 -17812 18670 -17796
rect 18082 -17829 18121 -17812
rect 17613 -17846 17838 -17829
rect 16878 -17884 17838 -17846
rect 17896 -17846 18121 -17829
rect 18155 -17846 18189 -17812
rect 18223 -17846 18257 -17812
rect 18291 -17846 18325 -17812
rect 18359 -17846 18393 -17812
rect 18427 -17846 18461 -17812
rect 18495 -17846 18529 -17812
rect 18563 -17846 18597 -17812
rect 18631 -17829 18670 -17812
rect 19100 -17812 19688 -17796
rect 19100 -17829 19139 -17812
rect 18631 -17846 18856 -17829
rect 17896 -17884 18856 -17846
rect 18914 -17846 19139 -17829
rect 19173 -17846 19207 -17812
rect 19241 -17846 19275 -17812
rect 19309 -17846 19343 -17812
rect 19377 -17846 19411 -17812
rect 19445 -17846 19479 -17812
rect 19513 -17846 19547 -17812
rect 19581 -17846 19615 -17812
rect 19649 -17829 19688 -17812
rect 20118 -17812 20706 -17796
rect 20118 -17829 20157 -17812
rect 19649 -17846 19874 -17829
rect 18914 -17884 19874 -17846
rect 19932 -17846 20157 -17829
rect 20191 -17846 20225 -17812
rect 20259 -17846 20293 -17812
rect 20327 -17846 20361 -17812
rect 20395 -17846 20429 -17812
rect 20463 -17846 20497 -17812
rect 20531 -17846 20565 -17812
rect 20599 -17846 20633 -17812
rect 20667 -17829 20706 -17812
rect 21136 -17812 21724 -17796
rect 21136 -17829 21175 -17812
rect 20667 -17846 20892 -17829
rect 19932 -17884 20892 -17846
rect 20950 -17846 21175 -17829
rect 21209 -17846 21243 -17812
rect 21277 -17846 21311 -17812
rect 21345 -17846 21379 -17812
rect 21413 -17846 21447 -17812
rect 21481 -17846 21515 -17812
rect 21549 -17846 21583 -17812
rect 21617 -17846 21651 -17812
rect 21685 -17829 21724 -17812
rect 22154 -17812 22742 -17796
rect 22154 -17829 22193 -17812
rect 21685 -17846 21910 -17829
rect 20950 -17884 21910 -17846
rect 21968 -17846 22193 -17829
rect 22227 -17846 22261 -17812
rect 22295 -17846 22329 -17812
rect 22363 -17846 22397 -17812
rect 22431 -17846 22465 -17812
rect 22499 -17846 22533 -17812
rect 22567 -17846 22601 -17812
rect 22635 -17846 22669 -17812
rect 22703 -17829 22742 -17812
rect 22703 -17846 22928 -17829
rect 21968 -17884 22928 -17846
rect -9138 -18058 -8178 -18020
rect -9138 -18075 -8913 -18058
rect -8952 -18092 -8913 -18075
rect -8879 -18092 -8845 -18058
rect -8811 -18092 -8777 -18058
rect -8743 -18092 -8709 -18058
rect -8675 -18092 -8641 -18058
rect -8607 -18092 -8573 -18058
rect -8539 -18092 -8505 -18058
rect -8471 -18092 -8437 -18058
rect -8403 -18075 -8178 -18058
rect -8120 -18058 -7160 -18020
rect -8120 -18075 -7895 -18058
rect -8403 -18092 -8364 -18075
rect -8952 -18108 -8364 -18092
rect -7934 -18092 -7895 -18075
rect -7861 -18092 -7827 -18058
rect -7793 -18092 -7759 -18058
rect -7725 -18092 -7691 -18058
rect -7657 -18092 -7623 -18058
rect -7589 -18092 -7555 -18058
rect -7521 -18092 -7487 -18058
rect -7453 -18092 -7419 -18058
rect -7385 -18075 -7160 -18058
rect -7102 -18058 -6142 -18020
rect -7102 -18075 -6877 -18058
rect -7385 -18092 -7346 -18075
rect -7934 -18108 -7346 -18092
rect -6916 -18092 -6877 -18075
rect -6843 -18092 -6809 -18058
rect -6775 -18092 -6741 -18058
rect -6707 -18092 -6673 -18058
rect -6639 -18092 -6605 -18058
rect -6571 -18092 -6537 -18058
rect -6503 -18092 -6469 -18058
rect -6435 -18092 -6401 -18058
rect -6367 -18075 -6142 -18058
rect -6084 -18058 -5124 -18020
rect -6084 -18075 -5859 -18058
rect -6367 -18092 -6328 -18075
rect -6916 -18108 -6328 -18092
rect -5898 -18092 -5859 -18075
rect -5825 -18092 -5791 -18058
rect -5757 -18092 -5723 -18058
rect -5689 -18092 -5655 -18058
rect -5621 -18092 -5587 -18058
rect -5553 -18092 -5519 -18058
rect -5485 -18092 -5451 -18058
rect -5417 -18092 -5383 -18058
rect -5349 -18075 -5124 -18058
rect -5066 -18058 -4106 -18020
rect -5066 -18075 -4841 -18058
rect -5349 -18092 -5310 -18075
rect -5898 -18108 -5310 -18092
rect -4880 -18092 -4841 -18075
rect -4807 -18092 -4773 -18058
rect -4739 -18092 -4705 -18058
rect -4671 -18092 -4637 -18058
rect -4603 -18092 -4569 -18058
rect -4535 -18092 -4501 -18058
rect -4467 -18092 -4433 -18058
rect -4399 -18092 -4365 -18058
rect -4331 -18075 -4106 -18058
rect -4048 -18058 -3088 -18020
rect -4048 -18075 -3823 -18058
rect -4331 -18092 -4292 -18075
rect -4880 -18108 -4292 -18092
rect -3862 -18092 -3823 -18075
rect -3789 -18092 -3755 -18058
rect -3721 -18092 -3687 -18058
rect -3653 -18092 -3619 -18058
rect -3585 -18092 -3551 -18058
rect -3517 -18092 -3483 -18058
rect -3449 -18092 -3415 -18058
rect -3381 -18092 -3347 -18058
rect -3313 -18075 -3088 -18058
rect -3030 -18058 -2070 -18020
rect -3030 -18075 -2805 -18058
rect -3313 -18092 -3274 -18075
rect -3862 -18108 -3274 -18092
rect -2844 -18092 -2805 -18075
rect -2771 -18092 -2737 -18058
rect -2703 -18092 -2669 -18058
rect -2635 -18092 -2601 -18058
rect -2567 -18092 -2533 -18058
rect -2499 -18092 -2465 -18058
rect -2431 -18092 -2397 -18058
rect -2363 -18092 -2329 -18058
rect -2295 -18075 -2070 -18058
rect -2012 -18058 -1052 -18020
rect -2012 -18075 -1787 -18058
rect -2295 -18092 -2256 -18075
rect -2844 -18108 -2256 -18092
rect -1826 -18092 -1787 -18075
rect -1753 -18092 -1719 -18058
rect -1685 -18092 -1651 -18058
rect -1617 -18092 -1583 -18058
rect -1549 -18092 -1515 -18058
rect -1481 -18092 -1447 -18058
rect -1413 -18092 -1379 -18058
rect -1345 -18092 -1311 -18058
rect -1277 -18075 -1052 -18058
rect -994 -18058 -34 -18020
rect -994 -18075 -769 -18058
rect -1277 -18092 -1238 -18075
rect -1826 -18108 -1238 -18092
rect -808 -18092 -769 -18075
rect -735 -18092 -701 -18058
rect -667 -18092 -633 -18058
rect -599 -18092 -565 -18058
rect -531 -18092 -497 -18058
rect -463 -18092 -429 -18058
rect -395 -18092 -361 -18058
rect -327 -18092 -293 -18058
rect -259 -18075 -34 -18058
rect -259 -18092 -220 -18075
rect -808 -18108 -220 -18092
rect -8952 -18166 -8364 -18150
rect -8952 -18183 -8913 -18166
rect -9138 -18200 -8913 -18183
rect -8879 -18200 -8845 -18166
rect -8811 -18200 -8777 -18166
rect -8743 -18200 -8709 -18166
rect -8675 -18200 -8641 -18166
rect -8607 -18200 -8573 -18166
rect -8539 -18200 -8505 -18166
rect -8471 -18200 -8437 -18166
rect -8403 -18183 -8364 -18166
rect -7934 -18166 -7346 -18150
rect -7934 -18183 -7895 -18166
rect -8403 -18200 -8178 -18183
rect -9138 -18238 -8178 -18200
rect -8120 -18200 -7895 -18183
rect -7861 -18200 -7827 -18166
rect -7793 -18200 -7759 -18166
rect -7725 -18200 -7691 -18166
rect -7657 -18200 -7623 -18166
rect -7589 -18200 -7555 -18166
rect -7521 -18200 -7487 -18166
rect -7453 -18200 -7419 -18166
rect -7385 -18183 -7346 -18166
rect -6916 -18166 -6328 -18150
rect -6916 -18183 -6877 -18166
rect -7385 -18200 -7160 -18183
rect -8120 -18238 -7160 -18200
rect -7102 -18200 -6877 -18183
rect -6843 -18200 -6809 -18166
rect -6775 -18200 -6741 -18166
rect -6707 -18200 -6673 -18166
rect -6639 -18200 -6605 -18166
rect -6571 -18200 -6537 -18166
rect -6503 -18200 -6469 -18166
rect -6435 -18200 -6401 -18166
rect -6367 -18183 -6328 -18166
rect -5898 -18166 -5310 -18150
rect -5898 -18183 -5859 -18166
rect -6367 -18200 -6142 -18183
rect -7102 -18238 -6142 -18200
rect -6084 -18200 -5859 -18183
rect -5825 -18200 -5791 -18166
rect -5757 -18200 -5723 -18166
rect -5689 -18200 -5655 -18166
rect -5621 -18200 -5587 -18166
rect -5553 -18200 -5519 -18166
rect -5485 -18200 -5451 -18166
rect -5417 -18200 -5383 -18166
rect -5349 -18183 -5310 -18166
rect -4880 -18166 -4292 -18150
rect -4880 -18183 -4841 -18166
rect -5349 -18200 -5124 -18183
rect -6084 -18238 -5124 -18200
rect -5066 -18200 -4841 -18183
rect -4807 -18200 -4773 -18166
rect -4739 -18200 -4705 -18166
rect -4671 -18200 -4637 -18166
rect -4603 -18200 -4569 -18166
rect -4535 -18200 -4501 -18166
rect -4467 -18200 -4433 -18166
rect -4399 -18200 -4365 -18166
rect -4331 -18183 -4292 -18166
rect -3862 -18166 -3274 -18150
rect -3862 -18183 -3823 -18166
rect -4331 -18200 -4106 -18183
rect -5066 -18238 -4106 -18200
rect -4048 -18200 -3823 -18183
rect -3789 -18200 -3755 -18166
rect -3721 -18200 -3687 -18166
rect -3653 -18200 -3619 -18166
rect -3585 -18200 -3551 -18166
rect -3517 -18200 -3483 -18166
rect -3449 -18200 -3415 -18166
rect -3381 -18200 -3347 -18166
rect -3313 -18183 -3274 -18166
rect -2844 -18166 -2256 -18150
rect -2844 -18183 -2805 -18166
rect -3313 -18200 -3088 -18183
rect -4048 -18238 -3088 -18200
rect -3030 -18200 -2805 -18183
rect -2771 -18200 -2737 -18166
rect -2703 -18200 -2669 -18166
rect -2635 -18200 -2601 -18166
rect -2567 -18200 -2533 -18166
rect -2499 -18200 -2465 -18166
rect -2431 -18200 -2397 -18166
rect -2363 -18200 -2329 -18166
rect -2295 -18183 -2256 -18166
rect -1826 -18166 -1238 -18150
rect -1826 -18183 -1787 -18166
rect -2295 -18200 -2070 -18183
rect -3030 -18238 -2070 -18200
rect -2012 -18200 -1787 -18183
rect -1753 -18200 -1719 -18166
rect -1685 -18200 -1651 -18166
rect -1617 -18200 -1583 -18166
rect -1549 -18200 -1515 -18166
rect -1481 -18200 -1447 -18166
rect -1413 -18200 -1379 -18166
rect -1345 -18200 -1311 -18166
rect -1277 -18183 -1238 -18166
rect -808 -18166 -220 -18150
rect -808 -18183 -769 -18166
rect -1277 -18200 -1052 -18183
rect -2012 -18238 -1052 -18200
rect -994 -18200 -769 -18183
rect -735 -18200 -701 -18166
rect -667 -18200 -633 -18166
rect -599 -18200 -565 -18166
rect -531 -18200 -497 -18166
rect -463 -18200 -429 -18166
rect -395 -18200 -361 -18166
rect -327 -18200 -293 -18166
rect -259 -18183 -220 -18166
rect -259 -18200 -34 -18183
rect -994 -18238 -34 -18200
rect 2626 -18522 3586 -18484
rect 2626 -18539 2851 -18522
rect 2812 -18556 2851 -18539
rect 2885 -18556 2919 -18522
rect 2953 -18556 2987 -18522
rect 3021 -18556 3055 -18522
rect 3089 -18556 3123 -18522
rect 3157 -18556 3191 -18522
rect 3225 -18556 3259 -18522
rect 3293 -18556 3327 -18522
rect 3361 -18539 3586 -18522
rect 3644 -18522 4604 -18484
rect 3644 -18539 3869 -18522
rect 3361 -18556 3400 -18539
rect 2812 -18572 3400 -18556
rect 3830 -18556 3869 -18539
rect 3903 -18556 3937 -18522
rect 3971 -18556 4005 -18522
rect 4039 -18556 4073 -18522
rect 4107 -18556 4141 -18522
rect 4175 -18556 4209 -18522
rect 4243 -18556 4277 -18522
rect 4311 -18556 4345 -18522
rect 4379 -18539 4604 -18522
rect 4662 -18522 5622 -18484
rect 4662 -18539 4887 -18522
rect 4379 -18556 4418 -18539
rect 3830 -18572 4418 -18556
rect 4848 -18556 4887 -18539
rect 4921 -18556 4955 -18522
rect 4989 -18556 5023 -18522
rect 5057 -18556 5091 -18522
rect 5125 -18556 5159 -18522
rect 5193 -18556 5227 -18522
rect 5261 -18556 5295 -18522
rect 5329 -18556 5363 -18522
rect 5397 -18539 5622 -18522
rect 5680 -18522 6640 -18484
rect 5680 -18539 5905 -18522
rect 5397 -18556 5436 -18539
rect 4848 -18572 5436 -18556
rect 5866 -18556 5905 -18539
rect 5939 -18556 5973 -18522
rect 6007 -18556 6041 -18522
rect 6075 -18556 6109 -18522
rect 6143 -18556 6177 -18522
rect 6211 -18556 6245 -18522
rect 6279 -18556 6313 -18522
rect 6347 -18556 6381 -18522
rect 6415 -18539 6640 -18522
rect 6698 -18522 7658 -18484
rect 6698 -18539 6923 -18522
rect 6415 -18556 6454 -18539
rect 5866 -18572 6454 -18556
rect 6884 -18556 6923 -18539
rect 6957 -18556 6991 -18522
rect 7025 -18556 7059 -18522
rect 7093 -18556 7127 -18522
rect 7161 -18556 7195 -18522
rect 7229 -18556 7263 -18522
rect 7297 -18556 7331 -18522
rect 7365 -18556 7399 -18522
rect 7433 -18539 7658 -18522
rect 7716 -18522 8676 -18484
rect 7716 -18539 7941 -18522
rect 7433 -18556 7472 -18539
rect 6884 -18572 7472 -18556
rect 7902 -18556 7941 -18539
rect 7975 -18556 8009 -18522
rect 8043 -18556 8077 -18522
rect 8111 -18556 8145 -18522
rect 8179 -18556 8213 -18522
rect 8247 -18556 8281 -18522
rect 8315 -18556 8349 -18522
rect 8383 -18556 8417 -18522
rect 8451 -18539 8676 -18522
rect 8734 -18522 9694 -18484
rect 8734 -18539 8959 -18522
rect 8451 -18556 8490 -18539
rect 7902 -18572 8490 -18556
rect 8920 -18556 8959 -18539
rect 8993 -18556 9027 -18522
rect 9061 -18556 9095 -18522
rect 9129 -18556 9163 -18522
rect 9197 -18556 9231 -18522
rect 9265 -18556 9299 -18522
rect 9333 -18556 9367 -18522
rect 9401 -18556 9435 -18522
rect 9469 -18539 9694 -18522
rect 9752 -18522 10712 -18484
rect 9752 -18539 9977 -18522
rect 9469 -18556 9508 -18539
rect 8920 -18572 9508 -18556
rect 9938 -18556 9977 -18539
rect 10011 -18556 10045 -18522
rect 10079 -18556 10113 -18522
rect 10147 -18556 10181 -18522
rect 10215 -18556 10249 -18522
rect 10283 -18556 10317 -18522
rect 10351 -18556 10385 -18522
rect 10419 -18556 10453 -18522
rect 10487 -18539 10712 -18522
rect 10770 -18522 11730 -18484
rect 10770 -18539 10995 -18522
rect 10487 -18556 10526 -18539
rect 9938 -18572 10526 -18556
rect 10956 -18556 10995 -18539
rect 11029 -18556 11063 -18522
rect 11097 -18556 11131 -18522
rect 11165 -18556 11199 -18522
rect 11233 -18556 11267 -18522
rect 11301 -18556 11335 -18522
rect 11369 -18556 11403 -18522
rect 11437 -18556 11471 -18522
rect 11505 -18539 11730 -18522
rect 11788 -18522 12748 -18484
rect 11788 -18539 12013 -18522
rect 11505 -18556 11544 -18539
rect 10956 -18572 11544 -18556
rect 11974 -18556 12013 -18539
rect 12047 -18556 12081 -18522
rect 12115 -18556 12149 -18522
rect 12183 -18556 12217 -18522
rect 12251 -18556 12285 -18522
rect 12319 -18556 12353 -18522
rect 12387 -18556 12421 -18522
rect 12455 -18556 12489 -18522
rect 12523 -18539 12748 -18522
rect 12806 -18522 13766 -18484
rect 12806 -18539 13031 -18522
rect 12523 -18556 12562 -18539
rect 11974 -18572 12562 -18556
rect 12992 -18556 13031 -18539
rect 13065 -18556 13099 -18522
rect 13133 -18556 13167 -18522
rect 13201 -18556 13235 -18522
rect 13269 -18556 13303 -18522
rect 13337 -18556 13371 -18522
rect 13405 -18556 13439 -18522
rect 13473 -18556 13507 -18522
rect 13541 -18539 13766 -18522
rect 13824 -18522 14784 -18484
rect 13824 -18539 14049 -18522
rect 13541 -18556 13580 -18539
rect 12992 -18572 13580 -18556
rect 14010 -18556 14049 -18539
rect 14083 -18556 14117 -18522
rect 14151 -18556 14185 -18522
rect 14219 -18556 14253 -18522
rect 14287 -18556 14321 -18522
rect 14355 -18556 14389 -18522
rect 14423 -18556 14457 -18522
rect 14491 -18556 14525 -18522
rect 14559 -18539 14784 -18522
rect 14842 -18522 15802 -18484
rect 14842 -18539 15067 -18522
rect 14559 -18556 14598 -18539
rect 14010 -18572 14598 -18556
rect 15028 -18556 15067 -18539
rect 15101 -18556 15135 -18522
rect 15169 -18556 15203 -18522
rect 15237 -18556 15271 -18522
rect 15305 -18556 15339 -18522
rect 15373 -18556 15407 -18522
rect 15441 -18556 15475 -18522
rect 15509 -18556 15543 -18522
rect 15577 -18539 15802 -18522
rect 15860 -18522 16820 -18484
rect 15860 -18539 16085 -18522
rect 15577 -18556 15616 -18539
rect 15028 -18572 15616 -18556
rect 16046 -18556 16085 -18539
rect 16119 -18556 16153 -18522
rect 16187 -18556 16221 -18522
rect 16255 -18556 16289 -18522
rect 16323 -18556 16357 -18522
rect 16391 -18556 16425 -18522
rect 16459 -18556 16493 -18522
rect 16527 -18556 16561 -18522
rect 16595 -18539 16820 -18522
rect 16878 -18522 17838 -18484
rect 16878 -18539 17103 -18522
rect 16595 -18556 16634 -18539
rect 16046 -18572 16634 -18556
rect 17064 -18556 17103 -18539
rect 17137 -18556 17171 -18522
rect 17205 -18556 17239 -18522
rect 17273 -18556 17307 -18522
rect 17341 -18556 17375 -18522
rect 17409 -18556 17443 -18522
rect 17477 -18556 17511 -18522
rect 17545 -18556 17579 -18522
rect 17613 -18539 17838 -18522
rect 17896 -18522 18856 -18484
rect 17896 -18539 18121 -18522
rect 17613 -18556 17652 -18539
rect 17064 -18572 17652 -18556
rect 18082 -18556 18121 -18539
rect 18155 -18556 18189 -18522
rect 18223 -18556 18257 -18522
rect 18291 -18556 18325 -18522
rect 18359 -18556 18393 -18522
rect 18427 -18556 18461 -18522
rect 18495 -18556 18529 -18522
rect 18563 -18556 18597 -18522
rect 18631 -18539 18856 -18522
rect 18914 -18522 19874 -18484
rect 18914 -18539 19139 -18522
rect 18631 -18556 18670 -18539
rect 18082 -18572 18670 -18556
rect 19100 -18556 19139 -18539
rect 19173 -18556 19207 -18522
rect 19241 -18556 19275 -18522
rect 19309 -18556 19343 -18522
rect 19377 -18556 19411 -18522
rect 19445 -18556 19479 -18522
rect 19513 -18556 19547 -18522
rect 19581 -18556 19615 -18522
rect 19649 -18539 19874 -18522
rect 19932 -18522 20892 -18484
rect 19932 -18539 20157 -18522
rect 19649 -18556 19688 -18539
rect 19100 -18572 19688 -18556
rect 20118 -18556 20157 -18539
rect 20191 -18556 20225 -18522
rect 20259 -18556 20293 -18522
rect 20327 -18556 20361 -18522
rect 20395 -18556 20429 -18522
rect 20463 -18556 20497 -18522
rect 20531 -18556 20565 -18522
rect 20599 -18556 20633 -18522
rect 20667 -18539 20892 -18522
rect 20950 -18522 21910 -18484
rect 20950 -18539 21175 -18522
rect 20667 -18556 20706 -18539
rect 20118 -18572 20706 -18556
rect 21136 -18556 21175 -18539
rect 21209 -18556 21243 -18522
rect 21277 -18556 21311 -18522
rect 21345 -18556 21379 -18522
rect 21413 -18556 21447 -18522
rect 21481 -18556 21515 -18522
rect 21549 -18556 21583 -18522
rect 21617 -18556 21651 -18522
rect 21685 -18539 21910 -18522
rect 21968 -18522 22928 -18484
rect 21968 -18539 22193 -18522
rect 21685 -18556 21724 -18539
rect 21136 -18572 21724 -18556
rect 22154 -18556 22193 -18539
rect 22227 -18556 22261 -18522
rect 22295 -18556 22329 -18522
rect 22363 -18556 22397 -18522
rect 22431 -18556 22465 -18522
rect 22499 -18556 22533 -18522
rect 22567 -18556 22601 -18522
rect 22635 -18556 22669 -18522
rect 22703 -18539 22928 -18522
rect 22703 -18556 22742 -18539
rect 22154 -18572 22742 -18556
rect -9138 -18876 -8178 -18838
rect -9138 -18893 -8913 -18876
rect -8952 -18910 -8913 -18893
rect -8879 -18910 -8845 -18876
rect -8811 -18910 -8777 -18876
rect -8743 -18910 -8709 -18876
rect -8675 -18910 -8641 -18876
rect -8607 -18910 -8573 -18876
rect -8539 -18910 -8505 -18876
rect -8471 -18910 -8437 -18876
rect -8403 -18893 -8178 -18876
rect -8120 -18876 -7160 -18838
rect -8120 -18893 -7895 -18876
rect -8403 -18910 -8364 -18893
rect -8952 -18926 -8364 -18910
rect -7934 -18910 -7895 -18893
rect -7861 -18910 -7827 -18876
rect -7793 -18910 -7759 -18876
rect -7725 -18910 -7691 -18876
rect -7657 -18910 -7623 -18876
rect -7589 -18910 -7555 -18876
rect -7521 -18910 -7487 -18876
rect -7453 -18910 -7419 -18876
rect -7385 -18893 -7160 -18876
rect -7102 -18876 -6142 -18838
rect -7102 -18893 -6877 -18876
rect -7385 -18910 -7346 -18893
rect -7934 -18926 -7346 -18910
rect -6916 -18910 -6877 -18893
rect -6843 -18910 -6809 -18876
rect -6775 -18910 -6741 -18876
rect -6707 -18910 -6673 -18876
rect -6639 -18910 -6605 -18876
rect -6571 -18910 -6537 -18876
rect -6503 -18910 -6469 -18876
rect -6435 -18910 -6401 -18876
rect -6367 -18893 -6142 -18876
rect -6084 -18876 -5124 -18838
rect -6084 -18893 -5859 -18876
rect -6367 -18910 -6328 -18893
rect -6916 -18926 -6328 -18910
rect -5898 -18910 -5859 -18893
rect -5825 -18910 -5791 -18876
rect -5757 -18910 -5723 -18876
rect -5689 -18910 -5655 -18876
rect -5621 -18910 -5587 -18876
rect -5553 -18910 -5519 -18876
rect -5485 -18910 -5451 -18876
rect -5417 -18910 -5383 -18876
rect -5349 -18893 -5124 -18876
rect -5066 -18876 -4106 -18838
rect -5066 -18893 -4841 -18876
rect -5349 -18910 -5310 -18893
rect -5898 -18926 -5310 -18910
rect -4880 -18910 -4841 -18893
rect -4807 -18910 -4773 -18876
rect -4739 -18910 -4705 -18876
rect -4671 -18910 -4637 -18876
rect -4603 -18910 -4569 -18876
rect -4535 -18910 -4501 -18876
rect -4467 -18910 -4433 -18876
rect -4399 -18910 -4365 -18876
rect -4331 -18893 -4106 -18876
rect -4048 -18876 -3088 -18838
rect -4048 -18893 -3823 -18876
rect -4331 -18910 -4292 -18893
rect -4880 -18926 -4292 -18910
rect -3862 -18910 -3823 -18893
rect -3789 -18910 -3755 -18876
rect -3721 -18910 -3687 -18876
rect -3653 -18910 -3619 -18876
rect -3585 -18910 -3551 -18876
rect -3517 -18910 -3483 -18876
rect -3449 -18910 -3415 -18876
rect -3381 -18910 -3347 -18876
rect -3313 -18893 -3088 -18876
rect -3030 -18876 -2070 -18838
rect -3030 -18893 -2805 -18876
rect -3313 -18910 -3274 -18893
rect -3862 -18926 -3274 -18910
rect -2844 -18910 -2805 -18893
rect -2771 -18910 -2737 -18876
rect -2703 -18910 -2669 -18876
rect -2635 -18910 -2601 -18876
rect -2567 -18910 -2533 -18876
rect -2499 -18910 -2465 -18876
rect -2431 -18910 -2397 -18876
rect -2363 -18910 -2329 -18876
rect -2295 -18893 -2070 -18876
rect -2012 -18876 -1052 -18838
rect -2012 -18893 -1787 -18876
rect -2295 -18910 -2256 -18893
rect -2844 -18926 -2256 -18910
rect -1826 -18910 -1787 -18893
rect -1753 -18910 -1719 -18876
rect -1685 -18910 -1651 -18876
rect -1617 -18910 -1583 -18876
rect -1549 -18910 -1515 -18876
rect -1481 -18910 -1447 -18876
rect -1413 -18910 -1379 -18876
rect -1345 -18910 -1311 -18876
rect -1277 -18893 -1052 -18876
rect -994 -18876 -34 -18838
rect -994 -18893 -769 -18876
rect -1277 -18910 -1238 -18893
rect -1826 -18926 -1238 -18910
rect -808 -18910 -769 -18893
rect -735 -18910 -701 -18876
rect -667 -18910 -633 -18876
rect -599 -18910 -565 -18876
rect -531 -18910 -497 -18876
rect -463 -18910 -429 -18876
rect -395 -18910 -361 -18876
rect -327 -18910 -293 -18876
rect -259 -18893 -34 -18876
rect -259 -18910 -220 -18893
rect -808 -18926 -220 -18910
rect 2812 -19046 3400 -19030
rect 2812 -19063 2851 -19046
rect 2626 -19080 2851 -19063
rect 2885 -19080 2919 -19046
rect 2953 -19080 2987 -19046
rect 3021 -19080 3055 -19046
rect 3089 -19080 3123 -19046
rect 3157 -19080 3191 -19046
rect 3225 -19080 3259 -19046
rect 3293 -19080 3327 -19046
rect 3361 -19063 3400 -19046
rect 3830 -19046 4418 -19030
rect 3830 -19063 3869 -19046
rect 3361 -19080 3586 -19063
rect 2626 -19118 3586 -19080
rect 3644 -19080 3869 -19063
rect 3903 -19080 3937 -19046
rect 3971 -19080 4005 -19046
rect 4039 -19080 4073 -19046
rect 4107 -19080 4141 -19046
rect 4175 -19080 4209 -19046
rect 4243 -19080 4277 -19046
rect 4311 -19080 4345 -19046
rect 4379 -19063 4418 -19046
rect 4848 -19046 5436 -19030
rect 4848 -19063 4887 -19046
rect 4379 -19080 4604 -19063
rect 3644 -19118 4604 -19080
rect 4662 -19080 4887 -19063
rect 4921 -19080 4955 -19046
rect 4989 -19080 5023 -19046
rect 5057 -19080 5091 -19046
rect 5125 -19080 5159 -19046
rect 5193 -19080 5227 -19046
rect 5261 -19080 5295 -19046
rect 5329 -19080 5363 -19046
rect 5397 -19063 5436 -19046
rect 5866 -19046 6454 -19030
rect 5866 -19063 5905 -19046
rect 5397 -19080 5622 -19063
rect 4662 -19118 5622 -19080
rect 5680 -19080 5905 -19063
rect 5939 -19080 5973 -19046
rect 6007 -19080 6041 -19046
rect 6075 -19080 6109 -19046
rect 6143 -19080 6177 -19046
rect 6211 -19080 6245 -19046
rect 6279 -19080 6313 -19046
rect 6347 -19080 6381 -19046
rect 6415 -19063 6454 -19046
rect 6884 -19046 7472 -19030
rect 6884 -19063 6923 -19046
rect 6415 -19080 6640 -19063
rect 5680 -19118 6640 -19080
rect 6698 -19080 6923 -19063
rect 6957 -19080 6991 -19046
rect 7025 -19080 7059 -19046
rect 7093 -19080 7127 -19046
rect 7161 -19080 7195 -19046
rect 7229 -19080 7263 -19046
rect 7297 -19080 7331 -19046
rect 7365 -19080 7399 -19046
rect 7433 -19063 7472 -19046
rect 7902 -19046 8490 -19030
rect 7902 -19063 7941 -19046
rect 7433 -19080 7658 -19063
rect 6698 -19118 7658 -19080
rect 7716 -19080 7941 -19063
rect 7975 -19080 8009 -19046
rect 8043 -19080 8077 -19046
rect 8111 -19080 8145 -19046
rect 8179 -19080 8213 -19046
rect 8247 -19080 8281 -19046
rect 8315 -19080 8349 -19046
rect 8383 -19080 8417 -19046
rect 8451 -19063 8490 -19046
rect 8920 -19046 9508 -19030
rect 8920 -19063 8959 -19046
rect 8451 -19080 8676 -19063
rect 7716 -19118 8676 -19080
rect 8734 -19080 8959 -19063
rect 8993 -19080 9027 -19046
rect 9061 -19080 9095 -19046
rect 9129 -19080 9163 -19046
rect 9197 -19080 9231 -19046
rect 9265 -19080 9299 -19046
rect 9333 -19080 9367 -19046
rect 9401 -19080 9435 -19046
rect 9469 -19063 9508 -19046
rect 9938 -19046 10526 -19030
rect 9938 -19063 9977 -19046
rect 9469 -19080 9694 -19063
rect 8734 -19118 9694 -19080
rect 9752 -19080 9977 -19063
rect 10011 -19080 10045 -19046
rect 10079 -19080 10113 -19046
rect 10147 -19080 10181 -19046
rect 10215 -19080 10249 -19046
rect 10283 -19080 10317 -19046
rect 10351 -19080 10385 -19046
rect 10419 -19080 10453 -19046
rect 10487 -19063 10526 -19046
rect 10956 -19046 11544 -19030
rect 10956 -19063 10995 -19046
rect 10487 -19080 10712 -19063
rect 9752 -19118 10712 -19080
rect 10770 -19080 10995 -19063
rect 11029 -19080 11063 -19046
rect 11097 -19080 11131 -19046
rect 11165 -19080 11199 -19046
rect 11233 -19080 11267 -19046
rect 11301 -19080 11335 -19046
rect 11369 -19080 11403 -19046
rect 11437 -19080 11471 -19046
rect 11505 -19063 11544 -19046
rect 11974 -19046 12562 -19030
rect 11974 -19063 12013 -19046
rect 11505 -19080 11730 -19063
rect 10770 -19118 11730 -19080
rect 11788 -19080 12013 -19063
rect 12047 -19080 12081 -19046
rect 12115 -19080 12149 -19046
rect 12183 -19080 12217 -19046
rect 12251 -19080 12285 -19046
rect 12319 -19080 12353 -19046
rect 12387 -19080 12421 -19046
rect 12455 -19080 12489 -19046
rect 12523 -19063 12562 -19046
rect 12992 -19046 13580 -19030
rect 12992 -19063 13031 -19046
rect 12523 -19080 12748 -19063
rect 11788 -19118 12748 -19080
rect 12806 -19080 13031 -19063
rect 13065 -19080 13099 -19046
rect 13133 -19080 13167 -19046
rect 13201 -19080 13235 -19046
rect 13269 -19080 13303 -19046
rect 13337 -19080 13371 -19046
rect 13405 -19080 13439 -19046
rect 13473 -19080 13507 -19046
rect 13541 -19063 13580 -19046
rect 14010 -19046 14598 -19030
rect 14010 -19063 14049 -19046
rect 13541 -19080 13766 -19063
rect 12806 -19118 13766 -19080
rect 13824 -19080 14049 -19063
rect 14083 -19080 14117 -19046
rect 14151 -19080 14185 -19046
rect 14219 -19080 14253 -19046
rect 14287 -19080 14321 -19046
rect 14355 -19080 14389 -19046
rect 14423 -19080 14457 -19046
rect 14491 -19080 14525 -19046
rect 14559 -19063 14598 -19046
rect 15028 -19046 15616 -19030
rect 15028 -19063 15067 -19046
rect 14559 -19080 14784 -19063
rect 13824 -19118 14784 -19080
rect 14842 -19080 15067 -19063
rect 15101 -19080 15135 -19046
rect 15169 -19080 15203 -19046
rect 15237 -19080 15271 -19046
rect 15305 -19080 15339 -19046
rect 15373 -19080 15407 -19046
rect 15441 -19080 15475 -19046
rect 15509 -19080 15543 -19046
rect 15577 -19063 15616 -19046
rect 16046 -19046 16634 -19030
rect 16046 -19063 16085 -19046
rect 15577 -19080 15802 -19063
rect 14842 -19118 15802 -19080
rect 15860 -19080 16085 -19063
rect 16119 -19080 16153 -19046
rect 16187 -19080 16221 -19046
rect 16255 -19080 16289 -19046
rect 16323 -19080 16357 -19046
rect 16391 -19080 16425 -19046
rect 16459 -19080 16493 -19046
rect 16527 -19080 16561 -19046
rect 16595 -19063 16634 -19046
rect 17064 -19046 17652 -19030
rect 17064 -19063 17103 -19046
rect 16595 -19080 16820 -19063
rect 15860 -19118 16820 -19080
rect 16878 -19080 17103 -19063
rect 17137 -19080 17171 -19046
rect 17205 -19080 17239 -19046
rect 17273 -19080 17307 -19046
rect 17341 -19080 17375 -19046
rect 17409 -19080 17443 -19046
rect 17477 -19080 17511 -19046
rect 17545 -19080 17579 -19046
rect 17613 -19063 17652 -19046
rect 18082 -19046 18670 -19030
rect 18082 -19063 18121 -19046
rect 17613 -19080 17838 -19063
rect 16878 -19118 17838 -19080
rect 17896 -19080 18121 -19063
rect 18155 -19080 18189 -19046
rect 18223 -19080 18257 -19046
rect 18291 -19080 18325 -19046
rect 18359 -19080 18393 -19046
rect 18427 -19080 18461 -19046
rect 18495 -19080 18529 -19046
rect 18563 -19080 18597 -19046
rect 18631 -19063 18670 -19046
rect 19100 -19046 19688 -19030
rect 19100 -19063 19139 -19046
rect 18631 -19080 18856 -19063
rect 17896 -19118 18856 -19080
rect 18914 -19080 19139 -19063
rect 19173 -19080 19207 -19046
rect 19241 -19080 19275 -19046
rect 19309 -19080 19343 -19046
rect 19377 -19080 19411 -19046
rect 19445 -19080 19479 -19046
rect 19513 -19080 19547 -19046
rect 19581 -19080 19615 -19046
rect 19649 -19063 19688 -19046
rect 20118 -19046 20706 -19030
rect 20118 -19063 20157 -19046
rect 19649 -19080 19874 -19063
rect 18914 -19118 19874 -19080
rect 19932 -19080 20157 -19063
rect 20191 -19080 20225 -19046
rect 20259 -19080 20293 -19046
rect 20327 -19080 20361 -19046
rect 20395 -19080 20429 -19046
rect 20463 -19080 20497 -19046
rect 20531 -19080 20565 -19046
rect 20599 -19080 20633 -19046
rect 20667 -19063 20706 -19046
rect 21136 -19046 21724 -19030
rect 21136 -19063 21175 -19046
rect 20667 -19080 20892 -19063
rect 19932 -19118 20892 -19080
rect 20950 -19080 21175 -19063
rect 21209 -19080 21243 -19046
rect 21277 -19080 21311 -19046
rect 21345 -19080 21379 -19046
rect 21413 -19080 21447 -19046
rect 21481 -19080 21515 -19046
rect 21549 -19080 21583 -19046
rect 21617 -19080 21651 -19046
rect 21685 -19063 21724 -19046
rect 22154 -19046 22742 -19030
rect 22154 -19063 22193 -19046
rect 21685 -19080 21910 -19063
rect 20950 -19118 21910 -19080
rect 21968 -19080 22193 -19063
rect 22227 -19080 22261 -19046
rect 22295 -19080 22329 -19046
rect 22363 -19080 22397 -19046
rect 22431 -19080 22465 -19046
rect 22499 -19080 22533 -19046
rect 22567 -19080 22601 -19046
rect 22635 -19080 22669 -19046
rect 22703 -19063 22742 -19046
rect 22703 -19080 22928 -19063
rect 21968 -19118 22928 -19080
rect -2252 -19550 -2144 -19534
rect -2252 -19567 -2215 -19550
rect -2278 -19584 -2215 -19567
rect -2181 -19567 -2144 -19550
rect -2034 -19550 -1926 -19534
rect -2034 -19567 -1997 -19550
rect -2181 -19584 -2118 -19567
rect -2278 -19622 -2118 -19584
rect -2060 -19584 -1997 -19567
rect -1963 -19567 -1926 -19550
rect -1816 -19550 -1708 -19534
rect -1816 -19567 -1779 -19550
rect -1963 -19584 -1900 -19567
rect -2060 -19622 -1900 -19584
rect -1842 -19584 -1779 -19567
rect -1745 -19567 -1708 -19550
rect -1598 -19550 -1490 -19534
rect -1598 -19567 -1561 -19550
rect -1745 -19584 -1682 -19567
rect -1842 -19622 -1682 -19584
rect -1624 -19584 -1561 -19567
rect -1527 -19567 -1490 -19550
rect -1380 -19550 -1272 -19534
rect -1380 -19567 -1343 -19550
rect -1527 -19584 -1464 -19567
rect -1624 -19622 -1464 -19584
rect -1406 -19584 -1343 -19567
rect -1309 -19567 -1272 -19550
rect -1162 -19550 -1054 -19534
rect -1162 -19567 -1125 -19550
rect -1309 -19584 -1246 -19567
rect -1406 -19622 -1246 -19584
rect -1188 -19584 -1125 -19567
rect -1091 -19567 -1054 -19550
rect -944 -19550 -836 -19534
rect -944 -19567 -907 -19550
rect -1091 -19584 -1028 -19567
rect -1188 -19622 -1028 -19584
rect -970 -19584 -907 -19567
rect -873 -19567 -836 -19550
rect -726 -19550 -618 -19534
rect -726 -19567 -689 -19550
rect -873 -19584 -810 -19567
rect -970 -19622 -810 -19584
rect -752 -19584 -689 -19567
rect -655 -19567 -618 -19550
rect -508 -19550 -400 -19534
rect -508 -19567 -471 -19550
rect -655 -19584 -592 -19567
rect -752 -19622 -592 -19584
rect -534 -19584 -471 -19567
rect -437 -19567 -400 -19550
rect -290 -19550 -182 -19534
rect -290 -19567 -253 -19550
rect -437 -19584 -374 -19567
rect -534 -19622 -374 -19584
rect -316 -19584 -253 -19567
rect -219 -19567 -182 -19550
rect -219 -19584 -156 -19567
rect -316 -19622 -156 -19584
rect 2626 -19756 3586 -19718
rect 2626 -19773 2851 -19756
rect 2812 -19790 2851 -19773
rect 2885 -19790 2919 -19756
rect 2953 -19790 2987 -19756
rect 3021 -19790 3055 -19756
rect 3089 -19790 3123 -19756
rect 3157 -19790 3191 -19756
rect 3225 -19790 3259 -19756
rect 3293 -19790 3327 -19756
rect 3361 -19773 3586 -19756
rect 3644 -19756 4604 -19718
rect 3644 -19773 3869 -19756
rect 3361 -19790 3400 -19773
rect 2812 -19806 3400 -19790
rect 3830 -19790 3869 -19773
rect 3903 -19790 3937 -19756
rect 3971 -19790 4005 -19756
rect 4039 -19790 4073 -19756
rect 4107 -19790 4141 -19756
rect 4175 -19790 4209 -19756
rect 4243 -19790 4277 -19756
rect 4311 -19790 4345 -19756
rect 4379 -19773 4604 -19756
rect 4662 -19756 5622 -19718
rect 4662 -19773 4887 -19756
rect 4379 -19790 4418 -19773
rect 3830 -19806 4418 -19790
rect 4848 -19790 4887 -19773
rect 4921 -19790 4955 -19756
rect 4989 -19790 5023 -19756
rect 5057 -19790 5091 -19756
rect 5125 -19790 5159 -19756
rect 5193 -19790 5227 -19756
rect 5261 -19790 5295 -19756
rect 5329 -19790 5363 -19756
rect 5397 -19773 5622 -19756
rect 5680 -19756 6640 -19718
rect 5680 -19773 5905 -19756
rect 5397 -19790 5436 -19773
rect 4848 -19806 5436 -19790
rect 5866 -19790 5905 -19773
rect 5939 -19790 5973 -19756
rect 6007 -19790 6041 -19756
rect 6075 -19790 6109 -19756
rect 6143 -19790 6177 -19756
rect 6211 -19790 6245 -19756
rect 6279 -19790 6313 -19756
rect 6347 -19790 6381 -19756
rect 6415 -19773 6640 -19756
rect 6698 -19756 7658 -19718
rect 6698 -19773 6923 -19756
rect 6415 -19790 6454 -19773
rect 5866 -19806 6454 -19790
rect 6884 -19790 6923 -19773
rect 6957 -19790 6991 -19756
rect 7025 -19790 7059 -19756
rect 7093 -19790 7127 -19756
rect 7161 -19790 7195 -19756
rect 7229 -19790 7263 -19756
rect 7297 -19790 7331 -19756
rect 7365 -19790 7399 -19756
rect 7433 -19773 7658 -19756
rect 7716 -19756 8676 -19718
rect 7716 -19773 7941 -19756
rect 7433 -19790 7472 -19773
rect 6884 -19806 7472 -19790
rect 7902 -19790 7941 -19773
rect 7975 -19790 8009 -19756
rect 8043 -19790 8077 -19756
rect 8111 -19790 8145 -19756
rect 8179 -19790 8213 -19756
rect 8247 -19790 8281 -19756
rect 8315 -19790 8349 -19756
rect 8383 -19790 8417 -19756
rect 8451 -19773 8676 -19756
rect 8734 -19756 9694 -19718
rect 8734 -19773 8959 -19756
rect 8451 -19790 8490 -19773
rect 7902 -19806 8490 -19790
rect 8920 -19790 8959 -19773
rect 8993 -19790 9027 -19756
rect 9061 -19790 9095 -19756
rect 9129 -19790 9163 -19756
rect 9197 -19790 9231 -19756
rect 9265 -19790 9299 -19756
rect 9333 -19790 9367 -19756
rect 9401 -19790 9435 -19756
rect 9469 -19773 9694 -19756
rect 9752 -19756 10712 -19718
rect 9752 -19773 9977 -19756
rect 9469 -19790 9508 -19773
rect 8920 -19806 9508 -19790
rect 9938 -19790 9977 -19773
rect 10011 -19790 10045 -19756
rect 10079 -19790 10113 -19756
rect 10147 -19790 10181 -19756
rect 10215 -19790 10249 -19756
rect 10283 -19790 10317 -19756
rect 10351 -19790 10385 -19756
rect 10419 -19790 10453 -19756
rect 10487 -19773 10712 -19756
rect 10770 -19756 11730 -19718
rect 10770 -19773 10995 -19756
rect 10487 -19790 10526 -19773
rect 9938 -19806 10526 -19790
rect 10956 -19790 10995 -19773
rect 11029 -19790 11063 -19756
rect 11097 -19790 11131 -19756
rect 11165 -19790 11199 -19756
rect 11233 -19790 11267 -19756
rect 11301 -19790 11335 -19756
rect 11369 -19790 11403 -19756
rect 11437 -19790 11471 -19756
rect 11505 -19773 11730 -19756
rect 11788 -19756 12748 -19718
rect 11788 -19773 12013 -19756
rect 11505 -19790 11544 -19773
rect 10956 -19806 11544 -19790
rect 11974 -19790 12013 -19773
rect 12047 -19790 12081 -19756
rect 12115 -19790 12149 -19756
rect 12183 -19790 12217 -19756
rect 12251 -19790 12285 -19756
rect 12319 -19790 12353 -19756
rect 12387 -19790 12421 -19756
rect 12455 -19790 12489 -19756
rect 12523 -19773 12748 -19756
rect 12806 -19756 13766 -19718
rect 12806 -19773 13031 -19756
rect 12523 -19790 12562 -19773
rect 11974 -19806 12562 -19790
rect 12992 -19790 13031 -19773
rect 13065 -19790 13099 -19756
rect 13133 -19790 13167 -19756
rect 13201 -19790 13235 -19756
rect 13269 -19790 13303 -19756
rect 13337 -19790 13371 -19756
rect 13405 -19790 13439 -19756
rect 13473 -19790 13507 -19756
rect 13541 -19773 13766 -19756
rect 13824 -19756 14784 -19718
rect 13824 -19773 14049 -19756
rect 13541 -19790 13580 -19773
rect 12992 -19806 13580 -19790
rect 14010 -19790 14049 -19773
rect 14083 -19790 14117 -19756
rect 14151 -19790 14185 -19756
rect 14219 -19790 14253 -19756
rect 14287 -19790 14321 -19756
rect 14355 -19790 14389 -19756
rect 14423 -19790 14457 -19756
rect 14491 -19790 14525 -19756
rect 14559 -19773 14784 -19756
rect 14842 -19756 15802 -19718
rect 14842 -19773 15067 -19756
rect 14559 -19790 14598 -19773
rect 14010 -19806 14598 -19790
rect 15028 -19790 15067 -19773
rect 15101 -19790 15135 -19756
rect 15169 -19790 15203 -19756
rect 15237 -19790 15271 -19756
rect 15305 -19790 15339 -19756
rect 15373 -19790 15407 -19756
rect 15441 -19790 15475 -19756
rect 15509 -19790 15543 -19756
rect 15577 -19773 15802 -19756
rect 15860 -19756 16820 -19718
rect 15860 -19773 16085 -19756
rect 15577 -19790 15616 -19773
rect 15028 -19806 15616 -19790
rect 16046 -19790 16085 -19773
rect 16119 -19790 16153 -19756
rect 16187 -19790 16221 -19756
rect 16255 -19790 16289 -19756
rect 16323 -19790 16357 -19756
rect 16391 -19790 16425 -19756
rect 16459 -19790 16493 -19756
rect 16527 -19790 16561 -19756
rect 16595 -19773 16820 -19756
rect 16878 -19756 17838 -19718
rect 16878 -19773 17103 -19756
rect 16595 -19790 16634 -19773
rect 16046 -19806 16634 -19790
rect 17064 -19790 17103 -19773
rect 17137 -19790 17171 -19756
rect 17205 -19790 17239 -19756
rect 17273 -19790 17307 -19756
rect 17341 -19790 17375 -19756
rect 17409 -19790 17443 -19756
rect 17477 -19790 17511 -19756
rect 17545 -19790 17579 -19756
rect 17613 -19773 17838 -19756
rect 17896 -19756 18856 -19718
rect 17896 -19773 18121 -19756
rect 17613 -19790 17652 -19773
rect 17064 -19806 17652 -19790
rect 18082 -19790 18121 -19773
rect 18155 -19790 18189 -19756
rect 18223 -19790 18257 -19756
rect 18291 -19790 18325 -19756
rect 18359 -19790 18393 -19756
rect 18427 -19790 18461 -19756
rect 18495 -19790 18529 -19756
rect 18563 -19790 18597 -19756
rect 18631 -19773 18856 -19756
rect 18914 -19756 19874 -19718
rect 18914 -19773 19139 -19756
rect 18631 -19790 18670 -19773
rect 18082 -19806 18670 -19790
rect 19100 -19790 19139 -19773
rect 19173 -19790 19207 -19756
rect 19241 -19790 19275 -19756
rect 19309 -19790 19343 -19756
rect 19377 -19790 19411 -19756
rect 19445 -19790 19479 -19756
rect 19513 -19790 19547 -19756
rect 19581 -19790 19615 -19756
rect 19649 -19773 19874 -19756
rect 19932 -19756 20892 -19718
rect 19932 -19773 20157 -19756
rect 19649 -19790 19688 -19773
rect 19100 -19806 19688 -19790
rect 20118 -19790 20157 -19773
rect 20191 -19790 20225 -19756
rect 20259 -19790 20293 -19756
rect 20327 -19790 20361 -19756
rect 20395 -19790 20429 -19756
rect 20463 -19790 20497 -19756
rect 20531 -19790 20565 -19756
rect 20599 -19790 20633 -19756
rect 20667 -19773 20892 -19756
rect 20950 -19756 21910 -19718
rect 20950 -19773 21175 -19756
rect 20667 -19790 20706 -19773
rect 20118 -19806 20706 -19790
rect 21136 -19790 21175 -19773
rect 21209 -19790 21243 -19756
rect 21277 -19790 21311 -19756
rect 21345 -19790 21379 -19756
rect 21413 -19790 21447 -19756
rect 21481 -19790 21515 -19756
rect 21549 -19790 21583 -19756
rect 21617 -19790 21651 -19756
rect 21685 -19773 21910 -19756
rect 21968 -19756 22928 -19718
rect 21968 -19773 22193 -19756
rect 21685 -19790 21724 -19773
rect 21136 -19806 21724 -19790
rect 22154 -19790 22193 -19773
rect 22227 -19790 22261 -19756
rect 22295 -19790 22329 -19756
rect 22363 -19790 22397 -19756
rect 22431 -19790 22465 -19756
rect 22499 -19790 22533 -19756
rect 22567 -19790 22601 -19756
rect 22635 -19790 22669 -19756
rect 22703 -19773 22928 -19756
rect 22703 -19790 22742 -19773
rect 22154 -19806 22742 -19790
rect -2278 -19860 -2118 -19822
rect -2278 -19877 -2215 -19860
rect -2252 -19894 -2215 -19877
rect -2181 -19877 -2118 -19860
rect -2060 -19860 -1900 -19822
rect -2060 -19877 -1997 -19860
rect -2181 -19894 -2144 -19877
rect -2252 -19910 -2144 -19894
rect -2034 -19894 -1997 -19877
rect -1963 -19877 -1900 -19860
rect -1842 -19860 -1682 -19822
rect -1842 -19877 -1779 -19860
rect -1963 -19894 -1926 -19877
rect -2034 -19910 -1926 -19894
rect -1816 -19894 -1779 -19877
rect -1745 -19877 -1682 -19860
rect -1624 -19860 -1464 -19822
rect -1624 -19877 -1561 -19860
rect -1745 -19894 -1708 -19877
rect -1816 -19910 -1708 -19894
rect -1598 -19894 -1561 -19877
rect -1527 -19877 -1464 -19860
rect -1406 -19860 -1246 -19822
rect -1406 -19877 -1343 -19860
rect -1527 -19894 -1490 -19877
rect -1598 -19910 -1490 -19894
rect -1380 -19894 -1343 -19877
rect -1309 -19877 -1246 -19860
rect -1188 -19860 -1028 -19822
rect -1188 -19877 -1125 -19860
rect -1309 -19894 -1272 -19877
rect -1380 -19910 -1272 -19894
rect -1162 -19894 -1125 -19877
rect -1091 -19877 -1028 -19860
rect -970 -19860 -810 -19822
rect -970 -19877 -907 -19860
rect -1091 -19894 -1054 -19877
rect -1162 -19910 -1054 -19894
rect -944 -19894 -907 -19877
rect -873 -19877 -810 -19860
rect -752 -19860 -592 -19822
rect -752 -19877 -689 -19860
rect -873 -19894 -836 -19877
rect -944 -19910 -836 -19894
rect -726 -19894 -689 -19877
rect -655 -19877 -592 -19860
rect -534 -19860 -374 -19822
rect -534 -19877 -471 -19860
rect -655 -19894 -618 -19877
rect -726 -19910 -618 -19894
rect -508 -19894 -471 -19877
rect -437 -19877 -374 -19860
rect -316 -19860 -156 -19822
rect -316 -19877 -253 -19860
rect -437 -19894 -400 -19877
rect -508 -19910 -400 -19894
rect -290 -19894 -253 -19877
rect -219 -19877 -156 -19860
rect -219 -19894 -182 -19877
rect -290 -19910 -182 -19894
rect 2812 -20280 3400 -20264
rect 2812 -20297 2851 -20280
rect 2626 -20314 2851 -20297
rect 2885 -20314 2919 -20280
rect 2953 -20314 2987 -20280
rect 3021 -20314 3055 -20280
rect 3089 -20314 3123 -20280
rect 3157 -20314 3191 -20280
rect 3225 -20314 3259 -20280
rect 3293 -20314 3327 -20280
rect 3361 -20297 3400 -20280
rect 3830 -20280 4418 -20264
rect 3830 -20297 3869 -20280
rect 3361 -20314 3586 -20297
rect 2626 -20352 3586 -20314
rect 3644 -20314 3869 -20297
rect 3903 -20314 3937 -20280
rect 3971 -20314 4005 -20280
rect 4039 -20314 4073 -20280
rect 4107 -20314 4141 -20280
rect 4175 -20314 4209 -20280
rect 4243 -20314 4277 -20280
rect 4311 -20314 4345 -20280
rect 4379 -20297 4418 -20280
rect 4848 -20280 5436 -20264
rect 4848 -20297 4887 -20280
rect 4379 -20314 4604 -20297
rect 3644 -20352 4604 -20314
rect 4662 -20314 4887 -20297
rect 4921 -20314 4955 -20280
rect 4989 -20314 5023 -20280
rect 5057 -20314 5091 -20280
rect 5125 -20314 5159 -20280
rect 5193 -20314 5227 -20280
rect 5261 -20314 5295 -20280
rect 5329 -20314 5363 -20280
rect 5397 -20297 5436 -20280
rect 5866 -20280 6454 -20264
rect 5866 -20297 5905 -20280
rect 5397 -20314 5622 -20297
rect 4662 -20352 5622 -20314
rect 5680 -20314 5905 -20297
rect 5939 -20314 5973 -20280
rect 6007 -20314 6041 -20280
rect 6075 -20314 6109 -20280
rect 6143 -20314 6177 -20280
rect 6211 -20314 6245 -20280
rect 6279 -20314 6313 -20280
rect 6347 -20314 6381 -20280
rect 6415 -20297 6454 -20280
rect 6884 -20280 7472 -20264
rect 6884 -20297 6923 -20280
rect 6415 -20314 6640 -20297
rect 5680 -20352 6640 -20314
rect 6698 -20314 6923 -20297
rect 6957 -20314 6991 -20280
rect 7025 -20314 7059 -20280
rect 7093 -20314 7127 -20280
rect 7161 -20314 7195 -20280
rect 7229 -20314 7263 -20280
rect 7297 -20314 7331 -20280
rect 7365 -20314 7399 -20280
rect 7433 -20297 7472 -20280
rect 7902 -20280 8490 -20264
rect 7902 -20297 7941 -20280
rect 7433 -20314 7658 -20297
rect 6698 -20352 7658 -20314
rect 7716 -20314 7941 -20297
rect 7975 -20314 8009 -20280
rect 8043 -20314 8077 -20280
rect 8111 -20314 8145 -20280
rect 8179 -20314 8213 -20280
rect 8247 -20314 8281 -20280
rect 8315 -20314 8349 -20280
rect 8383 -20314 8417 -20280
rect 8451 -20297 8490 -20280
rect 8920 -20280 9508 -20264
rect 8920 -20297 8959 -20280
rect 8451 -20314 8676 -20297
rect 7716 -20352 8676 -20314
rect 8734 -20314 8959 -20297
rect 8993 -20314 9027 -20280
rect 9061 -20314 9095 -20280
rect 9129 -20314 9163 -20280
rect 9197 -20314 9231 -20280
rect 9265 -20314 9299 -20280
rect 9333 -20314 9367 -20280
rect 9401 -20314 9435 -20280
rect 9469 -20297 9508 -20280
rect 9938 -20280 10526 -20264
rect 9938 -20297 9977 -20280
rect 9469 -20314 9694 -20297
rect 8734 -20352 9694 -20314
rect 9752 -20314 9977 -20297
rect 10011 -20314 10045 -20280
rect 10079 -20314 10113 -20280
rect 10147 -20314 10181 -20280
rect 10215 -20314 10249 -20280
rect 10283 -20314 10317 -20280
rect 10351 -20314 10385 -20280
rect 10419 -20314 10453 -20280
rect 10487 -20297 10526 -20280
rect 10956 -20280 11544 -20264
rect 10956 -20297 10995 -20280
rect 10487 -20314 10712 -20297
rect 9752 -20352 10712 -20314
rect 10770 -20314 10995 -20297
rect 11029 -20314 11063 -20280
rect 11097 -20314 11131 -20280
rect 11165 -20314 11199 -20280
rect 11233 -20314 11267 -20280
rect 11301 -20314 11335 -20280
rect 11369 -20314 11403 -20280
rect 11437 -20314 11471 -20280
rect 11505 -20297 11544 -20280
rect 11974 -20280 12562 -20264
rect 11974 -20297 12013 -20280
rect 11505 -20314 11730 -20297
rect 10770 -20352 11730 -20314
rect 11788 -20314 12013 -20297
rect 12047 -20314 12081 -20280
rect 12115 -20314 12149 -20280
rect 12183 -20314 12217 -20280
rect 12251 -20314 12285 -20280
rect 12319 -20314 12353 -20280
rect 12387 -20314 12421 -20280
rect 12455 -20314 12489 -20280
rect 12523 -20297 12562 -20280
rect 12992 -20280 13580 -20264
rect 12992 -20297 13031 -20280
rect 12523 -20314 12748 -20297
rect 11788 -20352 12748 -20314
rect 12806 -20314 13031 -20297
rect 13065 -20314 13099 -20280
rect 13133 -20314 13167 -20280
rect 13201 -20314 13235 -20280
rect 13269 -20314 13303 -20280
rect 13337 -20314 13371 -20280
rect 13405 -20314 13439 -20280
rect 13473 -20314 13507 -20280
rect 13541 -20297 13580 -20280
rect 14010 -20280 14598 -20264
rect 14010 -20297 14049 -20280
rect 13541 -20314 13766 -20297
rect 12806 -20352 13766 -20314
rect 13824 -20314 14049 -20297
rect 14083 -20314 14117 -20280
rect 14151 -20314 14185 -20280
rect 14219 -20314 14253 -20280
rect 14287 -20314 14321 -20280
rect 14355 -20314 14389 -20280
rect 14423 -20314 14457 -20280
rect 14491 -20314 14525 -20280
rect 14559 -20297 14598 -20280
rect 15028 -20280 15616 -20264
rect 15028 -20297 15067 -20280
rect 14559 -20314 14784 -20297
rect 13824 -20352 14784 -20314
rect 14842 -20314 15067 -20297
rect 15101 -20314 15135 -20280
rect 15169 -20314 15203 -20280
rect 15237 -20314 15271 -20280
rect 15305 -20314 15339 -20280
rect 15373 -20314 15407 -20280
rect 15441 -20314 15475 -20280
rect 15509 -20314 15543 -20280
rect 15577 -20297 15616 -20280
rect 16046 -20280 16634 -20264
rect 16046 -20297 16085 -20280
rect 15577 -20314 15802 -20297
rect 14842 -20352 15802 -20314
rect 15860 -20314 16085 -20297
rect 16119 -20314 16153 -20280
rect 16187 -20314 16221 -20280
rect 16255 -20314 16289 -20280
rect 16323 -20314 16357 -20280
rect 16391 -20314 16425 -20280
rect 16459 -20314 16493 -20280
rect 16527 -20314 16561 -20280
rect 16595 -20297 16634 -20280
rect 17064 -20280 17652 -20264
rect 17064 -20297 17103 -20280
rect 16595 -20314 16820 -20297
rect 15860 -20352 16820 -20314
rect 16878 -20314 17103 -20297
rect 17137 -20314 17171 -20280
rect 17205 -20314 17239 -20280
rect 17273 -20314 17307 -20280
rect 17341 -20314 17375 -20280
rect 17409 -20314 17443 -20280
rect 17477 -20314 17511 -20280
rect 17545 -20314 17579 -20280
rect 17613 -20297 17652 -20280
rect 18082 -20280 18670 -20264
rect 18082 -20297 18121 -20280
rect 17613 -20314 17838 -20297
rect 16878 -20352 17838 -20314
rect 17896 -20314 18121 -20297
rect 18155 -20314 18189 -20280
rect 18223 -20314 18257 -20280
rect 18291 -20314 18325 -20280
rect 18359 -20314 18393 -20280
rect 18427 -20314 18461 -20280
rect 18495 -20314 18529 -20280
rect 18563 -20314 18597 -20280
rect 18631 -20297 18670 -20280
rect 19100 -20280 19688 -20264
rect 19100 -20297 19139 -20280
rect 18631 -20314 18856 -20297
rect 17896 -20352 18856 -20314
rect 18914 -20314 19139 -20297
rect 19173 -20314 19207 -20280
rect 19241 -20314 19275 -20280
rect 19309 -20314 19343 -20280
rect 19377 -20314 19411 -20280
rect 19445 -20314 19479 -20280
rect 19513 -20314 19547 -20280
rect 19581 -20314 19615 -20280
rect 19649 -20297 19688 -20280
rect 20118 -20280 20706 -20264
rect 20118 -20297 20157 -20280
rect 19649 -20314 19874 -20297
rect 18914 -20352 19874 -20314
rect 19932 -20314 20157 -20297
rect 20191 -20314 20225 -20280
rect 20259 -20314 20293 -20280
rect 20327 -20314 20361 -20280
rect 20395 -20314 20429 -20280
rect 20463 -20314 20497 -20280
rect 20531 -20314 20565 -20280
rect 20599 -20314 20633 -20280
rect 20667 -20297 20706 -20280
rect 21136 -20280 21724 -20264
rect 21136 -20297 21175 -20280
rect 20667 -20314 20892 -20297
rect 19932 -20352 20892 -20314
rect 20950 -20314 21175 -20297
rect 21209 -20314 21243 -20280
rect 21277 -20314 21311 -20280
rect 21345 -20314 21379 -20280
rect 21413 -20314 21447 -20280
rect 21481 -20314 21515 -20280
rect 21549 -20314 21583 -20280
rect 21617 -20314 21651 -20280
rect 21685 -20297 21724 -20280
rect 22154 -20280 22742 -20264
rect 22154 -20297 22193 -20280
rect 21685 -20314 21910 -20297
rect 20950 -20352 21910 -20314
rect 21968 -20314 22193 -20297
rect 22227 -20314 22261 -20280
rect 22295 -20314 22329 -20280
rect 22363 -20314 22397 -20280
rect 22431 -20314 22465 -20280
rect 22499 -20314 22533 -20280
rect 22567 -20314 22601 -20280
rect 22635 -20314 22669 -20280
rect 22703 -20297 22742 -20280
rect 22703 -20314 22928 -20297
rect 21968 -20352 22928 -20314
rect -2252 -20382 -2144 -20366
rect -2252 -20399 -2215 -20382
rect -2278 -20416 -2215 -20399
rect -2181 -20399 -2144 -20382
rect -2034 -20382 -1926 -20366
rect -2034 -20399 -1997 -20382
rect -2181 -20416 -2118 -20399
rect -2278 -20454 -2118 -20416
rect -2060 -20416 -1997 -20399
rect -1963 -20399 -1926 -20382
rect -1816 -20382 -1708 -20366
rect -1816 -20399 -1779 -20382
rect -1963 -20416 -1900 -20399
rect -2060 -20454 -1900 -20416
rect -1842 -20416 -1779 -20399
rect -1745 -20399 -1708 -20382
rect -1598 -20382 -1490 -20366
rect -1598 -20399 -1561 -20382
rect -1745 -20416 -1682 -20399
rect -1842 -20454 -1682 -20416
rect -1624 -20416 -1561 -20399
rect -1527 -20399 -1490 -20382
rect -1380 -20382 -1272 -20366
rect -1380 -20399 -1343 -20382
rect -1527 -20416 -1464 -20399
rect -1624 -20454 -1464 -20416
rect -1406 -20416 -1343 -20399
rect -1309 -20399 -1272 -20382
rect -1162 -20382 -1054 -20366
rect -1162 -20399 -1125 -20382
rect -1309 -20416 -1246 -20399
rect -1406 -20454 -1246 -20416
rect -1188 -20416 -1125 -20399
rect -1091 -20399 -1054 -20382
rect -944 -20382 -836 -20366
rect -944 -20399 -907 -20382
rect -1091 -20416 -1028 -20399
rect -1188 -20454 -1028 -20416
rect -970 -20416 -907 -20399
rect -873 -20399 -836 -20382
rect -726 -20382 -618 -20366
rect -726 -20399 -689 -20382
rect -873 -20416 -810 -20399
rect -970 -20454 -810 -20416
rect -752 -20416 -689 -20399
rect -655 -20399 -618 -20382
rect -508 -20382 -400 -20366
rect -508 -20399 -471 -20382
rect -655 -20416 -592 -20399
rect -752 -20454 -592 -20416
rect -534 -20416 -471 -20399
rect -437 -20399 -400 -20382
rect -290 -20382 -182 -20366
rect -290 -20399 -253 -20382
rect -437 -20416 -374 -20399
rect -534 -20454 -374 -20416
rect -316 -20416 -253 -20399
rect -219 -20399 -182 -20382
rect -219 -20416 -156 -20399
rect -316 -20454 -156 -20416
rect -2278 -20692 -2118 -20654
rect -2278 -20709 -2215 -20692
rect -2252 -20726 -2215 -20709
rect -2181 -20709 -2118 -20692
rect -2060 -20692 -1900 -20654
rect -2060 -20709 -1997 -20692
rect -2181 -20726 -2144 -20709
rect -2252 -20742 -2144 -20726
rect -2034 -20726 -1997 -20709
rect -1963 -20709 -1900 -20692
rect -1842 -20692 -1682 -20654
rect -1842 -20709 -1779 -20692
rect -1963 -20726 -1926 -20709
rect -2034 -20742 -1926 -20726
rect -1816 -20726 -1779 -20709
rect -1745 -20709 -1682 -20692
rect -1624 -20692 -1464 -20654
rect -1624 -20709 -1561 -20692
rect -1745 -20726 -1708 -20709
rect -1816 -20742 -1708 -20726
rect -1598 -20726 -1561 -20709
rect -1527 -20709 -1464 -20692
rect -1406 -20692 -1246 -20654
rect -1406 -20709 -1343 -20692
rect -1527 -20726 -1490 -20709
rect -1598 -20742 -1490 -20726
rect -1380 -20726 -1343 -20709
rect -1309 -20709 -1246 -20692
rect -1188 -20692 -1028 -20654
rect -1188 -20709 -1125 -20692
rect -1309 -20726 -1272 -20709
rect -1380 -20742 -1272 -20726
rect -1162 -20726 -1125 -20709
rect -1091 -20709 -1028 -20692
rect -970 -20692 -810 -20654
rect -970 -20709 -907 -20692
rect -1091 -20726 -1054 -20709
rect -1162 -20742 -1054 -20726
rect -944 -20726 -907 -20709
rect -873 -20709 -810 -20692
rect -752 -20692 -592 -20654
rect -752 -20709 -689 -20692
rect -873 -20726 -836 -20709
rect -944 -20742 -836 -20726
rect -726 -20726 -689 -20709
rect -655 -20709 -592 -20692
rect -534 -20692 -374 -20654
rect -534 -20709 -471 -20692
rect -655 -20726 -618 -20709
rect -726 -20742 -618 -20726
rect -508 -20726 -471 -20709
rect -437 -20709 -374 -20692
rect -316 -20692 -156 -20654
rect -316 -20709 -253 -20692
rect -437 -20726 -400 -20709
rect -508 -20742 -400 -20726
rect -290 -20726 -253 -20709
rect -219 -20709 -156 -20692
rect -219 -20726 -182 -20709
rect -290 -20742 -182 -20726
rect 2626 -20990 3586 -20952
rect 2626 -21007 2851 -20990
rect 2812 -21024 2851 -21007
rect 2885 -21024 2919 -20990
rect 2953 -21024 2987 -20990
rect 3021 -21024 3055 -20990
rect 3089 -21024 3123 -20990
rect 3157 -21024 3191 -20990
rect 3225 -21024 3259 -20990
rect 3293 -21024 3327 -20990
rect 3361 -21007 3586 -20990
rect 3644 -20990 4604 -20952
rect 3644 -21007 3869 -20990
rect 3361 -21024 3400 -21007
rect 2812 -21040 3400 -21024
rect 3830 -21024 3869 -21007
rect 3903 -21024 3937 -20990
rect 3971 -21024 4005 -20990
rect 4039 -21024 4073 -20990
rect 4107 -21024 4141 -20990
rect 4175 -21024 4209 -20990
rect 4243 -21024 4277 -20990
rect 4311 -21024 4345 -20990
rect 4379 -21007 4604 -20990
rect 4662 -20990 5622 -20952
rect 4662 -21007 4887 -20990
rect 4379 -21024 4418 -21007
rect 3830 -21040 4418 -21024
rect 4848 -21024 4887 -21007
rect 4921 -21024 4955 -20990
rect 4989 -21024 5023 -20990
rect 5057 -21024 5091 -20990
rect 5125 -21024 5159 -20990
rect 5193 -21024 5227 -20990
rect 5261 -21024 5295 -20990
rect 5329 -21024 5363 -20990
rect 5397 -21007 5622 -20990
rect 5680 -20990 6640 -20952
rect 5680 -21007 5905 -20990
rect 5397 -21024 5436 -21007
rect 4848 -21040 5436 -21024
rect 5866 -21024 5905 -21007
rect 5939 -21024 5973 -20990
rect 6007 -21024 6041 -20990
rect 6075 -21024 6109 -20990
rect 6143 -21024 6177 -20990
rect 6211 -21024 6245 -20990
rect 6279 -21024 6313 -20990
rect 6347 -21024 6381 -20990
rect 6415 -21007 6640 -20990
rect 6698 -20990 7658 -20952
rect 6698 -21007 6923 -20990
rect 6415 -21024 6454 -21007
rect 5866 -21040 6454 -21024
rect 6884 -21024 6923 -21007
rect 6957 -21024 6991 -20990
rect 7025 -21024 7059 -20990
rect 7093 -21024 7127 -20990
rect 7161 -21024 7195 -20990
rect 7229 -21024 7263 -20990
rect 7297 -21024 7331 -20990
rect 7365 -21024 7399 -20990
rect 7433 -21007 7658 -20990
rect 7716 -20990 8676 -20952
rect 7716 -21007 7941 -20990
rect 7433 -21024 7472 -21007
rect 6884 -21040 7472 -21024
rect 7902 -21024 7941 -21007
rect 7975 -21024 8009 -20990
rect 8043 -21024 8077 -20990
rect 8111 -21024 8145 -20990
rect 8179 -21024 8213 -20990
rect 8247 -21024 8281 -20990
rect 8315 -21024 8349 -20990
rect 8383 -21024 8417 -20990
rect 8451 -21007 8676 -20990
rect 8734 -20990 9694 -20952
rect 8734 -21007 8959 -20990
rect 8451 -21024 8490 -21007
rect 7902 -21040 8490 -21024
rect 8920 -21024 8959 -21007
rect 8993 -21024 9027 -20990
rect 9061 -21024 9095 -20990
rect 9129 -21024 9163 -20990
rect 9197 -21024 9231 -20990
rect 9265 -21024 9299 -20990
rect 9333 -21024 9367 -20990
rect 9401 -21024 9435 -20990
rect 9469 -21007 9694 -20990
rect 9752 -20990 10712 -20952
rect 9752 -21007 9977 -20990
rect 9469 -21024 9508 -21007
rect 8920 -21040 9508 -21024
rect 9938 -21024 9977 -21007
rect 10011 -21024 10045 -20990
rect 10079 -21024 10113 -20990
rect 10147 -21024 10181 -20990
rect 10215 -21024 10249 -20990
rect 10283 -21024 10317 -20990
rect 10351 -21024 10385 -20990
rect 10419 -21024 10453 -20990
rect 10487 -21007 10712 -20990
rect 10770 -20990 11730 -20952
rect 10770 -21007 10995 -20990
rect 10487 -21024 10526 -21007
rect 9938 -21040 10526 -21024
rect 10956 -21024 10995 -21007
rect 11029 -21024 11063 -20990
rect 11097 -21024 11131 -20990
rect 11165 -21024 11199 -20990
rect 11233 -21024 11267 -20990
rect 11301 -21024 11335 -20990
rect 11369 -21024 11403 -20990
rect 11437 -21024 11471 -20990
rect 11505 -21007 11730 -20990
rect 11788 -20990 12748 -20952
rect 11788 -21007 12013 -20990
rect 11505 -21024 11544 -21007
rect 10956 -21040 11544 -21024
rect 11974 -21024 12013 -21007
rect 12047 -21024 12081 -20990
rect 12115 -21024 12149 -20990
rect 12183 -21024 12217 -20990
rect 12251 -21024 12285 -20990
rect 12319 -21024 12353 -20990
rect 12387 -21024 12421 -20990
rect 12455 -21024 12489 -20990
rect 12523 -21007 12748 -20990
rect 12806 -20990 13766 -20952
rect 12806 -21007 13031 -20990
rect 12523 -21024 12562 -21007
rect 11974 -21040 12562 -21024
rect 12992 -21024 13031 -21007
rect 13065 -21024 13099 -20990
rect 13133 -21024 13167 -20990
rect 13201 -21024 13235 -20990
rect 13269 -21024 13303 -20990
rect 13337 -21024 13371 -20990
rect 13405 -21024 13439 -20990
rect 13473 -21024 13507 -20990
rect 13541 -21007 13766 -20990
rect 13824 -20990 14784 -20952
rect 13824 -21007 14049 -20990
rect 13541 -21024 13580 -21007
rect 12992 -21040 13580 -21024
rect 14010 -21024 14049 -21007
rect 14083 -21024 14117 -20990
rect 14151 -21024 14185 -20990
rect 14219 -21024 14253 -20990
rect 14287 -21024 14321 -20990
rect 14355 -21024 14389 -20990
rect 14423 -21024 14457 -20990
rect 14491 -21024 14525 -20990
rect 14559 -21007 14784 -20990
rect 14842 -20990 15802 -20952
rect 14842 -21007 15067 -20990
rect 14559 -21024 14598 -21007
rect 14010 -21040 14598 -21024
rect 15028 -21024 15067 -21007
rect 15101 -21024 15135 -20990
rect 15169 -21024 15203 -20990
rect 15237 -21024 15271 -20990
rect 15305 -21024 15339 -20990
rect 15373 -21024 15407 -20990
rect 15441 -21024 15475 -20990
rect 15509 -21024 15543 -20990
rect 15577 -21007 15802 -20990
rect 15860 -20990 16820 -20952
rect 15860 -21007 16085 -20990
rect 15577 -21024 15616 -21007
rect 15028 -21040 15616 -21024
rect 16046 -21024 16085 -21007
rect 16119 -21024 16153 -20990
rect 16187 -21024 16221 -20990
rect 16255 -21024 16289 -20990
rect 16323 -21024 16357 -20990
rect 16391 -21024 16425 -20990
rect 16459 -21024 16493 -20990
rect 16527 -21024 16561 -20990
rect 16595 -21007 16820 -20990
rect 16878 -20990 17838 -20952
rect 16878 -21007 17103 -20990
rect 16595 -21024 16634 -21007
rect 16046 -21040 16634 -21024
rect 17064 -21024 17103 -21007
rect 17137 -21024 17171 -20990
rect 17205 -21024 17239 -20990
rect 17273 -21024 17307 -20990
rect 17341 -21024 17375 -20990
rect 17409 -21024 17443 -20990
rect 17477 -21024 17511 -20990
rect 17545 -21024 17579 -20990
rect 17613 -21007 17838 -20990
rect 17896 -20990 18856 -20952
rect 17896 -21007 18121 -20990
rect 17613 -21024 17652 -21007
rect 17064 -21040 17652 -21024
rect 18082 -21024 18121 -21007
rect 18155 -21024 18189 -20990
rect 18223 -21024 18257 -20990
rect 18291 -21024 18325 -20990
rect 18359 -21024 18393 -20990
rect 18427 -21024 18461 -20990
rect 18495 -21024 18529 -20990
rect 18563 -21024 18597 -20990
rect 18631 -21007 18856 -20990
rect 18914 -20990 19874 -20952
rect 18914 -21007 19139 -20990
rect 18631 -21024 18670 -21007
rect 18082 -21040 18670 -21024
rect 19100 -21024 19139 -21007
rect 19173 -21024 19207 -20990
rect 19241 -21024 19275 -20990
rect 19309 -21024 19343 -20990
rect 19377 -21024 19411 -20990
rect 19445 -21024 19479 -20990
rect 19513 -21024 19547 -20990
rect 19581 -21024 19615 -20990
rect 19649 -21007 19874 -20990
rect 19932 -20990 20892 -20952
rect 19932 -21007 20157 -20990
rect 19649 -21024 19688 -21007
rect 19100 -21040 19688 -21024
rect 20118 -21024 20157 -21007
rect 20191 -21024 20225 -20990
rect 20259 -21024 20293 -20990
rect 20327 -21024 20361 -20990
rect 20395 -21024 20429 -20990
rect 20463 -21024 20497 -20990
rect 20531 -21024 20565 -20990
rect 20599 -21024 20633 -20990
rect 20667 -21007 20892 -20990
rect 20950 -20990 21910 -20952
rect 20950 -21007 21175 -20990
rect 20667 -21024 20706 -21007
rect 20118 -21040 20706 -21024
rect 21136 -21024 21175 -21007
rect 21209 -21024 21243 -20990
rect 21277 -21024 21311 -20990
rect 21345 -21024 21379 -20990
rect 21413 -21024 21447 -20990
rect 21481 -21024 21515 -20990
rect 21549 -21024 21583 -20990
rect 21617 -21024 21651 -20990
rect 21685 -21007 21910 -20990
rect 21968 -20990 22928 -20952
rect 21968 -21007 22193 -20990
rect 21685 -21024 21724 -21007
rect 21136 -21040 21724 -21024
rect 22154 -21024 22193 -21007
rect 22227 -21024 22261 -20990
rect 22295 -21024 22329 -20990
rect 22363 -21024 22397 -20990
rect 22431 -21024 22465 -20990
rect 22499 -21024 22533 -20990
rect 22567 -21024 22601 -20990
rect 22635 -21024 22669 -20990
rect 22703 -21007 22928 -20990
rect 22703 -21024 22742 -21007
rect 22154 -21040 22742 -21024
rect 2812 -21512 3400 -21496
rect 2812 -21529 2851 -21512
rect 2626 -21546 2851 -21529
rect 2885 -21546 2919 -21512
rect 2953 -21546 2987 -21512
rect 3021 -21546 3055 -21512
rect 3089 -21546 3123 -21512
rect 3157 -21546 3191 -21512
rect 3225 -21546 3259 -21512
rect 3293 -21546 3327 -21512
rect 3361 -21529 3400 -21512
rect 3830 -21512 4418 -21496
rect 3830 -21529 3869 -21512
rect 3361 -21546 3586 -21529
rect 2626 -21584 3586 -21546
rect 3644 -21546 3869 -21529
rect 3903 -21546 3937 -21512
rect 3971 -21546 4005 -21512
rect 4039 -21546 4073 -21512
rect 4107 -21546 4141 -21512
rect 4175 -21546 4209 -21512
rect 4243 -21546 4277 -21512
rect 4311 -21546 4345 -21512
rect 4379 -21529 4418 -21512
rect 4848 -21512 5436 -21496
rect 4848 -21529 4887 -21512
rect 4379 -21546 4604 -21529
rect 3644 -21584 4604 -21546
rect 4662 -21546 4887 -21529
rect 4921 -21546 4955 -21512
rect 4989 -21546 5023 -21512
rect 5057 -21546 5091 -21512
rect 5125 -21546 5159 -21512
rect 5193 -21546 5227 -21512
rect 5261 -21546 5295 -21512
rect 5329 -21546 5363 -21512
rect 5397 -21529 5436 -21512
rect 5866 -21512 6454 -21496
rect 5866 -21529 5905 -21512
rect 5397 -21546 5622 -21529
rect 4662 -21584 5622 -21546
rect 5680 -21546 5905 -21529
rect 5939 -21546 5973 -21512
rect 6007 -21546 6041 -21512
rect 6075 -21546 6109 -21512
rect 6143 -21546 6177 -21512
rect 6211 -21546 6245 -21512
rect 6279 -21546 6313 -21512
rect 6347 -21546 6381 -21512
rect 6415 -21529 6454 -21512
rect 6884 -21512 7472 -21496
rect 6884 -21529 6923 -21512
rect 6415 -21546 6640 -21529
rect 5680 -21584 6640 -21546
rect 6698 -21546 6923 -21529
rect 6957 -21546 6991 -21512
rect 7025 -21546 7059 -21512
rect 7093 -21546 7127 -21512
rect 7161 -21546 7195 -21512
rect 7229 -21546 7263 -21512
rect 7297 -21546 7331 -21512
rect 7365 -21546 7399 -21512
rect 7433 -21529 7472 -21512
rect 7902 -21512 8490 -21496
rect 7902 -21529 7941 -21512
rect 7433 -21546 7658 -21529
rect 6698 -21584 7658 -21546
rect 7716 -21546 7941 -21529
rect 7975 -21546 8009 -21512
rect 8043 -21546 8077 -21512
rect 8111 -21546 8145 -21512
rect 8179 -21546 8213 -21512
rect 8247 -21546 8281 -21512
rect 8315 -21546 8349 -21512
rect 8383 -21546 8417 -21512
rect 8451 -21529 8490 -21512
rect 8920 -21512 9508 -21496
rect 8920 -21529 8959 -21512
rect 8451 -21546 8676 -21529
rect 7716 -21584 8676 -21546
rect 8734 -21546 8959 -21529
rect 8993 -21546 9027 -21512
rect 9061 -21546 9095 -21512
rect 9129 -21546 9163 -21512
rect 9197 -21546 9231 -21512
rect 9265 -21546 9299 -21512
rect 9333 -21546 9367 -21512
rect 9401 -21546 9435 -21512
rect 9469 -21529 9508 -21512
rect 9938 -21512 10526 -21496
rect 9938 -21529 9977 -21512
rect 9469 -21546 9694 -21529
rect 8734 -21584 9694 -21546
rect 9752 -21546 9977 -21529
rect 10011 -21546 10045 -21512
rect 10079 -21546 10113 -21512
rect 10147 -21546 10181 -21512
rect 10215 -21546 10249 -21512
rect 10283 -21546 10317 -21512
rect 10351 -21546 10385 -21512
rect 10419 -21546 10453 -21512
rect 10487 -21529 10526 -21512
rect 10956 -21512 11544 -21496
rect 10956 -21529 10995 -21512
rect 10487 -21546 10712 -21529
rect 9752 -21584 10712 -21546
rect 10770 -21546 10995 -21529
rect 11029 -21546 11063 -21512
rect 11097 -21546 11131 -21512
rect 11165 -21546 11199 -21512
rect 11233 -21546 11267 -21512
rect 11301 -21546 11335 -21512
rect 11369 -21546 11403 -21512
rect 11437 -21546 11471 -21512
rect 11505 -21529 11544 -21512
rect 11974 -21512 12562 -21496
rect 11974 -21529 12013 -21512
rect 11505 -21546 11730 -21529
rect 10770 -21584 11730 -21546
rect 11788 -21546 12013 -21529
rect 12047 -21546 12081 -21512
rect 12115 -21546 12149 -21512
rect 12183 -21546 12217 -21512
rect 12251 -21546 12285 -21512
rect 12319 -21546 12353 -21512
rect 12387 -21546 12421 -21512
rect 12455 -21546 12489 -21512
rect 12523 -21529 12562 -21512
rect 12992 -21512 13580 -21496
rect 12992 -21529 13031 -21512
rect 12523 -21546 12748 -21529
rect 11788 -21584 12748 -21546
rect 12806 -21546 13031 -21529
rect 13065 -21546 13099 -21512
rect 13133 -21546 13167 -21512
rect 13201 -21546 13235 -21512
rect 13269 -21546 13303 -21512
rect 13337 -21546 13371 -21512
rect 13405 -21546 13439 -21512
rect 13473 -21546 13507 -21512
rect 13541 -21529 13580 -21512
rect 14010 -21512 14598 -21496
rect 14010 -21529 14049 -21512
rect 13541 -21546 13766 -21529
rect 12806 -21584 13766 -21546
rect 13824 -21546 14049 -21529
rect 14083 -21546 14117 -21512
rect 14151 -21546 14185 -21512
rect 14219 -21546 14253 -21512
rect 14287 -21546 14321 -21512
rect 14355 -21546 14389 -21512
rect 14423 -21546 14457 -21512
rect 14491 -21546 14525 -21512
rect 14559 -21529 14598 -21512
rect 15028 -21512 15616 -21496
rect 15028 -21529 15067 -21512
rect 14559 -21546 14784 -21529
rect 13824 -21584 14784 -21546
rect 14842 -21546 15067 -21529
rect 15101 -21546 15135 -21512
rect 15169 -21546 15203 -21512
rect 15237 -21546 15271 -21512
rect 15305 -21546 15339 -21512
rect 15373 -21546 15407 -21512
rect 15441 -21546 15475 -21512
rect 15509 -21546 15543 -21512
rect 15577 -21529 15616 -21512
rect 16046 -21512 16634 -21496
rect 16046 -21529 16085 -21512
rect 15577 -21546 15802 -21529
rect 14842 -21584 15802 -21546
rect 15860 -21546 16085 -21529
rect 16119 -21546 16153 -21512
rect 16187 -21546 16221 -21512
rect 16255 -21546 16289 -21512
rect 16323 -21546 16357 -21512
rect 16391 -21546 16425 -21512
rect 16459 -21546 16493 -21512
rect 16527 -21546 16561 -21512
rect 16595 -21529 16634 -21512
rect 17064 -21512 17652 -21496
rect 17064 -21529 17103 -21512
rect 16595 -21546 16820 -21529
rect 15860 -21584 16820 -21546
rect 16878 -21546 17103 -21529
rect 17137 -21546 17171 -21512
rect 17205 -21546 17239 -21512
rect 17273 -21546 17307 -21512
rect 17341 -21546 17375 -21512
rect 17409 -21546 17443 -21512
rect 17477 -21546 17511 -21512
rect 17545 -21546 17579 -21512
rect 17613 -21529 17652 -21512
rect 18082 -21512 18670 -21496
rect 18082 -21529 18121 -21512
rect 17613 -21546 17838 -21529
rect 16878 -21584 17838 -21546
rect 17896 -21546 18121 -21529
rect 18155 -21546 18189 -21512
rect 18223 -21546 18257 -21512
rect 18291 -21546 18325 -21512
rect 18359 -21546 18393 -21512
rect 18427 -21546 18461 -21512
rect 18495 -21546 18529 -21512
rect 18563 -21546 18597 -21512
rect 18631 -21529 18670 -21512
rect 19100 -21512 19688 -21496
rect 19100 -21529 19139 -21512
rect 18631 -21546 18856 -21529
rect 17896 -21584 18856 -21546
rect 18914 -21546 19139 -21529
rect 19173 -21546 19207 -21512
rect 19241 -21546 19275 -21512
rect 19309 -21546 19343 -21512
rect 19377 -21546 19411 -21512
rect 19445 -21546 19479 -21512
rect 19513 -21546 19547 -21512
rect 19581 -21546 19615 -21512
rect 19649 -21529 19688 -21512
rect 20118 -21512 20706 -21496
rect 20118 -21529 20157 -21512
rect 19649 -21546 19874 -21529
rect 18914 -21584 19874 -21546
rect 19932 -21546 20157 -21529
rect 20191 -21546 20225 -21512
rect 20259 -21546 20293 -21512
rect 20327 -21546 20361 -21512
rect 20395 -21546 20429 -21512
rect 20463 -21546 20497 -21512
rect 20531 -21546 20565 -21512
rect 20599 -21546 20633 -21512
rect 20667 -21529 20706 -21512
rect 21136 -21512 21724 -21496
rect 21136 -21529 21175 -21512
rect 20667 -21546 20892 -21529
rect 19932 -21584 20892 -21546
rect 20950 -21546 21175 -21529
rect 21209 -21546 21243 -21512
rect 21277 -21546 21311 -21512
rect 21345 -21546 21379 -21512
rect 21413 -21546 21447 -21512
rect 21481 -21546 21515 -21512
rect 21549 -21546 21583 -21512
rect 21617 -21546 21651 -21512
rect 21685 -21529 21724 -21512
rect 22154 -21512 22742 -21496
rect 22154 -21529 22193 -21512
rect 21685 -21546 21910 -21529
rect 20950 -21584 21910 -21546
rect 21968 -21546 22193 -21529
rect 22227 -21546 22261 -21512
rect 22295 -21546 22329 -21512
rect 22363 -21546 22397 -21512
rect 22431 -21546 22465 -21512
rect 22499 -21546 22533 -21512
rect 22567 -21546 22601 -21512
rect 22635 -21546 22669 -21512
rect 22703 -21529 22742 -21512
rect 22703 -21546 22928 -21529
rect 21968 -21584 22928 -21546
rect -9173 -21709 -8585 -21693
rect -9173 -21726 -9134 -21709
rect -9359 -21743 -9134 -21726
rect -9100 -21743 -9066 -21709
rect -9032 -21743 -8998 -21709
rect -8964 -21743 -8930 -21709
rect -8896 -21743 -8862 -21709
rect -8828 -21743 -8794 -21709
rect -8760 -21743 -8726 -21709
rect -8692 -21743 -8658 -21709
rect -8624 -21726 -8585 -21709
rect -8155 -21709 -7567 -21693
rect -8155 -21726 -8116 -21709
rect -8624 -21743 -8399 -21726
rect -9359 -21781 -8399 -21743
rect -8341 -21743 -8116 -21726
rect -8082 -21743 -8048 -21709
rect -8014 -21743 -7980 -21709
rect -7946 -21743 -7912 -21709
rect -7878 -21743 -7844 -21709
rect -7810 -21743 -7776 -21709
rect -7742 -21743 -7708 -21709
rect -7674 -21743 -7640 -21709
rect -7606 -21726 -7567 -21709
rect -7137 -21709 -6549 -21693
rect -7137 -21726 -7098 -21709
rect -7606 -21743 -7381 -21726
rect -8341 -21781 -7381 -21743
rect -7323 -21743 -7098 -21726
rect -7064 -21743 -7030 -21709
rect -6996 -21743 -6962 -21709
rect -6928 -21743 -6894 -21709
rect -6860 -21743 -6826 -21709
rect -6792 -21743 -6758 -21709
rect -6724 -21743 -6690 -21709
rect -6656 -21743 -6622 -21709
rect -6588 -21726 -6549 -21709
rect -6119 -21709 -5531 -21693
rect -6119 -21726 -6080 -21709
rect -6588 -21743 -6363 -21726
rect -7323 -21781 -6363 -21743
rect -6305 -21743 -6080 -21726
rect -6046 -21743 -6012 -21709
rect -5978 -21743 -5944 -21709
rect -5910 -21743 -5876 -21709
rect -5842 -21743 -5808 -21709
rect -5774 -21743 -5740 -21709
rect -5706 -21743 -5672 -21709
rect -5638 -21743 -5604 -21709
rect -5570 -21726 -5531 -21709
rect -5101 -21709 -4513 -21693
rect -5101 -21726 -5062 -21709
rect -5570 -21743 -5345 -21726
rect -6305 -21781 -5345 -21743
rect -5287 -21743 -5062 -21726
rect -5028 -21743 -4994 -21709
rect -4960 -21743 -4926 -21709
rect -4892 -21743 -4858 -21709
rect -4824 -21743 -4790 -21709
rect -4756 -21743 -4722 -21709
rect -4688 -21743 -4654 -21709
rect -4620 -21743 -4586 -21709
rect -4552 -21726 -4513 -21709
rect -4083 -21709 -3495 -21693
rect -4083 -21726 -4044 -21709
rect -4552 -21743 -4327 -21726
rect -5287 -21781 -4327 -21743
rect -4269 -21743 -4044 -21726
rect -4010 -21743 -3976 -21709
rect -3942 -21743 -3908 -21709
rect -3874 -21743 -3840 -21709
rect -3806 -21743 -3772 -21709
rect -3738 -21743 -3704 -21709
rect -3670 -21743 -3636 -21709
rect -3602 -21743 -3568 -21709
rect -3534 -21726 -3495 -21709
rect -2322 -21708 -2166 -21692
rect -2322 -21725 -2295 -21708
rect -3534 -21743 -3309 -21726
rect -4269 -21781 -3309 -21743
rect -2364 -21742 -2295 -21725
rect -2261 -21742 -2227 -21708
rect -2193 -21725 -2166 -21708
rect -2024 -21708 -1868 -21692
rect -2024 -21725 -1997 -21708
rect -2193 -21742 -2124 -21725
rect -2364 -21780 -2124 -21742
rect -2066 -21742 -1997 -21725
rect -1963 -21742 -1929 -21708
rect -1895 -21725 -1868 -21708
rect -1726 -21708 -1570 -21692
rect -1726 -21725 -1699 -21708
rect -1895 -21742 -1826 -21725
rect -2066 -21780 -1826 -21742
rect -1768 -21742 -1699 -21725
rect -1665 -21742 -1631 -21708
rect -1597 -21725 -1570 -21708
rect -1428 -21708 -1272 -21692
rect -1428 -21725 -1401 -21708
rect -1597 -21742 -1528 -21725
rect -1768 -21780 -1528 -21742
rect -1470 -21742 -1401 -21725
rect -1367 -21742 -1333 -21708
rect -1299 -21725 -1272 -21708
rect -1130 -21708 -974 -21692
rect -1130 -21725 -1103 -21708
rect -1299 -21742 -1230 -21725
rect -1470 -21780 -1230 -21742
rect -1172 -21742 -1103 -21725
rect -1069 -21742 -1035 -21708
rect -1001 -21725 -974 -21708
rect -832 -21708 -676 -21692
rect -832 -21725 -805 -21708
rect -1001 -21742 -932 -21725
rect -1172 -21780 -932 -21742
rect -874 -21742 -805 -21725
rect -771 -21742 -737 -21708
rect -703 -21725 -676 -21708
rect -534 -21708 -378 -21692
rect -534 -21725 -507 -21708
rect -703 -21742 -634 -21725
rect -874 -21780 -634 -21742
rect -576 -21742 -507 -21725
rect -473 -21742 -439 -21708
rect -405 -21725 -378 -21708
rect -236 -21708 -80 -21692
rect -236 -21725 -209 -21708
rect -405 -21742 -336 -21725
rect -576 -21780 -336 -21742
rect -278 -21742 -209 -21725
rect -175 -21742 -141 -21708
rect -107 -21725 -80 -21708
rect 62 -21708 218 -21692
rect 62 -21725 89 -21708
rect -107 -21742 -38 -21725
rect -278 -21780 -38 -21742
rect 20 -21742 89 -21725
rect 123 -21742 157 -21708
rect 191 -21725 218 -21708
rect 360 -21708 516 -21692
rect 360 -21725 387 -21708
rect 191 -21742 260 -21725
rect 20 -21780 260 -21742
rect 318 -21742 387 -21725
rect 421 -21742 455 -21708
rect 489 -21725 516 -21708
rect 658 -21708 814 -21692
rect 658 -21725 685 -21708
rect 489 -21742 558 -21725
rect 318 -21780 558 -21742
rect 616 -21742 685 -21725
rect 719 -21742 753 -21708
rect 787 -21725 814 -21708
rect 787 -21742 856 -21725
rect 616 -21780 856 -21742
rect 2626 -22222 3586 -22184
rect 2626 -22239 2851 -22222
rect 2812 -22256 2851 -22239
rect 2885 -22256 2919 -22222
rect 2953 -22256 2987 -22222
rect 3021 -22256 3055 -22222
rect 3089 -22256 3123 -22222
rect 3157 -22256 3191 -22222
rect 3225 -22256 3259 -22222
rect 3293 -22256 3327 -22222
rect 3361 -22239 3586 -22222
rect 3644 -22222 4604 -22184
rect 3644 -22239 3869 -22222
rect 3361 -22256 3400 -22239
rect 2812 -22272 3400 -22256
rect 3830 -22256 3869 -22239
rect 3903 -22256 3937 -22222
rect 3971 -22256 4005 -22222
rect 4039 -22256 4073 -22222
rect 4107 -22256 4141 -22222
rect 4175 -22256 4209 -22222
rect 4243 -22256 4277 -22222
rect 4311 -22256 4345 -22222
rect 4379 -22239 4604 -22222
rect 4662 -22222 5622 -22184
rect 4662 -22239 4887 -22222
rect 4379 -22256 4418 -22239
rect 3830 -22272 4418 -22256
rect 4848 -22256 4887 -22239
rect 4921 -22256 4955 -22222
rect 4989 -22256 5023 -22222
rect 5057 -22256 5091 -22222
rect 5125 -22256 5159 -22222
rect 5193 -22256 5227 -22222
rect 5261 -22256 5295 -22222
rect 5329 -22256 5363 -22222
rect 5397 -22239 5622 -22222
rect 5680 -22222 6640 -22184
rect 5680 -22239 5905 -22222
rect 5397 -22256 5436 -22239
rect 4848 -22272 5436 -22256
rect 5866 -22256 5905 -22239
rect 5939 -22256 5973 -22222
rect 6007 -22256 6041 -22222
rect 6075 -22256 6109 -22222
rect 6143 -22256 6177 -22222
rect 6211 -22256 6245 -22222
rect 6279 -22256 6313 -22222
rect 6347 -22256 6381 -22222
rect 6415 -22239 6640 -22222
rect 6698 -22222 7658 -22184
rect 6698 -22239 6923 -22222
rect 6415 -22256 6454 -22239
rect 5866 -22272 6454 -22256
rect 6884 -22256 6923 -22239
rect 6957 -22256 6991 -22222
rect 7025 -22256 7059 -22222
rect 7093 -22256 7127 -22222
rect 7161 -22256 7195 -22222
rect 7229 -22256 7263 -22222
rect 7297 -22256 7331 -22222
rect 7365 -22256 7399 -22222
rect 7433 -22239 7658 -22222
rect 7716 -22222 8676 -22184
rect 7716 -22239 7941 -22222
rect 7433 -22256 7472 -22239
rect 6884 -22272 7472 -22256
rect 7902 -22256 7941 -22239
rect 7975 -22256 8009 -22222
rect 8043 -22256 8077 -22222
rect 8111 -22256 8145 -22222
rect 8179 -22256 8213 -22222
rect 8247 -22256 8281 -22222
rect 8315 -22256 8349 -22222
rect 8383 -22256 8417 -22222
rect 8451 -22239 8676 -22222
rect 8734 -22222 9694 -22184
rect 8734 -22239 8959 -22222
rect 8451 -22256 8490 -22239
rect 7902 -22272 8490 -22256
rect 8920 -22256 8959 -22239
rect 8993 -22256 9027 -22222
rect 9061 -22256 9095 -22222
rect 9129 -22256 9163 -22222
rect 9197 -22256 9231 -22222
rect 9265 -22256 9299 -22222
rect 9333 -22256 9367 -22222
rect 9401 -22256 9435 -22222
rect 9469 -22239 9694 -22222
rect 9752 -22222 10712 -22184
rect 9752 -22239 9977 -22222
rect 9469 -22256 9508 -22239
rect 8920 -22272 9508 -22256
rect 9938 -22256 9977 -22239
rect 10011 -22256 10045 -22222
rect 10079 -22256 10113 -22222
rect 10147 -22256 10181 -22222
rect 10215 -22256 10249 -22222
rect 10283 -22256 10317 -22222
rect 10351 -22256 10385 -22222
rect 10419 -22256 10453 -22222
rect 10487 -22239 10712 -22222
rect 10770 -22222 11730 -22184
rect 10770 -22239 10995 -22222
rect 10487 -22256 10526 -22239
rect 9938 -22272 10526 -22256
rect 10956 -22256 10995 -22239
rect 11029 -22256 11063 -22222
rect 11097 -22256 11131 -22222
rect 11165 -22256 11199 -22222
rect 11233 -22256 11267 -22222
rect 11301 -22256 11335 -22222
rect 11369 -22256 11403 -22222
rect 11437 -22256 11471 -22222
rect 11505 -22239 11730 -22222
rect 11788 -22222 12748 -22184
rect 11788 -22239 12013 -22222
rect 11505 -22256 11544 -22239
rect 10956 -22272 11544 -22256
rect 11974 -22256 12013 -22239
rect 12047 -22256 12081 -22222
rect 12115 -22256 12149 -22222
rect 12183 -22256 12217 -22222
rect 12251 -22256 12285 -22222
rect 12319 -22256 12353 -22222
rect 12387 -22256 12421 -22222
rect 12455 -22256 12489 -22222
rect 12523 -22239 12748 -22222
rect 12806 -22222 13766 -22184
rect 12806 -22239 13031 -22222
rect 12523 -22256 12562 -22239
rect 11974 -22272 12562 -22256
rect 12992 -22256 13031 -22239
rect 13065 -22256 13099 -22222
rect 13133 -22256 13167 -22222
rect 13201 -22256 13235 -22222
rect 13269 -22256 13303 -22222
rect 13337 -22256 13371 -22222
rect 13405 -22256 13439 -22222
rect 13473 -22256 13507 -22222
rect 13541 -22239 13766 -22222
rect 13824 -22222 14784 -22184
rect 13824 -22239 14049 -22222
rect 13541 -22256 13580 -22239
rect 12992 -22272 13580 -22256
rect 14010 -22256 14049 -22239
rect 14083 -22256 14117 -22222
rect 14151 -22256 14185 -22222
rect 14219 -22256 14253 -22222
rect 14287 -22256 14321 -22222
rect 14355 -22256 14389 -22222
rect 14423 -22256 14457 -22222
rect 14491 -22256 14525 -22222
rect 14559 -22239 14784 -22222
rect 14842 -22222 15802 -22184
rect 14842 -22239 15067 -22222
rect 14559 -22256 14598 -22239
rect 14010 -22272 14598 -22256
rect 15028 -22256 15067 -22239
rect 15101 -22256 15135 -22222
rect 15169 -22256 15203 -22222
rect 15237 -22256 15271 -22222
rect 15305 -22256 15339 -22222
rect 15373 -22256 15407 -22222
rect 15441 -22256 15475 -22222
rect 15509 -22256 15543 -22222
rect 15577 -22239 15802 -22222
rect 15860 -22222 16820 -22184
rect 15860 -22239 16085 -22222
rect 15577 -22256 15616 -22239
rect 15028 -22272 15616 -22256
rect 16046 -22256 16085 -22239
rect 16119 -22256 16153 -22222
rect 16187 -22256 16221 -22222
rect 16255 -22256 16289 -22222
rect 16323 -22256 16357 -22222
rect 16391 -22256 16425 -22222
rect 16459 -22256 16493 -22222
rect 16527 -22256 16561 -22222
rect 16595 -22239 16820 -22222
rect 16878 -22222 17838 -22184
rect 16878 -22239 17103 -22222
rect 16595 -22256 16634 -22239
rect 16046 -22272 16634 -22256
rect 17064 -22256 17103 -22239
rect 17137 -22256 17171 -22222
rect 17205 -22256 17239 -22222
rect 17273 -22256 17307 -22222
rect 17341 -22256 17375 -22222
rect 17409 -22256 17443 -22222
rect 17477 -22256 17511 -22222
rect 17545 -22256 17579 -22222
rect 17613 -22239 17838 -22222
rect 17896 -22222 18856 -22184
rect 17896 -22239 18121 -22222
rect 17613 -22256 17652 -22239
rect 17064 -22272 17652 -22256
rect 18082 -22256 18121 -22239
rect 18155 -22256 18189 -22222
rect 18223 -22256 18257 -22222
rect 18291 -22256 18325 -22222
rect 18359 -22256 18393 -22222
rect 18427 -22256 18461 -22222
rect 18495 -22256 18529 -22222
rect 18563 -22256 18597 -22222
rect 18631 -22239 18856 -22222
rect 18914 -22222 19874 -22184
rect 18914 -22239 19139 -22222
rect 18631 -22256 18670 -22239
rect 18082 -22272 18670 -22256
rect 19100 -22256 19139 -22239
rect 19173 -22256 19207 -22222
rect 19241 -22256 19275 -22222
rect 19309 -22256 19343 -22222
rect 19377 -22256 19411 -22222
rect 19445 -22256 19479 -22222
rect 19513 -22256 19547 -22222
rect 19581 -22256 19615 -22222
rect 19649 -22239 19874 -22222
rect 19932 -22222 20892 -22184
rect 19932 -22239 20157 -22222
rect 19649 -22256 19688 -22239
rect 19100 -22272 19688 -22256
rect 20118 -22256 20157 -22239
rect 20191 -22256 20225 -22222
rect 20259 -22256 20293 -22222
rect 20327 -22256 20361 -22222
rect 20395 -22256 20429 -22222
rect 20463 -22256 20497 -22222
rect 20531 -22256 20565 -22222
rect 20599 -22256 20633 -22222
rect 20667 -22239 20892 -22222
rect 20950 -22222 21910 -22184
rect 20950 -22239 21175 -22222
rect 20667 -22256 20706 -22239
rect 20118 -22272 20706 -22256
rect 21136 -22256 21175 -22239
rect 21209 -22256 21243 -22222
rect 21277 -22256 21311 -22222
rect 21345 -22256 21379 -22222
rect 21413 -22256 21447 -22222
rect 21481 -22256 21515 -22222
rect 21549 -22256 21583 -22222
rect 21617 -22256 21651 -22222
rect 21685 -22239 21910 -22222
rect 21968 -22222 22928 -22184
rect 21968 -22239 22193 -22222
rect 21685 -22256 21724 -22239
rect 21136 -22272 21724 -22256
rect 22154 -22256 22193 -22239
rect 22227 -22256 22261 -22222
rect 22295 -22256 22329 -22222
rect 22363 -22256 22397 -22222
rect 22431 -22256 22465 -22222
rect 22499 -22256 22533 -22222
rect 22567 -22256 22601 -22222
rect 22635 -22256 22669 -22222
rect 22703 -22239 22928 -22222
rect 22703 -22256 22742 -22239
rect 22154 -22272 22742 -22256
rect -9359 -22419 -8399 -22381
rect -9359 -22436 -9134 -22419
rect -9173 -22453 -9134 -22436
rect -9100 -22453 -9066 -22419
rect -9032 -22453 -8998 -22419
rect -8964 -22453 -8930 -22419
rect -8896 -22453 -8862 -22419
rect -8828 -22453 -8794 -22419
rect -8760 -22453 -8726 -22419
rect -8692 -22453 -8658 -22419
rect -8624 -22436 -8399 -22419
rect -8341 -22419 -7381 -22381
rect -8341 -22436 -8116 -22419
rect -8624 -22453 -8585 -22436
rect -9173 -22469 -8585 -22453
rect -8155 -22453 -8116 -22436
rect -8082 -22453 -8048 -22419
rect -8014 -22453 -7980 -22419
rect -7946 -22453 -7912 -22419
rect -7878 -22453 -7844 -22419
rect -7810 -22453 -7776 -22419
rect -7742 -22453 -7708 -22419
rect -7674 -22453 -7640 -22419
rect -7606 -22436 -7381 -22419
rect -7323 -22419 -6363 -22381
rect -7323 -22436 -7098 -22419
rect -7606 -22453 -7567 -22436
rect -8155 -22469 -7567 -22453
rect -7137 -22453 -7098 -22436
rect -7064 -22453 -7030 -22419
rect -6996 -22453 -6962 -22419
rect -6928 -22453 -6894 -22419
rect -6860 -22453 -6826 -22419
rect -6792 -22453 -6758 -22419
rect -6724 -22453 -6690 -22419
rect -6656 -22453 -6622 -22419
rect -6588 -22436 -6363 -22419
rect -6305 -22419 -5345 -22381
rect -6305 -22436 -6080 -22419
rect -6588 -22453 -6549 -22436
rect -7137 -22469 -6549 -22453
rect -6119 -22453 -6080 -22436
rect -6046 -22453 -6012 -22419
rect -5978 -22453 -5944 -22419
rect -5910 -22453 -5876 -22419
rect -5842 -22453 -5808 -22419
rect -5774 -22453 -5740 -22419
rect -5706 -22453 -5672 -22419
rect -5638 -22453 -5604 -22419
rect -5570 -22436 -5345 -22419
rect -5287 -22419 -4327 -22381
rect -5287 -22436 -5062 -22419
rect -5570 -22453 -5531 -22436
rect -6119 -22469 -5531 -22453
rect -5101 -22453 -5062 -22436
rect -5028 -22453 -4994 -22419
rect -4960 -22453 -4926 -22419
rect -4892 -22453 -4858 -22419
rect -4824 -22453 -4790 -22419
rect -4756 -22453 -4722 -22419
rect -4688 -22453 -4654 -22419
rect -4620 -22453 -4586 -22419
rect -4552 -22436 -4327 -22419
rect -4269 -22419 -3309 -22381
rect -4269 -22436 -4044 -22419
rect -4552 -22453 -4513 -22436
rect -5101 -22469 -4513 -22453
rect -4083 -22453 -4044 -22436
rect -4010 -22453 -3976 -22419
rect -3942 -22453 -3908 -22419
rect -3874 -22453 -3840 -22419
rect -3806 -22453 -3772 -22419
rect -3738 -22453 -3704 -22419
rect -3670 -22453 -3636 -22419
rect -3602 -22453 -3568 -22419
rect -3534 -22436 -3309 -22419
rect -2364 -22418 -2124 -22380
rect -2364 -22435 -2295 -22418
rect -3534 -22453 -3495 -22436
rect -4083 -22469 -3495 -22453
rect -2322 -22452 -2295 -22435
rect -2261 -22452 -2227 -22418
rect -2193 -22435 -2124 -22418
rect -2066 -22418 -1826 -22380
rect -2066 -22435 -1997 -22418
rect -2193 -22452 -2166 -22435
rect -2322 -22468 -2166 -22452
rect -2024 -22452 -1997 -22435
rect -1963 -22452 -1929 -22418
rect -1895 -22435 -1826 -22418
rect -1768 -22418 -1528 -22380
rect -1768 -22435 -1699 -22418
rect -1895 -22452 -1868 -22435
rect -2024 -22468 -1868 -22452
rect -1726 -22452 -1699 -22435
rect -1665 -22452 -1631 -22418
rect -1597 -22435 -1528 -22418
rect -1470 -22418 -1230 -22380
rect -1470 -22435 -1401 -22418
rect -1597 -22452 -1570 -22435
rect -1726 -22468 -1570 -22452
rect -1428 -22452 -1401 -22435
rect -1367 -22452 -1333 -22418
rect -1299 -22435 -1230 -22418
rect -1172 -22418 -932 -22380
rect -1172 -22435 -1103 -22418
rect -1299 -22452 -1272 -22435
rect -1428 -22468 -1272 -22452
rect -1130 -22452 -1103 -22435
rect -1069 -22452 -1035 -22418
rect -1001 -22435 -932 -22418
rect -874 -22418 -634 -22380
rect -874 -22435 -805 -22418
rect -1001 -22452 -974 -22435
rect -1130 -22468 -974 -22452
rect -832 -22452 -805 -22435
rect -771 -22452 -737 -22418
rect -703 -22435 -634 -22418
rect -576 -22418 -336 -22380
rect -576 -22435 -507 -22418
rect -703 -22452 -676 -22435
rect -832 -22468 -676 -22452
rect -534 -22452 -507 -22435
rect -473 -22452 -439 -22418
rect -405 -22435 -336 -22418
rect -278 -22418 -38 -22380
rect -278 -22435 -209 -22418
rect -405 -22452 -378 -22435
rect -534 -22468 -378 -22452
rect -236 -22452 -209 -22435
rect -175 -22452 -141 -22418
rect -107 -22435 -38 -22418
rect 20 -22418 260 -22380
rect 20 -22435 89 -22418
rect -107 -22452 -80 -22435
rect -236 -22468 -80 -22452
rect 62 -22452 89 -22435
rect 123 -22452 157 -22418
rect 191 -22435 260 -22418
rect 318 -22418 558 -22380
rect 318 -22435 387 -22418
rect 191 -22452 218 -22435
rect 62 -22468 218 -22452
rect 360 -22452 387 -22435
rect 421 -22452 455 -22418
rect 489 -22435 558 -22418
rect 616 -22418 856 -22380
rect 616 -22435 685 -22418
rect 489 -22452 516 -22435
rect 360 -22468 516 -22452
rect 658 -22452 685 -22435
rect 719 -22452 753 -22418
rect 787 -22435 856 -22418
rect 787 -22452 814 -22435
rect 658 -22468 814 -22452
rect 2812 -22746 3400 -22730
rect 2812 -22763 2851 -22746
rect 2626 -22780 2851 -22763
rect 2885 -22780 2919 -22746
rect 2953 -22780 2987 -22746
rect 3021 -22780 3055 -22746
rect 3089 -22780 3123 -22746
rect 3157 -22780 3191 -22746
rect 3225 -22780 3259 -22746
rect 3293 -22780 3327 -22746
rect 3361 -22763 3400 -22746
rect 3830 -22746 4418 -22730
rect 3830 -22763 3869 -22746
rect 3361 -22780 3586 -22763
rect -9174 -22822 -8586 -22806
rect -9174 -22839 -9135 -22822
rect -9360 -22856 -9135 -22839
rect -9101 -22856 -9067 -22822
rect -9033 -22856 -8999 -22822
rect -8965 -22856 -8931 -22822
rect -8897 -22856 -8863 -22822
rect -8829 -22856 -8795 -22822
rect -8761 -22856 -8727 -22822
rect -8693 -22856 -8659 -22822
rect -8625 -22839 -8586 -22822
rect -8156 -22822 -7568 -22806
rect -8156 -22839 -8117 -22822
rect -8625 -22856 -8400 -22839
rect -9360 -22894 -8400 -22856
rect -8342 -22856 -8117 -22839
rect -8083 -22856 -8049 -22822
rect -8015 -22856 -7981 -22822
rect -7947 -22856 -7913 -22822
rect -7879 -22856 -7845 -22822
rect -7811 -22856 -7777 -22822
rect -7743 -22856 -7709 -22822
rect -7675 -22856 -7641 -22822
rect -7607 -22839 -7568 -22822
rect -7138 -22822 -6550 -22806
rect -7138 -22839 -7099 -22822
rect -7607 -22856 -7382 -22839
rect -8342 -22894 -7382 -22856
rect -7324 -22856 -7099 -22839
rect -7065 -22856 -7031 -22822
rect -6997 -22856 -6963 -22822
rect -6929 -22856 -6895 -22822
rect -6861 -22856 -6827 -22822
rect -6793 -22856 -6759 -22822
rect -6725 -22856 -6691 -22822
rect -6657 -22856 -6623 -22822
rect -6589 -22839 -6550 -22822
rect -6120 -22822 -5532 -22806
rect -6120 -22839 -6081 -22822
rect -6589 -22856 -6364 -22839
rect -7324 -22894 -6364 -22856
rect -6306 -22856 -6081 -22839
rect -6047 -22856 -6013 -22822
rect -5979 -22856 -5945 -22822
rect -5911 -22856 -5877 -22822
rect -5843 -22856 -5809 -22822
rect -5775 -22856 -5741 -22822
rect -5707 -22856 -5673 -22822
rect -5639 -22856 -5605 -22822
rect -5571 -22839 -5532 -22822
rect -5102 -22822 -4514 -22806
rect -5102 -22839 -5063 -22822
rect -5571 -22856 -5346 -22839
rect -6306 -22894 -5346 -22856
rect -5288 -22856 -5063 -22839
rect -5029 -22856 -4995 -22822
rect -4961 -22856 -4927 -22822
rect -4893 -22856 -4859 -22822
rect -4825 -22856 -4791 -22822
rect -4757 -22856 -4723 -22822
rect -4689 -22856 -4655 -22822
rect -4621 -22856 -4587 -22822
rect -4553 -22839 -4514 -22822
rect -4084 -22822 -3496 -22806
rect -4084 -22839 -4045 -22822
rect -4553 -22856 -4328 -22839
rect -5288 -22894 -4328 -22856
rect -4270 -22856 -4045 -22839
rect -4011 -22856 -3977 -22822
rect -3943 -22856 -3909 -22822
rect -3875 -22856 -3841 -22822
rect -3807 -22856 -3773 -22822
rect -3739 -22856 -3705 -22822
rect -3671 -22856 -3637 -22822
rect -3603 -22856 -3569 -22822
rect -3535 -22839 -3496 -22822
rect -2322 -22820 -2166 -22804
rect -2322 -22837 -2295 -22820
rect -3535 -22856 -3310 -22839
rect -4270 -22894 -3310 -22856
rect -2364 -22854 -2295 -22837
rect -2261 -22854 -2227 -22820
rect -2193 -22837 -2166 -22820
rect -2024 -22820 -1868 -22804
rect -2024 -22837 -1997 -22820
rect -2193 -22854 -2124 -22837
rect -2364 -22892 -2124 -22854
rect -2066 -22854 -1997 -22837
rect -1963 -22854 -1929 -22820
rect -1895 -22837 -1868 -22820
rect -1726 -22820 -1570 -22804
rect -1726 -22837 -1699 -22820
rect -1895 -22854 -1826 -22837
rect -2066 -22892 -1826 -22854
rect -1768 -22854 -1699 -22837
rect -1665 -22854 -1631 -22820
rect -1597 -22837 -1570 -22820
rect -1428 -22820 -1272 -22804
rect -1428 -22837 -1401 -22820
rect -1597 -22854 -1528 -22837
rect -1768 -22892 -1528 -22854
rect -1470 -22854 -1401 -22837
rect -1367 -22854 -1333 -22820
rect -1299 -22837 -1272 -22820
rect -1130 -22820 -974 -22804
rect -1130 -22837 -1103 -22820
rect -1299 -22854 -1230 -22837
rect -1470 -22892 -1230 -22854
rect -1172 -22854 -1103 -22837
rect -1069 -22854 -1035 -22820
rect -1001 -22837 -974 -22820
rect -832 -22820 -676 -22804
rect -832 -22837 -805 -22820
rect -1001 -22854 -932 -22837
rect -1172 -22892 -932 -22854
rect -874 -22854 -805 -22837
rect -771 -22854 -737 -22820
rect -703 -22837 -676 -22820
rect -534 -22820 -378 -22804
rect -534 -22837 -507 -22820
rect -703 -22854 -634 -22837
rect -874 -22892 -634 -22854
rect -576 -22854 -507 -22837
rect -473 -22854 -439 -22820
rect -405 -22837 -378 -22820
rect -236 -22820 -80 -22804
rect -236 -22837 -209 -22820
rect -405 -22854 -336 -22837
rect -576 -22892 -336 -22854
rect -278 -22854 -209 -22837
rect -175 -22854 -141 -22820
rect -107 -22837 -80 -22820
rect 62 -22820 218 -22804
rect 62 -22837 89 -22820
rect -107 -22854 -38 -22837
rect -278 -22892 -38 -22854
rect 20 -22854 89 -22837
rect 123 -22854 157 -22820
rect 191 -22837 218 -22820
rect 360 -22820 516 -22804
rect 360 -22837 387 -22820
rect 191 -22854 260 -22837
rect 20 -22892 260 -22854
rect 318 -22854 387 -22837
rect 421 -22854 455 -22820
rect 489 -22837 516 -22820
rect 658 -22820 814 -22804
rect 2626 -22818 3586 -22780
rect 3644 -22780 3869 -22763
rect 3903 -22780 3937 -22746
rect 3971 -22780 4005 -22746
rect 4039 -22780 4073 -22746
rect 4107 -22780 4141 -22746
rect 4175 -22780 4209 -22746
rect 4243 -22780 4277 -22746
rect 4311 -22780 4345 -22746
rect 4379 -22763 4418 -22746
rect 4848 -22746 5436 -22730
rect 4848 -22763 4887 -22746
rect 4379 -22780 4604 -22763
rect 3644 -22818 4604 -22780
rect 4662 -22780 4887 -22763
rect 4921 -22780 4955 -22746
rect 4989 -22780 5023 -22746
rect 5057 -22780 5091 -22746
rect 5125 -22780 5159 -22746
rect 5193 -22780 5227 -22746
rect 5261 -22780 5295 -22746
rect 5329 -22780 5363 -22746
rect 5397 -22763 5436 -22746
rect 5866 -22746 6454 -22730
rect 5866 -22763 5905 -22746
rect 5397 -22780 5622 -22763
rect 4662 -22818 5622 -22780
rect 5680 -22780 5905 -22763
rect 5939 -22780 5973 -22746
rect 6007 -22780 6041 -22746
rect 6075 -22780 6109 -22746
rect 6143 -22780 6177 -22746
rect 6211 -22780 6245 -22746
rect 6279 -22780 6313 -22746
rect 6347 -22780 6381 -22746
rect 6415 -22763 6454 -22746
rect 6884 -22746 7472 -22730
rect 6884 -22763 6923 -22746
rect 6415 -22780 6640 -22763
rect 5680 -22818 6640 -22780
rect 6698 -22780 6923 -22763
rect 6957 -22780 6991 -22746
rect 7025 -22780 7059 -22746
rect 7093 -22780 7127 -22746
rect 7161 -22780 7195 -22746
rect 7229 -22780 7263 -22746
rect 7297 -22780 7331 -22746
rect 7365 -22780 7399 -22746
rect 7433 -22763 7472 -22746
rect 7902 -22746 8490 -22730
rect 7902 -22763 7941 -22746
rect 7433 -22780 7658 -22763
rect 6698 -22818 7658 -22780
rect 7716 -22780 7941 -22763
rect 7975 -22780 8009 -22746
rect 8043 -22780 8077 -22746
rect 8111 -22780 8145 -22746
rect 8179 -22780 8213 -22746
rect 8247 -22780 8281 -22746
rect 8315 -22780 8349 -22746
rect 8383 -22780 8417 -22746
rect 8451 -22763 8490 -22746
rect 8920 -22746 9508 -22730
rect 8920 -22763 8959 -22746
rect 8451 -22780 8676 -22763
rect 7716 -22818 8676 -22780
rect 8734 -22780 8959 -22763
rect 8993 -22780 9027 -22746
rect 9061 -22780 9095 -22746
rect 9129 -22780 9163 -22746
rect 9197 -22780 9231 -22746
rect 9265 -22780 9299 -22746
rect 9333 -22780 9367 -22746
rect 9401 -22780 9435 -22746
rect 9469 -22763 9508 -22746
rect 9938 -22746 10526 -22730
rect 9938 -22763 9977 -22746
rect 9469 -22780 9694 -22763
rect 8734 -22818 9694 -22780
rect 9752 -22780 9977 -22763
rect 10011 -22780 10045 -22746
rect 10079 -22780 10113 -22746
rect 10147 -22780 10181 -22746
rect 10215 -22780 10249 -22746
rect 10283 -22780 10317 -22746
rect 10351 -22780 10385 -22746
rect 10419 -22780 10453 -22746
rect 10487 -22763 10526 -22746
rect 10956 -22746 11544 -22730
rect 10956 -22763 10995 -22746
rect 10487 -22780 10712 -22763
rect 9752 -22818 10712 -22780
rect 10770 -22780 10995 -22763
rect 11029 -22780 11063 -22746
rect 11097 -22780 11131 -22746
rect 11165 -22780 11199 -22746
rect 11233 -22780 11267 -22746
rect 11301 -22780 11335 -22746
rect 11369 -22780 11403 -22746
rect 11437 -22780 11471 -22746
rect 11505 -22763 11544 -22746
rect 11974 -22746 12562 -22730
rect 11974 -22763 12013 -22746
rect 11505 -22780 11730 -22763
rect 10770 -22818 11730 -22780
rect 11788 -22780 12013 -22763
rect 12047 -22780 12081 -22746
rect 12115 -22780 12149 -22746
rect 12183 -22780 12217 -22746
rect 12251 -22780 12285 -22746
rect 12319 -22780 12353 -22746
rect 12387 -22780 12421 -22746
rect 12455 -22780 12489 -22746
rect 12523 -22763 12562 -22746
rect 12992 -22746 13580 -22730
rect 12992 -22763 13031 -22746
rect 12523 -22780 12748 -22763
rect 11788 -22818 12748 -22780
rect 12806 -22780 13031 -22763
rect 13065 -22780 13099 -22746
rect 13133 -22780 13167 -22746
rect 13201 -22780 13235 -22746
rect 13269 -22780 13303 -22746
rect 13337 -22780 13371 -22746
rect 13405 -22780 13439 -22746
rect 13473 -22780 13507 -22746
rect 13541 -22763 13580 -22746
rect 14010 -22746 14598 -22730
rect 14010 -22763 14049 -22746
rect 13541 -22780 13766 -22763
rect 12806 -22818 13766 -22780
rect 13824 -22780 14049 -22763
rect 14083 -22780 14117 -22746
rect 14151 -22780 14185 -22746
rect 14219 -22780 14253 -22746
rect 14287 -22780 14321 -22746
rect 14355 -22780 14389 -22746
rect 14423 -22780 14457 -22746
rect 14491 -22780 14525 -22746
rect 14559 -22763 14598 -22746
rect 15028 -22746 15616 -22730
rect 15028 -22763 15067 -22746
rect 14559 -22780 14784 -22763
rect 13824 -22818 14784 -22780
rect 14842 -22780 15067 -22763
rect 15101 -22780 15135 -22746
rect 15169 -22780 15203 -22746
rect 15237 -22780 15271 -22746
rect 15305 -22780 15339 -22746
rect 15373 -22780 15407 -22746
rect 15441 -22780 15475 -22746
rect 15509 -22780 15543 -22746
rect 15577 -22763 15616 -22746
rect 16046 -22746 16634 -22730
rect 16046 -22763 16085 -22746
rect 15577 -22780 15802 -22763
rect 14842 -22818 15802 -22780
rect 15860 -22780 16085 -22763
rect 16119 -22780 16153 -22746
rect 16187 -22780 16221 -22746
rect 16255 -22780 16289 -22746
rect 16323 -22780 16357 -22746
rect 16391 -22780 16425 -22746
rect 16459 -22780 16493 -22746
rect 16527 -22780 16561 -22746
rect 16595 -22763 16634 -22746
rect 17064 -22746 17652 -22730
rect 17064 -22763 17103 -22746
rect 16595 -22780 16820 -22763
rect 15860 -22818 16820 -22780
rect 16878 -22780 17103 -22763
rect 17137 -22780 17171 -22746
rect 17205 -22780 17239 -22746
rect 17273 -22780 17307 -22746
rect 17341 -22780 17375 -22746
rect 17409 -22780 17443 -22746
rect 17477 -22780 17511 -22746
rect 17545 -22780 17579 -22746
rect 17613 -22763 17652 -22746
rect 18082 -22746 18670 -22730
rect 18082 -22763 18121 -22746
rect 17613 -22780 17838 -22763
rect 16878 -22818 17838 -22780
rect 17896 -22780 18121 -22763
rect 18155 -22780 18189 -22746
rect 18223 -22780 18257 -22746
rect 18291 -22780 18325 -22746
rect 18359 -22780 18393 -22746
rect 18427 -22780 18461 -22746
rect 18495 -22780 18529 -22746
rect 18563 -22780 18597 -22746
rect 18631 -22763 18670 -22746
rect 19100 -22746 19688 -22730
rect 19100 -22763 19139 -22746
rect 18631 -22780 18856 -22763
rect 17896 -22818 18856 -22780
rect 18914 -22780 19139 -22763
rect 19173 -22780 19207 -22746
rect 19241 -22780 19275 -22746
rect 19309 -22780 19343 -22746
rect 19377 -22780 19411 -22746
rect 19445 -22780 19479 -22746
rect 19513 -22780 19547 -22746
rect 19581 -22780 19615 -22746
rect 19649 -22763 19688 -22746
rect 20118 -22746 20706 -22730
rect 20118 -22763 20157 -22746
rect 19649 -22780 19874 -22763
rect 18914 -22818 19874 -22780
rect 19932 -22780 20157 -22763
rect 20191 -22780 20225 -22746
rect 20259 -22780 20293 -22746
rect 20327 -22780 20361 -22746
rect 20395 -22780 20429 -22746
rect 20463 -22780 20497 -22746
rect 20531 -22780 20565 -22746
rect 20599 -22780 20633 -22746
rect 20667 -22763 20706 -22746
rect 21136 -22746 21724 -22730
rect 21136 -22763 21175 -22746
rect 20667 -22780 20892 -22763
rect 19932 -22818 20892 -22780
rect 20950 -22780 21175 -22763
rect 21209 -22780 21243 -22746
rect 21277 -22780 21311 -22746
rect 21345 -22780 21379 -22746
rect 21413 -22780 21447 -22746
rect 21481 -22780 21515 -22746
rect 21549 -22780 21583 -22746
rect 21617 -22780 21651 -22746
rect 21685 -22763 21724 -22746
rect 22154 -22746 22742 -22730
rect 22154 -22763 22193 -22746
rect 21685 -22780 21910 -22763
rect 20950 -22818 21910 -22780
rect 21968 -22780 22193 -22763
rect 22227 -22780 22261 -22746
rect 22295 -22780 22329 -22746
rect 22363 -22780 22397 -22746
rect 22431 -22780 22465 -22746
rect 22499 -22780 22533 -22746
rect 22567 -22780 22601 -22746
rect 22635 -22780 22669 -22746
rect 22703 -22763 22742 -22746
rect 22703 -22780 22928 -22763
rect 21968 -22818 22928 -22780
rect 658 -22837 685 -22820
rect 489 -22854 558 -22837
rect 318 -22892 558 -22854
rect 616 -22854 685 -22837
rect 719 -22854 753 -22820
rect 787 -22837 814 -22820
rect 787 -22854 856 -22837
rect 616 -22892 856 -22854
rect 2626 -23456 3586 -23418
rect 2626 -23473 2851 -23456
rect 2812 -23490 2851 -23473
rect 2885 -23490 2919 -23456
rect 2953 -23490 2987 -23456
rect 3021 -23490 3055 -23456
rect 3089 -23490 3123 -23456
rect 3157 -23490 3191 -23456
rect 3225 -23490 3259 -23456
rect 3293 -23490 3327 -23456
rect 3361 -23473 3586 -23456
rect 3644 -23456 4604 -23418
rect 3644 -23473 3869 -23456
rect 3361 -23490 3400 -23473
rect -9360 -23532 -8400 -23494
rect -9360 -23549 -9135 -23532
rect -9174 -23566 -9135 -23549
rect -9101 -23566 -9067 -23532
rect -9033 -23566 -8999 -23532
rect -8965 -23566 -8931 -23532
rect -8897 -23566 -8863 -23532
rect -8829 -23566 -8795 -23532
rect -8761 -23566 -8727 -23532
rect -8693 -23566 -8659 -23532
rect -8625 -23549 -8400 -23532
rect -8342 -23532 -7382 -23494
rect -8342 -23549 -8117 -23532
rect -8625 -23566 -8586 -23549
rect -9174 -23582 -8586 -23566
rect -8156 -23566 -8117 -23549
rect -8083 -23566 -8049 -23532
rect -8015 -23566 -7981 -23532
rect -7947 -23566 -7913 -23532
rect -7879 -23566 -7845 -23532
rect -7811 -23566 -7777 -23532
rect -7743 -23566 -7709 -23532
rect -7675 -23566 -7641 -23532
rect -7607 -23549 -7382 -23532
rect -7324 -23532 -6364 -23494
rect -7324 -23549 -7099 -23532
rect -7607 -23566 -7568 -23549
rect -8156 -23582 -7568 -23566
rect -7138 -23566 -7099 -23549
rect -7065 -23566 -7031 -23532
rect -6997 -23566 -6963 -23532
rect -6929 -23566 -6895 -23532
rect -6861 -23566 -6827 -23532
rect -6793 -23566 -6759 -23532
rect -6725 -23566 -6691 -23532
rect -6657 -23566 -6623 -23532
rect -6589 -23549 -6364 -23532
rect -6306 -23532 -5346 -23494
rect -6306 -23549 -6081 -23532
rect -6589 -23566 -6550 -23549
rect -7138 -23582 -6550 -23566
rect -6120 -23566 -6081 -23549
rect -6047 -23566 -6013 -23532
rect -5979 -23566 -5945 -23532
rect -5911 -23566 -5877 -23532
rect -5843 -23566 -5809 -23532
rect -5775 -23566 -5741 -23532
rect -5707 -23566 -5673 -23532
rect -5639 -23566 -5605 -23532
rect -5571 -23549 -5346 -23532
rect -5288 -23532 -4328 -23494
rect -5288 -23549 -5063 -23532
rect -5571 -23566 -5532 -23549
rect -6120 -23582 -5532 -23566
rect -5102 -23566 -5063 -23549
rect -5029 -23566 -4995 -23532
rect -4961 -23566 -4927 -23532
rect -4893 -23566 -4859 -23532
rect -4825 -23566 -4791 -23532
rect -4757 -23566 -4723 -23532
rect -4689 -23566 -4655 -23532
rect -4621 -23566 -4587 -23532
rect -4553 -23549 -4328 -23532
rect -4270 -23532 -3310 -23494
rect -4270 -23549 -4045 -23532
rect -4553 -23566 -4514 -23549
rect -5102 -23582 -4514 -23566
rect -4084 -23566 -4045 -23549
rect -4011 -23566 -3977 -23532
rect -3943 -23566 -3909 -23532
rect -3875 -23566 -3841 -23532
rect -3807 -23566 -3773 -23532
rect -3739 -23566 -3705 -23532
rect -3671 -23566 -3637 -23532
rect -3603 -23566 -3569 -23532
rect -3535 -23549 -3310 -23532
rect -2364 -23530 -2124 -23492
rect -2364 -23547 -2295 -23530
rect -3535 -23566 -3496 -23549
rect -4084 -23582 -3496 -23566
rect -2322 -23564 -2295 -23547
rect -2261 -23564 -2227 -23530
rect -2193 -23547 -2124 -23530
rect -2066 -23530 -1826 -23492
rect -2066 -23547 -1997 -23530
rect -2193 -23564 -2166 -23547
rect -2322 -23580 -2166 -23564
rect -2024 -23564 -1997 -23547
rect -1963 -23564 -1929 -23530
rect -1895 -23547 -1826 -23530
rect -1768 -23530 -1528 -23492
rect -1768 -23547 -1699 -23530
rect -1895 -23564 -1868 -23547
rect -2024 -23580 -1868 -23564
rect -1726 -23564 -1699 -23547
rect -1665 -23564 -1631 -23530
rect -1597 -23547 -1528 -23530
rect -1470 -23530 -1230 -23492
rect -1470 -23547 -1401 -23530
rect -1597 -23564 -1570 -23547
rect -1726 -23580 -1570 -23564
rect -1428 -23564 -1401 -23547
rect -1367 -23564 -1333 -23530
rect -1299 -23547 -1230 -23530
rect -1172 -23530 -932 -23492
rect -1172 -23547 -1103 -23530
rect -1299 -23564 -1272 -23547
rect -1428 -23580 -1272 -23564
rect -1130 -23564 -1103 -23547
rect -1069 -23564 -1035 -23530
rect -1001 -23547 -932 -23530
rect -874 -23530 -634 -23492
rect -874 -23547 -805 -23530
rect -1001 -23564 -974 -23547
rect -1130 -23580 -974 -23564
rect -832 -23564 -805 -23547
rect -771 -23564 -737 -23530
rect -703 -23547 -634 -23530
rect -576 -23530 -336 -23492
rect -576 -23547 -507 -23530
rect -703 -23564 -676 -23547
rect -832 -23580 -676 -23564
rect -534 -23564 -507 -23547
rect -473 -23564 -439 -23530
rect -405 -23547 -336 -23530
rect -278 -23530 -38 -23492
rect -278 -23547 -209 -23530
rect -405 -23564 -378 -23547
rect -534 -23580 -378 -23564
rect -236 -23564 -209 -23547
rect -175 -23564 -141 -23530
rect -107 -23547 -38 -23530
rect 20 -23530 260 -23492
rect 20 -23547 89 -23530
rect -107 -23564 -80 -23547
rect -236 -23580 -80 -23564
rect 62 -23564 89 -23547
rect 123 -23564 157 -23530
rect 191 -23547 260 -23530
rect 318 -23530 558 -23492
rect 318 -23547 387 -23530
rect 191 -23564 218 -23547
rect 62 -23580 218 -23564
rect 360 -23564 387 -23547
rect 421 -23564 455 -23530
rect 489 -23547 558 -23530
rect 616 -23530 856 -23492
rect 2812 -23506 3400 -23490
rect 3830 -23490 3869 -23473
rect 3903 -23490 3937 -23456
rect 3971 -23490 4005 -23456
rect 4039 -23490 4073 -23456
rect 4107 -23490 4141 -23456
rect 4175 -23490 4209 -23456
rect 4243 -23490 4277 -23456
rect 4311 -23490 4345 -23456
rect 4379 -23473 4604 -23456
rect 4662 -23456 5622 -23418
rect 4662 -23473 4887 -23456
rect 4379 -23490 4418 -23473
rect 3830 -23506 4418 -23490
rect 4848 -23490 4887 -23473
rect 4921 -23490 4955 -23456
rect 4989 -23490 5023 -23456
rect 5057 -23490 5091 -23456
rect 5125 -23490 5159 -23456
rect 5193 -23490 5227 -23456
rect 5261 -23490 5295 -23456
rect 5329 -23490 5363 -23456
rect 5397 -23473 5622 -23456
rect 5680 -23456 6640 -23418
rect 5680 -23473 5905 -23456
rect 5397 -23490 5436 -23473
rect 4848 -23506 5436 -23490
rect 5866 -23490 5905 -23473
rect 5939 -23490 5973 -23456
rect 6007 -23490 6041 -23456
rect 6075 -23490 6109 -23456
rect 6143 -23490 6177 -23456
rect 6211 -23490 6245 -23456
rect 6279 -23490 6313 -23456
rect 6347 -23490 6381 -23456
rect 6415 -23473 6640 -23456
rect 6698 -23456 7658 -23418
rect 6698 -23473 6923 -23456
rect 6415 -23490 6454 -23473
rect 5866 -23506 6454 -23490
rect 6884 -23490 6923 -23473
rect 6957 -23490 6991 -23456
rect 7025 -23490 7059 -23456
rect 7093 -23490 7127 -23456
rect 7161 -23490 7195 -23456
rect 7229 -23490 7263 -23456
rect 7297 -23490 7331 -23456
rect 7365 -23490 7399 -23456
rect 7433 -23473 7658 -23456
rect 7716 -23456 8676 -23418
rect 7716 -23473 7941 -23456
rect 7433 -23490 7472 -23473
rect 6884 -23506 7472 -23490
rect 7902 -23490 7941 -23473
rect 7975 -23490 8009 -23456
rect 8043 -23490 8077 -23456
rect 8111 -23490 8145 -23456
rect 8179 -23490 8213 -23456
rect 8247 -23490 8281 -23456
rect 8315 -23490 8349 -23456
rect 8383 -23490 8417 -23456
rect 8451 -23473 8676 -23456
rect 8734 -23456 9694 -23418
rect 8734 -23473 8959 -23456
rect 8451 -23490 8490 -23473
rect 7902 -23506 8490 -23490
rect 8920 -23490 8959 -23473
rect 8993 -23490 9027 -23456
rect 9061 -23490 9095 -23456
rect 9129 -23490 9163 -23456
rect 9197 -23490 9231 -23456
rect 9265 -23490 9299 -23456
rect 9333 -23490 9367 -23456
rect 9401 -23490 9435 -23456
rect 9469 -23473 9694 -23456
rect 9752 -23456 10712 -23418
rect 9752 -23473 9977 -23456
rect 9469 -23490 9508 -23473
rect 8920 -23506 9508 -23490
rect 9938 -23490 9977 -23473
rect 10011 -23490 10045 -23456
rect 10079 -23490 10113 -23456
rect 10147 -23490 10181 -23456
rect 10215 -23490 10249 -23456
rect 10283 -23490 10317 -23456
rect 10351 -23490 10385 -23456
rect 10419 -23490 10453 -23456
rect 10487 -23473 10712 -23456
rect 10770 -23456 11730 -23418
rect 10770 -23473 10995 -23456
rect 10487 -23490 10526 -23473
rect 9938 -23506 10526 -23490
rect 10956 -23490 10995 -23473
rect 11029 -23490 11063 -23456
rect 11097 -23490 11131 -23456
rect 11165 -23490 11199 -23456
rect 11233 -23490 11267 -23456
rect 11301 -23490 11335 -23456
rect 11369 -23490 11403 -23456
rect 11437 -23490 11471 -23456
rect 11505 -23473 11730 -23456
rect 11788 -23456 12748 -23418
rect 11788 -23473 12013 -23456
rect 11505 -23490 11544 -23473
rect 10956 -23506 11544 -23490
rect 11974 -23490 12013 -23473
rect 12047 -23490 12081 -23456
rect 12115 -23490 12149 -23456
rect 12183 -23490 12217 -23456
rect 12251 -23490 12285 -23456
rect 12319 -23490 12353 -23456
rect 12387 -23490 12421 -23456
rect 12455 -23490 12489 -23456
rect 12523 -23473 12748 -23456
rect 12806 -23456 13766 -23418
rect 12806 -23473 13031 -23456
rect 12523 -23490 12562 -23473
rect 11974 -23506 12562 -23490
rect 12992 -23490 13031 -23473
rect 13065 -23490 13099 -23456
rect 13133 -23490 13167 -23456
rect 13201 -23490 13235 -23456
rect 13269 -23490 13303 -23456
rect 13337 -23490 13371 -23456
rect 13405 -23490 13439 -23456
rect 13473 -23490 13507 -23456
rect 13541 -23473 13766 -23456
rect 13824 -23456 14784 -23418
rect 13824 -23473 14049 -23456
rect 13541 -23490 13580 -23473
rect 12992 -23506 13580 -23490
rect 14010 -23490 14049 -23473
rect 14083 -23490 14117 -23456
rect 14151 -23490 14185 -23456
rect 14219 -23490 14253 -23456
rect 14287 -23490 14321 -23456
rect 14355 -23490 14389 -23456
rect 14423 -23490 14457 -23456
rect 14491 -23490 14525 -23456
rect 14559 -23473 14784 -23456
rect 14842 -23456 15802 -23418
rect 14842 -23473 15067 -23456
rect 14559 -23490 14598 -23473
rect 14010 -23506 14598 -23490
rect 15028 -23490 15067 -23473
rect 15101 -23490 15135 -23456
rect 15169 -23490 15203 -23456
rect 15237 -23490 15271 -23456
rect 15305 -23490 15339 -23456
rect 15373 -23490 15407 -23456
rect 15441 -23490 15475 -23456
rect 15509 -23490 15543 -23456
rect 15577 -23473 15802 -23456
rect 15860 -23456 16820 -23418
rect 15860 -23473 16085 -23456
rect 15577 -23490 15616 -23473
rect 15028 -23506 15616 -23490
rect 16046 -23490 16085 -23473
rect 16119 -23490 16153 -23456
rect 16187 -23490 16221 -23456
rect 16255 -23490 16289 -23456
rect 16323 -23490 16357 -23456
rect 16391 -23490 16425 -23456
rect 16459 -23490 16493 -23456
rect 16527 -23490 16561 -23456
rect 16595 -23473 16820 -23456
rect 16878 -23456 17838 -23418
rect 16878 -23473 17103 -23456
rect 16595 -23490 16634 -23473
rect 16046 -23506 16634 -23490
rect 17064 -23490 17103 -23473
rect 17137 -23490 17171 -23456
rect 17205 -23490 17239 -23456
rect 17273 -23490 17307 -23456
rect 17341 -23490 17375 -23456
rect 17409 -23490 17443 -23456
rect 17477 -23490 17511 -23456
rect 17545 -23490 17579 -23456
rect 17613 -23473 17838 -23456
rect 17896 -23456 18856 -23418
rect 17896 -23473 18121 -23456
rect 17613 -23490 17652 -23473
rect 17064 -23506 17652 -23490
rect 18082 -23490 18121 -23473
rect 18155 -23490 18189 -23456
rect 18223 -23490 18257 -23456
rect 18291 -23490 18325 -23456
rect 18359 -23490 18393 -23456
rect 18427 -23490 18461 -23456
rect 18495 -23490 18529 -23456
rect 18563 -23490 18597 -23456
rect 18631 -23473 18856 -23456
rect 18914 -23456 19874 -23418
rect 18914 -23473 19139 -23456
rect 18631 -23490 18670 -23473
rect 18082 -23506 18670 -23490
rect 19100 -23490 19139 -23473
rect 19173 -23490 19207 -23456
rect 19241 -23490 19275 -23456
rect 19309 -23490 19343 -23456
rect 19377 -23490 19411 -23456
rect 19445 -23490 19479 -23456
rect 19513 -23490 19547 -23456
rect 19581 -23490 19615 -23456
rect 19649 -23473 19874 -23456
rect 19932 -23456 20892 -23418
rect 19932 -23473 20157 -23456
rect 19649 -23490 19688 -23473
rect 19100 -23506 19688 -23490
rect 20118 -23490 20157 -23473
rect 20191 -23490 20225 -23456
rect 20259 -23490 20293 -23456
rect 20327 -23490 20361 -23456
rect 20395 -23490 20429 -23456
rect 20463 -23490 20497 -23456
rect 20531 -23490 20565 -23456
rect 20599 -23490 20633 -23456
rect 20667 -23473 20892 -23456
rect 20950 -23456 21910 -23418
rect 20950 -23473 21175 -23456
rect 20667 -23490 20706 -23473
rect 20118 -23506 20706 -23490
rect 21136 -23490 21175 -23473
rect 21209 -23490 21243 -23456
rect 21277 -23490 21311 -23456
rect 21345 -23490 21379 -23456
rect 21413 -23490 21447 -23456
rect 21481 -23490 21515 -23456
rect 21549 -23490 21583 -23456
rect 21617 -23490 21651 -23456
rect 21685 -23473 21910 -23456
rect 21968 -23456 22928 -23418
rect 21968 -23473 22193 -23456
rect 21685 -23490 21724 -23473
rect 21136 -23506 21724 -23490
rect 22154 -23490 22193 -23473
rect 22227 -23490 22261 -23456
rect 22295 -23490 22329 -23456
rect 22363 -23490 22397 -23456
rect 22431 -23490 22465 -23456
rect 22499 -23490 22533 -23456
rect 22567 -23490 22601 -23456
rect 22635 -23490 22669 -23456
rect 22703 -23473 22928 -23456
rect 22703 -23490 22742 -23473
rect 22154 -23506 22742 -23490
rect 616 -23547 685 -23530
rect 489 -23564 516 -23547
rect 360 -23580 516 -23564
rect 658 -23564 685 -23547
rect 719 -23564 753 -23530
rect 787 -23547 856 -23530
rect 787 -23564 814 -23547
rect 658 -23580 814 -23564
rect -9173 -23933 -8585 -23917
rect -9173 -23950 -9134 -23933
rect -9359 -23967 -9134 -23950
rect -9100 -23967 -9066 -23933
rect -9032 -23967 -8998 -23933
rect -8964 -23967 -8930 -23933
rect -8896 -23967 -8862 -23933
rect -8828 -23967 -8794 -23933
rect -8760 -23967 -8726 -23933
rect -8692 -23967 -8658 -23933
rect -8624 -23950 -8585 -23933
rect -8155 -23933 -7567 -23917
rect -8155 -23950 -8116 -23933
rect -8624 -23967 -8399 -23950
rect -9359 -24005 -8399 -23967
rect -8341 -23967 -8116 -23950
rect -8082 -23967 -8048 -23933
rect -8014 -23967 -7980 -23933
rect -7946 -23967 -7912 -23933
rect -7878 -23967 -7844 -23933
rect -7810 -23967 -7776 -23933
rect -7742 -23967 -7708 -23933
rect -7674 -23967 -7640 -23933
rect -7606 -23950 -7567 -23933
rect -7137 -23933 -6549 -23917
rect -7137 -23950 -7098 -23933
rect -7606 -23967 -7381 -23950
rect -8341 -24005 -7381 -23967
rect -7323 -23967 -7098 -23950
rect -7064 -23967 -7030 -23933
rect -6996 -23967 -6962 -23933
rect -6928 -23967 -6894 -23933
rect -6860 -23967 -6826 -23933
rect -6792 -23967 -6758 -23933
rect -6724 -23967 -6690 -23933
rect -6656 -23967 -6622 -23933
rect -6588 -23950 -6549 -23933
rect -6119 -23933 -5531 -23917
rect -6119 -23950 -6080 -23933
rect -6588 -23967 -6363 -23950
rect -7323 -24005 -6363 -23967
rect -6305 -23967 -6080 -23950
rect -6046 -23967 -6012 -23933
rect -5978 -23967 -5944 -23933
rect -5910 -23967 -5876 -23933
rect -5842 -23967 -5808 -23933
rect -5774 -23967 -5740 -23933
rect -5706 -23967 -5672 -23933
rect -5638 -23967 -5604 -23933
rect -5570 -23950 -5531 -23933
rect -5101 -23933 -4513 -23917
rect -5101 -23950 -5062 -23933
rect -5570 -23967 -5345 -23950
rect -6305 -24005 -5345 -23967
rect -5287 -23967 -5062 -23950
rect -5028 -23967 -4994 -23933
rect -4960 -23967 -4926 -23933
rect -4892 -23967 -4858 -23933
rect -4824 -23967 -4790 -23933
rect -4756 -23967 -4722 -23933
rect -4688 -23967 -4654 -23933
rect -4620 -23967 -4586 -23933
rect -4552 -23950 -4513 -23933
rect -4083 -23933 -3495 -23917
rect -4083 -23950 -4044 -23933
rect -4552 -23967 -4327 -23950
rect -5287 -24005 -4327 -23967
rect -4269 -23967 -4044 -23950
rect -4010 -23967 -3976 -23933
rect -3942 -23967 -3908 -23933
rect -3874 -23967 -3840 -23933
rect -3806 -23967 -3772 -23933
rect -3738 -23967 -3704 -23933
rect -3670 -23967 -3636 -23933
rect -3602 -23967 -3568 -23933
rect -3534 -23950 -3495 -23933
rect -2324 -23932 -2168 -23916
rect -2324 -23949 -2297 -23932
rect -3534 -23967 -3309 -23950
rect -4269 -24005 -3309 -23967
rect -2366 -23966 -2297 -23949
rect -2263 -23966 -2229 -23932
rect -2195 -23949 -2168 -23932
rect -2026 -23932 -1870 -23916
rect -2026 -23949 -1999 -23932
rect -2195 -23966 -2126 -23949
rect -2366 -24004 -2126 -23966
rect -2068 -23966 -1999 -23949
rect -1965 -23966 -1931 -23932
rect -1897 -23949 -1870 -23932
rect -1728 -23932 -1572 -23916
rect -1728 -23949 -1701 -23932
rect -1897 -23966 -1828 -23949
rect -2068 -24004 -1828 -23966
rect -1770 -23966 -1701 -23949
rect -1667 -23966 -1633 -23932
rect -1599 -23949 -1572 -23932
rect -1430 -23932 -1274 -23916
rect -1430 -23949 -1403 -23932
rect -1599 -23966 -1530 -23949
rect -1770 -24004 -1530 -23966
rect -1472 -23966 -1403 -23949
rect -1369 -23966 -1335 -23932
rect -1301 -23949 -1274 -23932
rect -1132 -23932 -976 -23916
rect -1132 -23949 -1105 -23932
rect -1301 -23966 -1232 -23949
rect -1472 -24004 -1232 -23966
rect -1174 -23966 -1105 -23949
rect -1071 -23966 -1037 -23932
rect -1003 -23949 -976 -23932
rect -834 -23932 -678 -23916
rect -834 -23949 -807 -23932
rect -1003 -23966 -934 -23949
rect -1174 -24004 -934 -23966
rect -876 -23966 -807 -23949
rect -773 -23966 -739 -23932
rect -705 -23949 -678 -23932
rect -536 -23932 -380 -23916
rect -536 -23949 -509 -23932
rect -705 -23966 -636 -23949
rect -876 -24004 -636 -23966
rect -578 -23966 -509 -23949
rect -475 -23966 -441 -23932
rect -407 -23949 -380 -23932
rect -238 -23932 -82 -23916
rect -238 -23949 -211 -23932
rect -407 -23966 -338 -23949
rect -578 -24004 -338 -23966
rect -280 -23966 -211 -23949
rect -177 -23966 -143 -23932
rect -109 -23949 -82 -23932
rect 60 -23932 216 -23916
rect 60 -23949 87 -23932
rect -109 -23966 -40 -23949
rect -280 -24004 -40 -23966
rect 18 -23966 87 -23949
rect 121 -23966 155 -23932
rect 189 -23949 216 -23932
rect 358 -23932 514 -23916
rect 358 -23949 385 -23932
rect 189 -23966 258 -23949
rect 18 -24004 258 -23966
rect 316 -23966 385 -23949
rect 419 -23966 453 -23932
rect 487 -23949 514 -23932
rect 656 -23932 812 -23916
rect 656 -23949 683 -23932
rect 487 -23966 556 -23949
rect 316 -24004 556 -23966
rect 614 -23966 683 -23949
rect 717 -23966 751 -23932
rect 785 -23949 812 -23932
rect 785 -23966 854 -23949
rect 614 -24004 854 -23966
rect 2812 -23980 3400 -23964
rect 2812 -23997 2851 -23980
rect 2626 -24014 2851 -23997
rect 2885 -24014 2919 -23980
rect 2953 -24014 2987 -23980
rect 3021 -24014 3055 -23980
rect 3089 -24014 3123 -23980
rect 3157 -24014 3191 -23980
rect 3225 -24014 3259 -23980
rect 3293 -24014 3327 -23980
rect 3361 -23997 3400 -23980
rect 3830 -23980 4418 -23964
rect 3830 -23997 3869 -23980
rect 3361 -24014 3586 -23997
rect 2626 -24052 3586 -24014
rect 3644 -24014 3869 -23997
rect 3903 -24014 3937 -23980
rect 3971 -24014 4005 -23980
rect 4039 -24014 4073 -23980
rect 4107 -24014 4141 -23980
rect 4175 -24014 4209 -23980
rect 4243 -24014 4277 -23980
rect 4311 -24014 4345 -23980
rect 4379 -23997 4418 -23980
rect 4848 -23980 5436 -23964
rect 4848 -23997 4887 -23980
rect 4379 -24014 4604 -23997
rect 3644 -24052 4604 -24014
rect 4662 -24014 4887 -23997
rect 4921 -24014 4955 -23980
rect 4989 -24014 5023 -23980
rect 5057 -24014 5091 -23980
rect 5125 -24014 5159 -23980
rect 5193 -24014 5227 -23980
rect 5261 -24014 5295 -23980
rect 5329 -24014 5363 -23980
rect 5397 -23997 5436 -23980
rect 5866 -23980 6454 -23964
rect 5866 -23997 5905 -23980
rect 5397 -24014 5622 -23997
rect 4662 -24052 5622 -24014
rect 5680 -24014 5905 -23997
rect 5939 -24014 5973 -23980
rect 6007 -24014 6041 -23980
rect 6075 -24014 6109 -23980
rect 6143 -24014 6177 -23980
rect 6211 -24014 6245 -23980
rect 6279 -24014 6313 -23980
rect 6347 -24014 6381 -23980
rect 6415 -23997 6454 -23980
rect 6884 -23980 7472 -23964
rect 6884 -23997 6923 -23980
rect 6415 -24014 6640 -23997
rect 5680 -24052 6640 -24014
rect 6698 -24014 6923 -23997
rect 6957 -24014 6991 -23980
rect 7025 -24014 7059 -23980
rect 7093 -24014 7127 -23980
rect 7161 -24014 7195 -23980
rect 7229 -24014 7263 -23980
rect 7297 -24014 7331 -23980
rect 7365 -24014 7399 -23980
rect 7433 -23997 7472 -23980
rect 7902 -23980 8490 -23964
rect 7902 -23997 7941 -23980
rect 7433 -24014 7658 -23997
rect 6698 -24052 7658 -24014
rect 7716 -24014 7941 -23997
rect 7975 -24014 8009 -23980
rect 8043 -24014 8077 -23980
rect 8111 -24014 8145 -23980
rect 8179 -24014 8213 -23980
rect 8247 -24014 8281 -23980
rect 8315 -24014 8349 -23980
rect 8383 -24014 8417 -23980
rect 8451 -23997 8490 -23980
rect 8920 -23980 9508 -23964
rect 8920 -23997 8959 -23980
rect 8451 -24014 8676 -23997
rect 7716 -24052 8676 -24014
rect 8734 -24014 8959 -23997
rect 8993 -24014 9027 -23980
rect 9061 -24014 9095 -23980
rect 9129 -24014 9163 -23980
rect 9197 -24014 9231 -23980
rect 9265 -24014 9299 -23980
rect 9333 -24014 9367 -23980
rect 9401 -24014 9435 -23980
rect 9469 -23997 9508 -23980
rect 9938 -23980 10526 -23964
rect 9938 -23997 9977 -23980
rect 9469 -24014 9694 -23997
rect 8734 -24052 9694 -24014
rect 9752 -24014 9977 -23997
rect 10011 -24014 10045 -23980
rect 10079 -24014 10113 -23980
rect 10147 -24014 10181 -23980
rect 10215 -24014 10249 -23980
rect 10283 -24014 10317 -23980
rect 10351 -24014 10385 -23980
rect 10419 -24014 10453 -23980
rect 10487 -23997 10526 -23980
rect 10956 -23980 11544 -23964
rect 10956 -23997 10995 -23980
rect 10487 -24014 10712 -23997
rect 9752 -24052 10712 -24014
rect 10770 -24014 10995 -23997
rect 11029 -24014 11063 -23980
rect 11097 -24014 11131 -23980
rect 11165 -24014 11199 -23980
rect 11233 -24014 11267 -23980
rect 11301 -24014 11335 -23980
rect 11369 -24014 11403 -23980
rect 11437 -24014 11471 -23980
rect 11505 -23997 11544 -23980
rect 11974 -23980 12562 -23964
rect 11974 -23997 12013 -23980
rect 11505 -24014 11730 -23997
rect 10770 -24052 11730 -24014
rect 11788 -24014 12013 -23997
rect 12047 -24014 12081 -23980
rect 12115 -24014 12149 -23980
rect 12183 -24014 12217 -23980
rect 12251 -24014 12285 -23980
rect 12319 -24014 12353 -23980
rect 12387 -24014 12421 -23980
rect 12455 -24014 12489 -23980
rect 12523 -23997 12562 -23980
rect 12992 -23980 13580 -23964
rect 12992 -23997 13031 -23980
rect 12523 -24014 12748 -23997
rect 11788 -24052 12748 -24014
rect 12806 -24014 13031 -23997
rect 13065 -24014 13099 -23980
rect 13133 -24014 13167 -23980
rect 13201 -24014 13235 -23980
rect 13269 -24014 13303 -23980
rect 13337 -24014 13371 -23980
rect 13405 -24014 13439 -23980
rect 13473 -24014 13507 -23980
rect 13541 -23997 13580 -23980
rect 14010 -23980 14598 -23964
rect 14010 -23997 14049 -23980
rect 13541 -24014 13766 -23997
rect 12806 -24052 13766 -24014
rect 13824 -24014 14049 -23997
rect 14083 -24014 14117 -23980
rect 14151 -24014 14185 -23980
rect 14219 -24014 14253 -23980
rect 14287 -24014 14321 -23980
rect 14355 -24014 14389 -23980
rect 14423 -24014 14457 -23980
rect 14491 -24014 14525 -23980
rect 14559 -23997 14598 -23980
rect 15028 -23980 15616 -23964
rect 15028 -23997 15067 -23980
rect 14559 -24014 14784 -23997
rect 13824 -24052 14784 -24014
rect 14842 -24014 15067 -23997
rect 15101 -24014 15135 -23980
rect 15169 -24014 15203 -23980
rect 15237 -24014 15271 -23980
rect 15305 -24014 15339 -23980
rect 15373 -24014 15407 -23980
rect 15441 -24014 15475 -23980
rect 15509 -24014 15543 -23980
rect 15577 -23997 15616 -23980
rect 16046 -23980 16634 -23964
rect 16046 -23997 16085 -23980
rect 15577 -24014 15802 -23997
rect 14842 -24052 15802 -24014
rect 15860 -24014 16085 -23997
rect 16119 -24014 16153 -23980
rect 16187 -24014 16221 -23980
rect 16255 -24014 16289 -23980
rect 16323 -24014 16357 -23980
rect 16391 -24014 16425 -23980
rect 16459 -24014 16493 -23980
rect 16527 -24014 16561 -23980
rect 16595 -23997 16634 -23980
rect 17064 -23980 17652 -23964
rect 17064 -23997 17103 -23980
rect 16595 -24014 16820 -23997
rect 15860 -24052 16820 -24014
rect 16878 -24014 17103 -23997
rect 17137 -24014 17171 -23980
rect 17205 -24014 17239 -23980
rect 17273 -24014 17307 -23980
rect 17341 -24014 17375 -23980
rect 17409 -24014 17443 -23980
rect 17477 -24014 17511 -23980
rect 17545 -24014 17579 -23980
rect 17613 -23997 17652 -23980
rect 18082 -23980 18670 -23964
rect 18082 -23997 18121 -23980
rect 17613 -24014 17838 -23997
rect 16878 -24052 17838 -24014
rect 17896 -24014 18121 -23997
rect 18155 -24014 18189 -23980
rect 18223 -24014 18257 -23980
rect 18291 -24014 18325 -23980
rect 18359 -24014 18393 -23980
rect 18427 -24014 18461 -23980
rect 18495 -24014 18529 -23980
rect 18563 -24014 18597 -23980
rect 18631 -23997 18670 -23980
rect 19100 -23980 19688 -23964
rect 19100 -23997 19139 -23980
rect 18631 -24014 18856 -23997
rect 17896 -24052 18856 -24014
rect 18914 -24014 19139 -23997
rect 19173 -24014 19207 -23980
rect 19241 -24014 19275 -23980
rect 19309 -24014 19343 -23980
rect 19377 -24014 19411 -23980
rect 19445 -24014 19479 -23980
rect 19513 -24014 19547 -23980
rect 19581 -24014 19615 -23980
rect 19649 -23997 19688 -23980
rect 20118 -23980 20706 -23964
rect 20118 -23997 20157 -23980
rect 19649 -24014 19874 -23997
rect 18914 -24052 19874 -24014
rect 19932 -24014 20157 -23997
rect 20191 -24014 20225 -23980
rect 20259 -24014 20293 -23980
rect 20327 -24014 20361 -23980
rect 20395 -24014 20429 -23980
rect 20463 -24014 20497 -23980
rect 20531 -24014 20565 -23980
rect 20599 -24014 20633 -23980
rect 20667 -23997 20706 -23980
rect 21136 -23980 21724 -23964
rect 21136 -23997 21175 -23980
rect 20667 -24014 20892 -23997
rect 19932 -24052 20892 -24014
rect 20950 -24014 21175 -23997
rect 21209 -24014 21243 -23980
rect 21277 -24014 21311 -23980
rect 21345 -24014 21379 -23980
rect 21413 -24014 21447 -23980
rect 21481 -24014 21515 -23980
rect 21549 -24014 21583 -23980
rect 21617 -24014 21651 -23980
rect 21685 -23997 21724 -23980
rect 22154 -23980 22742 -23964
rect 22154 -23997 22193 -23980
rect 21685 -24014 21910 -23997
rect 20950 -24052 21910 -24014
rect 21968 -24014 22193 -23997
rect 22227 -24014 22261 -23980
rect 22295 -24014 22329 -23980
rect 22363 -24014 22397 -23980
rect 22431 -24014 22465 -23980
rect 22499 -24014 22533 -23980
rect 22567 -24014 22601 -23980
rect 22635 -24014 22669 -23980
rect 22703 -23997 22742 -23980
rect 22703 -24014 22928 -23997
rect 21968 -24052 22928 -24014
rect -9359 -24643 -8399 -24605
rect -9359 -24660 -9134 -24643
rect -9173 -24677 -9134 -24660
rect -9100 -24677 -9066 -24643
rect -9032 -24677 -8998 -24643
rect -8964 -24677 -8930 -24643
rect -8896 -24677 -8862 -24643
rect -8828 -24677 -8794 -24643
rect -8760 -24677 -8726 -24643
rect -8692 -24677 -8658 -24643
rect -8624 -24660 -8399 -24643
rect -8341 -24643 -7381 -24605
rect -8341 -24660 -8116 -24643
rect -8624 -24677 -8585 -24660
rect -9173 -24693 -8585 -24677
rect -8155 -24677 -8116 -24660
rect -8082 -24677 -8048 -24643
rect -8014 -24677 -7980 -24643
rect -7946 -24677 -7912 -24643
rect -7878 -24677 -7844 -24643
rect -7810 -24677 -7776 -24643
rect -7742 -24677 -7708 -24643
rect -7674 -24677 -7640 -24643
rect -7606 -24660 -7381 -24643
rect -7323 -24643 -6363 -24605
rect -7323 -24660 -7098 -24643
rect -7606 -24677 -7567 -24660
rect -8155 -24693 -7567 -24677
rect -7137 -24677 -7098 -24660
rect -7064 -24677 -7030 -24643
rect -6996 -24677 -6962 -24643
rect -6928 -24677 -6894 -24643
rect -6860 -24677 -6826 -24643
rect -6792 -24677 -6758 -24643
rect -6724 -24677 -6690 -24643
rect -6656 -24677 -6622 -24643
rect -6588 -24660 -6363 -24643
rect -6305 -24643 -5345 -24605
rect -6305 -24660 -6080 -24643
rect -6588 -24677 -6549 -24660
rect -7137 -24693 -6549 -24677
rect -6119 -24677 -6080 -24660
rect -6046 -24677 -6012 -24643
rect -5978 -24677 -5944 -24643
rect -5910 -24677 -5876 -24643
rect -5842 -24677 -5808 -24643
rect -5774 -24677 -5740 -24643
rect -5706 -24677 -5672 -24643
rect -5638 -24677 -5604 -24643
rect -5570 -24660 -5345 -24643
rect -5287 -24643 -4327 -24605
rect -5287 -24660 -5062 -24643
rect -5570 -24677 -5531 -24660
rect -6119 -24693 -5531 -24677
rect -5101 -24677 -5062 -24660
rect -5028 -24677 -4994 -24643
rect -4960 -24677 -4926 -24643
rect -4892 -24677 -4858 -24643
rect -4824 -24677 -4790 -24643
rect -4756 -24677 -4722 -24643
rect -4688 -24677 -4654 -24643
rect -4620 -24677 -4586 -24643
rect -4552 -24660 -4327 -24643
rect -4269 -24643 -3309 -24605
rect -4269 -24660 -4044 -24643
rect -4552 -24677 -4513 -24660
rect -5101 -24693 -4513 -24677
rect -4083 -24677 -4044 -24660
rect -4010 -24677 -3976 -24643
rect -3942 -24677 -3908 -24643
rect -3874 -24677 -3840 -24643
rect -3806 -24677 -3772 -24643
rect -3738 -24677 -3704 -24643
rect -3670 -24677 -3636 -24643
rect -3602 -24677 -3568 -24643
rect -3534 -24660 -3309 -24643
rect -2366 -24642 -2126 -24604
rect -2366 -24659 -2297 -24642
rect -3534 -24677 -3495 -24660
rect -4083 -24693 -3495 -24677
rect -2324 -24676 -2297 -24659
rect -2263 -24676 -2229 -24642
rect -2195 -24659 -2126 -24642
rect -2068 -24642 -1828 -24604
rect -2068 -24659 -1999 -24642
rect -2195 -24676 -2168 -24659
rect -2324 -24692 -2168 -24676
rect -2026 -24676 -1999 -24659
rect -1965 -24676 -1931 -24642
rect -1897 -24659 -1828 -24642
rect -1770 -24642 -1530 -24604
rect -1770 -24659 -1701 -24642
rect -1897 -24676 -1870 -24659
rect -2026 -24692 -1870 -24676
rect -1728 -24676 -1701 -24659
rect -1667 -24676 -1633 -24642
rect -1599 -24659 -1530 -24642
rect -1472 -24642 -1232 -24604
rect -1472 -24659 -1403 -24642
rect -1599 -24676 -1572 -24659
rect -1728 -24692 -1572 -24676
rect -1430 -24676 -1403 -24659
rect -1369 -24676 -1335 -24642
rect -1301 -24659 -1232 -24642
rect -1174 -24642 -934 -24604
rect -1174 -24659 -1105 -24642
rect -1301 -24676 -1274 -24659
rect -1430 -24692 -1274 -24676
rect -1132 -24676 -1105 -24659
rect -1071 -24676 -1037 -24642
rect -1003 -24659 -934 -24642
rect -876 -24642 -636 -24604
rect -876 -24659 -807 -24642
rect -1003 -24676 -976 -24659
rect -1132 -24692 -976 -24676
rect -834 -24676 -807 -24659
rect -773 -24676 -739 -24642
rect -705 -24659 -636 -24642
rect -578 -24642 -338 -24604
rect -578 -24659 -509 -24642
rect -705 -24676 -678 -24659
rect -834 -24692 -678 -24676
rect -536 -24676 -509 -24659
rect -475 -24676 -441 -24642
rect -407 -24659 -338 -24642
rect -280 -24642 -40 -24604
rect -280 -24659 -211 -24642
rect -407 -24676 -380 -24659
rect -536 -24692 -380 -24676
rect -238 -24676 -211 -24659
rect -177 -24676 -143 -24642
rect -109 -24659 -40 -24642
rect 18 -24642 258 -24604
rect 18 -24659 87 -24642
rect -109 -24676 -82 -24659
rect -238 -24692 -82 -24676
rect 60 -24676 87 -24659
rect 121 -24676 155 -24642
rect 189 -24659 258 -24642
rect 316 -24642 556 -24604
rect 316 -24659 385 -24642
rect 189 -24676 216 -24659
rect 60 -24692 216 -24676
rect 358 -24676 385 -24659
rect 419 -24676 453 -24642
rect 487 -24659 556 -24642
rect 614 -24642 854 -24604
rect 614 -24659 683 -24642
rect 487 -24676 514 -24659
rect 358 -24692 514 -24676
rect 656 -24676 683 -24659
rect 717 -24676 751 -24642
rect 785 -24659 854 -24642
rect 785 -24676 812 -24659
rect 656 -24692 812 -24676
rect 2626 -24690 3586 -24652
rect 2626 -24707 2851 -24690
rect 2812 -24724 2851 -24707
rect 2885 -24724 2919 -24690
rect 2953 -24724 2987 -24690
rect 3021 -24724 3055 -24690
rect 3089 -24724 3123 -24690
rect 3157 -24724 3191 -24690
rect 3225 -24724 3259 -24690
rect 3293 -24724 3327 -24690
rect 3361 -24707 3586 -24690
rect 3644 -24690 4604 -24652
rect 3644 -24707 3869 -24690
rect 3361 -24724 3400 -24707
rect 2812 -24740 3400 -24724
rect 3830 -24724 3869 -24707
rect 3903 -24724 3937 -24690
rect 3971 -24724 4005 -24690
rect 4039 -24724 4073 -24690
rect 4107 -24724 4141 -24690
rect 4175 -24724 4209 -24690
rect 4243 -24724 4277 -24690
rect 4311 -24724 4345 -24690
rect 4379 -24707 4604 -24690
rect 4662 -24690 5622 -24652
rect 4662 -24707 4887 -24690
rect 4379 -24724 4418 -24707
rect 3830 -24740 4418 -24724
rect 4848 -24724 4887 -24707
rect 4921 -24724 4955 -24690
rect 4989 -24724 5023 -24690
rect 5057 -24724 5091 -24690
rect 5125 -24724 5159 -24690
rect 5193 -24724 5227 -24690
rect 5261 -24724 5295 -24690
rect 5329 -24724 5363 -24690
rect 5397 -24707 5622 -24690
rect 5680 -24690 6640 -24652
rect 5680 -24707 5905 -24690
rect 5397 -24724 5436 -24707
rect 4848 -24740 5436 -24724
rect 5866 -24724 5905 -24707
rect 5939 -24724 5973 -24690
rect 6007 -24724 6041 -24690
rect 6075 -24724 6109 -24690
rect 6143 -24724 6177 -24690
rect 6211 -24724 6245 -24690
rect 6279 -24724 6313 -24690
rect 6347 -24724 6381 -24690
rect 6415 -24707 6640 -24690
rect 6698 -24690 7658 -24652
rect 6698 -24707 6923 -24690
rect 6415 -24724 6454 -24707
rect 5866 -24740 6454 -24724
rect 6884 -24724 6923 -24707
rect 6957 -24724 6991 -24690
rect 7025 -24724 7059 -24690
rect 7093 -24724 7127 -24690
rect 7161 -24724 7195 -24690
rect 7229 -24724 7263 -24690
rect 7297 -24724 7331 -24690
rect 7365 -24724 7399 -24690
rect 7433 -24707 7658 -24690
rect 7716 -24690 8676 -24652
rect 7716 -24707 7941 -24690
rect 7433 -24724 7472 -24707
rect 6884 -24740 7472 -24724
rect 7902 -24724 7941 -24707
rect 7975 -24724 8009 -24690
rect 8043 -24724 8077 -24690
rect 8111 -24724 8145 -24690
rect 8179 -24724 8213 -24690
rect 8247 -24724 8281 -24690
rect 8315 -24724 8349 -24690
rect 8383 -24724 8417 -24690
rect 8451 -24707 8676 -24690
rect 8734 -24690 9694 -24652
rect 8734 -24707 8959 -24690
rect 8451 -24724 8490 -24707
rect 7902 -24740 8490 -24724
rect 8920 -24724 8959 -24707
rect 8993 -24724 9027 -24690
rect 9061 -24724 9095 -24690
rect 9129 -24724 9163 -24690
rect 9197 -24724 9231 -24690
rect 9265 -24724 9299 -24690
rect 9333 -24724 9367 -24690
rect 9401 -24724 9435 -24690
rect 9469 -24707 9694 -24690
rect 9752 -24690 10712 -24652
rect 9752 -24707 9977 -24690
rect 9469 -24724 9508 -24707
rect 8920 -24740 9508 -24724
rect 9938 -24724 9977 -24707
rect 10011 -24724 10045 -24690
rect 10079 -24724 10113 -24690
rect 10147 -24724 10181 -24690
rect 10215 -24724 10249 -24690
rect 10283 -24724 10317 -24690
rect 10351 -24724 10385 -24690
rect 10419 -24724 10453 -24690
rect 10487 -24707 10712 -24690
rect 10770 -24690 11730 -24652
rect 10770 -24707 10995 -24690
rect 10487 -24724 10526 -24707
rect 9938 -24740 10526 -24724
rect 10956 -24724 10995 -24707
rect 11029 -24724 11063 -24690
rect 11097 -24724 11131 -24690
rect 11165 -24724 11199 -24690
rect 11233 -24724 11267 -24690
rect 11301 -24724 11335 -24690
rect 11369 -24724 11403 -24690
rect 11437 -24724 11471 -24690
rect 11505 -24707 11730 -24690
rect 11788 -24690 12748 -24652
rect 11788 -24707 12013 -24690
rect 11505 -24724 11544 -24707
rect 10956 -24740 11544 -24724
rect 11974 -24724 12013 -24707
rect 12047 -24724 12081 -24690
rect 12115 -24724 12149 -24690
rect 12183 -24724 12217 -24690
rect 12251 -24724 12285 -24690
rect 12319 -24724 12353 -24690
rect 12387 -24724 12421 -24690
rect 12455 -24724 12489 -24690
rect 12523 -24707 12748 -24690
rect 12806 -24690 13766 -24652
rect 12806 -24707 13031 -24690
rect 12523 -24724 12562 -24707
rect 11974 -24740 12562 -24724
rect 12992 -24724 13031 -24707
rect 13065 -24724 13099 -24690
rect 13133 -24724 13167 -24690
rect 13201 -24724 13235 -24690
rect 13269 -24724 13303 -24690
rect 13337 -24724 13371 -24690
rect 13405 -24724 13439 -24690
rect 13473 -24724 13507 -24690
rect 13541 -24707 13766 -24690
rect 13824 -24690 14784 -24652
rect 13824 -24707 14049 -24690
rect 13541 -24724 13580 -24707
rect 12992 -24740 13580 -24724
rect 14010 -24724 14049 -24707
rect 14083 -24724 14117 -24690
rect 14151 -24724 14185 -24690
rect 14219 -24724 14253 -24690
rect 14287 -24724 14321 -24690
rect 14355 -24724 14389 -24690
rect 14423 -24724 14457 -24690
rect 14491 -24724 14525 -24690
rect 14559 -24707 14784 -24690
rect 14842 -24690 15802 -24652
rect 14842 -24707 15067 -24690
rect 14559 -24724 14598 -24707
rect 14010 -24740 14598 -24724
rect 15028 -24724 15067 -24707
rect 15101 -24724 15135 -24690
rect 15169 -24724 15203 -24690
rect 15237 -24724 15271 -24690
rect 15305 -24724 15339 -24690
rect 15373 -24724 15407 -24690
rect 15441 -24724 15475 -24690
rect 15509 -24724 15543 -24690
rect 15577 -24707 15802 -24690
rect 15860 -24690 16820 -24652
rect 15860 -24707 16085 -24690
rect 15577 -24724 15616 -24707
rect 15028 -24740 15616 -24724
rect 16046 -24724 16085 -24707
rect 16119 -24724 16153 -24690
rect 16187 -24724 16221 -24690
rect 16255 -24724 16289 -24690
rect 16323 -24724 16357 -24690
rect 16391 -24724 16425 -24690
rect 16459 -24724 16493 -24690
rect 16527 -24724 16561 -24690
rect 16595 -24707 16820 -24690
rect 16878 -24690 17838 -24652
rect 16878 -24707 17103 -24690
rect 16595 -24724 16634 -24707
rect 16046 -24740 16634 -24724
rect 17064 -24724 17103 -24707
rect 17137 -24724 17171 -24690
rect 17205 -24724 17239 -24690
rect 17273 -24724 17307 -24690
rect 17341 -24724 17375 -24690
rect 17409 -24724 17443 -24690
rect 17477 -24724 17511 -24690
rect 17545 -24724 17579 -24690
rect 17613 -24707 17838 -24690
rect 17896 -24690 18856 -24652
rect 17896 -24707 18121 -24690
rect 17613 -24724 17652 -24707
rect 17064 -24740 17652 -24724
rect 18082 -24724 18121 -24707
rect 18155 -24724 18189 -24690
rect 18223 -24724 18257 -24690
rect 18291 -24724 18325 -24690
rect 18359 -24724 18393 -24690
rect 18427 -24724 18461 -24690
rect 18495 -24724 18529 -24690
rect 18563 -24724 18597 -24690
rect 18631 -24707 18856 -24690
rect 18914 -24690 19874 -24652
rect 18914 -24707 19139 -24690
rect 18631 -24724 18670 -24707
rect 18082 -24740 18670 -24724
rect 19100 -24724 19139 -24707
rect 19173 -24724 19207 -24690
rect 19241 -24724 19275 -24690
rect 19309 -24724 19343 -24690
rect 19377 -24724 19411 -24690
rect 19445 -24724 19479 -24690
rect 19513 -24724 19547 -24690
rect 19581 -24724 19615 -24690
rect 19649 -24707 19874 -24690
rect 19932 -24690 20892 -24652
rect 19932 -24707 20157 -24690
rect 19649 -24724 19688 -24707
rect 19100 -24740 19688 -24724
rect 20118 -24724 20157 -24707
rect 20191 -24724 20225 -24690
rect 20259 -24724 20293 -24690
rect 20327 -24724 20361 -24690
rect 20395 -24724 20429 -24690
rect 20463 -24724 20497 -24690
rect 20531 -24724 20565 -24690
rect 20599 -24724 20633 -24690
rect 20667 -24707 20892 -24690
rect 20950 -24690 21910 -24652
rect 20950 -24707 21175 -24690
rect 20667 -24724 20706 -24707
rect 20118 -24740 20706 -24724
rect 21136 -24724 21175 -24707
rect 21209 -24724 21243 -24690
rect 21277 -24724 21311 -24690
rect 21345 -24724 21379 -24690
rect 21413 -24724 21447 -24690
rect 21481 -24724 21515 -24690
rect 21549 -24724 21583 -24690
rect 21617 -24724 21651 -24690
rect 21685 -24707 21910 -24690
rect 21968 -24690 22928 -24652
rect 21968 -24707 22193 -24690
rect 21685 -24724 21724 -24707
rect 21136 -24740 21724 -24724
rect 22154 -24724 22193 -24707
rect 22227 -24724 22261 -24690
rect 22295 -24724 22329 -24690
rect 22363 -24724 22397 -24690
rect 22431 -24724 22465 -24690
rect 22499 -24724 22533 -24690
rect 22567 -24724 22601 -24690
rect 22635 -24724 22669 -24690
rect 22703 -24707 22928 -24690
rect 22703 -24724 22742 -24707
rect 22154 -24740 22742 -24724
rect -9174 -25046 -8586 -25030
rect -9174 -25063 -9135 -25046
rect -9360 -25080 -9135 -25063
rect -9101 -25080 -9067 -25046
rect -9033 -25080 -8999 -25046
rect -8965 -25080 -8931 -25046
rect -8897 -25080 -8863 -25046
rect -8829 -25080 -8795 -25046
rect -8761 -25080 -8727 -25046
rect -8693 -25080 -8659 -25046
rect -8625 -25063 -8586 -25046
rect -8156 -25046 -7568 -25030
rect -8156 -25063 -8117 -25046
rect -8625 -25080 -8400 -25063
rect -9360 -25118 -8400 -25080
rect -8342 -25080 -8117 -25063
rect -8083 -25080 -8049 -25046
rect -8015 -25080 -7981 -25046
rect -7947 -25080 -7913 -25046
rect -7879 -25080 -7845 -25046
rect -7811 -25080 -7777 -25046
rect -7743 -25080 -7709 -25046
rect -7675 -25080 -7641 -25046
rect -7607 -25063 -7568 -25046
rect -7138 -25046 -6550 -25030
rect -7138 -25063 -7099 -25046
rect -7607 -25080 -7382 -25063
rect -8342 -25118 -7382 -25080
rect -7324 -25080 -7099 -25063
rect -7065 -25080 -7031 -25046
rect -6997 -25080 -6963 -25046
rect -6929 -25080 -6895 -25046
rect -6861 -25080 -6827 -25046
rect -6793 -25080 -6759 -25046
rect -6725 -25080 -6691 -25046
rect -6657 -25080 -6623 -25046
rect -6589 -25063 -6550 -25046
rect -6120 -25046 -5532 -25030
rect -6120 -25063 -6081 -25046
rect -6589 -25080 -6364 -25063
rect -7324 -25118 -6364 -25080
rect -6306 -25080 -6081 -25063
rect -6047 -25080 -6013 -25046
rect -5979 -25080 -5945 -25046
rect -5911 -25080 -5877 -25046
rect -5843 -25080 -5809 -25046
rect -5775 -25080 -5741 -25046
rect -5707 -25080 -5673 -25046
rect -5639 -25080 -5605 -25046
rect -5571 -25063 -5532 -25046
rect -5102 -25046 -4514 -25030
rect -5102 -25063 -5063 -25046
rect -5571 -25080 -5346 -25063
rect -6306 -25118 -5346 -25080
rect -5288 -25080 -5063 -25063
rect -5029 -25080 -4995 -25046
rect -4961 -25080 -4927 -25046
rect -4893 -25080 -4859 -25046
rect -4825 -25080 -4791 -25046
rect -4757 -25080 -4723 -25046
rect -4689 -25080 -4655 -25046
rect -4621 -25080 -4587 -25046
rect -4553 -25063 -4514 -25046
rect -4084 -25046 -3496 -25030
rect -4084 -25063 -4045 -25046
rect -4553 -25080 -4328 -25063
rect -5288 -25118 -4328 -25080
rect -4270 -25080 -4045 -25063
rect -4011 -25080 -3977 -25046
rect -3943 -25080 -3909 -25046
rect -3875 -25080 -3841 -25046
rect -3807 -25080 -3773 -25046
rect -3739 -25080 -3705 -25046
rect -3671 -25080 -3637 -25046
rect -3603 -25080 -3569 -25046
rect -3535 -25063 -3496 -25046
rect -2324 -25042 -2168 -25026
rect -2324 -25059 -2297 -25042
rect -3535 -25080 -3310 -25063
rect -4270 -25118 -3310 -25080
rect -2366 -25076 -2297 -25059
rect -2263 -25076 -2229 -25042
rect -2195 -25059 -2168 -25042
rect -2026 -25042 -1870 -25026
rect -2026 -25059 -1999 -25042
rect -2195 -25076 -2126 -25059
rect -2366 -25114 -2126 -25076
rect -2068 -25076 -1999 -25059
rect -1965 -25076 -1931 -25042
rect -1897 -25059 -1870 -25042
rect -1728 -25042 -1572 -25026
rect -1728 -25059 -1701 -25042
rect -1897 -25076 -1828 -25059
rect -2068 -25114 -1828 -25076
rect -1770 -25076 -1701 -25059
rect -1667 -25076 -1633 -25042
rect -1599 -25059 -1572 -25042
rect -1430 -25042 -1274 -25026
rect -1430 -25059 -1403 -25042
rect -1599 -25076 -1530 -25059
rect -1770 -25114 -1530 -25076
rect -1472 -25076 -1403 -25059
rect -1369 -25076 -1335 -25042
rect -1301 -25059 -1274 -25042
rect -1132 -25042 -976 -25026
rect -1132 -25059 -1105 -25042
rect -1301 -25076 -1232 -25059
rect -1472 -25114 -1232 -25076
rect -1174 -25076 -1105 -25059
rect -1071 -25076 -1037 -25042
rect -1003 -25059 -976 -25042
rect -834 -25042 -678 -25026
rect -834 -25059 -807 -25042
rect -1003 -25076 -934 -25059
rect -1174 -25114 -934 -25076
rect -876 -25076 -807 -25059
rect -773 -25076 -739 -25042
rect -705 -25059 -678 -25042
rect -536 -25042 -380 -25026
rect -536 -25059 -509 -25042
rect -705 -25076 -636 -25059
rect -876 -25114 -636 -25076
rect -578 -25076 -509 -25059
rect -475 -25076 -441 -25042
rect -407 -25059 -380 -25042
rect -238 -25042 -82 -25026
rect -238 -25059 -211 -25042
rect -407 -25076 -338 -25059
rect -578 -25114 -338 -25076
rect -280 -25076 -211 -25059
rect -177 -25076 -143 -25042
rect -109 -25059 -82 -25042
rect 60 -25042 216 -25026
rect 60 -25059 87 -25042
rect -109 -25076 -40 -25059
rect -280 -25114 -40 -25076
rect 18 -25076 87 -25059
rect 121 -25076 155 -25042
rect 189 -25059 216 -25042
rect 358 -25042 514 -25026
rect 358 -25059 385 -25042
rect 189 -25076 258 -25059
rect 18 -25114 258 -25076
rect 316 -25076 385 -25059
rect 419 -25076 453 -25042
rect 487 -25059 514 -25042
rect 656 -25042 812 -25026
rect 656 -25059 683 -25042
rect 487 -25076 556 -25059
rect 316 -25114 556 -25076
rect 614 -25076 683 -25059
rect 717 -25076 751 -25042
rect 785 -25059 812 -25042
rect 785 -25076 854 -25059
rect 614 -25114 854 -25076
rect 2812 -25212 3400 -25196
rect 2812 -25229 2851 -25212
rect 2626 -25246 2851 -25229
rect 2885 -25246 2919 -25212
rect 2953 -25246 2987 -25212
rect 3021 -25246 3055 -25212
rect 3089 -25246 3123 -25212
rect 3157 -25246 3191 -25212
rect 3225 -25246 3259 -25212
rect 3293 -25246 3327 -25212
rect 3361 -25229 3400 -25212
rect 3830 -25212 4418 -25196
rect 3830 -25229 3869 -25212
rect 3361 -25246 3586 -25229
rect 2626 -25284 3586 -25246
rect 3644 -25246 3869 -25229
rect 3903 -25246 3937 -25212
rect 3971 -25246 4005 -25212
rect 4039 -25246 4073 -25212
rect 4107 -25246 4141 -25212
rect 4175 -25246 4209 -25212
rect 4243 -25246 4277 -25212
rect 4311 -25246 4345 -25212
rect 4379 -25229 4418 -25212
rect 4848 -25212 5436 -25196
rect 4848 -25229 4887 -25212
rect 4379 -25246 4604 -25229
rect 3644 -25284 4604 -25246
rect 4662 -25246 4887 -25229
rect 4921 -25246 4955 -25212
rect 4989 -25246 5023 -25212
rect 5057 -25246 5091 -25212
rect 5125 -25246 5159 -25212
rect 5193 -25246 5227 -25212
rect 5261 -25246 5295 -25212
rect 5329 -25246 5363 -25212
rect 5397 -25229 5436 -25212
rect 5866 -25212 6454 -25196
rect 5866 -25229 5905 -25212
rect 5397 -25246 5622 -25229
rect 4662 -25284 5622 -25246
rect 5680 -25246 5905 -25229
rect 5939 -25246 5973 -25212
rect 6007 -25246 6041 -25212
rect 6075 -25246 6109 -25212
rect 6143 -25246 6177 -25212
rect 6211 -25246 6245 -25212
rect 6279 -25246 6313 -25212
rect 6347 -25246 6381 -25212
rect 6415 -25229 6454 -25212
rect 6884 -25212 7472 -25196
rect 6884 -25229 6923 -25212
rect 6415 -25246 6640 -25229
rect 5680 -25284 6640 -25246
rect 6698 -25246 6923 -25229
rect 6957 -25246 6991 -25212
rect 7025 -25246 7059 -25212
rect 7093 -25246 7127 -25212
rect 7161 -25246 7195 -25212
rect 7229 -25246 7263 -25212
rect 7297 -25246 7331 -25212
rect 7365 -25246 7399 -25212
rect 7433 -25229 7472 -25212
rect 7902 -25212 8490 -25196
rect 7902 -25229 7941 -25212
rect 7433 -25246 7658 -25229
rect 6698 -25284 7658 -25246
rect 7716 -25246 7941 -25229
rect 7975 -25246 8009 -25212
rect 8043 -25246 8077 -25212
rect 8111 -25246 8145 -25212
rect 8179 -25246 8213 -25212
rect 8247 -25246 8281 -25212
rect 8315 -25246 8349 -25212
rect 8383 -25246 8417 -25212
rect 8451 -25229 8490 -25212
rect 8920 -25212 9508 -25196
rect 8920 -25229 8959 -25212
rect 8451 -25246 8676 -25229
rect 7716 -25284 8676 -25246
rect 8734 -25246 8959 -25229
rect 8993 -25246 9027 -25212
rect 9061 -25246 9095 -25212
rect 9129 -25246 9163 -25212
rect 9197 -25246 9231 -25212
rect 9265 -25246 9299 -25212
rect 9333 -25246 9367 -25212
rect 9401 -25246 9435 -25212
rect 9469 -25229 9508 -25212
rect 9938 -25212 10526 -25196
rect 9938 -25229 9977 -25212
rect 9469 -25246 9694 -25229
rect 8734 -25284 9694 -25246
rect 9752 -25246 9977 -25229
rect 10011 -25246 10045 -25212
rect 10079 -25246 10113 -25212
rect 10147 -25246 10181 -25212
rect 10215 -25246 10249 -25212
rect 10283 -25246 10317 -25212
rect 10351 -25246 10385 -25212
rect 10419 -25246 10453 -25212
rect 10487 -25229 10526 -25212
rect 10956 -25212 11544 -25196
rect 10956 -25229 10995 -25212
rect 10487 -25246 10712 -25229
rect 9752 -25284 10712 -25246
rect 10770 -25246 10995 -25229
rect 11029 -25246 11063 -25212
rect 11097 -25246 11131 -25212
rect 11165 -25246 11199 -25212
rect 11233 -25246 11267 -25212
rect 11301 -25246 11335 -25212
rect 11369 -25246 11403 -25212
rect 11437 -25246 11471 -25212
rect 11505 -25229 11544 -25212
rect 11974 -25212 12562 -25196
rect 11974 -25229 12013 -25212
rect 11505 -25246 11730 -25229
rect 10770 -25284 11730 -25246
rect 11788 -25246 12013 -25229
rect 12047 -25246 12081 -25212
rect 12115 -25246 12149 -25212
rect 12183 -25246 12217 -25212
rect 12251 -25246 12285 -25212
rect 12319 -25246 12353 -25212
rect 12387 -25246 12421 -25212
rect 12455 -25246 12489 -25212
rect 12523 -25229 12562 -25212
rect 12992 -25212 13580 -25196
rect 12992 -25229 13031 -25212
rect 12523 -25246 12748 -25229
rect 11788 -25284 12748 -25246
rect 12806 -25246 13031 -25229
rect 13065 -25246 13099 -25212
rect 13133 -25246 13167 -25212
rect 13201 -25246 13235 -25212
rect 13269 -25246 13303 -25212
rect 13337 -25246 13371 -25212
rect 13405 -25246 13439 -25212
rect 13473 -25246 13507 -25212
rect 13541 -25229 13580 -25212
rect 14010 -25212 14598 -25196
rect 14010 -25229 14049 -25212
rect 13541 -25246 13766 -25229
rect 12806 -25284 13766 -25246
rect 13824 -25246 14049 -25229
rect 14083 -25246 14117 -25212
rect 14151 -25246 14185 -25212
rect 14219 -25246 14253 -25212
rect 14287 -25246 14321 -25212
rect 14355 -25246 14389 -25212
rect 14423 -25246 14457 -25212
rect 14491 -25246 14525 -25212
rect 14559 -25229 14598 -25212
rect 15028 -25212 15616 -25196
rect 15028 -25229 15067 -25212
rect 14559 -25246 14784 -25229
rect 13824 -25284 14784 -25246
rect 14842 -25246 15067 -25229
rect 15101 -25246 15135 -25212
rect 15169 -25246 15203 -25212
rect 15237 -25246 15271 -25212
rect 15305 -25246 15339 -25212
rect 15373 -25246 15407 -25212
rect 15441 -25246 15475 -25212
rect 15509 -25246 15543 -25212
rect 15577 -25229 15616 -25212
rect 16046 -25212 16634 -25196
rect 16046 -25229 16085 -25212
rect 15577 -25246 15802 -25229
rect 14842 -25284 15802 -25246
rect 15860 -25246 16085 -25229
rect 16119 -25246 16153 -25212
rect 16187 -25246 16221 -25212
rect 16255 -25246 16289 -25212
rect 16323 -25246 16357 -25212
rect 16391 -25246 16425 -25212
rect 16459 -25246 16493 -25212
rect 16527 -25246 16561 -25212
rect 16595 -25229 16634 -25212
rect 17064 -25212 17652 -25196
rect 17064 -25229 17103 -25212
rect 16595 -25246 16820 -25229
rect 15860 -25284 16820 -25246
rect 16878 -25246 17103 -25229
rect 17137 -25246 17171 -25212
rect 17205 -25246 17239 -25212
rect 17273 -25246 17307 -25212
rect 17341 -25246 17375 -25212
rect 17409 -25246 17443 -25212
rect 17477 -25246 17511 -25212
rect 17545 -25246 17579 -25212
rect 17613 -25229 17652 -25212
rect 18082 -25212 18670 -25196
rect 18082 -25229 18121 -25212
rect 17613 -25246 17838 -25229
rect 16878 -25284 17838 -25246
rect 17896 -25246 18121 -25229
rect 18155 -25246 18189 -25212
rect 18223 -25246 18257 -25212
rect 18291 -25246 18325 -25212
rect 18359 -25246 18393 -25212
rect 18427 -25246 18461 -25212
rect 18495 -25246 18529 -25212
rect 18563 -25246 18597 -25212
rect 18631 -25229 18670 -25212
rect 19100 -25212 19688 -25196
rect 19100 -25229 19139 -25212
rect 18631 -25246 18856 -25229
rect 17896 -25284 18856 -25246
rect 18914 -25246 19139 -25229
rect 19173 -25246 19207 -25212
rect 19241 -25246 19275 -25212
rect 19309 -25246 19343 -25212
rect 19377 -25246 19411 -25212
rect 19445 -25246 19479 -25212
rect 19513 -25246 19547 -25212
rect 19581 -25246 19615 -25212
rect 19649 -25229 19688 -25212
rect 20118 -25212 20706 -25196
rect 20118 -25229 20157 -25212
rect 19649 -25246 19874 -25229
rect 18914 -25284 19874 -25246
rect 19932 -25246 20157 -25229
rect 20191 -25246 20225 -25212
rect 20259 -25246 20293 -25212
rect 20327 -25246 20361 -25212
rect 20395 -25246 20429 -25212
rect 20463 -25246 20497 -25212
rect 20531 -25246 20565 -25212
rect 20599 -25246 20633 -25212
rect 20667 -25229 20706 -25212
rect 21136 -25212 21724 -25196
rect 21136 -25229 21175 -25212
rect 20667 -25246 20892 -25229
rect 19932 -25284 20892 -25246
rect 20950 -25246 21175 -25229
rect 21209 -25246 21243 -25212
rect 21277 -25246 21311 -25212
rect 21345 -25246 21379 -25212
rect 21413 -25246 21447 -25212
rect 21481 -25246 21515 -25212
rect 21549 -25246 21583 -25212
rect 21617 -25246 21651 -25212
rect 21685 -25229 21724 -25212
rect 22154 -25212 22742 -25196
rect 22154 -25229 22193 -25212
rect 21685 -25246 21910 -25229
rect 20950 -25284 21910 -25246
rect 21968 -25246 22193 -25229
rect 22227 -25246 22261 -25212
rect 22295 -25246 22329 -25212
rect 22363 -25246 22397 -25212
rect 22431 -25246 22465 -25212
rect 22499 -25246 22533 -25212
rect 22567 -25246 22601 -25212
rect 22635 -25246 22669 -25212
rect 22703 -25229 22742 -25212
rect 22703 -25246 22928 -25229
rect 21968 -25284 22928 -25246
rect -9360 -25756 -8400 -25718
rect -9360 -25773 -9135 -25756
rect -9174 -25790 -9135 -25773
rect -9101 -25790 -9067 -25756
rect -9033 -25790 -8999 -25756
rect -8965 -25790 -8931 -25756
rect -8897 -25790 -8863 -25756
rect -8829 -25790 -8795 -25756
rect -8761 -25790 -8727 -25756
rect -8693 -25790 -8659 -25756
rect -8625 -25773 -8400 -25756
rect -8342 -25756 -7382 -25718
rect -8342 -25773 -8117 -25756
rect -8625 -25790 -8586 -25773
rect -9174 -25806 -8586 -25790
rect -8156 -25790 -8117 -25773
rect -8083 -25790 -8049 -25756
rect -8015 -25790 -7981 -25756
rect -7947 -25790 -7913 -25756
rect -7879 -25790 -7845 -25756
rect -7811 -25790 -7777 -25756
rect -7743 -25790 -7709 -25756
rect -7675 -25790 -7641 -25756
rect -7607 -25773 -7382 -25756
rect -7324 -25756 -6364 -25718
rect -7324 -25773 -7099 -25756
rect -7607 -25790 -7568 -25773
rect -8156 -25806 -7568 -25790
rect -7138 -25790 -7099 -25773
rect -7065 -25790 -7031 -25756
rect -6997 -25790 -6963 -25756
rect -6929 -25790 -6895 -25756
rect -6861 -25790 -6827 -25756
rect -6793 -25790 -6759 -25756
rect -6725 -25790 -6691 -25756
rect -6657 -25790 -6623 -25756
rect -6589 -25773 -6364 -25756
rect -6306 -25756 -5346 -25718
rect -6306 -25773 -6081 -25756
rect -6589 -25790 -6550 -25773
rect -7138 -25806 -6550 -25790
rect -6120 -25790 -6081 -25773
rect -6047 -25790 -6013 -25756
rect -5979 -25790 -5945 -25756
rect -5911 -25790 -5877 -25756
rect -5843 -25790 -5809 -25756
rect -5775 -25790 -5741 -25756
rect -5707 -25790 -5673 -25756
rect -5639 -25790 -5605 -25756
rect -5571 -25773 -5346 -25756
rect -5288 -25756 -4328 -25718
rect -5288 -25773 -5063 -25756
rect -5571 -25790 -5532 -25773
rect -6120 -25806 -5532 -25790
rect -5102 -25790 -5063 -25773
rect -5029 -25790 -4995 -25756
rect -4961 -25790 -4927 -25756
rect -4893 -25790 -4859 -25756
rect -4825 -25790 -4791 -25756
rect -4757 -25790 -4723 -25756
rect -4689 -25790 -4655 -25756
rect -4621 -25790 -4587 -25756
rect -4553 -25773 -4328 -25756
rect -4270 -25756 -3310 -25718
rect -4270 -25773 -4045 -25756
rect -4553 -25790 -4514 -25773
rect -5102 -25806 -4514 -25790
rect -4084 -25790 -4045 -25773
rect -4011 -25790 -3977 -25756
rect -3943 -25790 -3909 -25756
rect -3875 -25790 -3841 -25756
rect -3807 -25790 -3773 -25756
rect -3739 -25790 -3705 -25756
rect -3671 -25790 -3637 -25756
rect -3603 -25790 -3569 -25756
rect -3535 -25773 -3310 -25756
rect -2366 -25752 -2126 -25714
rect -2366 -25769 -2297 -25752
rect -3535 -25790 -3496 -25773
rect -4084 -25806 -3496 -25790
rect -2324 -25786 -2297 -25769
rect -2263 -25786 -2229 -25752
rect -2195 -25769 -2126 -25752
rect -2068 -25752 -1828 -25714
rect -2068 -25769 -1999 -25752
rect -2195 -25786 -2168 -25769
rect -2324 -25802 -2168 -25786
rect -2026 -25786 -1999 -25769
rect -1965 -25786 -1931 -25752
rect -1897 -25769 -1828 -25752
rect -1770 -25752 -1530 -25714
rect -1770 -25769 -1701 -25752
rect -1897 -25786 -1870 -25769
rect -2026 -25802 -1870 -25786
rect -1728 -25786 -1701 -25769
rect -1667 -25786 -1633 -25752
rect -1599 -25769 -1530 -25752
rect -1472 -25752 -1232 -25714
rect -1472 -25769 -1403 -25752
rect -1599 -25786 -1572 -25769
rect -1728 -25802 -1572 -25786
rect -1430 -25786 -1403 -25769
rect -1369 -25786 -1335 -25752
rect -1301 -25769 -1232 -25752
rect -1174 -25752 -934 -25714
rect -1174 -25769 -1105 -25752
rect -1301 -25786 -1274 -25769
rect -1430 -25802 -1274 -25786
rect -1132 -25786 -1105 -25769
rect -1071 -25786 -1037 -25752
rect -1003 -25769 -934 -25752
rect -876 -25752 -636 -25714
rect -876 -25769 -807 -25752
rect -1003 -25786 -976 -25769
rect -1132 -25802 -976 -25786
rect -834 -25786 -807 -25769
rect -773 -25786 -739 -25752
rect -705 -25769 -636 -25752
rect -578 -25752 -338 -25714
rect -578 -25769 -509 -25752
rect -705 -25786 -678 -25769
rect -834 -25802 -678 -25786
rect -536 -25786 -509 -25769
rect -475 -25786 -441 -25752
rect -407 -25769 -338 -25752
rect -280 -25752 -40 -25714
rect -280 -25769 -211 -25752
rect -407 -25786 -380 -25769
rect -536 -25802 -380 -25786
rect -238 -25786 -211 -25769
rect -177 -25786 -143 -25752
rect -109 -25769 -40 -25752
rect 18 -25752 258 -25714
rect 18 -25769 87 -25752
rect -109 -25786 -82 -25769
rect -238 -25802 -82 -25786
rect 60 -25786 87 -25769
rect 121 -25786 155 -25752
rect 189 -25769 258 -25752
rect 316 -25752 556 -25714
rect 316 -25769 385 -25752
rect 189 -25786 216 -25769
rect 60 -25802 216 -25786
rect 358 -25786 385 -25769
rect 419 -25786 453 -25752
rect 487 -25769 556 -25752
rect 614 -25752 854 -25714
rect 614 -25769 683 -25752
rect 487 -25786 514 -25769
rect 358 -25802 514 -25786
rect 656 -25786 683 -25769
rect 717 -25786 751 -25752
rect 785 -25769 854 -25752
rect 785 -25786 812 -25769
rect 656 -25802 812 -25786
rect 2626 -25922 3586 -25884
rect 2626 -25939 2851 -25922
rect 2812 -25956 2851 -25939
rect 2885 -25956 2919 -25922
rect 2953 -25956 2987 -25922
rect 3021 -25956 3055 -25922
rect 3089 -25956 3123 -25922
rect 3157 -25956 3191 -25922
rect 3225 -25956 3259 -25922
rect 3293 -25956 3327 -25922
rect 3361 -25939 3586 -25922
rect 3644 -25922 4604 -25884
rect 3644 -25939 3869 -25922
rect 3361 -25956 3400 -25939
rect 2812 -25972 3400 -25956
rect 3830 -25956 3869 -25939
rect 3903 -25956 3937 -25922
rect 3971 -25956 4005 -25922
rect 4039 -25956 4073 -25922
rect 4107 -25956 4141 -25922
rect 4175 -25956 4209 -25922
rect 4243 -25956 4277 -25922
rect 4311 -25956 4345 -25922
rect 4379 -25939 4604 -25922
rect 4662 -25922 5622 -25884
rect 4662 -25939 4887 -25922
rect 4379 -25956 4418 -25939
rect 3830 -25972 4418 -25956
rect 4848 -25956 4887 -25939
rect 4921 -25956 4955 -25922
rect 4989 -25956 5023 -25922
rect 5057 -25956 5091 -25922
rect 5125 -25956 5159 -25922
rect 5193 -25956 5227 -25922
rect 5261 -25956 5295 -25922
rect 5329 -25956 5363 -25922
rect 5397 -25939 5622 -25922
rect 5680 -25922 6640 -25884
rect 5680 -25939 5905 -25922
rect 5397 -25956 5436 -25939
rect 4848 -25972 5436 -25956
rect 5866 -25956 5905 -25939
rect 5939 -25956 5973 -25922
rect 6007 -25956 6041 -25922
rect 6075 -25956 6109 -25922
rect 6143 -25956 6177 -25922
rect 6211 -25956 6245 -25922
rect 6279 -25956 6313 -25922
rect 6347 -25956 6381 -25922
rect 6415 -25939 6640 -25922
rect 6698 -25922 7658 -25884
rect 6698 -25939 6923 -25922
rect 6415 -25956 6454 -25939
rect 5866 -25972 6454 -25956
rect 6884 -25956 6923 -25939
rect 6957 -25956 6991 -25922
rect 7025 -25956 7059 -25922
rect 7093 -25956 7127 -25922
rect 7161 -25956 7195 -25922
rect 7229 -25956 7263 -25922
rect 7297 -25956 7331 -25922
rect 7365 -25956 7399 -25922
rect 7433 -25939 7658 -25922
rect 7716 -25922 8676 -25884
rect 7716 -25939 7941 -25922
rect 7433 -25956 7472 -25939
rect 6884 -25972 7472 -25956
rect 7902 -25956 7941 -25939
rect 7975 -25956 8009 -25922
rect 8043 -25956 8077 -25922
rect 8111 -25956 8145 -25922
rect 8179 -25956 8213 -25922
rect 8247 -25956 8281 -25922
rect 8315 -25956 8349 -25922
rect 8383 -25956 8417 -25922
rect 8451 -25939 8676 -25922
rect 8734 -25922 9694 -25884
rect 8734 -25939 8959 -25922
rect 8451 -25956 8490 -25939
rect 7902 -25972 8490 -25956
rect 8920 -25956 8959 -25939
rect 8993 -25956 9027 -25922
rect 9061 -25956 9095 -25922
rect 9129 -25956 9163 -25922
rect 9197 -25956 9231 -25922
rect 9265 -25956 9299 -25922
rect 9333 -25956 9367 -25922
rect 9401 -25956 9435 -25922
rect 9469 -25939 9694 -25922
rect 9752 -25922 10712 -25884
rect 9752 -25939 9977 -25922
rect 9469 -25956 9508 -25939
rect 8920 -25972 9508 -25956
rect 9938 -25956 9977 -25939
rect 10011 -25956 10045 -25922
rect 10079 -25956 10113 -25922
rect 10147 -25956 10181 -25922
rect 10215 -25956 10249 -25922
rect 10283 -25956 10317 -25922
rect 10351 -25956 10385 -25922
rect 10419 -25956 10453 -25922
rect 10487 -25939 10712 -25922
rect 10770 -25922 11730 -25884
rect 10770 -25939 10995 -25922
rect 10487 -25956 10526 -25939
rect 9938 -25972 10526 -25956
rect 10956 -25956 10995 -25939
rect 11029 -25956 11063 -25922
rect 11097 -25956 11131 -25922
rect 11165 -25956 11199 -25922
rect 11233 -25956 11267 -25922
rect 11301 -25956 11335 -25922
rect 11369 -25956 11403 -25922
rect 11437 -25956 11471 -25922
rect 11505 -25939 11730 -25922
rect 11788 -25922 12748 -25884
rect 11788 -25939 12013 -25922
rect 11505 -25956 11544 -25939
rect 10956 -25972 11544 -25956
rect 11974 -25956 12013 -25939
rect 12047 -25956 12081 -25922
rect 12115 -25956 12149 -25922
rect 12183 -25956 12217 -25922
rect 12251 -25956 12285 -25922
rect 12319 -25956 12353 -25922
rect 12387 -25956 12421 -25922
rect 12455 -25956 12489 -25922
rect 12523 -25939 12748 -25922
rect 12806 -25922 13766 -25884
rect 12806 -25939 13031 -25922
rect 12523 -25956 12562 -25939
rect 11974 -25972 12562 -25956
rect 12992 -25956 13031 -25939
rect 13065 -25956 13099 -25922
rect 13133 -25956 13167 -25922
rect 13201 -25956 13235 -25922
rect 13269 -25956 13303 -25922
rect 13337 -25956 13371 -25922
rect 13405 -25956 13439 -25922
rect 13473 -25956 13507 -25922
rect 13541 -25939 13766 -25922
rect 13824 -25922 14784 -25884
rect 13824 -25939 14049 -25922
rect 13541 -25956 13580 -25939
rect 12992 -25972 13580 -25956
rect 14010 -25956 14049 -25939
rect 14083 -25956 14117 -25922
rect 14151 -25956 14185 -25922
rect 14219 -25956 14253 -25922
rect 14287 -25956 14321 -25922
rect 14355 -25956 14389 -25922
rect 14423 -25956 14457 -25922
rect 14491 -25956 14525 -25922
rect 14559 -25939 14784 -25922
rect 14842 -25922 15802 -25884
rect 14842 -25939 15067 -25922
rect 14559 -25956 14598 -25939
rect 14010 -25972 14598 -25956
rect 15028 -25956 15067 -25939
rect 15101 -25956 15135 -25922
rect 15169 -25956 15203 -25922
rect 15237 -25956 15271 -25922
rect 15305 -25956 15339 -25922
rect 15373 -25956 15407 -25922
rect 15441 -25956 15475 -25922
rect 15509 -25956 15543 -25922
rect 15577 -25939 15802 -25922
rect 15860 -25922 16820 -25884
rect 15860 -25939 16085 -25922
rect 15577 -25956 15616 -25939
rect 15028 -25972 15616 -25956
rect 16046 -25956 16085 -25939
rect 16119 -25956 16153 -25922
rect 16187 -25956 16221 -25922
rect 16255 -25956 16289 -25922
rect 16323 -25956 16357 -25922
rect 16391 -25956 16425 -25922
rect 16459 -25956 16493 -25922
rect 16527 -25956 16561 -25922
rect 16595 -25939 16820 -25922
rect 16878 -25922 17838 -25884
rect 16878 -25939 17103 -25922
rect 16595 -25956 16634 -25939
rect 16046 -25972 16634 -25956
rect 17064 -25956 17103 -25939
rect 17137 -25956 17171 -25922
rect 17205 -25956 17239 -25922
rect 17273 -25956 17307 -25922
rect 17341 -25956 17375 -25922
rect 17409 -25956 17443 -25922
rect 17477 -25956 17511 -25922
rect 17545 -25956 17579 -25922
rect 17613 -25939 17838 -25922
rect 17896 -25922 18856 -25884
rect 17896 -25939 18121 -25922
rect 17613 -25956 17652 -25939
rect 17064 -25972 17652 -25956
rect 18082 -25956 18121 -25939
rect 18155 -25956 18189 -25922
rect 18223 -25956 18257 -25922
rect 18291 -25956 18325 -25922
rect 18359 -25956 18393 -25922
rect 18427 -25956 18461 -25922
rect 18495 -25956 18529 -25922
rect 18563 -25956 18597 -25922
rect 18631 -25939 18856 -25922
rect 18914 -25922 19874 -25884
rect 18914 -25939 19139 -25922
rect 18631 -25956 18670 -25939
rect 18082 -25972 18670 -25956
rect 19100 -25956 19139 -25939
rect 19173 -25956 19207 -25922
rect 19241 -25956 19275 -25922
rect 19309 -25956 19343 -25922
rect 19377 -25956 19411 -25922
rect 19445 -25956 19479 -25922
rect 19513 -25956 19547 -25922
rect 19581 -25956 19615 -25922
rect 19649 -25939 19874 -25922
rect 19932 -25922 20892 -25884
rect 19932 -25939 20157 -25922
rect 19649 -25956 19688 -25939
rect 19100 -25972 19688 -25956
rect 20118 -25956 20157 -25939
rect 20191 -25956 20225 -25922
rect 20259 -25956 20293 -25922
rect 20327 -25956 20361 -25922
rect 20395 -25956 20429 -25922
rect 20463 -25956 20497 -25922
rect 20531 -25956 20565 -25922
rect 20599 -25956 20633 -25922
rect 20667 -25939 20892 -25922
rect 20950 -25922 21910 -25884
rect 20950 -25939 21175 -25922
rect 20667 -25956 20706 -25939
rect 20118 -25972 20706 -25956
rect 21136 -25956 21175 -25939
rect 21209 -25956 21243 -25922
rect 21277 -25956 21311 -25922
rect 21345 -25956 21379 -25922
rect 21413 -25956 21447 -25922
rect 21481 -25956 21515 -25922
rect 21549 -25956 21583 -25922
rect 21617 -25956 21651 -25922
rect 21685 -25939 21910 -25922
rect 21968 -25922 22928 -25884
rect 21968 -25939 22193 -25922
rect 21685 -25956 21724 -25939
rect 21136 -25972 21724 -25956
rect 22154 -25956 22193 -25939
rect 22227 -25956 22261 -25922
rect 22295 -25956 22329 -25922
rect 22363 -25956 22397 -25922
rect 22431 -25956 22465 -25922
rect 22499 -25956 22533 -25922
rect 22567 -25956 22601 -25922
rect 22635 -25956 22669 -25922
rect 22703 -25939 22928 -25922
rect 22703 -25956 22742 -25939
rect 22154 -25972 22742 -25956
<< polycont >>
rect 3735 -4643 3769 -4609
rect 3953 -4643 3987 -4609
rect 4171 -4643 4205 -4609
rect 4389 -4643 4423 -4609
rect 4607 -4643 4641 -4609
rect 4825 -4643 4859 -4609
rect 5043 -4643 5077 -4609
rect 5261 -4643 5295 -4609
rect 5479 -4643 5513 -4609
rect 5697 -4643 5731 -4609
rect 3735 -5171 3769 -5137
rect 3953 -5171 3987 -5137
rect 4171 -5171 4205 -5137
rect 4389 -5171 4423 -5137
rect 4607 -5171 4641 -5137
rect 4825 -5171 4859 -5137
rect 5043 -5171 5077 -5137
rect 5261 -5171 5295 -5137
rect 5479 -5171 5513 -5137
rect 5697 -5171 5731 -5137
rect 3735 -5581 3769 -5547
rect 3953 -5581 3987 -5547
rect 4171 -5581 4205 -5547
rect 4389 -5581 4423 -5547
rect 4607 -5581 4641 -5547
rect 4825 -5581 4859 -5547
rect 5043 -5581 5077 -5547
rect 5261 -5581 5295 -5547
rect 5479 -5581 5513 -5547
rect 5697 -5581 5731 -5547
rect 3735 -6109 3769 -6075
rect 3953 -6109 3987 -6075
rect 4171 -6109 4205 -6075
rect 4389 -6109 4423 -6075
rect 4607 -6109 4641 -6075
rect 4825 -6109 4859 -6075
rect 5043 -6109 5077 -6075
rect 5261 -6109 5295 -6075
rect 5479 -6109 5513 -6075
rect 5697 -6109 5731 -6075
rect 3735 -6519 3769 -6485
rect 3953 -6519 3987 -6485
rect 4171 -6519 4205 -6485
rect 4389 -6519 4423 -6485
rect 4607 -6519 4641 -6485
rect 4825 -6519 4859 -6485
rect 5043 -6519 5077 -6485
rect 5261 -6519 5295 -6485
rect 5479 -6519 5513 -6485
rect 5697 -6519 5731 -6485
rect 3735 -7047 3769 -7013
rect 3953 -7047 3987 -7013
rect 4171 -7047 4205 -7013
rect 4389 -7047 4423 -7013
rect 4607 -7047 4641 -7013
rect 4825 -7047 4859 -7013
rect 5043 -7047 5077 -7013
rect 5261 -7047 5295 -7013
rect 5479 -7047 5513 -7013
rect 5697 -7047 5731 -7013
rect 3735 -7457 3769 -7423
rect 3953 -7457 3987 -7423
rect 4171 -7457 4205 -7423
rect 4389 -7457 4423 -7423
rect 4607 -7457 4641 -7423
rect 4825 -7457 4859 -7423
rect 5043 -7457 5077 -7423
rect 5261 -7457 5295 -7423
rect 5479 -7457 5513 -7423
rect 5697 -7457 5731 -7423
rect 3735 -7985 3769 -7951
rect 3953 -7985 3987 -7951
rect 4171 -7985 4205 -7951
rect 4389 -7985 4423 -7951
rect 4607 -7985 4641 -7951
rect 4825 -7985 4859 -7951
rect 5043 -7985 5077 -7951
rect 5261 -7985 5295 -7951
rect 5479 -7985 5513 -7951
rect 5697 -7985 5731 -7951
rect 2853 -11680 2887 -11646
rect 2921 -11680 2955 -11646
rect 2989 -11680 3023 -11646
rect 3057 -11680 3091 -11646
rect 3125 -11680 3159 -11646
rect 3193 -11680 3227 -11646
rect 3261 -11680 3295 -11646
rect 3329 -11680 3363 -11646
rect 3871 -11680 3905 -11646
rect 3939 -11680 3973 -11646
rect 4007 -11680 4041 -11646
rect 4075 -11680 4109 -11646
rect 4143 -11680 4177 -11646
rect 4211 -11680 4245 -11646
rect 4279 -11680 4313 -11646
rect 4347 -11680 4381 -11646
rect 4889 -11680 4923 -11646
rect 4957 -11680 4991 -11646
rect 5025 -11680 5059 -11646
rect 5093 -11680 5127 -11646
rect 5161 -11680 5195 -11646
rect 5229 -11680 5263 -11646
rect 5297 -11680 5331 -11646
rect 5365 -11680 5399 -11646
rect 5907 -11680 5941 -11646
rect 5975 -11680 6009 -11646
rect 6043 -11680 6077 -11646
rect 6111 -11680 6145 -11646
rect 6179 -11680 6213 -11646
rect 6247 -11680 6281 -11646
rect 6315 -11680 6349 -11646
rect 6383 -11680 6417 -11646
rect 6925 -11680 6959 -11646
rect 6993 -11680 7027 -11646
rect 7061 -11680 7095 -11646
rect 7129 -11680 7163 -11646
rect 7197 -11680 7231 -11646
rect 7265 -11680 7299 -11646
rect 7333 -11680 7367 -11646
rect 7401 -11680 7435 -11646
rect 7943 -11680 7977 -11646
rect 8011 -11680 8045 -11646
rect 8079 -11680 8113 -11646
rect 8147 -11680 8181 -11646
rect 8215 -11680 8249 -11646
rect 8283 -11680 8317 -11646
rect 8351 -11680 8385 -11646
rect 8419 -11680 8453 -11646
rect 8961 -11680 8995 -11646
rect 9029 -11680 9063 -11646
rect 9097 -11680 9131 -11646
rect 9165 -11680 9199 -11646
rect 9233 -11680 9267 -11646
rect 9301 -11680 9335 -11646
rect 9369 -11680 9403 -11646
rect 9437 -11680 9471 -11646
rect 9979 -11680 10013 -11646
rect 10047 -11680 10081 -11646
rect 10115 -11680 10149 -11646
rect 10183 -11680 10217 -11646
rect 10251 -11680 10285 -11646
rect 10319 -11680 10353 -11646
rect 10387 -11680 10421 -11646
rect 10455 -11680 10489 -11646
rect 10997 -11680 11031 -11646
rect 11065 -11680 11099 -11646
rect 11133 -11680 11167 -11646
rect 11201 -11680 11235 -11646
rect 11269 -11680 11303 -11646
rect 11337 -11680 11371 -11646
rect 11405 -11680 11439 -11646
rect 11473 -11680 11507 -11646
rect 12015 -11680 12049 -11646
rect 12083 -11680 12117 -11646
rect 12151 -11680 12185 -11646
rect 12219 -11680 12253 -11646
rect 12287 -11680 12321 -11646
rect 12355 -11680 12389 -11646
rect 12423 -11680 12457 -11646
rect 12491 -11680 12525 -11646
rect 13033 -11680 13067 -11646
rect 13101 -11680 13135 -11646
rect 13169 -11680 13203 -11646
rect 13237 -11680 13271 -11646
rect 13305 -11680 13339 -11646
rect 13373 -11680 13407 -11646
rect 13441 -11680 13475 -11646
rect 13509 -11680 13543 -11646
rect 14051 -11680 14085 -11646
rect 14119 -11680 14153 -11646
rect 14187 -11680 14221 -11646
rect 14255 -11680 14289 -11646
rect 14323 -11680 14357 -11646
rect 14391 -11680 14425 -11646
rect 14459 -11680 14493 -11646
rect 14527 -11680 14561 -11646
rect 15069 -11680 15103 -11646
rect 15137 -11680 15171 -11646
rect 15205 -11680 15239 -11646
rect 15273 -11680 15307 -11646
rect 15341 -11680 15375 -11646
rect 15409 -11680 15443 -11646
rect 15477 -11680 15511 -11646
rect 15545 -11680 15579 -11646
rect 16087 -11680 16121 -11646
rect 16155 -11680 16189 -11646
rect 16223 -11680 16257 -11646
rect 16291 -11680 16325 -11646
rect 16359 -11680 16393 -11646
rect 16427 -11680 16461 -11646
rect 16495 -11680 16529 -11646
rect 16563 -11680 16597 -11646
rect 17105 -11680 17139 -11646
rect 17173 -11680 17207 -11646
rect 17241 -11680 17275 -11646
rect 17309 -11680 17343 -11646
rect 17377 -11680 17411 -11646
rect 17445 -11680 17479 -11646
rect 17513 -11680 17547 -11646
rect 17581 -11680 17615 -11646
rect 18123 -11680 18157 -11646
rect 18191 -11680 18225 -11646
rect 18259 -11680 18293 -11646
rect 18327 -11680 18361 -11646
rect 18395 -11680 18429 -11646
rect 18463 -11680 18497 -11646
rect 18531 -11680 18565 -11646
rect 18599 -11680 18633 -11646
rect 19141 -11680 19175 -11646
rect 19209 -11680 19243 -11646
rect 19277 -11680 19311 -11646
rect 19345 -11680 19379 -11646
rect 19413 -11680 19447 -11646
rect 19481 -11680 19515 -11646
rect 19549 -11680 19583 -11646
rect 19617 -11680 19651 -11646
rect 20159 -11680 20193 -11646
rect 20227 -11680 20261 -11646
rect 20295 -11680 20329 -11646
rect 20363 -11680 20397 -11646
rect 20431 -11680 20465 -11646
rect 20499 -11680 20533 -11646
rect 20567 -11680 20601 -11646
rect 20635 -11680 20669 -11646
rect 21177 -11680 21211 -11646
rect 21245 -11680 21279 -11646
rect 21313 -11680 21347 -11646
rect 21381 -11680 21415 -11646
rect 21449 -11680 21483 -11646
rect 21517 -11680 21551 -11646
rect 21585 -11680 21619 -11646
rect 21653 -11680 21687 -11646
rect 22195 -11680 22229 -11646
rect 22263 -11680 22297 -11646
rect 22331 -11680 22365 -11646
rect 22399 -11680 22433 -11646
rect 22467 -11680 22501 -11646
rect 22535 -11680 22569 -11646
rect 22603 -11680 22637 -11646
rect 22671 -11680 22705 -11646
rect 2853 -12390 2887 -12356
rect 2921 -12390 2955 -12356
rect 2989 -12390 3023 -12356
rect 3057 -12390 3091 -12356
rect 3125 -12390 3159 -12356
rect 3193 -12390 3227 -12356
rect 3261 -12390 3295 -12356
rect 3329 -12390 3363 -12356
rect 3871 -12390 3905 -12356
rect 3939 -12390 3973 -12356
rect 4007 -12390 4041 -12356
rect 4075 -12390 4109 -12356
rect 4143 -12390 4177 -12356
rect 4211 -12390 4245 -12356
rect 4279 -12390 4313 -12356
rect 4347 -12390 4381 -12356
rect 4889 -12390 4923 -12356
rect 4957 -12390 4991 -12356
rect 5025 -12390 5059 -12356
rect 5093 -12390 5127 -12356
rect 5161 -12390 5195 -12356
rect 5229 -12390 5263 -12356
rect 5297 -12390 5331 -12356
rect 5365 -12390 5399 -12356
rect 5907 -12390 5941 -12356
rect 5975 -12390 6009 -12356
rect 6043 -12390 6077 -12356
rect 6111 -12390 6145 -12356
rect 6179 -12390 6213 -12356
rect 6247 -12390 6281 -12356
rect 6315 -12390 6349 -12356
rect 6383 -12390 6417 -12356
rect 6925 -12390 6959 -12356
rect 6993 -12390 7027 -12356
rect 7061 -12390 7095 -12356
rect 7129 -12390 7163 -12356
rect 7197 -12390 7231 -12356
rect 7265 -12390 7299 -12356
rect 7333 -12390 7367 -12356
rect 7401 -12390 7435 -12356
rect 7943 -12390 7977 -12356
rect 8011 -12390 8045 -12356
rect 8079 -12390 8113 -12356
rect 8147 -12390 8181 -12356
rect 8215 -12390 8249 -12356
rect 8283 -12390 8317 -12356
rect 8351 -12390 8385 -12356
rect 8419 -12390 8453 -12356
rect 8961 -12390 8995 -12356
rect 9029 -12390 9063 -12356
rect 9097 -12390 9131 -12356
rect 9165 -12390 9199 -12356
rect 9233 -12390 9267 -12356
rect 9301 -12390 9335 -12356
rect 9369 -12390 9403 -12356
rect 9437 -12390 9471 -12356
rect 9979 -12390 10013 -12356
rect 10047 -12390 10081 -12356
rect 10115 -12390 10149 -12356
rect 10183 -12390 10217 -12356
rect 10251 -12390 10285 -12356
rect 10319 -12390 10353 -12356
rect 10387 -12390 10421 -12356
rect 10455 -12390 10489 -12356
rect 10997 -12390 11031 -12356
rect 11065 -12390 11099 -12356
rect 11133 -12390 11167 -12356
rect 11201 -12390 11235 -12356
rect 11269 -12390 11303 -12356
rect 11337 -12390 11371 -12356
rect 11405 -12390 11439 -12356
rect 11473 -12390 11507 -12356
rect 12015 -12390 12049 -12356
rect 12083 -12390 12117 -12356
rect 12151 -12390 12185 -12356
rect 12219 -12390 12253 -12356
rect 12287 -12390 12321 -12356
rect 12355 -12390 12389 -12356
rect 12423 -12390 12457 -12356
rect 12491 -12390 12525 -12356
rect 13033 -12390 13067 -12356
rect 13101 -12390 13135 -12356
rect 13169 -12390 13203 -12356
rect 13237 -12390 13271 -12356
rect 13305 -12390 13339 -12356
rect 13373 -12390 13407 -12356
rect 13441 -12390 13475 -12356
rect 13509 -12390 13543 -12356
rect 14051 -12390 14085 -12356
rect 14119 -12390 14153 -12356
rect 14187 -12390 14221 -12356
rect 14255 -12390 14289 -12356
rect 14323 -12390 14357 -12356
rect 14391 -12390 14425 -12356
rect 14459 -12390 14493 -12356
rect 14527 -12390 14561 -12356
rect 15069 -12390 15103 -12356
rect 15137 -12390 15171 -12356
rect 15205 -12390 15239 -12356
rect 15273 -12390 15307 -12356
rect 15341 -12390 15375 -12356
rect 15409 -12390 15443 -12356
rect 15477 -12390 15511 -12356
rect 15545 -12390 15579 -12356
rect 16087 -12390 16121 -12356
rect 16155 -12390 16189 -12356
rect 16223 -12390 16257 -12356
rect 16291 -12390 16325 -12356
rect 16359 -12390 16393 -12356
rect 16427 -12390 16461 -12356
rect 16495 -12390 16529 -12356
rect 16563 -12390 16597 -12356
rect 17105 -12390 17139 -12356
rect 17173 -12390 17207 -12356
rect 17241 -12390 17275 -12356
rect 17309 -12390 17343 -12356
rect 17377 -12390 17411 -12356
rect 17445 -12390 17479 -12356
rect 17513 -12390 17547 -12356
rect 17581 -12390 17615 -12356
rect 18123 -12390 18157 -12356
rect 18191 -12390 18225 -12356
rect 18259 -12390 18293 -12356
rect 18327 -12390 18361 -12356
rect 18395 -12390 18429 -12356
rect 18463 -12390 18497 -12356
rect 18531 -12390 18565 -12356
rect 18599 -12390 18633 -12356
rect 19141 -12390 19175 -12356
rect 19209 -12390 19243 -12356
rect 19277 -12390 19311 -12356
rect 19345 -12390 19379 -12356
rect 19413 -12390 19447 -12356
rect 19481 -12390 19515 -12356
rect 19549 -12390 19583 -12356
rect 19617 -12390 19651 -12356
rect 20159 -12390 20193 -12356
rect 20227 -12390 20261 -12356
rect 20295 -12390 20329 -12356
rect 20363 -12390 20397 -12356
rect 20431 -12390 20465 -12356
rect 20499 -12390 20533 -12356
rect 20567 -12390 20601 -12356
rect 20635 -12390 20669 -12356
rect 21177 -12390 21211 -12356
rect 21245 -12390 21279 -12356
rect 21313 -12390 21347 -12356
rect 21381 -12390 21415 -12356
rect 21449 -12390 21483 -12356
rect 21517 -12390 21551 -12356
rect 21585 -12390 21619 -12356
rect 21653 -12390 21687 -12356
rect 22195 -12390 22229 -12356
rect 22263 -12390 22297 -12356
rect 22331 -12390 22365 -12356
rect 22399 -12390 22433 -12356
rect 22467 -12390 22501 -12356
rect 22535 -12390 22569 -12356
rect 22603 -12390 22637 -12356
rect 22671 -12390 22705 -12356
rect -8913 -12474 -8879 -12440
rect -8845 -12474 -8811 -12440
rect -8777 -12474 -8743 -12440
rect -8709 -12474 -8675 -12440
rect -8641 -12474 -8607 -12440
rect -8573 -12474 -8539 -12440
rect -8505 -12474 -8471 -12440
rect -8437 -12474 -8403 -12440
rect -7895 -12474 -7861 -12440
rect -7827 -12474 -7793 -12440
rect -7759 -12474 -7725 -12440
rect -7691 -12474 -7657 -12440
rect -7623 -12474 -7589 -12440
rect -7555 -12474 -7521 -12440
rect -7487 -12474 -7453 -12440
rect -7419 -12474 -7385 -12440
rect -6877 -12474 -6843 -12440
rect -6809 -12474 -6775 -12440
rect -6741 -12474 -6707 -12440
rect -6673 -12474 -6639 -12440
rect -6605 -12474 -6571 -12440
rect -6537 -12474 -6503 -12440
rect -6469 -12474 -6435 -12440
rect -6401 -12474 -6367 -12440
rect -5859 -12474 -5825 -12440
rect -5791 -12474 -5757 -12440
rect -5723 -12474 -5689 -12440
rect -5655 -12474 -5621 -12440
rect -5587 -12474 -5553 -12440
rect -5519 -12474 -5485 -12440
rect -5451 -12474 -5417 -12440
rect -5383 -12474 -5349 -12440
rect -4841 -12474 -4807 -12440
rect -4773 -12474 -4739 -12440
rect -4705 -12474 -4671 -12440
rect -4637 -12474 -4603 -12440
rect -4569 -12474 -4535 -12440
rect -4501 -12474 -4467 -12440
rect -4433 -12474 -4399 -12440
rect -4365 -12474 -4331 -12440
rect -3823 -12474 -3789 -12440
rect -3755 -12474 -3721 -12440
rect -3687 -12474 -3653 -12440
rect -3619 -12474 -3585 -12440
rect -3551 -12474 -3517 -12440
rect -3483 -12474 -3449 -12440
rect -3415 -12474 -3381 -12440
rect -3347 -12474 -3313 -12440
rect -2805 -12474 -2771 -12440
rect -2737 -12474 -2703 -12440
rect -2669 -12474 -2635 -12440
rect -2601 -12474 -2567 -12440
rect -2533 -12474 -2499 -12440
rect -2465 -12474 -2431 -12440
rect -2397 -12474 -2363 -12440
rect -2329 -12474 -2295 -12440
rect -1787 -12474 -1753 -12440
rect -1719 -12474 -1685 -12440
rect -1651 -12474 -1617 -12440
rect -1583 -12474 -1549 -12440
rect -1515 -12474 -1481 -12440
rect -1447 -12474 -1413 -12440
rect -1379 -12474 -1345 -12440
rect -1311 -12474 -1277 -12440
rect -769 -12474 -735 -12440
rect -701 -12474 -667 -12440
rect -633 -12474 -599 -12440
rect -565 -12474 -531 -12440
rect -497 -12474 -463 -12440
rect -429 -12474 -395 -12440
rect -361 -12474 -327 -12440
rect -293 -12474 -259 -12440
rect 2853 -12914 2887 -12880
rect 2921 -12914 2955 -12880
rect 2989 -12914 3023 -12880
rect 3057 -12914 3091 -12880
rect 3125 -12914 3159 -12880
rect 3193 -12914 3227 -12880
rect 3261 -12914 3295 -12880
rect 3329 -12914 3363 -12880
rect 3871 -12914 3905 -12880
rect 3939 -12914 3973 -12880
rect 4007 -12914 4041 -12880
rect 4075 -12914 4109 -12880
rect 4143 -12914 4177 -12880
rect 4211 -12914 4245 -12880
rect 4279 -12914 4313 -12880
rect 4347 -12914 4381 -12880
rect 4889 -12914 4923 -12880
rect 4957 -12914 4991 -12880
rect 5025 -12914 5059 -12880
rect 5093 -12914 5127 -12880
rect 5161 -12914 5195 -12880
rect 5229 -12914 5263 -12880
rect 5297 -12914 5331 -12880
rect 5365 -12914 5399 -12880
rect 5907 -12914 5941 -12880
rect 5975 -12914 6009 -12880
rect 6043 -12914 6077 -12880
rect 6111 -12914 6145 -12880
rect 6179 -12914 6213 -12880
rect 6247 -12914 6281 -12880
rect 6315 -12914 6349 -12880
rect 6383 -12914 6417 -12880
rect 6925 -12914 6959 -12880
rect 6993 -12914 7027 -12880
rect 7061 -12914 7095 -12880
rect 7129 -12914 7163 -12880
rect 7197 -12914 7231 -12880
rect 7265 -12914 7299 -12880
rect 7333 -12914 7367 -12880
rect 7401 -12914 7435 -12880
rect 7943 -12914 7977 -12880
rect 8011 -12914 8045 -12880
rect 8079 -12914 8113 -12880
rect 8147 -12914 8181 -12880
rect 8215 -12914 8249 -12880
rect 8283 -12914 8317 -12880
rect 8351 -12914 8385 -12880
rect 8419 -12914 8453 -12880
rect 8961 -12914 8995 -12880
rect 9029 -12914 9063 -12880
rect 9097 -12914 9131 -12880
rect 9165 -12914 9199 -12880
rect 9233 -12914 9267 -12880
rect 9301 -12914 9335 -12880
rect 9369 -12914 9403 -12880
rect 9437 -12914 9471 -12880
rect 9979 -12914 10013 -12880
rect 10047 -12914 10081 -12880
rect 10115 -12914 10149 -12880
rect 10183 -12914 10217 -12880
rect 10251 -12914 10285 -12880
rect 10319 -12914 10353 -12880
rect 10387 -12914 10421 -12880
rect 10455 -12914 10489 -12880
rect 10997 -12914 11031 -12880
rect 11065 -12914 11099 -12880
rect 11133 -12914 11167 -12880
rect 11201 -12914 11235 -12880
rect 11269 -12914 11303 -12880
rect 11337 -12914 11371 -12880
rect 11405 -12914 11439 -12880
rect 11473 -12914 11507 -12880
rect 12015 -12914 12049 -12880
rect 12083 -12914 12117 -12880
rect 12151 -12914 12185 -12880
rect 12219 -12914 12253 -12880
rect 12287 -12914 12321 -12880
rect 12355 -12914 12389 -12880
rect 12423 -12914 12457 -12880
rect 12491 -12914 12525 -12880
rect 13033 -12914 13067 -12880
rect 13101 -12914 13135 -12880
rect 13169 -12914 13203 -12880
rect 13237 -12914 13271 -12880
rect 13305 -12914 13339 -12880
rect 13373 -12914 13407 -12880
rect 13441 -12914 13475 -12880
rect 13509 -12914 13543 -12880
rect 14051 -12914 14085 -12880
rect 14119 -12914 14153 -12880
rect 14187 -12914 14221 -12880
rect 14255 -12914 14289 -12880
rect 14323 -12914 14357 -12880
rect 14391 -12914 14425 -12880
rect 14459 -12914 14493 -12880
rect 14527 -12914 14561 -12880
rect 15069 -12914 15103 -12880
rect 15137 -12914 15171 -12880
rect 15205 -12914 15239 -12880
rect 15273 -12914 15307 -12880
rect 15341 -12914 15375 -12880
rect 15409 -12914 15443 -12880
rect 15477 -12914 15511 -12880
rect 15545 -12914 15579 -12880
rect 16087 -12914 16121 -12880
rect 16155 -12914 16189 -12880
rect 16223 -12914 16257 -12880
rect 16291 -12914 16325 -12880
rect 16359 -12914 16393 -12880
rect 16427 -12914 16461 -12880
rect 16495 -12914 16529 -12880
rect 16563 -12914 16597 -12880
rect 17105 -12914 17139 -12880
rect 17173 -12914 17207 -12880
rect 17241 -12914 17275 -12880
rect 17309 -12914 17343 -12880
rect 17377 -12914 17411 -12880
rect 17445 -12914 17479 -12880
rect 17513 -12914 17547 -12880
rect 17581 -12914 17615 -12880
rect 18123 -12914 18157 -12880
rect 18191 -12914 18225 -12880
rect 18259 -12914 18293 -12880
rect 18327 -12914 18361 -12880
rect 18395 -12914 18429 -12880
rect 18463 -12914 18497 -12880
rect 18531 -12914 18565 -12880
rect 18599 -12914 18633 -12880
rect 19141 -12914 19175 -12880
rect 19209 -12914 19243 -12880
rect 19277 -12914 19311 -12880
rect 19345 -12914 19379 -12880
rect 19413 -12914 19447 -12880
rect 19481 -12914 19515 -12880
rect 19549 -12914 19583 -12880
rect 19617 -12914 19651 -12880
rect 20159 -12914 20193 -12880
rect 20227 -12914 20261 -12880
rect 20295 -12914 20329 -12880
rect 20363 -12914 20397 -12880
rect 20431 -12914 20465 -12880
rect 20499 -12914 20533 -12880
rect 20567 -12914 20601 -12880
rect 20635 -12914 20669 -12880
rect 21177 -12914 21211 -12880
rect 21245 -12914 21279 -12880
rect 21313 -12914 21347 -12880
rect 21381 -12914 21415 -12880
rect 21449 -12914 21483 -12880
rect 21517 -12914 21551 -12880
rect 21585 -12914 21619 -12880
rect 21653 -12914 21687 -12880
rect 22195 -12914 22229 -12880
rect 22263 -12914 22297 -12880
rect 22331 -12914 22365 -12880
rect 22399 -12914 22433 -12880
rect 22467 -12914 22501 -12880
rect 22535 -12914 22569 -12880
rect 22603 -12914 22637 -12880
rect 22671 -12914 22705 -12880
rect -8913 -13184 -8879 -13150
rect -8845 -13184 -8811 -13150
rect -8777 -13184 -8743 -13150
rect -8709 -13184 -8675 -13150
rect -8641 -13184 -8607 -13150
rect -8573 -13184 -8539 -13150
rect -8505 -13184 -8471 -13150
rect -8437 -13184 -8403 -13150
rect -7895 -13184 -7861 -13150
rect -7827 -13184 -7793 -13150
rect -7759 -13184 -7725 -13150
rect -7691 -13184 -7657 -13150
rect -7623 -13184 -7589 -13150
rect -7555 -13184 -7521 -13150
rect -7487 -13184 -7453 -13150
rect -7419 -13184 -7385 -13150
rect -6877 -13184 -6843 -13150
rect -6809 -13184 -6775 -13150
rect -6741 -13184 -6707 -13150
rect -6673 -13184 -6639 -13150
rect -6605 -13184 -6571 -13150
rect -6537 -13184 -6503 -13150
rect -6469 -13184 -6435 -13150
rect -6401 -13184 -6367 -13150
rect -5859 -13184 -5825 -13150
rect -5791 -13184 -5757 -13150
rect -5723 -13184 -5689 -13150
rect -5655 -13184 -5621 -13150
rect -5587 -13184 -5553 -13150
rect -5519 -13184 -5485 -13150
rect -5451 -13184 -5417 -13150
rect -5383 -13184 -5349 -13150
rect -4841 -13184 -4807 -13150
rect -4773 -13184 -4739 -13150
rect -4705 -13184 -4671 -13150
rect -4637 -13184 -4603 -13150
rect -4569 -13184 -4535 -13150
rect -4501 -13184 -4467 -13150
rect -4433 -13184 -4399 -13150
rect -4365 -13184 -4331 -13150
rect -3823 -13184 -3789 -13150
rect -3755 -13184 -3721 -13150
rect -3687 -13184 -3653 -13150
rect -3619 -13184 -3585 -13150
rect -3551 -13184 -3517 -13150
rect -3483 -13184 -3449 -13150
rect -3415 -13184 -3381 -13150
rect -3347 -13184 -3313 -13150
rect -2805 -13184 -2771 -13150
rect -2737 -13184 -2703 -13150
rect -2669 -13184 -2635 -13150
rect -2601 -13184 -2567 -13150
rect -2533 -13184 -2499 -13150
rect -2465 -13184 -2431 -13150
rect -2397 -13184 -2363 -13150
rect -2329 -13184 -2295 -13150
rect -1787 -13184 -1753 -13150
rect -1719 -13184 -1685 -13150
rect -1651 -13184 -1617 -13150
rect -1583 -13184 -1549 -13150
rect -1515 -13184 -1481 -13150
rect -1447 -13184 -1413 -13150
rect -1379 -13184 -1345 -13150
rect -1311 -13184 -1277 -13150
rect -769 -13184 -735 -13150
rect -701 -13184 -667 -13150
rect -633 -13184 -599 -13150
rect -565 -13184 -531 -13150
rect -497 -13184 -463 -13150
rect -429 -13184 -395 -13150
rect -361 -13184 -327 -13150
rect -293 -13184 -259 -13150
rect -8913 -13292 -8879 -13258
rect -8845 -13292 -8811 -13258
rect -8777 -13292 -8743 -13258
rect -8709 -13292 -8675 -13258
rect -8641 -13292 -8607 -13258
rect -8573 -13292 -8539 -13258
rect -8505 -13292 -8471 -13258
rect -8437 -13292 -8403 -13258
rect -7895 -13292 -7861 -13258
rect -7827 -13292 -7793 -13258
rect -7759 -13292 -7725 -13258
rect -7691 -13292 -7657 -13258
rect -7623 -13292 -7589 -13258
rect -7555 -13292 -7521 -13258
rect -7487 -13292 -7453 -13258
rect -7419 -13292 -7385 -13258
rect -6877 -13292 -6843 -13258
rect -6809 -13292 -6775 -13258
rect -6741 -13292 -6707 -13258
rect -6673 -13292 -6639 -13258
rect -6605 -13292 -6571 -13258
rect -6537 -13292 -6503 -13258
rect -6469 -13292 -6435 -13258
rect -6401 -13292 -6367 -13258
rect -5859 -13292 -5825 -13258
rect -5791 -13292 -5757 -13258
rect -5723 -13292 -5689 -13258
rect -5655 -13292 -5621 -13258
rect -5587 -13292 -5553 -13258
rect -5519 -13292 -5485 -13258
rect -5451 -13292 -5417 -13258
rect -5383 -13292 -5349 -13258
rect -4841 -13292 -4807 -13258
rect -4773 -13292 -4739 -13258
rect -4705 -13292 -4671 -13258
rect -4637 -13292 -4603 -13258
rect -4569 -13292 -4535 -13258
rect -4501 -13292 -4467 -13258
rect -4433 -13292 -4399 -13258
rect -4365 -13292 -4331 -13258
rect -3823 -13292 -3789 -13258
rect -3755 -13292 -3721 -13258
rect -3687 -13292 -3653 -13258
rect -3619 -13292 -3585 -13258
rect -3551 -13292 -3517 -13258
rect -3483 -13292 -3449 -13258
rect -3415 -13292 -3381 -13258
rect -3347 -13292 -3313 -13258
rect -2805 -13292 -2771 -13258
rect -2737 -13292 -2703 -13258
rect -2669 -13292 -2635 -13258
rect -2601 -13292 -2567 -13258
rect -2533 -13292 -2499 -13258
rect -2465 -13292 -2431 -13258
rect -2397 -13292 -2363 -13258
rect -2329 -13292 -2295 -13258
rect -1787 -13292 -1753 -13258
rect -1719 -13292 -1685 -13258
rect -1651 -13292 -1617 -13258
rect -1583 -13292 -1549 -13258
rect -1515 -13292 -1481 -13258
rect -1447 -13292 -1413 -13258
rect -1379 -13292 -1345 -13258
rect -1311 -13292 -1277 -13258
rect -769 -13292 -735 -13258
rect -701 -13292 -667 -13258
rect -633 -13292 -599 -13258
rect -565 -13292 -531 -13258
rect -497 -13292 -463 -13258
rect -429 -13292 -395 -13258
rect -361 -13292 -327 -13258
rect -293 -13292 -259 -13258
rect 2853 -13624 2887 -13590
rect 2921 -13624 2955 -13590
rect 2989 -13624 3023 -13590
rect 3057 -13624 3091 -13590
rect 3125 -13624 3159 -13590
rect 3193 -13624 3227 -13590
rect 3261 -13624 3295 -13590
rect 3329 -13624 3363 -13590
rect 3871 -13624 3905 -13590
rect 3939 -13624 3973 -13590
rect 4007 -13624 4041 -13590
rect 4075 -13624 4109 -13590
rect 4143 -13624 4177 -13590
rect 4211 -13624 4245 -13590
rect 4279 -13624 4313 -13590
rect 4347 -13624 4381 -13590
rect 4889 -13624 4923 -13590
rect 4957 -13624 4991 -13590
rect 5025 -13624 5059 -13590
rect 5093 -13624 5127 -13590
rect 5161 -13624 5195 -13590
rect 5229 -13624 5263 -13590
rect 5297 -13624 5331 -13590
rect 5365 -13624 5399 -13590
rect 5907 -13624 5941 -13590
rect 5975 -13624 6009 -13590
rect 6043 -13624 6077 -13590
rect 6111 -13624 6145 -13590
rect 6179 -13624 6213 -13590
rect 6247 -13624 6281 -13590
rect 6315 -13624 6349 -13590
rect 6383 -13624 6417 -13590
rect 6925 -13624 6959 -13590
rect 6993 -13624 7027 -13590
rect 7061 -13624 7095 -13590
rect 7129 -13624 7163 -13590
rect 7197 -13624 7231 -13590
rect 7265 -13624 7299 -13590
rect 7333 -13624 7367 -13590
rect 7401 -13624 7435 -13590
rect 7943 -13624 7977 -13590
rect 8011 -13624 8045 -13590
rect 8079 -13624 8113 -13590
rect 8147 -13624 8181 -13590
rect 8215 -13624 8249 -13590
rect 8283 -13624 8317 -13590
rect 8351 -13624 8385 -13590
rect 8419 -13624 8453 -13590
rect 8961 -13624 8995 -13590
rect 9029 -13624 9063 -13590
rect 9097 -13624 9131 -13590
rect 9165 -13624 9199 -13590
rect 9233 -13624 9267 -13590
rect 9301 -13624 9335 -13590
rect 9369 -13624 9403 -13590
rect 9437 -13624 9471 -13590
rect 9979 -13624 10013 -13590
rect 10047 -13624 10081 -13590
rect 10115 -13624 10149 -13590
rect 10183 -13624 10217 -13590
rect 10251 -13624 10285 -13590
rect 10319 -13624 10353 -13590
rect 10387 -13624 10421 -13590
rect 10455 -13624 10489 -13590
rect 10997 -13624 11031 -13590
rect 11065 -13624 11099 -13590
rect 11133 -13624 11167 -13590
rect 11201 -13624 11235 -13590
rect 11269 -13624 11303 -13590
rect 11337 -13624 11371 -13590
rect 11405 -13624 11439 -13590
rect 11473 -13624 11507 -13590
rect 12015 -13624 12049 -13590
rect 12083 -13624 12117 -13590
rect 12151 -13624 12185 -13590
rect 12219 -13624 12253 -13590
rect 12287 -13624 12321 -13590
rect 12355 -13624 12389 -13590
rect 12423 -13624 12457 -13590
rect 12491 -13624 12525 -13590
rect 13033 -13624 13067 -13590
rect 13101 -13624 13135 -13590
rect 13169 -13624 13203 -13590
rect 13237 -13624 13271 -13590
rect 13305 -13624 13339 -13590
rect 13373 -13624 13407 -13590
rect 13441 -13624 13475 -13590
rect 13509 -13624 13543 -13590
rect 14051 -13624 14085 -13590
rect 14119 -13624 14153 -13590
rect 14187 -13624 14221 -13590
rect 14255 -13624 14289 -13590
rect 14323 -13624 14357 -13590
rect 14391 -13624 14425 -13590
rect 14459 -13624 14493 -13590
rect 14527 -13624 14561 -13590
rect 15069 -13624 15103 -13590
rect 15137 -13624 15171 -13590
rect 15205 -13624 15239 -13590
rect 15273 -13624 15307 -13590
rect 15341 -13624 15375 -13590
rect 15409 -13624 15443 -13590
rect 15477 -13624 15511 -13590
rect 15545 -13624 15579 -13590
rect 16087 -13624 16121 -13590
rect 16155 -13624 16189 -13590
rect 16223 -13624 16257 -13590
rect 16291 -13624 16325 -13590
rect 16359 -13624 16393 -13590
rect 16427 -13624 16461 -13590
rect 16495 -13624 16529 -13590
rect 16563 -13624 16597 -13590
rect 17105 -13624 17139 -13590
rect 17173 -13624 17207 -13590
rect 17241 -13624 17275 -13590
rect 17309 -13624 17343 -13590
rect 17377 -13624 17411 -13590
rect 17445 -13624 17479 -13590
rect 17513 -13624 17547 -13590
rect 17581 -13624 17615 -13590
rect 18123 -13624 18157 -13590
rect 18191 -13624 18225 -13590
rect 18259 -13624 18293 -13590
rect 18327 -13624 18361 -13590
rect 18395 -13624 18429 -13590
rect 18463 -13624 18497 -13590
rect 18531 -13624 18565 -13590
rect 18599 -13624 18633 -13590
rect 19141 -13624 19175 -13590
rect 19209 -13624 19243 -13590
rect 19277 -13624 19311 -13590
rect 19345 -13624 19379 -13590
rect 19413 -13624 19447 -13590
rect 19481 -13624 19515 -13590
rect 19549 -13624 19583 -13590
rect 19617 -13624 19651 -13590
rect 20159 -13624 20193 -13590
rect 20227 -13624 20261 -13590
rect 20295 -13624 20329 -13590
rect 20363 -13624 20397 -13590
rect 20431 -13624 20465 -13590
rect 20499 -13624 20533 -13590
rect 20567 -13624 20601 -13590
rect 20635 -13624 20669 -13590
rect 21177 -13624 21211 -13590
rect 21245 -13624 21279 -13590
rect 21313 -13624 21347 -13590
rect 21381 -13624 21415 -13590
rect 21449 -13624 21483 -13590
rect 21517 -13624 21551 -13590
rect 21585 -13624 21619 -13590
rect 21653 -13624 21687 -13590
rect 22195 -13624 22229 -13590
rect 22263 -13624 22297 -13590
rect 22331 -13624 22365 -13590
rect 22399 -13624 22433 -13590
rect 22467 -13624 22501 -13590
rect 22535 -13624 22569 -13590
rect 22603 -13624 22637 -13590
rect 22671 -13624 22705 -13590
rect -8913 -14002 -8879 -13968
rect -8845 -14002 -8811 -13968
rect -8777 -14002 -8743 -13968
rect -8709 -14002 -8675 -13968
rect -8641 -14002 -8607 -13968
rect -8573 -14002 -8539 -13968
rect -8505 -14002 -8471 -13968
rect -8437 -14002 -8403 -13968
rect -7895 -14002 -7861 -13968
rect -7827 -14002 -7793 -13968
rect -7759 -14002 -7725 -13968
rect -7691 -14002 -7657 -13968
rect -7623 -14002 -7589 -13968
rect -7555 -14002 -7521 -13968
rect -7487 -14002 -7453 -13968
rect -7419 -14002 -7385 -13968
rect -6877 -14002 -6843 -13968
rect -6809 -14002 -6775 -13968
rect -6741 -14002 -6707 -13968
rect -6673 -14002 -6639 -13968
rect -6605 -14002 -6571 -13968
rect -6537 -14002 -6503 -13968
rect -6469 -14002 -6435 -13968
rect -6401 -14002 -6367 -13968
rect -5859 -14002 -5825 -13968
rect -5791 -14002 -5757 -13968
rect -5723 -14002 -5689 -13968
rect -5655 -14002 -5621 -13968
rect -5587 -14002 -5553 -13968
rect -5519 -14002 -5485 -13968
rect -5451 -14002 -5417 -13968
rect -5383 -14002 -5349 -13968
rect -4841 -14002 -4807 -13968
rect -4773 -14002 -4739 -13968
rect -4705 -14002 -4671 -13968
rect -4637 -14002 -4603 -13968
rect -4569 -14002 -4535 -13968
rect -4501 -14002 -4467 -13968
rect -4433 -14002 -4399 -13968
rect -4365 -14002 -4331 -13968
rect -3823 -14002 -3789 -13968
rect -3755 -14002 -3721 -13968
rect -3687 -14002 -3653 -13968
rect -3619 -14002 -3585 -13968
rect -3551 -14002 -3517 -13968
rect -3483 -14002 -3449 -13968
rect -3415 -14002 -3381 -13968
rect -3347 -14002 -3313 -13968
rect -2805 -14002 -2771 -13968
rect -2737 -14002 -2703 -13968
rect -2669 -14002 -2635 -13968
rect -2601 -14002 -2567 -13968
rect -2533 -14002 -2499 -13968
rect -2465 -14002 -2431 -13968
rect -2397 -14002 -2363 -13968
rect -2329 -14002 -2295 -13968
rect -1787 -14002 -1753 -13968
rect -1719 -14002 -1685 -13968
rect -1651 -14002 -1617 -13968
rect -1583 -14002 -1549 -13968
rect -1515 -14002 -1481 -13968
rect -1447 -14002 -1413 -13968
rect -1379 -14002 -1345 -13968
rect -1311 -14002 -1277 -13968
rect -769 -14002 -735 -13968
rect -701 -14002 -667 -13968
rect -633 -14002 -599 -13968
rect -565 -14002 -531 -13968
rect -497 -14002 -463 -13968
rect -429 -14002 -395 -13968
rect -361 -14002 -327 -13968
rect -293 -14002 -259 -13968
rect -8913 -14110 -8879 -14076
rect -8845 -14110 -8811 -14076
rect -8777 -14110 -8743 -14076
rect -8709 -14110 -8675 -14076
rect -8641 -14110 -8607 -14076
rect -8573 -14110 -8539 -14076
rect -8505 -14110 -8471 -14076
rect -8437 -14110 -8403 -14076
rect -7895 -14110 -7861 -14076
rect -7827 -14110 -7793 -14076
rect -7759 -14110 -7725 -14076
rect -7691 -14110 -7657 -14076
rect -7623 -14110 -7589 -14076
rect -7555 -14110 -7521 -14076
rect -7487 -14110 -7453 -14076
rect -7419 -14110 -7385 -14076
rect -6877 -14110 -6843 -14076
rect -6809 -14110 -6775 -14076
rect -6741 -14110 -6707 -14076
rect -6673 -14110 -6639 -14076
rect -6605 -14110 -6571 -14076
rect -6537 -14110 -6503 -14076
rect -6469 -14110 -6435 -14076
rect -6401 -14110 -6367 -14076
rect -5859 -14110 -5825 -14076
rect -5791 -14110 -5757 -14076
rect -5723 -14110 -5689 -14076
rect -5655 -14110 -5621 -14076
rect -5587 -14110 -5553 -14076
rect -5519 -14110 -5485 -14076
rect -5451 -14110 -5417 -14076
rect -5383 -14110 -5349 -14076
rect -4841 -14110 -4807 -14076
rect -4773 -14110 -4739 -14076
rect -4705 -14110 -4671 -14076
rect -4637 -14110 -4603 -14076
rect -4569 -14110 -4535 -14076
rect -4501 -14110 -4467 -14076
rect -4433 -14110 -4399 -14076
rect -4365 -14110 -4331 -14076
rect -3823 -14110 -3789 -14076
rect -3755 -14110 -3721 -14076
rect -3687 -14110 -3653 -14076
rect -3619 -14110 -3585 -14076
rect -3551 -14110 -3517 -14076
rect -3483 -14110 -3449 -14076
rect -3415 -14110 -3381 -14076
rect -3347 -14110 -3313 -14076
rect -2805 -14110 -2771 -14076
rect -2737 -14110 -2703 -14076
rect -2669 -14110 -2635 -14076
rect -2601 -14110 -2567 -14076
rect -2533 -14110 -2499 -14076
rect -2465 -14110 -2431 -14076
rect -2397 -14110 -2363 -14076
rect -2329 -14110 -2295 -14076
rect -1787 -14110 -1753 -14076
rect -1719 -14110 -1685 -14076
rect -1651 -14110 -1617 -14076
rect -1583 -14110 -1549 -14076
rect -1515 -14110 -1481 -14076
rect -1447 -14110 -1413 -14076
rect -1379 -14110 -1345 -14076
rect -1311 -14110 -1277 -14076
rect -769 -14110 -735 -14076
rect -701 -14110 -667 -14076
rect -633 -14110 -599 -14076
rect -565 -14110 -531 -14076
rect -497 -14110 -463 -14076
rect -429 -14110 -395 -14076
rect -361 -14110 -327 -14076
rect -293 -14110 -259 -14076
rect 2853 -14146 2887 -14112
rect 2921 -14146 2955 -14112
rect 2989 -14146 3023 -14112
rect 3057 -14146 3091 -14112
rect 3125 -14146 3159 -14112
rect 3193 -14146 3227 -14112
rect 3261 -14146 3295 -14112
rect 3329 -14146 3363 -14112
rect 3871 -14146 3905 -14112
rect 3939 -14146 3973 -14112
rect 4007 -14146 4041 -14112
rect 4075 -14146 4109 -14112
rect 4143 -14146 4177 -14112
rect 4211 -14146 4245 -14112
rect 4279 -14146 4313 -14112
rect 4347 -14146 4381 -14112
rect 4889 -14146 4923 -14112
rect 4957 -14146 4991 -14112
rect 5025 -14146 5059 -14112
rect 5093 -14146 5127 -14112
rect 5161 -14146 5195 -14112
rect 5229 -14146 5263 -14112
rect 5297 -14146 5331 -14112
rect 5365 -14146 5399 -14112
rect 5907 -14146 5941 -14112
rect 5975 -14146 6009 -14112
rect 6043 -14146 6077 -14112
rect 6111 -14146 6145 -14112
rect 6179 -14146 6213 -14112
rect 6247 -14146 6281 -14112
rect 6315 -14146 6349 -14112
rect 6383 -14146 6417 -14112
rect 6925 -14146 6959 -14112
rect 6993 -14146 7027 -14112
rect 7061 -14146 7095 -14112
rect 7129 -14146 7163 -14112
rect 7197 -14146 7231 -14112
rect 7265 -14146 7299 -14112
rect 7333 -14146 7367 -14112
rect 7401 -14146 7435 -14112
rect 7943 -14146 7977 -14112
rect 8011 -14146 8045 -14112
rect 8079 -14146 8113 -14112
rect 8147 -14146 8181 -14112
rect 8215 -14146 8249 -14112
rect 8283 -14146 8317 -14112
rect 8351 -14146 8385 -14112
rect 8419 -14146 8453 -14112
rect 8961 -14146 8995 -14112
rect 9029 -14146 9063 -14112
rect 9097 -14146 9131 -14112
rect 9165 -14146 9199 -14112
rect 9233 -14146 9267 -14112
rect 9301 -14146 9335 -14112
rect 9369 -14146 9403 -14112
rect 9437 -14146 9471 -14112
rect 9979 -14146 10013 -14112
rect 10047 -14146 10081 -14112
rect 10115 -14146 10149 -14112
rect 10183 -14146 10217 -14112
rect 10251 -14146 10285 -14112
rect 10319 -14146 10353 -14112
rect 10387 -14146 10421 -14112
rect 10455 -14146 10489 -14112
rect 10997 -14146 11031 -14112
rect 11065 -14146 11099 -14112
rect 11133 -14146 11167 -14112
rect 11201 -14146 11235 -14112
rect 11269 -14146 11303 -14112
rect 11337 -14146 11371 -14112
rect 11405 -14146 11439 -14112
rect 11473 -14146 11507 -14112
rect 12015 -14146 12049 -14112
rect 12083 -14146 12117 -14112
rect 12151 -14146 12185 -14112
rect 12219 -14146 12253 -14112
rect 12287 -14146 12321 -14112
rect 12355 -14146 12389 -14112
rect 12423 -14146 12457 -14112
rect 12491 -14146 12525 -14112
rect 13033 -14146 13067 -14112
rect 13101 -14146 13135 -14112
rect 13169 -14146 13203 -14112
rect 13237 -14146 13271 -14112
rect 13305 -14146 13339 -14112
rect 13373 -14146 13407 -14112
rect 13441 -14146 13475 -14112
rect 13509 -14146 13543 -14112
rect 14051 -14146 14085 -14112
rect 14119 -14146 14153 -14112
rect 14187 -14146 14221 -14112
rect 14255 -14146 14289 -14112
rect 14323 -14146 14357 -14112
rect 14391 -14146 14425 -14112
rect 14459 -14146 14493 -14112
rect 14527 -14146 14561 -14112
rect 15069 -14146 15103 -14112
rect 15137 -14146 15171 -14112
rect 15205 -14146 15239 -14112
rect 15273 -14146 15307 -14112
rect 15341 -14146 15375 -14112
rect 15409 -14146 15443 -14112
rect 15477 -14146 15511 -14112
rect 15545 -14146 15579 -14112
rect 16087 -14146 16121 -14112
rect 16155 -14146 16189 -14112
rect 16223 -14146 16257 -14112
rect 16291 -14146 16325 -14112
rect 16359 -14146 16393 -14112
rect 16427 -14146 16461 -14112
rect 16495 -14146 16529 -14112
rect 16563 -14146 16597 -14112
rect 17105 -14146 17139 -14112
rect 17173 -14146 17207 -14112
rect 17241 -14146 17275 -14112
rect 17309 -14146 17343 -14112
rect 17377 -14146 17411 -14112
rect 17445 -14146 17479 -14112
rect 17513 -14146 17547 -14112
rect 17581 -14146 17615 -14112
rect 18123 -14146 18157 -14112
rect 18191 -14146 18225 -14112
rect 18259 -14146 18293 -14112
rect 18327 -14146 18361 -14112
rect 18395 -14146 18429 -14112
rect 18463 -14146 18497 -14112
rect 18531 -14146 18565 -14112
rect 18599 -14146 18633 -14112
rect 19141 -14146 19175 -14112
rect 19209 -14146 19243 -14112
rect 19277 -14146 19311 -14112
rect 19345 -14146 19379 -14112
rect 19413 -14146 19447 -14112
rect 19481 -14146 19515 -14112
rect 19549 -14146 19583 -14112
rect 19617 -14146 19651 -14112
rect 20159 -14146 20193 -14112
rect 20227 -14146 20261 -14112
rect 20295 -14146 20329 -14112
rect 20363 -14146 20397 -14112
rect 20431 -14146 20465 -14112
rect 20499 -14146 20533 -14112
rect 20567 -14146 20601 -14112
rect 20635 -14146 20669 -14112
rect 21177 -14146 21211 -14112
rect 21245 -14146 21279 -14112
rect 21313 -14146 21347 -14112
rect 21381 -14146 21415 -14112
rect 21449 -14146 21483 -14112
rect 21517 -14146 21551 -14112
rect 21585 -14146 21619 -14112
rect 21653 -14146 21687 -14112
rect 22195 -14146 22229 -14112
rect 22263 -14146 22297 -14112
rect 22331 -14146 22365 -14112
rect 22399 -14146 22433 -14112
rect 22467 -14146 22501 -14112
rect 22535 -14146 22569 -14112
rect 22603 -14146 22637 -14112
rect 22671 -14146 22705 -14112
rect -8913 -14820 -8879 -14786
rect -8845 -14820 -8811 -14786
rect -8777 -14820 -8743 -14786
rect -8709 -14820 -8675 -14786
rect -8641 -14820 -8607 -14786
rect -8573 -14820 -8539 -14786
rect -8505 -14820 -8471 -14786
rect -8437 -14820 -8403 -14786
rect -7895 -14820 -7861 -14786
rect -7827 -14820 -7793 -14786
rect -7759 -14820 -7725 -14786
rect -7691 -14820 -7657 -14786
rect -7623 -14820 -7589 -14786
rect -7555 -14820 -7521 -14786
rect -7487 -14820 -7453 -14786
rect -7419 -14820 -7385 -14786
rect -6877 -14820 -6843 -14786
rect -6809 -14820 -6775 -14786
rect -6741 -14820 -6707 -14786
rect -6673 -14820 -6639 -14786
rect -6605 -14820 -6571 -14786
rect -6537 -14820 -6503 -14786
rect -6469 -14820 -6435 -14786
rect -6401 -14820 -6367 -14786
rect -5859 -14820 -5825 -14786
rect -5791 -14820 -5757 -14786
rect -5723 -14820 -5689 -14786
rect -5655 -14820 -5621 -14786
rect -5587 -14820 -5553 -14786
rect -5519 -14820 -5485 -14786
rect -5451 -14820 -5417 -14786
rect -5383 -14820 -5349 -14786
rect -4841 -14820 -4807 -14786
rect -4773 -14820 -4739 -14786
rect -4705 -14820 -4671 -14786
rect -4637 -14820 -4603 -14786
rect -4569 -14820 -4535 -14786
rect -4501 -14820 -4467 -14786
rect -4433 -14820 -4399 -14786
rect -4365 -14820 -4331 -14786
rect -3823 -14820 -3789 -14786
rect -3755 -14820 -3721 -14786
rect -3687 -14820 -3653 -14786
rect -3619 -14820 -3585 -14786
rect -3551 -14820 -3517 -14786
rect -3483 -14820 -3449 -14786
rect -3415 -14820 -3381 -14786
rect -3347 -14820 -3313 -14786
rect -2805 -14820 -2771 -14786
rect -2737 -14820 -2703 -14786
rect -2669 -14820 -2635 -14786
rect -2601 -14820 -2567 -14786
rect -2533 -14820 -2499 -14786
rect -2465 -14820 -2431 -14786
rect -2397 -14820 -2363 -14786
rect -2329 -14820 -2295 -14786
rect -1787 -14820 -1753 -14786
rect -1719 -14820 -1685 -14786
rect -1651 -14820 -1617 -14786
rect -1583 -14820 -1549 -14786
rect -1515 -14820 -1481 -14786
rect -1447 -14820 -1413 -14786
rect -1379 -14820 -1345 -14786
rect -1311 -14820 -1277 -14786
rect -769 -14820 -735 -14786
rect -701 -14820 -667 -14786
rect -633 -14820 -599 -14786
rect -565 -14820 -531 -14786
rect -497 -14820 -463 -14786
rect -429 -14820 -395 -14786
rect -361 -14820 -327 -14786
rect -293 -14820 -259 -14786
rect 2853 -14856 2887 -14822
rect 2921 -14856 2955 -14822
rect 2989 -14856 3023 -14822
rect 3057 -14856 3091 -14822
rect 3125 -14856 3159 -14822
rect 3193 -14856 3227 -14822
rect 3261 -14856 3295 -14822
rect 3329 -14856 3363 -14822
rect 3871 -14856 3905 -14822
rect 3939 -14856 3973 -14822
rect 4007 -14856 4041 -14822
rect 4075 -14856 4109 -14822
rect 4143 -14856 4177 -14822
rect 4211 -14856 4245 -14822
rect 4279 -14856 4313 -14822
rect 4347 -14856 4381 -14822
rect 4889 -14856 4923 -14822
rect 4957 -14856 4991 -14822
rect 5025 -14856 5059 -14822
rect 5093 -14856 5127 -14822
rect 5161 -14856 5195 -14822
rect 5229 -14856 5263 -14822
rect 5297 -14856 5331 -14822
rect 5365 -14856 5399 -14822
rect 5907 -14856 5941 -14822
rect 5975 -14856 6009 -14822
rect 6043 -14856 6077 -14822
rect 6111 -14856 6145 -14822
rect 6179 -14856 6213 -14822
rect 6247 -14856 6281 -14822
rect 6315 -14856 6349 -14822
rect 6383 -14856 6417 -14822
rect 6925 -14856 6959 -14822
rect 6993 -14856 7027 -14822
rect 7061 -14856 7095 -14822
rect 7129 -14856 7163 -14822
rect 7197 -14856 7231 -14822
rect 7265 -14856 7299 -14822
rect 7333 -14856 7367 -14822
rect 7401 -14856 7435 -14822
rect 7943 -14856 7977 -14822
rect 8011 -14856 8045 -14822
rect 8079 -14856 8113 -14822
rect 8147 -14856 8181 -14822
rect 8215 -14856 8249 -14822
rect 8283 -14856 8317 -14822
rect 8351 -14856 8385 -14822
rect 8419 -14856 8453 -14822
rect 8961 -14856 8995 -14822
rect 9029 -14856 9063 -14822
rect 9097 -14856 9131 -14822
rect 9165 -14856 9199 -14822
rect 9233 -14856 9267 -14822
rect 9301 -14856 9335 -14822
rect 9369 -14856 9403 -14822
rect 9437 -14856 9471 -14822
rect 9979 -14856 10013 -14822
rect 10047 -14856 10081 -14822
rect 10115 -14856 10149 -14822
rect 10183 -14856 10217 -14822
rect 10251 -14856 10285 -14822
rect 10319 -14856 10353 -14822
rect 10387 -14856 10421 -14822
rect 10455 -14856 10489 -14822
rect 10997 -14856 11031 -14822
rect 11065 -14856 11099 -14822
rect 11133 -14856 11167 -14822
rect 11201 -14856 11235 -14822
rect 11269 -14856 11303 -14822
rect 11337 -14856 11371 -14822
rect 11405 -14856 11439 -14822
rect 11473 -14856 11507 -14822
rect 12015 -14856 12049 -14822
rect 12083 -14856 12117 -14822
rect 12151 -14856 12185 -14822
rect 12219 -14856 12253 -14822
rect 12287 -14856 12321 -14822
rect 12355 -14856 12389 -14822
rect 12423 -14856 12457 -14822
rect 12491 -14856 12525 -14822
rect 13033 -14856 13067 -14822
rect 13101 -14856 13135 -14822
rect 13169 -14856 13203 -14822
rect 13237 -14856 13271 -14822
rect 13305 -14856 13339 -14822
rect 13373 -14856 13407 -14822
rect 13441 -14856 13475 -14822
rect 13509 -14856 13543 -14822
rect 14051 -14856 14085 -14822
rect 14119 -14856 14153 -14822
rect 14187 -14856 14221 -14822
rect 14255 -14856 14289 -14822
rect 14323 -14856 14357 -14822
rect 14391 -14856 14425 -14822
rect 14459 -14856 14493 -14822
rect 14527 -14856 14561 -14822
rect 15069 -14856 15103 -14822
rect 15137 -14856 15171 -14822
rect 15205 -14856 15239 -14822
rect 15273 -14856 15307 -14822
rect 15341 -14856 15375 -14822
rect 15409 -14856 15443 -14822
rect 15477 -14856 15511 -14822
rect 15545 -14856 15579 -14822
rect 16087 -14856 16121 -14822
rect 16155 -14856 16189 -14822
rect 16223 -14856 16257 -14822
rect 16291 -14856 16325 -14822
rect 16359 -14856 16393 -14822
rect 16427 -14856 16461 -14822
rect 16495 -14856 16529 -14822
rect 16563 -14856 16597 -14822
rect 17105 -14856 17139 -14822
rect 17173 -14856 17207 -14822
rect 17241 -14856 17275 -14822
rect 17309 -14856 17343 -14822
rect 17377 -14856 17411 -14822
rect 17445 -14856 17479 -14822
rect 17513 -14856 17547 -14822
rect 17581 -14856 17615 -14822
rect 18123 -14856 18157 -14822
rect 18191 -14856 18225 -14822
rect 18259 -14856 18293 -14822
rect 18327 -14856 18361 -14822
rect 18395 -14856 18429 -14822
rect 18463 -14856 18497 -14822
rect 18531 -14856 18565 -14822
rect 18599 -14856 18633 -14822
rect 19141 -14856 19175 -14822
rect 19209 -14856 19243 -14822
rect 19277 -14856 19311 -14822
rect 19345 -14856 19379 -14822
rect 19413 -14856 19447 -14822
rect 19481 -14856 19515 -14822
rect 19549 -14856 19583 -14822
rect 19617 -14856 19651 -14822
rect 20159 -14856 20193 -14822
rect 20227 -14856 20261 -14822
rect 20295 -14856 20329 -14822
rect 20363 -14856 20397 -14822
rect 20431 -14856 20465 -14822
rect 20499 -14856 20533 -14822
rect 20567 -14856 20601 -14822
rect 20635 -14856 20669 -14822
rect 21177 -14856 21211 -14822
rect 21245 -14856 21279 -14822
rect 21313 -14856 21347 -14822
rect 21381 -14856 21415 -14822
rect 21449 -14856 21483 -14822
rect 21517 -14856 21551 -14822
rect 21585 -14856 21619 -14822
rect 21653 -14856 21687 -14822
rect 22195 -14856 22229 -14822
rect 22263 -14856 22297 -14822
rect 22331 -14856 22365 -14822
rect 22399 -14856 22433 -14822
rect 22467 -14856 22501 -14822
rect 22535 -14856 22569 -14822
rect 22603 -14856 22637 -14822
rect 22671 -14856 22705 -14822
rect -8913 -14928 -8879 -14894
rect -8845 -14928 -8811 -14894
rect -8777 -14928 -8743 -14894
rect -8709 -14928 -8675 -14894
rect -8641 -14928 -8607 -14894
rect -8573 -14928 -8539 -14894
rect -8505 -14928 -8471 -14894
rect -8437 -14928 -8403 -14894
rect -7895 -14928 -7861 -14894
rect -7827 -14928 -7793 -14894
rect -7759 -14928 -7725 -14894
rect -7691 -14928 -7657 -14894
rect -7623 -14928 -7589 -14894
rect -7555 -14928 -7521 -14894
rect -7487 -14928 -7453 -14894
rect -7419 -14928 -7385 -14894
rect -6877 -14928 -6843 -14894
rect -6809 -14928 -6775 -14894
rect -6741 -14928 -6707 -14894
rect -6673 -14928 -6639 -14894
rect -6605 -14928 -6571 -14894
rect -6537 -14928 -6503 -14894
rect -6469 -14928 -6435 -14894
rect -6401 -14928 -6367 -14894
rect -5859 -14928 -5825 -14894
rect -5791 -14928 -5757 -14894
rect -5723 -14928 -5689 -14894
rect -5655 -14928 -5621 -14894
rect -5587 -14928 -5553 -14894
rect -5519 -14928 -5485 -14894
rect -5451 -14928 -5417 -14894
rect -5383 -14928 -5349 -14894
rect -4841 -14928 -4807 -14894
rect -4773 -14928 -4739 -14894
rect -4705 -14928 -4671 -14894
rect -4637 -14928 -4603 -14894
rect -4569 -14928 -4535 -14894
rect -4501 -14928 -4467 -14894
rect -4433 -14928 -4399 -14894
rect -4365 -14928 -4331 -14894
rect -3823 -14928 -3789 -14894
rect -3755 -14928 -3721 -14894
rect -3687 -14928 -3653 -14894
rect -3619 -14928 -3585 -14894
rect -3551 -14928 -3517 -14894
rect -3483 -14928 -3449 -14894
rect -3415 -14928 -3381 -14894
rect -3347 -14928 -3313 -14894
rect -2805 -14928 -2771 -14894
rect -2737 -14928 -2703 -14894
rect -2669 -14928 -2635 -14894
rect -2601 -14928 -2567 -14894
rect -2533 -14928 -2499 -14894
rect -2465 -14928 -2431 -14894
rect -2397 -14928 -2363 -14894
rect -2329 -14928 -2295 -14894
rect -1787 -14928 -1753 -14894
rect -1719 -14928 -1685 -14894
rect -1651 -14928 -1617 -14894
rect -1583 -14928 -1549 -14894
rect -1515 -14928 -1481 -14894
rect -1447 -14928 -1413 -14894
rect -1379 -14928 -1345 -14894
rect -1311 -14928 -1277 -14894
rect -769 -14928 -735 -14894
rect -701 -14928 -667 -14894
rect -633 -14928 -599 -14894
rect -565 -14928 -531 -14894
rect -497 -14928 -463 -14894
rect -429 -14928 -395 -14894
rect -361 -14928 -327 -14894
rect -293 -14928 -259 -14894
rect 2851 -15380 2885 -15346
rect 2919 -15380 2953 -15346
rect 2987 -15380 3021 -15346
rect 3055 -15380 3089 -15346
rect 3123 -15380 3157 -15346
rect 3191 -15380 3225 -15346
rect 3259 -15380 3293 -15346
rect 3327 -15380 3361 -15346
rect 3869 -15380 3903 -15346
rect 3937 -15380 3971 -15346
rect 4005 -15380 4039 -15346
rect 4073 -15380 4107 -15346
rect 4141 -15380 4175 -15346
rect 4209 -15380 4243 -15346
rect 4277 -15380 4311 -15346
rect 4345 -15380 4379 -15346
rect 4887 -15380 4921 -15346
rect 4955 -15380 4989 -15346
rect 5023 -15380 5057 -15346
rect 5091 -15380 5125 -15346
rect 5159 -15380 5193 -15346
rect 5227 -15380 5261 -15346
rect 5295 -15380 5329 -15346
rect 5363 -15380 5397 -15346
rect 5905 -15380 5939 -15346
rect 5973 -15380 6007 -15346
rect 6041 -15380 6075 -15346
rect 6109 -15380 6143 -15346
rect 6177 -15380 6211 -15346
rect 6245 -15380 6279 -15346
rect 6313 -15380 6347 -15346
rect 6381 -15380 6415 -15346
rect 6923 -15380 6957 -15346
rect 6991 -15380 7025 -15346
rect 7059 -15380 7093 -15346
rect 7127 -15380 7161 -15346
rect 7195 -15380 7229 -15346
rect 7263 -15380 7297 -15346
rect 7331 -15380 7365 -15346
rect 7399 -15380 7433 -15346
rect 7941 -15380 7975 -15346
rect 8009 -15380 8043 -15346
rect 8077 -15380 8111 -15346
rect 8145 -15380 8179 -15346
rect 8213 -15380 8247 -15346
rect 8281 -15380 8315 -15346
rect 8349 -15380 8383 -15346
rect 8417 -15380 8451 -15346
rect 8959 -15380 8993 -15346
rect 9027 -15380 9061 -15346
rect 9095 -15380 9129 -15346
rect 9163 -15380 9197 -15346
rect 9231 -15380 9265 -15346
rect 9299 -15380 9333 -15346
rect 9367 -15380 9401 -15346
rect 9435 -15380 9469 -15346
rect 9977 -15380 10011 -15346
rect 10045 -15380 10079 -15346
rect 10113 -15380 10147 -15346
rect 10181 -15380 10215 -15346
rect 10249 -15380 10283 -15346
rect 10317 -15380 10351 -15346
rect 10385 -15380 10419 -15346
rect 10453 -15380 10487 -15346
rect 10995 -15380 11029 -15346
rect 11063 -15380 11097 -15346
rect 11131 -15380 11165 -15346
rect 11199 -15380 11233 -15346
rect 11267 -15380 11301 -15346
rect 11335 -15380 11369 -15346
rect 11403 -15380 11437 -15346
rect 11471 -15380 11505 -15346
rect 12013 -15380 12047 -15346
rect 12081 -15380 12115 -15346
rect 12149 -15380 12183 -15346
rect 12217 -15380 12251 -15346
rect 12285 -15380 12319 -15346
rect 12353 -15380 12387 -15346
rect 12421 -15380 12455 -15346
rect 12489 -15380 12523 -15346
rect 13031 -15380 13065 -15346
rect 13099 -15380 13133 -15346
rect 13167 -15380 13201 -15346
rect 13235 -15380 13269 -15346
rect 13303 -15380 13337 -15346
rect 13371 -15380 13405 -15346
rect 13439 -15380 13473 -15346
rect 13507 -15380 13541 -15346
rect 14049 -15380 14083 -15346
rect 14117 -15380 14151 -15346
rect 14185 -15380 14219 -15346
rect 14253 -15380 14287 -15346
rect 14321 -15380 14355 -15346
rect 14389 -15380 14423 -15346
rect 14457 -15380 14491 -15346
rect 14525 -15380 14559 -15346
rect 15067 -15380 15101 -15346
rect 15135 -15380 15169 -15346
rect 15203 -15380 15237 -15346
rect 15271 -15380 15305 -15346
rect 15339 -15380 15373 -15346
rect 15407 -15380 15441 -15346
rect 15475 -15380 15509 -15346
rect 15543 -15380 15577 -15346
rect 16085 -15380 16119 -15346
rect 16153 -15380 16187 -15346
rect 16221 -15380 16255 -15346
rect 16289 -15380 16323 -15346
rect 16357 -15380 16391 -15346
rect 16425 -15380 16459 -15346
rect 16493 -15380 16527 -15346
rect 16561 -15380 16595 -15346
rect 17103 -15380 17137 -15346
rect 17171 -15380 17205 -15346
rect 17239 -15380 17273 -15346
rect 17307 -15380 17341 -15346
rect 17375 -15380 17409 -15346
rect 17443 -15380 17477 -15346
rect 17511 -15380 17545 -15346
rect 17579 -15380 17613 -15346
rect 18121 -15380 18155 -15346
rect 18189 -15380 18223 -15346
rect 18257 -15380 18291 -15346
rect 18325 -15380 18359 -15346
rect 18393 -15380 18427 -15346
rect 18461 -15380 18495 -15346
rect 18529 -15380 18563 -15346
rect 18597 -15380 18631 -15346
rect 19139 -15380 19173 -15346
rect 19207 -15380 19241 -15346
rect 19275 -15380 19309 -15346
rect 19343 -15380 19377 -15346
rect 19411 -15380 19445 -15346
rect 19479 -15380 19513 -15346
rect 19547 -15380 19581 -15346
rect 19615 -15380 19649 -15346
rect 20157 -15380 20191 -15346
rect 20225 -15380 20259 -15346
rect 20293 -15380 20327 -15346
rect 20361 -15380 20395 -15346
rect 20429 -15380 20463 -15346
rect 20497 -15380 20531 -15346
rect 20565 -15380 20599 -15346
rect 20633 -15380 20667 -15346
rect 21175 -15380 21209 -15346
rect 21243 -15380 21277 -15346
rect 21311 -15380 21345 -15346
rect 21379 -15380 21413 -15346
rect 21447 -15380 21481 -15346
rect 21515 -15380 21549 -15346
rect 21583 -15380 21617 -15346
rect 21651 -15380 21685 -15346
rect 22193 -15380 22227 -15346
rect 22261 -15380 22295 -15346
rect 22329 -15380 22363 -15346
rect 22397 -15380 22431 -15346
rect 22465 -15380 22499 -15346
rect 22533 -15380 22567 -15346
rect 22601 -15380 22635 -15346
rect 22669 -15380 22703 -15346
rect -8913 -15638 -8879 -15604
rect -8845 -15638 -8811 -15604
rect -8777 -15638 -8743 -15604
rect -8709 -15638 -8675 -15604
rect -8641 -15638 -8607 -15604
rect -8573 -15638 -8539 -15604
rect -8505 -15638 -8471 -15604
rect -8437 -15638 -8403 -15604
rect -7895 -15638 -7861 -15604
rect -7827 -15638 -7793 -15604
rect -7759 -15638 -7725 -15604
rect -7691 -15638 -7657 -15604
rect -7623 -15638 -7589 -15604
rect -7555 -15638 -7521 -15604
rect -7487 -15638 -7453 -15604
rect -7419 -15638 -7385 -15604
rect -6877 -15638 -6843 -15604
rect -6809 -15638 -6775 -15604
rect -6741 -15638 -6707 -15604
rect -6673 -15638 -6639 -15604
rect -6605 -15638 -6571 -15604
rect -6537 -15638 -6503 -15604
rect -6469 -15638 -6435 -15604
rect -6401 -15638 -6367 -15604
rect -5859 -15638 -5825 -15604
rect -5791 -15638 -5757 -15604
rect -5723 -15638 -5689 -15604
rect -5655 -15638 -5621 -15604
rect -5587 -15638 -5553 -15604
rect -5519 -15638 -5485 -15604
rect -5451 -15638 -5417 -15604
rect -5383 -15638 -5349 -15604
rect -4841 -15638 -4807 -15604
rect -4773 -15638 -4739 -15604
rect -4705 -15638 -4671 -15604
rect -4637 -15638 -4603 -15604
rect -4569 -15638 -4535 -15604
rect -4501 -15638 -4467 -15604
rect -4433 -15638 -4399 -15604
rect -4365 -15638 -4331 -15604
rect -3823 -15638 -3789 -15604
rect -3755 -15638 -3721 -15604
rect -3687 -15638 -3653 -15604
rect -3619 -15638 -3585 -15604
rect -3551 -15638 -3517 -15604
rect -3483 -15638 -3449 -15604
rect -3415 -15638 -3381 -15604
rect -3347 -15638 -3313 -15604
rect -2805 -15638 -2771 -15604
rect -2737 -15638 -2703 -15604
rect -2669 -15638 -2635 -15604
rect -2601 -15638 -2567 -15604
rect -2533 -15638 -2499 -15604
rect -2465 -15638 -2431 -15604
rect -2397 -15638 -2363 -15604
rect -2329 -15638 -2295 -15604
rect -1787 -15638 -1753 -15604
rect -1719 -15638 -1685 -15604
rect -1651 -15638 -1617 -15604
rect -1583 -15638 -1549 -15604
rect -1515 -15638 -1481 -15604
rect -1447 -15638 -1413 -15604
rect -1379 -15638 -1345 -15604
rect -1311 -15638 -1277 -15604
rect -769 -15638 -735 -15604
rect -701 -15638 -667 -15604
rect -633 -15638 -599 -15604
rect -565 -15638 -531 -15604
rect -497 -15638 -463 -15604
rect -429 -15638 -395 -15604
rect -361 -15638 -327 -15604
rect -293 -15638 -259 -15604
rect -8913 -15746 -8879 -15712
rect -8845 -15746 -8811 -15712
rect -8777 -15746 -8743 -15712
rect -8709 -15746 -8675 -15712
rect -8641 -15746 -8607 -15712
rect -8573 -15746 -8539 -15712
rect -8505 -15746 -8471 -15712
rect -8437 -15746 -8403 -15712
rect -7895 -15746 -7861 -15712
rect -7827 -15746 -7793 -15712
rect -7759 -15746 -7725 -15712
rect -7691 -15746 -7657 -15712
rect -7623 -15746 -7589 -15712
rect -7555 -15746 -7521 -15712
rect -7487 -15746 -7453 -15712
rect -7419 -15746 -7385 -15712
rect -6877 -15746 -6843 -15712
rect -6809 -15746 -6775 -15712
rect -6741 -15746 -6707 -15712
rect -6673 -15746 -6639 -15712
rect -6605 -15746 -6571 -15712
rect -6537 -15746 -6503 -15712
rect -6469 -15746 -6435 -15712
rect -6401 -15746 -6367 -15712
rect -5859 -15746 -5825 -15712
rect -5791 -15746 -5757 -15712
rect -5723 -15746 -5689 -15712
rect -5655 -15746 -5621 -15712
rect -5587 -15746 -5553 -15712
rect -5519 -15746 -5485 -15712
rect -5451 -15746 -5417 -15712
rect -5383 -15746 -5349 -15712
rect -4841 -15746 -4807 -15712
rect -4773 -15746 -4739 -15712
rect -4705 -15746 -4671 -15712
rect -4637 -15746 -4603 -15712
rect -4569 -15746 -4535 -15712
rect -4501 -15746 -4467 -15712
rect -4433 -15746 -4399 -15712
rect -4365 -15746 -4331 -15712
rect -3823 -15746 -3789 -15712
rect -3755 -15746 -3721 -15712
rect -3687 -15746 -3653 -15712
rect -3619 -15746 -3585 -15712
rect -3551 -15746 -3517 -15712
rect -3483 -15746 -3449 -15712
rect -3415 -15746 -3381 -15712
rect -3347 -15746 -3313 -15712
rect -2805 -15746 -2771 -15712
rect -2737 -15746 -2703 -15712
rect -2669 -15746 -2635 -15712
rect -2601 -15746 -2567 -15712
rect -2533 -15746 -2499 -15712
rect -2465 -15746 -2431 -15712
rect -2397 -15746 -2363 -15712
rect -2329 -15746 -2295 -15712
rect -1787 -15746 -1753 -15712
rect -1719 -15746 -1685 -15712
rect -1651 -15746 -1617 -15712
rect -1583 -15746 -1549 -15712
rect -1515 -15746 -1481 -15712
rect -1447 -15746 -1413 -15712
rect -1379 -15746 -1345 -15712
rect -1311 -15746 -1277 -15712
rect -769 -15746 -735 -15712
rect -701 -15746 -667 -15712
rect -633 -15746 -599 -15712
rect -565 -15746 -531 -15712
rect -497 -15746 -463 -15712
rect -429 -15746 -395 -15712
rect -361 -15746 -327 -15712
rect -293 -15746 -259 -15712
rect 2851 -16090 2885 -16056
rect 2919 -16090 2953 -16056
rect 2987 -16090 3021 -16056
rect 3055 -16090 3089 -16056
rect 3123 -16090 3157 -16056
rect 3191 -16090 3225 -16056
rect 3259 -16090 3293 -16056
rect 3327 -16090 3361 -16056
rect 3869 -16090 3903 -16056
rect 3937 -16090 3971 -16056
rect 4005 -16090 4039 -16056
rect 4073 -16090 4107 -16056
rect 4141 -16090 4175 -16056
rect 4209 -16090 4243 -16056
rect 4277 -16090 4311 -16056
rect 4345 -16090 4379 -16056
rect 4887 -16090 4921 -16056
rect 4955 -16090 4989 -16056
rect 5023 -16090 5057 -16056
rect 5091 -16090 5125 -16056
rect 5159 -16090 5193 -16056
rect 5227 -16090 5261 -16056
rect 5295 -16090 5329 -16056
rect 5363 -16090 5397 -16056
rect 5905 -16090 5939 -16056
rect 5973 -16090 6007 -16056
rect 6041 -16090 6075 -16056
rect 6109 -16090 6143 -16056
rect 6177 -16090 6211 -16056
rect 6245 -16090 6279 -16056
rect 6313 -16090 6347 -16056
rect 6381 -16090 6415 -16056
rect 6923 -16090 6957 -16056
rect 6991 -16090 7025 -16056
rect 7059 -16090 7093 -16056
rect 7127 -16090 7161 -16056
rect 7195 -16090 7229 -16056
rect 7263 -16090 7297 -16056
rect 7331 -16090 7365 -16056
rect 7399 -16090 7433 -16056
rect 7941 -16090 7975 -16056
rect 8009 -16090 8043 -16056
rect 8077 -16090 8111 -16056
rect 8145 -16090 8179 -16056
rect 8213 -16090 8247 -16056
rect 8281 -16090 8315 -16056
rect 8349 -16090 8383 -16056
rect 8417 -16090 8451 -16056
rect 8959 -16090 8993 -16056
rect 9027 -16090 9061 -16056
rect 9095 -16090 9129 -16056
rect 9163 -16090 9197 -16056
rect 9231 -16090 9265 -16056
rect 9299 -16090 9333 -16056
rect 9367 -16090 9401 -16056
rect 9435 -16090 9469 -16056
rect 9977 -16090 10011 -16056
rect 10045 -16090 10079 -16056
rect 10113 -16090 10147 -16056
rect 10181 -16090 10215 -16056
rect 10249 -16090 10283 -16056
rect 10317 -16090 10351 -16056
rect 10385 -16090 10419 -16056
rect 10453 -16090 10487 -16056
rect 10995 -16090 11029 -16056
rect 11063 -16090 11097 -16056
rect 11131 -16090 11165 -16056
rect 11199 -16090 11233 -16056
rect 11267 -16090 11301 -16056
rect 11335 -16090 11369 -16056
rect 11403 -16090 11437 -16056
rect 11471 -16090 11505 -16056
rect 12013 -16090 12047 -16056
rect 12081 -16090 12115 -16056
rect 12149 -16090 12183 -16056
rect 12217 -16090 12251 -16056
rect 12285 -16090 12319 -16056
rect 12353 -16090 12387 -16056
rect 12421 -16090 12455 -16056
rect 12489 -16090 12523 -16056
rect 13031 -16090 13065 -16056
rect 13099 -16090 13133 -16056
rect 13167 -16090 13201 -16056
rect 13235 -16090 13269 -16056
rect 13303 -16090 13337 -16056
rect 13371 -16090 13405 -16056
rect 13439 -16090 13473 -16056
rect 13507 -16090 13541 -16056
rect 14049 -16090 14083 -16056
rect 14117 -16090 14151 -16056
rect 14185 -16090 14219 -16056
rect 14253 -16090 14287 -16056
rect 14321 -16090 14355 -16056
rect 14389 -16090 14423 -16056
rect 14457 -16090 14491 -16056
rect 14525 -16090 14559 -16056
rect 15067 -16090 15101 -16056
rect 15135 -16090 15169 -16056
rect 15203 -16090 15237 -16056
rect 15271 -16090 15305 -16056
rect 15339 -16090 15373 -16056
rect 15407 -16090 15441 -16056
rect 15475 -16090 15509 -16056
rect 15543 -16090 15577 -16056
rect 16085 -16090 16119 -16056
rect 16153 -16090 16187 -16056
rect 16221 -16090 16255 -16056
rect 16289 -16090 16323 -16056
rect 16357 -16090 16391 -16056
rect 16425 -16090 16459 -16056
rect 16493 -16090 16527 -16056
rect 16561 -16090 16595 -16056
rect 17103 -16090 17137 -16056
rect 17171 -16090 17205 -16056
rect 17239 -16090 17273 -16056
rect 17307 -16090 17341 -16056
rect 17375 -16090 17409 -16056
rect 17443 -16090 17477 -16056
rect 17511 -16090 17545 -16056
rect 17579 -16090 17613 -16056
rect 18121 -16090 18155 -16056
rect 18189 -16090 18223 -16056
rect 18257 -16090 18291 -16056
rect 18325 -16090 18359 -16056
rect 18393 -16090 18427 -16056
rect 18461 -16090 18495 -16056
rect 18529 -16090 18563 -16056
rect 18597 -16090 18631 -16056
rect 19139 -16090 19173 -16056
rect 19207 -16090 19241 -16056
rect 19275 -16090 19309 -16056
rect 19343 -16090 19377 -16056
rect 19411 -16090 19445 -16056
rect 19479 -16090 19513 -16056
rect 19547 -16090 19581 -16056
rect 19615 -16090 19649 -16056
rect 20157 -16090 20191 -16056
rect 20225 -16090 20259 -16056
rect 20293 -16090 20327 -16056
rect 20361 -16090 20395 -16056
rect 20429 -16090 20463 -16056
rect 20497 -16090 20531 -16056
rect 20565 -16090 20599 -16056
rect 20633 -16090 20667 -16056
rect 21175 -16090 21209 -16056
rect 21243 -16090 21277 -16056
rect 21311 -16090 21345 -16056
rect 21379 -16090 21413 -16056
rect 21447 -16090 21481 -16056
rect 21515 -16090 21549 -16056
rect 21583 -16090 21617 -16056
rect 21651 -16090 21685 -16056
rect 22193 -16090 22227 -16056
rect 22261 -16090 22295 -16056
rect 22329 -16090 22363 -16056
rect 22397 -16090 22431 -16056
rect 22465 -16090 22499 -16056
rect 22533 -16090 22567 -16056
rect 22601 -16090 22635 -16056
rect 22669 -16090 22703 -16056
rect -8913 -16456 -8879 -16422
rect -8845 -16456 -8811 -16422
rect -8777 -16456 -8743 -16422
rect -8709 -16456 -8675 -16422
rect -8641 -16456 -8607 -16422
rect -8573 -16456 -8539 -16422
rect -8505 -16456 -8471 -16422
rect -8437 -16456 -8403 -16422
rect -7895 -16456 -7861 -16422
rect -7827 -16456 -7793 -16422
rect -7759 -16456 -7725 -16422
rect -7691 -16456 -7657 -16422
rect -7623 -16456 -7589 -16422
rect -7555 -16456 -7521 -16422
rect -7487 -16456 -7453 -16422
rect -7419 -16456 -7385 -16422
rect -6877 -16456 -6843 -16422
rect -6809 -16456 -6775 -16422
rect -6741 -16456 -6707 -16422
rect -6673 -16456 -6639 -16422
rect -6605 -16456 -6571 -16422
rect -6537 -16456 -6503 -16422
rect -6469 -16456 -6435 -16422
rect -6401 -16456 -6367 -16422
rect -5859 -16456 -5825 -16422
rect -5791 -16456 -5757 -16422
rect -5723 -16456 -5689 -16422
rect -5655 -16456 -5621 -16422
rect -5587 -16456 -5553 -16422
rect -5519 -16456 -5485 -16422
rect -5451 -16456 -5417 -16422
rect -5383 -16456 -5349 -16422
rect -4841 -16456 -4807 -16422
rect -4773 -16456 -4739 -16422
rect -4705 -16456 -4671 -16422
rect -4637 -16456 -4603 -16422
rect -4569 -16456 -4535 -16422
rect -4501 -16456 -4467 -16422
rect -4433 -16456 -4399 -16422
rect -4365 -16456 -4331 -16422
rect -3823 -16456 -3789 -16422
rect -3755 -16456 -3721 -16422
rect -3687 -16456 -3653 -16422
rect -3619 -16456 -3585 -16422
rect -3551 -16456 -3517 -16422
rect -3483 -16456 -3449 -16422
rect -3415 -16456 -3381 -16422
rect -3347 -16456 -3313 -16422
rect -2805 -16456 -2771 -16422
rect -2737 -16456 -2703 -16422
rect -2669 -16456 -2635 -16422
rect -2601 -16456 -2567 -16422
rect -2533 -16456 -2499 -16422
rect -2465 -16456 -2431 -16422
rect -2397 -16456 -2363 -16422
rect -2329 -16456 -2295 -16422
rect -1787 -16456 -1753 -16422
rect -1719 -16456 -1685 -16422
rect -1651 -16456 -1617 -16422
rect -1583 -16456 -1549 -16422
rect -1515 -16456 -1481 -16422
rect -1447 -16456 -1413 -16422
rect -1379 -16456 -1345 -16422
rect -1311 -16456 -1277 -16422
rect -769 -16456 -735 -16422
rect -701 -16456 -667 -16422
rect -633 -16456 -599 -16422
rect -565 -16456 -531 -16422
rect -497 -16456 -463 -16422
rect -429 -16456 -395 -16422
rect -361 -16456 -327 -16422
rect -293 -16456 -259 -16422
rect -8913 -16564 -8879 -16530
rect -8845 -16564 -8811 -16530
rect -8777 -16564 -8743 -16530
rect -8709 -16564 -8675 -16530
rect -8641 -16564 -8607 -16530
rect -8573 -16564 -8539 -16530
rect -8505 -16564 -8471 -16530
rect -8437 -16564 -8403 -16530
rect -7895 -16564 -7861 -16530
rect -7827 -16564 -7793 -16530
rect -7759 -16564 -7725 -16530
rect -7691 -16564 -7657 -16530
rect -7623 -16564 -7589 -16530
rect -7555 -16564 -7521 -16530
rect -7487 -16564 -7453 -16530
rect -7419 -16564 -7385 -16530
rect -6877 -16564 -6843 -16530
rect -6809 -16564 -6775 -16530
rect -6741 -16564 -6707 -16530
rect -6673 -16564 -6639 -16530
rect -6605 -16564 -6571 -16530
rect -6537 -16564 -6503 -16530
rect -6469 -16564 -6435 -16530
rect -6401 -16564 -6367 -16530
rect -5859 -16564 -5825 -16530
rect -5791 -16564 -5757 -16530
rect -5723 -16564 -5689 -16530
rect -5655 -16564 -5621 -16530
rect -5587 -16564 -5553 -16530
rect -5519 -16564 -5485 -16530
rect -5451 -16564 -5417 -16530
rect -5383 -16564 -5349 -16530
rect -4841 -16564 -4807 -16530
rect -4773 -16564 -4739 -16530
rect -4705 -16564 -4671 -16530
rect -4637 -16564 -4603 -16530
rect -4569 -16564 -4535 -16530
rect -4501 -16564 -4467 -16530
rect -4433 -16564 -4399 -16530
rect -4365 -16564 -4331 -16530
rect -3823 -16564 -3789 -16530
rect -3755 -16564 -3721 -16530
rect -3687 -16564 -3653 -16530
rect -3619 -16564 -3585 -16530
rect -3551 -16564 -3517 -16530
rect -3483 -16564 -3449 -16530
rect -3415 -16564 -3381 -16530
rect -3347 -16564 -3313 -16530
rect -2805 -16564 -2771 -16530
rect -2737 -16564 -2703 -16530
rect -2669 -16564 -2635 -16530
rect -2601 -16564 -2567 -16530
rect -2533 -16564 -2499 -16530
rect -2465 -16564 -2431 -16530
rect -2397 -16564 -2363 -16530
rect -2329 -16564 -2295 -16530
rect -1787 -16564 -1753 -16530
rect -1719 -16564 -1685 -16530
rect -1651 -16564 -1617 -16530
rect -1583 -16564 -1549 -16530
rect -1515 -16564 -1481 -16530
rect -1447 -16564 -1413 -16530
rect -1379 -16564 -1345 -16530
rect -1311 -16564 -1277 -16530
rect -769 -16564 -735 -16530
rect -701 -16564 -667 -16530
rect -633 -16564 -599 -16530
rect -565 -16564 -531 -16530
rect -497 -16564 -463 -16530
rect -429 -16564 -395 -16530
rect -361 -16564 -327 -16530
rect -293 -16564 -259 -16530
rect 2851 -16614 2885 -16580
rect 2919 -16614 2953 -16580
rect 2987 -16614 3021 -16580
rect 3055 -16614 3089 -16580
rect 3123 -16614 3157 -16580
rect 3191 -16614 3225 -16580
rect 3259 -16614 3293 -16580
rect 3327 -16614 3361 -16580
rect 3869 -16614 3903 -16580
rect 3937 -16614 3971 -16580
rect 4005 -16614 4039 -16580
rect 4073 -16614 4107 -16580
rect 4141 -16614 4175 -16580
rect 4209 -16614 4243 -16580
rect 4277 -16614 4311 -16580
rect 4345 -16614 4379 -16580
rect 4887 -16614 4921 -16580
rect 4955 -16614 4989 -16580
rect 5023 -16614 5057 -16580
rect 5091 -16614 5125 -16580
rect 5159 -16614 5193 -16580
rect 5227 -16614 5261 -16580
rect 5295 -16614 5329 -16580
rect 5363 -16614 5397 -16580
rect 5905 -16614 5939 -16580
rect 5973 -16614 6007 -16580
rect 6041 -16614 6075 -16580
rect 6109 -16614 6143 -16580
rect 6177 -16614 6211 -16580
rect 6245 -16614 6279 -16580
rect 6313 -16614 6347 -16580
rect 6381 -16614 6415 -16580
rect 6923 -16614 6957 -16580
rect 6991 -16614 7025 -16580
rect 7059 -16614 7093 -16580
rect 7127 -16614 7161 -16580
rect 7195 -16614 7229 -16580
rect 7263 -16614 7297 -16580
rect 7331 -16614 7365 -16580
rect 7399 -16614 7433 -16580
rect 7941 -16614 7975 -16580
rect 8009 -16614 8043 -16580
rect 8077 -16614 8111 -16580
rect 8145 -16614 8179 -16580
rect 8213 -16614 8247 -16580
rect 8281 -16614 8315 -16580
rect 8349 -16614 8383 -16580
rect 8417 -16614 8451 -16580
rect 8959 -16614 8993 -16580
rect 9027 -16614 9061 -16580
rect 9095 -16614 9129 -16580
rect 9163 -16614 9197 -16580
rect 9231 -16614 9265 -16580
rect 9299 -16614 9333 -16580
rect 9367 -16614 9401 -16580
rect 9435 -16614 9469 -16580
rect 9977 -16614 10011 -16580
rect 10045 -16614 10079 -16580
rect 10113 -16614 10147 -16580
rect 10181 -16614 10215 -16580
rect 10249 -16614 10283 -16580
rect 10317 -16614 10351 -16580
rect 10385 -16614 10419 -16580
rect 10453 -16614 10487 -16580
rect 10995 -16614 11029 -16580
rect 11063 -16614 11097 -16580
rect 11131 -16614 11165 -16580
rect 11199 -16614 11233 -16580
rect 11267 -16614 11301 -16580
rect 11335 -16614 11369 -16580
rect 11403 -16614 11437 -16580
rect 11471 -16614 11505 -16580
rect 12013 -16614 12047 -16580
rect 12081 -16614 12115 -16580
rect 12149 -16614 12183 -16580
rect 12217 -16614 12251 -16580
rect 12285 -16614 12319 -16580
rect 12353 -16614 12387 -16580
rect 12421 -16614 12455 -16580
rect 12489 -16614 12523 -16580
rect 13031 -16614 13065 -16580
rect 13099 -16614 13133 -16580
rect 13167 -16614 13201 -16580
rect 13235 -16614 13269 -16580
rect 13303 -16614 13337 -16580
rect 13371 -16614 13405 -16580
rect 13439 -16614 13473 -16580
rect 13507 -16614 13541 -16580
rect 14049 -16614 14083 -16580
rect 14117 -16614 14151 -16580
rect 14185 -16614 14219 -16580
rect 14253 -16614 14287 -16580
rect 14321 -16614 14355 -16580
rect 14389 -16614 14423 -16580
rect 14457 -16614 14491 -16580
rect 14525 -16614 14559 -16580
rect 15067 -16614 15101 -16580
rect 15135 -16614 15169 -16580
rect 15203 -16614 15237 -16580
rect 15271 -16614 15305 -16580
rect 15339 -16614 15373 -16580
rect 15407 -16614 15441 -16580
rect 15475 -16614 15509 -16580
rect 15543 -16614 15577 -16580
rect 16085 -16614 16119 -16580
rect 16153 -16614 16187 -16580
rect 16221 -16614 16255 -16580
rect 16289 -16614 16323 -16580
rect 16357 -16614 16391 -16580
rect 16425 -16614 16459 -16580
rect 16493 -16614 16527 -16580
rect 16561 -16614 16595 -16580
rect 17103 -16614 17137 -16580
rect 17171 -16614 17205 -16580
rect 17239 -16614 17273 -16580
rect 17307 -16614 17341 -16580
rect 17375 -16614 17409 -16580
rect 17443 -16614 17477 -16580
rect 17511 -16614 17545 -16580
rect 17579 -16614 17613 -16580
rect 18121 -16614 18155 -16580
rect 18189 -16614 18223 -16580
rect 18257 -16614 18291 -16580
rect 18325 -16614 18359 -16580
rect 18393 -16614 18427 -16580
rect 18461 -16614 18495 -16580
rect 18529 -16614 18563 -16580
rect 18597 -16614 18631 -16580
rect 19139 -16614 19173 -16580
rect 19207 -16614 19241 -16580
rect 19275 -16614 19309 -16580
rect 19343 -16614 19377 -16580
rect 19411 -16614 19445 -16580
rect 19479 -16614 19513 -16580
rect 19547 -16614 19581 -16580
rect 19615 -16614 19649 -16580
rect 20157 -16614 20191 -16580
rect 20225 -16614 20259 -16580
rect 20293 -16614 20327 -16580
rect 20361 -16614 20395 -16580
rect 20429 -16614 20463 -16580
rect 20497 -16614 20531 -16580
rect 20565 -16614 20599 -16580
rect 20633 -16614 20667 -16580
rect 21175 -16614 21209 -16580
rect 21243 -16614 21277 -16580
rect 21311 -16614 21345 -16580
rect 21379 -16614 21413 -16580
rect 21447 -16614 21481 -16580
rect 21515 -16614 21549 -16580
rect 21583 -16614 21617 -16580
rect 21651 -16614 21685 -16580
rect 22193 -16614 22227 -16580
rect 22261 -16614 22295 -16580
rect 22329 -16614 22363 -16580
rect 22397 -16614 22431 -16580
rect 22465 -16614 22499 -16580
rect 22533 -16614 22567 -16580
rect 22601 -16614 22635 -16580
rect 22669 -16614 22703 -16580
rect -8913 -17274 -8879 -17240
rect -8845 -17274 -8811 -17240
rect -8777 -17274 -8743 -17240
rect -8709 -17274 -8675 -17240
rect -8641 -17274 -8607 -17240
rect -8573 -17274 -8539 -17240
rect -8505 -17274 -8471 -17240
rect -8437 -17274 -8403 -17240
rect -7895 -17274 -7861 -17240
rect -7827 -17274 -7793 -17240
rect -7759 -17274 -7725 -17240
rect -7691 -17274 -7657 -17240
rect -7623 -17274 -7589 -17240
rect -7555 -17274 -7521 -17240
rect -7487 -17274 -7453 -17240
rect -7419 -17274 -7385 -17240
rect -6877 -17274 -6843 -17240
rect -6809 -17274 -6775 -17240
rect -6741 -17274 -6707 -17240
rect -6673 -17274 -6639 -17240
rect -6605 -17274 -6571 -17240
rect -6537 -17274 -6503 -17240
rect -6469 -17274 -6435 -17240
rect -6401 -17274 -6367 -17240
rect -5859 -17274 -5825 -17240
rect -5791 -17274 -5757 -17240
rect -5723 -17274 -5689 -17240
rect -5655 -17274 -5621 -17240
rect -5587 -17274 -5553 -17240
rect -5519 -17274 -5485 -17240
rect -5451 -17274 -5417 -17240
rect -5383 -17274 -5349 -17240
rect -4841 -17274 -4807 -17240
rect -4773 -17274 -4739 -17240
rect -4705 -17274 -4671 -17240
rect -4637 -17274 -4603 -17240
rect -4569 -17274 -4535 -17240
rect -4501 -17274 -4467 -17240
rect -4433 -17274 -4399 -17240
rect -4365 -17274 -4331 -17240
rect -3823 -17274 -3789 -17240
rect -3755 -17274 -3721 -17240
rect -3687 -17274 -3653 -17240
rect -3619 -17274 -3585 -17240
rect -3551 -17274 -3517 -17240
rect -3483 -17274 -3449 -17240
rect -3415 -17274 -3381 -17240
rect -3347 -17274 -3313 -17240
rect -2805 -17274 -2771 -17240
rect -2737 -17274 -2703 -17240
rect -2669 -17274 -2635 -17240
rect -2601 -17274 -2567 -17240
rect -2533 -17274 -2499 -17240
rect -2465 -17274 -2431 -17240
rect -2397 -17274 -2363 -17240
rect -2329 -17274 -2295 -17240
rect -1787 -17274 -1753 -17240
rect -1719 -17274 -1685 -17240
rect -1651 -17274 -1617 -17240
rect -1583 -17274 -1549 -17240
rect -1515 -17274 -1481 -17240
rect -1447 -17274 -1413 -17240
rect -1379 -17274 -1345 -17240
rect -1311 -17274 -1277 -17240
rect -769 -17274 -735 -17240
rect -701 -17274 -667 -17240
rect -633 -17274 -599 -17240
rect -565 -17274 -531 -17240
rect -497 -17274 -463 -17240
rect -429 -17274 -395 -17240
rect -361 -17274 -327 -17240
rect -293 -17274 -259 -17240
rect 2851 -17324 2885 -17290
rect 2919 -17324 2953 -17290
rect 2987 -17324 3021 -17290
rect 3055 -17324 3089 -17290
rect 3123 -17324 3157 -17290
rect 3191 -17324 3225 -17290
rect 3259 -17324 3293 -17290
rect 3327 -17324 3361 -17290
rect -8913 -17382 -8879 -17348
rect -8845 -17382 -8811 -17348
rect -8777 -17382 -8743 -17348
rect -8709 -17382 -8675 -17348
rect -8641 -17382 -8607 -17348
rect -8573 -17382 -8539 -17348
rect -8505 -17382 -8471 -17348
rect -8437 -17382 -8403 -17348
rect -7895 -17382 -7861 -17348
rect -7827 -17382 -7793 -17348
rect -7759 -17382 -7725 -17348
rect -7691 -17382 -7657 -17348
rect -7623 -17382 -7589 -17348
rect -7555 -17382 -7521 -17348
rect -7487 -17382 -7453 -17348
rect -7419 -17382 -7385 -17348
rect -6877 -17382 -6843 -17348
rect -6809 -17382 -6775 -17348
rect -6741 -17382 -6707 -17348
rect -6673 -17382 -6639 -17348
rect -6605 -17382 -6571 -17348
rect -6537 -17382 -6503 -17348
rect -6469 -17382 -6435 -17348
rect -6401 -17382 -6367 -17348
rect -5859 -17382 -5825 -17348
rect -5791 -17382 -5757 -17348
rect -5723 -17382 -5689 -17348
rect -5655 -17382 -5621 -17348
rect -5587 -17382 -5553 -17348
rect -5519 -17382 -5485 -17348
rect -5451 -17382 -5417 -17348
rect -5383 -17382 -5349 -17348
rect -4841 -17382 -4807 -17348
rect -4773 -17382 -4739 -17348
rect -4705 -17382 -4671 -17348
rect -4637 -17382 -4603 -17348
rect -4569 -17382 -4535 -17348
rect -4501 -17382 -4467 -17348
rect -4433 -17382 -4399 -17348
rect -4365 -17382 -4331 -17348
rect -3823 -17382 -3789 -17348
rect -3755 -17382 -3721 -17348
rect -3687 -17382 -3653 -17348
rect -3619 -17382 -3585 -17348
rect -3551 -17382 -3517 -17348
rect -3483 -17382 -3449 -17348
rect -3415 -17382 -3381 -17348
rect -3347 -17382 -3313 -17348
rect -2805 -17382 -2771 -17348
rect -2737 -17382 -2703 -17348
rect -2669 -17382 -2635 -17348
rect -2601 -17382 -2567 -17348
rect -2533 -17382 -2499 -17348
rect -2465 -17382 -2431 -17348
rect -2397 -17382 -2363 -17348
rect -2329 -17382 -2295 -17348
rect -1787 -17382 -1753 -17348
rect -1719 -17382 -1685 -17348
rect -1651 -17382 -1617 -17348
rect -1583 -17382 -1549 -17348
rect -1515 -17382 -1481 -17348
rect -1447 -17382 -1413 -17348
rect -1379 -17382 -1345 -17348
rect -1311 -17382 -1277 -17348
rect 3869 -17324 3903 -17290
rect 3937 -17324 3971 -17290
rect 4005 -17324 4039 -17290
rect 4073 -17324 4107 -17290
rect 4141 -17324 4175 -17290
rect 4209 -17324 4243 -17290
rect 4277 -17324 4311 -17290
rect 4345 -17324 4379 -17290
rect 4887 -17324 4921 -17290
rect 4955 -17324 4989 -17290
rect 5023 -17324 5057 -17290
rect 5091 -17324 5125 -17290
rect 5159 -17324 5193 -17290
rect 5227 -17324 5261 -17290
rect 5295 -17324 5329 -17290
rect 5363 -17324 5397 -17290
rect 5905 -17324 5939 -17290
rect 5973 -17324 6007 -17290
rect 6041 -17324 6075 -17290
rect 6109 -17324 6143 -17290
rect 6177 -17324 6211 -17290
rect 6245 -17324 6279 -17290
rect 6313 -17324 6347 -17290
rect 6381 -17324 6415 -17290
rect 6923 -17324 6957 -17290
rect 6991 -17324 7025 -17290
rect 7059 -17324 7093 -17290
rect 7127 -17324 7161 -17290
rect 7195 -17324 7229 -17290
rect 7263 -17324 7297 -17290
rect 7331 -17324 7365 -17290
rect 7399 -17324 7433 -17290
rect 7941 -17324 7975 -17290
rect 8009 -17324 8043 -17290
rect 8077 -17324 8111 -17290
rect 8145 -17324 8179 -17290
rect 8213 -17324 8247 -17290
rect 8281 -17324 8315 -17290
rect 8349 -17324 8383 -17290
rect 8417 -17324 8451 -17290
rect 8959 -17324 8993 -17290
rect 9027 -17324 9061 -17290
rect 9095 -17324 9129 -17290
rect 9163 -17324 9197 -17290
rect 9231 -17324 9265 -17290
rect 9299 -17324 9333 -17290
rect 9367 -17324 9401 -17290
rect 9435 -17324 9469 -17290
rect 9977 -17324 10011 -17290
rect 10045 -17324 10079 -17290
rect 10113 -17324 10147 -17290
rect 10181 -17324 10215 -17290
rect 10249 -17324 10283 -17290
rect 10317 -17324 10351 -17290
rect 10385 -17324 10419 -17290
rect 10453 -17324 10487 -17290
rect 10995 -17324 11029 -17290
rect 11063 -17324 11097 -17290
rect 11131 -17324 11165 -17290
rect 11199 -17324 11233 -17290
rect 11267 -17324 11301 -17290
rect 11335 -17324 11369 -17290
rect 11403 -17324 11437 -17290
rect 11471 -17324 11505 -17290
rect 12013 -17324 12047 -17290
rect 12081 -17324 12115 -17290
rect 12149 -17324 12183 -17290
rect 12217 -17324 12251 -17290
rect 12285 -17324 12319 -17290
rect 12353 -17324 12387 -17290
rect 12421 -17324 12455 -17290
rect 12489 -17324 12523 -17290
rect 13031 -17324 13065 -17290
rect 13099 -17324 13133 -17290
rect 13167 -17324 13201 -17290
rect 13235 -17324 13269 -17290
rect 13303 -17324 13337 -17290
rect 13371 -17324 13405 -17290
rect 13439 -17324 13473 -17290
rect 13507 -17324 13541 -17290
rect 14049 -17324 14083 -17290
rect 14117 -17324 14151 -17290
rect 14185 -17324 14219 -17290
rect 14253 -17324 14287 -17290
rect 14321 -17324 14355 -17290
rect 14389 -17324 14423 -17290
rect 14457 -17324 14491 -17290
rect 14525 -17324 14559 -17290
rect 15067 -17324 15101 -17290
rect 15135 -17324 15169 -17290
rect 15203 -17324 15237 -17290
rect 15271 -17324 15305 -17290
rect 15339 -17324 15373 -17290
rect 15407 -17324 15441 -17290
rect 15475 -17324 15509 -17290
rect 15543 -17324 15577 -17290
rect 16085 -17324 16119 -17290
rect 16153 -17324 16187 -17290
rect 16221 -17324 16255 -17290
rect 16289 -17324 16323 -17290
rect 16357 -17324 16391 -17290
rect 16425 -17324 16459 -17290
rect 16493 -17324 16527 -17290
rect 16561 -17324 16595 -17290
rect 17103 -17324 17137 -17290
rect 17171 -17324 17205 -17290
rect 17239 -17324 17273 -17290
rect 17307 -17324 17341 -17290
rect 17375 -17324 17409 -17290
rect 17443 -17324 17477 -17290
rect 17511 -17324 17545 -17290
rect 17579 -17324 17613 -17290
rect 18121 -17324 18155 -17290
rect 18189 -17324 18223 -17290
rect 18257 -17324 18291 -17290
rect 18325 -17324 18359 -17290
rect 18393 -17324 18427 -17290
rect 18461 -17324 18495 -17290
rect 18529 -17324 18563 -17290
rect 18597 -17324 18631 -17290
rect 19139 -17324 19173 -17290
rect 19207 -17324 19241 -17290
rect 19275 -17324 19309 -17290
rect 19343 -17324 19377 -17290
rect 19411 -17324 19445 -17290
rect 19479 -17324 19513 -17290
rect 19547 -17324 19581 -17290
rect 19615 -17324 19649 -17290
rect 20157 -17324 20191 -17290
rect 20225 -17324 20259 -17290
rect 20293 -17324 20327 -17290
rect 20361 -17324 20395 -17290
rect 20429 -17324 20463 -17290
rect 20497 -17324 20531 -17290
rect 20565 -17324 20599 -17290
rect 20633 -17324 20667 -17290
rect 21175 -17324 21209 -17290
rect 21243 -17324 21277 -17290
rect 21311 -17324 21345 -17290
rect 21379 -17324 21413 -17290
rect 21447 -17324 21481 -17290
rect 21515 -17324 21549 -17290
rect 21583 -17324 21617 -17290
rect 21651 -17324 21685 -17290
rect 22193 -17324 22227 -17290
rect 22261 -17324 22295 -17290
rect 22329 -17324 22363 -17290
rect 22397 -17324 22431 -17290
rect 22465 -17324 22499 -17290
rect 22533 -17324 22567 -17290
rect 22601 -17324 22635 -17290
rect 22669 -17324 22703 -17290
rect -769 -17382 -735 -17348
rect -701 -17382 -667 -17348
rect -633 -17382 -599 -17348
rect -565 -17382 -531 -17348
rect -497 -17382 -463 -17348
rect -429 -17382 -395 -17348
rect -361 -17382 -327 -17348
rect -293 -17382 -259 -17348
rect 2851 -17846 2885 -17812
rect 2919 -17846 2953 -17812
rect 2987 -17846 3021 -17812
rect 3055 -17846 3089 -17812
rect 3123 -17846 3157 -17812
rect 3191 -17846 3225 -17812
rect 3259 -17846 3293 -17812
rect 3327 -17846 3361 -17812
rect 3869 -17846 3903 -17812
rect 3937 -17846 3971 -17812
rect 4005 -17846 4039 -17812
rect 4073 -17846 4107 -17812
rect 4141 -17846 4175 -17812
rect 4209 -17846 4243 -17812
rect 4277 -17846 4311 -17812
rect 4345 -17846 4379 -17812
rect 4887 -17846 4921 -17812
rect 4955 -17846 4989 -17812
rect 5023 -17846 5057 -17812
rect 5091 -17846 5125 -17812
rect 5159 -17846 5193 -17812
rect 5227 -17846 5261 -17812
rect 5295 -17846 5329 -17812
rect 5363 -17846 5397 -17812
rect 5905 -17846 5939 -17812
rect 5973 -17846 6007 -17812
rect 6041 -17846 6075 -17812
rect 6109 -17846 6143 -17812
rect 6177 -17846 6211 -17812
rect 6245 -17846 6279 -17812
rect 6313 -17846 6347 -17812
rect 6381 -17846 6415 -17812
rect 6923 -17846 6957 -17812
rect 6991 -17846 7025 -17812
rect 7059 -17846 7093 -17812
rect 7127 -17846 7161 -17812
rect 7195 -17846 7229 -17812
rect 7263 -17846 7297 -17812
rect 7331 -17846 7365 -17812
rect 7399 -17846 7433 -17812
rect 7941 -17846 7975 -17812
rect 8009 -17846 8043 -17812
rect 8077 -17846 8111 -17812
rect 8145 -17846 8179 -17812
rect 8213 -17846 8247 -17812
rect 8281 -17846 8315 -17812
rect 8349 -17846 8383 -17812
rect 8417 -17846 8451 -17812
rect 8959 -17846 8993 -17812
rect 9027 -17846 9061 -17812
rect 9095 -17846 9129 -17812
rect 9163 -17846 9197 -17812
rect 9231 -17846 9265 -17812
rect 9299 -17846 9333 -17812
rect 9367 -17846 9401 -17812
rect 9435 -17846 9469 -17812
rect 9977 -17846 10011 -17812
rect 10045 -17846 10079 -17812
rect 10113 -17846 10147 -17812
rect 10181 -17846 10215 -17812
rect 10249 -17846 10283 -17812
rect 10317 -17846 10351 -17812
rect 10385 -17846 10419 -17812
rect 10453 -17846 10487 -17812
rect 10995 -17846 11029 -17812
rect 11063 -17846 11097 -17812
rect 11131 -17846 11165 -17812
rect 11199 -17846 11233 -17812
rect 11267 -17846 11301 -17812
rect 11335 -17846 11369 -17812
rect 11403 -17846 11437 -17812
rect 11471 -17846 11505 -17812
rect 12013 -17846 12047 -17812
rect 12081 -17846 12115 -17812
rect 12149 -17846 12183 -17812
rect 12217 -17846 12251 -17812
rect 12285 -17846 12319 -17812
rect 12353 -17846 12387 -17812
rect 12421 -17846 12455 -17812
rect 12489 -17846 12523 -17812
rect 13031 -17846 13065 -17812
rect 13099 -17846 13133 -17812
rect 13167 -17846 13201 -17812
rect 13235 -17846 13269 -17812
rect 13303 -17846 13337 -17812
rect 13371 -17846 13405 -17812
rect 13439 -17846 13473 -17812
rect 13507 -17846 13541 -17812
rect 14049 -17846 14083 -17812
rect 14117 -17846 14151 -17812
rect 14185 -17846 14219 -17812
rect 14253 -17846 14287 -17812
rect 14321 -17846 14355 -17812
rect 14389 -17846 14423 -17812
rect 14457 -17846 14491 -17812
rect 14525 -17846 14559 -17812
rect 15067 -17846 15101 -17812
rect 15135 -17846 15169 -17812
rect 15203 -17846 15237 -17812
rect 15271 -17846 15305 -17812
rect 15339 -17846 15373 -17812
rect 15407 -17846 15441 -17812
rect 15475 -17846 15509 -17812
rect 15543 -17846 15577 -17812
rect 16085 -17846 16119 -17812
rect 16153 -17846 16187 -17812
rect 16221 -17846 16255 -17812
rect 16289 -17846 16323 -17812
rect 16357 -17846 16391 -17812
rect 16425 -17846 16459 -17812
rect 16493 -17846 16527 -17812
rect 16561 -17846 16595 -17812
rect 17103 -17846 17137 -17812
rect 17171 -17846 17205 -17812
rect 17239 -17846 17273 -17812
rect 17307 -17846 17341 -17812
rect 17375 -17846 17409 -17812
rect 17443 -17846 17477 -17812
rect 17511 -17846 17545 -17812
rect 17579 -17846 17613 -17812
rect 18121 -17846 18155 -17812
rect 18189 -17846 18223 -17812
rect 18257 -17846 18291 -17812
rect 18325 -17846 18359 -17812
rect 18393 -17846 18427 -17812
rect 18461 -17846 18495 -17812
rect 18529 -17846 18563 -17812
rect 18597 -17846 18631 -17812
rect 19139 -17846 19173 -17812
rect 19207 -17846 19241 -17812
rect 19275 -17846 19309 -17812
rect 19343 -17846 19377 -17812
rect 19411 -17846 19445 -17812
rect 19479 -17846 19513 -17812
rect 19547 -17846 19581 -17812
rect 19615 -17846 19649 -17812
rect 20157 -17846 20191 -17812
rect 20225 -17846 20259 -17812
rect 20293 -17846 20327 -17812
rect 20361 -17846 20395 -17812
rect 20429 -17846 20463 -17812
rect 20497 -17846 20531 -17812
rect 20565 -17846 20599 -17812
rect 20633 -17846 20667 -17812
rect 21175 -17846 21209 -17812
rect 21243 -17846 21277 -17812
rect 21311 -17846 21345 -17812
rect 21379 -17846 21413 -17812
rect 21447 -17846 21481 -17812
rect 21515 -17846 21549 -17812
rect 21583 -17846 21617 -17812
rect 21651 -17846 21685 -17812
rect 22193 -17846 22227 -17812
rect 22261 -17846 22295 -17812
rect 22329 -17846 22363 -17812
rect 22397 -17846 22431 -17812
rect 22465 -17846 22499 -17812
rect 22533 -17846 22567 -17812
rect 22601 -17846 22635 -17812
rect 22669 -17846 22703 -17812
rect -8913 -18092 -8879 -18058
rect -8845 -18092 -8811 -18058
rect -8777 -18092 -8743 -18058
rect -8709 -18092 -8675 -18058
rect -8641 -18092 -8607 -18058
rect -8573 -18092 -8539 -18058
rect -8505 -18092 -8471 -18058
rect -8437 -18092 -8403 -18058
rect -7895 -18092 -7861 -18058
rect -7827 -18092 -7793 -18058
rect -7759 -18092 -7725 -18058
rect -7691 -18092 -7657 -18058
rect -7623 -18092 -7589 -18058
rect -7555 -18092 -7521 -18058
rect -7487 -18092 -7453 -18058
rect -7419 -18092 -7385 -18058
rect -6877 -18092 -6843 -18058
rect -6809 -18092 -6775 -18058
rect -6741 -18092 -6707 -18058
rect -6673 -18092 -6639 -18058
rect -6605 -18092 -6571 -18058
rect -6537 -18092 -6503 -18058
rect -6469 -18092 -6435 -18058
rect -6401 -18092 -6367 -18058
rect -5859 -18092 -5825 -18058
rect -5791 -18092 -5757 -18058
rect -5723 -18092 -5689 -18058
rect -5655 -18092 -5621 -18058
rect -5587 -18092 -5553 -18058
rect -5519 -18092 -5485 -18058
rect -5451 -18092 -5417 -18058
rect -5383 -18092 -5349 -18058
rect -4841 -18092 -4807 -18058
rect -4773 -18092 -4739 -18058
rect -4705 -18092 -4671 -18058
rect -4637 -18092 -4603 -18058
rect -4569 -18092 -4535 -18058
rect -4501 -18092 -4467 -18058
rect -4433 -18092 -4399 -18058
rect -4365 -18092 -4331 -18058
rect -3823 -18092 -3789 -18058
rect -3755 -18092 -3721 -18058
rect -3687 -18092 -3653 -18058
rect -3619 -18092 -3585 -18058
rect -3551 -18092 -3517 -18058
rect -3483 -18092 -3449 -18058
rect -3415 -18092 -3381 -18058
rect -3347 -18092 -3313 -18058
rect -2805 -18092 -2771 -18058
rect -2737 -18092 -2703 -18058
rect -2669 -18092 -2635 -18058
rect -2601 -18092 -2567 -18058
rect -2533 -18092 -2499 -18058
rect -2465 -18092 -2431 -18058
rect -2397 -18092 -2363 -18058
rect -2329 -18092 -2295 -18058
rect -1787 -18092 -1753 -18058
rect -1719 -18092 -1685 -18058
rect -1651 -18092 -1617 -18058
rect -1583 -18092 -1549 -18058
rect -1515 -18092 -1481 -18058
rect -1447 -18092 -1413 -18058
rect -1379 -18092 -1345 -18058
rect -1311 -18092 -1277 -18058
rect -769 -18092 -735 -18058
rect -701 -18092 -667 -18058
rect -633 -18092 -599 -18058
rect -565 -18092 -531 -18058
rect -497 -18092 -463 -18058
rect -429 -18092 -395 -18058
rect -361 -18092 -327 -18058
rect -293 -18092 -259 -18058
rect -8913 -18200 -8879 -18166
rect -8845 -18200 -8811 -18166
rect -8777 -18200 -8743 -18166
rect -8709 -18200 -8675 -18166
rect -8641 -18200 -8607 -18166
rect -8573 -18200 -8539 -18166
rect -8505 -18200 -8471 -18166
rect -8437 -18200 -8403 -18166
rect -7895 -18200 -7861 -18166
rect -7827 -18200 -7793 -18166
rect -7759 -18200 -7725 -18166
rect -7691 -18200 -7657 -18166
rect -7623 -18200 -7589 -18166
rect -7555 -18200 -7521 -18166
rect -7487 -18200 -7453 -18166
rect -7419 -18200 -7385 -18166
rect -6877 -18200 -6843 -18166
rect -6809 -18200 -6775 -18166
rect -6741 -18200 -6707 -18166
rect -6673 -18200 -6639 -18166
rect -6605 -18200 -6571 -18166
rect -6537 -18200 -6503 -18166
rect -6469 -18200 -6435 -18166
rect -6401 -18200 -6367 -18166
rect -5859 -18200 -5825 -18166
rect -5791 -18200 -5757 -18166
rect -5723 -18200 -5689 -18166
rect -5655 -18200 -5621 -18166
rect -5587 -18200 -5553 -18166
rect -5519 -18200 -5485 -18166
rect -5451 -18200 -5417 -18166
rect -5383 -18200 -5349 -18166
rect -4841 -18200 -4807 -18166
rect -4773 -18200 -4739 -18166
rect -4705 -18200 -4671 -18166
rect -4637 -18200 -4603 -18166
rect -4569 -18200 -4535 -18166
rect -4501 -18200 -4467 -18166
rect -4433 -18200 -4399 -18166
rect -4365 -18200 -4331 -18166
rect -3823 -18200 -3789 -18166
rect -3755 -18200 -3721 -18166
rect -3687 -18200 -3653 -18166
rect -3619 -18200 -3585 -18166
rect -3551 -18200 -3517 -18166
rect -3483 -18200 -3449 -18166
rect -3415 -18200 -3381 -18166
rect -3347 -18200 -3313 -18166
rect -2805 -18200 -2771 -18166
rect -2737 -18200 -2703 -18166
rect -2669 -18200 -2635 -18166
rect -2601 -18200 -2567 -18166
rect -2533 -18200 -2499 -18166
rect -2465 -18200 -2431 -18166
rect -2397 -18200 -2363 -18166
rect -2329 -18200 -2295 -18166
rect -1787 -18200 -1753 -18166
rect -1719 -18200 -1685 -18166
rect -1651 -18200 -1617 -18166
rect -1583 -18200 -1549 -18166
rect -1515 -18200 -1481 -18166
rect -1447 -18200 -1413 -18166
rect -1379 -18200 -1345 -18166
rect -1311 -18200 -1277 -18166
rect -769 -18200 -735 -18166
rect -701 -18200 -667 -18166
rect -633 -18200 -599 -18166
rect -565 -18200 -531 -18166
rect -497 -18200 -463 -18166
rect -429 -18200 -395 -18166
rect -361 -18200 -327 -18166
rect -293 -18200 -259 -18166
rect 2851 -18556 2885 -18522
rect 2919 -18556 2953 -18522
rect 2987 -18556 3021 -18522
rect 3055 -18556 3089 -18522
rect 3123 -18556 3157 -18522
rect 3191 -18556 3225 -18522
rect 3259 -18556 3293 -18522
rect 3327 -18556 3361 -18522
rect 3869 -18556 3903 -18522
rect 3937 -18556 3971 -18522
rect 4005 -18556 4039 -18522
rect 4073 -18556 4107 -18522
rect 4141 -18556 4175 -18522
rect 4209 -18556 4243 -18522
rect 4277 -18556 4311 -18522
rect 4345 -18556 4379 -18522
rect 4887 -18556 4921 -18522
rect 4955 -18556 4989 -18522
rect 5023 -18556 5057 -18522
rect 5091 -18556 5125 -18522
rect 5159 -18556 5193 -18522
rect 5227 -18556 5261 -18522
rect 5295 -18556 5329 -18522
rect 5363 -18556 5397 -18522
rect 5905 -18556 5939 -18522
rect 5973 -18556 6007 -18522
rect 6041 -18556 6075 -18522
rect 6109 -18556 6143 -18522
rect 6177 -18556 6211 -18522
rect 6245 -18556 6279 -18522
rect 6313 -18556 6347 -18522
rect 6381 -18556 6415 -18522
rect 6923 -18556 6957 -18522
rect 6991 -18556 7025 -18522
rect 7059 -18556 7093 -18522
rect 7127 -18556 7161 -18522
rect 7195 -18556 7229 -18522
rect 7263 -18556 7297 -18522
rect 7331 -18556 7365 -18522
rect 7399 -18556 7433 -18522
rect 7941 -18556 7975 -18522
rect 8009 -18556 8043 -18522
rect 8077 -18556 8111 -18522
rect 8145 -18556 8179 -18522
rect 8213 -18556 8247 -18522
rect 8281 -18556 8315 -18522
rect 8349 -18556 8383 -18522
rect 8417 -18556 8451 -18522
rect 8959 -18556 8993 -18522
rect 9027 -18556 9061 -18522
rect 9095 -18556 9129 -18522
rect 9163 -18556 9197 -18522
rect 9231 -18556 9265 -18522
rect 9299 -18556 9333 -18522
rect 9367 -18556 9401 -18522
rect 9435 -18556 9469 -18522
rect 9977 -18556 10011 -18522
rect 10045 -18556 10079 -18522
rect 10113 -18556 10147 -18522
rect 10181 -18556 10215 -18522
rect 10249 -18556 10283 -18522
rect 10317 -18556 10351 -18522
rect 10385 -18556 10419 -18522
rect 10453 -18556 10487 -18522
rect 10995 -18556 11029 -18522
rect 11063 -18556 11097 -18522
rect 11131 -18556 11165 -18522
rect 11199 -18556 11233 -18522
rect 11267 -18556 11301 -18522
rect 11335 -18556 11369 -18522
rect 11403 -18556 11437 -18522
rect 11471 -18556 11505 -18522
rect 12013 -18556 12047 -18522
rect 12081 -18556 12115 -18522
rect 12149 -18556 12183 -18522
rect 12217 -18556 12251 -18522
rect 12285 -18556 12319 -18522
rect 12353 -18556 12387 -18522
rect 12421 -18556 12455 -18522
rect 12489 -18556 12523 -18522
rect 13031 -18556 13065 -18522
rect 13099 -18556 13133 -18522
rect 13167 -18556 13201 -18522
rect 13235 -18556 13269 -18522
rect 13303 -18556 13337 -18522
rect 13371 -18556 13405 -18522
rect 13439 -18556 13473 -18522
rect 13507 -18556 13541 -18522
rect 14049 -18556 14083 -18522
rect 14117 -18556 14151 -18522
rect 14185 -18556 14219 -18522
rect 14253 -18556 14287 -18522
rect 14321 -18556 14355 -18522
rect 14389 -18556 14423 -18522
rect 14457 -18556 14491 -18522
rect 14525 -18556 14559 -18522
rect 15067 -18556 15101 -18522
rect 15135 -18556 15169 -18522
rect 15203 -18556 15237 -18522
rect 15271 -18556 15305 -18522
rect 15339 -18556 15373 -18522
rect 15407 -18556 15441 -18522
rect 15475 -18556 15509 -18522
rect 15543 -18556 15577 -18522
rect 16085 -18556 16119 -18522
rect 16153 -18556 16187 -18522
rect 16221 -18556 16255 -18522
rect 16289 -18556 16323 -18522
rect 16357 -18556 16391 -18522
rect 16425 -18556 16459 -18522
rect 16493 -18556 16527 -18522
rect 16561 -18556 16595 -18522
rect 17103 -18556 17137 -18522
rect 17171 -18556 17205 -18522
rect 17239 -18556 17273 -18522
rect 17307 -18556 17341 -18522
rect 17375 -18556 17409 -18522
rect 17443 -18556 17477 -18522
rect 17511 -18556 17545 -18522
rect 17579 -18556 17613 -18522
rect 18121 -18556 18155 -18522
rect 18189 -18556 18223 -18522
rect 18257 -18556 18291 -18522
rect 18325 -18556 18359 -18522
rect 18393 -18556 18427 -18522
rect 18461 -18556 18495 -18522
rect 18529 -18556 18563 -18522
rect 18597 -18556 18631 -18522
rect 19139 -18556 19173 -18522
rect 19207 -18556 19241 -18522
rect 19275 -18556 19309 -18522
rect 19343 -18556 19377 -18522
rect 19411 -18556 19445 -18522
rect 19479 -18556 19513 -18522
rect 19547 -18556 19581 -18522
rect 19615 -18556 19649 -18522
rect 20157 -18556 20191 -18522
rect 20225 -18556 20259 -18522
rect 20293 -18556 20327 -18522
rect 20361 -18556 20395 -18522
rect 20429 -18556 20463 -18522
rect 20497 -18556 20531 -18522
rect 20565 -18556 20599 -18522
rect 20633 -18556 20667 -18522
rect 21175 -18556 21209 -18522
rect 21243 -18556 21277 -18522
rect 21311 -18556 21345 -18522
rect 21379 -18556 21413 -18522
rect 21447 -18556 21481 -18522
rect 21515 -18556 21549 -18522
rect 21583 -18556 21617 -18522
rect 21651 -18556 21685 -18522
rect 22193 -18556 22227 -18522
rect 22261 -18556 22295 -18522
rect 22329 -18556 22363 -18522
rect 22397 -18556 22431 -18522
rect 22465 -18556 22499 -18522
rect 22533 -18556 22567 -18522
rect 22601 -18556 22635 -18522
rect 22669 -18556 22703 -18522
rect -8913 -18910 -8879 -18876
rect -8845 -18910 -8811 -18876
rect -8777 -18910 -8743 -18876
rect -8709 -18910 -8675 -18876
rect -8641 -18910 -8607 -18876
rect -8573 -18910 -8539 -18876
rect -8505 -18910 -8471 -18876
rect -8437 -18910 -8403 -18876
rect -7895 -18910 -7861 -18876
rect -7827 -18910 -7793 -18876
rect -7759 -18910 -7725 -18876
rect -7691 -18910 -7657 -18876
rect -7623 -18910 -7589 -18876
rect -7555 -18910 -7521 -18876
rect -7487 -18910 -7453 -18876
rect -7419 -18910 -7385 -18876
rect -6877 -18910 -6843 -18876
rect -6809 -18910 -6775 -18876
rect -6741 -18910 -6707 -18876
rect -6673 -18910 -6639 -18876
rect -6605 -18910 -6571 -18876
rect -6537 -18910 -6503 -18876
rect -6469 -18910 -6435 -18876
rect -6401 -18910 -6367 -18876
rect -5859 -18910 -5825 -18876
rect -5791 -18910 -5757 -18876
rect -5723 -18910 -5689 -18876
rect -5655 -18910 -5621 -18876
rect -5587 -18910 -5553 -18876
rect -5519 -18910 -5485 -18876
rect -5451 -18910 -5417 -18876
rect -5383 -18910 -5349 -18876
rect -4841 -18910 -4807 -18876
rect -4773 -18910 -4739 -18876
rect -4705 -18910 -4671 -18876
rect -4637 -18910 -4603 -18876
rect -4569 -18910 -4535 -18876
rect -4501 -18910 -4467 -18876
rect -4433 -18910 -4399 -18876
rect -4365 -18910 -4331 -18876
rect -3823 -18910 -3789 -18876
rect -3755 -18910 -3721 -18876
rect -3687 -18910 -3653 -18876
rect -3619 -18910 -3585 -18876
rect -3551 -18910 -3517 -18876
rect -3483 -18910 -3449 -18876
rect -3415 -18910 -3381 -18876
rect -3347 -18910 -3313 -18876
rect -2805 -18910 -2771 -18876
rect -2737 -18910 -2703 -18876
rect -2669 -18910 -2635 -18876
rect -2601 -18910 -2567 -18876
rect -2533 -18910 -2499 -18876
rect -2465 -18910 -2431 -18876
rect -2397 -18910 -2363 -18876
rect -2329 -18910 -2295 -18876
rect -1787 -18910 -1753 -18876
rect -1719 -18910 -1685 -18876
rect -1651 -18910 -1617 -18876
rect -1583 -18910 -1549 -18876
rect -1515 -18910 -1481 -18876
rect -1447 -18910 -1413 -18876
rect -1379 -18910 -1345 -18876
rect -1311 -18910 -1277 -18876
rect -769 -18910 -735 -18876
rect -701 -18910 -667 -18876
rect -633 -18910 -599 -18876
rect -565 -18910 -531 -18876
rect -497 -18910 -463 -18876
rect -429 -18910 -395 -18876
rect -361 -18910 -327 -18876
rect -293 -18910 -259 -18876
rect 2851 -19080 2885 -19046
rect 2919 -19080 2953 -19046
rect 2987 -19080 3021 -19046
rect 3055 -19080 3089 -19046
rect 3123 -19080 3157 -19046
rect 3191 -19080 3225 -19046
rect 3259 -19080 3293 -19046
rect 3327 -19080 3361 -19046
rect 3869 -19080 3903 -19046
rect 3937 -19080 3971 -19046
rect 4005 -19080 4039 -19046
rect 4073 -19080 4107 -19046
rect 4141 -19080 4175 -19046
rect 4209 -19080 4243 -19046
rect 4277 -19080 4311 -19046
rect 4345 -19080 4379 -19046
rect 4887 -19080 4921 -19046
rect 4955 -19080 4989 -19046
rect 5023 -19080 5057 -19046
rect 5091 -19080 5125 -19046
rect 5159 -19080 5193 -19046
rect 5227 -19080 5261 -19046
rect 5295 -19080 5329 -19046
rect 5363 -19080 5397 -19046
rect 5905 -19080 5939 -19046
rect 5973 -19080 6007 -19046
rect 6041 -19080 6075 -19046
rect 6109 -19080 6143 -19046
rect 6177 -19080 6211 -19046
rect 6245 -19080 6279 -19046
rect 6313 -19080 6347 -19046
rect 6381 -19080 6415 -19046
rect 6923 -19080 6957 -19046
rect 6991 -19080 7025 -19046
rect 7059 -19080 7093 -19046
rect 7127 -19080 7161 -19046
rect 7195 -19080 7229 -19046
rect 7263 -19080 7297 -19046
rect 7331 -19080 7365 -19046
rect 7399 -19080 7433 -19046
rect 7941 -19080 7975 -19046
rect 8009 -19080 8043 -19046
rect 8077 -19080 8111 -19046
rect 8145 -19080 8179 -19046
rect 8213 -19080 8247 -19046
rect 8281 -19080 8315 -19046
rect 8349 -19080 8383 -19046
rect 8417 -19080 8451 -19046
rect 8959 -19080 8993 -19046
rect 9027 -19080 9061 -19046
rect 9095 -19080 9129 -19046
rect 9163 -19080 9197 -19046
rect 9231 -19080 9265 -19046
rect 9299 -19080 9333 -19046
rect 9367 -19080 9401 -19046
rect 9435 -19080 9469 -19046
rect 9977 -19080 10011 -19046
rect 10045 -19080 10079 -19046
rect 10113 -19080 10147 -19046
rect 10181 -19080 10215 -19046
rect 10249 -19080 10283 -19046
rect 10317 -19080 10351 -19046
rect 10385 -19080 10419 -19046
rect 10453 -19080 10487 -19046
rect 10995 -19080 11029 -19046
rect 11063 -19080 11097 -19046
rect 11131 -19080 11165 -19046
rect 11199 -19080 11233 -19046
rect 11267 -19080 11301 -19046
rect 11335 -19080 11369 -19046
rect 11403 -19080 11437 -19046
rect 11471 -19080 11505 -19046
rect 12013 -19080 12047 -19046
rect 12081 -19080 12115 -19046
rect 12149 -19080 12183 -19046
rect 12217 -19080 12251 -19046
rect 12285 -19080 12319 -19046
rect 12353 -19080 12387 -19046
rect 12421 -19080 12455 -19046
rect 12489 -19080 12523 -19046
rect 13031 -19080 13065 -19046
rect 13099 -19080 13133 -19046
rect 13167 -19080 13201 -19046
rect 13235 -19080 13269 -19046
rect 13303 -19080 13337 -19046
rect 13371 -19080 13405 -19046
rect 13439 -19080 13473 -19046
rect 13507 -19080 13541 -19046
rect 14049 -19080 14083 -19046
rect 14117 -19080 14151 -19046
rect 14185 -19080 14219 -19046
rect 14253 -19080 14287 -19046
rect 14321 -19080 14355 -19046
rect 14389 -19080 14423 -19046
rect 14457 -19080 14491 -19046
rect 14525 -19080 14559 -19046
rect 15067 -19080 15101 -19046
rect 15135 -19080 15169 -19046
rect 15203 -19080 15237 -19046
rect 15271 -19080 15305 -19046
rect 15339 -19080 15373 -19046
rect 15407 -19080 15441 -19046
rect 15475 -19080 15509 -19046
rect 15543 -19080 15577 -19046
rect 16085 -19080 16119 -19046
rect 16153 -19080 16187 -19046
rect 16221 -19080 16255 -19046
rect 16289 -19080 16323 -19046
rect 16357 -19080 16391 -19046
rect 16425 -19080 16459 -19046
rect 16493 -19080 16527 -19046
rect 16561 -19080 16595 -19046
rect 17103 -19080 17137 -19046
rect 17171 -19080 17205 -19046
rect 17239 -19080 17273 -19046
rect 17307 -19080 17341 -19046
rect 17375 -19080 17409 -19046
rect 17443 -19080 17477 -19046
rect 17511 -19080 17545 -19046
rect 17579 -19080 17613 -19046
rect 18121 -19080 18155 -19046
rect 18189 -19080 18223 -19046
rect 18257 -19080 18291 -19046
rect 18325 -19080 18359 -19046
rect 18393 -19080 18427 -19046
rect 18461 -19080 18495 -19046
rect 18529 -19080 18563 -19046
rect 18597 -19080 18631 -19046
rect 19139 -19080 19173 -19046
rect 19207 -19080 19241 -19046
rect 19275 -19080 19309 -19046
rect 19343 -19080 19377 -19046
rect 19411 -19080 19445 -19046
rect 19479 -19080 19513 -19046
rect 19547 -19080 19581 -19046
rect 19615 -19080 19649 -19046
rect 20157 -19080 20191 -19046
rect 20225 -19080 20259 -19046
rect 20293 -19080 20327 -19046
rect 20361 -19080 20395 -19046
rect 20429 -19080 20463 -19046
rect 20497 -19080 20531 -19046
rect 20565 -19080 20599 -19046
rect 20633 -19080 20667 -19046
rect 21175 -19080 21209 -19046
rect 21243 -19080 21277 -19046
rect 21311 -19080 21345 -19046
rect 21379 -19080 21413 -19046
rect 21447 -19080 21481 -19046
rect 21515 -19080 21549 -19046
rect 21583 -19080 21617 -19046
rect 21651 -19080 21685 -19046
rect 22193 -19080 22227 -19046
rect 22261 -19080 22295 -19046
rect 22329 -19080 22363 -19046
rect 22397 -19080 22431 -19046
rect 22465 -19080 22499 -19046
rect 22533 -19080 22567 -19046
rect 22601 -19080 22635 -19046
rect 22669 -19080 22703 -19046
rect -2215 -19584 -2181 -19550
rect -1997 -19584 -1963 -19550
rect -1779 -19584 -1745 -19550
rect -1561 -19584 -1527 -19550
rect -1343 -19584 -1309 -19550
rect -1125 -19584 -1091 -19550
rect -907 -19584 -873 -19550
rect -689 -19584 -655 -19550
rect -471 -19584 -437 -19550
rect -253 -19584 -219 -19550
rect 2851 -19790 2885 -19756
rect 2919 -19790 2953 -19756
rect 2987 -19790 3021 -19756
rect 3055 -19790 3089 -19756
rect 3123 -19790 3157 -19756
rect 3191 -19790 3225 -19756
rect 3259 -19790 3293 -19756
rect 3327 -19790 3361 -19756
rect 3869 -19790 3903 -19756
rect 3937 -19790 3971 -19756
rect 4005 -19790 4039 -19756
rect 4073 -19790 4107 -19756
rect 4141 -19790 4175 -19756
rect 4209 -19790 4243 -19756
rect 4277 -19790 4311 -19756
rect 4345 -19790 4379 -19756
rect 4887 -19790 4921 -19756
rect 4955 -19790 4989 -19756
rect 5023 -19790 5057 -19756
rect 5091 -19790 5125 -19756
rect 5159 -19790 5193 -19756
rect 5227 -19790 5261 -19756
rect 5295 -19790 5329 -19756
rect 5363 -19790 5397 -19756
rect 5905 -19790 5939 -19756
rect 5973 -19790 6007 -19756
rect 6041 -19790 6075 -19756
rect 6109 -19790 6143 -19756
rect 6177 -19790 6211 -19756
rect 6245 -19790 6279 -19756
rect 6313 -19790 6347 -19756
rect 6381 -19790 6415 -19756
rect 6923 -19790 6957 -19756
rect 6991 -19790 7025 -19756
rect 7059 -19790 7093 -19756
rect 7127 -19790 7161 -19756
rect 7195 -19790 7229 -19756
rect 7263 -19790 7297 -19756
rect 7331 -19790 7365 -19756
rect 7399 -19790 7433 -19756
rect 7941 -19790 7975 -19756
rect 8009 -19790 8043 -19756
rect 8077 -19790 8111 -19756
rect 8145 -19790 8179 -19756
rect 8213 -19790 8247 -19756
rect 8281 -19790 8315 -19756
rect 8349 -19790 8383 -19756
rect 8417 -19790 8451 -19756
rect 8959 -19790 8993 -19756
rect 9027 -19790 9061 -19756
rect 9095 -19790 9129 -19756
rect 9163 -19790 9197 -19756
rect 9231 -19790 9265 -19756
rect 9299 -19790 9333 -19756
rect 9367 -19790 9401 -19756
rect 9435 -19790 9469 -19756
rect 9977 -19790 10011 -19756
rect 10045 -19790 10079 -19756
rect 10113 -19790 10147 -19756
rect 10181 -19790 10215 -19756
rect 10249 -19790 10283 -19756
rect 10317 -19790 10351 -19756
rect 10385 -19790 10419 -19756
rect 10453 -19790 10487 -19756
rect 10995 -19790 11029 -19756
rect 11063 -19790 11097 -19756
rect 11131 -19790 11165 -19756
rect 11199 -19790 11233 -19756
rect 11267 -19790 11301 -19756
rect 11335 -19790 11369 -19756
rect 11403 -19790 11437 -19756
rect 11471 -19790 11505 -19756
rect 12013 -19790 12047 -19756
rect 12081 -19790 12115 -19756
rect 12149 -19790 12183 -19756
rect 12217 -19790 12251 -19756
rect 12285 -19790 12319 -19756
rect 12353 -19790 12387 -19756
rect 12421 -19790 12455 -19756
rect 12489 -19790 12523 -19756
rect 13031 -19790 13065 -19756
rect 13099 -19790 13133 -19756
rect 13167 -19790 13201 -19756
rect 13235 -19790 13269 -19756
rect 13303 -19790 13337 -19756
rect 13371 -19790 13405 -19756
rect 13439 -19790 13473 -19756
rect 13507 -19790 13541 -19756
rect 14049 -19790 14083 -19756
rect 14117 -19790 14151 -19756
rect 14185 -19790 14219 -19756
rect 14253 -19790 14287 -19756
rect 14321 -19790 14355 -19756
rect 14389 -19790 14423 -19756
rect 14457 -19790 14491 -19756
rect 14525 -19790 14559 -19756
rect 15067 -19790 15101 -19756
rect 15135 -19790 15169 -19756
rect 15203 -19790 15237 -19756
rect 15271 -19790 15305 -19756
rect 15339 -19790 15373 -19756
rect 15407 -19790 15441 -19756
rect 15475 -19790 15509 -19756
rect 15543 -19790 15577 -19756
rect 16085 -19790 16119 -19756
rect 16153 -19790 16187 -19756
rect 16221 -19790 16255 -19756
rect 16289 -19790 16323 -19756
rect 16357 -19790 16391 -19756
rect 16425 -19790 16459 -19756
rect 16493 -19790 16527 -19756
rect 16561 -19790 16595 -19756
rect 17103 -19790 17137 -19756
rect 17171 -19790 17205 -19756
rect 17239 -19790 17273 -19756
rect 17307 -19790 17341 -19756
rect 17375 -19790 17409 -19756
rect 17443 -19790 17477 -19756
rect 17511 -19790 17545 -19756
rect 17579 -19790 17613 -19756
rect 18121 -19790 18155 -19756
rect 18189 -19790 18223 -19756
rect 18257 -19790 18291 -19756
rect 18325 -19790 18359 -19756
rect 18393 -19790 18427 -19756
rect 18461 -19790 18495 -19756
rect 18529 -19790 18563 -19756
rect 18597 -19790 18631 -19756
rect 19139 -19790 19173 -19756
rect 19207 -19790 19241 -19756
rect 19275 -19790 19309 -19756
rect 19343 -19790 19377 -19756
rect 19411 -19790 19445 -19756
rect 19479 -19790 19513 -19756
rect 19547 -19790 19581 -19756
rect 19615 -19790 19649 -19756
rect 20157 -19790 20191 -19756
rect 20225 -19790 20259 -19756
rect 20293 -19790 20327 -19756
rect 20361 -19790 20395 -19756
rect 20429 -19790 20463 -19756
rect 20497 -19790 20531 -19756
rect 20565 -19790 20599 -19756
rect 20633 -19790 20667 -19756
rect 21175 -19790 21209 -19756
rect 21243 -19790 21277 -19756
rect 21311 -19790 21345 -19756
rect 21379 -19790 21413 -19756
rect 21447 -19790 21481 -19756
rect 21515 -19790 21549 -19756
rect 21583 -19790 21617 -19756
rect 21651 -19790 21685 -19756
rect 22193 -19790 22227 -19756
rect 22261 -19790 22295 -19756
rect 22329 -19790 22363 -19756
rect 22397 -19790 22431 -19756
rect 22465 -19790 22499 -19756
rect 22533 -19790 22567 -19756
rect 22601 -19790 22635 -19756
rect 22669 -19790 22703 -19756
rect -2215 -19894 -2181 -19860
rect -1997 -19894 -1963 -19860
rect -1779 -19894 -1745 -19860
rect -1561 -19894 -1527 -19860
rect -1343 -19894 -1309 -19860
rect -1125 -19894 -1091 -19860
rect -907 -19894 -873 -19860
rect -689 -19894 -655 -19860
rect -471 -19894 -437 -19860
rect -253 -19894 -219 -19860
rect 2851 -20314 2885 -20280
rect 2919 -20314 2953 -20280
rect 2987 -20314 3021 -20280
rect 3055 -20314 3089 -20280
rect 3123 -20314 3157 -20280
rect 3191 -20314 3225 -20280
rect 3259 -20314 3293 -20280
rect 3327 -20314 3361 -20280
rect 3869 -20314 3903 -20280
rect 3937 -20314 3971 -20280
rect 4005 -20314 4039 -20280
rect 4073 -20314 4107 -20280
rect 4141 -20314 4175 -20280
rect 4209 -20314 4243 -20280
rect 4277 -20314 4311 -20280
rect 4345 -20314 4379 -20280
rect 4887 -20314 4921 -20280
rect 4955 -20314 4989 -20280
rect 5023 -20314 5057 -20280
rect 5091 -20314 5125 -20280
rect 5159 -20314 5193 -20280
rect 5227 -20314 5261 -20280
rect 5295 -20314 5329 -20280
rect 5363 -20314 5397 -20280
rect 5905 -20314 5939 -20280
rect 5973 -20314 6007 -20280
rect 6041 -20314 6075 -20280
rect 6109 -20314 6143 -20280
rect 6177 -20314 6211 -20280
rect 6245 -20314 6279 -20280
rect 6313 -20314 6347 -20280
rect 6381 -20314 6415 -20280
rect 6923 -20314 6957 -20280
rect 6991 -20314 7025 -20280
rect 7059 -20314 7093 -20280
rect 7127 -20314 7161 -20280
rect 7195 -20314 7229 -20280
rect 7263 -20314 7297 -20280
rect 7331 -20314 7365 -20280
rect 7399 -20314 7433 -20280
rect 7941 -20314 7975 -20280
rect 8009 -20314 8043 -20280
rect 8077 -20314 8111 -20280
rect 8145 -20314 8179 -20280
rect 8213 -20314 8247 -20280
rect 8281 -20314 8315 -20280
rect 8349 -20314 8383 -20280
rect 8417 -20314 8451 -20280
rect 8959 -20314 8993 -20280
rect 9027 -20314 9061 -20280
rect 9095 -20314 9129 -20280
rect 9163 -20314 9197 -20280
rect 9231 -20314 9265 -20280
rect 9299 -20314 9333 -20280
rect 9367 -20314 9401 -20280
rect 9435 -20314 9469 -20280
rect 9977 -20314 10011 -20280
rect 10045 -20314 10079 -20280
rect 10113 -20314 10147 -20280
rect 10181 -20314 10215 -20280
rect 10249 -20314 10283 -20280
rect 10317 -20314 10351 -20280
rect 10385 -20314 10419 -20280
rect 10453 -20314 10487 -20280
rect 10995 -20314 11029 -20280
rect 11063 -20314 11097 -20280
rect 11131 -20314 11165 -20280
rect 11199 -20314 11233 -20280
rect 11267 -20314 11301 -20280
rect 11335 -20314 11369 -20280
rect 11403 -20314 11437 -20280
rect 11471 -20314 11505 -20280
rect 12013 -20314 12047 -20280
rect 12081 -20314 12115 -20280
rect 12149 -20314 12183 -20280
rect 12217 -20314 12251 -20280
rect 12285 -20314 12319 -20280
rect 12353 -20314 12387 -20280
rect 12421 -20314 12455 -20280
rect 12489 -20314 12523 -20280
rect 13031 -20314 13065 -20280
rect 13099 -20314 13133 -20280
rect 13167 -20314 13201 -20280
rect 13235 -20314 13269 -20280
rect 13303 -20314 13337 -20280
rect 13371 -20314 13405 -20280
rect 13439 -20314 13473 -20280
rect 13507 -20314 13541 -20280
rect 14049 -20314 14083 -20280
rect 14117 -20314 14151 -20280
rect 14185 -20314 14219 -20280
rect 14253 -20314 14287 -20280
rect 14321 -20314 14355 -20280
rect 14389 -20314 14423 -20280
rect 14457 -20314 14491 -20280
rect 14525 -20314 14559 -20280
rect 15067 -20314 15101 -20280
rect 15135 -20314 15169 -20280
rect 15203 -20314 15237 -20280
rect 15271 -20314 15305 -20280
rect 15339 -20314 15373 -20280
rect 15407 -20314 15441 -20280
rect 15475 -20314 15509 -20280
rect 15543 -20314 15577 -20280
rect 16085 -20314 16119 -20280
rect 16153 -20314 16187 -20280
rect 16221 -20314 16255 -20280
rect 16289 -20314 16323 -20280
rect 16357 -20314 16391 -20280
rect 16425 -20314 16459 -20280
rect 16493 -20314 16527 -20280
rect 16561 -20314 16595 -20280
rect 17103 -20314 17137 -20280
rect 17171 -20314 17205 -20280
rect 17239 -20314 17273 -20280
rect 17307 -20314 17341 -20280
rect 17375 -20314 17409 -20280
rect 17443 -20314 17477 -20280
rect 17511 -20314 17545 -20280
rect 17579 -20314 17613 -20280
rect 18121 -20314 18155 -20280
rect 18189 -20314 18223 -20280
rect 18257 -20314 18291 -20280
rect 18325 -20314 18359 -20280
rect 18393 -20314 18427 -20280
rect 18461 -20314 18495 -20280
rect 18529 -20314 18563 -20280
rect 18597 -20314 18631 -20280
rect 19139 -20314 19173 -20280
rect 19207 -20314 19241 -20280
rect 19275 -20314 19309 -20280
rect 19343 -20314 19377 -20280
rect 19411 -20314 19445 -20280
rect 19479 -20314 19513 -20280
rect 19547 -20314 19581 -20280
rect 19615 -20314 19649 -20280
rect 20157 -20314 20191 -20280
rect 20225 -20314 20259 -20280
rect 20293 -20314 20327 -20280
rect 20361 -20314 20395 -20280
rect 20429 -20314 20463 -20280
rect 20497 -20314 20531 -20280
rect 20565 -20314 20599 -20280
rect 20633 -20314 20667 -20280
rect 21175 -20314 21209 -20280
rect 21243 -20314 21277 -20280
rect 21311 -20314 21345 -20280
rect 21379 -20314 21413 -20280
rect 21447 -20314 21481 -20280
rect 21515 -20314 21549 -20280
rect 21583 -20314 21617 -20280
rect 21651 -20314 21685 -20280
rect 22193 -20314 22227 -20280
rect 22261 -20314 22295 -20280
rect 22329 -20314 22363 -20280
rect 22397 -20314 22431 -20280
rect 22465 -20314 22499 -20280
rect 22533 -20314 22567 -20280
rect 22601 -20314 22635 -20280
rect 22669 -20314 22703 -20280
rect -2215 -20416 -2181 -20382
rect -1997 -20416 -1963 -20382
rect -1779 -20416 -1745 -20382
rect -1561 -20416 -1527 -20382
rect -1343 -20416 -1309 -20382
rect -1125 -20416 -1091 -20382
rect -907 -20416 -873 -20382
rect -689 -20416 -655 -20382
rect -471 -20416 -437 -20382
rect -253 -20416 -219 -20382
rect -2215 -20726 -2181 -20692
rect -1997 -20726 -1963 -20692
rect -1779 -20726 -1745 -20692
rect -1561 -20726 -1527 -20692
rect -1343 -20726 -1309 -20692
rect -1125 -20726 -1091 -20692
rect -907 -20726 -873 -20692
rect -689 -20726 -655 -20692
rect -471 -20726 -437 -20692
rect -253 -20726 -219 -20692
rect 2851 -21024 2885 -20990
rect 2919 -21024 2953 -20990
rect 2987 -21024 3021 -20990
rect 3055 -21024 3089 -20990
rect 3123 -21024 3157 -20990
rect 3191 -21024 3225 -20990
rect 3259 -21024 3293 -20990
rect 3327 -21024 3361 -20990
rect 3869 -21024 3903 -20990
rect 3937 -21024 3971 -20990
rect 4005 -21024 4039 -20990
rect 4073 -21024 4107 -20990
rect 4141 -21024 4175 -20990
rect 4209 -21024 4243 -20990
rect 4277 -21024 4311 -20990
rect 4345 -21024 4379 -20990
rect 4887 -21024 4921 -20990
rect 4955 -21024 4989 -20990
rect 5023 -21024 5057 -20990
rect 5091 -21024 5125 -20990
rect 5159 -21024 5193 -20990
rect 5227 -21024 5261 -20990
rect 5295 -21024 5329 -20990
rect 5363 -21024 5397 -20990
rect 5905 -21024 5939 -20990
rect 5973 -21024 6007 -20990
rect 6041 -21024 6075 -20990
rect 6109 -21024 6143 -20990
rect 6177 -21024 6211 -20990
rect 6245 -21024 6279 -20990
rect 6313 -21024 6347 -20990
rect 6381 -21024 6415 -20990
rect 6923 -21024 6957 -20990
rect 6991 -21024 7025 -20990
rect 7059 -21024 7093 -20990
rect 7127 -21024 7161 -20990
rect 7195 -21024 7229 -20990
rect 7263 -21024 7297 -20990
rect 7331 -21024 7365 -20990
rect 7399 -21024 7433 -20990
rect 7941 -21024 7975 -20990
rect 8009 -21024 8043 -20990
rect 8077 -21024 8111 -20990
rect 8145 -21024 8179 -20990
rect 8213 -21024 8247 -20990
rect 8281 -21024 8315 -20990
rect 8349 -21024 8383 -20990
rect 8417 -21024 8451 -20990
rect 8959 -21024 8993 -20990
rect 9027 -21024 9061 -20990
rect 9095 -21024 9129 -20990
rect 9163 -21024 9197 -20990
rect 9231 -21024 9265 -20990
rect 9299 -21024 9333 -20990
rect 9367 -21024 9401 -20990
rect 9435 -21024 9469 -20990
rect 9977 -21024 10011 -20990
rect 10045 -21024 10079 -20990
rect 10113 -21024 10147 -20990
rect 10181 -21024 10215 -20990
rect 10249 -21024 10283 -20990
rect 10317 -21024 10351 -20990
rect 10385 -21024 10419 -20990
rect 10453 -21024 10487 -20990
rect 10995 -21024 11029 -20990
rect 11063 -21024 11097 -20990
rect 11131 -21024 11165 -20990
rect 11199 -21024 11233 -20990
rect 11267 -21024 11301 -20990
rect 11335 -21024 11369 -20990
rect 11403 -21024 11437 -20990
rect 11471 -21024 11505 -20990
rect 12013 -21024 12047 -20990
rect 12081 -21024 12115 -20990
rect 12149 -21024 12183 -20990
rect 12217 -21024 12251 -20990
rect 12285 -21024 12319 -20990
rect 12353 -21024 12387 -20990
rect 12421 -21024 12455 -20990
rect 12489 -21024 12523 -20990
rect 13031 -21024 13065 -20990
rect 13099 -21024 13133 -20990
rect 13167 -21024 13201 -20990
rect 13235 -21024 13269 -20990
rect 13303 -21024 13337 -20990
rect 13371 -21024 13405 -20990
rect 13439 -21024 13473 -20990
rect 13507 -21024 13541 -20990
rect 14049 -21024 14083 -20990
rect 14117 -21024 14151 -20990
rect 14185 -21024 14219 -20990
rect 14253 -21024 14287 -20990
rect 14321 -21024 14355 -20990
rect 14389 -21024 14423 -20990
rect 14457 -21024 14491 -20990
rect 14525 -21024 14559 -20990
rect 15067 -21024 15101 -20990
rect 15135 -21024 15169 -20990
rect 15203 -21024 15237 -20990
rect 15271 -21024 15305 -20990
rect 15339 -21024 15373 -20990
rect 15407 -21024 15441 -20990
rect 15475 -21024 15509 -20990
rect 15543 -21024 15577 -20990
rect 16085 -21024 16119 -20990
rect 16153 -21024 16187 -20990
rect 16221 -21024 16255 -20990
rect 16289 -21024 16323 -20990
rect 16357 -21024 16391 -20990
rect 16425 -21024 16459 -20990
rect 16493 -21024 16527 -20990
rect 16561 -21024 16595 -20990
rect 17103 -21024 17137 -20990
rect 17171 -21024 17205 -20990
rect 17239 -21024 17273 -20990
rect 17307 -21024 17341 -20990
rect 17375 -21024 17409 -20990
rect 17443 -21024 17477 -20990
rect 17511 -21024 17545 -20990
rect 17579 -21024 17613 -20990
rect 18121 -21024 18155 -20990
rect 18189 -21024 18223 -20990
rect 18257 -21024 18291 -20990
rect 18325 -21024 18359 -20990
rect 18393 -21024 18427 -20990
rect 18461 -21024 18495 -20990
rect 18529 -21024 18563 -20990
rect 18597 -21024 18631 -20990
rect 19139 -21024 19173 -20990
rect 19207 -21024 19241 -20990
rect 19275 -21024 19309 -20990
rect 19343 -21024 19377 -20990
rect 19411 -21024 19445 -20990
rect 19479 -21024 19513 -20990
rect 19547 -21024 19581 -20990
rect 19615 -21024 19649 -20990
rect 20157 -21024 20191 -20990
rect 20225 -21024 20259 -20990
rect 20293 -21024 20327 -20990
rect 20361 -21024 20395 -20990
rect 20429 -21024 20463 -20990
rect 20497 -21024 20531 -20990
rect 20565 -21024 20599 -20990
rect 20633 -21024 20667 -20990
rect 21175 -21024 21209 -20990
rect 21243 -21024 21277 -20990
rect 21311 -21024 21345 -20990
rect 21379 -21024 21413 -20990
rect 21447 -21024 21481 -20990
rect 21515 -21024 21549 -20990
rect 21583 -21024 21617 -20990
rect 21651 -21024 21685 -20990
rect 22193 -21024 22227 -20990
rect 22261 -21024 22295 -20990
rect 22329 -21024 22363 -20990
rect 22397 -21024 22431 -20990
rect 22465 -21024 22499 -20990
rect 22533 -21024 22567 -20990
rect 22601 -21024 22635 -20990
rect 22669 -21024 22703 -20990
rect 2851 -21546 2885 -21512
rect 2919 -21546 2953 -21512
rect 2987 -21546 3021 -21512
rect 3055 -21546 3089 -21512
rect 3123 -21546 3157 -21512
rect 3191 -21546 3225 -21512
rect 3259 -21546 3293 -21512
rect 3327 -21546 3361 -21512
rect 3869 -21546 3903 -21512
rect 3937 -21546 3971 -21512
rect 4005 -21546 4039 -21512
rect 4073 -21546 4107 -21512
rect 4141 -21546 4175 -21512
rect 4209 -21546 4243 -21512
rect 4277 -21546 4311 -21512
rect 4345 -21546 4379 -21512
rect 4887 -21546 4921 -21512
rect 4955 -21546 4989 -21512
rect 5023 -21546 5057 -21512
rect 5091 -21546 5125 -21512
rect 5159 -21546 5193 -21512
rect 5227 -21546 5261 -21512
rect 5295 -21546 5329 -21512
rect 5363 -21546 5397 -21512
rect 5905 -21546 5939 -21512
rect 5973 -21546 6007 -21512
rect 6041 -21546 6075 -21512
rect 6109 -21546 6143 -21512
rect 6177 -21546 6211 -21512
rect 6245 -21546 6279 -21512
rect 6313 -21546 6347 -21512
rect 6381 -21546 6415 -21512
rect 6923 -21546 6957 -21512
rect 6991 -21546 7025 -21512
rect 7059 -21546 7093 -21512
rect 7127 -21546 7161 -21512
rect 7195 -21546 7229 -21512
rect 7263 -21546 7297 -21512
rect 7331 -21546 7365 -21512
rect 7399 -21546 7433 -21512
rect 7941 -21546 7975 -21512
rect 8009 -21546 8043 -21512
rect 8077 -21546 8111 -21512
rect 8145 -21546 8179 -21512
rect 8213 -21546 8247 -21512
rect 8281 -21546 8315 -21512
rect 8349 -21546 8383 -21512
rect 8417 -21546 8451 -21512
rect 8959 -21546 8993 -21512
rect 9027 -21546 9061 -21512
rect 9095 -21546 9129 -21512
rect 9163 -21546 9197 -21512
rect 9231 -21546 9265 -21512
rect 9299 -21546 9333 -21512
rect 9367 -21546 9401 -21512
rect 9435 -21546 9469 -21512
rect 9977 -21546 10011 -21512
rect 10045 -21546 10079 -21512
rect 10113 -21546 10147 -21512
rect 10181 -21546 10215 -21512
rect 10249 -21546 10283 -21512
rect 10317 -21546 10351 -21512
rect 10385 -21546 10419 -21512
rect 10453 -21546 10487 -21512
rect 10995 -21546 11029 -21512
rect 11063 -21546 11097 -21512
rect 11131 -21546 11165 -21512
rect 11199 -21546 11233 -21512
rect 11267 -21546 11301 -21512
rect 11335 -21546 11369 -21512
rect 11403 -21546 11437 -21512
rect 11471 -21546 11505 -21512
rect 12013 -21546 12047 -21512
rect 12081 -21546 12115 -21512
rect 12149 -21546 12183 -21512
rect 12217 -21546 12251 -21512
rect 12285 -21546 12319 -21512
rect 12353 -21546 12387 -21512
rect 12421 -21546 12455 -21512
rect 12489 -21546 12523 -21512
rect 13031 -21546 13065 -21512
rect 13099 -21546 13133 -21512
rect 13167 -21546 13201 -21512
rect 13235 -21546 13269 -21512
rect 13303 -21546 13337 -21512
rect 13371 -21546 13405 -21512
rect 13439 -21546 13473 -21512
rect 13507 -21546 13541 -21512
rect 14049 -21546 14083 -21512
rect 14117 -21546 14151 -21512
rect 14185 -21546 14219 -21512
rect 14253 -21546 14287 -21512
rect 14321 -21546 14355 -21512
rect 14389 -21546 14423 -21512
rect 14457 -21546 14491 -21512
rect 14525 -21546 14559 -21512
rect 15067 -21546 15101 -21512
rect 15135 -21546 15169 -21512
rect 15203 -21546 15237 -21512
rect 15271 -21546 15305 -21512
rect 15339 -21546 15373 -21512
rect 15407 -21546 15441 -21512
rect 15475 -21546 15509 -21512
rect 15543 -21546 15577 -21512
rect 16085 -21546 16119 -21512
rect 16153 -21546 16187 -21512
rect 16221 -21546 16255 -21512
rect 16289 -21546 16323 -21512
rect 16357 -21546 16391 -21512
rect 16425 -21546 16459 -21512
rect 16493 -21546 16527 -21512
rect 16561 -21546 16595 -21512
rect 17103 -21546 17137 -21512
rect 17171 -21546 17205 -21512
rect 17239 -21546 17273 -21512
rect 17307 -21546 17341 -21512
rect 17375 -21546 17409 -21512
rect 17443 -21546 17477 -21512
rect 17511 -21546 17545 -21512
rect 17579 -21546 17613 -21512
rect 18121 -21546 18155 -21512
rect 18189 -21546 18223 -21512
rect 18257 -21546 18291 -21512
rect 18325 -21546 18359 -21512
rect 18393 -21546 18427 -21512
rect 18461 -21546 18495 -21512
rect 18529 -21546 18563 -21512
rect 18597 -21546 18631 -21512
rect 19139 -21546 19173 -21512
rect 19207 -21546 19241 -21512
rect 19275 -21546 19309 -21512
rect 19343 -21546 19377 -21512
rect 19411 -21546 19445 -21512
rect 19479 -21546 19513 -21512
rect 19547 -21546 19581 -21512
rect 19615 -21546 19649 -21512
rect 20157 -21546 20191 -21512
rect 20225 -21546 20259 -21512
rect 20293 -21546 20327 -21512
rect 20361 -21546 20395 -21512
rect 20429 -21546 20463 -21512
rect 20497 -21546 20531 -21512
rect 20565 -21546 20599 -21512
rect 20633 -21546 20667 -21512
rect 21175 -21546 21209 -21512
rect 21243 -21546 21277 -21512
rect 21311 -21546 21345 -21512
rect 21379 -21546 21413 -21512
rect 21447 -21546 21481 -21512
rect 21515 -21546 21549 -21512
rect 21583 -21546 21617 -21512
rect 21651 -21546 21685 -21512
rect 22193 -21546 22227 -21512
rect 22261 -21546 22295 -21512
rect 22329 -21546 22363 -21512
rect 22397 -21546 22431 -21512
rect 22465 -21546 22499 -21512
rect 22533 -21546 22567 -21512
rect 22601 -21546 22635 -21512
rect 22669 -21546 22703 -21512
rect -9134 -21743 -9100 -21709
rect -9066 -21743 -9032 -21709
rect -8998 -21743 -8964 -21709
rect -8930 -21743 -8896 -21709
rect -8862 -21743 -8828 -21709
rect -8794 -21743 -8760 -21709
rect -8726 -21743 -8692 -21709
rect -8658 -21743 -8624 -21709
rect -8116 -21743 -8082 -21709
rect -8048 -21743 -8014 -21709
rect -7980 -21743 -7946 -21709
rect -7912 -21743 -7878 -21709
rect -7844 -21743 -7810 -21709
rect -7776 -21743 -7742 -21709
rect -7708 -21743 -7674 -21709
rect -7640 -21743 -7606 -21709
rect -7098 -21743 -7064 -21709
rect -7030 -21743 -6996 -21709
rect -6962 -21743 -6928 -21709
rect -6894 -21743 -6860 -21709
rect -6826 -21743 -6792 -21709
rect -6758 -21743 -6724 -21709
rect -6690 -21743 -6656 -21709
rect -6622 -21743 -6588 -21709
rect -6080 -21743 -6046 -21709
rect -6012 -21743 -5978 -21709
rect -5944 -21743 -5910 -21709
rect -5876 -21743 -5842 -21709
rect -5808 -21743 -5774 -21709
rect -5740 -21743 -5706 -21709
rect -5672 -21743 -5638 -21709
rect -5604 -21743 -5570 -21709
rect -5062 -21743 -5028 -21709
rect -4994 -21743 -4960 -21709
rect -4926 -21743 -4892 -21709
rect -4858 -21743 -4824 -21709
rect -4790 -21743 -4756 -21709
rect -4722 -21743 -4688 -21709
rect -4654 -21743 -4620 -21709
rect -4586 -21743 -4552 -21709
rect -4044 -21743 -4010 -21709
rect -3976 -21743 -3942 -21709
rect -3908 -21743 -3874 -21709
rect -3840 -21743 -3806 -21709
rect -3772 -21743 -3738 -21709
rect -3704 -21743 -3670 -21709
rect -3636 -21743 -3602 -21709
rect -3568 -21743 -3534 -21709
rect -2295 -21742 -2261 -21708
rect -2227 -21742 -2193 -21708
rect -1997 -21742 -1963 -21708
rect -1929 -21742 -1895 -21708
rect -1699 -21742 -1665 -21708
rect -1631 -21742 -1597 -21708
rect -1401 -21742 -1367 -21708
rect -1333 -21742 -1299 -21708
rect -1103 -21742 -1069 -21708
rect -1035 -21742 -1001 -21708
rect -805 -21742 -771 -21708
rect -737 -21742 -703 -21708
rect -507 -21742 -473 -21708
rect -439 -21742 -405 -21708
rect -209 -21742 -175 -21708
rect -141 -21742 -107 -21708
rect 89 -21742 123 -21708
rect 157 -21742 191 -21708
rect 387 -21742 421 -21708
rect 455 -21742 489 -21708
rect 685 -21742 719 -21708
rect 753 -21742 787 -21708
rect 2851 -22256 2885 -22222
rect 2919 -22256 2953 -22222
rect 2987 -22256 3021 -22222
rect 3055 -22256 3089 -22222
rect 3123 -22256 3157 -22222
rect 3191 -22256 3225 -22222
rect 3259 -22256 3293 -22222
rect 3327 -22256 3361 -22222
rect 3869 -22256 3903 -22222
rect 3937 -22256 3971 -22222
rect 4005 -22256 4039 -22222
rect 4073 -22256 4107 -22222
rect 4141 -22256 4175 -22222
rect 4209 -22256 4243 -22222
rect 4277 -22256 4311 -22222
rect 4345 -22256 4379 -22222
rect 4887 -22256 4921 -22222
rect 4955 -22256 4989 -22222
rect 5023 -22256 5057 -22222
rect 5091 -22256 5125 -22222
rect 5159 -22256 5193 -22222
rect 5227 -22256 5261 -22222
rect 5295 -22256 5329 -22222
rect 5363 -22256 5397 -22222
rect 5905 -22256 5939 -22222
rect 5973 -22256 6007 -22222
rect 6041 -22256 6075 -22222
rect 6109 -22256 6143 -22222
rect 6177 -22256 6211 -22222
rect 6245 -22256 6279 -22222
rect 6313 -22256 6347 -22222
rect 6381 -22256 6415 -22222
rect 6923 -22256 6957 -22222
rect 6991 -22256 7025 -22222
rect 7059 -22256 7093 -22222
rect 7127 -22256 7161 -22222
rect 7195 -22256 7229 -22222
rect 7263 -22256 7297 -22222
rect 7331 -22256 7365 -22222
rect 7399 -22256 7433 -22222
rect 7941 -22256 7975 -22222
rect 8009 -22256 8043 -22222
rect 8077 -22256 8111 -22222
rect 8145 -22256 8179 -22222
rect 8213 -22256 8247 -22222
rect 8281 -22256 8315 -22222
rect 8349 -22256 8383 -22222
rect 8417 -22256 8451 -22222
rect 8959 -22256 8993 -22222
rect 9027 -22256 9061 -22222
rect 9095 -22256 9129 -22222
rect 9163 -22256 9197 -22222
rect 9231 -22256 9265 -22222
rect 9299 -22256 9333 -22222
rect 9367 -22256 9401 -22222
rect 9435 -22256 9469 -22222
rect 9977 -22256 10011 -22222
rect 10045 -22256 10079 -22222
rect 10113 -22256 10147 -22222
rect 10181 -22256 10215 -22222
rect 10249 -22256 10283 -22222
rect 10317 -22256 10351 -22222
rect 10385 -22256 10419 -22222
rect 10453 -22256 10487 -22222
rect 10995 -22256 11029 -22222
rect 11063 -22256 11097 -22222
rect 11131 -22256 11165 -22222
rect 11199 -22256 11233 -22222
rect 11267 -22256 11301 -22222
rect 11335 -22256 11369 -22222
rect 11403 -22256 11437 -22222
rect 11471 -22256 11505 -22222
rect 12013 -22256 12047 -22222
rect 12081 -22256 12115 -22222
rect 12149 -22256 12183 -22222
rect 12217 -22256 12251 -22222
rect 12285 -22256 12319 -22222
rect 12353 -22256 12387 -22222
rect 12421 -22256 12455 -22222
rect 12489 -22256 12523 -22222
rect 13031 -22256 13065 -22222
rect 13099 -22256 13133 -22222
rect 13167 -22256 13201 -22222
rect 13235 -22256 13269 -22222
rect 13303 -22256 13337 -22222
rect 13371 -22256 13405 -22222
rect 13439 -22256 13473 -22222
rect 13507 -22256 13541 -22222
rect 14049 -22256 14083 -22222
rect 14117 -22256 14151 -22222
rect 14185 -22256 14219 -22222
rect 14253 -22256 14287 -22222
rect 14321 -22256 14355 -22222
rect 14389 -22256 14423 -22222
rect 14457 -22256 14491 -22222
rect 14525 -22256 14559 -22222
rect 15067 -22256 15101 -22222
rect 15135 -22256 15169 -22222
rect 15203 -22256 15237 -22222
rect 15271 -22256 15305 -22222
rect 15339 -22256 15373 -22222
rect 15407 -22256 15441 -22222
rect 15475 -22256 15509 -22222
rect 15543 -22256 15577 -22222
rect 16085 -22256 16119 -22222
rect 16153 -22256 16187 -22222
rect 16221 -22256 16255 -22222
rect 16289 -22256 16323 -22222
rect 16357 -22256 16391 -22222
rect 16425 -22256 16459 -22222
rect 16493 -22256 16527 -22222
rect 16561 -22256 16595 -22222
rect 17103 -22256 17137 -22222
rect 17171 -22256 17205 -22222
rect 17239 -22256 17273 -22222
rect 17307 -22256 17341 -22222
rect 17375 -22256 17409 -22222
rect 17443 -22256 17477 -22222
rect 17511 -22256 17545 -22222
rect 17579 -22256 17613 -22222
rect 18121 -22256 18155 -22222
rect 18189 -22256 18223 -22222
rect 18257 -22256 18291 -22222
rect 18325 -22256 18359 -22222
rect 18393 -22256 18427 -22222
rect 18461 -22256 18495 -22222
rect 18529 -22256 18563 -22222
rect 18597 -22256 18631 -22222
rect 19139 -22256 19173 -22222
rect 19207 -22256 19241 -22222
rect 19275 -22256 19309 -22222
rect 19343 -22256 19377 -22222
rect 19411 -22256 19445 -22222
rect 19479 -22256 19513 -22222
rect 19547 -22256 19581 -22222
rect 19615 -22256 19649 -22222
rect 20157 -22256 20191 -22222
rect 20225 -22256 20259 -22222
rect 20293 -22256 20327 -22222
rect 20361 -22256 20395 -22222
rect 20429 -22256 20463 -22222
rect 20497 -22256 20531 -22222
rect 20565 -22256 20599 -22222
rect 20633 -22256 20667 -22222
rect 21175 -22256 21209 -22222
rect 21243 -22256 21277 -22222
rect 21311 -22256 21345 -22222
rect 21379 -22256 21413 -22222
rect 21447 -22256 21481 -22222
rect 21515 -22256 21549 -22222
rect 21583 -22256 21617 -22222
rect 21651 -22256 21685 -22222
rect 22193 -22256 22227 -22222
rect 22261 -22256 22295 -22222
rect 22329 -22256 22363 -22222
rect 22397 -22256 22431 -22222
rect 22465 -22256 22499 -22222
rect 22533 -22256 22567 -22222
rect 22601 -22256 22635 -22222
rect 22669 -22256 22703 -22222
rect -9134 -22453 -9100 -22419
rect -9066 -22453 -9032 -22419
rect -8998 -22453 -8964 -22419
rect -8930 -22453 -8896 -22419
rect -8862 -22453 -8828 -22419
rect -8794 -22453 -8760 -22419
rect -8726 -22453 -8692 -22419
rect -8658 -22453 -8624 -22419
rect -8116 -22453 -8082 -22419
rect -8048 -22453 -8014 -22419
rect -7980 -22453 -7946 -22419
rect -7912 -22453 -7878 -22419
rect -7844 -22453 -7810 -22419
rect -7776 -22453 -7742 -22419
rect -7708 -22453 -7674 -22419
rect -7640 -22453 -7606 -22419
rect -7098 -22453 -7064 -22419
rect -7030 -22453 -6996 -22419
rect -6962 -22453 -6928 -22419
rect -6894 -22453 -6860 -22419
rect -6826 -22453 -6792 -22419
rect -6758 -22453 -6724 -22419
rect -6690 -22453 -6656 -22419
rect -6622 -22453 -6588 -22419
rect -6080 -22453 -6046 -22419
rect -6012 -22453 -5978 -22419
rect -5944 -22453 -5910 -22419
rect -5876 -22453 -5842 -22419
rect -5808 -22453 -5774 -22419
rect -5740 -22453 -5706 -22419
rect -5672 -22453 -5638 -22419
rect -5604 -22453 -5570 -22419
rect -5062 -22453 -5028 -22419
rect -4994 -22453 -4960 -22419
rect -4926 -22453 -4892 -22419
rect -4858 -22453 -4824 -22419
rect -4790 -22453 -4756 -22419
rect -4722 -22453 -4688 -22419
rect -4654 -22453 -4620 -22419
rect -4586 -22453 -4552 -22419
rect -4044 -22453 -4010 -22419
rect -3976 -22453 -3942 -22419
rect -3908 -22453 -3874 -22419
rect -3840 -22453 -3806 -22419
rect -3772 -22453 -3738 -22419
rect -3704 -22453 -3670 -22419
rect -3636 -22453 -3602 -22419
rect -3568 -22453 -3534 -22419
rect -2295 -22452 -2261 -22418
rect -2227 -22452 -2193 -22418
rect -1997 -22452 -1963 -22418
rect -1929 -22452 -1895 -22418
rect -1699 -22452 -1665 -22418
rect -1631 -22452 -1597 -22418
rect -1401 -22452 -1367 -22418
rect -1333 -22452 -1299 -22418
rect -1103 -22452 -1069 -22418
rect -1035 -22452 -1001 -22418
rect -805 -22452 -771 -22418
rect -737 -22452 -703 -22418
rect -507 -22452 -473 -22418
rect -439 -22452 -405 -22418
rect -209 -22452 -175 -22418
rect -141 -22452 -107 -22418
rect 89 -22452 123 -22418
rect 157 -22452 191 -22418
rect 387 -22452 421 -22418
rect 455 -22452 489 -22418
rect 685 -22452 719 -22418
rect 753 -22452 787 -22418
rect 2851 -22780 2885 -22746
rect 2919 -22780 2953 -22746
rect 2987 -22780 3021 -22746
rect 3055 -22780 3089 -22746
rect 3123 -22780 3157 -22746
rect 3191 -22780 3225 -22746
rect 3259 -22780 3293 -22746
rect 3327 -22780 3361 -22746
rect -9135 -22856 -9101 -22822
rect -9067 -22856 -9033 -22822
rect -8999 -22856 -8965 -22822
rect -8931 -22856 -8897 -22822
rect -8863 -22856 -8829 -22822
rect -8795 -22856 -8761 -22822
rect -8727 -22856 -8693 -22822
rect -8659 -22856 -8625 -22822
rect -8117 -22856 -8083 -22822
rect -8049 -22856 -8015 -22822
rect -7981 -22856 -7947 -22822
rect -7913 -22856 -7879 -22822
rect -7845 -22856 -7811 -22822
rect -7777 -22856 -7743 -22822
rect -7709 -22856 -7675 -22822
rect -7641 -22856 -7607 -22822
rect -7099 -22856 -7065 -22822
rect -7031 -22856 -6997 -22822
rect -6963 -22856 -6929 -22822
rect -6895 -22856 -6861 -22822
rect -6827 -22856 -6793 -22822
rect -6759 -22856 -6725 -22822
rect -6691 -22856 -6657 -22822
rect -6623 -22856 -6589 -22822
rect -6081 -22856 -6047 -22822
rect -6013 -22856 -5979 -22822
rect -5945 -22856 -5911 -22822
rect -5877 -22856 -5843 -22822
rect -5809 -22856 -5775 -22822
rect -5741 -22856 -5707 -22822
rect -5673 -22856 -5639 -22822
rect -5605 -22856 -5571 -22822
rect -5063 -22856 -5029 -22822
rect -4995 -22856 -4961 -22822
rect -4927 -22856 -4893 -22822
rect -4859 -22856 -4825 -22822
rect -4791 -22856 -4757 -22822
rect -4723 -22856 -4689 -22822
rect -4655 -22856 -4621 -22822
rect -4587 -22856 -4553 -22822
rect -4045 -22856 -4011 -22822
rect -3977 -22856 -3943 -22822
rect -3909 -22856 -3875 -22822
rect -3841 -22856 -3807 -22822
rect -3773 -22856 -3739 -22822
rect -3705 -22856 -3671 -22822
rect -3637 -22856 -3603 -22822
rect -3569 -22856 -3535 -22822
rect -2295 -22854 -2261 -22820
rect -2227 -22854 -2193 -22820
rect -1997 -22854 -1963 -22820
rect -1929 -22854 -1895 -22820
rect -1699 -22854 -1665 -22820
rect -1631 -22854 -1597 -22820
rect -1401 -22854 -1367 -22820
rect -1333 -22854 -1299 -22820
rect -1103 -22854 -1069 -22820
rect -1035 -22854 -1001 -22820
rect -805 -22854 -771 -22820
rect -737 -22854 -703 -22820
rect -507 -22854 -473 -22820
rect -439 -22854 -405 -22820
rect -209 -22854 -175 -22820
rect -141 -22854 -107 -22820
rect 89 -22854 123 -22820
rect 157 -22854 191 -22820
rect 387 -22854 421 -22820
rect 455 -22854 489 -22820
rect 3869 -22780 3903 -22746
rect 3937 -22780 3971 -22746
rect 4005 -22780 4039 -22746
rect 4073 -22780 4107 -22746
rect 4141 -22780 4175 -22746
rect 4209 -22780 4243 -22746
rect 4277 -22780 4311 -22746
rect 4345 -22780 4379 -22746
rect 4887 -22780 4921 -22746
rect 4955 -22780 4989 -22746
rect 5023 -22780 5057 -22746
rect 5091 -22780 5125 -22746
rect 5159 -22780 5193 -22746
rect 5227 -22780 5261 -22746
rect 5295 -22780 5329 -22746
rect 5363 -22780 5397 -22746
rect 5905 -22780 5939 -22746
rect 5973 -22780 6007 -22746
rect 6041 -22780 6075 -22746
rect 6109 -22780 6143 -22746
rect 6177 -22780 6211 -22746
rect 6245 -22780 6279 -22746
rect 6313 -22780 6347 -22746
rect 6381 -22780 6415 -22746
rect 6923 -22780 6957 -22746
rect 6991 -22780 7025 -22746
rect 7059 -22780 7093 -22746
rect 7127 -22780 7161 -22746
rect 7195 -22780 7229 -22746
rect 7263 -22780 7297 -22746
rect 7331 -22780 7365 -22746
rect 7399 -22780 7433 -22746
rect 7941 -22780 7975 -22746
rect 8009 -22780 8043 -22746
rect 8077 -22780 8111 -22746
rect 8145 -22780 8179 -22746
rect 8213 -22780 8247 -22746
rect 8281 -22780 8315 -22746
rect 8349 -22780 8383 -22746
rect 8417 -22780 8451 -22746
rect 8959 -22780 8993 -22746
rect 9027 -22780 9061 -22746
rect 9095 -22780 9129 -22746
rect 9163 -22780 9197 -22746
rect 9231 -22780 9265 -22746
rect 9299 -22780 9333 -22746
rect 9367 -22780 9401 -22746
rect 9435 -22780 9469 -22746
rect 9977 -22780 10011 -22746
rect 10045 -22780 10079 -22746
rect 10113 -22780 10147 -22746
rect 10181 -22780 10215 -22746
rect 10249 -22780 10283 -22746
rect 10317 -22780 10351 -22746
rect 10385 -22780 10419 -22746
rect 10453 -22780 10487 -22746
rect 10995 -22780 11029 -22746
rect 11063 -22780 11097 -22746
rect 11131 -22780 11165 -22746
rect 11199 -22780 11233 -22746
rect 11267 -22780 11301 -22746
rect 11335 -22780 11369 -22746
rect 11403 -22780 11437 -22746
rect 11471 -22780 11505 -22746
rect 12013 -22780 12047 -22746
rect 12081 -22780 12115 -22746
rect 12149 -22780 12183 -22746
rect 12217 -22780 12251 -22746
rect 12285 -22780 12319 -22746
rect 12353 -22780 12387 -22746
rect 12421 -22780 12455 -22746
rect 12489 -22780 12523 -22746
rect 13031 -22780 13065 -22746
rect 13099 -22780 13133 -22746
rect 13167 -22780 13201 -22746
rect 13235 -22780 13269 -22746
rect 13303 -22780 13337 -22746
rect 13371 -22780 13405 -22746
rect 13439 -22780 13473 -22746
rect 13507 -22780 13541 -22746
rect 14049 -22780 14083 -22746
rect 14117 -22780 14151 -22746
rect 14185 -22780 14219 -22746
rect 14253 -22780 14287 -22746
rect 14321 -22780 14355 -22746
rect 14389 -22780 14423 -22746
rect 14457 -22780 14491 -22746
rect 14525 -22780 14559 -22746
rect 15067 -22780 15101 -22746
rect 15135 -22780 15169 -22746
rect 15203 -22780 15237 -22746
rect 15271 -22780 15305 -22746
rect 15339 -22780 15373 -22746
rect 15407 -22780 15441 -22746
rect 15475 -22780 15509 -22746
rect 15543 -22780 15577 -22746
rect 16085 -22780 16119 -22746
rect 16153 -22780 16187 -22746
rect 16221 -22780 16255 -22746
rect 16289 -22780 16323 -22746
rect 16357 -22780 16391 -22746
rect 16425 -22780 16459 -22746
rect 16493 -22780 16527 -22746
rect 16561 -22780 16595 -22746
rect 17103 -22780 17137 -22746
rect 17171 -22780 17205 -22746
rect 17239 -22780 17273 -22746
rect 17307 -22780 17341 -22746
rect 17375 -22780 17409 -22746
rect 17443 -22780 17477 -22746
rect 17511 -22780 17545 -22746
rect 17579 -22780 17613 -22746
rect 18121 -22780 18155 -22746
rect 18189 -22780 18223 -22746
rect 18257 -22780 18291 -22746
rect 18325 -22780 18359 -22746
rect 18393 -22780 18427 -22746
rect 18461 -22780 18495 -22746
rect 18529 -22780 18563 -22746
rect 18597 -22780 18631 -22746
rect 19139 -22780 19173 -22746
rect 19207 -22780 19241 -22746
rect 19275 -22780 19309 -22746
rect 19343 -22780 19377 -22746
rect 19411 -22780 19445 -22746
rect 19479 -22780 19513 -22746
rect 19547 -22780 19581 -22746
rect 19615 -22780 19649 -22746
rect 20157 -22780 20191 -22746
rect 20225 -22780 20259 -22746
rect 20293 -22780 20327 -22746
rect 20361 -22780 20395 -22746
rect 20429 -22780 20463 -22746
rect 20497 -22780 20531 -22746
rect 20565 -22780 20599 -22746
rect 20633 -22780 20667 -22746
rect 21175 -22780 21209 -22746
rect 21243 -22780 21277 -22746
rect 21311 -22780 21345 -22746
rect 21379 -22780 21413 -22746
rect 21447 -22780 21481 -22746
rect 21515 -22780 21549 -22746
rect 21583 -22780 21617 -22746
rect 21651 -22780 21685 -22746
rect 22193 -22780 22227 -22746
rect 22261 -22780 22295 -22746
rect 22329 -22780 22363 -22746
rect 22397 -22780 22431 -22746
rect 22465 -22780 22499 -22746
rect 22533 -22780 22567 -22746
rect 22601 -22780 22635 -22746
rect 22669 -22780 22703 -22746
rect 685 -22854 719 -22820
rect 753 -22854 787 -22820
rect 2851 -23490 2885 -23456
rect 2919 -23490 2953 -23456
rect 2987 -23490 3021 -23456
rect 3055 -23490 3089 -23456
rect 3123 -23490 3157 -23456
rect 3191 -23490 3225 -23456
rect 3259 -23490 3293 -23456
rect 3327 -23490 3361 -23456
rect -9135 -23566 -9101 -23532
rect -9067 -23566 -9033 -23532
rect -8999 -23566 -8965 -23532
rect -8931 -23566 -8897 -23532
rect -8863 -23566 -8829 -23532
rect -8795 -23566 -8761 -23532
rect -8727 -23566 -8693 -23532
rect -8659 -23566 -8625 -23532
rect -8117 -23566 -8083 -23532
rect -8049 -23566 -8015 -23532
rect -7981 -23566 -7947 -23532
rect -7913 -23566 -7879 -23532
rect -7845 -23566 -7811 -23532
rect -7777 -23566 -7743 -23532
rect -7709 -23566 -7675 -23532
rect -7641 -23566 -7607 -23532
rect -7099 -23566 -7065 -23532
rect -7031 -23566 -6997 -23532
rect -6963 -23566 -6929 -23532
rect -6895 -23566 -6861 -23532
rect -6827 -23566 -6793 -23532
rect -6759 -23566 -6725 -23532
rect -6691 -23566 -6657 -23532
rect -6623 -23566 -6589 -23532
rect -6081 -23566 -6047 -23532
rect -6013 -23566 -5979 -23532
rect -5945 -23566 -5911 -23532
rect -5877 -23566 -5843 -23532
rect -5809 -23566 -5775 -23532
rect -5741 -23566 -5707 -23532
rect -5673 -23566 -5639 -23532
rect -5605 -23566 -5571 -23532
rect -5063 -23566 -5029 -23532
rect -4995 -23566 -4961 -23532
rect -4927 -23566 -4893 -23532
rect -4859 -23566 -4825 -23532
rect -4791 -23566 -4757 -23532
rect -4723 -23566 -4689 -23532
rect -4655 -23566 -4621 -23532
rect -4587 -23566 -4553 -23532
rect -4045 -23566 -4011 -23532
rect -3977 -23566 -3943 -23532
rect -3909 -23566 -3875 -23532
rect -3841 -23566 -3807 -23532
rect -3773 -23566 -3739 -23532
rect -3705 -23566 -3671 -23532
rect -3637 -23566 -3603 -23532
rect -3569 -23566 -3535 -23532
rect -2295 -23564 -2261 -23530
rect -2227 -23564 -2193 -23530
rect -1997 -23564 -1963 -23530
rect -1929 -23564 -1895 -23530
rect -1699 -23564 -1665 -23530
rect -1631 -23564 -1597 -23530
rect -1401 -23564 -1367 -23530
rect -1333 -23564 -1299 -23530
rect -1103 -23564 -1069 -23530
rect -1035 -23564 -1001 -23530
rect -805 -23564 -771 -23530
rect -737 -23564 -703 -23530
rect -507 -23564 -473 -23530
rect -439 -23564 -405 -23530
rect -209 -23564 -175 -23530
rect -141 -23564 -107 -23530
rect 89 -23564 123 -23530
rect 157 -23564 191 -23530
rect 387 -23564 421 -23530
rect 455 -23564 489 -23530
rect 3869 -23490 3903 -23456
rect 3937 -23490 3971 -23456
rect 4005 -23490 4039 -23456
rect 4073 -23490 4107 -23456
rect 4141 -23490 4175 -23456
rect 4209 -23490 4243 -23456
rect 4277 -23490 4311 -23456
rect 4345 -23490 4379 -23456
rect 4887 -23490 4921 -23456
rect 4955 -23490 4989 -23456
rect 5023 -23490 5057 -23456
rect 5091 -23490 5125 -23456
rect 5159 -23490 5193 -23456
rect 5227 -23490 5261 -23456
rect 5295 -23490 5329 -23456
rect 5363 -23490 5397 -23456
rect 5905 -23490 5939 -23456
rect 5973 -23490 6007 -23456
rect 6041 -23490 6075 -23456
rect 6109 -23490 6143 -23456
rect 6177 -23490 6211 -23456
rect 6245 -23490 6279 -23456
rect 6313 -23490 6347 -23456
rect 6381 -23490 6415 -23456
rect 6923 -23490 6957 -23456
rect 6991 -23490 7025 -23456
rect 7059 -23490 7093 -23456
rect 7127 -23490 7161 -23456
rect 7195 -23490 7229 -23456
rect 7263 -23490 7297 -23456
rect 7331 -23490 7365 -23456
rect 7399 -23490 7433 -23456
rect 7941 -23490 7975 -23456
rect 8009 -23490 8043 -23456
rect 8077 -23490 8111 -23456
rect 8145 -23490 8179 -23456
rect 8213 -23490 8247 -23456
rect 8281 -23490 8315 -23456
rect 8349 -23490 8383 -23456
rect 8417 -23490 8451 -23456
rect 8959 -23490 8993 -23456
rect 9027 -23490 9061 -23456
rect 9095 -23490 9129 -23456
rect 9163 -23490 9197 -23456
rect 9231 -23490 9265 -23456
rect 9299 -23490 9333 -23456
rect 9367 -23490 9401 -23456
rect 9435 -23490 9469 -23456
rect 9977 -23490 10011 -23456
rect 10045 -23490 10079 -23456
rect 10113 -23490 10147 -23456
rect 10181 -23490 10215 -23456
rect 10249 -23490 10283 -23456
rect 10317 -23490 10351 -23456
rect 10385 -23490 10419 -23456
rect 10453 -23490 10487 -23456
rect 10995 -23490 11029 -23456
rect 11063 -23490 11097 -23456
rect 11131 -23490 11165 -23456
rect 11199 -23490 11233 -23456
rect 11267 -23490 11301 -23456
rect 11335 -23490 11369 -23456
rect 11403 -23490 11437 -23456
rect 11471 -23490 11505 -23456
rect 12013 -23490 12047 -23456
rect 12081 -23490 12115 -23456
rect 12149 -23490 12183 -23456
rect 12217 -23490 12251 -23456
rect 12285 -23490 12319 -23456
rect 12353 -23490 12387 -23456
rect 12421 -23490 12455 -23456
rect 12489 -23490 12523 -23456
rect 13031 -23490 13065 -23456
rect 13099 -23490 13133 -23456
rect 13167 -23490 13201 -23456
rect 13235 -23490 13269 -23456
rect 13303 -23490 13337 -23456
rect 13371 -23490 13405 -23456
rect 13439 -23490 13473 -23456
rect 13507 -23490 13541 -23456
rect 14049 -23490 14083 -23456
rect 14117 -23490 14151 -23456
rect 14185 -23490 14219 -23456
rect 14253 -23490 14287 -23456
rect 14321 -23490 14355 -23456
rect 14389 -23490 14423 -23456
rect 14457 -23490 14491 -23456
rect 14525 -23490 14559 -23456
rect 15067 -23490 15101 -23456
rect 15135 -23490 15169 -23456
rect 15203 -23490 15237 -23456
rect 15271 -23490 15305 -23456
rect 15339 -23490 15373 -23456
rect 15407 -23490 15441 -23456
rect 15475 -23490 15509 -23456
rect 15543 -23490 15577 -23456
rect 16085 -23490 16119 -23456
rect 16153 -23490 16187 -23456
rect 16221 -23490 16255 -23456
rect 16289 -23490 16323 -23456
rect 16357 -23490 16391 -23456
rect 16425 -23490 16459 -23456
rect 16493 -23490 16527 -23456
rect 16561 -23490 16595 -23456
rect 17103 -23490 17137 -23456
rect 17171 -23490 17205 -23456
rect 17239 -23490 17273 -23456
rect 17307 -23490 17341 -23456
rect 17375 -23490 17409 -23456
rect 17443 -23490 17477 -23456
rect 17511 -23490 17545 -23456
rect 17579 -23490 17613 -23456
rect 18121 -23490 18155 -23456
rect 18189 -23490 18223 -23456
rect 18257 -23490 18291 -23456
rect 18325 -23490 18359 -23456
rect 18393 -23490 18427 -23456
rect 18461 -23490 18495 -23456
rect 18529 -23490 18563 -23456
rect 18597 -23490 18631 -23456
rect 19139 -23490 19173 -23456
rect 19207 -23490 19241 -23456
rect 19275 -23490 19309 -23456
rect 19343 -23490 19377 -23456
rect 19411 -23490 19445 -23456
rect 19479 -23490 19513 -23456
rect 19547 -23490 19581 -23456
rect 19615 -23490 19649 -23456
rect 20157 -23490 20191 -23456
rect 20225 -23490 20259 -23456
rect 20293 -23490 20327 -23456
rect 20361 -23490 20395 -23456
rect 20429 -23490 20463 -23456
rect 20497 -23490 20531 -23456
rect 20565 -23490 20599 -23456
rect 20633 -23490 20667 -23456
rect 21175 -23490 21209 -23456
rect 21243 -23490 21277 -23456
rect 21311 -23490 21345 -23456
rect 21379 -23490 21413 -23456
rect 21447 -23490 21481 -23456
rect 21515 -23490 21549 -23456
rect 21583 -23490 21617 -23456
rect 21651 -23490 21685 -23456
rect 22193 -23490 22227 -23456
rect 22261 -23490 22295 -23456
rect 22329 -23490 22363 -23456
rect 22397 -23490 22431 -23456
rect 22465 -23490 22499 -23456
rect 22533 -23490 22567 -23456
rect 22601 -23490 22635 -23456
rect 22669 -23490 22703 -23456
rect 685 -23564 719 -23530
rect 753 -23564 787 -23530
rect -9134 -23967 -9100 -23933
rect -9066 -23967 -9032 -23933
rect -8998 -23967 -8964 -23933
rect -8930 -23967 -8896 -23933
rect -8862 -23967 -8828 -23933
rect -8794 -23967 -8760 -23933
rect -8726 -23967 -8692 -23933
rect -8658 -23967 -8624 -23933
rect -8116 -23967 -8082 -23933
rect -8048 -23967 -8014 -23933
rect -7980 -23967 -7946 -23933
rect -7912 -23967 -7878 -23933
rect -7844 -23967 -7810 -23933
rect -7776 -23967 -7742 -23933
rect -7708 -23967 -7674 -23933
rect -7640 -23967 -7606 -23933
rect -7098 -23967 -7064 -23933
rect -7030 -23967 -6996 -23933
rect -6962 -23967 -6928 -23933
rect -6894 -23967 -6860 -23933
rect -6826 -23967 -6792 -23933
rect -6758 -23967 -6724 -23933
rect -6690 -23967 -6656 -23933
rect -6622 -23967 -6588 -23933
rect -6080 -23967 -6046 -23933
rect -6012 -23967 -5978 -23933
rect -5944 -23967 -5910 -23933
rect -5876 -23967 -5842 -23933
rect -5808 -23967 -5774 -23933
rect -5740 -23967 -5706 -23933
rect -5672 -23967 -5638 -23933
rect -5604 -23967 -5570 -23933
rect -5062 -23967 -5028 -23933
rect -4994 -23967 -4960 -23933
rect -4926 -23967 -4892 -23933
rect -4858 -23967 -4824 -23933
rect -4790 -23967 -4756 -23933
rect -4722 -23967 -4688 -23933
rect -4654 -23967 -4620 -23933
rect -4586 -23967 -4552 -23933
rect -4044 -23967 -4010 -23933
rect -3976 -23967 -3942 -23933
rect -3908 -23967 -3874 -23933
rect -3840 -23967 -3806 -23933
rect -3772 -23967 -3738 -23933
rect -3704 -23967 -3670 -23933
rect -3636 -23967 -3602 -23933
rect -3568 -23967 -3534 -23933
rect -2297 -23966 -2263 -23932
rect -2229 -23966 -2195 -23932
rect -1999 -23966 -1965 -23932
rect -1931 -23966 -1897 -23932
rect -1701 -23966 -1667 -23932
rect -1633 -23966 -1599 -23932
rect -1403 -23966 -1369 -23932
rect -1335 -23966 -1301 -23932
rect -1105 -23966 -1071 -23932
rect -1037 -23966 -1003 -23932
rect -807 -23966 -773 -23932
rect -739 -23966 -705 -23932
rect -509 -23966 -475 -23932
rect -441 -23966 -407 -23932
rect -211 -23966 -177 -23932
rect -143 -23966 -109 -23932
rect 87 -23966 121 -23932
rect 155 -23966 189 -23932
rect 385 -23966 419 -23932
rect 453 -23966 487 -23932
rect 683 -23966 717 -23932
rect 751 -23966 785 -23932
rect 2851 -24014 2885 -23980
rect 2919 -24014 2953 -23980
rect 2987 -24014 3021 -23980
rect 3055 -24014 3089 -23980
rect 3123 -24014 3157 -23980
rect 3191 -24014 3225 -23980
rect 3259 -24014 3293 -23980
rect 3327 -24014 3361 -23980
rect 3869 -24014 3903 -23980
rect 3937 -24014 3971 -23980
rect 4005 -24014 4039 -23980
rect 4073 -24014 4107 -23980
rect 4141 -24014 4175 -23980
rect 4209 -24014 4243 -23980
rect 4277 -24014 4311 -23980
rect 4345 -24014 4379 -23980
rect 4887 -24014 4921 -23980
rect 4955 -24014 4989 -23980
rect 5023 -24014 5057 -23980
rect 5091 -24014 5125 -23980
rect 5159 -24014 5193 -23980
rect 5227 -24014 5261 -23980
rect 5295 -24014 5329 -23980
rect 5363 -24014 5397 -23980
rect 5905 -24014 5939 -23980
rect 5973 -24014 6007 -23980
rect 6041 -24014 6075 -23980
rect 6109 -24014 6143 -23980
rect 6177 -24014 6211 -23980
rect 6245 -24014 6279 -23980
rect 6313 -24014 6347 -23980
rect 6381 -24014 6415 -23980
rect 6923 -24014 6957 -23980
rect 6991 -24014 7025 -23980
rect 7059 -24014 7093 -23980
rect 7127 -24014 7161 -23980
rect 7195 -24014 7229 -23980
rect 7263 -24014 7297 -23980
rect 7331 -24014 7365 -23980
rect 7399 -24014 7433 -23980
rect 7941 -24014 7975 -23980
rect 8009 -24014 8043 -23980
rect 8077 -24014 8111 -23980
rect 8145 -24014 8179 -23980
rect 8213 -24014 8247 -23980
rect 8281 -24014 8315 -23980
rect 8349 -24014 8383 -23980
rect 8417 -24014 8451 -23980
rect 8959 -24014 8993 -23980
rect 9027 -24014 9061 -23980
rect 9095 -24014 9129 -23980
rect 9163 -24014 9197 -23980
rect 9231 -24014 9265 -23980
rect 9299 -24014 9333 -23980
rect 9367 -24014 9401 -23980
rect 9435 -24014 9469 -23980
rect 9977 -24014 10011 -23980
rect 10045 -24014 10079 -23980
rect 10113 -24014 10147 -23980
rect 10181 -24014 10215 -23980
rect 10249 -24014 10283 -23980
rect 10317 -24014 10351 -23980
rect 10385 -24014 10419 -23980
rect 10453 -24014 10487 -23980
rect 10995 -24014 11029 -23980
rect 11063 -24014 11097 -23980
rect 11131 -24014 11165 -23980
rect 11199 -24014 11233 -23980
rect 11267 -24014 11301 -23980
rect 11335 -24014 11369 -23980
rect 11403 -24014 11437 -23980
rect 11471 -24014 11505 -23980
rect 12013 -24014 12047 -23980
rect 12081 -24014 12115 -23980
rect 12149 -24014 12183 -23980
rect 12217 -24014 12251 -23980
rect 12285 -24014 12319 -23980
rect 12353 -24014 12387 -23980
rect 12421 -24014 12455 -23980
rect 12489 -24014 12523 -23980
rect 13031 -24014 13065 -23980
rect 13099 -24014 13133 -23980
rect 13167 -24014 13201 -23980
rect 13235 -24014 13269 -23980
rect 13303 -24014 13337 -23980
rect 13371 -24014 13405 -23980
rect 13439 -24014 13473 -23980
rect 13507 -24014 13541 -23980
rect 14049 -24014 14083 -23980
rect 14117 -24014 14151 -23980
rect 14185 -24014 14219 -23980
rect 14253 -24014 14287 -23980
rect 14321 -24014 14355 -23980
rect 14389 -24014 14423 -23980
rect 14457 -24014 14491 -23980
rect 14525 -24014 14559 -23980
rect 15067 -24014 15101 -23980
rect 15135 -24014 15169 -23980
rect 15203 -24014 15237 -23980
rect 15271 -24014 15305 -23980
rect 15339 -24014 15373 -23980
rect 15407 -24014 15441 -23980
rect 15475 -24014 15509 -23980
rect 15543 -24014 15577 -23980
rect 16085 -24014 16119 -23980
rect 16153 -24014 16187 -23980
rect 16221 -24014 16255 -23980
rect 16289 -24014 16323 -23980
rect 16357 -24014 16391 -23980
rect 16425 -24014 16459 -23980
rect 16493 -24014 16527 -23980
rect 16561 -24014 16595 -23980
rect 17103 -24014 17137 -23980
rect 17171 -24014 17205 -23980
rect 17239 -24014 17273 -23980
rect 17307 -24014 17341 -23980
rect 17375 -24014 17409 -23980
rect 17443 -24014 17477 -23980
rect 17511 -24014 17545 -23980
rect 17579 -24014 17613 -23980
rect 18121 -24014 18155 -23980
rect 18189 -24014 18223 -23980
rect 18257 -24014 18291 -23980
rect 18325 -24014 18359 -23980
rect 18393 -24014 18427 -23980
rect 18461 -24014 18495 -23980
rect 18529 -24014 18563 -23980
rect 18597 -24014 18631 -23980
rect 19139 -24014 19173 -23980
rect 19207 -24014 19241 -23980
rect 19275 -24014 19309 -23980
rect 19343 -24014 19377 -23980
rect 19411 -24014 19445 -23980
rect 19479 -24014 19513 -23980
rect 19547 -24014 19581 -23980
rect 19615 -24014 19649 -23980
rect 20157 -24014 20191 -23980
rect 20225 -24014 20259 -23980
rect 20293 -24014 20327 -23980
rect 20361 -24014 20395 -23980
rect 20429 -24014 20463 -23980
rect 20497 -24014 20531 -23980
rect 20565 -24014 20599 -23980
rect 20633 -24014 20667 -23980
rect 21175 -24014 21209 -23980
rect 21243 -24014 21277 -23980
rect 21311 -24014 21345 -23980
rect 21379 -24014 21413 -23980
rect 21447 -24014 21481 -23980
rect 21515 -24014 21549 -23980
rect 21583 -24014 21617 -23980
rect 21651 -24014 21685 -23980
rect 22193 -24014 22227 -23980
rect 22261 -24014 22295 -23980
rect 22329 -24014 22363 -23980
rect 22397 -24014 22431 -23980
rect 22465 -24014 22499 -23980
rect 22533 -24014 22567 -23980
rect 22601 -24014 22635 -23980
rect 22669 -24014 22703 -23980
rect -9134 -24677 -9100 -24643
rect -9066 -24677 -9032 -24643
rect -8998 -24677 -8964 -24643
rect -8930 -24677 -8896 -24643
rect -8862 -24677 -8828 -24643
rect -8794 -24677 -8760 -24643
rect -8726 -24677 -8692 -24643
rect -8658 -24677 -8624 -24643
rect -8116 -24677 -8082 -24643
rect -8048 -24677 -8014 -24643
rect -7980 -24677 -7946 -24643
rect -7912 -24677 -7878 -24643
rect -7844 -24677 -7810 -24643
rect -7776 -24677 -7742 -24643
rect -7708 -24677 -7674 -24643
rect -7640 -24677 -7606 -24643
rect -7098 -24677 -7064 -24643
rect -7030 -24677 -6996 -24643
rect -6962 -24677 -6928 -24643
rect -6894 -24677 -6860 -24643
rect -6826 -24677 -6792 -24643
rect -6758 -24677 -6724 -24643
rect -6690 -24677 -6656 -24643
rect -6622 -24677 -6588 -24643
rect -6080 -24677 -6046 -24643
rect -6012 -24677 -5978 -24643
rect -5944 -24677 -5910 -24643
rect -5876 -24677 -5842 -24643
rect -5808 -24677 -5774 -24643
rect -5740 -24677 -5706 -24643
rect -5672 -24677 -5638 -24643
rect -5604 -24677 -5570 -24643
rect -5062 -24677 -5028 -24643
rect -4994 -24677 -4960 -24643
rect -4926 -24677 -4892 -24643
rect -4858 -24677 -4824 -24643
rect -4790 -24677 -4756 -24643
rect -4722 -24677 -4688 -24643
rect -4654 -24677 -4620 -24643
rect -4586 -24677 -4552 -24643
rect -4044 -24677 -4010 -24643
rect -3976 -24677 -3942 -24643
rect -3908 -24677 -3874 -24643
rect -3840 -24677 -3806 -24643
rect -3772 -24677 -3738 -24643
rect -3704 -24677 -3670 -24643
rect -3636 -24677 -3602 -24643
rect -3568 -24677 -3534 -24643
rect -2297 -24676 -2263 -24642
rect -2229 -24676 -2195 -24642
rect -1999 -24676 -1965 -24642
rect -1931 -24676 -1897 -24642
rect -1701 -24676 -1667 -24642
rect -1633 -24676 -1599 -24642
rect -1403 -24676 -1369 -24642
rect -1335 -24676 -1301 -24642
rect -1105 -24676 -1071 -24642
rect -1037 -24676 -1003 -24642
rect -807 -24676 -773 -24642
rect -739 -24676 -705 -24642
rect -509 -24676 -475 -24642
rect -441 -24676 -407 -24642
rect -211 -24676 -177 -24642
rect -143 -24676 -109 -24642
rect 87 -24676 121 -24642
rect 155 -24676 189 -24642
rect 385 -24676 419 -24642
rect 453 -24676 487 -24642
rect 683 -24676 717 -24642
rect 751 -24676 785 -24642
rect 2851 -24724 2885 -24690
rect 2919 -24724 2953 -24690
rect 2987 -24724 3021 -24690
rect 3055 -24724 3089 -24690
rect 3123 -24724 3157 -24690
rect 3191 -24724 3225 -24690
rect 3259 -24724 3293 -24690
rect 3327 -24724 3361 -24690
rect 3869 -24724 3903 -24690
rect 3937 -24724 3971 -24690
rect 4005 -24724 4039 -24690
rect 4073 -24724 4107 -24690
rect 4141 -24724 4175 -24690
rect 4209 -24724 4243 -24690
rect 4277 -24724 4311 -24690
rect 4345 -24724 4379 -24690
rect 4887 -24724 4921 -24690
rect 4955 -24724 4989 -24690
rect 5023 -24724 5057 -24690
rect 5091 -24724 5125 -24690
rect 5159 -24724 5193 -24690
rect 5227 -24724 5261 -24690
rect 5295 -24724 5329 -24690
rect 5363 -24724 5397 -24690
rect 5905 -24724 5939 -24690
rect 5973 -24724 6007 -24690
rect 6041 -24724 6075 -24690
rect 6109 -24724 6143 -24690
rect 6177 -24724 6211 -24690
rect 6245 -24724 6279 -24690
rect 6313 -24724 6347 -24690
rect 6381 -24724 6415 -24690
rect 6923 -24724 6957 -24690
rect 6991 -24724 7025 -24690
rect 7059 -24724 7093 -24690
rect 7127 -24724 7161 -24690
rect 7195 -24724 7229 -24690
rect 7263 -24724 7297 -24690
rect 7331 -24724 7365 -24690
rect 7399 -24724 7433 -24690
rect 7941 -24724 7975 -24690
rect 8009 -24724 8043 -24690
rect 8077 -24724 8111 -24690
rect 8145 -24724 8179 -24690
rect 8213 -24724 8247 -24690
rect 8281 -24724 8315 -24690
rect 8349 -24724 8383 -24690
rect 8417 -24724 8451 -24690
rect 8959 -24724 8993 -24690
rect 9027 -24724 9061 -24690
rect 9095 -24724 9129 -24690
rect 9163 -24724 9197 -24690
rect 9231 -24724 9265 -24690
rect 9299 -24724 9333 -24690
rect 9367 -24724 9401 -24690
rect 9435 -24724 9469 -24690
rect 9977 -24724 10011 -24690
rect 10045 -24724 10079 -24690
rect 10113 -24724 10147 -24690
rect 10181 -24724 10215 -24690
rect 10249 -24724 10283 -24690
rect 10317 -24724 10351 -24690
rect 10385 -24724 10419 -24690
rect 10453 -24724 10487 -24690
rect 10995 -24724 11029 -24690
rect 11063 -24724 11097 -24690
rect 11131 -24724 11165 -24690
rect 11199 -24724 11233 -24690
rect 11267 -24724 11301 -24690
rect 11335 -24724 11369 -24690
rect 11403 -24724 11437 -24690
rect 11471 -24724 11505 -24690
rect 12013 -24724 12047 -24690
rect 12081 -24724 12115 -24690
rect 12149 -24724 12183 -24690
rect 12217 -24724 12251 -24690
rect 12285 -24724 12319 -24690
rect 12353 -24724 12387 -24690
rect 12421 -24724 12455 -24690
rect 12489 -24724 12523 -24690
rect 13031 -24724 13065 -24690
rect 13099 -24724 13133 -24690
rect 13167 -24724 13201 -24690
rect 13235 -24724 13269 -24690
rect 13303 -24724 13337 -24690
rect 13371 -24724 13405 -24690
rect 13439 -24724 13473 -24690
rect 13507 -24724 13541 -24690
rect 14049 -24724 14083 -24690
rect 14117 -24724 14151 -24690
rect 14185 -24724 14219 -24690
rect 14253 -24724 14287 -24690
rect 14321 -24724 14355 -24690
rect 14389 -24724 14423 -24690
rect 14457 -24724 14491 -24690
rect 14525 -24724 14559 -24690
rect 15067 -24724 15101 -24690
rect 15135 -24724 15169 -24690
rect 15203 -24724 15237 -24690
rect 15271 -24724 15305 -24690
rect 15339 -24724 15373 -24690
rect 15407 -24724 15441 -24690
rect 15475 -24724 15509 -24690
rect 15543 -24724 15577 -24690
rect 16085 -24724 16119 -24690
rect 16153 -24724 16187 -24690
rect 16221 -24724 16255 -24690
rect 16289 -24724 16323 -24690
rect 16357 -24724 16391 -24690
rect 16425 -24724 16459 -24690
rect 16493 -24724 16527 -24690
rect 16561 -24724 16595 -24690
rect 17103 -24724 17137 -24690
rect 17171 -24724 17205 -24690
rect 17239 -24724 17273 -24690
rect 17307 -24724 17341 -24690
rect 17375 -24724 17409 -24690
rect 17443 -24724 17477 -24690
rect 17511 -24724 17545 -24690
rect 17579 -24724 17613 -24690
rect 18121 -24724 18155 -24690
rect 18189 -24724 18223 -24690
rect 18257 -24724 18291 -24690
rect 18325 -24724 18359 -24690
rect 18393 -24724 18427 -24690
rect 18461 -24724 18495 -24690
rect 18529 -24724 18563 -24690
rect 18597 -24724 18631 -24690
rect 19139 -24724 19173 -24690
rect 19207 -24724 19241 -24690
rect 19275 -24724 19309 -24690
rect 19343 -24724 19377 -24690
rect 19411 -24724 19445 -24690
rect 19479 -24724 19513 -24690
rect 19547 -24724 19581 -24690
rect 19615 -24724 19649 -24690
rect 20157 -24724 20191 -24690
rect 20225 -24724 20259 -24690
rect 20293 -24724 20327 -24690
rect 20361 -24724 20395 -24690
rect 20429 -24724 20463 -24690
rect 20497 -24724 20531 -24690
rect 20565 -24724 20599 -24690
rect 20633 -24724 20667 -24690
rect 21175 -24724 21209 -24690
rect 21243 -24724 21277 -24690
rect 21311 -24724 21345 -24690
rect 21379 -24724 21413 -24690
rect 21447 -24724 21481 -24690
rect 21515 -24724 21549 -24690
rect 21583 -24724 21617 -24690
rect 21651 -24724 21685 -24690
rect 22193 -24724 22227 -24690
rect 22261 -24724 22295 -24690
rect 22329 -24724 22363 -24690
rect 22397 -24724 22431 -24690
rect 22465 -24724 22499 -24690
rect 22533 -24724 22567 -24690
rect 22601 -24724 22635 -24690
rect 22669 -24724 22703 -24690
rect -9135 -25080 -9101 -25046
rect -9067 -25080 -9033 -25046
rect -8999 -25080 -8965 -25046
rect -8931 -25080 -8897 -25046
rect -8863 -25080 -8829 -25046
rect -8795 -25080 -8761 -25046
rect -8727 -25080 -8693 -25046
rect -8659 -25080 -8625 -25046
rect -8117 -25080 -8083 -25046
rect -8049 -25080 -8015 -25046
rect -7981 -25080 -7947 -25046
rect -7913 -25080 -7879 -25046
rect -7845 -25080 -7811 -25046
rect -7777 -25080 -7743 -25046
rect -7709 -25080 -7675 -25046
rect -7641 -25080 -7607 -25046
rect -7099 -25080 -7065 -25046
rect -7031 -25080 -6997 -25046
rect -6963 -25080 -6929 -25046
rect -6895 -25080 -6861 -25046
rect -6827 -25080 -6793 -25046
rect -6759 -25080 -6725 -25046
rect -6691 -25080 -6657 -25046
rect -6623 -25080 -6589 -25046
rect -6081 -25080 -6047 -25046
rect -6013 -25080 -5979 -25046
rect -5945 -25080 -5911 -25046
rect -5877 -25080 -5843 -25046
rect -5809 -25080 -5775 -25046
rect -5741 -25080 -5707 -25046
rect -5673 -25080 -5639 -25046
rect -5605 -25080 -5571 -25046
rect -5063 -25080 -5029 -25046
rect -4995 -25080 -4961 -25046
rect -4927 -25080 -4893 -25046
rect -4859 -25080 -4825 -25046
rect -4791 -25080 -4757 -25046
rect -4723 -25080 -4689 -25046
rect -4655 -25080 -4621 -25046
rect -4587 -25080 -4553 -25046
rect -4045 -25080 -4011 -25046
rect -3977 -25080 -3943 -25046
rect -3909 -25080 -3875 -25046
rect -3841 -25080 -3807 -25046
rect -3773 -25080 -3739 -25046
rect -3705 -25080 -3671 -25046
rect -3637 -25080 -3603 -25046
rect -3569 -25080 -3535 -25046
rect -2297 -25076 -2263 -25042
rect -2229 -25076 -2195 -25042
rect -1999 -25076 -1965 -25042
rect -1931 -25076 -1897 -25042
rect -1701 -25076 -1667 -25042
rect -1633 -25076 -1599 -25042
rect -1403 -25076 -1369 -25042
rect -1335 -25076 -1301 -25042
rect -1105 -25076 -1071 -25042
rect -1037 -25076 -1003 -25042
rect -807 -25076 -773 -25042
rect -739 -25076 -705 -25042
rect -509 -25076 -475 -25042
rect -441 -25076 -407 -25042
rect -211 -25076 -177 -25042
rect -143 -25076 -109 -25042
rect 87 -25076 121 -25042
rect 155 -25076 189 -25042
rect 385 -25076 419 -25042
rect 453 -25076 487 -25042
rect 683 -25076 717 -25042
rect 751 -25076 785 -25042
rect 2851 -25246 2885 -25212
rect 2919 -25246 2953 -25212
rect 2987 -25246 3021 -25212
rect 3055 -25246 3089 -25212
rect 3123 -25246 3157 -25212
rect 3191 -25246 3225 -25212
rect 3259 -25246 3293 -25212
rect 3327 -25246 3361 -25212
rect 3869 -25246 3903 -25212
rect 3937 -25246 3971 -25212
rect 4005 -25246 4039 -25212
rect 4073 -25246 4107 -25212
rect 4141 -25246 4175 -25212
rect 4209 -25246 4243 -25212
rect 4277 -25246 4311 -25212
rect 4345 -25246 4379 -25212
rect 4887 -25246 4921 -25212
rect 4955 -25246 4989 -25212
rect 5023 -25246 5057 -25212
rect 5091 -25246 5125 -25212
rect 5159 -25246 5193 -25212
rect 5227 -25246 5261 -25212
rect 5295 -25246 5329 -25212
rect 5363 -25246 5397 -25212
rect 5905 -25246 5939 -25212
rect 5973 -25246 6007 -25212
rect 6041 -25246 6075 -25212
rect 6109 -25246 6143 -25212
rect 6177 -25246 6211 -25212
rect 6245 -25246 6279 -25212
rect 6313 -25246 6347 -25212
rect 6381 -25246 6415 -25212
rect 6923 -25246 6957 -25212
rect 6991 -25246 7025 -25212
rect 7059 -25246 7093 -25212
rect 7127 -25246 7161 -25212
rect 7195 -25246 7229 -25212
rect 7263 -25246 7297 -25212
rect 7331 -25246 7365 -25212
rect 7399 -25246 7433 -25212
rect 7941 -25246 7975 -25212
rect 8009 -25246 8043 -25212
rect 8077 -25246 8111 -25212
rect 8145 -25246 8179 -25212
rect 8213 -25246 8247 -25212
rect 8281 -25246 8315 -25212
rect 8349 -25246 8383 -25212
rect 8417 -25246 8451 -25212
rect 8959 -25246 8993 -25212
rect 9027 -25246 9061 -25212
rect 9095 -25246 9129 -25212
rect 9163 -25246 9197 -25212
rect 9231 -25246 9265 -25212
rect 9299 -25246 9333 -25212
rect 9367 -25246 9401 -25212
rect 9435 -25246 9469 -25212
rect 9977 -25246 10011 -25212
rect 10045 -25246 10079 -25212
rect 10113 -25246 10147 -25212
rect 10181 -25246 10215 -25212
rect 10249 -25246 10283 -25212
rect 10317 -25246 10351 -25212
rect 10385 -25246 10419 -25212
rect 10453 -25246 10487 -25212
rect 10995 -25246 11029 -25212
rect 11063 -25246 11097 -25212
rect 11131 -25246 11165 -25212
rect 11199 -25246 11233 -25212
rect 11267 -25246 11301 -25212
rect 11335 -25246 11369 -25212
rect 11403 -25246 11437 -25212
rect 11471 -25246 11505 -25212
rect 12013 -25246 12047 -25212
rect 12081 -25246 12115 -25212
rect 12149 -25246 12183 -25212
rect 12217 -25246 12251 -25212
rect 12285 -25246 12319 -25212
rect 12353 -25246 12387 -25212
rect 12421 -25246 12455 -25212
rect 12489 -25246 12523 -25212
rect 13031 -25246 13065 -25212
rect 13099 -25246 13133 -25212
rect 13167 -25246 13201 -25212
rect 13235 -25246 13269 -25212
rect 13303 -25246 13337 -25212
rect 13371 -25246 13405 -25212
rect 13439 -25246 13473 -25212
rect 13507 -25246 13541 -25212
rect 14049 -25246 14083 -25212
rect 14117 -25246 14151 -25212
rect 14185 -25246 14219 -25212
rect 14253 -25246 14287 -25212
rect 14321 -25246 14355 -25212
rect 14389 -25246 14423 -25212
rect 14457 -25246 14491 -25212
rect 14525 -25246 14559 -25212
rect 15067 -25246 15101 -25212
rect 15135 -25246 15169 -25212
rect 15203 -25246 15237 -25212
rect 15271 -25246 15305 -25212
rect 15339 -25246 15373 -25212
rect 15407 -25246 15441 -25212
rect 15475 -25246 15509 -25212
rect 15543 -25246 15577 -25212
rect 16085 -25246 16119 -25212
rect 16153 -25246 16187 -25212
rect 16221 -25246 16255 -25212
rect 16289 -25246 16323 -25212
rect 16357 -25246 16391 -25212
rect 16425 -25246 16459 -25212
rect 16493 -25246 16527 -25212
rect 16561 -25246 16595 -25212
rect 17103 -25246 17137 -25212
rect 17171 -25246 17205 -25212
rect 17239 -25246 17273 -25212
rect 17307 -25246 17341 -25212
rect 17375 -25246 17409 -25212
rect 17443 -25246 17477 -25212
rect 17511 -25246 17545 -25212
rect 17579 -25246 17613 -25212
rect 18121 -25246 18155 -25212
rect 18189 -25246 18223 -25212
rect 18257 -25246 18291 -25212
rect 18325 -25246 18359 -25212
rect 18393 -25246 18427 -25212
rect 18461 -25246 18495 -25212
rect 18529 -25246 18563 -25212
rect 18597 -25246 18631 -25212
rect 19139 -25246 19173 -25212
rect 19207 -25246 19241 -25212
rect 19275 -25246 19309 -25212
rect 19343 -25246 19377 -25212
rect 19411 -25246 19445 -25212
rect 19479 -25246 19513 -25212
rect 19547 -25246 19581 -25212
rect 19615 -25246 19649 -25212
rect 20157 -25246 20191 -25212
rect 20225 -25246 20259 -25212
rect 20293 -25246 20327 -25212
rect 20361 -25246 20395 -25212
rect 20429 -25246 20463 -25212
rect 20497 -25246 20531 -25212
rect 20565 -25246 20599 -25212
rect 20633 -25246 20667 -25212
rect 21175 -25246 21209 -25212
rect 21243 -25246 21277 -25212
rect 21311 -25246 21345 -25212
rect 21379 -25246 21413 -25212
rect 21447 -25246 21481 -25212
rect 21515 -25246 21549 -25212
rect 21583 -25246 21617 -25212
rect 21651 -25246 21685 -25212
rect 22193 -25246 22227 -25212
rect 22261 -25246 22295 -25212
rect 22329 -25246 22363 -25212
rect 22397 -25246 22431 -25212
rect 22465 -25246 22499 -25212
rect 22533 -25246 22567 -25212
rect 22601 -25246 22635 -25212
rect 22669 -25246 22703 -25212
rect -9135 -25790 -9101 -25756
rect -9067 -25790 -9033 -25756
rect -8999 -25790 -8965 -25756
rect -8931 -25790 -8897 -25756
rect -8863 -25790 -8829 -25756
rect -8795 -25790 -8761 -25756
rect -8727 -25790 -8693 -25756
rect -8659 -25790 -8625 -25756
rect -8117 -25790 -8083 -25756
rect -8049 -25790 -8015 -25756
rect -7981 -25790 -7947 -25756
rect -7913 -25790 -7879 -25756
rect -7845 -25790 -7811 -25756
rect -7777 -25790 -7743 -25756
rect -7709 -25790 -7675 -25756
rect -7641 -25790 -7607 -25756
rect -7099 -25790 -7065 -25756
rect -7031 -25790 -6997 -25756
rect -6963 -25790 -6929 -25756
rect -6895 -25790 -6861 -25756
rect -6827 -25790 -6793 -25756
rect -6759 -25790 -6725 -25756
rect -6691 -25790 -6657 -25756
rect -6623 -25790 -6589 -25756
rect -6081 -25790 -6047 -25756
rect -6013 -25790 -5979 -25756
rect -5945 -25790 -5911 -25756
rect -5877 -25790 -5843 -25756
rect -5809 -25790 -5775 -25756
rect -5741 -25790 -5707 -25756
rect -5673 -25790 -5639 -25756
rect -5605 -25790 -5571 -25756
rect -5063 -25790 -5029 -25756
rect -4995 -25790 -4961 -25756
rect -4927 -25790 -4893 -25756
rect -4859 -25790 -4825 -25756
rect -4791 -25790 -4757 -25756
rect -4723 -25790 -4689 -25756
rect -4655 -25790 -4621 -25756
rect -4587 -25790 -4553 -25756
rect -4045 -25790 -4011 -25756
rect -3977 -25790 -3943 -25756
rect -3909 -25790 -3875 -25756
rect -3841 -25790 -3807 -25756
rect -3773 -25790 -3739 -25756
rect -3705 -25790 -3671 -25756
rect -3637 -25790 -3603 -25756
rect -3569 -25790 -3535 -25756
rect -2297 -25786 -2263 -25752
rect -2229 -25786 -2195 -25752
rect -1999 -25786 -1965 -25752
rect -1931 -25786 -1897 -25752
rect -1701 -25786 -1667 -25752
rect -1633 -25786 -1599 -25752
rect -1403 -25786 -1369 -25752
rect -1335 -25786 -1301 -25752
rect -1105 -25786 -1071 -25752
rect -1037 -25786 -1003 -25752
rect -807 -25786 -773 -25752
rect -739 -25786 -705 -25752
rect -509 -25786 -475 -25752
rect -441 -25786 -407 -25752
rect -211 -25786 -177 -25752
rect -143 -25786 -109 -25752
rect 87 -25786 121 -25752
rect 155 -25786 189 -25752
rect 385 -25786 419 -25752
rect 453 -25786 487 -25752
rect 683 -25786 717 -25752
rect 751 -25786 785 -25752
rect 2851 -25956 2885 -25922
rect 2919 -25956 2953 -25922
rect 2987 -25956 3021 -25922
rect 3055 -25956 3089 -25922
rect 3123 -25956 3157 -25922
rect 3191 -25956 3225 -25922
rect 3259 -25956 3293 -25922
rect 3327 -25956 3361 -25922
rect 3869 -25956 3903 -25922
rect 3937 -25956 3971 -25922
rect 4005 -25956 4039 -25922
rect 4073 -25956 4107 -25922
rect 4141 -25956 4175 -25922
rect 4209 -25956 4243 -25922
rect 4277 -25956 4311 -25922
rect 4345 -25956 4379 -25922
rect 4887 -25956 4921 -25922
rect 4955 -25956 4989 -25922
rect 5023 -25956 5057 -25922
rect 5091 -25956 5125 -25922
rect 5159 -25956 5193 -25922
rect 5227 -25956 5261 -25922
rect 5295 -25956 5329 -25922
rect 5363 -25956 5397 -25922
rect 5905 -25956 5939 -25922
rect 5973 -25956 6007 -25922
rect 6041 -25956 6075 -25922
rect 6109 -25956 6143 -25922
rect 6177 -25956 6211 -25922
rect 6245 -25956 6279 -25922
rect 6313 -25956 6347 -25922
rect 6381 -25956 6415 -25922
rect 6923 -25956 6957 -25922
rect 6991 -25956 7025 -25922
rect 7059 -25956 7093 -25922
rect 7127 -25956 7161 -25922
rect 7195 -25956 7229 -25922
rect 7263 -25956 7297 -25922
rect 7331 -25956 7365 -25922
rect 7399 -25956 7433 -25922
rect 7941 -25956 7975 -25922
rect 8009 -25956 8043 -25922
rect 8077 -25956 8111 -25922
rect 8145 -25956 8179 -25922
rect 8213 -25956 8247 -25922
rect 8281 -25956 8315 -25922
rect 8349 -25956 8383 -25922
rect 8417 -25956 8451 -25922
rect 8959 -25956 8993 -25922
rect 9027 -25956 9061 -25922
rect 9095 -25956 9129 -25922
rect 9163 -25956 9197 -25922
rect 9231 -25956 9265 -25922
rect 9299 -25956 9333 -25922
rect 9367 -25956 9401 -25922
rect 9435 -25956 9469 -25922
rect 9977 -25956 10011 -25922
rect 10045 -25956 10079 -25922
rect 10113 -25956 10147 -25922
rect 10181 -25956 10215 -25922
rect 10249 -25956 10283 -25922
rect 10317 -25956 10351 -25922
rect 10385 -25956 10419 -25922
rect 10453 -25956 10487 -25922
rect 10995 -25956 11029 -25922
rect 11063 -25956 11097 -25922
rect 11131 -25956 11165 -25922
rect 11199 -25956 11233 -25922
rect 11267 -25956 11301 -25922
rect 11335 -25956 11369 -25922
rect 11403 -25956 11437 -25922
rect 11471 -25956 11505 -25922
rect 12013 -25956 12047 -25922
rect 12081 -25956 12115 -25922
rect 12149 -25956 12183 -25922
rect 12217 -25956 12251 -25922
rect 12285 -25956 12319 -25922
rect 12353 -25956 12387 -25922
rect 12421 -25956 12455 -25922
rect 12489 -25956 12523 -25922
rect 13031 -25956 13065 -25922
rect 13099 -25956 13133 -25922
rect 13167 -25956 13201 -25922
rect 13235 -25956 13269 -25922
rect 13303 -25956 13337 -25922
rect 13371 -25956 13405 -25922
rect 13439 -25956 13473 -25922
rect 13507 -25956 13541 -25922
rect 14049 -25956 14083 -25922
rect 14117 -25956 14151 -25922
rect 14185 -25956 14219 -25922
rect 14253 -25956 14287 -25922
rect 14321 -25956 14355 -25922
rect 14389 -25956 14423 -25922
rect 14457 -25956 14491 -25922
rect 14525 -25956 14559 -25922
rect 15067 -25956 15101 -25922
rect 15135 -25956 15169 -25922
rect 15203 -25956 15237 -25922
rect 15271 -25956 15305 -25922
rect 15339 -25956 15373 -25922
rect 15407 -25956 15441 -25922
rect 15475 -25956 15509 -25922
rect 15543 -25956 15577 -25922
rect 16085 -25956 16119 -25922
rect 16153 -25956 16187 -25922
rect 16221 -25956 16255 -25922
rect 16289 -25956 16323 -25922
rect 16357 -25956 16391 -25922
rect 16425 -25956 16459 -25922
rect 16493 -25956 16527 -25922
rect 16561 -25956 16595 -25922
rect 17103 -25956 17137 -25922
rect 17171 -25956 17205 -25922
rect 17239 -25956 17273 -25922
rect 17307 -25956 17341 -25922
rect 17375 -25956 17409 -25922
rect 17443 -25956 17477 -25922
rect 17511 -25956 17545 -25922
rect 17579 -25956 17613 -25922
rect 18121 -25956 18155 -25922
rect 18189 -25956 18223 -25922
rect 18257 -25956 18291 -25922
rect 18325 -25956 18359 -25922
rect 18393 -25956 18427 -25922
rect 18461 -25956 18495 -25922
rect 18529 -25956 18563 -25922
rect 18597 -25956 18631 -25922
rect 19139 -25956 19173 -25922
rect 19207 -25956 19241 -25922
rect 19275 -25956 19309 -25922
rect 19343 -25956 19377 -25922
rect 19411 -25956 19445 -25922
rect 19479 -25956 19513 -25922
rect 19547 -25956 19581 -25922
rect 19615 -25956 19649 -25922
rect 20157 -25956 20191 -25922
rect 20225 -25956 20259 -25922
rect 20293 -25956 20327 -25922
rect 20361 -25956 20395 -25922
rect 20429 -25956 20463 -25922
rect 20497 -25956 20531 -25922
rect 20565 -25956 20599 -25922
rect 20633 -25956 20667 -25922
rect 21175 -25956 21209 -25922
rect 21243 -25956 21277 -25922
rect 21311 -25956 21345 -25922
rect 21379 -25956 21413 -25922
rect 21447 -25956 21481 -25922
rect 21515 -25956 21549 -25922
rect 21583 -25956 21617 -25922
rect 21651 -25956 21685 -25922
rect 22193 -25956 22227 -25922
rect 22261 -25956 22295 -25922
rect 22329 -25956 22363 -25922
rect 22397 -25956 22431 -25922
rect 22465 -25956 22499 -25922
rect 22533 -25956 22567 -25922
rect 22601 -25956 22635 -25922
rect 22669 -25956 22703 -25922
<< locali >>
rect 378 1689 24822 1722
rect 378 1655 487 1689
rect 521 1655 547 1689
rect 593 1655 615 1689
rect 665 1655 683 1689
rect 737 1655 751 1689
rect 809 1655 819 1689
rect 881 1655 887 1689
rect 953 1655 955 1689
rect 989 1655 991 1689
rect 1057 1655 1063 1689
rect 1125 1655 1135 1689
rect 1193 1655 1207 1689
rect 1261 1655 1279 1689
rect 1329 1655 1351 1689
rect 1397 1655 1423 1689
rect 1465 1655 1495 1689
rect 1533 1655 1567 1689
rect 1601 1655 1635 1689
rect 1673 1655 1703 1689
rect 1745 1655 1771 1689
rect 1817 1655 1839 1689
rect 1889 1655 1907 1689
rect 1961 1655 1975 1689
rect 2033 1655 2043 1689
rect 2105 1655 2111 1689
rect 2177 1655 2179 1689
rect 2213 1655 2215 1689
rect 2281 1655 2287 1689
rect 2349 1655 2359 1689
rect 2417 1655 2431 1689
rect 2485 1655 2503 1689
rect 2553 1655 2575 1689
rect 2621 1655 2647 1689
rect 2689 1655 2719 1689
rect 2757 1655 2791 1689
rect 2825 1655 2859 1689
rect 2897 1655 2927 1689
rect 2969 1655 2995 1689
rect 3041 1655 3063 1689
rect 3113 1655 3131 1689
rect 3185 1655 3199 1689
rect 3257 1655 3267 1689
rect 3329 1655 3335 1689
rect 3401 1655 3403 1689
rect 3437 1655 3439 1689
rect 3505 1655 3511 1689
rect 3573 1655 3583 1689
rect 3641 1655 3655 1689
rect 3709 1655 3727 1689
rect 3777 1655 3799 1689
rect 3845 1655 3871 1689
rect 3913 1655 3943 1689
rect 3981 1655 4015 1689
rect 4049 1655 4083 1689
rect 4121 1655 4151 1689
rect 4193 1655 4219 1689
rect 4265 1655 4287 1689
rect 4337 1655 4355 1689
rect 4409 1655 4423 1689
rect 4481 1655 4491 1689
rect 4553 1655 4559 1689
rect 4625 1655 4627 1689
rect 4661 1655 4663 1689
rect 4729 1655 4735 1689
rect 4797 1655 4807 1689
rect 4865 1655 4879 1689
rect 4933 1655 4951 1689
rect 5001 1655 5023 1689
rect 5069 1655 5095 1689
rect 5137 1655 5167 1689
rect 5205 1655 5239 1689
rect 5273 1655 5307 1689
rect 5345 1655 5375 1689
rect 5417 1655 5443 1689
rect 5489 1655 5511 1689
rect 5561 1655 5579 1689
rect 5633 1655 5647 1689
rect 5705 1655 5715 1689
rect 5777 1655 5783 1689
rect 5849 1655 5851 1689
rect 5885 1655 5887 1689
rect 5953 1655 5959 1689
rect 6021 1655 6031 1689
rect 6089 1655 6103 1689
rect 6157 1655 6175 1689
rect 6225 1655 6247 1689
rect 6293 1655 6319 1689
rect 6361 1655 6391 1689
rect 6429 1655 6463 1689
rect 6497 1655 6531 1689
rect 6569 1655 6599 1689
rect 6641 1655 6667 1689
rect 6713 1655 6735 1689
rect 6785 1655 6803 1689
rect 6857 1655 6871 1689
rect 6929 1655 6939 1689
rect 7001 1655 7007 1689
rect 7073 1655 7075 1689
rect 7109 1655 7111 1689
rect 7177 1655 7183 1689
rect 7245 1655 7255 1689
rect 7313 1655 7327 1689
rect 7381 1655 7399 1689
rect 7449 1655 7471 1689
rect 7517 1655 7543 1689
rect 7585 1655 7615 1689
rect 7653 1655 7687 1689
rect 7721 1655 7755 1689
rect 7793 1655 7823 1689
rect 7865 1655 7891 1689
rect 7937 1655 7959 1689
rect 8009 1655 8027 1689
rect 8081 1655 8095 1689
rect 8153 1655 8163 1689
rect 8225 1655 8231 1689
rect 8297 1655 8299 1689
rect 8333 1655 8335 1689
rect 8401 1655 8407 1689
rect 8469 1655 8479 1689
rect 8537 1655 8551 1689
rect 8605 1655 8623 1689
rect 8673 1655 8695 1689
rect 8741 1655 8767 1689
rect 8809 1655 8839 1689
rect 8877 1655 8911 1689
rect 8945 1655 8979 1689
rect 9017 1655 9047 1689
rect 9089 1655 9115 1689
rect 9161 1655 9183 1689
rect 9233 1655 9251 1689
rect 9305 1655 9319 1689
rect 9377 1655 9387 1689
rect 9449 1655 9455 1689
rect 9521 1655 9523 1689
rect 9557 1655 9559 1689
rect 9625 1655 9631 1689
rect 9693 1655 9703 1689
rect 9761 1655 9775 1689
rect 9829 1655 9847 1689
rect 9897 1655 9919 1689
rect 9965 1655 9991 1689
rect 10033 1655 10063 1689
rect 10101 1655 10135 1689
rect 10169 1655 10203 1689
rect 10241 1655 10271 1689
rect 10313 1655 10339 1689
rect 10385 1655 10407 1689
rect 10457 1655 10475 1689
rect 10529 1655 10543 1689
rect 10601 1655 10611 1689
rect 10673 1655 10679 1689
rect 10745 1655 10747 1689
rect 10781 1655 10783 1689
rect 10849 1655 10855 1689
rect 10917 1655 10927 1689
rect 10985 1655 10999 1689
rect 11053 1655 11071 1689
rect 11121 1655 11143 1689
rect 11189 1655 11215 1689
rect 11257 1655 11287 1689
rect 11325 1655 11359 1689
rect 11393 1655 11427 1689
rect 11465 1655 11495 1689
rect 11537 1655 11563 1689
rect 11609 1655 11631 1689
rect 11681 1655 11699 1689
rect 11753 1655 11767 1689
rect 11825 1655 11835 1689
rect 11897 1655 11903 1689
rect 11969 1655 11971 1689
rect 12005 1655 12007 1689
rect 12073 1655 12079 1689
rect 12141 1655 12151 1689
rect 12209 1655 12223 1689
rect 12277 1655 12295 1689
rect 12345 1655 12367 1689
rect 12413 1655 12439 1689
rect 12481 1655 12511 1689
rect 12549 1655 12583 1689
rect 12617 1655 12651 1689
rect 12689 1655 12719 1689
rect 12761 1655 12787 1689
rect 12833 1655 12855 1689
rect 12905 1655 12923 1689
rect 12977 1655 12991 1689
rect 13049 1655 13059 1689
rect 13121 1655 13127 1689
rect 13193 1655 13195 1689
rect 13229 1655 13231 1689
rect 13297 1655 13303 1689
rect 13365 1655 13375 1689
rect 13433 1655 13447 1689
rect 13501 1655 13519 1689
rect 13569 1655 13591 1689
rect 13637 1655 13663 1689
rect 13705 1655 13735 1689
rect 13773 1655 13807 1689
rect 13841 1655 13875 1689
rect 13913 1655 13943 1689
rect 13985 1655 14011 1689
rect 14057 1655 14079 1689
rect 14129 1655 14147 1689
rect 14201 1655 14215 1689
rect 14273 1655 14283 1689
rect 14345 1655 14351 1689
rect 14417 1655 14419 1689
rect 14453 1655 14455 1689
rect 14521 1655 14527 1689
rect 14589 1655 14599 1689
rect 14657 1655 14671 1689
rect 14725 1655 14743 1689
rect 14793 1655 14815 1689
rect 14861 1655 14887 1689
rect 14929 1655 14959 1689
rect 14997 1655 15031 1689
rect 15065 1655 15099 1689
rect 15137 1655 15167 1689
rect 15209 1655 15235 1689
rect 15281 1655 15303 1689
rect 15353 1655 15371 1689
rect 15425 1655 15439 1689
rect 15497 1655 15507 1689
rect 15569 1655 15575 1689
rect 15641 1655 15643 1689
rect 15677 1655 15679 1689
rect 15745 1655 15751 1689
rect 15813 1655 15823 1689
rect 15881 1655 15895 1689
rect 15949 1655 15967 1689
rect 16017 1655 16039 1689
rect 16085 1655 16111 1689
rect 16153 1655 16183 1689
rect 16221 1655 16255 1689
rect 16289 1655 16323 1689
rect 16361 1655 16391 1689
rect 16433 1655 16459 1689
rect 16505 1655 16527 1689
rect 16577 1655 16595 1689
rect 16649 1655 16663 1689
rect 16721 1655 16731 1689
rect 16793 1655 16799 1689
rect 16865 1655 16867 1689
rect 16901 1655 16903 1689
rect 16969 1655 16975 1689
rect 17037 1655 17047 1689
rect 17105 1655 17119 1689
rect 17173 1655 17191 1689
rect 17241 1655 17263 1689
rect 17309 1655 17335 1689
rect 17377 1655 17407 1689
rect 17445 1655 17479 1689
rect 17513 1655 17547 1689
rect 17585 1655 17615 1689
rect 17657 1655 17683 1689
rect 17729 1655 17751 1689
rect 17801 1655 17819 1689
rect 17873 1655 17887 1689
rect 17945 1655 17955 1689
rect 18017 1655 18023 1689
rect 18089 1655 18091 1689
rect 18125 1655 18127 1689
rect 18193 1655 18199 1689
rect 18261 1655 18271 1689
rect 18329 1655 18343 1689
rect 18397 1655 18415 1689
rect 18465 1655 18487 1689
rect 18533 1655 18559 1689
rect 18601 1655 18631 1689
rect 18669 1655 18703 1689
rect 18737 1655 18771 1689
rect 18809 1655 18839 1689
rect 18881 1655 18907 1689
rect 18953 1655 18975 1689
rect 19025 1655 19043 1689
rect 19097 1655 19111 1689
rect 19169 1655 19179 1689
rect 19241 1655 19247 1689
rect 19313 1655 19315 1689
rect 19349 1655 19351 1689
rect 19417 1655 19423 1689
rect 19485 1655 19495 1689
rect 19553 1655 19567 1689
rect 19621 1655 19639 1689
rect 19689 1655 19711 1689
rect 19757 1655 19783 1689
rect 19825 1655 19855 1689
rect 19893 1655 19927 1689
rect 19961 1655 19995 1689
rect 20033 1655 20063 1689
rect 20105 1655 20131 1689
rect 20177 1655 20199 1689
rect 20249 1655 20267 1689
rect 20321 1655 20335 1689
rect 20393 1655 20403 1689
rect 20465 1655 20471 1689
rect 20537 1655 20539 1689
rect 20573 1655 20575 1689
rect 20641 1655 20647 1689
rect 20709 1655 20719 1689
rect 20777 1655 20791 1689
rect 20845 1655 20863 1689
rect 20913 1655 20935 1689
rect 20981 1655 21007 1689
rect 21049 1655 21079 1689
rect 21117 1655 21151 1689
rect 21185 1655 21219 1689
rect 21257 1655 21287 1689
rect 21329 1655 21355 1689
rect 21401 1655 21423 1689
rect 21473 1655 21491 1689
rect 21545 1655 21559 1689
rect 21617 1655 21627 1689
rect 21689 1655 21695 1689
rect 21761 1655 21763 1689
rect 21797 1655 21799 1689
rect 21865 1655 21871 1689
rect 21933 1655 21943 1689
rect 22001 1655 22015 1689
rect 22069 1655 22087 1689
rect 22137 1655 22159 1689
rect 22205 1655 22231 1689
rect 22273 1655 22303 1689
rect 22341 1655 22375 1689
rect 22409 1655 22443 1689
rect 22481 1655 22511 1689
rect 22553 1655 22579 1689
rect 22625 1655 22647 1689
rect 22697 1655 22715 1689
rect 22769 1655 22783 1689
rect 22841 1655 22851 1689
rect 22913 1655 22919 1689
rect 22985 1655 22987 1689
rect 23021 1655 23023 1689
rect 23089 1655 23095 1689
rect 23157 1655 23167 1689
rect 23225 1655 23239 1689
rect 23293 1655 23311 1689
rect 23361 1655 23383 1689
rect 23429 1655 23455 1689
rect 23497 1655 23527 1689
rect 23565 1655 23599 1689
rect 23633 1655 23667 1689
rect 23705 1655 23735 1689
rect 23777 1655 23803 1689
rect 23849 1655 23871 1689
rect 23921 1655 23939 1689
rect 23993 1655 24007 1689
rect 24065 1655 24075 1689
rect 24137 1655 24143 1689
rect 24209 1655 24211 1689
rect 24245 1655 24247 1689
rect 24313 1655 24319 1689
rect 24381 1655 24391 1689
rect 24449 1655 24463 1689
rect 24517 1655 24535 1689
rect 24585 1655 24607 1689
rect 24653 1655 24679 1689
rect 24713 1655 24822 1689
rect 378 1622 24822 1655
rect 378 1537 478 1622
rect 378 1503 411 1537
rect 445 1503 478 1537
rect 378 1469 478 1503
rect 378 1435 411 1469
rect 445 1435 478 1469
rect 378 1401 478 1435
rect 378 1367 411 1401
rect 445 1367 478 1401
rect 378 1333 478 1367
rect 378 1299 411 1333
rect 445 1299 478 1333
rect 378 1265 478 1299
rect 378 1231 411 1265
rect 445 1231 478 1265
rect 378 1197 478 1231
rect 378 1163 411 1197
rect 445 1163 478 1197
rect 378 1129 478 1163
rect 378 1095 411 1129
rect 445 1095 478 1129
rect 378 1081 478 1095
rect 378 1027 411 1081
rect 445 1027 478 1081
rect 378 1009 478 1027
rect 378 959 411 1009
rect 445 959 478 1009
rect 378 937 478 959
rect 378 891 411 937
rect 445 891 478 937
rect 378 865 478 891
rect 378 823 411 865
rect 445 823 478 865
rect 378 793 478 823
rect 378 755 411 793
rect 445 755 478 793
rect 378 721 478 755
rect 378 687 411 721
rect 445 687 478 721
rect 378 653 478 687
rect 378 615 411 653
rect 445 615 478 653
rect 378 585 478 615
rect 378 543 411 585
rect 445 543 478 585
rect 378 517 478 543
rect 378 471 411 517
rect 445 471 478 517
rect 378 449 478 471
rect 378 399 411 449
rect 445 399 478 449
rect 378 381 478 399
rect 378 327 411 381
rect 445 327 478 381
rect 378 313 478 327
rect 378 255 411 313
rect 445 255 478 313
rect 378 245 478 255
rect 378 183 411 245
rect 445 183 478 245
rect 378 177 478 183
rect 378 111 411 177
rect 445 111 478 177
rect 378 109 478 111
rect 378 75 411 109
rect 445 75 478 109
rect 378 73 478 75
rect 378 7 411 73
rect 445 7 478 73
rect 378 1 478 7
rect 378 -61 411 1
rect 445 -61 478 1
rect 378 -71 478 -61
rect 378 -129 411 -71
rect 445 -129 478 -71
rect 378 -143 478 -129
rect 378 -197 411 -143
rect 445 -197 478 -143
rect 378 -215 478 -197
rect 378 -265 411 -215
rect 445 -265 478 -215
rect 378 -287 478 -265
rect 378 -333 411 -287
rect 445 -333 478 -287
rect 378 -359 478 -333
rect 378 -401 411 -359
rect 445 -401 478 -359
rect 378 -431 478 -401
rect 378 -469 411 -431
rect 445 -469 478 -431
rect 378 -503 478 -469
rect 378 -537 411 -503
rect 445 -537 478 -503
rect 378 -571 478 -537
rect 378 -609 411 -571
rect 445 -609 478 -571
rect 378 -639 478 -609
rect 378 -681 411 -639
rect 445 -681 478 -639
rect 378 -707 478 -681
rect 378 -753 411 -707
rect 445 -753 478 -707
rect 378 -775 478 -753
rect 378 -825 411 -775
rect 445 -825 478 -775
rect 378 -843 478 -825
rect 378 -897 411 -843
rect 445 -897 478 -843
rect 378 -911 478 -897
rect 378 -969 411 -911
rect 445 -969 478 -911
rect 378 -979 478 -969
rect 378 -1041 411 -979
rect 445 -1041 478 -979
rect 378 -1047 478 -1041
rect 378 -1113 411 -1047
rect 445 -1113 478 -1047
rect 378 -1115 478 -1113
rect 378 -1149 411 -1115
rect 445 -1149 478 -1115
rect 378 -1151 478 -1149
rect 378 -1217 411 -1151
rect 445 -1217 478 -1151
rect 378 -1223 478 -1217
rect 378 -1285 411 -1223
rect 445 -1285 478 -1223
rect 378 -1295 478 -1285
rect 378 -1353 411 -1295
rect 445 -1353 478 -1295
rect 378 -1367 478 -1353
rect 378 -1421 411 -1367
rect 445 -1421 478 -1367
rect 378 -1439 478 -1421
rect 378 -1489 411 -1439
rect 445 -1489 478 -1439
rect 378 -1511 478 -1489
rect 378 -1557 411 -1511
rect 445 -1557 478 -1511
rect 378 -1583 478 -1557
rect 378 -1625 411 -1583
rect 445 -1625 478 -1583
rect 378 -1655 478 -1625
rect 378 -1693 411 -1655
rect 445 -1693 478 -1655
rect 378 -1727 478 -1693
rect 378 -1761 411 -1727
rect 445 -1761 478 -1727
rect 378 -1795 478 -1761
rect 378 -1833 411 -1795
rect 445 -1833 478 -1795
rect 378 -1863 478 -1833
rect 378 -1905 411 -1863
rect 445 -1905 478 -1863
rect 378 -1931 478 -1905
rect 378 -1977 411 -1931
rect 445 -1977 478 -1931
rect 378 -1999 478 -1977
rect 378 -2049 411 -1999
rect 445 -2049 478 -1999
rect 378 -2067 478 -2049
rect 378 -2121 411 -2067
rect 445 -2121 478 -2067
rect 378 -2135 478 -2121
rect 378 -2193 411 -2135
rect 445 -2193 478 -2135
rect 378 -2203 478 -2193
rect 378 -2265 411 -2203
rect 445 -2265 478 -2203
rect 378 -2271 478 -2265
rect 378 -2337 411 -2271
rect 445 -2337 478 -2271
rect 378 -2339 478 -2337
rect 378 -2373 411 -2339
rect 445 -2373 478 -2339
rect 378 -2375 478 -2373
rect 378 -2441 411 -2375
rect 445 -2441 478 -2375
rect 378 -2447 478 -2441
rect 378 -2509 411 -2447
rect 445 -2509 478 -2447
rect 378 -2519 478 -2509
rect 378 -2577 411 -2519
rect 445 -2577 478 -2519
rect 378 -2591 478 -2577
rect 378 -2645 411 -2591
rect 445 -2645 478 -2591
rect 378 -2663 478 -2645
rect 378 -2713 411 -2663
rect 445 -2713 478 -2663
rect 378 -2735 478 -2713
rect 378 -2781 411 -2735
rect 445 -2781 478 -2735
rect 378 -2807 478 -2781
rect 378 -2849 411 -2807
rect 445 -2849 478 -2807
rect 378 -2879 478 -2849
rect 378 -2917 411 -2879
rect 445 -2917 478 -2879
rect 378 -2951 478 -2917
rect 378 -2985 411 -2951
rect 445 -2985 478 -2951
rect 378 -3019 478 -2985
rect 378 -3057 411 -3019
rect 445 -3057 478 -3019
rect 378 -3087 478 -3057
rect 378 -3129 411 -3087
rect 445 -3129 478 -3087
rect 378 -3155 478 -3129
rect 378 -3201 411 -3155
rect 445 -3201 478 -3155
rect 378 -3223 478 -3201
rect 378 -3273 411 -3223
rect 445 -3273 478 -3223
rect 378 -3291 478 -3273
rect 378 -3345 411 -3291
rect 445 -3345 478 -3291
rect 378 -3359 478 -3345
rect 378 -3417 411 -3359
rect 445 -3417 478 -3359
rect 378 -3427 478 -3417
rect 378 -3489 411 -3427
rect 445 -3489 478 -3427
rect 378 -3495 478 -3489
rect 378 -3561 411 -3495
rect 445 -3561 478 -3495
rect 378 -3563 478 -3561
rect 378 -3597 411 -3563
rect 445 -3597 478 -3563
rect 378 -3599 478 -3597
rect 378 -3665 411 -3599
rect 445 -3665 478 -3599
rect 378 -3671 478 -3665
rect 378 -3733 411 -3671
rect 445 -3733 478 -3671
rect 378 -3743 478 -3733
rect 378 -3801 411 -3743
rect 445 -3801 478 -3743
rect 378 -3815 478 -3801
rect 378 -3869 411 -3815
rect 445 -3869 478 -3815
rect 378 -3887 478 -3869
rect 378 -3937 411 -3887
rect 445 -3937 478 -3887
rect 378 -3959 478 -3937
rect 378 -4005 411 -3959
rect 445 -4005 478 -3959
rect 378 -4031 478 -4005
rect 378 -4073 411 -4031
rect 445 -4073 478 -4031
rect 378 -4103 478 -4073
rect 378 -4141 411 -4103
rect 445 -4141 478 -4103
rect 378 -4175 478 -4141
rect 378 -4209 411 -4175
rect 445 -4209 478 -4175
rect 378 -4243 478 -4209
rect 378 -4281 411 -4243
rect 445 -4281 478 -4243
rect 378 -4311 478 -4281
rect 378 -4353 411 -4311
rect 445 -4353 478 -4311
rect 378 -4379 478 -4353
rect 378 -4425 411 -4379
rect 445 -4425 478 -4379
rect 378 -4447 478 -4425
rect 378 -4497 411 -4447
rect 445 -4497 478 -4447
rect 378 -4515 478 -4497
rect 378 -4569 411 -4515
rect 445 -4569 478 -4515
rect 378 -4583 478 -4569
rect 378 -4641 411 -4583
rect 445 -4641 478 -4583
rect 24722 1537 24822 1622
rect 24722 1503 24755 1537
rect 24789 1503 24822 1537
rect 24722 1469 24822 1503
rect 24722 1435 24755 1469
rect 24789 1435 24822 1469
rect 24722 1401 24822 1435
rect 24722 1367 24755 1401
rect 24789 1367 24822 1401
rect 24722 1333 24822 1367
rect 24722 1299 24755 1333
rect 24789 1299 24822 1333
rect 24722 1265 24822 1299
rect 24722 1231 24755 1265
rect 24789 1231 24822 1265
rect 24722 1197 24822 1231
rect 24722 1163 24755 1197
rect 24789 1163 24822 1197
rect 24722 1129 24822 1163
rect 24722 1095 24755 1129
rect 24789 1095 24822 1129
rect 24722 1081 24822 1095
rect 24722 1027 24755 1081
rect 24789 1027 24822 1081
rect 24722 1009 24822 1027
rect 24722 959 24755 1009
rect 24789 959 24822 1009
rect 24722 937 24822 959
rect 24722 891 24755 937
rect 24789 891 24822 937
rect 24722 865 24822 891
rect 24722 823 24755 865
rect 24789 823 24822 865
rect 24722 793 24822 823
rect 24722 755 24755 793
rect 24789 755 24822 793
rect 24722 721 24822 755
rect 24722 687 24755 721
rect 24789 687 24822 721
rect 24722 653 24822 687
rect 24722 615 24755 653
rect 24789 615 24822 653
rect 24722 585 24822 615
rect 24722 543 24755 585
rect 24789 543 24822 585
rect 24722 517 24822 543
rect 24722 471 24755 517
rect 24789 471 24822 517
rect 24722 449 24822 471
rect 24722 399 24755 449
rect 24789 399 24822 449
rect 24722 381 24822 399
rect 24722 327 24755 381
rect 24789 327 24822 381
rect 24722 313 24822 327
rect 24722 255 24755 313
rect 24789 255 24822 313
rect 24722 245 24822 255
rect 24722 183 24755 245
rect 24789 183 24822 245
rect 24722 177 24822 183
rect 24722 111 24755 177
rect 24789 111 24822 177
rect 24722 109 24822 111
rect 24722 75 24755 109
rect 24789 75 24822 109
rect 24722 73 24822 75
rect 24722 7 24755 73
rect 24789 7 24822 73
rect 24722 1 24822 7
rect 24722 -61 24755 1
rect 24789 -61 24822 1
rect 24722 -71 24822 -61
rect 24722 -129 24755 -71
rect 24789 -129 24822 -71
rect 24722 -143 24822 -129
rect 24722 -197 24755 -143
rect 24789 -197 24822 -143
rect 24722 -215 24822 -197
rect 24722 -265 24755 -215
rect 24789 -265 24822 -215
rect 24722 -287 24822 -265
rect 24722 -333 24755 -287
rect 24789 -333 24822 -287
rect 24722 -359 24822 -333
rect 24722 -401 24755 -359
rect 24789 -401 24822 -359
rect 24722 -431 24822 -401
rect 24722 -469 24755 -431
rect 24789 -469 24822 -431
rect 24722 -503 24822 -469
rect 24722 -537 24755 -503
rect 24789 -537 24822 -503
rect 24722 -571 24822 -537
rect 24722 -609 24755 -571
rect 24789 -609 24822 -571
rect 24722 -639 24822 -609
rect 24722 -681 24755 -639
rect 24789 -681 24822 -639
rect 24722 -707 24822 -681
rect 24722 -753 24755 -707
rect 24789 -753 24822 -707
rect 24722 -775 24822 -753
rect 24722 -825 24755 -775
rect 24789 -825 24822 -775
rect 24722 -843 24822 -825
rect 24722 -897 24755 -843
rect 24789 -897 24822 -843
rect 24722 -911 24822 -897
rect 24722 -969 24755 -911
rect 24789 -969 24822 -911
rect 24722 -979 24822 -969
rect 24722 -1041 24755 -979
rect 24789 -1041 24822 -979
rect 24722 -1047 24822 -1041
rect 24722 -1113 24755 -1047
rect 24789 -1113 24822 -1047
rect 24722 -1115 24822 -1113
rect 24722 -1149 24755 -1115
rect 24789 -1149 24822 -1115
rect 24722 -1151 24822 -1149
rect 24722 -1217 24755 -1151
rect 24789 -1217 24822 -1151
rect 24722 -1223 24822 -1217
rect 24722 -1285 24755 -1223
rect 24789 -1285 24822 -1223
rect 24722 -1295 24822 -1285
rect 24722 -1353 24755 -1295
rect 24789 -1353 24822 -1295
rect 24722 -1367 24822 -1353
rect 24722 -1421 24755 -1367
rect 24789 -1421 24822 -1367
rect 24722 -1439 24822 -1421
rect 24722 -1489 24755 -1439
rect 24789 -1489 24822 -1439
rect 24722 -1511 24822 -1489
rect 24722 -1557 24755 -1511
rect 24789 -1557 24822 -1511
rect 24722 -1583 24822 -1557
rect 24722 -1625 24755 -1583
rect 24789 -1625 24822 -1583
rect 24722 -1655 24822 -1625
rect 24722 -1693 24755 -1655
rect 24789 -1693 24822 -1655
rect 24722 -1727 24822 -1693
rect 24722 -1761 24755 -1727
rect 24789 -1761 24822 -1727
rect 24722 -1795 24822 -1761
rect 24722 -1833 24755 -1795
rect 24789 -1833 24822 -1795
rect 24722 -1863 24822 -1833
rect 24722 -1905 24755 -1863
rect 24789 -1905 24822 -1863
rect 24722 -1931 24822 -1905
rect 24722 -1977 24755 -1931
rect 24789 -1977 24822 -1931
rect 24722 -1999 24822 -1977
rect 24722 -2049 24755 -1999
rect 24789 -2049 24822 -1999
rect 24722 -2067 24822 -2049
rect 24722 -2121 24755 -2067
rect 24789 -2121 24822 -2067
rect 24722 -2135 24822 -2121
rect 24722 -2193 24755 -2135
rect 24789 -2193 24822 -2135
rect 24722 -2203 24822 -2193
rect 24722 -2265 24755 -2203
rect 24789 -2265 24822 -2203
rect 24722 -2271 24822 -2265
rect 24722 -2337 24755 -2271
rect 24789 -2337 24822 -2271
rect 24722 -2339 24822 -2337
rect 24722 -2373 24755 -2339
rect 24789 -2373 24822 -2339
rect 24722 -2375 24822 -2373
rect 24722 -2441 24755 -2375
rect 24789 -2441 24822 -2375
rect 24722 -2447 24822 -2441
rect 24722 -2509 24755 -2447
rect 24789 -2509 24822 -2447
rect 24722 -2519 24822 -2509
rect 24722 -2577 24755 -2519
rect 24789 -2577 24822 -2519
rect 24722 -2591 24822 -2577
rect 24722 -2645 24755 -2591
rect 24789 -2645 24822 -2591
rect 24722 -2663 24822 -2645
rect 24722 -2713 24755 -2663
rect 24789 -2713 24822 -2663
rect 24722 -2735 24822 -2713
rect 24722 -2781 24755 -2735
rect 24789 -2781 24822 -2735
rect 24722 -2807 24822 -2781
rect 24722 -2849 24755 -2807
rect 24789 -2849 24822 -2807
rect 24722 -2879 24822 -2849
rect 24722 -2917 24755 -2879
rect 24789 -2917 24822 -2879
rect 24722 -2951 24822 -2917
rect 24722 -2985 24755 -2951
rect 24789 -2985 24822 -2951
rect 24722 -3019 24822 -2985
rect 24722 -3057 24755 -3019
rect 24789 -3057 24822 -3019
rect 24722 -3087 24822 -3057
rect 24722 -3129 24755 -3087
rect 24789 -3129 24822 -3087
rect 24722 -3155 24822 -3129
rect 24722 -3201 24755 -3155
rect 24789 -3201 24822 -3155
rect 24722 -3223 24822 -3201
rect 24722 -3273 24755 -3223
rect 24789 -3273 24822 -3223
rect 24722 -3291 24822 -3273
rect 24722 -3345 24755 -3291
rect 24789 -3345 24822 -3291
rect 24722 -3359 24822 -3345
rect 24722 -3417 24755 -3359
rect 24789 -3417 24822 -3359
rect 24722 -3427 24822 -3417
rect 24722 -3489 24755 -3427
rect 24789 -3489 24822 -3427
rect 24722 -3495 24822 -3489
rect 24722 -3561 24755 -3495
rect 24789 -3561 24822 -3495
rect 24722 -3563 24822 -3561
rect 24722 -3597 24755 -3563
rect 24789 -3597 24822 -3563
rect 24722 -3599 24822 -3597
rect 24722 -3665 24755 -3599
rect 24789 -3665 24822 -3599
rect 24722 -3671 24822 -3665
rect 24722 -3733 24755 -3671
rect 24789 -3733 24822 -3671
rect 24722 -3743 24822 -3733
rect 24722 -3801 24755 -3743
rect 24789 -3801 24822 -3743
rect 24722 -3815 24822 -3801
rect 24722 -3869 24755 -3815
rect 24789 -3869 24822 -3815
rect 24722 -3887 24822 -3869
rect 24722 -3937 24755 -3887
rect 24789 -3937 24822 -3887
rect 24722 -3959 24822 -3937
rect 24722 -4005 24755 -3959
rect 24789 -4005 24822 -3959
rect 24722 -4031 24822 -4005
rect 24722 -4073 24755 -4031
rect 24789 -4073 24822 -4031
rect 24722 -4103 24822 -4073
rect 24722 -4141 24755 -4103
rect 24789 -4141 24822 -4103
rect 24722 -4175 24822 -4141
rect 24722 -4209 24755 -4175
rect 24789 -4209 24822 -4175
rect 24722 -4243 24822 -4209
rect 24722 -4281 24755 -4243
rect 24789 -4281 24822 -4243
rect 24722 -4311 24822 -4281
rect 24722 -4353 24755 -4311
rect 24789 -4353 24822 -4311
rect 24722 -4379 24822 -4353
rect 24722 -4425 24755 -4379
rect 24789 -4425 24822 -4379
rect 24722 -4447 24822 -4425
rect 24722 -4497 24755 -4447
rect 24789 -4497 24822 -4447
rect 24722 -4515 24822 -4497
rect 24722 -4569 24755 -4515
rect 24789 -4569 24822 -4515
rect 24722 -4583 24822 -4569
rect 378 -4651 478 -4641
rect 3698 -4643 3735 -4609
rect 3769 -4643 3806 -4609
rect 3916 -4643 3953 -4609
rect 3987 -4643 4024 -4609
rect 4134 -4643 4171 -4609
rect 4205 -4643 4242 -4609
rect 4352 -4643 4389 -4609
rect 4423 -4643 4460 -4609
rect 4570 -4643 4607 -4609
rect 4641 -4643 4678 -4609
rect 4788 -4643 4825 -4609
rect 4859 -4643 4896 -4609
rect 5006 -4643 5043 -4609
rect 5077 -4643 5114 -4609
rect 5224 -4643 5261 -4609
rect 5295 -4643 5332 -4609
rect 5442 -4643 5479 -4609
rect 5513 -4643 5550 -4609
rect 5660 -4643 5697 -4609
rect 5731 -4643 5768 -4609
rect 24722 -4641 24755 -4583
rect 24789 -4641 24822 -4583
rect 378 -4713 411 -4651
rect 445 -4713 478 -4651
rect 24722 -4651 24822 -4641
rect 378 -4719 478 -4713
rect 378 -4785 411 -4719
rect 445 -4785 478 -4719
rect 378 -4787 478 -4785
rect 378 -4821 411 -4787
rect 445 -4821 478 -4787
rect 378 -4823 478 -4821
rect 378 -4889 411 -4823
rect 445 -4889 478 -4823
rect 378 -4895 478 -4889
rect 378 -4957 411 -4895
rect 445 -4957 478 -4895
rect 378 -4967 478 -4957
rect 378 -5025 411 -4967
rect 445 -5025 478 -4967
rect 378 -5039 478 -5025
rect 378 -5093 411 -5039
rect 445 -5093 478 -5039
rect 378 -5111 478 -5093
rect 3626 -4703 3660 -4686
rect 3626 -4771 3660 -4763
rect 3626 -4839 3660 -4835
rect 3626 -4945 3660 -4941
rect 3626 -5017 3660 -5009
rect 3626 -5094 3660 -5077
rect 3844 -4703 3878 -4686
rect 3844 -4771 3878 -4763
rect 3844 -4839 3878 -4835
rect 3844 -4945 3878 -4941
rect 3844 -5017 3878 -5009
rect 3844 -5094 3878 -5077
rect 4062 -4703 4096 -4686
rect 4062 -4771 4096 -4763
rect 4062 -4839 4096 -4835
rect 4062 -4945 4096 -4941
rect 4062 -5017 4096 -5009
rect 4062 -5094 4096 -5077
rect 4280 -4703 4314 -4686
rect 4280 -4771 4314 -4763
rect 4280 -4839 4314 -4835
rect 4280 -4945 4314 -4941
rect 4280 -5017 4314 -5009
rect 4280 -5094 4314 -5077
rect 4498 -4703 4532 -4686
rect 4498 -4771 4532 -4763
rect 4498 -4839 4532 -4835
rect 4498 -4945 4532 -4941
rect 4498 -5017 4532 -5009
rect 4498 -5094 4532 -5077
rect 4716 -4703 4750 -4686
rect 4716 -4771 4750 -4763
rect 4716 -4839 4750 -4835
rect 4716 -4945 4750 -4941
rect 4716 -5017 4750 -5009
rect 4716 -5094 4750 -5077
rect 4934 -4703 4968 -4686
rect 4934 -4771 4968 -4763
rect 4934 -4839 4968 -4835
rect 4934 -4945 4968 -4941
rect 4934 -5017 4968 -5009
rect 4934 -5094 4968 -5077
rect 5152 -4703 5186 -4686
rect 5152 -4771 5186 -4763
rect 5152 -4839 5186 -4835
rect 5152 -4945 5186 -4941
rect 5152 -5017 5186 -5009
rect 5152 -5094 5186 -5077
rect 5370 -4703 5404 -4686
rect 5370 -4771 5404 -4763
rect 5370 -4839 5404 -4835
rect 5370 -4945 5404 -4941
rect 5370 -5017 5404 -5009
rect 5370 -5094 5404 -5077
rect 5588 -4703 5622 -4686
rect 5588 -4771 5622 -4763
rect 5588 -4839 5622 -4835
rect 5588 -4945 5622 -4941
rect 5588 -5017 5622 -5009
rect 5588 -5094 5622 -5077
rect 5806 -4703 5840 -4686
rect 5806 -4771 5840 -4763
rect 5806 -4839 5840 -4835
rect 5806 -4945 5840 -4941
rect 5806 -5017 5840 -5009
rect 5806 -5094 5840 -5077
rect 24722 -4713 24755 -4651
rect 24789 -4713 24822 -4651
rect 24722 -4719 24822 -4713
rect 24722 -4785 24755 -4719
rect 24789 -4785 24822 -4719
rect 24722 -4787 24822 -4785
rect 24722 -4821 24755 -4787
rect 24789 -4821 24822 -4787
rect 24722 -4823 24822 -4821
rect 24722 -4889 24755 -4823
rect 24789 -4889 24822 -4823
rect 24722 -4895 24822 -4889
rect 24722 -4957 24755 -4895
rect 24789 -4957 24822 -4895
rect 24722 -4967 24822 -4957
rect 24722 -5025 24755 -4967
rect 24789 -5025 24822 -4967
rect 24722 -5039 24822 -5025
rect 24722 -5093 24755 -5039
rect 24789 -5093 24822 -5039
rect 378 -5161 411 -5111
rect 445 -5161 478 -5111
rect 24722 -5111 24822 -5093
rect 3944 -5137 4004 -5136
rect 378 -5183 478 -5161
rect 3698 -5171 3735 -5137
rect 3769 -5171 3806 -5137
rect 3916 -5171 3953 -5137
rect 3987 -5171 4024 -5137
rect 4134 -5171 4171 -5137
rect 4205 -5171 4242 -5137
rect 4352 -5171 4389 -5137
rect 4423 -5171 4460 -5137
rect 4570 -5171 4607 -5137
rect 4641 -5171 4678 -5137
rect 4788 -5171 4825 -5137
rect 4859 -5171 4896 -5137
rect 5006 -5171 5043 -5137
rect 5077 -5171 5114 -5137
rect 5224 -5171 5261 -5137
rect 5295 -5171 5332 -5137
rect 5442 -5171 5479 -5137
rect 5513 -5171 5550 -5137
rect 5660 -5171 5697 -5137
rect 5731 -5171 5768 -5137
rect 24722 -5161 24755 -5111
rect 24789 -5161 24822 -5111
rect 378 -5229 411 -5183
rect 445 -5229 478 -5183
rect 378 -5255 478 -5229
rect 378 -5297 411 -5255
rect 445 -5297 478 -5255
rect 378 -5327 478 -5297
rect 378 -5365 411 -5327
rect 445 -5365 478 -5327
rect 378 -5399 478 -5365
rect 378 -5433 411 -5399
rect 445 -5433 478 -5399
rect 378 -5467 478 -5433
rect 378 -5505 411 -5467
rect 445 -5505 478 -5467
rect 378 -5535 478 -5505
rect 378 -5577 411 -5535
rect 445 -5577 478 -5535
rect 24722 -5183 24822 -5161
rect 24722 -5229 24755 -5183
rect 24789 -5229 24822 -5183
rect 24722 -5255 24822 -5229
rect 24722 -5297 24755 -5255
rect 24789 -5297 24822 -5255
rect 24722 -5327 24822 -5297
rect 24722 -5365 24755 -5327
rect 24789 -5365 24822 -5327
rect 24722 -5399 24822 -5365
rect 24722 -5433 24755 -5399
rect 24789 -5433 24822 -5399
rect 24722 -5467 24822 -5433
rect 24722 -5505 24755 -5467
rect 24789 -5505 24822 -5467
rect 24722 -5535 24822 -5505
rect 378 -5603 478 -5577
rect 3698 -5581 3735 -5547
rect 3769 -5581 3806 -5547
rect 3916 -5581 3953 -5547
rect 3987 -5581 4024 -5547
rect 4134 -5581 4171 -5547
rect 4205 -5581 4242 -5547
rect 4352 -5581 4389 -5547
rect 4423 -5581 4460 -5547
rect 4570 -5581 4607 -5547
rect 4641 -5581 4678 -5547
rect 4788 -5581 4825 -5547
rect 4859 -5581 4896 -5547
rect 5006 -5581 5043 -5547
rect 5077 -5581 5114 -5547
rect 5224 -5581 5261 -5547
rect 5295 -5581 5332 -5547
rect 5442 -5581 5479 -5547
rect 5513 -5581 5550 -5547
rect 5660 -5581 5697 -5547
rect 5731 -5581 5768 -5547
rect 24722 -5577 24755 -5535
rect 24789 -5577 24822 -5535
rect 378 -5649 411 -5603
rect 445 -5649 478 -5603
rect 24722 -5603 24822 -5577
rect 378 -5671 478 -5649
rect 378 -5721 411 -5671
rect 445 -5721 478 -5671
rect 378 -5739 478 -5721
rect 378 -5793 411 -5739
rect 445 -5793 478 -5739
rect 378 -5807 478 -5793
rect 378 -5865 411 -5807
rect 445 -5865 478 -5807
rect 378 -5875 478 -5865
rect 378 -5937 411 -5875
rect 445 -5937 478 -5875
rect 378 -5943 478 -5937
rect 378 -6009 411 -5943
rect 445 -6009 478 -5943
rect 378 -6011 478 -6009
rect 378 -6045 411 -6011
rect 445 -6045 478 -6011
rect 3626 -5641 3660 -5624
rect 3626 -5709 3660 -5701
rect 3626 -5777 3660 -5773
rect 3626 -5883 3660 -5879
rect 3626 -5955 3660 -5947
rect 3626 -6032 3660 -6015
rect 3844 -5641 3878 -5624
rect 3844 -5709 3878 -5701
rect 3844 -5777 3878 -5773
rect 3844 -5883 3878 -5879
rect 3844 -5955 3878 -5947
rect 3844 -6032 3878 -6015
rect 4062 -5641 4096 -5624
rect 4062 -5709 4096 -5701
rect 4062 -5777 4096 -5773
rect 4062 -5883 4096 -5879
rect 4062 -5955 4096 -5947
rect 4062 -6032 4096 -6015
rect 4280 -5641 4314 -5624
rect 4280 -5709 4314 -5701
rect 4280 -5777 4314 -5773
rect 4280 -5883 4314 -5879
rect 4280 -5955 4314 -5947
rect 4280 -6032 4314 -6015
rect 4498 -5641 4532 -5624
rect 4498 -5709 4532 -5701
rect 4498 -5777 4532 -5773
rect 4498 -5883 4532 -5879
rect 4498 -5955 4532 -5947
rect 4498 -6032 4532 -6015
rect 4716 -5641 4750 -5624
rect 4716 -5709 4750 -5701
rect 4716 -5777 4750 -5773
rect 4716 -5883 4750 -5879
rect 4716 -5955 4750 -5947
rect 4716 -6032 4750 -6015
rect 4934 -5641 4968 -5624
rect 4934 -5709 4968 -5701
rect 4934 -5777 4968 -5773
rect 4934 -5883 4968 -5879
rect 4934 -5955 4968 -5947
rect 4934 -6032 4968 -6015
rect 5152 -5641 5186 -5624
rect 5152 -5709 5186 -5701
rect 5152 -5777 5186 -5773
rect 5152 -5883 5186 -5879
rect 5152 -5955 5186 -5947
rect 5152 -6032 5186 -6015
rect 5370 -5641 5404 -5624
rect 5370 -5709 5404 -5701
rect 5370 -5777 5404 -5773
rect 5370 -5883 5404 -5879
rect 5370 -5955 5404 -5947
rect 5370 -6032 5404 -6015
rect 5588 -5641 5622 -5624
rect 5588 -5709 5622 -5701
rect 5588 -5777 5622 -5773
rect 5588 -5883 5622 -5879
rect 5588 -5955 5622 -5947
rect 5588 -6032 5622 -6015
rect 5806 -5641 5840 -5624
rect 5806 -5709 5840 -5701
rect 5806 -5777 5840 -5773
rect 5806 -5883 5840 -5879
rect 5806 -5955 5840 -5947
rect 5806 -6032 5840 -6015
rect 24722 -5649 24755 -5603
rect 24789 -5649 24822 -5603
rect 24722 -5671 24822 -5649
rect 24722 -5721 24755 -5671
rect 24789 -5721 24822 -5671
rect 24722 -5739 24822 -5721
rect 24722 -5793 24755 -5739
rect 24789 -5793 24822 -5739
rect 24722 -5807 24822 -5793
rect 24722 -5865 24755 -5807
rect 24789 -5865 24822 -5807
rect 24722 -5875 24822 -5865
rect 24722 -5937 24755 -5875
rect 24789 -5937 24822 -5875
rect 24722 -5943 24822 -5937
rect 24722 -6009 24755 -5943
rect 24789 -6009 24822 -5943
rect 24722 -6011 24822 -6009
rect 378 -6047 478 -6045
rect 378 -6113 411 -6047
rect 445 -6113 478 -6047
rect 24722 -6045 24755 -6011
rect 24789 -6045 24822 -6011
rect 24722 -6047 24822 -6045
rect 4376 -6075 4436 -6074
rect 5248 -6075 5308 -6074
rect 3698 -6109 3735 -6075
rect 3769 -6109 3806 -6075
rect 3916 -6109 3953 -6075
rect 3987 -6109 4024 -6075
rect 4134 -6109 4171 -6075
rect 4205 -6109 4242 -6075
rect 4352 -6109 4389 -6075
rect 4423 -6109 4460 -6075
rect 4570 -6109 4607 -6075
rect 4641 -6109 4678 -6075
rect 4788 -6109 4825 -6075
rect 4859 -6109 4896 -6075
rect 5006 -6109 5043 -6075
rect 5077 -6109 5114 -6075
rect 5224 -6109 5261 -6075
rect 5295 -6109 5332 -6075
rect 5442 -6109 5479 -6075
rect 5513 -6109 5550 -6075
rect 5660 -6109 5697 -6075
rect 5731 -6109 5768 -6075
rect 378 -6119 478 -6113
rect 378 -6181 411 -6119
rect 445 -6181 478 -6119
rect 378 -6191 478 -6181
rect 378 -6249 411 -6191
rect 445 -6249 478 -6191
rect 378 -6263 478 -6249
rect 378 -6317 411 -6263
rect 445 -6317 478 -6263
rect 378 -6335 478 -6317
rect 378 -6385 411 -6335
rect 445 -6385 478 -6335
rect 378 -6407 478 -6385
rect 378 -6453 411 -6407
rect 445 -6453 478 -6407
rect 378 -6479 478 -6453
rect 378 -6521 411 -6479
rect 445 -6521 478 -6479
rect 24722 -6113 24755 -6047
rect 24789 -6113 24822 -6047
rect 24722 -6119 24822 -6113
rect 24722 -6181 24755 -6119
rect 24789 -6181 24822 -6119
rect 24722 -6191 24822 -6181
rect 24722 -6249 24755 -6191
rect 24789 -6249 24822 -6191
rect 24722 -6263 24822 -6249
rect 24722 -6317 24755 -6263
rect 24789 -6317 24822 -6263
rect 24722 -6335 24822 -6317
rect 24722 -6385 24755 -6335
rect 24789 -6385 24822 -6335
rect 24722 -6407 24822 -6385
rect 24722 -6453 24755 -6407
rect 24789 -6453 24822 -6407
rect 24722 -6479 24822 -6453
rect 3698 -6519 3735 -6485
rect 3769 -6519 3806 -6485
rect 3916 -6519 3953 -6485
rect 3987 -6519 4024 -6485
rect 4134 -6519 4171 -6485
rect 4205 -6519 4242 -6485
rect 4352 -6519 4389 -6485
rect 4423 -6519 4460 -6485
rect 4570 -6519 4607 -6485
rect 4641 -6519 4678 -6485
rect 4788 -6519 4825 -6485
rect 4859 -6519 4896 -6485
rect 5006 -6519 5043 -6485
rect 5077 -6519 5114 -6485
rect 5224 -6519 5261 -6485
rect 5295 -6519 5332 -6485
rect 5442 -6519 5479 -6485
rect 5513 -6519 5550 -6485
rect 5660 -6519 5697 -6485
rect 5731 -6519 5768 -6485
rect 3938 -6520 3998 -6519
rect 4376 -6520 4436 -6519
rect 378 -6551 478 -6521
rect 378 -6589 411 -6551
rect 445 -6589 478 -6551
rect 24722 -6521 24755 -6479
rect 24789 -6521 24822 -6479
rect 24722 -6551 24822 -6521
rect 378 -6623 478 -6589
rect 378 -6657 411 -6623
rect 445 -6657 478 -6623
rect 378 -6691 478 -6657
rect 378 -6729 411 -6691
rect 445 -6729 478 -6691
rect 378 -6759 478 -6729
rect 378 -6801 411 -6759
rect 445 -6801 478 -6759
rect 378 -6827 478 -6801
rect 378 -6873 411 -6827
rect 445 -6873 478 -6827
rect 378 -6895 478 -6873
rect 378 -6945 411 -6895
rect 445 -6945 478 -6895
rect 378 -6963 478 -6945
rect 378 -7017 411 -6963
rect 445 -7017 478 -6963
rect 3626 -6579 3660 -6562
rect 3626 -6647 3660 -6639
rect 3626 -6715 3660 -6711
rect 3626 -6821 3660 -6817
rect 3626 -6893 3660 -6885
rect 3626 -6970 3660 -6953
rect 3844 -6579 3878 -6562
rect 3844 -6647 3878 -6639
rect 3844 -6715 3878 -6711
rect 3844 -6821 3878 -6817
rect 3844 -6893 3878 -6885
rect 3844 -6970 3878 -6953
rect 4062 -6579 4096 -6562
rect 4062 -6647 4096 -6639
rect 4062 -6715 4096 -6711
rect 4062 -6821 4096 -6817
rect 4062 -6893 4096 -6885
rect 4062 -6970 4096 -6953
rect 4280 -6579 4314 -6562
rect 4280 -6647 4314 -6639
rect 4280 -6715 4314 -6711
rect 4280 -6821 4314 -6817
rect 4280 -6893 4314 -6885
rect 4280 -6970 4314 -6953
rect 4498 -6579 4532 -6562
rect 4498 -6647 4532 -6639
rect 4498 -6715 4532 -6711
rect 4498 -6821 4532 -6817
rect 4498 -6893 4532 -6885
rect 4498 -6970 4532 -6953
rect 4716 -6579 4750 -6562
rect 4716 -6647 4750 -6639
rect 4716 -6715 4750 -6711
rect 4716 -6821 4750 -6817
rect 4716 -6893 4750 -6885
rect 4716 -6970 4750 -6953
rect 4934 -6579 4968 -6562
rect 4934 -6647 4968 -6639
rect 4934 -6715 4968 -6711
rect 4934 -6821 4968 -6817
rect 4934 -6893 4968 -6885
rect 4934 -6970 4968 -6953
rect 5152 -6579 5186 -6562
rect 5152 -6647 5186 -6639
rect 5152 -6715 5186 -6711
rect 5152 -6821 5186 -6817
rect 5152 -6893 5186 -6885
rect 5152 -6970 5186 -6953
rect 5370 -6579 5404 -6562
rect 5370 -6647 5404 -6639
rect 5370 -6715 5404 -6711
rect 5370 -6821 5404 -6817
rect 5370 -6893 5404 -6885
rect 5370 -6970 5404 -6953
rect 5588 -6579 5622 -6562
rect 5588 -6647 5622 -6639
rect 5588 -6715 5622 -6711
rect 5588 -6821 5622 -6817
rect 5588 -6893 5622 -6885
rect 5588 -6970 5622 -6953
rect 5806 -6579 5840 -6562
rect 5806 -6647 5840 -6639
rect 5806 -6715 5840 -6711
rect 5806 -6821 5840 -6817
rect 5806 -6893 5840 -6885
rect 5806 -6970 5840 -6953
rect 24722 -6589 24755 -6551
rect 24789 -6589 24822 -6551
rect 24722 -6623 24822 -6589
rect 24722 -6657 24755 -6623
rect 24789 -6657 24822 -6623
rect 24722 -6691 24822 -6657
rect 24722 -6729 24755 -6691
rect 24789 -6729 24822 -6691
rect 24722 -6759 24822 -6729
rect 24722 -6801 24755 -6759
rect 24789 -6801 24822 -6759
rect 24722 -6827 24822 -6801
rect 24722 -6873 24755 -6827
rect 24789 -6873 24822 -6827
rect 24722 -6895 24822 -6873
rect 24722 -6945 24755 -6895
rect 24789 -6945 24822 -6895
rect 24722 -6963 24822 -6945
rect 378 -7031 478 -7017
rect 378 -7089 411 -7031
rect 445 -7089 478 -7031
rect 3698 -7047 3735 -7013
rect 3769 -7047 3806 -7013
rect 3916 -7047 3953 -7013
rect 3987 -7047 4024 -7013
rect 4134 -7047 4171 -7013
rect 4205 -7047 4242 -7013
rect 4352 -7047 4389 -7013
rect 4423 -7047 4460 -7013
rect 4570 -7047 4607 -7013
rect 4641 -7047 4678 -7013
rect 4788 -7047 4825 -7013
rect 4859 -7047 4896 -7013
rect 5006 -7047 5043 -7013
rect 5077 -7047 5114 -7013
rect 5224 -7047 5261 -7013
rect 5295 -7047 5332 -7013
rect 5442 -7047 5479 -7013
rect 5513 -7047 5550 -7013
rect 5660 -7047 5697 -7013
rect 5731 -7047 5768 -7013
rect 24722 -7017 24755 -6963
rect 24789 -7017 24822 -6963
rect 24722 -7031 24822 -7017
rect 378 -7099 478 -7089
rect 378 -7161 411 -7099
rect 445 -7161 478 -7099
rect 378 -7167 478 -7161
rect 378 -7233 411 -7167
rect 445 -7233 478 -7167
rect 378 -7235 478 -7233
rect 378 -7269 411 -7235
rect 445 -7269 478 -7235
rect 378 -7271 478 -7269
rect 378 -7337 411 -7271
rect 445 -7337 478 -7271
rect 378 -7343 478 -7337
rect 378 -7405 411 -7343
rect 445 -7405 478 -7343
rect 378 -7415 478 -7405
rect 378 -7473 411 -7415
rect 445 -7473 478 -7415
rect 24722 -7089 24755 -7031
rect 24789 -7089 24822 -7031
rect 24722 -7099 24822 -7089
rect 24722 -7161 24755 -7099
rect 24789 -7161 24822 -7099
rect 24722 -7167 24822 -7161
rect 24722 -7233 24755 -7167
rect 24789 -7233 24822 -7167
rect 24722 -7235 24822 -7233
rect 24722 -7269 24755 -7235
rect 24789 -7269 24822 -7235
rect 24722 -7271 24822 -7269
rect 24722 -7337 24755 -7271
rect 24789 -7337 24822 -7271
rect 24722 -7343 24822 -7337
rect 24722 -7405 24755 -7343
rect 24789 -7405 24822 -7343
rect 24722 -7415 24822 -7405
rect 3698 -7457 3735 -7423
rect 3769 -7457 3806 -7423
rect 3916 -7457 3953 -7423
rect 3987 -7457 4024 -7423
rect 4134 -7457 4171 -7423
rect 4205 -7457 4242 -7423
rect 4352 -7457 4389 -7423
rect 4423 -7457 4460 -7423
rect 4570 -7457 4607 -7423
rect 4641 -7457 4678 -7423
rect 4788 -7457 4825 -7423
rect 4859 -7457 4896 -7423
rect 5006 -7457 5043 -7423
rect 5077 -7457 5114 -7423
rect 5224 -7457 5261 -7423
rect 5295 -7457 5332 -7423
rect 5442 -7457 5479 -7423
rect 5513 -7457 5550 -7423
rect 5660 -7457 5697 -7423
rect 5731 -7457 5768 -7423
rect 4380 -7458 4440 -7457
rect 378 -7487 478 -7473
rect 378 -7541 411 -7487
rect 445 -7541 478 -7487
rect 24722 -7473 24755 -7415
rect 24789 -7473 24822 -7415
rect 24722 -7487 24822 -7473
rect 378 -7559 478 -7541
rect 378 -7609 411 -7559
rect 445 -7609 478 -7559
rect 378 -7631 478 -7609
rect 378 -7677 411 -7631
rect 445 -7677 478 -7631
rect 378 -7703 478 -7677
rect 378 -7745 411 -7703
rect 445 -7745 478 -7703
rect 378 -7775 478 -7745
rect 378 -7813 411 -7775
rect 445 -7813 478 -7775
rect 378 -7847 478 -7813
rect 378 -7881 411 -7847
rect 445 -7881 478 -7847
rect 378 -7915 478 -7881
rect 3626 -7517 3660 -7500
rect 3626 -7585 3660 -7577
rect 3626 -7653 3660 -7649
rect 3626 -7759 3660 -7755
rect 3626 -7831 3660 -7823
rect 3626 -7908 3660 -7891
rect 3844 -7517 3878 -7500
rect 3844 -7585 3878 -7577
rect 3844 -7653 3878 -7649
rect 3844 -7759 3878 -7755
rect 3844 -7831 3878 -7823
rect 3844 -7908 3878 -7891
rect 4062 -7517 4096 -7500
rect 4062 -7585 4096 -7577
rect 4062 -7653 4096 -7649
rect 4062 -7759 4096 -7755
rect 4062 -7831 4096 -7823
rect 4062 -7908 4096 -7891
rect 4280 -7517 4314 -7500
rect 4280 -7585 4314 -7577
rect 4280 -7653 4314 -7649
rect 4280 -7759 4314 -7755
rect 4280 -7831 4314 -7823
rect 4280 -7908 4314 -7891
rect 4498 -7517 4532 -7500
rect 4498 -7585 4532 -7577
rect 4498 -7653 4532 -7649
rect 4498 -7759 4532 -7755
rect 4498 -7831 4532 -7823
rect 4498 -7908 4532 -7891
rect 4716 -7517 4750 -7500
rect 4716 -7585 4750 -7577
rect 4716 -7653 4750 -7649
rect 4716 -7759 4750 -7755
rect 4716 -7831 4750 -7823
rect 4716 -7908 4750 -7891
rect 4934 -7517 4968 -7500
rect 4934 -7585 4968 -7577
rect 4934 -7653 4968 -7649
rect 4934 -7759 4968 -7755
rect 4934 -7831 4968 -7823
rect 4934 -7908 4968 -7891
rect 5152 -7517 5186 -7500
rect 5152 -7585 5186 -7577
rect 5152 -7653 5186 -7649
rect 5152 -7759 5186 -7755
rect 5152 -7831 5186 -7823
rect 5152 -7908 5186 -7891
rect 5370 -7517 5404 -7500
rect 5370 -7585 5404 -7577
rect 5370 -7653 5404 -7649
rect 5370 -7759 5404 -7755
rect 5370 -7831 5404 -7823
rect 5370 -7908 5404 -7891
rect 5588 -7517 5622 -7500
rect 5588 -7585 5622 -7577
rect 5588 -7653 5622 -7649
rect 5588 -7759 5622 -7755
rect 5588 -7831 5622 -7823
rect 5588 -7908 5622 -7891
rect 5806 -7517 5840 -7500
rect 5806 -7585 5840 -7577
rect 5806 -7653 5840 -7649
rect 5806 -7759 5840 -7755
rect 5806 -7831 5840 -7823
rect 5806 -7908 5840 -7891
rect 24722 -7541 24755 -7487
rect 24789 -7541 24822 -7487
rect 24722 -7559 24822 -7541
rect 24722 -7609 24755 -7559
rect 24789 -7609 24822 -7559
rect 24722 -7631 24822 -7609
rect 24722 -7677 24755 -7631
rect 24789 -7677 24822 -7631
rect 24722 -7703 24822 -7677
rect 24722 -7745 24755 -7703
rect 24789 -7745 24822 -7703
rect 24722 -7775 24822 -7745
rect 24722 -7813 24755 -7775
rect 24789 -7813 24822 -7775
rect 24722 -7847 24822 -7813
rect 24722 -7881 24755 -7847
rect 24789 -7881 24822 -7847
rect 378 -7953 411 -7915
rect 445 -7953 478 -7915
rect 24722 -7915 24822 -7881
rect 378 -7983 478 -7953
rect 378 -8025 411 -7983
rect 445 -8025 478 -7983
rect 3698 -7985 3735 -7951
rect 3769 -7985 3806 -7951
rect 3916 -7985 3953 -7951
rect 3987 -7985 4024 -7951
rect 4134 -7985 4171 -7951
rect 4205 -7985 4242 -7951
rect 4352 -7985 4389 -7951
rect 4423 -7985 4460 -7951
rect 4570 -7985 4607 -7951
rect 4641 -7985 4678 -7951
rect 4788 -7985 4825 -7951
rect 4859 -7985 4896 -7951
rect 5006 -7985 5043 -7951
rect 5077 -7985 5114 -7951
rect 5224 -7985 5261 -7951
rect 5295 -7985 5332 -7951
rect 5442 -7985 5479 -7951
rect 5513 -7985 5550 -7951
rect 5660 -7985 5697 -7951
rect 5731 -7985 5768 -7951
rect 24722 -7953 24755 -7915
rect 24789 -7953 24822 -7915
rect 24722 -7983 24822 -7953
rect 378 -8051 478 -8025
rect 378 -8097 411 -8051
rect 445 -8097 478 -8051
rect 378 -8119 478 -8097
rect 378 -8169 411 -8119
rect 445 -8169 478 -8119
rect 378 -8187 478 -8169
rect 378 -8241 411 -8187
rect 445 -8241 478 -8187
rect 378 -8255 478 -8241
rect 378 -8289 411 -8255
rect 445 -8289 478 -8255
rect 378 -8323 478 -8289
rect 378 -8357 411 -8323
rect 445 -8357 478 -8323
rect 378 -8391 478 -8357
rect 378 -8425 411 -8391
rect 445 -8425 478 -8391
rect 378 -8459 478 -8425
rect 378 -8493 411 -8459
rect 445 -8493 478 -8459
rect 378 -8527 478 -8493
rect 378 -8561 411 -8527
rect 445 -8561 478 -8527
rect 378 -8595 478 -8561
rect 378 -8629 411 -8595
rect 445 -8629 478 -8595
rect 378 -8663 478 -8629
rect 378 -8697 411 -8663
rect 445 -8697 478 -8663
rect 378 -8782 478 -8697
rect 24722 -8025 24755 -7983
rect 24789 -8025 24822 -7983
rect 24722 -8051 24822 -8025
rect 24722 -8097 24755 -8051
rect 24789 -8097 24822 -8051
rect 24722 -8119 24822 -8097
rect 24722 -8169 24755 -8119
rect 24789 -8169 24822 -8119
rect 24722 -8187 24822 -8169
rect 24722 -8241 24755 -8187
rect 24789 -8241 24822 -8187
rect 24722 -8255 24822 -8241
rect 24722 -8289 24755 -8255
rect 24789 -8289 24822 -8255
rect 24722 -8323 24822 -8289
rect 24722 -8357 24755 -8323
rect 24789 -8357 24822 -8323
rect 24722 -8391 24822 -8357
rect 24722 -8425 24755 -8391
rect 24789 -8425 24822 -8391
rect 24722 -8459 24822 -8425
rect 24722 -8493 24755 -8459
rect 24789 -8493 24822 -8459
rect 24722 -8527 24822 -8493
rect 24722 -8561 24755 -8527
rect 24789 -8561 24822 -8527
rect 24722 -8595 24822 -8561
rect 24722 -8629 24755 -8595
rect 24789 -8629 24822 -8595
rect 24722 -8663 24822 -8629
rect 24722 -8697 24755 -8663
rect 24789 -8697 24822 -8663
rect 24722 -8782 24822 -8697
rect 378 -8815 24822 -8782
rect 378 -8849 487 -8815
rect 521 -8849 547 -8815
rect 593 -8849 615 -8815
rect 665 -8849 683 -8815
rect 737 -8849 751 -8815
rect 809 -8849 819 -8815
rect 881 -8849 887 -8815
rect 953 -8849 955 -8815
rect 989 -8849 991 -8815
rect 1057 -8849 1063 -8815
rect 1125 -8849 1135 -8815
rect 1193 -8849 1207 -8815
rect 1261 -8849 1279 -8815
rect 1329 -8849 1351 -8815
rect 1397 -8849 1423 -8815
rect 1465 -8849 1495 -8815
rect 1533 -8849 1567 -8815
rect 1601 -8849 1635 -8815
rect 1673 -8849 1703 -8815
rect 1745 -8849 1771 -8815
rect 1817 -8849 1839 -8815
rect 1889 -8849 1907 -8815
rect 1961 -8849 1975 -8815
rect 2033 -8849 2043 -8815
rect 2105 -8849 2111 -8815
rect 2177 -8849 2179 -8815
rect 2213 -8849 2215 -8815
rect 2281 -8849 2287 -8815
rect 2349 -8849 2359 -8815
rect 2417 -8849 2431 -8815
rect 2485 -8849 2503 -8815
rect 2553 -8849 2575 -8815
rect 2621 -8849 2647 -8815
rect 2689 -8849 2719 -8815
rect 2757 -8849 2791 -8815
rect 2825 -8849 2859 -8815
rect 2897 -8849 2927 -8815
rect 2969 -8849 2995 -8815
rect 3041 -8849 3063 -8815
rect 3113 -8849 3131 -8815
rect 3185 -8849 3199 -8815
rect 3257 -8849 3267 -8815
rect 3329 -8849 3335 -8815
rect 3401 -8849 3403 -8815
rect 3437 -8849 3439 -8815
rect 3505 -8849 3511 -8815
rect 3573 -8849 3583 -8815
rect 3641 -8849 3655 -8815
rect 3709 -8849 3727 -8815
rect 3777 -8849 3799 -8815
rect 3845 -8849 3871 -8815
rect 3913 -8849 3943 -8815
rect 3981 -8849 4015 -8815
rect 4049 -8849 4083 -8815
rect 4121 -8849 4151 -8815
rect 4193 -8849 4219 -8815
rect 4265 -8849 4287 -8815
rect 4337 -8849 4355 -8815
rect 4409 -8849 4423 -8815
rect 4481 -8849 4491 -8815
rect 4553 -8849 4559 -8815
rect 4625 -8849 4627 -8815
rect 4661 -8849 4663 -8815
rect 4729 -8849 4735 -8815
rect 4797 -8849 4807 -8815
rect 4865 -8849 4879 -8815
rect 4933 -8849 4951 -8815
rect 5001 -8849 5023 -8815
rect 5069 -8849 5095 -8815
rect 5137 -8849 5167 -8815
rect 5205 -8849 5239 -8815
rect 5273 -8849 5307 -8815
rect 5345 -8849 5375 -8815
rect 5417 -8849 5443 -8815
rect 5489 -8849 5511 -8815
rect 5561 -8849 5579 -8815
rect 5633 -8849 5647 -8815
rect 5705 -8849 5715 -8815
rect 5777 -8849 5783 -8815
rect 5849 -8849 5851 -8815
rect 5885 -8849 5887 -8815
rect 5953 -8849 5959 -8815
rect 6021 -8849 6031 -8815
rect 6089 -8849 6103 -8815
rect 6157 -8849 6175 -8815
rect 6225 -8849 6247 -8815
rect 6293 -8849 6319 -8815
rect 6361 -8849 6391 -8815
rect 6429 -8849 6463 -8815
rect 6497 -8849 6531 -8815
rect 6569 -8849 6599 -8815
rect 6641 -8849 6667 -8815
rect 6713 -8849 6735 -8815
rect 6785 -8849 6803 -8815
rect 6857 -8849 6871 -8815
rect 6929 -8849 6939 -8815
rect 7001 -8849 7007 -8815
rect 7073 -8849 7075 -8815
rect 7109 -8849 7111 -8815
rect 7177 -8849 7183 -8815
rect 7245 -8849 7255 -8815
rect 7313 -8849 7327 -8815
rect 7381 -8849 7399 -8815
rect 7449 -8849 7471 -8815
rect 7517 -8849 7543 -8815
rect 7585 -8849 7615 -8815
rect 7653 -8849 7687 -8815
rect 7721 -8849 7755 -8815
rect 7793 -8849 7823 -8815
rect 7865 -8849 7891 -8815
rect 7937 -8849 7959 -8815
rect 8009 -8849 8027 -8815
rect 8081 -8849 8095 -8815
rect 8153 -8849 8163 -8815
rect 8225 -8849 8231 -8815
rect 8297 -8849 8299 -8815
rect 8333 -8849 8335 -8815
rect 8401 -8849 8407 -8815
rect 8469 -8849 8479 -8815
rect 8537 -8849 8551 -8815
rect 8605 -8849 8623 -8815
rect 8673 -8849 8695 -8815
rect 8741 -8849 8767 -8815
rect 8809 -8849 8839 -8815
rect 8877 -8849 8911 -8815
rect 8945 -8849 8979 -8815
rect 9017 -8849 9047 -8815
rect 9089 -8849 9115 -8815
rect 9161 -8849 9183 -8815
rect 9233 -8849 9251 -8815
rect 9305 -8849 9319 -8815
rect 9377 -8849 9387 -8815
rect 9449 -8849 9455 -8815
rect 9521 -8849 9523 -8815
rect 9557 -8849 9559 -8815
rect 9625 -8849 9631 -8815
rect 9693 -8849 9703 -8815
rect 9761 -8849 9775 -8815
rect 9829 -8849 9847 -8815
rect 9897 -8849 9919 -8815
rect 9965 -8849 9991 -8815
rect 10033 -8849 10063 -8815
rect 10101 -8849 10135 -8815
rect 10169 -8849 10203 -8815
rect 10241 -8849 10271 -8815
rect 10313 -8849 10339 -8815
rect 10385 -8849 10407 -8815
rect 10457 -8849 10475 -8815
rect 10529 -8849 10543 -8815
rect 10601 -8849 10611 -8815
rect 10673 -8849 10679 -8815
rect 10745 -8849 10747 -8815
rect 10781 -8849 10783 -8815
rect 10849 -8849 10855 -8815
rect 10917 -8849 10927 -8815
rect 10985 -8849 10999 -8815
rect 11053 -8849 11071 -8815
rect 11121 -8849 11143 -8815
rect 11189 -8849 11215 -8815
rect 11257 -8849 11287 -8815
rect 11325 -8849 11359 -8815
rect 11393 -8849 11427 -8815
rect 11465 -8849 11495 -8815
rect 11537 -8849 11563 -8815
rect 11609 -8849 11631 -8815
rect 11681 -8849 11699 -8815
rect 11753 -8849 11767 -8815
rect 11825 -8849 11835 -8815
rect 11897 -8849 11903 -8815
rect 11969 -8849 11971 -8815
rect 12005 -8849 12007 -8815
rect 12073 -8849 12079 -8815
rect 12141 -8849 12151 -8815
rect 12209 -8849 12223 -8815
rect 12277 -8849 12295 -8815
rect 12345 -8849 12367 -8815
rect 12413 -8849 12439 -8815
rect 12481 -8849 12511 -8815
rect 12549 -8849 12583 -8815
rect 12617 -8849 12651 -8815
rect 12689 -8849 12719 -8815
rect 12761 -8849 12787 -8815
rect 12833 -8849 12855 -8815
rect 12905 -8849 12923 -8815
rect 12977 -8849 12991 -8815
rect 13049 -8849 13059 -8815
rect 13121 -8849 13127 -8815
rect 13193 -8849 13195 -8815
rect 13229 -8849 13231 -8815
rect 13297 -8849 13303 -8815
rect 13365 -8849 13375 -8815
rect 13433 -8849 13447 -8815
rect 13501 -8849 13519 -8815
rect 13569 -8849 13591 -8815
rect 13637 -8849 13663 -8815
rect 13705 -8849 13735 -8815
rect 13773 -8849 13807 -8815
rect 13841 -8849 13875 -8815
rect 13913 -8849 13943 -8815
rect 13985 -8849 14011 -8815
rect 14057 -8849 14079 -8815
rect 14129 -8849 14147 -8815
rect 14201 -8849 14215 -8815
rect 14273 -8849 14283 -8815
rect 14345 -8849 14351 -8815
rect 14417 -8849 14419 -8815
rect 14453 -8849 14455 -8815
rect 14521 -8849 14527 -8815
rect 14589 -8849 14599 -8815
rect 14657 -8849 14671 -8815
rect 14725 -8849 14743 -8815
rect 14793 -8849 14815 -8815
rect 14861 -8849 14887 -8815
rect 14929 -8849 14959 -8815
rect 14997 -8849 15031 -8815
rect 15065 -8849 15099 -8815
rect 15137 -8849 15167 -8815
rect 15209 -8849 15235 -8815
rect 15281 -8849 15303 -8815
rect 15353 -8849 15371 -8815
rect 15425 -8849 15439 -8815
rect 15497 -8849 15507 -8815
rect 15569 -8849 15575 -8815
rect 15641 -8849 15643 -8815
rect 15677 -8849 15679 -8815
rect 15745 -8849 15751 -8815
rect 15813 -8849 15823 -8815
rect 15881 -8849 15895 -8815
rect 15949 -8849 15967 -8815
rect 16017 -8849 16039 -8815
rect 16085 -8849 16111 -8815
rect 16153 -8849 16183 -8815
rect 16221 -8849 16255 -8815
rect 16289 -8849 16323 -8815
rect 16361 -8849 16391 -8815
rect 16433 -8849 16459 -8815
rect 16505 -8849 16527 -8815
rect 16577 -8849 16595 -8815
rect 16649 -8849 16663 -8815
rect 16721 -8849 16731 -8815
rect 16793 -8849 16799 -8815
rect 16865 -8849 16867 -8815
rect 16901 -8849 16903 -8815
rect 16969 -8849 16975 -8815
rect 17037 -8849 17047 -8815
rect 17105 -8849 17119 -8815
rect 17173 -8849 17191 -8815
rect 17241 -8849 17263 -8815
rect 17309 -8849 17335 -8815
rect 17377 -8849 17407 -8815
rect 17445 -8849 17479 -8815
rect 17513 -8849 17547 -8815
rect 17585 -8849 17615 -8815
rect 17657 -8849 17683 -8815
rect 17729 -8849 17751 -8815
rect 17801 -8849 17819 -8815
rect 17873 -8849 17887 -8815
rect 17945 -8849 17955 -8815
rect 18017 -8849 18023 -8815
rect 18089 -8849 18091 -8815
rect 18125 -8849 18127 -8815
rect 18193 -8849 18199 -8815
rect 18261 -8849 18271 -8815
rect 18329 -8849 18343 -8815
rect 18397 -8849 18415 -8815
rect 18465 -8849 18487 -8815
rect 18533 -8849 18559 -8815
rect 18601 -8849 18631 -8815
rect 18669 -8849 18703 -8815
rect 18737 -8849 18771 -8815
rect 18809 -8849 18839 -8815
rect 18881 -8849 18907 -8815
rect 18953 -8849 18975 -8815
rect 19025 -8849 19043 -8815
rect 19097 -8849 19111 -8815
rect 19169 -8849 19179 -8815
rect 19241 -8849 19247 -8815
rect 19313 -8849 19315 -8815
rect 19349 -8849 19351 -8815
rect 19417 -8849 19423 -8815
rect 19485 -8849 19495 -8815
rect 19553 -8849 19567 -8815
rect 19621 -8849 19639 -8815
rect 19689 -8849 19711 -8815
rect 19757 -8849 19783 -8815
rect 19825 -8849 19855 -8815
rect 19893 -8849 19927 -8815
rect 19961 -8849 19995 -8815
rect 20033 -8849 20063 -8815
rect 20105 -8849 20131 -8815
rect 20177 -8849 20199 -8815
rect 20249 -8849 20267 -8815
rect 20321 -8849 20335 -8815
rect 20393 -8849 20403 -8815
rect 20465 -8849 20471 -8815
rect 20537 -8849 20539 -8815
rect 20573 -8849 20575 -8815
rect 20641 -8849 20647 -8815
rect 20709 -8849 20719 -8815
rect 20777 -8849 20791 -8815
rect 20845 -8849 20863 -8815
rect 20913 -8849 20935 -8815
rect 20981 -8849 21007 -8815
rect 21049 -8849 21079 -8815
rect 21117 -8849 21151 -8815
rect 21185 -8849 21219 -8815
rect 21257 -8849 21287 -8815
rect 21329 -8849 21355 -8815
rect 21401 -8849 21423 -8815
rect 21473 -8849 21491 -8815
rect 21545 -8849 21559 -8815
rect 21617 -8849 21627 -8815
rect 21689 -8849 21695 -8815
rect 21761 -8849 21763 -8815
rect 21797 -8849 21799 -8815
rect 21865 -8849 21871 -8815
rect 21933 -8849 21943 -8815
rect 22001 -8849 22015 -8815
rect 22069 -8849 22087 -8815
rect 22137 -8849 22159 -8815
rect 22205 -8849 22231 -8815
rect 22273 -8849 22303 -8815
rect 22341 -8849 22375 -8815
rect 22409 -8849 22443 -8815
rect 22481 -8849 22511 -8815
rect 22553 -8849 22579 -8815
rect 22625 -8849 22647 -8815
rect 22697 -8849 22715 -8815
rect 22769 -8849 22783 -8815
rect 22841 -8849 22851 -8815
rect 22913 -8849 22919 -8815
rect 22985 -8849 22987 -8815
rect 23021 -8849 23023 -8815
rect 23089 -8849 23095 -8815
rect 23157 -8849 23167 -8815
rect 23225 -8849 23239 -8815
rect 23293 -8849 23311 -8815
rect 23361 -8849 23383 -8815
rect 23429 -8849 23455 -8815
rect 23497 -8849 23527 -8815
rect 23565 -8849 23599 -8815
rect 23633 -8849 23667 -8815
rect 23705 -8849 23735 -8815
rect 23777 -8849 23803 -8815
rect 23849 -8849 23871 -8815
rect 23921 -8849 23939 -8815
rect 23993 -8849 24007 -8815
rect 24065 -8849 24075 -8815
rect 24137 -8849 24143 -8815
rect 24209 -8849 24211 -8815
rect 24245 -8849 24247 -8815
rect 24313 -8849 24319 -8815
rect 24381 -8849 24391 -8815
rect 24449 -8849 24463 -8815
rect 24517 -8849 24535 -8815
rect 24585 -8849 24607 -8815
rect 24653 -8849 24679 -8815
rect 24713 -8849 24822 -8815
rect 378 -8882 24822 -8849
rect -12322 -11211 24922 -11178
rect -12322 -11245 -12221 -11211
rect -12187 -11245 -12149 -11211
rect -12111 -11245 -12077 -11211
rect -12043 -11245 -12009 -11211
rect -11971 -11245 -11941 -11211
rect -11899 -11245 -11873 -11211
rect -11827 -11245 -11805 -11211
rect -11755 -11245 -11737 -11211
rect -11683 -11245 -11669 -11211
rect -11611 -11245 -11601 -11211
rect -11539 -11245 -11533 -11211
rect -11467 -11245 -11465 -11211
rect -11431 -11245 -11429 -11211
rect -11363 -11245 -11357 -11211
rect -11295 -11245 -11285 -11211
rect -11227 -11245 -11213 -11211
rect -11159 -11245 -11141 -11211
rect -11091 -11245 -11069 -11211
rect -11023 -11245 -10997 -11211
rect -10955 -11245 -10925 -11211
rect -10887 -11245 -10853 -11211
rect -10819 -11245 -10785 -11211
rect -10747 -11245 -10717 -11211
rect -10675 -11245 -10649 -11211
rect -10603 -11245 -10581 -11211
rect -10531 -11245 -10513 -11211
rect -10459 -11245 -10445 -11211
rect -10387 -11245 -10377 -11211
rect -10315 -11245 -10309 -11211
rect -10243 -11245 -10241 -11211
rect -10207 -11245 -10205 -11211
rect -10139 -11245 -10133 -11211
rect -10071 -11245 -10061 -11211
rect -10003 -11245 -9989 -11211
rect -9935 -11245 -9917 -11211
rect -9867 -11245 -9845 -11211
rect -9799 -11245 -9773 -11211
rect -9731 -11245 -9701 -11211
rect -9663 -11245 -9629 -11211
rect -9595 -11245 -9561 -11211
rect -9523 -11245 -9493 -11211
rect -9451 -11245 -9425 -11211
rect -9379 -11245 -9357 -11211
rect -9307 -11245 -9289 -11211
rect -9235 -11245 -9221 -11211
rect -9163 -11245 -9153 -11211
rect -9091 -11245 -9085 -11211
rect -9019 -11245 -9017 -11211
rect -8983 -11245 -8981 -11211
rect -8915 -11245 -8909 -11211
rect -8847 -11245 -8837 -11211
rect -8779 -11245 -8765 -11211
rect -8711 -11245 -8693 -11211
rect -8643 -11245 -8621 -11211
rect -8575 -11245 -8549 -11211
rect -8507 -11245 -8477 -11211
rect -8439 -11245 -8405 -11211
rect -8371 -11245 -8337 -11211
rect -8299 -11245 -8269 -11211
rect -8227 -11245 -8201 -11211
rect -8155 -11245 -8133 -11211
rect -8083 -11245 -8065 -11211
rect -8011 -11245 -7997 -11211
rect -7939 -11245 -7929 -11211
rect -7867 -11245 -7861 -11211
rect -7795 -11245 -7793 -11211
rect -7759 -11245 -7757 -11211
rect -7691 -11245 -7685 -11211
rect -7623 -11245 -7613 -11211
rect -7555 -11245 -7541 -11211
rect -7487 -11245 -7469 -11211
rect -7419 -11245 -7397 -11211
rect -7351 -11245 -7325 -11211
rect -7283 -11245 -7253 -11211
rect -7215 -11245 -7181 -11211
rect -7147 -11245 -7113 -11211
rect -7075 -11245 -7045 -11211
rect -7003 -11245 -6977 -11211
rect -6931 -11245 -6909 -11211
rect -6859 -11245 -6841 -11211
rect -6787 -11245 -6773 -11211
rect -6715 -11245 -6705 -11211
rect -6643 -11245 -6637 -11211
rect -6571 -11245 -6569 -11211
rect -6535 -11245 -6533 -11211
rect -6467 -11245 -6461 -11211
rect -6399 -11245 -6389 -11211
rect -6331 -11245 -6317 -11211
rect -6263 -11245 -6245 -11211
rect -6195 -11245 -6173 -11211
rect -6127 -11245 -6101 -11211
rect -6059 -11245 -6029 -11211
rect -5991 -11245 -5957 -11211
rect -5923 -11245 -5889 -11211
rect -5851 -11245 -5821 -11211
rect -5779 -11245 -5753 -11211
rect -5707 -11245 -5685 -11211
rect -5635 -11245 -5617 -11211
rect -5563 -11245 -5549 -11211
rect -5491 -11245 -5481 -11211
rect -5419 -11245 -5413 -11211
rect -5347 -11245 -5345 -11211
rect -5311 -11245 -5309 -11211
rect -5243 -11245 -5237 -11211
rect -5175 -11245 -5165 -11211
rect -5107 -11245 -5093 -11211
rect -5039 -11245 -5021 -11211
rect -4971 -11245 -4949 -11211
rect -4903 -11245 -4877 -11211
rect -4835 -11245 -4805 -11211
rect -4767 -11245 -4733 -11211
rect -4699 -11245 -4665 -11211
rect -4627 -11245 -4597 -11211
rect -4555 -11245 -4529 -11211
rect -4483 -11245 -4461 -11211
rect -4411 -11245 -4393 -11211
rect -4339 -11245 -4325 -11211
rect -4267 -11245 -4257 -11211
rect -4195 -11245 -4189 -11211
rect -4123 -11245 -4121 -11211
rect -4087 -11245 -4085 -11211
rect -4019 -11245 -4013 -11211
rect -3951 -11245 -3941 -11211
rect -3883 -11245 -3869 -11211
rect -3815 -11245 -3797 -11211
rect -3747 -11245 -3725 -11211
rect -3679 -11245 -3653 -11211
rect -3611 -11245 -3581 -11211
rect -3543 -11245 -3509 -11211
rect -3475 -11245 -3441 -11211
rect -3403 -11245 -3373 -11211
rect -3331 -11245 -3305 -11211
rect -3259 -11245 -3237 -11211
rect -3187 -11245 -3169 -11211
rect -3115 -11245 -3101 -11211
rect -3043 -11245 -3033 -11211
rect -2971 -11245 -2965 -11211
rect -2899 -11245 -2897 -11211
rect -2863 -11245 -2861 -11211
rect -2795 -11245 -2789 -11211
rect -2727 -11245 -2717 -11211
rect -2659 -11245 -2645 -11211
rect -2591 -11245 -2573 -11211
rect -2523 -11245 -2501 -11211
rect -2455 -11245 -2429 -11211
rect -2387 -11245 -2357 -11211
rect -2319 -11245 -2285 -11211
rect -2251 -11245 -2217 -11211
rect -2179 -11245 -2149 -11211
rect -2107 -11245 -2081 -11211
rect -2035 -11245 -2013 -11211
rect -1963 -11245 -1945 -11211
rect -1891 -11245 -1877 -11211
rect -1819 -11245 -1809 -11211
rect -1747 -11245 -1741 -11211
rect -1675 -11245 -1673 -11211
rect -1639 -11245 -1637 -11211
rect -1571 -11245 -1565 -11211
rect -1503 -11245 -1493 -11211
rect -1435 -11245 -1421 -11211
rect -1367 -11245 -1349 -11211
rect -1299 -11245 -1277 -11211
rect -1231 -11245 -1205 -11211
rect -1163 -11245 -1133 -11211
rect -1095 -11245 -1061 -11211
rect -1027 -11245 -993 -11211
rect -955 -11245 -925 -11211
rect -883 -11245 -857 -11211
rect -811 -11245 -789 -11211
rect -739 -11245 -721 -11211
rect -667 -11245 -653 -11211
rect -595 -11245 -585 -11211
rect -523 -11245 -517 -11211
rect -451 -11245 -449 -11211
rect -415 -11245 -413 -11211
rect -347 -11245 -341 -11211
rect -279 -11245 -269 -11211
rect -211 -11245 -197 -11211
rect -143 -11245 -125 -11211
rect -75 -11245 -53 -11211
rect -7 -11245 19 -11211
rect 61 -11245 91 -11211
rect 129 -11245 163 -11211
rect 197 -11245 231 -11211
rect 269 -11245 299 -11211
rect 341 -11245 367 -11211
rect 413 -11245 435 -11211
rect 485 -11245 503 -11211
rect 557 -11245 571 -11211
rect 629 -11245 639 -11211
rect 701 -11245 707 -11211
rect 773 -11245 775 -11211
rect 809 -11245 811 -11211
rect 877 -11245 883 -11211
rect 945 -11245 955 -11211
rect 1013 -11245 1027 -11211
rect 1081 -11245 1099 -11211
rect 1149 -11245 1171 -11211
rect 1217 -11245 1243 -11211
rect 1285 -11245 1315 -11211
rect 1353 -11245 1387 -11211
rect 1421 -11245 1455 -11211
rect 1493 -11245 1523 -11211
rect 1565 -11245 1591 -11211
rect 1637 -11245 1659 -11211
rect 1709 -11245 1727 -11211
rect 1781 -11245 1795 -11211
rect 1853 -11245 1863 -11211
rect 1925 -11245 1931 -11211
rect 1997 -11245 1999 -11211
rect 2033 -11245 2035 -11211
rect 2101 -11245 2107 -11211
rect 2169 -11245 2179 -11211
rect 2237 -11245 2251 -11211
rect 2305 -11245 2323 -11211
rect 2373 -11245 2395 -11211
rect 2441 -11245 2467 -11211
rect 2509 -11245 2539 -11211
rect 2577 -11245 2611 -11211
rect 2645 -11245 2679 -11211
rect 2717 -11245 2747 -11211
rect 2789 -11245 2815 -11211
rect 2861 -11245 2883 -11211
rect 2933 -11245 2951 -11211
rect 3005 -11245 3019 -11211
rect 3077 -11245 3087 -11211
rect 3149 -11245 3155 -11211
rect 3221 -11245 3223 -11211
rect 3257 -11245 3259 -11211
rect 3325 -11245 3331 -11211
rect 3393 -11245 3403 -11211
rect 3461 -11245 3475 -11211
rect 3529 -11245 3547 -11211
rect 3597 -11245 3619 -11211
rect 3665 -11245 3691 -11211
rect 3733 -11245 3763 -11211
rect 3801 -11245 3835 -11211
rect 3869 -11245 3903 -11211
rect 3941 -11245 3971 -11211
rect 4013 -11245 4039 -11211
rect 4085 -11245 4107 -11211
rect 4157 -11245 4175 -11211
rect 4229 -11245 4243 -11211
rect 4301 -11245 4311 -11211
rect 4373 -11245 4379 -11211
rect 4445 -11245 4447 -11211
rect 4481 -11245 4483 -11211
rect 4549 -11245 4555 -11211
rect 4617 -11245 4627 -11211
rect 4685 -11245 4699 -11211
rect 4753 -11245 4771 -11211
rect 4821 -11245 4843 -11211
rect 4889 -11245 4915 -11211
rect 4957 -11245 4987 -11211
rect 5025 -11245 5059 -11211
rect 5093 -11245 5127 -11211
rect 5165 -11245 5195 -11211
rect 5237 -11245 5263 -11211
rect 5309 -11245 5331 -11211
rect 5381 -11245 5399 -11211
rect 5453 -11245 5467 -11211
rect 5525 -11245 5535 -11211
rect 5597 -11245 5603 -11211
rect 5669 -11245 5671 -11211
rect 5705 -11245 5707 -11211
rect 5773 -11245 5779 -11211
rect 5841 -11245 5851 -11211
rect 5909 -11245 5923 -11211
rect 5977 -11245 5995 -11211
rect 6045 -11245 6067 -11211
rect 6113 -11245 6139 -11211
rect 6181 -11245 6211 -11211
rect 6249 -11245 6283 -11211
rect 6317 -11245 6351 -11211
rect 6389 -11245 6419 -11211
rect 6461 -11245 6487 -11211
rect 6533 -11245 6555 -11211
rect 6605 -11245 6623 -11211
rect 6677 -11245 6691 -11211
rect 6749 -11245 6759 -11211
rect 6821 -11245 6827 -11211
rect 6893 -11245 6895 -11211
rect 6929 -11245 6931 -11211
rect 6997 -11245 7003 -11211
rect 7065 -11245 7075 -11211
rect 7133 -11245 7147 -11211
rect 7201 -11245 7219 -11211
rect 7269 -11245 7291 -11211
rect 7337 -11245 7363 -11211
rect 7405 -11245 7435 -11211
rect 7473 -11245 7507 -11211
rect 7541 -11245 7575 -11211
rect 7613 -11245 7643 -11211
rect 7685 -11245 7711 -11211
rect 7757 -11245 7779 -11211
rect 7829 -11245 7847 -11211
rect 7901 -11245 7915 -11211
rect 7973 -11245 7983 -11211
rect 8045 -11245 8051 -11211
rect 8117 -11245 8119 -11211
rect 8153 -11245 8155 -11211
rect 8221 -11245 8227 -11211
rect 8289 -11245 8299 -11211
rect 8357 -11245 8371 -11211
rect 8425 -11245 8443 -11211
rect 8493 -11245 8515 -11211
rect 8561 -11245 8587 -11211
rect 8629 -11245 8659 -11211
rect 8697 -11245 8731 -11211
rect 8765 -11245 8799 -11211
rect 8837 -11245 8867 -11211
rect 8909 -11245 8935 -11211
rect 8981 -11245 9003 -11211
rect 9053 -11245 9071 -11211
rect 9125 -11245 9139 -11211
rect 9197 -11245 9207 -11211
rect 9269 -11245 9275 -11211
rect 9341 -11245 9343 -11211
rect 9377 -11245 9379 -11211
rect 9445 -11245 9451 -11211
rect 9513 -11245 9523 -11211
rect 9581 -11245 9595 -11211
rect 9649 -11245 9667 -11211
rect 9717 -11245 9739 -11211
rect 9785 -11245 9811 -11211
rect 9853 -11245 9883 -11211
rect 9921 -11245 9955 -11211
rect 9989 -11245 10023 -11211
rect 10061 -11245 10091 -11211
rect 10133 -11245 10159 -11211
rect 10205 -11245 10227 -11211
rect 10277 -11245 10295 -11211
rect 10349 -11245 10363 -11211
rect 10421 -11245 10431 -11211
rect 10493 -11245 10499 -11211
rect 10565 -11245 10567 -11211
rect 10601 -11245 10603 -11211
rect 10669 -11245 10675 -11211
rect 10737 -11245 10747 -11211
rect 10805 -11245 10819 -11211
rect 10873 -11245 10891 -11211
rect 10941 -11245 10963 -11211
rect 11009 -11245 11035 -11211
rect 11077 -11245 11107 -11211
rect 11145 -11245 11179 -11211
rect 11213 -11245 11247 -11211
rect 11285 -11245 11315 -11211
rect 11357 -11245 11383 -11211
rect 11429 -11245 11451 -11211
rect 11501 -11245 11519 -11211
rect 11573 -11245 11587 -11211
rect 11645 -11245 11655 -11211
rect 11717 -11245 11723 -11211
rect 11789 -11245 11791 -11211
rect 11825 -11245 11827 -11211
rect 11893 -11245 11899 -11211
rect 11961 -11245 11971 -11211
rect 12029 -11245 12043 -11211
rect 12097 -11245 12115 -11211
rect 12165 -11245 12187 -11211
rect 12233 -11245 12259 -11211
rect 12301 -11245 12331 -11211
rect 12369 -11245 12403 -11211
rect 12437 -11245 12471 -11211
rect 12509 -11245 12539 -11211
rect 12581 -11245 12607 -11211
rect 12653 -11245 12675 -11211
rect 12725 -11245 12743 -11211
rect 12797 -11245 12811 -11211
rect 12869 -11245 12879 -11211
rect 12941 -11245 12947 -11211
rect 13013 -11245 13015 -11211
rect 13049 -11245 13051 -11211
rect 13117 -11245 13123 -11211
rect 13185 -11245 13195 -11211
rect 13253 -11245 13267 -11211
rect 13321 -11245 13339 -11211
rect 13389 -11245 13411 -11211
rect 13457 -11245 13483 -11211
rect 13525 -11245 13555 -11211
rect 13593 -11245 13627 -11211
rect 13661 -11245 13695 -11211
rect 13733 -11245 13763 -11211
rect 13805 -11245 13831 -11211
rect 13877 -11245 13899 -11211
rect 13949 -11245 13967 -11211
rect 14021 -11245 14035 -11211
rect 14093 -11245 14103 -11211
rect 14165 -11245 14171 -11211
rect 14237 -11245 14239 -11211
rect 14273 -11245 14275 -11211
rect 14341 -11245 14347 -11211
rect 14409 -11245 14419 -11211
rect 14477 -11245 14491 -11211
rect 14545 -11245 14563 -11211
rect 14613 -11245 14635 -11211
rect 14681 -11245 14707 -11211
rect 14749 -11245 14779 -11211
rect 14817 -11245 14851 -11211
rect 14885 -11245 14919 -11211
rect 14957 -11245 14987 -11211
rect 15029 -11245 15055 -11211
rect 15101 -11245 15123 -11211
rect 15173 -11245 15191 -11211
rect 15245 -11245 15259 -11211
rect 15317 -11245 15327 -11211
rect 15389 -11245 15395 -11211
rect 15461 -11245 15463 -11211
rect 15497 -11245 15499 -11211
rect 15565 -11245 15571 -11211
rect 15633 -11245 15643 -11211
rect 15701 -11245 15715 -11211
rect 15769 -11245 15787 -11211
rect 15837 -11245 15859 -11211
rect 15905 -11245 15931 -11211
rect 15973 -11245 16003 -11211
rect 16041 -11245 16075 -11211
rect 16109 -11245 16143 -11211
rect 16181 -11245 16211 -11211
rect 16253 -11245 16279 -11211
rect 16325 -11245 16347 -11211
rect 16397 -11245 16415 -11211
rect 16469 -11245 16483 -11211
rect 16541 -11245 16551 -11211
rect 16613 -11245 16619 -11211
rect 16685 -11245 16687 -11211
rect 16721 -11245 16723 -11211
rect 16789 -11245 16795 -11211
rect 16857 -11245 16867 -11211
rect 16925 -11245 16939 -11211
rect 16993 -11245 17011 -11211
rect 17061 -11245 17083 -11211
rect 17129 -11245 17155 -11211
rect 17197 -11245 17227 -11211
rect 17265 -11245 17299 -11211
rect 17333 -11245 17367 -11211
rect 17405 -11245 17435 -11211
rect 17477 -11245 17503 -11211
rect 17549 -11245 17571 -11211
rect 17621 -11245 17639 -11211
rect 17693 -11245 17707 -11211
rect 17765 -11245 17775 -11211
rect 17837 -11245 17843 -11211
rect 17909 -11245 17911 -11211
rect 17945 -11245 17947 -11211
rect 18013 -11245 18019 -11211
rect 18081 -11245 18091 -11211
rect 18149 -11245 18163 -11211
rect 18217 -11245 18235 -11211
rect 18285 -11245 18307 -11211
rect 18353 -11245 18379 -11211
rect 18421 -11245 18451 -11211
rect 18489 -11245 18523 -11211
rect 18557 -11245 18591 -11211
rect 18629 -11245 18659 -11211
rect 18701 -11245 18727 -11211
rect 18773 -11245 18795 -11211
rect 18845 -11245 18863 -11211
rect 18917 -11245 18931 -11211
rect 18989 -11245 18999 -11211
rect 19061 -11245 19067 -11211
rect 19133 -11245 19135 -11211
rect 19169 -11245 19171 -11211
rect 19237 -11245 19243 -11211
rect 19305 -11245 19315 -11211
rect 19373 -11245 19387 -11211
rect 19441 -11245 19459 -11211
rect 19509 -11245 19531 -11211
rect 19577 -11245 19603 -11211
rect 19645 -11245 19675 -11211
rect 19713 -11245 19747 -11211
rect 19781 -11245 19815 -11211
rect 19853 -11245 19883 -11211
rect 19925 -11245 19951 -11211
rect 19997 -11245 20019 -11211
rect 20069 -11245 20087 -11211
rect 20141 -11245 20155 -11211
rect 20213 -11245 20223 -11211
rect 20285 -11245 20291 -11211
rect 20357 -11245 20359 -11211
rect 20393 -11245 20395 -11211
rect 20461 -11245 20467 -11211
rect 20529 -11245 20539 -11211
rect 20597 -11245 20611 -11211
rect 20665 -11245 20683 -11211
rect 20733 -11245 20755 -11211
rect 20801 -11245 20827 -11211
rect 20869 -11245 20899 -11211
rect 20937 -11245 20971 -11211
rect 21005 -11245 21039 -11211
rect 21077 -11245 21107 -11211
rect 21149 -11245 21175 -11211
rect 21221 -11245 21243 -11211
rect 21293 -11245 21311 -11211
rect 21365 -11245 21379 -11211
rect 21437 -11245 21447 -11211
rect 21509 -11245 21515 -11211
rect 21581 -11245 21583 -11211
rect 21617 -11245 21619 -11211
rect 21685 -11245 21691 -11211
rect 21753 -11245 21763 -11211
rect 21821 -11245 21835 -11211
rect 21889 -11245 21907 -11211
rect 21957 -11245 21979 -11211
rect 22025 -11245 22051 -11211
rect 22093 -11245 22123 -11211
rect 22161 -11245 22195 -11211
rect 22229 -11245 22263 -11211
rect 22301 -11245 22331 -11211
rect 22373 -11245 22399 -11211
rect 22445 -11245 22467 -11211
rect 22517 -11245 22535 -11211
rect 22589 -11245 22603 -11211
rect 22661 -11245 22671 -11211
rect 22733 -11245 22739 -11211
rect 22805 -11245 22807 -11211
rect 22841 -11245 22843 -11211
rect 22909 -11245 22915 -11211
rect 22977 -11245 22987 -11211
rect 23045 -11245 23059 -11211
rect 23113 -11245 23131 -11211
rect 23181 -11245 23203 -11211
rect 23249 -11245 23275 -11211
rect 23317 -11245 23347 -11211
rect 23385 -11245 23419 -11211
rect 23453 -11245 23487 -11211
rect 23525 -11245 23555 -11211
rect 23597 -11245 23623 -11211
rect 23669 -11245 23691 -11211
rect 23741 -11245 23759 -11211
rect 23813 -11245 23827 -11211
rect 23885 -11245 23895 -11211
rect 23957 -11245 23963 -11211
rect 24029 -11245 24031 -11211
rect 24065 -11245 24067 -11211
rect 24133 -11245 24139 -11211
rect 24201 -11245 24211 -11211
rect 24269 -11245 24283 -11211
rect 24337 -11245 24355 -11211
rect 24405 -11245 24427 -11211
rect 24473 -11245 24499 -11211
rect 24541 -11245 24571 -11211
rect 24609 -11245 24643 -11211
rect 24677 -11245 24711 -11211
rect 24749 -11245 24787 -11211
rect 24821 -11245 24922 -11211
rect -12322 -11278 24922 -11245
rect -12322 -11363 -12222 -11278
rect -12322 -11397 -12289 -11363
rect -12255 -11397 -12222 -11363
rect -12322 -11431 -12222 -11397
rect -12322 -11465 -12289 -11431
rect -12255 -11465 -12222 -11431
rect -12322 -11499 -12222 -11465
rect -12322 -11533 -12289 -11499
rect -12255 -11533 -12222 -11499
rect -12322 -11567 -12222 -11533
rect -12322 -11601 -12289 -11567
rect -12255 -11601 -12222 -11567
rect -12322 -11635 -12222 -11601
rect -12322 -11669 -12289 -11635
rect -12255 -11669 -12222 -11635
rect 24822 -11363 24922 -11278
rect 24822 -11397 24855 -11363
rect 24889 -11397 24922 -11363
rect 24822 -11431 24922 -11397
rect 24822 -11465 24855 -11431
rect 24889 -11465 24922 -11431
rect 24822 -11499 24922 -11465
rect 24822 -11533 24855 -11499
rect 24889 -11533 24922 -11499
rect 24822 -11567 24922 -11533
rect 24822 -11601 24855 -11567
rect 24889 -11601 24922 -11567
rect 24822 -11635 24922 -11601
rect -12322 -11703 -12222 -11669
rect 2814 -11680 2853 -11646
rect 2887 -11680 2911 -11646
rect 2955 -11680 2983 -11646
rect 3023 -11680 3055 -11646
rect 3091 -11680 3125 -11646
rect 3161 -11680 3193 -11646
rect 3233 -11680 3261 -11646
rect 3305 -11680 3329 -11646
rect 3363 -11680 3402 -11646
rect 3848 -11680 3871 -11646
rect 3905 -11680 3929 -11646
rect 3973 -11680 4001 -11646
rect 4041 -11680 4073 -11646
rect 4109 -11680 4143 -11646
rect 4179 -11680 4211 -11646
rect 4251 -11680 4279 -11646
rect 4323 -11680 4347 -11646
rect 4381 -11680 4404 -11646
rect 4866 -11680 4889 -11646
rect 4923 -11680 4947 -11646
rect 4991 -11680 5019 -11646
rect 5059 -11680 5091 -11646
rect 5127 -11680 5161 -11646
rect 5197 -11680 5229 -11646
rect 5269 -11680 5297 -11646
rect 5341 -11680 5365 -11646
rect 5399 -11680 5422 -11646
rect 5884 -11680 5907 -11646
rect 5941 -11680 5965 -11646
rect 6009 -11680 6037 -11646
rect 6077 -11680 6109 -11646
rect 6145 -11680 6179 -11646
rect 6215 -11680 6247 -11646
rect 6287 -11680 6315 -11646
rect 6359 -11680 6383 -11646
rect 6417 -11680 6440 -11646
rect 6902 -11680 6925 -11646
rect 6959 -11680 6983 -11646
rect 7027 -11680 7055 -11646
rect 7095 -11680 7127 -11646
rect 7163 -11680 7197 -11646
rect 7233 -11680 7265 -11646
rect 7305 -11680 7333 -11646
rect 7377 -11680 7401 -11646
rect 7435 -11680 7458 -11646
rect 7920 -11680 7943 -11646
rect 7977 -11680 8001 -11646
rect 8045 -11680 8073 -11646
rect 8113 -11680 8145 -11646
rect 8181 -11680 8215 -11646
rect 8251 -11680 8283 -11646
rect 8323 -11680 8351 -11646
rect 8395 -11680 8419 -11646
rect 8453 -11680 8476 -11646
rect 8938 -11680 8961 -11646
rect 8995 -11680 9019 -11646
rect 9063 -11680 9091 -11646
rect 9131 -11680 9163 -11646
rect 9199 -11680 9233 -11646
rect 9269 -11680 9301 -11646
rect 9341 -11680 9369 -11646
rect 9413 -11680 9437 -11646
rect 9471 -11680 9494 -11646
rect 9956 -11680 9979 -11646
rect 10013 -11680 10037 -11646
rect 10081 -11680 10109 -11646
rect 10149 -11680 10181 -11646
rect 10217 -11680 10251 -11646
rect 10287 -11680 10319 -11646
rect 10359 -11680 10387 -11646
rect 10431 -11680 10455 -11646
rect 10489 -11680 10512 -11646
rect 10974 -11680 10997 -11646
rect 11031 -11680 11055 -11646
rect 11099 -11680 11127 -11646
rect 11167 -11680 11199 -11646
rect 11235 -11680 11269 -11646
rect 11305 -11680 11337 -11646
rect 11377 -11680 11405 -11646
rect 11449 -11680 11473 -11646
rect 11507 -11680 11530 -11646
rect 11992 -11680 12015 -11646
rect 12049 -11680 12073 -11646
rect 12117 -11680 12145 -11646
rect 12185 -11680 12217 -11646
rect 12253 -11680 12287 -11646
rect 12323 -11680 12355 -11646
rect 12395 -11680 12423 -11646
rect 12467 -11680 12491 -11646
rect 12525 -11680 12548 -11646
rect 13010 -11680 13033 -11646
rect 13067 -11680 13091 -11646
rect 13135 -11680 13163 -11646
rect 13203 -11680 13235 -11646
rect 13271 -11680 13305 -11646
rect 13341 -11680 13373 -11646
rect 13413 -11680 13441 -11646
rect 13485 -11680 13509 -11646
rect 13543 -11680 13566 -11646
rect 14028 -11680 14051 -11646
rect 14085 -11680 14109 -11646
rect 14153 -11680 14181 -11646
rect 14221 -11680 14253 -11646
rect 14289 -11680 14323 -11646
rect 14359 -11680 14391 -11646
rect 14431 -11680 14459 -11646
rect 14503 -11680 14527 -11646
rect 14561 -11680 14584 -11646
rect 15046 -11680 15069 -11646
rect 15103 -11680 15127 -11646
rect 15171 -11680 15199 -11646
rect 15239 -11680 15271 -11646
rect 15307 -11680 15341 -11646
rect 15377 -11680 15409 -11646
rect 15449 -11680 15477 -11646
rect 15521 -11680 15545 -11646
rect 15579 -11680 15602 -11646
rect 16064 -11680 16087 -11646
rect 16121 -11680 16145 -11646
rect 16189 -11680 16217 -11646
rect 16257 -11680 16289 -11646
rect 16325 -11680 16359 -11646
rect 16395 -11680 16427 -11646
rect 16467 -11680 16495 -11646
rect 16539 -11680 16563 -11646
rect 16597 -11680 16620 -11646
rect 17082 -11680 17105 -11646
rect 17139 -11680 17163 -11646
rect 17207 -11680 17235 -11646
rect 17275 -11680 17307 -11646
rect 17343 -11680 17377 -11646
rect 17413 -11680 17445 -11646
rect 17485 -11680 17513 -11646
rect 17557 -11680 17581 -11646
rect 17615 -11680 17638 -11646
rect 18100 -11680 18123 -11646
rect 18157 -11680 18181 -11646
rect 18225 -11680 18253 -11646
rect 18293 -11680 18325 -11646
rect 18361 -11680 18395 -11646
rect 18431 -11680 18463 -11646
rect 18503 -11680 18531 -11646
rect 18575 -11680 18599 -11646
rect 18633 -11680 18656 -11646
rect 19118 -11680 19141 -11646
rect 19175 -11680 19199 -11646
rect 19243 -11680 19271 -11646
rect 19311 -11680 19343 -11646
rect 19379 -11680 19413 -11646
rect 19449 -11680 19481 -11646
rect 19521 -11680 19549 -11646
rect 19593 -11680 19617 -11646
rect 19651 -11680 19674 -11646
rect 20136 -11680 20159 -11646
rect 20193 -11680 20217 -11646
rect 20261 -11680 20289 -11646
rect 20329 -11680 20361 -11646
rect 20397 -11680 20431 -11646
rect 20467 -11680 20499 -11646
rect 20539 -11680 20567 -11646
rect 20611 -11680 20635 -11646
rect 20669 -11680 20692 -11646
rect 21154 -11680 21177 -11646
rect 21211 -11680 21235 -11646
rect 21279 -11680 21307 -11646
rect 21347 -11680 21379 -11646
rect 21415 -11680 21449 -11646
rect 21485 -11680 21517 -11646
rect 21557 -11680 21585 -11646
rect 21629 -11680 21653 -11646
rect 21687 -11680 21710 -11646
rect 22172 -11680 22195 -11646
rect 22229 -11680 22253 -11646
rect 22297 -11680 22325 -11646
rect 22365 -11680 22397 -11646
rect 22433 -11680 22467 -11646
rect 22503 -11680 22535 -11646
rect 22575 -11680 22603 -11646
rect 22647 -11680 22671 -11646
rect 22705 -11680 22728 -11646
rect 24822 -11669 24855 -11635
rect 24889 -11669 24922 -11635
rect -12322 -11737 -12289 -11703
rect -12255 -11737 -12222 -11703
rect 24822 -11703 24922 -11669
rect -12322 -11771 -12222 -11737
rect -12322 -11805 -12289 -11771
rect -12255 -11805 -12222 -11771
rect -12322 -11839 -12222 -11805
rect -12322 -11873 -12289 -11839
rect -12255 -11873 -12222 -11839
rect -12322 -11907 -12222 -11873
rect -12322 -11941 -12289 -11907
rect -12255 -11941 -12222 -11907
rect -12322 -11975 -12222 -11941
rect -12322 -12009 -12289 -11975
rect -12255 -12009 -12222 -11975
rect -12322 -12043 -12222 -12009
rect -12322 -12077 -12289 -12043
rect -12255 -12077 -12222 -12043
rect -12322 -12091 -12222 -12077
rect -12322 -12145 -12289 -12091
rect -12255 -12145 -12222 -12091
rect -12322 -12163 -12222 -12145
rect -12322 -12213 -12289 -12163
rect -12255 -12213 -12222 -12163
rect -12322 -12235 -12222 -12213
rect -12322 -12281 -12289 -12235
rect -12255 -12281 -12222 -12235
rect -12322 -12307 -12222 -12281
rect -12322 -12349 -12289 -12307
rect -12255 -12349 -12222 -12307
rect 2582 -11749 2616 -11714
rect 2582 -11821 2616 -11797
rect 2582 -11893 2616 -11865
rect 2582 -11965 2616 -11933
rect 2582 -12035 2616 -12001
rect 2582 -12103 2616 -12071
rect 2582 -12171 2616 -12143
rect 2582 -12239 2616 -12215
rect 2582 -12322 2616 -12287
rect 3600 -11749 3634 -11730
rect 3600 -11821 3634 -11797
rect 3600 -11893 3634 -11865
rect 3600 -11965 3634 -11933
rect 3600 -12035 3634 -12001
rect 3600 -12103 3634 -12071
rect 3600 -12171 3634 -12143
rect 3600 -12239 3634 -12215
rect 3600 -12322 3634 -12287
rect 4618 -11749 4652 -11730
rect 4618 -11821 4652 -11797
rect 4618 -11893 4652 -11865
rect 4618 -11965 4652 -11933
rect 4618 -12035 4652 -12001
rect 4618 -12103 4652 -12071
rect 4618 -12171 4652 -12143
rect 4618 -12239 4652 -12215
rect 4618 -12322 4652 -12287
rect 5636 -11749 5670 -11730
rect 5636 -11821 5670 -11797
rect 5636 -11893 5670 -11865
rect 5636 -11965 5670 -11933
rect 5636 -12035 5670 -12001
rect 5636 -12103 5670 -12071
rect 5636 -12171 5670 -12143
rect 5636 -12239 5670 -12215
rect 5636 -12322 5670 -12287
rect 6654 -11749 6688 -11730
rect 6654 -11821 6688 -11797
rect 6654 -11893 6688 -11865
rect 6654 -11965 6688 -11933
rect 6654 -12035 6688 -12001
rect 6654 -12103 6688 -12071
rect 6654 -12171 6688 -12143
rect 6654 -12239 6688 -12215
rect 6654 -12322 6688 -12287
rect 7672 -11749 7706 -11730
rect 7672 -11821 7706 -11797
rect 7672 -11893 7706 -11865
rect 7672 -11965 7706 -11933
rect 7672 -12035 7706 -12001
rect 7672 -12103 7706 -12071
rect 7672 -12171 7706 -12143
rect 7672 -12239 7706 -12215
rect 7672 -12322 7706 -12287
rect 8690 -11749 8724 -11730
rect 8690 -11821 8724 -11797
rect 8690 -11893 8724 -11865
rect 8690 -11965 8724 -11933
rect 8690 -12035 8724 -12001
rect 8690 -12103 8724 -12071
rect 8690 -12171 8724 -12143
rect 8690 -12239 8724 -12215
rect 8690 -12322 8724 -12287
rect 9708 -11749 9742 -11730
rect 9708 -11821 9742 -11797
rect 9708 -11893 9742 -11865
rect 9708 -11965 9742 -11933
rect 9708 -12035 9742 -12001
rect 9708 -12103 9742 -12071
rect 9708 -12171 9742 -12143
rect 9708 -12239 9742 -12215
rect 9708 -12322 9742 -12287
rect 10726 -11749 10760 -11730
rect 10726 -11821 10760 -11797
rect 10726 -11893 10760 -11865
rect 10726 -11965 10760 -11933
rect 10726 -12035 10760 -12001
rect 10726 -12103 10760 -12071
rect 10726 -12171 10760 -12143
rect 10726 -12239 10760 -12215
rect 10726 -12322 10760 -12287
rect 11744 -11749 11778 -11730
rect 11744 -11821 11778 -11797
rect 11744 -11893 11778 -11865
rect 11744 -11965 11778 -11933
rect 11744 -12035 11778 -12001
rect 11744 -12103 11778 -12071
rect 11744 -12171 11778 -12143
rect 11744 -12239 11778 -12215
rect 11744 -12322 11778 -12287
rect 12762 -11749 12796 -11730
rect 12762 -11821 12796 -11797
rect 12762 -11893 12796 -11865
rect 12762 -11965 12796 -11933
rect 12762 -12035 12796 -12001
rect 12762 -12103 12796 -12071
rect 12762 -12171 12796 -12143
rect 12762 -12239 12796 -12215
rect 12762 -12322 12796 -12287
rect 13780 -11749 13814 -11730
rect 13780 -11821 13814 -11797
rect 13780 -11893 13814 -11865
rect 13780 -11965 13814 -11933
rect 13780 -12035 13814 -12001
rect 13780 -12103 13814 -12071
rect 13780 -12171 13814 -12143
rect 13780 -12239 13814 -12215
rect 13780 -12322 13814 -12287
rect 14798 -11749 14832 -11730
rect 14798 -11821 14832 -11797
rect 14798 -11893 14832 -11865
rect 14798 -11965 14832 -11933
rect 14798 -12035 14832 -12001
rect 14798 -12103 14832 -12071
rect 14798 -12171 14832 -12143
rect 14798 -12239 14832 -12215
rect 14798 -12322 14832 -12287
rect 15816 -11749 15850 -11730
rect 15816 -11821 15850 -11797
rect 15816 -11893 15850 -11865
rect 15816 -11965 15850 -11933
rect 15816 -12035 15850 -12001
rect 15816 -12103 15850 -12071
rect 15816 -12171 15850 -12143
rect 15816 -12239 15850 -12215
rect 15816 -12322 15850 -12287
rect 16834 -11749 16868 -11730
rect 16834 -11821 16868 -11797
rect 16834 -11893 16868 -11865
rect 16834 -11965 16868 -11933
rect 16834 -12035 16868 -12001
rect 16834 -12103 16868 -12071
rect 16834 -12171 16868 -12143
rect 16834 -12239 16868 -12215
rect 16834 -12322 16868 -12287
rect 17852 -11749 17886 -11730
rect 17852 -11821 17886 -11797
rect 17852 -11893 17886 -11865
rect 17852 -11965 17886 -11933
rect 17852 -12035 17886 -12001
rect 17852 -12103 17886 -12071
rect 17852 -12171 17886 -12143
rect 17852 -12239 17886 -12215
rect 17852 -12322 17886 -12287
rect 18870 -11749 18904 -11730
rect 18870 -11821 18904 -11797
rect 18870 -11893 18904 -11865
rect 18870 -11965 18904 -11933
rect 18870 -12035 18904 -12001
rect 18870 -12103 18904 -12071
rect 18870 -12171 18904 -12143
rect 18870 -12239 18904 -12215
rect 18870 -12322 18904 -12287
rect 19888 -11749 19922 -11730
rect 19888 -11821 19922 -11797
rect 19888 -11893 19922 -11865
rect 19888 -11965 19922 -11933
rect 19888 -12035 19922 -12001
rect 19888 -12103 19922 -12071
rect 19888 -12171 19922 -12143
rect 19888 -12239 19922 -12215
rect 19888 -12322 19922 -12287
rect 20906 -11749 20940 -11730
rect 20906 -11821 20940 -11797
rect 20906 -11893 20940 -11865
rect 20906 -11965 20940 -11933
rect 20906 -12035 20940 -12001
rect 20906 -12103 20940 -12071
rect 20906 -12171 20940 -12143
rect 20906 -12239 20940 -12215
rect 20906 -12322 20940 -12287
rect 21924 -11749 21958 -11730
rect 21924 -11821 21958 -11797
rect 21924 -11893 21958 -11865
rect 21924 -11965 21958 -11933
rect 21924 -12035 21958 -12001
rect 21924 -12103 21958 -12071
rect 21924 -12171 21958 -12143
rect 21924 -12239 21958 -12215
rect 21924 -12322 21958 -12287
rect 22942 -11749 22976 -11730
rect 22942 -11821 22976 -11797
rect 22942 -11893 22976 -11865
rect 22942 -11965 22976 -11933
rect 22942 -12035 22976 -12001
rect 22942 -12103 22976 -12071
rect 22942 -12171 22976 -12143
rect 22942 -12239 22976 -12215
rect 22942 -12322 22976 -12287
rect 24822 -11737 24855 -11703
rect 24889 -11737 24922 -11703
rect 24822 -11771 24922 -11737
rect 24822 -11805 24855 -11771
rect 24889 -11805 24922 -11771
rect 24822 -11839 24922 -11805
rect 24822 -11873 24855 -11839
rect 24889 -11873 24922 -11839
rect 24822 -11907 24922 -11873
rect 24822 -11941 24855 -11907
rect 24889 -11941 24922 -11907
rect 24822 -11975 24922 -11941
rect 24822 -12009 24855 -11975
rect 24889 -12009 24922 -11975
rect 24822 -12043 24922 -12009
rect 24822 -12077 24855 -12043
rect 24889 -12077 24922 -12043
rect 24822 -12091 24922 -12077
rect 24822 -12145 24855 -12091
rect 24889 -12145 24922 -12091
rect 24822 -12163 24922 -12145
rect 24822 -12213 24855 -12163
rect 24889 -12213 24922 -12163
rect 24822 -12235 24922 -12213
rect 24822 -12281 24855 -12235
rect 24889 -12281 24922 -12235
rect 24822 -12307 24922 -12281
rect -12322 -12379 -12222 -12349
rect 4100 -12356 4160 -12354
rect 5114 -12356 5174 -12348
rect 6118 -12356 6178 -12342
rect 7144 -12356 7204 -12354
rect 8168 -12356 8228 -12348
rect 9188 -12356 9248 -12354
rect 11214 -12356 11274 -12348
rect 12238 -12356 12298 -12354
rect 13248 -12356 13308 -12354
rect 14268 -12356 14328 -12348
rect 15298 -12356 15358 -12354
rect 16302 -12356 16362 -12348
rect 17318 -12356 17378 -12348
rect 24822 -12349 24855 -12307
rect 24889 -12349 24922 -12307
rect 18348 -12356 18408 -12354
rect 19362 -12356 19422 -12354
rect 20378 -12356 20438 -12354
rect 21404 -12356 21464 -12354
rect 22426 -12356 22486 -12354
rect -12322 -12417 -12289 -12379
rect -12255 -12417 -12222 -12379
rect 2814 -12390 2853 -12356
rect 2887 -12390 2911 -12356
rect 2955 -12390 2983 -12356
rect 3023 -12390 3055 -12356
rect 3091 -12390 3125 -12356
rect 3161 -12390 3193 -12356
rect 3233 -12390 3261 -12356
rect 3305 -12390 3329 -12356
rect 3363 -12390 3402 -12356
rect 3832 -12390 3871 -12356
rect 3905 -12390 3929 -12356
rect 3973 -12390 4001 -12356
rect 4041 -12390 4073 -12356
rect 4109 -12390 4143 -12356
rect 4179 -12390 4211 -12356
rect 4251 -12390 4279 -12356
rect 4323 -12390 4347 -12356
rect 4381 -12390 4420 -12356
rect 4850 -12390 4889 -12356
rect 4923 -12390 4947 -12356
rect 4991 -12390 5019 -12356
rect 5059 -12390 5091 -12356
rect 5127 -12390 5161 -12356
rect 5197 -12390 5229 -12356
rect 5269 -12390 5297 -12356
rect 5341 -12390 5365 -12356
rect 5399 -12390 5438 -12356
rect 5868 -12390 5907 -12356
rect 5941 -12390 5965 -12356
rect 6009 -12390 6037 -12356
rect 6077 -12390 6109 -12356
rect 6145 -12390 6179 -12356
rect 6215 -12390 6247 -12356
rect 6287 -12390 6315 -12356
rect 6359 -12390 6383 -12356
rect 6417 -12390 6456 -12356
rect 6886 -12390 6925 -12356
rect 6959 -12390 6983 -12356
rect 7027 -12390 7055 -12356
rect 7095 -12390 7127 -12356
rect 7163 -12390 7197 -12356
rect 7233 -12390 7265 -12356
rect 7305 -12390 7333 -12356
rect 7377 -12390 7401 -12356
rect 7435 -12390 7474 -12356
rect 7904 -12390 7943 -12356
rect 7977 -12390 8001 -12356
rect 8045 -12390 8073 -12356
rect 8113 -12390 8145 -12356
rect 8181 -12390 8215 -12356
rect 8251 -12390 8283 -12356
rect 8323 -12390 8351 -12356
rect 8395 -12390 8419 -12356
rect 8453 -12390 8492 -12356
rect 8922 -12390 8961 -12356
rect 8995 -12390 9019 -12356
rect 9063 -12390 9091 -12356
rect 9131 -12390 9163 -12356
rect 9199 -12390 9233 -12356
rect 9269 -12390 9301 -12356
rect 9341 -12390 9369 -12356
rect 9413 -12390 9437 -12356
rect 9471 -12390 9510 -12356
rect 9940 -12390 9979 -12356
rect 10013 -12390 10037 -12356
rect 10081 -12390 10109 -12356
rect 10149 -12390 10181 -12356
rect 10217 -12390 10251 -12356
rect 10287 -12390 10319 -12356
rect 10359 -12390 10387 -12356
rect 10431 -12390 10455 -12356
rect 10489 -12390 10528 -12356
rect 10958 -12390 10997 -12356
rect 11031 -12390 11055 -12356
rect 11099 -12390 11127 -12356
rect 11167 -12390 11199 -12356
rect 11235 -12390 11269 -12356
rect 11305 -12390 11337 -12356
rect 11377 -12390 11405 -12356
rect 11449 -12390 11473 -12356
rect 11507 -12390 11546 -12356
rect 11976 -12390 12015 -12356
rect 12049 -12390 12073 -12356
rect 12117 -12390 12145 -12356
rect 12185 -12390 12217 -12356
rect 12253 -12390 12287 -12356
rect 12323 -12390 12355 -12356
rect 12395 -12390 12423 -12356
rect 12467 -12390 12491 -12356
rect 12525 -12390 12564 -12356
rect 12994 -12390 13033 -12356
rect 13067 -12390 13091 -12356
rect 13135 -12390 13163 -12356
rect 13203 -12390 13235 -12356
rect 13271 -12390 13305 -12356
rect 13341 -12390 13373 -12356
rect 13413 -12390 13441 -12356
rect 13485 -12390 13509 -12356
rect 13543 -12390 13582 -12356
rect 14012 -12390 14051 -12356
rect 14085 -12390 14109 -12356
rect 14153 -12390 14181 -12356
rect 14221 -12390 14253 -12356
rect 14289 -12390 14323 -12356
rect 14359 -12390 14391 -12356
rect 14431 -12390 14459 -12356
rect 14503 -12390 14527 -12356
rect 14561 -12390 14600 -12356
rect 15030 -12390 15069 -12356
rect 15103 -12390 15127 -12356
rect 15171 -12390 15199 -12356
rect 15239 -12390 15271 -12356
rect 15307 -12390 15341 -12356
rect 15377 -12390 15409 -12356
rect 15449 -12390 15477 -12356
rect 15521 -12390 15545 -12356
rect 15579 -12390 15618 -12356
rect 16048 -12390 16087 -12356
rect 16121 -12390 16145 -12356
rect 16189 -12390 16217 -12356
rect 16257 -12390 16289 -12356
rect 16325 -12390 16359 -12356
rect 16395 -12390 16427 -12356
rect 16467 -12390 16495 -12356
rect 16539 -12390 16563 -12356
rect 16597 -12390 16636 -12356
rect 17066 -12390 17105 -12356
rect 17139 -12390 17163 -12356
rect 17207 -12390 17235 -12356
rect 17275 -12390 17307 -12356
rect 17343 -12390 17377 -12356
rect 17413 -12390 17445 -12356
rect 17485 -12390 17513 -12356
rect 17557 -12390 17581 -12356
rect 17615 -12390 17654 -12356
rect 18084 -12390 18123 -12356
rect 18157 -12390 18181 -12356
rect 18225 -12390 18253 -12356
rect 18293 -12390 18325 -12356
rect 18361 -12390 18395 -12356
rect 18431 -12390 18463 -12356
rect 18503 -12390 18531 -12356
rect 18575 -12390 18599 -12356
rect 18633 -12390 18672 -12356
rect 19102 -12390 19141 -12356
rect 19175 -12390 19199 -12356
rect 19243 -12390 19271 -12356
rect 19311 -12390 19343 -12356
rect 19379 -12390 19413 -12356
rect 19449 -12390 19481 -12356
rect 19521 -12390 19549 -12356
rect 19593 -12390 19617 -12356
rect 19651 -12390 19690 -12356
rect 20120 -12390 20159 -12356
rect 20193 -12390 20217 -12356
rect 20261 -12390 20289 -12356
rect 20329 -12390 20361 -12356
rect 20397 -12390 20431 -12356
rect 20467 -12390 20499 -12356
rect 20539 -12390 20567 -12356
rect 20611 -12390 20635 -12356
rect 20669 -12390 20708 -12356
rect 21138 -12390 21177 -12356
rect 21211 -12390 21235 -12356
rect 21279 -12390 21307 -12356
rect 21347 -12390 21379 -12356
rect 21415 -12390 21449 -12356
rect 21485 -12390 21517 -12356
rect 21557 -12390 21585 -12356
rect 21629 -12390 21653 -12356
rect 21687 -12390 21726 -12356
rect 22156 -12390 22195 -12356
rect 22229 -12390 22253 -12356
rect 22297 -12390 22325 -12356
rect 22365 -12390 22397 -12356
rect 22433 -12390 22467 -12356
rect 22503 -12390 22535 -12356
rect 22575 -12390 22603 -12356
rect 22647 -12390 22671 -12356
rect 22705 -12390 22744 -12356
rect 24822 -12379 24922 -12349
rect -12322 -12451 -12222 -12417
rect 24822 -12417 24855 -12379
rect 24889 -12417 24922 -12379
rect -12322 -12485 -12289 -12451
rect -12255 -12485 -12222 -12451
rect -8952 -12474 -8913 -12440
rect -8879 -12474 -8855 -12440
rect -8811 -12474 -8783 -12440
rect -8743 -12474 -8711 -12440
rect -8675 -12474 -8641 -12440
rect -8605 -12474 -8573 -12440
rect -8533 -12474 -8505 -12440
rect -8461 -12474 -8437 -12440
rect -8403 -12474 -8364 -12440
rect -7934 -12474 -7895 -12440
rect -7861 -12474 -7837 -12440
rect -7793 -12474 -7765 -12440
rect -7725 -12474 -7693 -12440
rect -7657 -12474 -7623 -12440
rect -7587 -12474 -7555 -12440
rect -7515 -12474 -7487 -12440
rect -7443 -12474 -7419 -12440
rect -7385 -12474 -7346 -12440
rect -6916 -12474 -6877 -12440
rect -6843 -12474 -6819 -12440
rect -6775 -12474 -6747 -12440
rect -6707 -12474 -6675 -12440
rect -6639 -12474 -6605 -12440
rect -6569 -12474 -6537 -12440
rect -6497 -12474 -6469 -12440
rect -6425 -12474 -6401 -12440
rect -6367 -12474 -6328 -12440
rect -5898 -12474 -5859 -12440
rect -5825 -12474 -5801 -12440
rect -5757 -12474 -5729 -12440
rect -5689 -12474 -5657 -12440
rect -5621 -12474 -5587 -12440
rect -5551 -12474 -5519 -12440
rect -5479 -12474 -5451 -12440
rect -5407 -12474 -5383 -12440
rect -5349 -12474 -5310 -12440
rect -4880 -12474 -4841 -12440
rect -4807 -12474 -4783 -12440
rect -4739 -12474 -4711 -12440
rect -4671 -12474 -4639 -12440
rect -4603 -12474 -4569 -12440
rect -4533 -12474 -4501 -12440
rect -4461 -12474 -4433 -12440
rect -4389 -12474 -4365 -12440
rect -4331 -12474 -4292 -12440
rect -3862 -12474 -3823 -12440
rect -3789 -12474 -3765 -12440
rect -3721 -12474 -3693 -12440
rect -3653 -12474 -3621 -12440
rect -3585 -12474 -3551 -12440
rect -3515 -12474 -3483 -12440
rect -3443 -12474 -3415 -12440
rect -3371 -12474 -3347 -12440
rect -3313 -12474 -3274 -12440
rect -2844 -12474 -2805 -12440
rect -2771 -12474 -2747 -12440
rect -2703 -12474 -2675 -12440
rect -2635 -12474 -2603 -12440
rect -2567 -12474 -2533 -12440
rect -2497 -12474 -2465 -12440
rect -2425 -12474 -2397 -12440
rect -2353 -12474 -2329 -12440
rect -2295 -12474 -2256 -12440
rect -1826 -12474 -1787 -12440
rect -1753 -12474 -1729 -12440
rect -1685 -12474 -1657 -12440
rect -1617 -12474 -1585 -12440
rect -1549 -12474 -1515 -12440
rect -1479 -12474 -1447 -12440
rect -1407 -12474 -1379 -12440
rect -1335 -12474 -1311 -12440
rect -1277 -12474 -1238 -12440
rect -808 -12474 -769 -12440
rect -735 -12474 -711 -12440
rect -667 -12474 -639 -12440
rect -599 -12474 -567 -12440
rect -531 -12474 -497 -12440
rect -461 -12474 -429 -12440
rect -389 -12474 -361 -12440
rect -317 -12474 -293 -12440
rect -259 -12474 -220 -12440
rect 24822 -12451 24922 -12417
rect -12322 -12519 -12222 -12485
rect 24822 -12485 24855 -12451
rect 24889 -12485 24922 -12451
rect -12322 -12557 -12289 -12519
rect -12255 -12557 -12222 -12519
rect -12322 -12587 -12222 -12557
rect -12322 -12629 -12289 -12587
rect -12255 -12629 -12222 -12587
rect -12322 -12655 -12222 -12629
rect -12322 -12701 -12289 -12655
rect -12255 -12701 -12222 -12655
rect -12322 -12723 -12222 -12701
rect -12322 -12773 -12289 -12723
rect -12255 -12773 -12222 -12723
rect -12322 -12791 -12222 -12773
rect -12322 -12845 -12289 -12791
rect -12255 -12845 -12222 -12791
rect -12322 -12859 -12222 -12845
rect -12322 -12917 -12289 -12859
rect -12255 -12917 -12222 -12859
rect -12322 -12927 -12222 -12917
rect -12322 -12989 -12289 -12927
rect -12255 -12989 -12222 -12927
rect -12322 -12995 -12222 -12989
rect -12322 -13061 -12289 -12995
rect -12255 -13061 -12222 -12995
rect -12322 -13063 -12222 -13061
rect -12322 -13097 -12289 -13063
rect -12255 -13097 -12222 -13063
rect -12322 -13099 -12222 -13097
rect -12322 -13165 -12289 -13099
rect -12255 -13165 -12222 -13099
rect -9184 -12543 -9150 -12508
rect -9184 -12615 -9150 -12591
rect -9184 -12687 -9150 -12659
rect -9184 -12759 -9150 -12727
rect -9184 -12829 -9150 -12795
rect -9184 -12897 -9150 -12865
rect -9184 -12965 -9150 -12937
rect -9184 -13033 -9150 -13009
rect -9184 -13116 -9150 -13081
rect -8166 -12543 -8132 -12508
rect -8166 -12615 -8132 -12591
rect -8166 -12687 -8132 -12659
rect -8166 -12759 -8132 -12727
rect -8166 -12829 -8132 -12795
rect -8166 -12897 -8132 -12865
rect -8166 -12965 -8132 -12937
rect -8166 -13033 -8132 -13009
rect -8166 -13116 -8132 -13081
rect -7148 -12543 -7114 -12508
rect -7148 -12615 -7114 -12591
rect -7148 -12687 -7114 -12659
rect -7148 -12759 -7114 -12727
rect -7148 -12829 -7114 -12795
rect -7148 -12897 -7114 -12865
rect -7148 -12965 -7114 -12937
rect -7148 -13033 -7114 -13009
rect -7148 -13116 -7114 -13081
rect -6130 -12543 -6096 -12508
rect -6130 -12615 -6096 -12591
rect -6130 -12687 -6096 -12659
rect -6130 -12759 -6096 -12727
rect -6130 -12829 -6096 -12795
rect -6130 -12897 -6096 -12865
rect -6130 -12965 -6096 -12937
rect -6130 -13033 -6096 -13009
rect -6130 -13116 -6096 -13081
rect -5112 -12543 -5078 -12508
rect -5112 -12615 -5078 -12591
rect -5112 -12687 -5078 -12659
rect -5112 -12759 -5078 -12727
rect -5112 -12829 -5078 -12795
rect -5112 -12897 -5078 -12865
rect -5112 -12965 -5078 -12937
rect -5112 -13033 -5078 -13009
rect -5112 -13116 -5078 -13081
rect -4094 -12543 -4060 -12508
rect -4094 -12615 -4060 -12591
rect -4094 -12687 -4060 -12659
rect -4094 -12759 -4060 -12727
rect -4094 -12829 -4060 -12795
rect -4094 -12897 -4060 -12865
rect -4094 -12965 -4060 -12937
rect -4094 -13033 -4060 -13009
rect -4094 -13116 -4060 -13081
rect -3076 -12543 -3042 -12508
rect -3076 -12615 -3042 -12591
rect -3076 -12687 -3042 -12659
rect -3076 -12759 -3042 -12727
rect -3076 -12829 -3042 -12795
rect -3076 -12897 -3042 -12865
rect -3076 -12965 -3042 -12937
rect -3076 -13033 -3042 -13009
rect -3076 -13116 -3042 -13081
rect -2058 -12543 -2024 -12508
rect -2058 -12615 -2024 -12591
rect -2058 -12687 -2024 -12659
rect -2058 -12759 -2024 -12727
rect -2058 -12829 -2024 -12795
rect -2058 -12897 -2024 -12865
rect -2058 -12965 -2024 -12937
rect -2058 -13033 -2024 -13009
rect -2058 -13116 -2024 -13081
rect -1040 -12543 -1006 -12508
rect -1040 -12615 -1006 -12591
rect -1040 -12687 -1006 -12659
rect -1040 -12759 -1006 -12727
rect -1040 -12829 -1006 -12795
rect -1040 -12897 -1006 -12865
rect -1040 -12965 -1006 -12937
rect -1040 -13033 -1006 -13009
rect -1040 -13116 -1006 -13081
rect -22 -12543 12 -12508
rect -22 -12615 12 -12591
rect -22 -12687 12 -12659
rect -22 -12759 12 -12727
rect -22 -12829 12 -12795
rect -22 -12897 12 -12865
rect 24822 -12519 24922 -12485
rect 24822 -12557 24855 -12519
rect 24889 -12557 24922 -12519
rect 24822 -12587 24922 -12557
rect 24822 -12629 24855 -12587
rect 24889 -12629 24922 -12587
rect 24822 -12655 24922 -12629
rect 24822 -12701 24855 -12655
rect 24889 -12701 24922 -12655
rect 24822 -12723 24922 -12701
rect 24822 -12773 24855 -12723
rect 24889 -12773 24922 -12723
rect 24822 -12791 24922 -12773
rect 24822 -12845 24855 -12791
rect 24889 -12845 24922 -12791
rect 24822 -12859 24922 -12845
rect 2814 -12914 2853 -12880
rect 2887 -12914 2911 -12880
rect 2955 -12914 2983 -12880
rect 3023 -12914 3055 -12880
rect 3091 -12914 3125 -12880
rect 3161 -12914 3193 -12880
rect 3233 -12914 3261 -12880
rect 3305 -12914 3329 -12880
rect 3363 -12914 3402 -12880
rect 3832 -12914 3871 -12880
rect 3905 -12914 3929 -12880
rect 3973 -12914 4001 -12880
rect 4041 -12914 4073 -12880
rect 4109 -12914 4143 -12880
rect 4179 -12914 4211 -12880
rect 4251 -12914 4279 -12880
rect 4323 -12914 4347 -12880
rect 4381 -12914 4420 -12880
rect 4850 -12914 4889 -12880
rect 4923 -12914 4947 -12880
rect 4991 -12914 5019 -12880
rect 5059 -12914 5091 -12880
rect 5127 -12914 5161 -12880
rect 5197 -12914 5229 -12880
rect 5269 -12914 5297 -12880
rect 5341 -12914 5365 -12880
rect 5399 -12914 5438 -12880
rect 5868 -12914 5907 -12880
rect 5941 -12914 5965 -12880
rect 6009 -12914 6037 -12880
rect 6077 -12914 6109 -12880
rect 6145 -12914 6179 -12880
rect 6215 -12914 6247 -12880
rect 6287 -12914 6315 -12880
rect 6359 -12914 6383 -12880
rect 6417 -12914 6456 -12880
rect 6886 -12914 6925 -12880
rect 6959 -12914 6983 -12880
rect 7027 -12914 7055 -12880
rect 7095 -12914 7127 -12880
rect 7163 -12914 7197 -12880
rect 7233 -12914 7265 -12880
rect 7305 -12914 7333 -12880
rect 7377 -12914 7401 -12880
rect 7435 -12914 7474 -12880
rect 7904 -12914 7943 -12880
rect 7977 -12914 8001 -12880
rect 8045 -12914 8073 -12880
rect 8113 -12914 8145 -12880
rect 8181 -12914 8215 -12880
rect 8251 -12914 8283 -12880
rect 8323 -12914 8351 -12880
rect 8395 -12914 8419 -12880
rect 8453 -12914 8492 -12880
rect 8922 -12914 8961 -12880
rect 8995 -12914 9019 -12880
rect 9063 -12914 9091 -12880
rect 9131 -12914 9163 -12880
rect 9199 -12914 9233 -12880
rect 9269 -12914 9301 -12880
rect 9341 -12914 9369 -12880
rect 9413 -12914 9437 -12880
rect 9471 -12914 9510 -12880
rect 9940 -12914 9979 -12880
rect 10013 -12914 10037 -12880
rect 10081 -12914 10109 -12880
rect 10149 -12914 10181 -12880
rect 10217 -12914 10251 -12880
rect 10287 -12914 10319 -12880
rect 10359 -12914 10387 -12880
rect 10431 -12914 10455 -12880
rect 10489 -12914 10528 -12880
rect 10958 -12914 10997 -12880
rect 11031 -12914 11055 -12880
rect 11099 -12914 11127 -12880
rect 11167 -12914 11199 -12880
rect 11235 -12914 11269 -12880
rect 11305 -12914 11337 -12880
rect 11377 -12914 11405 -12880
rect 11449 -12914 11473 -12880
rect 11507 -12914 11546 -12880
rect 11976 -12914 12015 -12880
rect 12049 -12914 12073 -12880
rect 12117 -12914 12145 -12880
rect 12185 -12914 12217 -12880
rect 12253 -12914 12287 -12880
rect 12323 -12914 12355 -12880
rect 12395 -12914 12423 -12880
rect 12467 -12914 12491 -12880
rect 12525 -12914 12564 -12880
rect 12994 -12914 13033 -12880
rect 13067 -12914 13091 -12880
rect 13135 -12914 13163 -12880
rect 13203 -12914 13235 -12880
rect 13271 -12914 13305 -12880
rect 13341 -12914 13373 -12880
rect 13413 -12914 13441 -12880
rect 13485 -12914 13509 -12880
rect 13543 -12914 13582 -12880
rect 14012 -12914 14051 -12880
rect 14085 -12914 14109 -12880
rect 14153 -12914 14181 -12880
rect 14221 -12914 14253 -12880
rect 14289 -12914 14323 -12880
rect 14359 -12914 14391 -12880
rect 14431 -12914 14459 -12880
rect 14503 -12914 14527 -12880
rect 14561 -12914 14600 -12880
rect 15030 -12914 15069 -12880
rect 15103 -12914 15127 -12880
rect 15171 -12914 15199 -12880
rect 15239 -12914 15271 -12880
rect 15307 -12914 15341 -12880
rect 15377 -12914 15409 -12880
rect 15449 -12914 15477 -12880
rect 15521 -12914 15545 -12880
rect 15579 -12914 15618 -12880
rect 16048 -12914 16087 -12880
rect 16121 -12914 16145 -12880
rect 16189 -12914 16217 -12880
rect 16257 -12914 16289 -12880
rect 16325 -12914 16359 -12880
rect 16395 -12914 16427 -12880
rect 16467 -12914 16495 -12880
rect 16539 -12914 16563 -12880
rect 16597 -12914 16636 -12880
rect 17066 -12914 17105 -12880
rect 17139 -12914 17163 -12880
rect 17207 -12914 17235 -12880
rect 17275 -12914 17307 -12880
rect 17343 -12914 17377 -12880
rect 17413 -12914 17445 -12880
rect 17485 -12914 17513 -12880
rect 17557 -12914 17581 -12880
rect 17615 -12914 17654 -12880
rect 18084 -12914 18123 -12880
rect 18157 -12914 18181 -12880
rect 18225 -12914 18253 -12880
rect 18293 -12914 18325 -12880
rect 18361 -12914 18395 -12880
rect 18431 -12914 18463 -12880
rect 18503 -12914 18531 -12880
rect 18575 -12914 18599 -12880
rect 18633 -12914 18672 -12880
rect 19102 -12914 19141 -12880
rect 19175 -12914 19199 -12880
rect 19243 -12914 19271 -12880
rect 19311 -12914 19343 -12880
rect 19379 -12914 19413 -12880
rect 19449 -12914 19481 -12880
rect 19521 -12914 19549 -12880
rect 19593 -12914 19617 -12880
rect 19651 -12914 19690 -12880
rect 20120 -12914 20159 -12880
rect 20193 -12914 20217 -12880
rect 20261 -12914 20289 -12880
rect 20329 -12914 20361 -12880
rect 20397 -12914 20431 -12880
rect 20467 -12914 20499 -12880
rect 20539 -12914 20567 -12880
rect 20611 -12914 20635 -12880
rect 20669 -12914 20708 -12880
rect 21138 -12914 21177 -12880
rect 21211 -12914 21235 -12880
rect 21279 -12914 21307 -12880
rect 21347 -12914 21379 -12880
rect 21415 -12914 21449 -12880
rect 21485 -12914 21517 -12880
rect 21557 -12914 21585 -12880
rect 21629 -12914 21653 -12880
rect 21687 -12914 21726 -12880
rect 22156 -12914 22195 -12880
rect 22229 -12914 22253 -12880
rect 22297 -12914 22325 -12880
rect 22365 -12914 22397 -12880
rect 22433 -12914 22467 -12880
rect 22503 -12914 22535 -12880
rect 22575 -12914 22603 -12880
rect 22647 -12914 22671 -12880
rect 22705 -12914 22744 -12880
rect 12238 -12920 12298 -12914
rect 24822 -12917 24855 -12859
rect 24889 -12917 24922 -12859
rect -22 -12965 12 -12937
rect 24822 -12927 24922 -12917
rect -22 -13033 12 -13009
rect -22 -13116 12 -13081
rect 2582 -12983 2616 -12948
rect 2582 -13055 2616 -13031
rect 2582 -13127 2616 -13099
rect -12322 -13171 -12222 -13165
rect -12322 -13233 -12289 -13171
rect -12255 -13233 -12222 -13171
rect -8952 -13184 -8913 -13150
rect -8879 -13184 -8855 -13150
rect -8811 -13184 -8783 -13150
rect -8743 -13184 -8711 -13150
rect -8675 -13184 -8641 -13150
rect -8605 -13184 -8573 -13150
rect -8533 -13184 -8505 -13150
rect -8461 -13184 -8437 -13150
rect -8403 -13184 -8364 -13150
rect -7934 -13184 -7895 -13150
rect -7861 -13184 -7837 -13150
rect -7793 -13184 -7765 -13150
rect -7725 -13184 -7693 -13150
rect -7657 -13184 -7623 -13150
rect -7587 -13184 -7555 -13150
rect -7515 -13184 -7487 -13150
rect -7443 -13184 -7419 -13150
rect -7385 -13184 -7346 -13150
rect -6916 -13184 -6877 -13150
rect -6843 -13184 -6819 -13150
rect -6775 -13184 -6747 -13150
rect -6707 -13184 -6675 -13150
rect -6639 -13184 -6605 -13150
rect -6569 -13184 -6537 -13150
rect -6497 -13184 -6469 -13150
rect -6425 -13184 -6401 -13150
rect -6367 -13184 -6328 -13150
rect -5898 -13184 -5859 -13150
rect -5825 -13184 -5801 -13150
rect -5757 -13184 -5729 -13150
rect -5689 -13184 -5657 -13150
rect -5621 -13184 -5587 -13150
rect -5551 -13184 -5519 -13150
rect -5479 -13184 -5451 -13150
rect -5407 -13184 -5383 -13150
rect -5349 -13184 -5310 -13150
rect -4880 -13184 -4841 -13150
rect -4807 -13184 -4783 -13150
rect -4739 -13184 -4711 -13150
rect -4671 -13184 -4639 -13150
rect -4603 -13184 -4569 -13150
rect -4533 -13184 -4501 -13150
rect -4461 -13184 -4433 -13150
rect -4389 -13184 -4365 -13150
rect -4331 -13184 -4292 -13150
rect -3862 -13184 -3823 -13150
rect -3789 -13184 -3765 -13150
rect -3721 -13184 -3693 -13150
rect -3653 -13184 -3621 -13150
rect -3585 -13184 -3551 -13150
rect -3515 -13184 -3483 -13150
rect -3443 -13184 -3415 -13150
rect -3371 -13184 -3347 -13150
rect -3313 -13184 -3274 -13150
rect -2844 -13184 -2805 -13150
rect -2771 -13184 -2747 -13150
rect -2703 -13184 -2675 -13150
rect -2635 -13184 -2603 -13150
rect -2567 -13184 -2533 -13150
rect -2497 -13184 -2465 -13150
rect -2425 -13184 -2397 -13150
rect -2353 -13184 -2329 -13150
rect -2295 -13184 -2256 -13150
rect -1826 -13184 -1787 -13150
rect -1753 -13184 -1729 -13150
rect -1685 -13184 -1657 -13150
rect -1617 -13184 -1585 -13150
rect -1549 -13184 -1515 -13150
rect -1479 -13184 -1447 -13150
rect -1407 -13184 -1379 -13150
rect -1335 -13184 -1311 -13150
rect -1277 -13184 -1238 -13150
rect -808 -13184 -769 -13150
rect -735 -13184 -711 -13150
rect -667 -13184 -639 -13150
rect -599 -13184 -567 -13150
rect -531 -13184 -497 -13150
rect -461 -13184 -429 -13150
rect -389 -13184 -361 -13150
rect -317 -13184 -293 -13150
rect -259 -13184 -220 -13150
rect -12322 -13243 -12222 -13233
rect -12322 -13301 -12289 -13243
rect -12255 -13301 -12222 -13243
rect 2582 -13199 2616 -13167
rect -8952 -13292 -8913 -13258
rect -8879 -13292 -8855 -13258
rect -8811 -13292 -8783 -13258
rect -8743 -13292 -8711 -13258
rect -8675 -13292 -8641 -13258
rect -8605 -13292 -8573 -13258
rect -8533 -13292 -8505 -13258
rect -8461 -13292 -8437 -13258
rect -8403 -13292 -8364 -13258
rect -7934 -13292 -7895 -13258
rect -7861 -13292 -7837 -13258
rect -7793 -13292 -7765 -13258
rect -7725 -13292 -7693 -13258
rect -7657 -13292 -7623 -13258
rect -7587 -13292 -7555 -13258
rect -7515 -13292 -7487 -13258
rect -7443 -13292 -7419 -13258
rect -7385 -13292 -7346 -13258
rect -6916 -13292 -6877 -13258
rect -6843 -13292 -6819 -13258
rect -6775 -13292 -6747 -13258
rect -6707 -13292 -6675 -13258
rect -6639 -13292 -6605 -13258
rect -6569 -13292 -6537 -13258
rect -6497 -13292 -6469 -13258
rect -6425 -13292 -6401 -13258
rect -6367 -13292 -6328 -13258
rect -5898 -13292 -5859 -13258
rect -5825 -13292 -5801 -13258
rect -5757 -13292 -5729 -13258
rect -5689 -13292 -5657 -13258
rect -5621 -13292 -5587 -13258
rect -5551 -13292 -5519 -13258
rect -5479 -13292 -5451 -13258
rect -5407 -13292 -5383 -13258
rect -5349 -13292 -5310 -13258
rect -4880 -13292 -4841 -13258
rect -4807 -13292 -4783 -13258
rect -4739 -13292 -4711 -13258
rect -4671 -13292 -4639 -13258
rect -4603 -13292 -4569 -13258
rect -4533 -13292 -4501 -13258
rect -4461 -13292 -4433 -13258
rect -4389 -13292 -4365 -13258
rect -4331 -13292 -4292 -13258
rect -3862 -13292 -3823 -13258
rect -3789 -13292 -3765 -13258
rect -3721 -13292 -3693 -13258
rect -3653 -13292 -3621 -13258
rect -3585 -13292 -3551 -13258
rect -3515 -13292 -3483 -13258
rect -3443 -13292 -3415 -13258
rect -3371 -13292 -3347 -13258
rect -3313 -13292 -3274 -13258
rect -2844 -13292 -2805 -13258
rect -2771 -13292 -2747 -13258
rect -2703 -13292 -2675 -13258
rect -2635 -13292 -2603 -13258
rect -2567 -13292 -2533 -13258
rect -2497 -13292 -2465 -13258
rect -2425 -13292 -2397 -13258
rect -2353 -13292 -2329 -13258
rect -2295 -13292 -2256 -13258
rect -1826 -13292 -1787 -13258
rect -1753 -13292 -1729 -13258
rect -1685 -13292 -1657 -13258
rect -1617 -13292 -1585 -13258
rect -1549 -13292 -1515 -13258
rect -1479 -13292 -1447 -13258
rect -1407 -13292 -1379 -13258
rect -1335 -13292 -1311 -13258
rect -1277 -13292 -1238 -13258
rect -808 -13292 -769 -13258
rect -735 -13292 -711 -13258
rect -667 -13292 -639 -13258
rect -599 -13292 -567 -13258
rect -531 -13292 -497 -13258
rect -461 -13292 -429 -13258
rect -389 -13292 -361 -13258
rect -317 -13292 -293 -13258
rect -259 -13292 -220 -13258
rect 2582 -13269 2616 -13235
rect -3592 -13294 -3532 -13292
rect -12322 -13315 -12222 -13301
rect -12322 -13369 -12289 -13315
rect -12255 -13369 -12222 -13315
rect -12322 -13387 -12222 -13369
rect -12322 -13437 -12289 -13387
rect -12255 -13437 -12222 -13387
rect -12322 -13459 -12222 -13437
rect -12322 -13505 -12289 -13459
rect -12255 -13505 -12222 -13459
rect -12322 -13531 -12222 -13505
rect -12322 -13573 -12289 -13531
rect -12255 -13573 -12222 -13531
rect -12322 -13603 -12222 -13573
rect -12322 -13641 -12289 -13603
rect -12255 -13641 -12222 -13603
rect -12322 -13675 -12222 -13641
rect -12322 -13709 -12289 -13675
rect -12255 -13709 -12222 -13675
rect -12322 -13743 -12222 -13709
rect -12322 -13781 -12289 -13743
rect -12255 -13781 -12222 -13743
rect -12322 -13811 -12222 -13781
rect -12322 -13853 -12289 -13811
rect -12255 -13853 -12222 -13811
rect -12322 -13879 -12222 -13853
rect -12322 -13925 -12289 -13879
rect -12255 -13925 -12222 -13879
rect -12322 -13947 -12222 -13925
rect -9184 -13361 -9150 -13326
rect -9184 -13433 -9150 -13409
rect -9184 -13505 -9150 -13477
rect -9184 -13577 -9150 -13545
rect -9184 -13647 -9150 -13613
rect -9184 -13715 -9150 -13683
rect -9184 -13783 -9150 -13755
rect -9184 -13851 -9150 -13827
rect -9184 -13934 -9150 -13899
rect -8166 -13361 -8132 -13326
rect -8166 -13433 -8132 -13409
rect -8166 -13505 -8132 -13477
rect -8166 -13577 -8132 -13545
rect -8166 -13647 -8132 -13613
rect -8166 -13715 -8132 -13683
rect -8166 -13783 -8132 -13755
rect -8166 -13851 -8132 -13827
rect -8166 -13934 -8132 -13899
rect -7148 -13361 -7114 -13326
rect -7148 -13433 -7114 -13409
rect -7148 -13505 -7114 -13477
rect -7148 -13577 -7114 -13545
rect -7148 -13647 -7114 -13613
rect -7148 -13715 -7114 -13683
rect -7148 -13783 -7114 -13755
rect -7148 -13851 -7114 -13827
rect -7148 -13934 -7114 -13899
rect -6130 -13361 -6096 -13326
rect -6130 -13433 -6096 -13409
rect -6130 -13505 -6096 -13477
rect -6130 -13577 -6096 -13545
rect -6130 -13647 -6096 -13613
rect -6130 -13715 -6096 -13683
rect -6130 -13783 -6096 -13755
rect -6130 -13851 -6096 -13827
rect -6130 -13934 -6096 -13899
rect -5112 -13361 -5078 -13326
rect -5112 -13433 -5078 -13409
rect -5112 -13505 -5078 -13477
rect -5112 -13577 -5078 -13545
rect -5112 -13647 -5078 -13613
rect -5112 -13715 -5078 -13683
rect -5112 -13783 -5078 -13755
rect -5112 -13851 -5078 -13827
rect -5112 -13934 -5078 -13899
rect -4094 -13361 -4060 -13326
rect -4094 -13433 -4060 -13409
rect -4094 -13505 -4060 -13477
rect -4094 -13577 -4060 -13545
rect -4094 -13647 -4060 -13613
rect -4094 -13715 -4060 -13683
rect -4094 -13783 -4060 -13755
rect -4094 -13851 -4060 -13827
rect -4094 -13934 -4060 -13899
rect -3076 -13361 -3042 -13326
rect -3076 -13433 -3042 -13409
rect -3076 -13505 -3042 -13477
rect -3076 -13577 -3042 -13545
rect -3076 -13647 -3042 -13613
rect -3076 -13715 -3042 -13683
rect -3076 -13783 -3042 -13755
rect -3076 -13851 -3042 -13827
rect -3076 -13934 -3042 -13899
rect -2058 -13361 -2024 -13326
rect -2058 -13433 -2024 -13409
rect -2058 -13505 -2024 -13477
rect -2058 -13577 -2024 -13545
rect -2058 -13647 -2024 -13613
rect -2058 -13715 -2024 -13683
rect -2058 -13783 -2024 -13755
rect -2058 -13851 -2024 -13827
rect -2058 -13934 -2024 -13899
rect -1040 -13361 -1006 -13326
rect -1040 -13433 -1006 -13409
rect -1040 -13505 -1006 -13477
rect -1040 -13577 -1006 -13545
rect -1040 -13647 -1006 -13613
rect -1040 -13715 -1006 -13683
rect -1040 -13783 -1006 -13755
rect -1040 -13851 -1006 -13827
rect -1040 -13934 -1006 -13899
rect -22 -13361 12 -13326
rect -22 -13433 12 -13409
rect -22 -13505 12 -13477
rect -22 -13577 12 -13545
rect 2582 -13337 2616 -13305
rect 2582 -13405 2616 -13377
rect 2582 -13473 2616 -13449
rect 2582 -13556 2616 -13521
rect 3600 -12983 3634 -12948
rect 3600 -13055 3634 -13031
rect 3600 -13127 3634 -13099
rect 3600 -13199 3634 -13167
rect 3600 -13269 3634 -13235
rect 3600 -13337 3634 -13305
rect 3600 -13405 3634 -13377
rect 3600 -13473 3634 -13449
rect 3600 -13556 3634 -13521
rect 4618 -12983 4652 -12948
rect 4618 -13055 4652 -13031
rect 4618 -13127 4652 -13099
rect 4618 -13199 4652 -13167
rect 4618 -13269 4652 -13235
rect 4618 -13337 4652 -13305
rect 4618 -13405 4652 -13377
rect 4618 -13473 4652 -13449
rect 4618 -13556 4652 -13521
rect 5636 -12983 5670 -12948
rect 5636 -13055 5670 -13031
rect 5636 -13127 5670 -13099
rect 5636 -13199 5670 -13167
rect 5636 -13269 5670 -13235
rect 5636 -13337 5670 -13305
rect 5636 -13405 5670 -13377
rect 5636 -13473 5670 -13449
rect 5636 -13556 5670 -13521
rect 6654 -12983 6688 -12948
rect 6654 -13055 6688 -13031
rect 6654 -13127 6688 -13099
rect 6654 -13199 6688 -13167
rect 6654 -13269 6688 -13235
rect 6654 -13337 6688 -13305
rect 6654 -13405 6688 -13377
rect 6654 -13473 6688 -13449
rect 6654 -13556 6688 -13521
rect 7672 -12983 7706 -12948
rect 7672 -13055 7706 -13031
rect 7672 -13127 7706 -13099
rect 7672 -13199 7706 -13167
rect 7672 -13269 7706 -13235
rect 7672 -13337 7706 -13305
rect 7672 -13405 7706 -13377
rect 7672 -13473 7706 -13449
rect 7672 -13556 7706 -13521
rect 8690 -12983 8724 -12948
rect 8690 -13055 8724 -13031
rect 8690 -13127 8724 -13099
rect 8690 -13199 8724 -13167
rect 8690 -13269 8724 -13235
rect 8690 -13337 8724 -13305
rect 8690 -13405 8724 -13377
rect 8690 -13473 8724 -13449
rect 8690 -13556 8724 -13521
rect 9708 -12983 9742 -12948
rect 9708 -13055 9742 -13031
rect 9708 -13127 9742 -13099
rect 9708 -13199 9742 -13167
rect 9708 -13269 9742 -13235
rect 9708 -13337 9742 -13305
rect 9708 -13405 9742 -13377
rect 9708 -13473 9742 -13449
rect 9708 -13556 9742 -13521
rect 10726 -12983 10760 -12948
rect 10726 -13055 10760 -13031
rect 10726 -13127 10760 -13099
rect 10726 -13199 10760 -13167
rect 10726 -13269 10760 -13235
rect 10726 -13337 10760 -13305
rect 10726 -13405 10760 -13377
rect 10726 -13473 10760 -13449
rect 10726 -13556 10760 -13521
rect 11744 -12983 11778 -12948
rect 11744 -13055 11778 -13031
rect 11744 -13127 11778 -13099
rect 11744 -13199 11778 -13167
rect 11744 -13269 11778 -13235
rect 11744 -13337 11778 -13305
rect 11744 -13405 11778 -13377
rect 11744 -13473 11778 -13449
rect 11744 -13556 11778 -13521
rect 12762 -12983 12796 -12948
rect 12762 -13055 12796 -13031
rect 12762 -13127 12796 -13099
rect 12762 -13199 12796 -13167
rect 12762 -13269 12796 -13235
rect 12762 -13337 12796 -13305
rect 12762 -13405 12796 -13377
rect 12762 -13473 12796 -13449
rect 12762 -13556 12796 -13521
rect 13780 -12983 13814 -12948
rect 13780 -13055 13814 -13031
rect 13780 -13127 13814 -13099
rect 13780 -13199 13814 -13167
rect 13780 -13269 13814 -13235
rect 13780 -13337 13814 -13305
rect 13780 -13405 13814 -13377
rect 13780 -13473 13814 -13449
rect 13780 -13556 13814 -13521
rect 14798 -12983 14832 -12948
rect 14798 -13055 14832 -13031
rect 14798 -13127 14832 -13099
rect 14798 -13199 14832 -13167
rect 14798 -13269 14832 -13235
rect 14798 -13337 14832 -13305
rect 14798 -13405 14832 -13377
rect 14798 -13473 14832 -13449
rect 14798 -13556 14832 -13521
rect 15816 -12983 15850 -12948
rect 15816 -13055 15850 -13031
rect 15816 -13127 15850 -13099
rect 15816 -13199 15850 -13167
rect 15816 -13269 15850 -13235
rect 15816 -13337 15850 -13305
rect 15816 -13405 15850 -13377
rect 15816 -13473 15850 -13449
rect 15816 -13556 15850 -13521
rect 16834 -12983 16868 -12948
rect 16834 -13055 16868 -13031
rect 16834 -13127 16868 -13099
rect 16834 -13199 16868 -13167
rect 16834 -13269 16868 -13235
rect 16834 -13337 16868 -13305
rect 16834 -13405 16868 -13377
rect 16834 -13473 16868 -13449
rect 16834 -13556 16868 -13521
rect 17852 -12983 17886 -12948
rect 17852 -13055 17886 -13031
rect 17852 -13127 17886 -13099
rect 17852 -13199 17886 -13167
rect 17852 -13269 17886 -13235
rect 17852 -13337 17886 -13305
rect 17852 -13405 17886 -13377
rect 17852 -13473 17886 -13449
rect 17852 -13556 17886 -13521
rect 18870 -12983 18904 -12948
rect 18870 -13055 18904 -13031
rect 18870 -13127 18904 -13099
rect 18870 -13199 18904 -13167
rect 18870 -13269 18904 -13235
rect 18870 -13337 18904 -13305
rect 18870 -13405 18904 -13377
rect 18870 -13473 18904 -13449
rect 18870 -13556 18904 -13521
rect 19888 -12983 19922 -12948
rect 19888 -13055 19922 -13031
rect 19888 -13127 19922 -13099
rect 19888 -13199 19922 -13167
rect 19888 -13269 19922 -13235
rect 19888 -13337 19922 -13305
rect 19888 -13405 19922 -13377
rect 19888 -13473 19922 -13449
rect 19888 -13556 19922 -13521
rect 20906 -12983 20940 -12948
rect 20906 -13055 20940 -13031
rect 20906 -13127 20940 -13099
rect 20906 -13199 20940 -13167
rect 20906 -13269 20940 -13235
rect 20906 -13337 20940 -13305
rect 20906 -13405 20940 -13377
rect 20906 -13473 20940 -13449
rect 20906 -13556 20940 -13521
rect 21924 -12983 21958 -12948
rect 21924 -13055 21958 -13031
rect 21924 -13127 21958 -13099
rect 21924 -13199 21958 -13167
rect 21924 -13269 21958 -13235
rect 21924 -13337 21958 -13305
rect 21924 -13405 21958 -13377
rect 21924 -13473 21958 -13449
rect 21924 -13556 21958 -13521
rect 22942 -12983 22976 -12948
rect 22942 -13055 22976 -13031
rect 22942 -13127 22976 -13099
rect 22942 -13199 22976 -13167
rect 22942 -13269 22976 -13235
rect 22942 -13337 22976 -13305
rect 22942 -13405 22976 -13377
rect 22942 -13473 22976 -13449
rect 22942 -13556 22976 -13521
rect 24822 -12989 24855 -12927
rect 24889 -12989 24922 -12927
rect 24822 -12995 24922 -12989
rect 24822 -13061 24855 -12995
rect 24889 -13061 24922 -12995
rect 24822 -13063 24922 -13061
rect 24822 -13097 24855 -13063
rect 24889 -13097 24922 -13063
rect 24822 -13099 24922 -13097
rect 24822 -13165 24855 -13099
rect 24889 -13165 24922 -13099
rect 24822 -13171 24922 -13165
rect 24822 -13233 24855 -13171
rect 24889 -13233 24922 -13171
rect 24822 -13243 24922 -13233
rect 24822 -13301 24855 -13243
rect 24889 -13301 24922 -13243
rect 24822 -13315 24922 -13301
rect 24822 -13369 24855 -13315
rect 24889 -13369 24922 -13315
rect 24822 -13387 24922 -13369
rect 24822 -13437 24855 -13387
rect 24889 -13437 24922 -13387
rect 24822 -13459 24922 -13437
rect 24822 -13505 24855 -13459
rect 24889 -13505 24922 -13459
rect 24822 -13531 24922 -13505
rect 24822 -13573 24855 -13531
rect 24889 -13573 24922 -13531
rect 8166 -13590 8226 -13584
rect 10202 -13590 10262 -13584
rect 11222 -13590 11282 -13584
rect 16294 -13590 16354 -13584
rect -22 -13647 12 -13613
rect 2814 -13624 2853 -13590
rect 2887 -13624 2911 -13590
rect 2955 -13624 2983 -13590
rect 3023 -13624 3055 -13590
rect 3091 -13624 3125 -13590
rect 3161 -13624 3193 -13590
rect 3233 -13624 3261 -13590
rect 3305 -13624 3329 -13590
rect 3363 -13624 3402 -13590
rect 3832 -13624 3871 -13590
rect 3905 -13624 3929 -13590
rect 3973 -13624 4001 -13590
rect 4041 -13624 4073 -13590
rect 4109 -13624 4143 -13590
rect 4179 -13624 4211 -13590
rect 4251 -13624 4279 -13590
rect 4323 -13624 4347 -13590
rect 4381 -13624 4420 -13590
rect 4850 -13624 4889 -13590
rect 4923 -13624 4947 -13590
rect 4991 -13624 5019 -13590
rect 5059 -13624 5091 -13590
rect 5127 -13624 5161 -13590
rect 5197 -13624 5229 -13590
rect 5269 -13624 5297 -13590
rect 5341 -13624 5365 -13590
rect 5399 -13624 5438 -13590
rect 5868 -13624 5907 -13590
rect 5941 -13624 5965 -13590
rect 6009 -13624 6037 -13590
rect 6077 -13624 6109 -13590
rect 6145 -13624 6179 -13590
rect 6215 -13624 6247 -13590
rect 6287 -13624 6315 -13590
rect 6359 -13624 6383 -13590
rect 6417 -13624 6456 -13590
rect 6886 -13624 6925 -13590
rect 6959 -13624 6983 -13590
rect 7027 -13624 7055 -13590
rect 7095 -13624 7127 -13590
rect 7163 -13624 7197 -13590
rect 7233 -13624 7265 -13590
rect 7305 -13624 7333 -13590
rect 7377 -13624 7401 -13590
rect 7435 -13624 7474 -13590
rect 7904 -13624 7943 -13590
rect 7977 -13624 8001 -13590
rect 8045 -13624 8073 -13590
rect 8113 -13624 8145 -13590
rect 8181 -13624 8215 -13590
rect 8251 -13624 8283 -13590
rect 8323 -13624 8351 -13590
rect 8395 -13624 8419 -13590
rect 8453 -13624 8492 -13590
rect 8922 -13624 8961 -13590
rect 8995 -13624 9019 -13590
rect 9063 -13624 9091 -13590
rect 9131 -13624 9163 -13590
rect 9199 -13624 9233 -13590
rect 9269 -13624 9301 -13590
rect 9341 -13624 9369 -13590
rect 9413 -13624 9437 -13590
rect 9471 -13624 9510 -13590
rect 9940 -13624 9979 -13590
rect 10013 -13624 10037 -13590
rect 10081 -13624 10109 -13590
rect 10149 -13624 10181 -13590
rect 10217 -13624 10251 -13590
rect 10287 -13624 10319 -13590
rect 10359 -13624 10387 -13590
rect 10431 -13624 10455 -13590
rect 10489 -13624 10528 -13590
rect 10958 -13624 10997 -13590
rect 11031 -13624 11055 -13590
rect 11099 -13624 11127 -13590
rect 11167 -13624 11199 -13590
rect 11235 -13624 11269 -13590
rect 11305 -13624 11337 -13590
rect 11377 -13624 11405 -13590
rect 11449 -13624 11473 -13590
rect 11507 -13624 11546 -13590
rect 11976 -13624 12015 -13590
rect 12049 -13624 12073 -13590
rect 12117 -13624 12145 -13590
rect 12185 -13624 12217 -13590
rect 12253 -13624 12287 -13590
rect 12323 -13624 12355 -13590
rect 12395 -13624 12423 -13590
rect 12467 -13624 12491 -13590
rect 12525 -13624 12564 -13590
rect 12994 -13624 13033 -13590
rect 13067 -13624 13091 -13590
rect 13135 -13624 13163 -13590
rect 13203 -13624 13235 -13590
rect 13271 -13624 13305 -13590
rect 13341 -13624 13373 -13590
rect 13413 -13624 13441 -13590
rect 13485 -13624 13509 -13590
rect 13543 -13624 13582 -13590
rect 14012 -13624 14051 -13590
rect 14085 -13624 14109 -13590
rect 14153 -13624 14181 -13590
rect 14221 -13624 14253 -13590
rect 14289 -13624 14323 -13590
rect 14359 -13624 14391 -13590
rect 14431 -13624 14459 -13590
rect 14503 -13624 14527 -13590
rect 14561 -13624 14600 -13590
rect 15030 -13624 15069 -13590
rect 15103 -13624 15127 -13590
rect 15171 -13624 15199 -13590
rect 15239 -13624 15271 -13590
rect 15307 -13624 15341 -13590
rect 15377 -13624 15409 -13590
rect 15449 -13624 15477 -13590
rect 15521 -13624 15545 -13590
rect 15579 -13624 15618 -13590
rect 16048 -13624 16087 -13590
rect 16121 -13624 16145 -13590
rect 16189 -13624 16217 -13590
rect 16257 -13624 16289 -13590
rect 16325 -13624 16359 -13590
rect 16395 -13624 16427 -13590
rect 16467 -13624 16495 -13590
rect 16539 -13624 16563 -13590
rect 16597 -13624 16636 -13590
rect 17066 -13624 17105 -13590
rect 17139 -13624 17163 -13590
rect 17207 -13624 17235 -13590
rect 17275 -13624 17307 -13590
rect 17343 -13624 17377 -13590
rect 17413 -13624 17445 -13590
rect 17485 -13624 17513 -13590
rect 17557 -13624 17581 -13590
rect 17615 -13624 17654 -13590
rect 18084 -13624 18123 -13590
rect 18157 -13624 18181 -13590
rect 18225 -13624 18253 -13590
rect 18293 -13624 18325 -13590
rect 18361 -13624 18395 -13590
rect 18431 -13624 18463 -13590
rect 18503 -13624 18531 -13590
rect 18575 -13624 18599 -13590
rect 18633 -13624 18672 -13590
rect 19102 -13624 19141 -13590
rect 19175 -13624 19199 -13590
rect 19243 -13624 19271 -13590
rect 19311 -13624 19343 -13590
rect 19379 -13624 19413 -13590
rect 19449 -13624 19481 -13590
rect 19521 -13624 19549 -13590
rect 19593 -13624 19617 -13590
rect 19651 -13624 19690 -13590
rect 20120 -13624 20159 -13590
rect 20193 -13624 20217 -13590
rect 20261 -13624 20289 -13590
rect 20329 -13624 20361 -13590
rect 20397 -13624 20431 -13590
rect 20467 -13624 20499 -13590
rect 20539 -13624 20567 -13590
rect 20611 -13624 20635 -13590
rect 20669 -13624 20708 -13590
rect 21138 -13624 21177 -13590
rect 21211 -13624 21235 -13590
rect 21279 -13624 21307 -13590
rect 21347 -13624 21379 -13590
rect 21415 -13624 21449 -13590
rect 21485 -13624 21517 -13590
rect 21557 -13624 21585 -13590
rect 21629 -13624 21653 -13590
rect 21687 -13624 21726 -13590
rect 22156 -13624 22195 -13590
rect 22229 -13624 22253 -13590
rect 22297 -13624 22325 -13590
rect 22365 -13624 22397 -13590
rect 22433 -13624 22467 -13590
rect 22503 -13624 22535 -13590
rect 22575 -13624 22603 -13590
rect 22647 -13624 22671 -13590
rect 22705 -13624 22744 -13590
rect 24822 -13603 24922 -13573
rect -22 -13715 12 -13683
rect -22 -13783 12 -13755
rect -22 -13851 12 -13827
rect -22 -13934 12 -13899
rect 24822 -13641 24855 -13603
rect 24889 -13641 24922 -13603
rect 24822 -13675 24922 -13641
rect 24822 -13709 24855 -13675
rect 24889 -13709 24922 -13675
rect 24822 -13743 24922 -13709
rect 24822 -13781 24855 -13743
rect 24889 -13781 24922 -13743
rect 24822 -13811 24922 -13781
rect 24822 -13853 24855 -13811
rect 24889 -13853 24922 -13811
rect 24822 -13879 24922 -13853
rect 24822 -13925 24855 -13879
rect 24889 -13925 24922 -13879
rect -12322 -13997 -12289 -13947
rect -12255 -13997 -12222 -13947
rect 24822 -13947 24922 -13925
rect -7660 -13968 -7600 -13966
rect -6646 -13968 -6586 -13966
rect -2572 -13968 -2512 -13966
rect -1556 -13968 -1496 -13966
rect -12322 -14015 -12222 -13997
rect -8952 -14002 -8913 -13968
rect -8879 -14002 -8855 -13968
rect -8811 -14002 -8783 -13968
rect -8743 -14002 -8711 -13968
rect -8675 -14002 -8641 -13968
rect -8605 -14002 -8573 -13968
rect -8533 -14002 -8505 -13968
rect -8461 -14002 -8437 -13968
rect -8403 -14002 -8364 -13968
rect -7934 -14002 -7895 -13968
rect -7861 -14002 -7837 -13968
rect -7793 -14002 -7765 -13968
rect -7725 -14002 -7693 -13968
rect -7657 -14002 -7623 -13968
rect -7587 -14002 -7555 -13968
rect -7515 -14002 -7487 -13968
rect -7443 -14002 -7419 -13968
rect -7385 -14002 -7346 -13968
rect -6916 -14002 -6877 -13968
rect -6843 -14002 -6819 -13968
rect -6775 -14002 -6747 -13968
rect -6707 -14002 -6675 -13968
rect -6639 -14002 -6605 -13968
rect -6569 -14002 -6537 -13968
rect -6497 -14002 -6469 -13968
rect -6425 -14002 -6401 -13968
rect -6367 -14002 -6328 -13968
rect -5898 -14002 -5859 -13968
rect -5825 -14002 -5801 -13968
rect -5757 -14002 -5729 -13968
rect -5689 -14002 -5657 -13968
rect -5621 -14002 -5587 -13968
rect -5551 -14002 -5519 -13968
rect -5479 -14002 -5451 -13968
rect -5407 -14002 -5383 -13968
rect -5349 -14002 -5310 -13968
rect -4880 -14002 -4841 -13968
rect -4807 -14002 -4783 -13968
rect -4739 -14002 -4711 -13968
rect -4671 -14002 -4639 -13968
rect -4603 -14002 -4569 -13968
rect -4533 -14002 -4501 -13968
rect -4461 -14002 -4433 -13968
rect -4389 -14002 -4365 -13968
rect -4331 -14002 -4292 -13968
rect -3862 -14002 -3823 -13968
rect -3789 -14002 -3765 -13968
rect -3721 -14002 -3693 -13968
rect -3653 -14002 -3621 -13968
rect -3585 -14002 -3551 -13968
rect -3515 -14002 -3483 -13968
rect -3443 -14002 -3415 -13968
rect -3371 -14002 -3347 -13968
rect -3313 -14002 -3274 -13968
rect -2844 -14002 -2805 -13968
rect -2771 -14002 -2747 -13968
rect -2703 -14002 -2675 -13968
rect -2635 -14002 -2603 -13968
rect -2567 -14002 -2533 -13968
rect -2497 -14002 -2465 -13968
rect -2425 -14002 -2397 -13968
rect -2353 -14002 -2329 -13968
rect -2295 -14002 -2256 -13968
rect -1826 -14002 -1787 -13968
rect -1753 -14002 -1729 -13968
rect -1685 -14002 -1657 -13968
rect -1617 -14002 -1585 -13968
rect -1549 -14002 -1515 -13968
rect -1479 -14002 -1447 -13968
rect -1407 -14002 -1379 -13968
rect -1335 -14002 -1311 -13968
rect -1277 -14002 -1238 -13968
rect -808 -14002 -769 -13968
rect -735 -14002 -711 -13968
rect -667 -14002 -639 -13968
rect -599 -14002 -567 -13968
rect -531 -14002 -497 -13968
rect -461 -14002 -429 -13968
rect -389 -14002 -361 -13968
rect -317 -14002 -293 -13968
rect -259 -14002 -220 -13968
rect 24822 -13997 24855 -13947
rect 24889 -13997 24922 -13947
rect -12322 -14069 -12289 -14015
rect -12255 -14069 -12222 -14015
rect -12322 -14083 -12222 -14069
rect 24822 -14015 24922 -13997
rect 24822 -14069 24855 -14015
rect 24889 -14069 24922 -14015
rect -12322 -14141 -12289 -14083
rect -12255 -14141 -12222 -14083
rect -8952 -14110 -8913 -14076
rect -8879 -14110 -8855 -14076
rect -8811 -14110 -8783 -14076
rect -8743 -14110 -8711 -14076
rect -8675 -14110 -8641 -14076
rect -8605 -14110 -8573 -14076
rect -8533 -14110 -8505 -14076
rect -8461 -14110 -8437 -14076
rect -8403 -14110 -8364 -14076
rect -7934 -14110 -7895 -14076
rect -7861 -14110 -7837 -14076
rect -7793 -14110 -7765 -14076
rect -7725 -14110 -7693 -14076
rect -7657 -14110 -7623 -14076
rect -7587 -14110 -7555 -14076
rect -7515 -14110 -7487 -14076
rect -7443 -14110 -7419 -14076
rect -7385 -14110 -7346 -14076
rect -6916 -14110 -6877 -14076
rect -6843 -14110 -6819 -14076
rect -6775 -14110 -6747 -14076
rect -6707 -14110 -6675 -14076
rect -6639 -14110 -6605 -14076
rect -6569 -14110 -6537 -14076
rect -6497 -14110 -6469 -14076
rect -6425 -14110 -6401 -14076
rect -6367 -14110 -6328 -14076
rect -5898 -14110 -5859 -14076
rect -5825 -14110 -5801 -14076
rect -5757 -14110 -5729 -14076
rect -5689 -14110 -5657 -14076
rect -5621 -14110 -5587 -14076
rect -5551 -14110 -5519 -14076
rect -5479 -14110 -5451 -14076
rect -5407 -14110 -5383 -14076
rect -5349 -14110 -5310 -14076
rect -4880 -14110 -4841 -14076
rect -4807 -14110 -4783 -14076
rect -4739 -14110 -4711 -14076
rect -4671 -14110 -4639 -14076
rect -4603 -14110 -4569 -14076
rect -4533 -14110 -4501 -14076
rect -4461 -14110 -4433 -14076
rect -4389 -14110 -4365 -14076
rect -4331 -14110 -4292 -14076
rect -3862 -14110 -3823 -14076
rect -3789 -14110 -3765 -14076
rect -3721 -14110 -3693 -14076
rect -3653 -14110 -3621 -14076
rect -3585 -14110 -3551 -14076
rect -3515 -14110 -3483 -14076
rect -3443 -14110 -3415 -14076
rect -3371 -14110 -3347 -14076
rect -3313 -14110 -3274 -14076
rect -2844 -14110 -2805 -14076
rect -2771 -14110 -2747 -14076
rect -2703 -14110 -2675 -14076
rect -2635 -14110 -2603 -14076
rect -2567 -14110 -2533 -14076
rect -2497 -14110 -2465 -14076
rect -2425 -14110 -2397 -14076
rect -2353 -14110 -2329 -14076
rect -2295 -14110 -2256 -14076
rect -1826 -14110 -1787 -14076
rect -1753 -14110 -1729 -14076
rect -1685 -14110 -1657 -14076
rect -1617 -14110 -1585 -14076
rect -1549 -14110 -1515 -14076
rect -1479 -14110 -1447 -14076
rect -1407 -14110 -1379 -14076
rect -1335 -14110 -1311 -14076
rect -1277 -14110 -1238 -14076
rect -808 -14110 -769 -14076
rect -735 -14110 -711 -14076
rect -667 -14110 -639 -14076
rect -599 -14110 -567 -14076
rect -531 -14110 -497 -14076
rect -461 -14110 -429 -14076
rect -389 -14110 -361 -14076
rect -317 -14110 -293 -14076
rect -259 -14110 -220 -14076
rect 24822 -14083 24922 -14069
rect -12322 -14151 -12222 -14141
rect -12322 -14213 -12289 -14151
rect -12255 -14213 -12222 -14151
rect -12322 -14219 -12222 -14213
rect -12322 -14285 -12289 -14219
rect -12255 -14285 -12222 -14219
rect -12322 -14287 -12222 -14285
rect -12322 -14321 -12289 -14287
rect -12255 -14321 -12222 -14287
rect -12322 -14323 -12222 -14321
rect -12322 -14389 -12289 -14323
rect -12255 -14389 -12222 -14323
rect -12322 -14395 -12222 -14389
rect -12322 -14457 -12289 -14395
rect -12255 -14457 -12222 -14395
rect -12322 -14467 -12222 -14457
rect -12322 -14525 -12289 -14467
rect -12255 -14525 -12222 -14467
rect -12322 -14539 -12222 -14525
rect -12322 -14593 -12289 -14539
rect -12255 -14593 -12222 -14539
rect -12322 -14611 -12222 -14593
rect -12322 -14661 -12289 -14611
rect -12255 -14661 -12222 -14611
rect -12322 -14683 -12222 -14661
rect -12322 -14729 -12289 -14683
rect -12255 -14729 -12222 -14683
rect -12322 -14755 -12222 -14729
rect -9184 -14179 -9150 -14144
rect -9184 -14251 -9150 -14227
rect -9184 -14323 -9150 -14295
rect -9184 -14395 -9150 -14363
rect -9184 -14465 -9150 -14431
rect -9184 -14533 -9150 -14501
rect -9184 -14601 -9150 -14573
rect -9184 -14669 -9150 -14645
rect -9184 -14752 -9150 -14717
rect -8166 -14179 -8132 -14144
rect -8166 -14251 -8132 -14227
rect -8166 -14323 -8132 -14295
rect -8166 -14395 -8132 -14363
rect -8166 -14465 -8132 -14431
rect -8166 -14533 -8132 -14501
rect -8166 -14601 -8132 -14573
rect -8166 -14669 -8132 -14645
rect -8166 -14752 -8132 -14717
rect -7148 -14179 -7114 -14144
rect -7148 -14251 -7114 -14227
rect -7148 -14323 -7114 -14295
rect -7148 -14395 -7114 -14363
rect -7148 -14465 -7114 -14431
rect -7148 -14533 -7114 -14501
rect -7148 -14601 -7114 -14573
rect -7148 -14669 -7114 -14645
rect -7148 -14752 -7114 -14717
rect -6130 -14179 -6096 -14144
rect -6130 -14251 -6096 -14227
rect -6130 -14323 -6096 -14295
rect -6130 -14395 -6096 -14363
rect -6130 -14465 -6096 -14431
rect -6130 -14533 -6096 -14501
rect -6130 -14601 -6096 -14573
rect -6130 -14669 -6096 -14645
rect -6130 -14752 -6096 -14717
rect -5112 -14179 -5078 -14144
rect -5112 -14251 -5078 -14227
rect -5112 -14323 -5078 -14295
rect -5112 -14395 -5078 -14363
rect -5112 -14465 -5078 -14431
rect -5112 -14533 -5078 -14501
rect -5112 -14601 -5078 -14573
rect -5112 -14669 -5078 -14645
rect -5112 -14752 -5078 -14717
rect -4094 -14179 -4060 -14144
rect -4094 -14251 -4060 -14227
rect -4094 -14323 -4060 -14295
rect -4094 -14395 -4060 -14363
rect -4094 -14465 -4060 -14431
rect -4094 -14533 -4060 -14501
rect -4094 -14601 -4060 -14573
rect -4094 -14669 -4060 -14645
rect -4094 -14752 -4060 -14717
rect -3076 -14179 -3042 -14144
rect -3076 -14251 -3042 -14227
rect -3076 -14323 -3042 -14295
rect -3076 -14395 -3042 -14363
rect -3076 -14465 -3042 -14431
rect -3076 -14533 -3042 -14501
rect -3076 -14601 -3042 -14573
rect -3076 -14669 -3042 -14645
rect -3076 -14752 -3042 -14717
rect -2058 -14179 -2024 -14144
rect -2058 -14251 -2024 -14227
rect -2058 -14323 -2024 -14295
rect -2058 -14395 -2024 -14363
rect -2058 -14465 -2024 -14431
rect -2058 -14533 -2024 -14501
rect -2058 -14601 -2024 -14573
rect -2058 -14669 -2024 -14645
rect -2058 -14752 -2024 -14717
rect -1040 -14179 -1006 -14144
rect -1040 -14251 -1006 -14227
rect -1040 -14323 -1006 -14295
rect -1040 -14395 -1006 -14363
rect -1040 -14465 -1006 -14431
rect -1040 -14533 -1006 -14501
rect -1040 -14601 -1006 -14573
rect -1040 -14669 -1006 -14645
rect -1040 -14752 -1006 -14717
rect -22 -14179 12 -14144
rect 2814 -14146 2853 -14112
rect 2887 -14146 2911 -14112
rect 2955 -14146 2983 -14112
rect 3023 -14146 3055 -14112
rect 3091 -14146 3125 -14112
rect 3161 -14146 3193 -14112
rect 3233 -14146 3261 -14112
rect 3305 -14146 3329 -14112
rect 3363 -14146 3402 -14112
rect 3832 -14146 3871 -14112
rect 3905 -14146 3929 -14112
rect 3973 -14146 4001 -14112
rect 4041 -14146 4073 -14112
rect 4109 -14146 4143 -14112
rect 4179 -14146 4211 -14112
rect 4251 -14146 4279 -14112
rect 4323 -14146 4347 -14112
rect 4381 -14146 4420 -14112
rect 4850 -14146 4889 -14112
rect 4923 -14146 4947 -14112
rect 4991 -14146 5019 -14112
rect 5059 -14146 5091 -14112
rect 5127 -14146 5161 -14112
rect 5197 -14146 5229 -14112
rect 5269 -14146 5297 -14112
rect 5341 -14146 5365 -14112
rect 5399 -14146 5438 -14112
rect 5868 -14146 5907 -14112
rect 5941 -14146 5965 -14112
rect 6009 -14146 6037 -14112
rect 6077 -14146 6109 -14112
rect 6145 -14146 6179 -14112
rect 6215 -14146 6247 -14112
rect 6287 -14146 6315 -14112
rect 6359 -14146 6383 -14112
rect 6417 -14146 6456 -14112
rect 6886 -14146 6925 -14112
rect 6959 -14146 6983 -14112
rect 7027 -14146 7055 -14112
rect 7095 -14146 7127 -14112
rect 7163 -14146 7197 -14112
rect 7233 -14146 7265 -14112
rect 7305 -14146 7333 -14112
rect 7377 -14146 7401 -14112
rect 7435 -14146 7474 -14112
rect 7904 -14146 7943 -14112
rect 7977 -14146 8001 -14112
rect 8045 -14146 8073 -14112
rect 8113 -14146 8145 -14112
rect 8181 -14146 8215 -14112
rect 8251 -14146 8283 -14112
rect 8323 -14146 8351 -14112
rect 8395 -14146 8419 -14112
rect 8453 -14146 8492 -14112
rect 8922 -14146 8961 -14112
rect 8995 -14146 9019 -14112
rect 9063 -14146 9091 -14112
rect 9131 -14146 9163 -14112
rect 9199 -14146 9233 -14112
rect 9269 -14146 9301 -14112
rect 9341 -14146 9369 -14112
rect 9413 -14146 9437 -14112
rect 9471 -14146 9510 -14112
rect 9940 -14146 9979 -14112
rect 10013 -14146 10037 -14112
rect 10081 -14146 10109 -14112
rect 10149 -14146 10181 -14112
rect 10217 -14146 10251 -14112
rect 10287 -14146 10319 -14112
rect 10359 -14146 10387 -14112
rect 10431 -14146 10455 -14112
rect 10489 -14146 10528 -14112
rect 10958 -14146 10997 -14112
rect 11031 -14146 11055 -14112
rect 11099 -14146 11127 -14112
rect 11167 -14146 11199 -14112
rect 11235 -14146 11269 -14112
rect 11305 -14146 11337 -14112
rect 11377 -14146 11405 -14112
rect 11449 -14146 11473 -14112
rect 11507 -14146 11546 -14112
rect 11976 -14146 12015 -14112
rect 12049 -14146 12073 -14112
rect 12117 -14146 12145 -14112
rect 12185 -14146 12217 -14112
rect 12253 -14146 12287 -14112
rect 12323 -14146 12355 -14112
rect 12395 -14146 12423 -14112
rect 12467 -14146 12491 -14112
rect 12525 -14146 12564 -14112
rect 12994 -14146 13033 -14112
rect 13067 -14146 13091 -14112
rect 13135 -14146 13163 -14112
rect 13203 -14146 13235 -14112
rect 13271 -14146 13305 -14112
rect 13341 -14146 13373 -14112
rect 13413 -14146 13441 -14112
rect 13485 -14146 13509 -14112
rect 13543 -14146 13582 -14112
rect 14012 -14146 14051 -14112
rect 14085 -14146 14109 -14112
rect 14153 -14146 14181 -14112
rect 14221 -14146 14253 -14112
rect 14289 -14146 14323 -14112
rect 14359 -14146 14391 -14112
rect 14431 -14146 14459 -14112
rect 14503 -14146 14527 -14112
rect 14561 -14146 14600 -14112
rect 15030 -14146 15069 -14112
rect 15103 -14146 15127 -14112
rect 15171 -14146 15199 -14112
rect 15239 -14146 15271 -14112
rect 15307 -14146 15341 -14112
rect 15377 -14146 15409 -14112
rect 15449 -14146 15477 -14112
rect 15521 -14146 15545 -14112
rect 15579 -14146 15618 -14112
rect 16048 -14146 16087 -14112
rect 16121 -14146 16145 -14112
rect 16189 -14146 16217 -14112
rect 16257 -14146 16289 -14112
rect 16325 -14146 16359 -14112
rect 16395 -14146 16427 -14112
rect 16467 -14146 16495 -14112
rect 16539 -14146 16563 -14112
rect 16597 -14146 16636 -14112
rect 17066 -14146 17105 -14112
rect 17139 -14146 17163 -14112
rect 17207 -14146 17235 -14112
rect 17275 -14146 17307 -14112
rect 17343 -14146 17377 -14112
rect 17413 -14146 17445 -14112
rect 17485 -14146 17513 -14112
rect 17557 -14146 17581 -14112
rect 17615 -14146 17654 -14112
rect 18084 -14146 18123 -14112
rect 18157 -14146 18181 -14112
rect 18225 -14146 18253 -14112
rect 18293 -14146 18325 -14112
rect 18361 -14146 18395 -14112
rect 18431 -14146 18463 -14112
rect 18503 -14146 18531 -14112
rect 18575 -14146 18599 -14112
rect 18633 -14146 18672 -14112
rect 19102 -14146 19141 -14112
rect 19175 -14146 19199 -14112
rect 19243 -14146 19271 -14112
rect 19311 -14146 19343 -14112
rect 19379 -14146 19413 -14112
rect 19449 -14146 19481 -14112
rect 19521 -14146 19549 -14112
rect 19593 -14146 19617 -14112
rect 19651 -14146 19690 -14112
rect 20120 -14146 20159 -14112
rect 20193 -14146 20217 -14112
rect 20261 -14146 20289 -14112
rect 20329 -14146 20361 -14112
rect 20397 -14146 20431 -14112
rect 20467 -14146 20499 -14112
rect 20539 -14146 20567 -14112
rect 20611 -14146 20635 -14112
rect 20669 -14146 20708 -14112
rect 21138 -14146 21177 -14112
rect 21211 -14146 21235 -14112
rect 21279 -14146 21307 -14112
rect 21347 -14146 21379 -14112
rect 21415 -14146 21449 -14112
rect 21485 -14146 21517 -14112
rect 21557 -14146 21585 -14112
rect 21629 -14146 21653 -14112
rect 21687 -14146 21726 -14112
rect 22156 -14146 22195 -14112
rect 22229 -14146 22253 -14112
rect 22297 -14146 22325 -14112
rect 22365 -14146 22397 -14112
rect 22433 -14146 22467 -14112
rect 22503 -14146 22535 -14112
rect 22575 -14146 22603 -14112
rect 22647 -14146 22671 -14112
rect 22705 -14146 22744 -14112
rect 24822 -14141 24855 -14083
rect 24889 -14141 24922 -14083
rect 4100 -14150 4160 -14146
rect 5116 -14150 5176 -14146
rect 9192 -14154 9252 -14146
rect 13258 -14150 13318 -14146
rect 15292 -14150 15352 -14146
rect 21404 -14150 21464 -14146
rect 24822 -14151 24922 -14141
rect -22 -14251 12 -14227
rect -22 -14323 12 -14295
rect -22 -14395 12 -14363
rect -22 -14465 12 -14431
rect -22 -14533 12 -14501
rect -22 -14601 12 -14573
rect -22 -14669 12 -14645
rect -22 -14752 12 -14717
rect 2582 -14215 2616 -14180
rect 2582 -14287 2616 -14263
rect 2582 -14359 2616 -14331
rect 2582 -14431 2616 -14399
rect 2582 -14501 2616 -14467
rect 2582 -14569 2616 -14537
rect 2582 -14637 2616 -14609
rect 2582 -14705 2616 -14681
rect -12322 -14797 -12289 -14755
rect -12255 -14797 -12222 -14755
rect -7656 -14786 -7596 -14784
rect -6642 -14786 -6582 -14784
rect -2568 -14786 -2508 -14784
rect -1552 -14786 -1492 -14784
rect -12322 -14827 -12222 -14797
rect -8952 -14820 -8913 -14786
rect -8879 -14820 -8855 -14786
rect -8811 -14820 -8783 -14786
rect -8743 -14820 -8711 -14786
rect -8675 -14820 -8641 -14786
rect -8605 -14820 -8573 -14786
rect -8533 -14820 -8505 -14786
rect -8461 -14820 -8437 -14786
rect -8403 -14820 -8364 -14786
rect -7934 -14820 -7895 -14786
rect -7861 -14820 -7837 -14786
rect -7793 -14820 -7765 -14786
rect -7725 -14820 -7693 -14786
rect -7657 -14820 -7623 -14786
rect -7587 -14820 -7555 -14786
rect -7515 -14820 -7487 -14786
rect -7443 -14820 -7419 -14786
rect -7385 -14820 -7346 -14786
rect -6916 -14820 -6877 -14786
rect -6843 -14820 -6819 -14786
rect -6775 -14820 -6747 -14786
rect -6707 -14820 -6675 -14786
rect -6639 -14820 -6605 -14786
rect -6569 -14820 -6537 -14786
rect -6497 -14820 -6469 -14786
rect -6425 -14820 -6401 -14786
rect -6367 -14820 -6328 -14786
rect -5898 -14820 -5859 -14786
rect -5825 -14820 -5801 -14786
rect -5757 -14820 -5729 -14786
rect -5689 -14820 -5657 -14786
rect -5621 -14820 -5587 -14786
rect -5551 -14820 -5519 -14786
rect -5479 -14820 -5451 -14786
rect -5407 -14820 -5383 -14786
rect -5349 -14820 -5310 -14786
rect -4880 -14820 -4841 -14786
rect -4807 -14820 -4783 -14786
rect -4739 -14820 -4711 -14786
rect -4671 -14820 -4639 -14786
rect -4603 -14820 -4569 -14786
rect -4533 -14820 -4501 -14786
rect -4461 -14820 -4433 -14786
rect -4389 -14820 -4365 -14786
rect -4331 -14820 -4292 -14786
rect -3862 -14820 -3823 -14786
rect -3789 -14820 -3765 -14786
rect -3721 -14820 -3693 -14786
rect -3653 -14820 -3621 -14786
rect -3585 -14820 -3551 -14786
rect -3515 -14820 -3483 -14786
rect -3443 -14820 -3415 -14786
rect -3371 -14820 -3347 -14786
rect -3313 -14820 -3274 -14786
rect -2844 -14820 -2805 -14786
rect -2771 -14820 -2747 -14786
rect -2703 -14820 -2675 -14786
rect -2635 -14820 -2603 -14786
rect -2567 -14820 -2533 -14786
rect -2497 -14820 -2465 -14786
rect -2425 -14820 -2397 -14786
rect -2353 -14820 -2329 -14786
rect -2295 -14820 -2256 -14786
rect -1826 -14820 -1787 -14786
rect -1753 -14820 -1729 -14786
rect -1685 -14820 -1657 -14786
rect -1617 -14820 -1585 -14786
rect -1549 -14820 -1515 -14786
rect -1479 -14820 -1447 -14786
rect -1407 -14820 -1379 -14786
rect -1335 -14820 -1311 -14786
rect -1277 -14820 -1238 -14786
rect -808 -14820 -769 -14786
rect -735 -14820 -711 -14786
rect -667 -14820 -639 -14786
rect -599 -14820 -567 -14786
rect -531 -14820 -497 -14786
rect -461 -14820 -429 -14786
rect -389 -14820 -361 -14786
rect -317 -14820 -293 -14786
rect -259 -14820 -220 -14786
rect 2582 -14788 2616 -14753
rect 3600 -14215 3634 -14180
rect 3600 -14287 3634 -14263
rect 3600 -14359 3634 -14331
rect 3600 -14431 3634 -14399
rect 3600 -14501 3634 -14467
rect 3600 -14569 3634 -14537
rect 3600 -14637 3634 -14609
rect 3600 -14705 3634 -14681
rect 3600 -14788 3634 -14753
rect 4618 -14215 4652 -14180
rect 4618 -14287 4652 -14263
rect 4618 -14359 4652 -14331
rect 4618 -14431 4652 -14399
rect 4618 -14501 4652 -14467
rect 4618 -14569 4652 -14537
rect 4618 -14637 4652 -14609
rect 4618 -14705 4652 -14681
rect 4618 -14788 4652 -14753
rect 5636 -14215 5670 -14180
rect 5636 -14287 5670 -14263
rect 5636 -14359 5670 -14331
rect 5636 -14431 5670 -14399
rect 5636 -14501 5670 -14467
rect 5636 -14569 5670 -14537
rect 5636 -14637 5670 -14609
rect 5636 -14705 5670 -14681
rect 5636 -14788 5670 -14753
rect 6654 -14215 6688 -14180
rect 6654 -14287 6688 -14263
rect 6654 -14359 6688 -14331
rect 6654 -14431 6688 -14399
rect 6654 -14501 6688 -14467
rect 6654 -14569 6688 -14537
rect 6654 -14637 6688 -14609
rect 6654 -14705 6688 -14681
rect 6654 -14788 6688 -14753
rect 7672 -14215 7706 -14180
rect 7672 -14287 7706 -14263
rect 7672 -14359 7706 -14331
rect 7672 -14431 7706 -14399
rect 7672 -14501 7706 -14467
rect 7672 -14569 7706 -14537
rect 7672 -14637 7706 -14609
rect 7672 -14705 7706 -14681
rect 7672 -14788 7706 -14753
rect 8690 -14215 8724 -14180
rect 8690 -14287 8724 -14263
rect 8690 -14359 8724 -14331
rect 8690 -14431 8724 -14399
rect 8690 -14501 8724 -14467
rect 8690 -14569 8724 -14537
rect 8690 -14637 8724 -14609
rect 8690 -14705 8724 -14681
rect 8690 -14788 8724 -14753
rect 9708 -14215 9742 -14180
rect 9708 -14287 9742 -14263
rect 9708 -14359 9742 -14331
rect 9708 -14431 9742 -14399
rect 9708 -14501 9742 -14467
rect 9708 -14569 9742 -14537
rect 9708 -14637 9742 -14609
rect 9708 -14705 9742 -14681
rect 9708 -14788 9742 -14753
rect 10726 -14215 10760 -14180
rect 10726 -14287 10760 -14263
rect 10726 -14359 10760 -14331
rect 10726 -14431 10760 -14399
rect 10726 -14501 10760 -14467
rect 10726 -14569 10760 -14537
rect 10726 -14637 10760 -14609
rect 10726 -14705 10760 -14681
rect 10726 -14788 10760 -14753
rect 11744 -14215 11778 -14180
rect 11744 -14287 11778 -14263
rect 11744 -14359 11778 -14331
rect 11744 -14431 11778 -14399
rect 11744 -14501 11778 -14467
rect 11744 -14569 11778 -14537
rect 11744 -14637 11778 -14609
rect 11744 -14705 11778 -14681
rect 11744 -14788 11778 -14753
rect 12762 -14215 12796 -14180
rect 12762 -14287 12796 -14263
rect 12762 -14359 12796 -14331
rect 12762 -14431 12796 -14399
rect 12762 -14501 12796 -14467
rect 12762 -14569 12796 -14537
rect 12762 -14637 12796 -14609
rect 12762 -14705 12796 -14681
rect 12762 -14788 12796 -14753
rect 13780 -14215 13814 -14180
rect 13780 -14287 13814 -14263
rect 13780 -14359 13814 -14331
rect 13780 -14431 13814 -14399
rect 13780 -14501 13814 -14467
rect 13780 -14569 13814 -14537
rect 13780 -14637 13814 -14609
rect 13780 -14705 13814 -14681
rect 13780 -14788 13814 -14753
rect 14798 -14215 14832 -14180
rect 14798 -14287 14832 -14263
rect 14798 -14359 14832 -14331
rect 14798 -14431 14832 -14399
rect 14798 -14501 14832 -14467
rect 14798 -14569 14832 -14537
rect 14798 -14637 14832 -14609
rect 14798 -14705 14832 -14681
rect 14798 -14788 14832 -14753
rect 15816 -14215 15850 -14180
rect 15816 -14287 15850 -14263
rect 15816 -14359 15850 -14331
rect 15816 -14431 15850 -14399
rect 15816 -14501 15850 -14467
rect 15816 -14569 15850 -14537
rect 15816 -14637 15850 -14609
rect 15816 -14705 15850 -14681
rect 15816 -14788 15850 -14753
rect 16834 -14215 16868 -14180
rect 16834 -14287 16868 -14263
rect 16834 -14359 16868 -14331
rect 16834 -14431 16868 -14399
rect 16834 -14501 16868 -14467
rect 16834 -14569 16868 -14537
rect 16834 -14637 16868 -14609
rect 16834 -14705 16868 -14681
rect 16834 -14788 16868 -14753
rect 17852 -14215 17886 -14180
rect 17852 -14287 17886 -14263
rect 17852 -14359 17886 -14331
rect 17852 -14431 17886 -14399
rect 17852 -14501 17886 -14467
rect 17852 -14569 17886 -14537
rect 17852 -14637 17886 -14609
rect 17852 -14705 17886 -14681
rect 17852 -14788 17886 -14753
rect 18870 -14215 18904 -14180
rect 18870 -14287 18904 -14263
rect 18870 -14359 18904 -14331
rect 18870 -14431 18904 -14399
rect 18870 -14501 18904 -14467
rect 18870 -14569 18904 -14537
rect 18870 -14637 18904 -14609
rect 18870 -14705 18904 -14681
rect 18870 -14788 18904 -14753
rect 19888 -14215 19922 -14180
rect 19888 -14287 19922 -14263
rect 19888 -14359 19922 -14331
rect 19888 -14431 19922 -14399
rect 19888 -14501 19922 -14467
rect 19888 -14569 19922 -14537
rect 19888 -14637 19922 -14609
rect 19888 -14705 19922 -14681
rect 19888 -14788 19922 -14753
rect 20906 -14215 20940 -14180
rect 20906 -14287 20940 -14263
rect 20906 -14359 20940 -14331
rect 20906 -14431 20940 -14399
rect 20906 -14501 20940 -14467
rect 20906 -14569 20940 -14537
rect 20906 -14637 20940 -14609
rect 20906 -14705 20940 -14681
rect 20906 -14788 20940 -14753
rect 21924 -14215 21958 -14180
rect 21924 -14287 21958 -14263
rect 21924 -14359 21958 -14331
rect 21924 -14431 21958 -14399
rect 21924 -14501 21958 -14467
rect 21924 -14569 21958 -14537
rect 21924 -14637 21958 -14609
rect 21924 -14705 21958 -14681
rect 21924 -14788 21958 -14753
rect 22942 -14215 22976 -14180
rect 22942 -14287 22976 -14263
rect 22942 -14359 22976 -14331
rect 22942 -14431 22976 -14399
rect 22942 -14501 22976 -14467
rect 22942 -14569 22976 -14537
rect 22942 -14637 22976 -14609
rect 22942 -14705 22976 -14681
rect 22942 -14788 22976 -14753
rect 24822 -14213 24855 -14151
rect 24889 -14213 24922 -14151
rect 24822 -14219 24922 -14213
rect 24822 -14285 24855 -14219
rect 24889 -14285 24922 -14219
rect 24822 -14287 24922 -14285
rect 24822 -14321 24855 -14287
rect 24889 -14321 24922 -14287
rect 24822 -14323 24922 -14321
rect 24822 -14389 24855 -14323
rect 24889 -14389 24922 -14323
rect 24822 -14395 24922 -14389
rect 24822 -14457 24855 -14395
rect 24889 -14457 24922 -14395
rect 24822 -14467 24922 -14457
rect 24822 -14525 24855 -14467
rect 24889 -14525 24922 -14467
rect 24822 -14539 24922 -14525
rect 24822 -14593 24855 -14539
rect 24889 -14593 24922 -14539
rect 24822 -14611 24922 -14593
rect 24822 -14661 24855 -14611
rect 24889 -14661 24922 -14611
rect 24822 -14683 24922 -14661
rect 24822 -14729 24855 -14683
rect 24889 -14729 24922 -14683
rect 24822 -14755 24922 -14729
rect 24822 -14797 24855 -14755
rect 24889 -14797 24922 -14755
rect 6126 -14822 6186 -14820
rect -12322 -14865 -12289 -14827
rect -12255 -14865 -12222 -14827
rect 2814 -14856 2853 -14822
rect 2887 -14856 2911 -14822
rect 2955 -14856 2983 -14822
rect 3023 -14856 3055 -14822
rect 3091 -14856 3125 -14822
rect 3161 -14856 3193 -14822
rect 3233 -14856 3261 -14822
rect 3305 -14856 3329 -14822
rect 3363 -14856 3402 -14822
rect 3832 -14856 3871 -14822
rect 3905 -14856 3929 -14822
rect 3973 -14856 4001 -14822
rect 4041 -14856 4073 -14822
rect 4109 -14856 4143 -14822
rect 4179 -14856 4211 -14822
rect 4251 -14856 4279 -14822
rect 4323 -14856 4347 -14822
rect 4381 -14856 4420 -14822
rect 4850 -14856 4889 -14822
rect 4923 -14856 4947 -14822
rect 4991 -14856 5019 -14822
rect 5059 -14856 5091 -14822
rect 5127 -14856 5161 -14822
rect 5197 -14856 5229 -14822
rect 5269 -14856 5297 -14822
rect 5341 -14856 5365 -14822
rect 5399 -14856 5438 -14822
rect 5868 -14856 5907 -14822
rect 5941 -14856 5965 -14822
rect 6009 -14856 6037 -14822
rect 6077 -14856 6109 -14822
rect 6145 -14856 6179 -14822
rect 6215 -14856 6247 -14822
rect 6287 -14856 6315 -14822
rect 6359 -14856 6383 -14822
rect 6417 -14856 6456 -14822
rect 6886 -14856 6925 -14822
rect 6959 -14856 6983 -14822
rect 7027 -14856 7055 -14822
rect 7095 -14856 7127 -14822
rect 7163 -14856 7197 -14822
rect 7233 -14856 7265 -14822
rect 7305 -14856 7333 -14822
rect 7377 -14856 7401 -14822
rect 7435 -14856 7474 -14822
rect 7904 -14856 7943 -14822
rect 7977 -14856 8001 -14822
rect 8045 -14856 8073 -14822
rect 8113 -14856 8145 -14822
rect 8181 -14856 8215 -14822
rect 8251 -14856 8283 -14822
rect 8323 -14856 8351 -14822
rect 8395 -14856 8419 -14822
rect 8453 -14856 8492 -14822
rect 8922 -14856 8961 -14822
rect 8995 -14856 9019 -14822
rect 9063 -14856 9091 -14822
rect 9131 -14856 9163 -14822
rect 9199 -14856 9233 -14822
rect 9269 -14856 9301 -14822
rect 9341 -14856 9369 -14822
rect 9413 -14856 9437 -14822
rect 9471 -14856 9510 -14822
rect 9940 -14856 9979 -14822
rect 10013 -14856 10037 -14822
rect 10081 -14856 10109 -14822
rect 10149 -14856 10181 -14822
rect 10217 -14856 10251 -14822
rect 10287 -14856 10319 -14822
rect 10359 -14856 10387 -14822
rect 10431 -14856 10455 -14822
rect 10489 -14856 10528 -14822
rect 10958 -14856 10997 -14822
rect 11031 -14856 11055 -14822
rect 11099 -14856 11127 -14822
rect 11167 -14856 11199 -14822
rect 11235 -14856 11269 -14822
rect 11305 -14856 11337 -14822
rect 11377 -14856 11405 -14822
rect 11449 -14856 11473 -14822
rect 11507 -14856 11546 -14822
rect 11976 -14856 12015 -14822
rect 12049 -14856 12073 -14822
rect 12117 -14856 12145 -14822
rect 12185 -14856 12217 -14822
rect 12253 -14856 12287 -14822
rect 12323 -14856 12355 -14822
rect 12395 -14856 12423 -14822
rect 12467 -14856 12491 -14822
rect 12525 -14856 12564 -14822
rect 12994 -14856 13033 -14822
rect 13067 -14856 13091 -14822
rect 13135 -14856 13163 -14822
rect 13203 -14856 13235 -14822
rect 13271 -14856 13305 -14822
rect 13341 -14856 13373 -14822
rect 13413 -14856 13441 -14822
rect 13485 -14856 13509 -14822
rect 13543 -14856 13582 -14822
rect 14012 -14856 14051 -14822
rect 14085 -14856 14109 -14822
rect 14153 -14856 14181 -14822
rect 14221 -14856 14253 -14822
rect 14289 -14856 14323 -14822
rect 14359 -14856 14391 -14822
rect 14431 -14856 14459 -14822
rect 14503 -14856 14527 -14822
rect 14561 -14856 14600 -14822
rect 15030 -14856 15069 -14822
rect 15103 -14856 15127 -14822
rect 15171 -14856 15199 -14822
rect 15239 -14856 15271 -14822
rect 15307 -14856 15341 -14822
rect 15377 -14856 15409 -14822
rect 15449 -14856 15477 -14822
rect 15521 -14856 15545 -14822
rect 15579 -14856 15618 -14822
rect 16048 -14856 16087 -14822
rect 16121 -14856 16145 -14822
rect 16189 -14856 16217 -14822
rect 16257 -14856 16289 -14822
rect 16325 -14856 16359 -14822
rect 16395 -14856 16427 -14822
rect 16467 -14856 16495 -14822
rect 16539 -14856 16563 -14822
rect 16597 -14856 16636 -14822
rect 17066 -14856 17105 -14822
rect 17139 -14856 17163 -14822
rect 17207 -14856 17235 -14822
rect 17275 -14856 17309 -14822
rect 17343 -14856 17377 -14822
rect 17413 -14856 17445 -14822
rect 17485 -14856 17513 -14822
rect 17557 -14856 17581 -14822
rect 17615 -14856 17654 -14822
rect 18084 -14856 18123 -14822
rect 18157 -14856 18181 -14822
rect 18225 -14856 18253 -14822
rect 18293 -14856 18327 -14822
rect 18361 -14856 18395 -14822
rect 18429 -14856 18463 -14822
rect 18503 -14856 18531 -14822
rect 18575 -14856 18599 -14822
rect 18633 -14856 18672 -14822
rect 19102 -14856 19141 -14822
rect 19175 -14856 19199 -14822
rect 19243 -14856 19271 -14822
rect 19311 -14856 19343 -14822
rect 19379 -14856 19413 -14822
rect 19449 -14856 19481 -14822
rect 19521 -14856 19549 -14822
rect 19593 -14856 19617 -14822
rect 19651 -14856 19690 -14822
rect 20120 -14856 20159 -14822
rect 20193 -14856 20217 -14822
rect 20261 -14856 20289 -14822
rect 20329 -14856 20361 -14822
rect 20397 -14856 20431 -14822
rect 20467 -14856 20499 -14822
rect 20539 -14856 20567 -14822
rect 20611 -14856 20635 -14822
rect 20669 -14856 20708 -14822
rect 21138 -14856 21177 -14822
rect 21211 -14856 21235 -14822
rect 21279 -14856 21307 -14822
rect 21347 -14856 21379 -14822
rect 21415 -14856 21449 -14822
rect 21485 -14856 21517 -14822
rect 21557 -14856 21585 -14822
rect 21629 -14856 21653 -14822
rect 21687 -14856 21726 -14822
rect 22156 -14856 22195 -14822
rect 22229 -14856 22253 -14822
rect 22297 -14856 22325 -14822
rect 22365 -14856 22397 -14822
rect 22433 -14856 22467 -14822
rect 22503 -14856 22535 -14822
rect 22575 -14856 22603 -14822
rect 22647 -14856 22671 -14822
rect 22705 -14856 22744 -14822
rect 24822 -14827 24922 -14797
rect 8160 -14860 8220 -14856
rect -12322 -14899 -12222 -14865
rect 17318 -14870 17378 -14856
rect 18352 -14870 18412 -14856
rect 24822 -14865 24855 -14827
rect 24889 -14865 24922 -14827
rect -12322 -14933 -12289 -14899
rect -12255 -14933 -12222 -14899
rect -8952 -14928 -8913 -14894
rect -8879 -14928 -8855 -14894
rect -8811 -14928 -8783 -14894
rect -8743 -14928 -8711 -14894
rect -8675 -14928 -8641 -14894
rect -8605 -14928 -8573 -14894
rect -8533 -14928 -8505 -14894
rect -8461 -14928 -8437 -14894
rect -8403 -14928 -8364 -14894
rect -7934 -14928 -7895 -14894
rect -7861 -14928 -7837 -14894
rect -7793 -14928 -7765 -14894
rect -7725 -14928 -7693 -14894
rect -7657 -14928 -7623 -14894
rect -7587 -14928 -7555 -14894
rect -7515 -14928 -7487 -14894
rect -7443 -14928 -7419 -14894
rect -7385 -14928 -7346 -14894
rect -6916 -14928 -6877 -14894
rect -6843 -14928 -6819 -14894
rect -6775 -14928 -6747 -14894
rect -6707 -14928 -6675 -14894
rect -6639 -14928 -6605 -14894
rect -6569 -14928 -6537 -14894
rect -6497 -14928 -6469 -14894
rect -6425 -14928 -6401 -14894
rect -6367 -14928 -6328 -14894
rect -5898 -14928 -5859 -14894
rect -5825 -14928 -5801 -14894
rect -5757 -14928 -5729 -14894
rect -5689 -14928 -5657 -14894
rect -5621 -14928 -5587 -14894
rect -5551 -14928 -5519 -14894
rect -5479 -14928 -5451 -14894
rect -5407 -14928 -5383 -14894
rect -5349 -14928 -5310 -14894
rect -4880 -14928 -4841 -14894
rect -4807 -14928 -4783 -14894
rect -4739 -14928 -4711 -14894
rect -4671 -14928 -4639 -14894
rect -4603 -14928 -4569 -14894
rect -4533 -14928 -4501 -14894
rect -4461 -14928 -4433 -14894
rect -4389 -14928 -4365 -14894
rect -4331 -14928 -4292 -14894
rect -3862 -14928 -3823 -14894
rect -3789 -14928 -3765 -14894
rect -3721 -14928 -3693 -14894
rect -3653 -14928 -3621 -14894
rect -3585 -14928 -3551 -14894
rect -3515 -14928 -3483 -14894
rect -3443 -14928 -3415 -14894
rect -3371 -14928 -3347 -14894
rect -3313 -14928 -3274 -14894
rect -2844 -14928 -2805 -14894
rect -2771 -14928 -2747 -14894
rect -2703 -14928 -2675 -14894
rect -2635 -14928 -2603 -14894
rect -2567 -14928 -2533 -14894
rect -2497 -14928 -2465 -14894
rect -2425 -14928 -2397 -14894
rect -2353 -14928 -2329 -14894
rect -2295 -14928 -2256 -14894
rect -1826 -14928 -1787 -14894
rect -1753 -14928 -1729 -14894
rect -1685 -14928 -1657 -14894
rect -1617 -14928 -1585 -14894
rect -1549 -14928 -1515 -14894
rect -1479 -14928 -1447 -14894
rect -1407 -14928 -1379 -14894
rect -1335 -14928 -1311 -14894
rect -1277 -14928 -1238 -14894
rect -808 -14928 -769 -14894
rect -735 -14928 -711 -14894
rect -667 -14928 -639 -14894
rect -599 -14928 -567 -14894
rect -531 -14928 -497 -14894
rect -461 -14928 -429 -14894
rect -389 -14928 -361 -14894
rect -317 -14928 -293 -14894
rect -259 -14928 -220 -14894
rect 24822 -14899 24922 -14865
rect -12322 -14967 -12222 -14933
rect 24822 -14933 24855 -14899
rect 24889 -14933 24922 -14899
rect -12322 -15005 -12289 -14967
rect -12255 -15005 -12222 -14967
rect -12322 -15035 -12222 -15005
rect -12322 -15077 -12289 -15035
rect -12255 -15077 -12222 -15035
rect -12322 -15103 -12222 -15077
rect -12322 -15149 -12289 -15103
rect -12255 -15149 -12222 -15103
rect -12322 -15171 -12222 -15149
rect -12322 -15221 -12289 -15171
rect -12255 -15221 -12222 -15171
rect -12322 -15239 -12222 -15221
rect -12322 -15293 -12289 -15239
rect -12255 -15293 -12222 -15239
rect -12322 -15307 -12222 -15293
rect -12322 -15365 -12289 -15307
rect -12255 -15365 -12222 -15307
rect -12322 -15375 -12222 -15365
rect -12322 -15437 -12289 -15375
rect -12255 -15437 -12222 -15375
rect -12322 -15443 -12222 -15437
rect -12322 -15509 -12289 -15443
rect -12255 -15509 -12222 -15443
rect -12322 -15511 -12222 -15509
rect -12322 -15545 -12289 -15511
rect -12255 -15545 -12222 -15511
rect -12322 -15547 -12222 -15545
rect -12322 -15613 -12289 -15547
rect -12255 -15613 -12222 -15547
rect -9184 -14997 -9150 -14962
rect -9184 -15069 -9150 -15045
rect -9184 -15141 -9150 -15113
rect -9184 -15213 -9150 -15181
rect -9184 -15283 -9150 -15249
rect -9184 -15351 -9150 -15319
rect -9184 -15419 -9150 -15391
rect -9184 -15487 -9150 -15463
rect -9184 -15570 -9150 -15535
rect -8166 -14997 -8132 -14962
rect -8166 -15069 -8132 -15045
rect -8166 -15141 -8132 -15113
rect -8166 -15213 -8132 -15181
rect -8166 -15283 -8132 -15249
rect -8166 -15351 -8132 -15319
rect -8166 -15419 -8132 -15391
rect -8166 -15487 -8132 -15463
rect -8166 -15570 -8132 -15535
rect -7148 -14997 -7114 -14962
rect -7148 -15069 -7114 -15045
rect -7148 -15141 -7114 -15113
rect -7148 -15213 -7114 -15181
rect -7148 -15283 -7114 -15249
rect -7148 -15351 -7114 -15319
rect -7148 -15419 -7114 -15391
rect -7148 -15487 -7114 -15463
rect -7148 -15570 -7114 -15535
rect -6130 -14997 -6096 -14962
rect -6130 -15069 -6096 -15045
rect -6130 -15141 -6096 -15113
rect -6130 -15213 -6096 -15181
rect -6130 -15283 -6096 -15249
rect -6130 -15351 -6096 -15319
rect -6130 -15419 -6096 -15391
rect -6130 -15487 -6096 -15463
rect -6130 -15570 -6096 -15535
rect -5112 -14997 -5078 -14962
rect -5112 -15069 -5078 -15045
rect -5112 -15141 -5078 -15113
rect -5112 -15213 -5078 -15181
rect -5112 -15283 -5078 -15249
rect -5112 -15351 -5078 -15319
rect -5112 -15419 -5078 -15391
rect -5112 -15487 -5078 -15463
rect -5112 -15570 -5078 -15535
rect -4094 -14997 -4060 -14962
rect -4094 -15069 -4060 -15045
rect -4094 -15141 -4060 -15113
rect -4094 -15213 -4060 -15181
rect -4094 -15283 -4060 -15249
rect -4094 -15351 -4060 -15319
rect -4094 -15419 -4060 -15391
rect -4094 -15487 -4060 -15463
rect -4094 -15570 -4060 -15535
rect -3076 -14997 -3042 -14962
rect -3076 -15069 -3042 -15045
rect -3076 -15141 -3042 -15113
rect -3076 -15213 -3042 -15181
rect -3076 -15283 -3042 -15249
rect -3076 -15351 -3042 -15319
rect -3076 -15419 -3042 -15391
rect -3076 -15487 -3042 -15463
rect -3076 -15570 -3042 -15535
rect -2058 -14997 -2024 -14962
rect -2058 -15069 -2024 -15045
rect -2058 -15141 -2024 -15113
rect -2058 -15213 -2024 -15181
rect -2058 -15283 -2024 -15249
rect -2058 -15351 -2024 -15319
rect -2058 -15419 -2024 -15391
rect -2058 -15487 -2024 -15463
rect -2058 -15570 -2024 -15535
rect -1040 -14997 -1006 -14962
rect -1040 -15069 -1006 -15045
rect -1040 -15141 -1006 -15113
rect -1040 -15213 -1006 -15181
rect -1040 -15283 -1006 -15249
rect -1040 -15351 -1006 -15319
rect -1040 -15419 -1006 -15391
rect -1040 -15487 -1006 -15463
rect -1040 -15570 -1006 -15535
rect -22 -14997 12 -14962
rect -22 -15069 12 -15045
rect -22 -15141 12 -15113
rect -22 -15213 12 -15181
rect -22 -15283 12 -15249
rect -22 -15351 12 -15319
rect 24822 -14967 24922 -14933
rect 24822 -15005 24855 -14967
rect 24889 -15005 24922 -14967
rect 24822 -15035 24922 -15005
rect 24822 -15077 24855 -15035
rect 24889 -15077 24922 -15035
rect 24822 -15103 24922 -15077
rect 24822 -15149 24855 -15103
rect 24889 -15149 24922 -15103
rect 24822 -15171 24922 -15149
rect 24822 -15221 24855 -15171
rect 24889 -15221 24922 -15171
rect 24822 -15239 24922 -15221
rect 24822 -15293 24855 -15239
rect 24889 -15293 24922 -15239
rect 24822 -15307 24922 -15293
rect 2812 -15380 2851 -15346
rect 2885 -15380 2909 -15346
rect 2953 -15380 2981 -15346
rect 3021 -15380 3053 -15346
rect 3089 -15380 3123 -15346
rect 3159 -15380 3191 -15346
rect 3231 -15380 3259 -15346
rect 3303 -15380 3327 -15346
rect 3361 -15380 3400 -15346
rect 3830 -15380 3869 -15346
rect 3903 -15380 3927 -15346
rect 3971 -15380 3999 -15346
rect 4039 -15380 4071 -15346
rect 4107 -15380 4141 -15346
rect 4177 -15380 4209 -15346
rect 4249 -15380 4277 -15346
rect 4321 -15380 4345 -15346
rect 4379 -15380 4418 -15346
rect 4848 -15380 4887 -15346
rect 4921 -15380 4945 -15346
rect 4989 -15380 5017 -15346
rect 5057 -15380 5089 -15346
rect 5125 -15380 5159 -15346
rect 5195 -15380 5227 -15346
rect 5267 -15380 5295 -15346
rect 5339 -15380 5363 -15346
rect 5397 -15380 5436 -15346
rect 5866 -15380 5905 -15346
rect 5939 -15380 5963 -15346
rect 6007 -15380 6035 -15346
rect 6075 -15380 6107 -15346
rect 6143 -15380 6177 -15346
rect 6213 -15380 6245 -15346
rect 6285 -15380 6313 -15346
rect 6357 -15380 6381 -15346
rect 6415 -15380 6454 -15346
rect 6884 -15380 6923 -15346
rect 6957 -15380 6981 -15346
rect 7025 -15380 7053 -15346
rect 7093 -15380 7125 -15346
rect 7161 -15380 7195 -15346
rect 7231 -15380 7263 -15346
rect 7303 -15380 7331 -15346
rect 7375 -15380 7399 -15346
rect 7433 -15380 7472 -15346
rect 7902 -15380 7941 -15346
rect 7975 -15380 7999 -15346
rect 8043 -15380 8071 -15346
rect 8111 -15380 8143 -15346
rect 8179 -15380 8213 -15346
rect 8249 -15380 8281 -15346
rect 8321 -15380 8349 -15346
rect 8393 -15380 8417 -15346
rect 8451 -15380 8490 -15346
rect 8920 -15380 8959 -15346
rect 8993 -15380 9017 -15346
rect 9061 -15380 9089 -15346
rect 9129 -15380 9161 -15346
rect 9197 -15380 9231 -15346
rect 9267 -15380 9299 -15346
rect 9339 -15380 9367 -15346
rect 9411 -15380 9435 -15346
rect 9469 -15380 9508 -15346
rect 9938 -15380 9977 -15346
rect 10011 -15380 10035 -15346
rect 10079 -15380 10107 -15346
rect 10147 -15380 10179 -15346
rect 10215 -15380 10249 -15346
rect 10285 -15380 10317 -15346
rect 10357 -15380 10385 -15346
rect 10429 -15380 10453 -15346
rect 10487 -15380 10526 -15346
rect 10956 -15380 10995 -15346
rect 11029 -15380 11053 -15346
rect 11097 -15380 11125 -15346
rect 11165 -15380 11197 -15346
rect 11233 -15380 11267 -15346
rect 11303 -15380 11335 -15346
rect 11375 -15380 11403 -15346
rect 11447 -15380 11471 -15346
rect 11505 -15380 11544 -15346
rect 11974 -15380 12013 -15346
rect 12047 -15380 12071 -15346
rect 12115 -15380 12143 -15346
rect 12183 -15380 12215 -15346
rect 12251 -15380 12285 -15346
rect 12321 -15380 12353 -15346
rect 12393 -15380 12421 -15346
rect 12465 -15380 12489 -15346
rect 12523 -15380 12562 -15346
rect 12992 -15380 13031 -15346
rect 13065 -15380 13089 -15346
rect 13133 -15380 13161 -15346
rect 13201 -15380 13233 -15346
rect 13269 -15380 13303 -15346
rect 13339 -15380 13371 -15346
rect 13411 -15380 13439 -15346
rect 13483 -15380 13507 -15346
rect 13541 -15380 13580 -15346
rect 14010 -15380 14049 -15346
rect 14083 -15380 14107 -15346
rect 14151 -15380 14179 -15346
rect 14219 -15380 14251 -15346
rect 14287 -15380 14321 -15346
rect 14357 -15380 14389 -15346
rect 14429 -15380 14457 -15346
rect 14501 -15380 14525 -15346
rect 14559 -15380 14598 -15346
rect 15028 -15380 15067 -15346
rect 15101 -15380 15125 -15346
rect 15169 -15380 15197 -15346
rect 15237 -15380 15269 -15346
rect 15305 -15380 15339 -15346
rect 15375 -15380 15407 -15346
rect 15447 -15380 15475 -15346
rect 15519 -15380 15543 -15346
rect 15577 -15380 15616 -15346
rect 16046 -15380 16085 -15346
rect 16119 -15380 16143 -15346
rect 16187 -15380 16215 -15346
rect 16255 -15380 16287 -15346
rect 16323 -15380 16357 -15346
rect 16393 -15380 16425 -15346
rect 16465 -15380 16493 -15346
rect 16537 -15380 16561 -15346
rect 16595 -15380 16634 -15346
rect 17064 -15380 17103 -15346
rect 17137 -15380 17161 -15346
rect 17205 -15380 17233 -15346
rect 17273 -15380 17305 -15346
rect 17341 -15380 17375 -15346
rect 17411 -15380 17443 -15346
rect 17483 -15380 17511 -15346
rect 17555 -15380 17579 -15346
rect 17613 -15380 17652 -15346
rect 18082 -15380 18121 -15346
rect 18155 -15380 18179 -15346
rect 18223 -15380 18251 -15346
rect 18291 -15380 18323 -15346
rect 18359 -15380 18393 -15346
rect 18429 -15380 18461 -15346
rect 18501 -15380 18529 -15346
rect 18573 -15380 18597 -15346
rect 18631 -15380 18670 -15346
rect 19100 -15380 19139 -15346
rect 19173 -15380 19197 -15346
rect 19241 -15380 19269 -15346
rect 19309 -15380 19341 -15346
rect 19377 -15380 19411 -15346
rect 19447 -15380 19479 -15346
rect 19519 -15380 19547 -15346
rect 19591 -15380 19615 -15346
rect 19649 -15380 19688 -15346
rect 20118 -15380 20157 -15346
rect 20191 -15380 20215 -15346
rect 20259 -15380 20287 -15346
rect 20327 -15380 20359 -15346
rect 20395 -15380 20429 -15346
rect 20465 -15380 20497 -15346
rect 20537 -15380 20565 -15346
rect 20609 -15380 20633 -15346
rect 20667 -15380 20706 -15346
rect 21136 -15380 21175 -15346
rect 21209 -15380 21233 -15346
rect 21277 -15380 21305 -15346
rect 21345 -15380 21377 -15346
rect 21413 -15380 21447 -15346
rect 21483 -15380 21515 -15346
rect 21555 -15380 21583 -15346
rect 21627 -15380 21651 -15346
rect 21685 -15380 21724 -15346
rect 22154 -15380 22193 -15346
rect 22227 -15380 22251 -15346
rect 22295 -15380 22323 -15346
rect 22363 -15380 22395 -15346
rect 22431 -15380 22465 -15346
rect 22501 -15380 22533 -15346
rect 22573 -15380 22601 -15346
rect 22645 -15380 22669 -15346
rect 22703 -15380 22742 -15346
rect 24822 -15365 24855 -15307
rect 24889 -15365 24922 -15307
rect 24822 -15375 24922 -15365
rect 5122 -15384 5182 -15380
rect -22 -15419 12 -15391
rect -22 -15487 12 -15463
rect -22 -15570 12 -15535
rect 2580 -15449 2614 -15414
rect 2580 -15521 2614 -15497
rect 2580 -15593 2614 -15565
rect -12322 -15619 -12222 -15613
rect -12322 -15681 -12289 -15619
rect -12255 -15681 -12222 -15619
rect -8952 -15638 -8913 -15604
rect -8879 -15638 -8855 -15604
rect -8811 -15638 -8783 -15604
rect -8743 -15638 -8711 -15604
rect -8675 -15638 -8641 -15604
rect -8605 -15638 -8573 -15604
rect -8533 -15638 -8505 -15604
rect -8461 -15638 -8437 -15604
rect -8403 -15638 -8364 -15604
rect -7934 -15638 -7895 -15604
rect -7861 -15638 -7837 -15604
rect -7793 -15638 -7765 -15604
rect -7725 -15638 -7693 -15604
rect -7657 -15638 -7623 -15604
rect -7587 -15638 -7555 -15604
rect -7515 -15638 -7487 -15604
rect -7443 -15638 -7419 -15604
rect -7385 -15638 -7346 -15604
rect -6916 -15638 -6877 -15604
rect -6843 -15638 -6819 -15604
rect -6775 -15638 -6747 -15604
rect -6707 -15638 -6675 -15604
rect -6639 -15638 -6605 -15604
rect -6569 -15638 -6537 -15604
rect -6497 -15638 -6469 -15604
rect -6425 -15638 -6401 -15604
rect -6367 -15638 -6328 -15604
rect -5898 -15638 -5859 -15604
rect -5825 -15638 -5801 -15604
rect -5757 -15638 -5729 -15604
rect -5689 -15638 -5657 -15604
rect -5621 -15638 -5587 -15604
rect -5551 -15638 -5519 -15604
rect -5479 -15638 -5451 -15604
rect -5407 -15638 -5383 -15604
rect -5349 -15638 -5310 -15604
rect -4880 -15638 -4841 -15604
rect -4807 -15638 -4783 -15604
rect -4739 -15638 -4711 -15604
rect -4671 -15638 -4639 -15604
rect -4603 -15638 -4569 -15604
rect -4533 -15638 -4501 -15604
rect -4461 -15638 -4433 -15604
rect -4389 -15638 -4365 -15604
rect -4331 -15638 -4292 -15604
rect -3862 -15638 -3823 -15604
rect -3789 -15638 -3765 -15604
rect -3721 -15638 -3693 -15604
rect -3653 -15638 -3621 -15604
rect -3585 -15638 -3551 -15604
rect -3515 -15638 -3483 -15604
rect -3443 -15638 -3415 -15604
rect -3371 -15638 -3347 -15604
rect -3313 -15638 -3274 -15604
rect -2844 -15638 -2805 -15604
rect -2771 -15638 -2747 -15604
rect -2703 -15638 -2675 -15604
rect -2635 -15638 -2603 -15604
rect -2567 -15638 -2533 -15604
rect -2497 -15638 -2465 -15604
rect -2425 -15638 -2397 -15604
rect -2353 -15638 -2329 -15604
rect -2295 -15638 -2256 -15604
rect -1826 -15638 -1787 -15604
rect -1753 -15638 -1729 -15604
rect -1685 -15638 -1657 -15604
rect -1617 -15638 -1585 -15604
rect -1549 -15638 -1515 -15604
rect -1479 -15638 -1447 -15604
rect -1407 -15638 -1379 -15604
rect -1335 -15638 -1311 -15604
rect -1277 -15638 -1238 -15604
rect -808 -15638 -769 -15604
rect -735 -15638 -711 -15604
rect -667 -15638 -639 -15604
rect -599 -15638 -567 -15604
rect -531 -15638 -497 -15604
rect -461 -15638 -429 -15604
rect -389 -15638 -361 -15604
rect -317 -15638 -293 -15604
rect -259 -15638 -220 -15604
rect -12322 -15691 -12222 -15681
rect -12322 -15749 -12289 -15691
rect -12255 -15749 -12222 -15691
rect 2580 -15665 2614 -15633
rect -8952 -15746 -8913 -15712
rect -8879 -15746 -8855 -15712
rect -8811 -15746 -8783 -15712
rect -8743 -15746 -8711 -15712
rect -8675 -15746 -8641 -15712
rect -8605 -15746 -8573 -15712
rect -8533 -15746 -8505 -15712
rect -8461 -15746 -8437 -15712
rect -8403 -15746 -8364 -15712
rect -7934 -15746 -7895 -15712
rect -7861 -15746 -7837 -15712
rect -7793 -15746 -7765 -15712
rect -7725 -15746 -7693 -15712
rect -7657 -15746 -7623 -15712
rect -7587 -15746 -7555 -15712
rect -7515 -15746 -7487 -15712
rect -7443 -15746 -7419 -15712
rect -7385 -15746 -7346 -15712
rect -6916 -15746 -6877 -15712
rect -6843 -15746 -6819 -15712
rect -6775 -15746 -6747 -15712
rect -6707 -15746 -6675 -15712
rect -6639 -15746 -6605 -15712
rect -6569 -15746 -6537 -15712
rect -6497 -15746 -6469 -15712
rect -6425 -15746 -6401 -15712
rect -6367 -15746 -6328 -15712
rect -5898 -15746 -5859 -15712
rect -5825 -15746 -5801 -15712
rect -5757 -15746 -5729 -15712
rect -5689 -15746 -5657 -15712
rect -5621 -15746 -5587 -15712
rect -5551 -15746 -5519 -15712
rect -5479 -15746 -5451 -15712
rect -5407 -15746 -5383 -15712
rect -5349 -15746 -5310 -15712
rect -4880 -15746 -4841 -15712
rect -4807 -15746 -4783 -15712
rect -4739 -15746 -4711 -15712
rect -4671 -15746 -4639 -15712
rect -4603 -15746 -4569 -15712
rect -4533 -15746 -4501 -15712
rect -4461 -15746 -4433 -15712
rect -4389 -15746 -4365 -15712
rect -4331 -15746 -4292 -15712
rect -3862 -15746 -3823 -15712
rect -3789 -15746 -3765 -15712
rect -3721 -15746 -3693 -15712
rect -3653 -15746 -3621 -15712
rect -3585 -15746 -3551 -15712
rect -3515 -15746 -3483 -15712
rect -3443 -15746 -3415 -15712
rect -3371 -15746 -3347 -15712
rect -3313 -15746 -3274 -15712
rect -2844 -15746 -2805 -15712
rect -2771 -15746 -2747 -15712
rect -2703 -15746 -2675 -15712
rect -2635 -15746 -2603 -15712
rect -2567 -15746 -2533 -15712
rect -2497 -15746 -2465 -15712
rect -2425 -15746 -2397 -15712
rect -2353 -15746 -2329 -15712
rect -2295 -15746 -2256 -15712
rect -1826 -15746 -1787 -15712
rect -1753 -15746 -1729 -15712
rect -1685 -15746 -1657 -15712
rect -1617 -15746 -1585 -15712
rect -1549 -15746 -1515 -15712
rect -1479 -15746 -1447 -15712
rect -1407 -15746 -1379 -15712
rect -1335 -15746 -1311 -15712
rect -1277 -15746 -1238 -15712
rect -808 -15746 -769 -15712
rect -735 -15746 -711 -15712
rect -667 -15746 -639 -15712
rect -599 -15746 -567 -15712
rect -531 -15746 -497 -15712
rect -461 -15746 -429 -15712
rect -389 -15746 -361 -15712
rect -317 -15746 -293 -15712
rect -259 -15746 -220 -15712
rect 2580 -15735 2614 -15701
rect -3596 -15748 -3536 -15746
rect -12322 -15763 -12222 -15749
rect -12322 -15817 -12289 -15763
rect -12255 -15817 -12222 -15763
rect -12322 -15835 -12222 -15817
rect -12322 -15885 -12289 -15835
rect -12255 -15885 -12222 -15835
rect -12322 -15907 -12222 -15885
rect -12322 -15953 -12289 -15907
rect -12255 -15953 -12222 -15907
rect -12322 -15979 -12222 -15953
rect -12322 -16021 -12289 -15979
rect -12255 -16021 -12222 -15979
rect -12322 -16051 -12222 -16021
rect -12322 -16089 -12289 -16051
rect -12255 -16089 -12222 -16051
rect -12322 -16123 -12222 -16089
rect -12322 -16157 -12289 -16123
rect -12255 -16157 -12222 -16123
rect -12322 -16191 -12222 -16157
rect -12322 -16229 -12289 -16191
rect -12255 -16229 -12222 -16191
rect -12322 -16259 -12222 -16229
rect -12322 -16301 -12289 -16259
rect -12255 -16301 -12222 -16259
rect -12322 -16327 -12222 -16301
rect -12322 -16373 -12289 -16327
rect -12255 -16373 -12222 -16327
rect -12322 -16395 -12222 -16373
rect -9184 -15815 -9150 -15780
rect -9184 -15887 -9150 -15863
rect -9184 -15959 -9150 -15931
rect -9184 -16031 -9150 -15999
rect -9184 -16101 -9150 -16067
rect -9184 -16169 -9150 -16137
rect -9184 -16237 -9150 -16209
rect -9184 -16305 -9150 -16281
rect -9184 -16388 -9150 -16353
rect -8166 -15815 -8132 -15780
rect -8166 -15887 -8132 -15863
rect -8166 -15959 -8132 -15931
rect -8166 -16031 -8132 -15999
rect -8166 -16101 -8132 -16067
rect -8166 -16169 -8132 -16137
rect -8166 -16237 -8132 -16209
rect -8166 -16305 -8132 -16281
rect -8166 -16388 -8132 -16353
rect -7148 -15815 -7114 -15780
rect -7148 -15887 -7114 -15863
rect -7148 -15959 -7114 -15931
rect -7148 -16031 -7114 -15999
rect -7148 -16101 -7114 -16067
rect -7148 -16169 -7114 -16137
rect -7148 -16237 -7114 -16209
rect -7148 -16305 -7114 -16281
rect -7148 -16388 -7114 -16353
rect -6130 -15815 -6096 -15780
rect -6130 -15887 -6096 -15863
rect -6130 -15959 -6096 -15931
rect -6130 -16031 -6096 -15999
rect -6130 -16101 -6096 -16067
rect -6130 -16169 -6096 -16137
rect -6130 -16237 -6096 -16209
rect -6130 -16305 -6096 -16281
rect -6130 -16388 -6096 -16353
rect -5112 -15815 -5078 -15780
rect -5112 -15887 -5078 -15863
rect -5112 -15959 -5078 -15931
rect -5112 -16031 -5078 -15999
rect -5112 -16101 -5078 -16067
rect -5112 -16169 -5078 -16137
rect -5112 -16237 -5078 -16209
rect -5112 -16305 -5078 -16281
rect -5112 -16388 -5078 -16353
rect -4094 -15815 -4060 -15780
rect -4094 -15887 -4060 -15863
rect -4094 -15959 -4060 -15931
rect -4094 -16031 -4060 -15999
rect -4094 -16101 -4060 -16067
rect -4094 -16169 -4060 -16137
rect -4094 -16237 -4060 -16209
rect -4094 -16305 -4060 -16281
rect -4094 -16388 -4060 -16353
rect -3076 -15815 -3042 -15780
rect -3076 -15887 -3042 -15863
rect -3076 -15959 -3042 -15931
rect -3076 -16031 -3042 -15999
rect -3076 -16101 -3042 -16067
rect -3076 -16169 -3042 -16137
rect -3076 -16237 -3042 -16209
rect -3076 -16305 -3042 -16281
rect -3076 -16388 -3042 -16353
rect -2058 -15815 -2024 -15780
rect -2058 -15887 -2024 -15863
rect -2058 -15959 -2024 -15931
rect -2058 -16031 -2024 -15999
rect -2058 -16101 -2024 -16067
rect -2058 -16169 -2024 -16137
rect -2058 -16237 -2024 -16209
rect -2058 -16305 -2024 -16281
rect -2058 -16388 -2024 -16353
rect -1040 -15815 -1006 -15780
rect -1040 -15887 -1006 -15863
rect -1040 -15959 -1006 -15931
rect -1040 -16031 -1006 -15999
rect -1040 -16101 -1006 -16067
rect -1040 -16169 -1006 -16137
rect -1040 -16237 -1006 -16209
rect -1040 -16305 -1006 -16281
rect -1040 -16388 -1006 -16353
rect -22 -15815 12 -15780
rect -22 -15887 12 -15863
rect -22 -15959 12 -15931
rect -22 -16031 12 -15999
rect 2580 -15803 2614 -15771
rect 2580 -15871 2614 -15843
rect 2580 -15939 2614 -15915
rect 2580 -16022 2614 -15987
rect 3598 -15449 3632 -15414
rect 3598 -15521 3632 -15497
rect 3598 -15593 3632 -15565
rect 3598 -15665 3632 -15633
rect 3598 -15735 3632 -15701
rect 3598 -15803 3632 -15771
rect 3598 -15871 3632 -15843
rect 3598 -15939 3632 -15915
rect 3598 -16022 3632 -15987
rect 4616 -15449 4650 -15414
rect 4616 -15521 4650 -15497
rect 4616 -15593 4650 -15565
rect 4616 -15665 4650 -15633
rect 4616 -15735 4650 -15701
rect 4616 -15803 4650 -15771
rect 4616 -15871 4650 -15843
rect 4616 -15939 4650 -15915
rect 4616 -16022 4650 -15987
rect 5634 -15449 5668 -15414
rect 5634 -15521 5668 -15497
rect 5634 -15593 5668 -15565
rect 5634 -15665 5668 -15633
rect 5634 -15735 5668 -15701
rect 5634 -15803 5668 -15771
rect 5634 -15871 5668 -15843
rect 5634 -15939 5668 -15915
rect 5634 -16022 5668 -15987
rect 6652 -15449 6686 -15414
rect 6652 -15521 6686 -15497
rect 6652 -15593 6686 -15565
rect 6652 -15665 6686 -15633
rect 6652 -15735 6686 -15701
rect 6652 -15803 6686 -15771
rect 6652 -15871 6686 -15843
rect 6652 -15939 6686 -15915
rect 6652 -16022 6686 -15987
rect 7670 -15449 7704 -15414
rect 7670 -15521 7704 -15497
rect 7670 -15593 7704 -15565
rect 7670 -15665 7704 -15633
rect 7670 -15735 7704 -15701
rect 7670 -15803 7704 -15771
rect 7670 -15871 7704 -15843
rect 7670 -15939 7704 -15915
rect 7670 -16022 7704 -15987
rect 8688 -15449 8722 -15414
rect 8688 -15521 8722 -15497
rect 8688 -15593 8722 -15565
rect 8688 -15665 8722 -15633
rect 8688 -15735 8722 -15701
rect 8688 -15803 8722 -15771
rect 8688 -15871 8722 -15843
rect 8688 -15939 8722 -15915
rect 8688 -16022 8722 -15987
rect 9706 -15449 9740 -15414
rect 9706 -15521 9740 -15497
rect 9706 -15593 9740 -15565
rect 9706 -15665 9740 -15633
rect 9706 -15735 9740 -15701
rect 9706 -15803 9740 -15771
rect 9706 -15871 9740 -15843
rect 9706 -15939 9740 -15915
rect 9706 -16022 9740 -15987
rect 10724 -15449 10758 -15414
rect 10724 -15521 10758 -15497
rect 10724 -15593 10758 -15565
rect 10724 -15665 10758 -15633
rect 10724 -15735 10758 -15701
rect 10724 -15803 10758 -15771
rect 10724 -15871 10758 -15843
rect 10724 -15939 10758 -15915
rect 10724 -16022 10758 -15987
rect 11742 -15449 11776 -15414
rect 11742 -15521 11776 -15497
rect 11742 -15593 11776 -15565
rect 11742 -15665 11776 -15633
rect 11742 -15735 11776 -15701
rect 11742 -15803 11776 -15771
rect 11742 -15871 11776 -15843
rect 11742 -15939 11776 -15915
rect 11742 -16022 11776 -15987
rect 12760 -15449 12794 -15414
rect 12760 -15521 12794 -15497
rect 12760 -15593 12794 -15565
rect 12760 -15665 12794 -15633
rect 12760 -15735 12794 -15701
rect 12760 -15803 12794 -15771
rect 12760 -15871 12794 -15843
rect 12760 -15939 12794 -15915
rect 12760 -16022 12794 -15987
rect 13778 -15449 13812 -15414
rect 13778 -15521 13812 -15497
rect 13778 -15593 13812 -15565
rect 13778 -15665 13812 -15633
rect 13778 -15735 13812 -15701
rect 13778 -15803 13812 -15771
rect 13778 -15871 13812 -15843
rect 13778 -15939 13812 -15915
rect 13778 -16022 13812 -15987
rect 14796 -15449 14830 -15414
rect 14796 -15521 14830 -15497
rect 14796 -15593 14830 -15565
rect 14796 -15665 14830 -15633
rect 14796 -15735 14830 -15701
rect 14796 -15803 14830 -15771
rect 14796 -15871 14830 -15843
rect 14796 -15939 14830 -15915
rect 14796 -16022 14830 -15987
rect 15814 -15449 15848 -15414
rect 15814 -15521 15848 -15497
rect 15814 -15593 15848 -15565
rect 15814 -15665 15848 -15633
rect 15814 -15735 15848 -15701
rect 15814 -15803 15848 -15771
rect 15814 -15871 15848 -15843
rect 15814 -15939 15848 -15915
rect 15814 -16022 15848 -15987
rect 16832 -15449 16866 -15414
rect 16832 -15521 16866 -15497
rect 16832 -15593 16866 -15565
rect 16832 -15665 16866 -15633
rect 16832 -15735 16866 -15701
rect 16832 -15803 16866 -15771
rect 16832 -15871 16866 -15843
rect 16832 -15939 16866 -15915
rect 16832 -16022 16866 -15987
rect 17850 -15449 17884 -15414
rect 17850 -15521 17884 -15497
rect 17850 -15593 17884 -15565
rect 17850 -15665 17884 -15633
rect 17850 -15735 17884 -15701
rect 17850 -15803 17884 -15771
rect 17850 -15871 17884 -15843
rect 17850 -15939 17884 -15915
rect 17850 -16022 17884 -15987
rect 18868 -15449 18902 -15414
rect 18868 -15521 18902 -15497
rect 18868 -15593 18902 -15565
rect 18868 -15665 18902 -15633
rect 18868 -15735 18902 -15701
rect 18868 -15803 18902 -15771
rect 18868 -15871 18902 -15843
rect 18868 -15939 18902 -15915
rect 18868 -16022 18902 -15987
rect 19886 -15449 19920 -15414
rect 19886 -15521 19920 -15497
rect 19886 -15593 19920 -15565
rect 19886 -15665 19920 -15633
rect 19886 -15735 19920 -15701
rect 19886 -15803 19920 -15771
rect 19886 -15871 19920 -15843
rect 19886 -15939 19920 -15915
rect 19886 -16022 19920 -15987
rect 20904 -15449 20938 -15414
rect 20904 -15521 20938 -15497
rect 20904 -15593 20938 -15565
rect 20904 -15665 20938 -15633
rect 20904 -15735 20938 -15701
rect 20904 -15803 20938 -15771
rect 20904 -15871 20938 -15843
rect 20904 -15939 20938 -15915
rect 20904 -16022 20938 -15987
rect 21922 -15449 21956 -15414
rect 21922 -15521 21956 -15497
rect 21922 -15593 21956 -15565
rect 21922 -15665 21956 -15633
rect 21922 -15735 21956 -15701
rect 21922 -15803 21956 -15771
rect 21922 -15871 21956 -15843
rect 21922 -15939 21956 -15915
rect 21922 -16022 21956 -15987
rect 22940 -15449 22974 -15414
rect 22940 -15521 22974 -15497
rect 22940 -15593 22974 -15565
rect 22940 -15665 22974 -15633
rect 22940 -15735 22974 -15701
rect 22940 -15803 22974 -15771
rect 22940 -15871 22974 -15843
rect 22940 -15939 22974 -15915
rect 22940 -16022 22974 -15987
rect 24822 -15437 24855 -15375
rect 24889 -15437 24922 -15375
rect 24822 -15443 24922 -15437
rect 24822 -15509 24855 -15443
rect 24889 -15509 24922 -15443
rect 24822 -15511 24922 -15509
rect 24822 -15545 24855 -15511
rect 24889 -15545 24922 -15511
rect 24822 -15547 24922 -15545
rect 24822 -15613 24855 -15547
rect 24889 -15613 24922 -15547
rect 24822 -15619 24922 -15613
rect 24822 -15681 24855 -15619
rect 24889 -15681 24922 -15619
rect 24822 -15691 24922 -15681
rect 24822 -15749 24855 -15691
rect 24889 -15749 24922 -15691
rect 24822 -15763 24922 -15749
rect 24822 -15817 24855 -15763
rect 24889 -15817 24922 -15763
rect 24822 -15835 24922 -15817
rect 24822 -15885 24855 -15835
rect 24889 -15885 24922 -15835
rect 24822 -15907 24922 -15885
rect 24822 -15953 24855 -15907
rect 24889 -15953 24922 -15907
rect 24822 -15979 24922 -15953
rect 24822 -16021 24855 -15979
rect 24889 -16021 24922 -15979
rect 24822 -16051 24922 -16021
rect 10190 -16056 10250 -16052
rect 11218 -16056 11278 -16054
rect 13262 -16056 13322 -16052
rect -22 -16101 12 -16067
rect 2812 -16090 2851 -16056
rect 2885 -16090 2909 -16056
rect 2953 -16090 2981 -16056
rect 3021 -16090 3053 -16056
rect 3089 -16090 3123 -16056
rect 3159 -16090 3191 -16056
rect 3231 -16090 3259 -16056
rect 3303 -16090 3327 -16056
rect 3361 -16090 3400 -16056
rect 3830 -16090 3869 -16056
rect 3903 -16090 3927 -16056
rect 3971 -16090 3999 -16056
rect 4039 -16090 4071 -16056
rect 4107 -16090 4141 -16056
rect 4177 -16090 4209 -16056
rect 4249 -16090 4277 -16056
rect 4321 -16090 4345 -16056
rect 4379 -16090 4418 -16056
rect 4848 -16090 4887 -16056
rect 4921 -16090 4945 -16056
rect 4989 -16090 5017 -16056
rect 5057 -16090 5089 -16056
rect 5125 -16090 5159 -16056
rect 5195 -16090 5227 -16056
rect 5267 -16090 5295 -16056
rect 5339 -16090 5363 -16056
rect 5397 -16090 5436 -16056
rect 5866 -16090 5905 -16056
rect 5939 -16090 5963 -16056
rect 6007 -16090 6035 -16056
rect 6075 -16090 6107 -16056
rect 6143 -16090 6177 -16056
rect 6213 -16090 6245 -16056
rect 6285 -16090 6313 -16056
rect 6357 -16090 6381 -16056
rect 6415 -16090 6454 -16056
rect 6884 -16090 6923 -16056
rect 6957 -16090 6981 -16056
rect 7025 -16090 7053 -16056
rect 7093 -16090 7125 -16056
rect 7161 -16090 7195 -16056
rect 7231 -16090 7263 -16056
rect 7303 -16090 7331 -16056
rect 7375 -16090 7399 -16056
rect 7433 -16090 7472 -16056
rect 7902 -16090 7941 -16056
rect 7975 -16090 7999 -16056
rect 8043 -16090 8071 -16056
rect 8111 -16090 8143 -16056
rect 8179 -16090 8213 -16056
rect 8249 -16090 8281 -16056
rect 8321 -16090 8349 -16056
rect 8393 -16090 8417 -16056
rect 8451 -16090 8490 -16056
rect 8920 -16090 8959 -16056
rect 8993 -16090 9017 -16056
rect 9061 -16090 9089 -16056
rect 9129 -16090 9161 -16056
rect 9197 -16090 9231 -16056
rect 9267 -16090 9299 -16056
rect 9339 -16090 9367 -16056
rect 9411 -16090 9435 -16056
rect 9469 -16090 9508 -16056
rect 9938 -16090 9977 -16056
rect 10011 -16090 10035 -16056
rect 10079 -16090 10107 -16056
rect 10147 -16090 10179 -16056
rect 10215 -16090 10249 -16056
rect 10285 -16090 10317 -16056
rect 10357 -16090 10385 -16056
rect 10429 -16090 10453 -16056
rect 10487 -16090 10526 -16056
rect 10956 -16090 10995 -16056
rect 11029 -16090 11053 -16056
rect 11097 -16090 11125 -16056
rect 11165 -16090 11197 -16056
rect 11233 -16090 11267 -16056
rect 11303 -16090 11335 -16056
rect 11375 -16090 11403 -16056
rect 11447 -16090 11471 -16056
rect 11505 -16090 11544 -16056
rect 11974 -16090 12013 -16056
rect 12047 -16090 12071 -16056
rect 12115 -16090 12143 -16056
rect 12183 -16090 12215 -16056
rect 12251 -16090 12285 -16056
rect 12321 -16090 12353 -16056
rect 12393 -16090 12421 -16056
rect 12465 -16090 12489 -16056
rect 12523 -16090 12562 -16056
rect 12992 -16090 13031 -16056
rect 13065 -16090 13089 -16056
rect 13133 -16090 13161 -16056
rect 13201 -16090 13233 -16056
rect 13269 -16090 13303 -16056
rect 13339 -16090 13371 -16056
rect 13411 -16090 13439 -16056
rect 13483 -16090 13507 -16056
rect 13541 -16090 13580 -16056
rect 14010 -16090 14049 -16056
rect 14083 -16090 14107 -16056
rect 14151 -16090 14179 -16056
rect 14219 -16090 14251 -16056
rect 14287 -16090 14321 -16056
rect 14357 -16090 14389 -16056
rect 14429 -16090 14457 -16056
rect 14501 -16090 14525 -16056
rect 14559 -16090 14598 -16056
rect 15028 -16090 15067 -16056
rect 15101 -16090 15125 -16056
rect 15169 -16090 15197 -16056
rect 15237 -16090 15269 -16056
rect 15305 -16090 15339 -16056
rect 15375 -16090 15407 -16056
rect 15447 -16090 15475 -16056
rect 15519 -16090 15543 -16056
rect 15577 -16090 15616 -16056
rect 16046 -16090 16085 -16056
rect 16119 -16090 16143 -16056
rect 16187 -16090 16215 -16056
rect 16255 -16090 16287 -16056
rect 16323 -16090 16357 -16056
rect 16393 -16090 16425 -16056
rect 16465 -16090 16493 -16056
rect 16537 -16090 16561 -16056
rect 16595 -16090 16634 -16056
rect 17064 -16090 17103 -16056
rect 17137 -16090 17161 -16056
rect 17205 -16090 17233 -16056
rect 17273 -16090 17305 -16056
rect 17341 -16090 17375 -16056
rect 17411 -16090 17443 -16056
rect 17483 -16090 17511 -16056
rect 17555 -16090 17579 -16056
rect 17613 -16090 17652 -16056
rect 18082 -16090 18121 -16056
rect 18155 -16090 18179 -16056
rect 18223 -16090 18251 -16056
rect 18291 -16090 18323 -16056
rect 18359 -16090 18393 -16056
rect 18429 -16090 18461 -16056
rect 18501 -16090 18529 -16056
rect 18573 -16090 18597 -16056
rect 18631 -16090 18670 -16056
rect 19100 -16090 19139 -16056
rect 19173 -16090 19197 -16056
rect 19241 -16090 19269 -16056
rect 19309 -16090 19341 -16056
rect 19377 -16090 19411 -16056
rect 19447 -16090 19479 -16056
rect 19519 -16090 19547 -16056
rect 19591 -16090 19615 -16056
rect 19649 -16090 19688 -16056
rect 20118 -16090 20157 -16056
rect 20191 -16090 20215 -16056
rect 20259 -16090 20287 -16056
rect 20327 -16090 20359 -16056
rect 20395 -16090 20429 -16056
rect 20465 -16090 20497 -16056
rect 20537 -16090 20565 -16056
rect 20609 -16090 20633 -16056
rect 20667 -16090 20706 -16056
rect 21136 -16090 21175 -16056
rect 21209 -16090 21233 -16056
rect 21277 -16090 21305 -16056
rect 21345 -16090 21377 -16056
rect 21413 -16090 21447 -16056
rect 21483 -16090 21515 -16056
rect 21555 -16090 21583 -16056
rect 21627 -16090 21651 -16056
rect 21685 -16090 21724 -16056
rect 22154 -16090 22193 -16056
rect 22227 -16090 22251 -16056
rect 22295 -16090 22323 -16056
rect 22363 -16090 22395 -16056
rect 22431 -16090 22465 -16056
rect 22501 -16090 22533 -16056
rect 22573 -16090 22601 -16056
rect 22645 -16090 22669 -16056
rect 22703 -16090 22742 -16056
rect 24822 -16089 24855 -16051
rect 24889 -16089 24922 -16051
rect -22 -16169 12 -16137
rect -22 -16237 12 -16209
rect -22 -16305 12 -16281
rect -22 -16388 12 -16353
rect 24822 -16123 24922 -16089
rect 24822 -16157 24855 -16123
rect 24889 -16157 24922 -16123
rect 24822 -16191 24922 -16157
rect 24822 -16229 24855 -16191
rect 24889 -16229 24922 -16191
rect 24822 -16259 24922 -16229
rect 24822 -16301 24855 -16259
rect 24889 -16301 24922 -16259
rect 24822 -16327 24922 -16301
rect 24822 -16373 24855 -16327
rect 24889 -16373 24922 -16327
rect -12322 -16445 -12289 -16395
rect -12255 -16445 -12222 -16395
rect 24822 -16395 24922 -16373
rect -7670 -16422 -7610 -16420
rect -6656 -16422 -6596 -16420
rect -2582 -16422 -2522 -16420
rect -1566 -16422 -1506 -16420
rect -12322 -16463 -12222 -16445
rect -8952 -16456 -8913 -16422
rect -8879 -16456 -8855 -16422
rect -8811 -16456 -8783 -16422
rect -8743 -16456 -8711 -16422
rect -8675 -16456 -8641 -16422
rect -8605 -16456 -8573 -16422
rect -8533 -16456 -8505 -16422
rect -8461 -16456 -8437 -16422
rect -8403 -16456 -8364 -16422
rect -7934 -16456 -7895 -16422
rect -7861 -16456 -7837 -16422
rect -7793 -16456 -7765 -16422
rect -7725 -16456 -7693 -16422
rect -7657 -16456 -7623 -16422
rect -7587 -16456 -7555 -16422
rect -7515 -16456 -7487 -16422
rect -7443 -16456 -7419 -16422
rect -7385 -16456 -7346 -16422
rect -6916 -16456 -6877 -16422
rect -6843 -16456 -6819 -16422
rect -6775 -16456 -6747 -16422
rect -6707 -16456 -6675 -16422
rect -6639 -16456 -6605 -16422
rect -6569 -16456 -6537 -16422
rect -6497 -16456 -6469 -16422
rect -6425 -16456 -6401 -16422
rect -6367 -16456 -6328 -16422
rect -5898 -16456 -5859 -16422
rect -5825 -16456 -5801 -16422
rect -5757 -16456 -5729 -16422
rect -5689 -16456 -5657 -16422
rect -5621 -16456 -5587 -16422
rect -5551 -16456 -5519 -16422
rect -5479 -16456 -5451 -16422
rect -5407 -16456 -5383 -16422
rect -5349 -16456 -5310 -16422
rect -4880 -16456 -4841 -16422
rect -4807 -16456 -4783 -16422
rect -4739 -16456 -4711 -16422
rect -4671 -16456 -4639 -16422
rect -4603 -16456 -4569 -16422
rect -4533 -16456 -4501 -16422
rect -4461 -16456 -4433 -16422
rect -4389 -16456 -4365 -16422
rect -4331 -16456 -4292 -16422
rect -3862 -16456 -3823 -16422
rect -3789 -16456 -3765 -16422
rect -3721 -16456 -3693 -16422
rect -3653 -16456 -3621 -16422
rect -3585 -16456 -3551 -16422
rect -3515 -16456 -3483 -16422
rect -3443 -16456 -3415 -16422
rect -3371 -16456 -3347 -16422
rect -3313 -16456 -3274 -16422
rect -2844 -16456 -2805 -16422
rect -2771 -16456 -2747 -16422
rect -2703 -16456 -2675 -16422
rect -2635 -16456 -2603 -16422
rect -2567 -16456 -2533 -16422
rect -2497 -16456 -2465 -16422
rect -2425 -16456 -2397 -16422
rect -2353 -16456 -2329 -16422
rect -2295 -16456 -2256 -16422
rect -1826 -16456 -1787 -16422
rect -1753 -16456 -1729 -16422
rect -1685 -16456 -1657 -16422
rect -1617 -16456 -1585 -16422
rect -1549 -16456 -1515 -16422
rect -1479 -16456 -1447 -16422
rect -1407 -16456 -1379 -16422
rect -1335 -16456 -1311 -16422
rect -1277 -16456 -1238 -16422
rect -808 -16456 -769 -16422
rect -735 -16456 -711 -16422
rect -667 -16456 -639 -16422
rect -599 -16456 -567 -16422
rect -531 -16456 -497 -16422
rect -461 -16456 -429 -16422
rect -389 -16456 -361 -16422
rect -317 -16456 -293 -16422
rect -259 -16456 -220 -16422
rect 24822 -16445 24855 -16395
rect 24889 -16445 24922 -16395
rect -12322 -16517 -12289 -16463
rect -12255 -16517 -12222 -16463
rect -12322 -16531 -12222 -16517
rect 24822 -16463 24922 -16445
rect 24822 -16517 24855 -16463
rect 24889 -16517 24922 -16463
rect -12322 -16589 -12289 -16531
rect -12255 -16589 -12222 -16531
rect -8952 -16564 -8913 -16530
rect -8879 -16564 -8855 -16530
rect -8811 -16564 -8783 -16530
rect -8743 -16564 -8711 -16530
rect -8675 -16564 -8641 -16530
rect -8605 -16564 -8573 -16530
rect -8533 -16564 -8505 -16530
rect -8461 -16564 -8437 -16530
rect -8403 -16564 -8364 -16530
rect -7934 -16564 -7895 -16530
rect -7861 -16564 -7837 -16530
rect -7793 -16564 -7765 -16530
rect -7725 -16564 -7693 -16530
rect -7657 -16564 -7623 -16530
rect -7587 -16564 -7555 -16530
rect -7515 -16564 -7487 -16530
rect -7443 -16564 -7419 -16530
rect -7385 -16564 -7346 -16530
rect -6916 -16564 -6877 -16530
rect -6843 -16564 -6819 -16530
rect -6775 -16564 -6747 -16530
rect -6707 -16564 -6675 -16530
rect -6639 -16564 -6605 -16530
rect -6569 -16564 -6537 -16530
rect -6497 -16564 -6469 -16530
rect -6425 -16564 -6401 -16530
rect -6367 -16564 -6328 -16530
rect -5898 -16564 -5859 -16530
rect -5825 -16564 -5801 -16530
rect -5757 -16564 -5729 -16530
rect -5689 -16564 -5657 -16530
rect -5621 -16564 -5587 -16530
rect -5551 -16564 -5519 -16530
rect -5479 -16564 -5451 -16530
rect -5407 -16564 -5383 -16530
rect -5349 -16564 -5310 -16530
rect -4880 -16564 -4841 -16530
rect -4807 -16564 -4783 -16530
rect -4739 -16564 -4711 -16530
rect -4671 -16564 -4639 -16530
rect -4603 -16564 -4569 -16530
rect -4533 -16564 -4501 -16530
rect -4461 -16564 -4433 -16530
rect -4389 -16564 -4365 -16530
rect -4331 -16564 -4292 -16530
rect -3862 -16564 -3823 -16530
rect -3789 -16564 -3765 -16530
rect -3721 -16564 -3693 -16530
rect -3653 -16564 -3621 -16530
rect -3585 -16564 -3551 -16530
rect -3515 -16564 -3483 -16530
rect -3443 -16564 -3415 -16530
rect -3371 -16564 -3347 -16530
rect -3313 -16564 -3274 -16530
rect -2844 -16564 -2805 -16530
rect -2771 -16564 -2747 -16530
rect -2703 -16564 -2675 -16530
rect -2635 -16564 -2603 -16530
rect -2567 -16564 -2533 -16530
rect -2497 -16564 -2465 -16530
rect -2425 -16564 -2397 -16530
rect -2353 -16564 -2329 -16530
rect -2295 -16564 -2256 -16530
rect -1826 -16564 -1787 -16530
rect -1753 -16564 -1729 -16530
rect -1685 -16564 -1657 -16530
rect -1617 -16564 -1585 -16530
rect -1549 -16564 -1515 -16530
rect -1479 -16564 -1447 -16530
rect -1407 -16564 -1379 -16530
rect -1335 -16564 -1311 -16530
rect -1277 -16564 -1238 -16530
rect -808 -16564 -769 -16530
rect -735 -16564 -711 -16530
rect -667 -16564 -639 -16530
rect -599 -16564 -567 -16530
rect -531 -16564 -497 -16530
rect -461 -16564 -429 -16530
rect -389 -16564 -361 -16530
rect -317 -16564 -293 -16530
rect -259 -16564 -220 -16530
rect 24822 -16531 24922 -16517
rect -12322 -16599 -12222 -16589
rect -12322 -16661 -12289 -16599
rect -12255 -16661 -12222 -16599
rect -12322 -16667 -12222 -16661
rect -12322 -16733 -12289 -16667
rect -12255 -16733 -12222 -16667
rect -12322 -16735 -12222 -16733
rect -12322 -16769 -12289 -16735
rect -12255 -16769 -12222 -16735
rect -12322 -16771 -12222 -16769
rect -12322 -16837 -12289 -16771
rect -12255 -16837 -12222 -16771
rect -12322 -16843 -12222 -16837
rect -12322 -16905 -12289 -16843
rect -12255 -16905 -12222 -16843
rect -12322 -16915 -12222 -16905
rect -12322 -16973 -12289 -16915
rect -12255 -16973 -12222 -16915
rect -12322 -16987 -12222 -16973
rect -12322 -17041 -12289 -16987
rect -12255 -17041 -12222 -16987
rect -12322 -17059 -12222 -17041
rect -12322 -17109 -12289 -17059
rect -12255 -17109 -12222 -17059
rect -12322 -17131 -12222 -17109
rect -12322 -17177 -12289 -17131
rect -12255 -17177 -12222 -17131
rect -12322 -17203 -12222 -17177
rect -12322 -17245 -12289 -17203
rect -12255 -17245 -12222 -17203
rect -9184 -16633 -9150 -16598
rect -9184 -16705 -9150 -16681
rect -9184 -16777 -9150 -16749
rect -9184 -16849 -9150 -16817
rect -9184 -16919 -9150 -16885
rect -9184 -16987 -9150 -16955
rect -9184 -17055 -9150 -17027
rect -9184 -17123 -9150 -17099
rect -9184 -17206 -9150 -17171
rect -8166 -16633 -8132 -16598
rect -8166 -16705 -8132 -16681
rect -8166 -16777 -8132 -16749
rect -8166 -16849 -8132 -16817
rect -8166 -16919 -8132 -16885
rect -8166 -16987 -8132 -16955
rect -8166 -17055 -8132 -17027
rect -8166 -17123 -8132 -17099
rect -8166 -17206 -8132 -17171
rect -7148 -16633 -7114 -16598
rect -7148 -16705 -7114 -16681
rect -7148 -16777 -7114 -16749
rect -7148 -16849 -7114 -16817
rect -7148 -16919 -7114 -16885
rect -7148 -16987 -7114 -16955
rect -7148 -17055 -7114 -17027
rect -7148 -17123 -7114 -17099
rect -7148 -17206 -7114 -17171
rect -6130 -16633 -6096 -16598
rect -6130 -16705 -6096 -16681
rect -6130 -16777 -6096 -16749
rect -6130 -16849 -6096 -16817
rect -6130 -16919 -6096 -16885
rect -6130 -16987 -6096 -16955
rect -6130 -17055 -6096 -17027
rect -6130 -17123 -6096 -17099
rect -6130 -17206 -6096 -17171
rect -5112 -16633 -5078 -16598
rect -5112 -16705 -5078 -16681
rect -5112 -16777 -5078 -16749
rect -5112 -16849 -5078 -16817
rect -5112 -16919 -5078 -16885
rect -5112 -16987 -5078 -16955
rect -5112 -17055 -5078 -17027
rect -5112 -17123 -5078 -17099
rect -5112 -17206 -5078 -17171
rect -4094 -16633 -4060 -16598
rect -4094 -16705 -4060 -16681
rect -4094 -16777 -4060 -16749
rect -4094 -16849 -4060 -16817
rect -4094 -16919 -4060 -16885
rect -4094 -16987 -4060 -16955
rect -4094 -17055 -4060 -17027
rect -4094 -17123 -4060 -17099
rect -4094 -17206 -4060 -17171
rect -3076 -16633 -3042 -16598
rect -3076 -16705 -3042 -16681
rect -3076 -16777 -3042 -16749
rect -3076 -16849 -3042 -16817
rect -3076 -16919 -3042 -16885
rect -3076 -16987 -3042 -16955
rect -3076 -17055 -3042 -17027
rect -3076 -17123 -3042 -17099
rect -3076 -17206 -3042 -17171
rect -2058 -16633 -2024 -16598
rect -2058 -16705 -2024 -16681
rect -2058 -16777 -2024 -16749
rect -2058 -16849 -2024 -16817
rect -2058 -16919 -2024 -16885
rect -2058 -16987 -2024 -16955
rect -2058 -17055 -2024 -17027
rect -2058 -17123 -2024 -17099
rect -2058 -17206 -2024 -17171
rect -1040 -16633 -1006 -16598
rect -1040 -16705 -1006 -16681
rect -1040 -16777 -1006 -16749
rect -1040 -16849 -1006 -16817
rect -1040 -16919 -1006 -16885
rect -1040 -16987 -1006 -16955
rect -1040 -17055 -1006 -17027
rect -1040 -17123 -1006 -17099
rect -1040 -17206 -1006 -17171
rect -22 -16633 12 -16598
rect 2812 -16614 2851 -16580
rect 2885 -16614 2909 -16580
rect 2953 -16614 2981 -16580
rect 3021 -16614 3053 -16580
rect 3089 -16614 3123 -16580
rect 3159 -16614 3191 -16580
rect 3231 -16614 3259 -16580
rect 3303 -16614 3327 -16580
rect 3361 -16614 3400 -16580
rect 3830 -16614 3869 -16580
rect 3903 -16614 3927 -16580
rect 3971 -16614 3999 -16580
rect 4039 -16614 4071 -16580
rect 4107 -16614 4141 -16580
rect 4177 -16614 4209 -16580
rect 4249 -16614 4277 -16580
rect 4321 -16614 4345 -16580
rect 4379 -16614 4418 -16580
rect 4848 -16614 4887 -16580
rect 4921 -16614 4945 -16580
rect 4989 -16614 5017 -16580
rect 5057 -16614 5089 -16580
rect 5125 -16614 5159 -16580
rect 5195 -16614 5227 -16580
rect 5267 -16614 5295 -16580
rect 5339 -16614 5363 -16580
rect 5397 -16614 5436 -16580
rect 5866 -16614 5905 -16580
rect 5939 -16614 5963 -16580
rect 6007 -16614 6035 -16580
rect 6075 -16614 6107 -16580
rect 6143 -16614 6177 -16580
rect 6213 -16614 6245 -16580
rect 6285 -16614 6313 -16580
rect 6357 -16614 6381 -16580
rect 6415 -16614 6454 -16580
rect 6884 -16614 6923 -16580
rect 6957 -16614 6981 -16580
rect 7025 -16614 7053 -16580
rect 7093 -16614 7125 -16580
rect 7161 -16614 7195 -16580
rect 7231 -16614 7263 -16580
rect 7303 -16614 7331 -16580
rect 7375 -16614 7399 -16580
rect 7433 -16614 7472 -16580
rect 7902 -16614 7941 -16580
rect 7975 -16614 7999 -16580
rect 8043 -16614 8071 -16580
rect 8111 -16614 8143 -16580
rect 8179 -16614 8213 -16580
rect 8249 -16614 8281 -16580
rect 8321 -16614 8349 -16580
rect 8393 -16614 8417 -16580
rect 8451 -16614 8490 -16580
rect 8920 -16614 8959 -16580
rect 8993 -16614 9017 -16580
rect 9061 -16614 9089 -16580
rect 9129 -16614 9161 -16580
rect 9197 -16614 9231 -16580
rect 9267 -16614 9299 -16580
rect 9339 -16614 9367 -16580
rect 9411 -16614 9435 -16580
rect 9469 -16614 9508 -16580
rect 9938 -16614 9977 -16580
rect 10011 -16614 10035 -16580
rect 10079 -16614 10107 -16580
rect 10147 -16614 10179 -16580
rect 10215 -16614 10249 -16580
rect 10285 -16614 10317 -16580
rect 10357 -16614 10385 -16580
rect 10429 -16614 10453 -16580
rect 10487 -16614 10526 -16580
rect 10956 -16614 10995 -16580
rect 11029 -16614 11053 -16580
rect 11097 -16614 11125 -16580
rect 11165 -16614 11197 -16580
rect 11233 -16614 11267 -16580
rect 11303 -16614 11335 -16580
rect 11375 -16614 11403 -16580
rect 11447 -16614 11471 -16580
rect 11505 -16614 11544 -16580
rect 11974 -16614 12013 -16580
rect 12047 -16614 12071 -16580
rect 12115 -16614 12143 -16580
rect 12183 -16614 12215 -16580
rect 12251 -16614 12285 -16580
rect 12321 -16614 12353 -16580
rect 12393 -16614 12421 -16580
rect 12465 -16614 12489 -16580
rect 12523 -16614 12562 -16580
rect 12992 -16614 13031 -16580
rect 13065 -16614 13089 -16580
rect 13133 -16614 13161 -16580
rect 13201 -16614 13233 -16580
rect 13269 -16614 13303 -16580
rect 13339 -16614 13371 -16580
rect 13411 -16614 13439 -16580
rect 13483 -16614 13507 -16580
rect 13541 -16614 13580 -16580
rect 14010 -16614 14049 -16580
rect 14083 -16614 14107 -16580
rect 14151 -16614 14179 -16580
rect 14219 -16614 14251 -16580
rect 14287 -16614 14321 -16580
rect 14357 -16614 14389 -16580
rect 14429 -16614 14457 -16580
rect 14501 -16614 14525 -16580
rect 14559 -16614 14598 -16580
rect 15028 -16614 15067 -16580
rect 15101 -16614 15125 -16580
rect 15169 -16614 15197 -16580
rect 15237 -16614 15269 -16580
rect 15305 -16614 15339 -16580
rect 15375 -16614 15407 -16580
rect 15447 -16614 15475 -16580
rect 15519 -16614 15543 -16580
rect 15577 -16614 15616 -16580
rect 16046 -16614 16085 -16580
rect 16119 -16614 16143 -16580
rect 16187 -16614 16215 -16580
rect 16255 -16614 16287 -16580
rect 16323 -16614 16357 -16580
rect 16393 -16614 16425 -16580
rect 16465 -16614 16493 -16580
rect 16537 -16614 16561 -16580
rect 16595 -16614 16634 -16580
rect 17064 -16614 17103 -16580
rect 17137 -16614 17161 -16580
rect 17205 -16614 17233 -16580
rect 17273 -16614 17305 -16580
rect 17341 -16614 17375 -16580
rect 17411 -16614 17443 -16580
rect 17483 -16614 17511 -16580
rect 17555 -16614 17579 -16580
rect 17613 -16614 17652 -16580
rect 18082 -16614 18121 -16580
rect 18155 -16614 18179 -16580
rect 18223 -16614 18251 -16580
rect 18291 -16614 18323 -16580
rect 18359 -16614 18393 -16580
rect 18429 -16614 18461 -16580
rect 18501 -16614 18529 -16580
rect 18573 -16614 18597 -16580
rect 18631 -16614 18670 -16580
rect 19100 -16614 19139 -16580
rect 19173 -16614 19197 -16580
rect 19241 -16614 19269 -16580
rect 19309 -16614 19341 -16580
rect 19377 -16614 19411 -16580
rect 19447 -16614 19479 -16580
rect 19519 -16614 19547 -16580
rect 19591 -16614 19615 -16580
rect 19649 -16614 19688 -16580
rect 20118 -16614 20157 -16580
rect 20191 -16614 20215 -16580
rect 20259 -16614 20287 -16580
rect 20327 -16614 20359 -16580
rect 20395 -16614 20429 -16580
rect 20465 -16614 20497 -16580
rect 20537 -16614 20565 -16580
rect 20609 -16614 20633 -16580
rect 20667 -16614 20706 -16580
rect 21136 -16614 21175 -16580
rect 21209 -16614 21233 -16580
rect 21277 -16614 21305 -16580
rect 21345 -16614 21377 -16580
rect 21413 -16614 21447 -16580
rect 21483 -16614 21515 -16580
rect 21555 -16614 21583 -16580
rect 21627 -16614 21651 -16580
rect 21685 -16614 21724 -16580
rect 22154 -16614 22193 -16580
rect 22227 -16614 22251 -16580
rect 22295 -16614 22323 -16580
rect 22363 -16614 22395 -16580
rect 22431 -16614 22465 -16580
rect 22501 -16614 22533 -16580
rect 22573 -16614 22601 -16580
rect 22645 -16614 22669 -16580
rect 22703 -16614 22742 -16580
rect 24822 -16589 24855 -16531
rect 24889 -16589 24922 -16531
rect 24822 -16599 24922 -16589
rect -22 -16705 12 -16681
rect -22 -16777 12 -16749
rect -22 -16849 12 -16817
rect -22 -16919 12 -16885
rect -22 -16987 12 -16955
rect -22 -17055 12 -17027
rect -22 -17123 12 -17099
rect -22 -17206 12 -17171
rect 2580 -16683 2614 -16648
rect 2580 -16755 2614 -16731
rect 2580 -16827 2614 -16799
rect 2580 -16899 2614 -16867
rect 2580 -16969 2614 -16935
rect 2580 -17037 2614 -17005
rect 2580 -17105 2614 -17077
rect 2580 -17173 2614 -17149
rect -7666 -17240 -7606 -17238
rect -6652 -17240 -6592 -17238
rect -2578 -17240 -2518 -17238
rect -1562 -17240 -1502 -17238
rect -12322 -17275 -12222 -17245
rect -8952 -17274 -8913 -17240
rect -8879 -17274 -8855 -17240
rect -8811 -17274 -8783 -17240
rect -8743 -17274 -8711 -17240
rect -8675 -17274 -8641 -17240
rect -8605 -17274 -8573 -17240
rect -8533 -17274 -8505 -17240
rect -8461 -17274 -8437 -17240
rect -8403 -17274 -8364 -17240
rect -7934 -17274 -7895 -17240
rect -7861 -17274 -7837 -17240
rect -7793 -17274 -7765 -17240
rect -7725 -17274 -7693 -17240
rect -7657 -17274 -7623 -17240
rect -7587 -17274 -7555 -17240
rect -7515 -17274 -7487 -17240
rect -7443 -17274 -7419 -17240
rect -7385 -17274 -7346 -17240
rect -6916 -17274 -6877 -17240
rect -6843 -17274 -6819 -17240
rect -6775 -17274 -6747 -17240
rect -6707 -17274 -6675 -17240
rect -6639 -17274 -6605 -17240
rect -6569 -17274 -6537 -17240
rect -6497 -17274 -6469 -17240
rect -6425 -17274 -6401 -17240
rect -6367 -17274 -6328 -17240
rect -5898 -17274 -5859 -17240
rect -5825 -17274 -5801 -17240
rect -5757 -17274 -5729 -17240
rect -5689 -17274 -5657 -17240
rect -5621 -17274 -5587 -17240
rect -5551 -17274 -5519 -17240
rect -5479 -17274 -5451 -17240
rect -5407 -17274 -5383 -17240
rect -5349 -17274 -5310 -17240
rect -4880 -17274 -4841 -17240
rect -4807 -17274 -4783 -17240
rect -4739 -17274 -4711 -17240
rect -4671 -17274 -4639 -17240
rect -4603 -17274 -4569 -17240
rect -4533 -17274 -4501 -17240
rect -4461 -17274 -4433 -17240
rect -4389 -17274 -4365 -17240
rect -4331 -17274 -4292 -17240
rect -3862 -17274 -3823 -17240
rect -3789 -17274 -3765 -17240
rect -3721 -17274 -3693 -17240
rect -3653 -17274 -3621 -17240
rect -3585 -17274 -3551 -17240
rect -3515 -17274 -3483 -17240
rect -3443 -17274 -3415 -17240
rect -3371 -17274 -3347 -17240
rect -3313 -17274 -3274 -17240
rect -2844 -17274 -2805 -17240
rect -2771 -17274 -2747 -17240
rect -2703 -17274 -2675 -17240
rect -2635 -17274 -2603 -17240
rect -2567 -17274 -2533 -17240
rect -2497 -17274 -2465 -17240
rect -2425 -17274 -2397 -17240
rect -2353 -17274 -2329 -17240
rect -2295 -17274 -2256 -17240
rect -1826 -17274 -1787 -17240
rect -1753 -17274 -1729 -17240
rect -1685 -17274 -1657 -17240
rect -1617 -17274 -1585 -17240
rect -1549 -17274 -1515 -17240
rect -1479 -17274 -1447 -17240
rect -1407 -17274 -1379 -17240
rect -1335 -17274 -1311 -17240
rect -1277 -17274 -1238 -17240
rect -808 -17274 -769 -17240
rect -735 -17274 -711 -17240
rect -667 -17274 -639 -17240
rect -599 -17274 -567 -17240
rect -531 -17274 -497 -17240
rect -461 -17274 -429 -17240
rect -389 -17274 -361 -17240
rect -317 -17274 -293 -17240
rect -259 -17274 -220 -17240
rect 2580 -17256 2614 -17221
rect 3598 -16683 3632 -16648
rect 3598 -16755 3632 -16731
rect 3598 -16827 3632 -16799
rect 3598 -16899 3632 -16867
rect 3598 -16969 3632 -16935
rect 3598 -17037 3632 -17005
rect 3598 -17105 3632 -17077
rect 3598 -17173 3632 -17149
rect 3598 -17256 3632 -17221
rect 4616 -16683 4650 -16648
rect 4616 -16755 4650 -16731
rect 4616 -16827 4650 -16799
rect 4616 -16899 4650 -16867
rect 4616 -16969 4650 -16935
rect 4616 -17037 4650 -17005
rect 4616 -17105 4650 -17077
rect 4616 -17173 4650 -17149
rect 4616 -17256 4650 -17221
rect 5634 -16683 5668 -16648
rect 5634 -16755 5668 -16731
rect 5634 -16827 5668 -16799
rect 5634 -16899 5668 -16867
rect 5634 -16969 5668 -16935
rect 5634 -17037 5668 -17005
rect 5634 -17105 5668 -17077
rect 5634 -17173 5668 -17149
rect 5634 -17256 5668 -17221
rect 6652 -16683 6686 -16648
rect 6652 -16755 6686 -16731
rect 6652 -16827 6686 -16799
rect 6652 -16899 6686 -16867
rect 6652 -16969 6686 -16935
rect 6652 -17037 6686 -17005
rect 6652 -17105 6686 -17077
rect 6652 -17173 6686 -17149
rect 6652 -17256 6686 -17221
rect 7670 -16683 7704 -16648
rect 7670 -16755 7704 -16731
rect 7670 -16827 7704 -16799
rect 7670 -16899 7704 -16867
rect 7670 -16969 7704 -16935
rect 7670 -17037 7704 -17005
rect 7670 -17105 7704 -17077
rect 7670 -17173 7704 -17149
rect 7670 -17256 7704 -17221
rect 8688 -16683 8722 -16648
rect 8688 -16755 8722 -16731
rect 8688 -16827 8722 -16799
rect 8688 -16899 8722 -16867
rect 8688 -16969 8722 -16935
rect 8688 -17037 8722 -17005
rect 8688 -17105 8722 -17077
rect 8688 -17173 8722 -17149
rect 8688 -17256 8722 -17221
rect 9706 -16683 9740 -16648
rect 9706 -16755 9740 -16731
rect 9706 -16827 9740 -16799
rect 9706 -16899 9740 -16867
rect 9706 -16969 9740 -16935
rect 9706 -17037 9740 -17005
rect 9706 -17105 9740 -17077
rect 9706 -17173 9740 -17149
rect 9706 -17256 9740 -17221
rect 10724 -16683 10758 -16648
rect 10724 -16755 10758 -16731
rect 10724 -16827 10758 -16799
rect 10724 -16899 10758 -16867
rect 10724 -16969 10758 -16935
rect 10724 -17037 10758 -17005
rect 10724 -17105 10758 -17077
rect 10724 -17173 10758 -17149
rect 10724 -17256 10758 -17221
rect 11742 -16683 11776 -16648
rect 11742 -16755 11776 -16731
rect 11742 -16827 11776 -16799
rect 11742 -16899 11776 -16867
rect 11742 -16969 11776 -16935
rect 11742 -17037 11776 -17005
rect 11742 -17105 11776 -17077
rect 11742 -17173 11776 -17149
rect 11742 -17256 11776 -17221
rect 12760 -16683 12794 -16648
rect 12760 -16755 12794 -16731
rect 12760 -16827 12794 -16799
rect 12760 -16899 12794 -16867
rect 12760 -16969 12794 -16935
rect 12760 -17037 12794 -17005
rect 12760 -17105 12794 -17077
rect 12760 -17173 12794 -17149
rect 12760 -17256 12794 -17221
rect 13778 -16683 13812 -16648
rect 13778 -16755 13812 -16731
rect 13778 -16827 13812 -16799
rect 13778 -16899 13812 -16867
rect 13778 -16969 13812 -16935
rect 13778 -17037 13812 -17005
rect 13778 -17105 13812 -17077
rect 13778 -17173 13812 -17149
rect 13778 -17256 13812 -17221
rect 14796 -16683 14830 -16648
rect 14796 -16755 14830 -16731
rect 14796 -16827 14830 -16799
rect 14796 -16899 14830 -16867
rect 14796 -16969 14830 -16935
rect 14796 -17037 14830 -17005
rect 14796 -17105 14830 -17077
rect 14796 -17173 14830 -17149
rect 14796 -17256 14830 -17221
rect 15814 -16683 15848 -16648
rect 15814 -16755 15848 -16731
rect 15814 -16827 15848 -16799
rect 15814 -16899 15848 -16867
rect 15814 -16969 15848 -16935
rect 15814 -17037 15848 -17005
rect 15814 -17105 15848 -17077
rect 15814 -17173 15848 -17149
rect 15814 -17256 15848 -17221
rect 16832 -16683 16866 -16648
rect 16832 -16755 16866 -16731
rect 16832 -16827 16866 -16799
rect 16832 -16899 16866 -16867
rect 16832 -16969 16866 -16935
rect 16832 -17037 16866 -17005
rect 16832 -17105 16866 -17077
rect 16832 -17173 16866 -17149
rect 16832 -17256 16866 -17221
rect 17850 -16683 17884 -16648
rect 17850 -16755 17884 -16731
rect 17850 -16827 17884 -16799
rect 17850 -16899 17884 -16867
rect 17850 -16969 17884 -16935
rect 17850 -17037 17884 -17005
rect 17850 -17105 17884 -17077
rect 17850 -17173 17884 -17149
rect 17850 -17256 17884 -17221
rect 18868 -16683 18902 -16648
rect 18868 -16755 18902 -16731
rect 18868 -16827 18902 -16799
rect 18868 -16899 18902 -16867
rect 18868 -16969 18902 -16935
rect 18868 -17037 18902 -17005
rect 18868 -17105 18902 -17077
rect 18868 -17173 18902 -17149
rect 18868 -17256 18902 -17221
rect 19886 -16683 19920 -16648
rect 19886 -16755 19920 -16731
rect 19886 -16827 19920 -16799
rect 19886 -16899 19920 -16867
rect 19886 -16969 19920 -16935
rect 19886 -17037 19920 -17005
rect 19886 -17105 19920 -17077
rect 19886 -17173 19920 -17149
rect 19886 -17256 19920 -17221
rect 20904 -16683 20938 -16648
rect 20904 -16755 20938 -16731
rect 20904 -16827 20938 -16799
rect 20904 -16899 20938 -16867
rect 20904 -16969 20938 -16935
rect 20904 -17037 20938 -17005
rect 20904 -17105 20938 -17077
rect 20904 -17173 20938 -17149
rect 20904 -17256 20938 -17221
rect 21922 -16683 21956 -16648
rect 21922 -16755 21956 -16731
rect 21922 -16827 21956 -16799
rect 21922 -16899 21956 -16867
rect 21922 -16969 21956 -16935
rect 21922 -17037 21956 -17005
rect 21922 -17105 21956 -17077
rect 21922 -17173 21956 -17149
rect 21922 -17256 21956 -17221
rect 22940 -16683 22974 -16648
rect 22940 -16755 22974 -16731
rect 22940 -16827 22974 -16799
rect 22940 -16899 22974 -16867
rect 22940 -16969 22974 -16935
rect 22940 -17037 22974 -17005
rect 22940 -17105 22974 -17077
rect 22940 -17173 22974 -17149
rect 22940 -17256 22974 -17221
rect 24822 -16661 24855 -16599
rect 24889 -16661 24922 -16599
rect 24822 -16667 24922 -16661
rect 24822 -16733 24855 -16667
rect 24889 -16733 24922 -16667
rect 24822 -16735 24922 -16733
rect 24822 -16769 24855 -16735
rect 24889 -16769 24922 -16735
rect 24822 -16771 24922 -16769
rect 24822 -16837 24855 -16771
rect 24889 -16837 24922 -16771
rect 24822 -16843 24922 -16837
rect 24822 -16905 24855 -16843
rect 24889 -16905 24922 -16843
rect 24822 -16915 24922 -16905
rect 24822 -16973 24855 -16915
rect 24889 -16973 24922 -16915
rect 24822 -16987 24922 -16973
rect 24822 -17041 24855 -16987
rect 24889 -17041 24922 -16987
rect 24822 -17059 24922 -17041
rect 24822 -17109 24855 -17059
rect 24889 -17109 24922 -17059
rect 24822 -17131 24922 -17109
rect 24822 -17177 24855 -17131
rect 24889 -17177 24922 -17131
rect 24822 -17203 24922 -17177
rect 24822 -17245 24855 -17203
rect 24889 -17245 24922 -17203
rect -12322 -17313 -12289 -17275
rect -12255 -17313 -12222 -17275
rect 24822 -17275 24922 -17245
rect -12322 -17347 -12222 -17313
rect 2812 -17324 2851 -17290
rect 2885 -17324 2909 -17290
rect 2953 -17324 2981 -17290
rect 3021 -17324 3053 -17290
rect 3089 -17324 3123 -17290
rect 3159 -17324 3191 -17290
rect 3231 -17324 3259 -17290
rect 3303 -17324 3327 -17290
rect 3361 -17324 3400 -17290
rect 3830 -17324 3869 -17290
rect 3903 -17324 3927 -17290
rect 3971 -17324 3999 -17290
rect 4039 -17324 4071 -17290
rect 4107 -17324 4141 -17290
rect 4177 -17324 4209 -17290
rect 4249 -17324 4277 -17290
rect 4321 -17324 4345 -17290
rect 4379 -17324 4418 -17290
rect 4848 -17324 4887 -17290
rect 4921 -17324 4945 -17290
rect 4989 -17324 5017 -17290
rect 5057 -17324 5089 -17290
rect 5125 -17324 5159 -17290
rect 5195 -17324 5227 -17290
rect 5267 -17324 5295 -17290
rect 5339 -17324 5363 -17290
rect 5397 -17324 5436 -17290
rect 5866 -17324 5905 -17290
rect 5939 -17324 5963 -17290
rect 6007 -17324 6035 -17290
rect 6075 -17324 6107 -17290
rect 6143 -17324 6177 -17290
rect 6213 -17324 6245 -17290
rect 6285 -17324 6313 -17290
rect 6357 -17324 6381 -17290
rect 6415 -17324 6454 -17290
rect 6884 -17324 6923 -17290
rect 6957 -17324 6981 -17290
rect 7025 -17324 7053 -17290
rect 7093 -17324 7125 -17290
rect 7161 -17324 7195 -17290
rect 7231 -17324 7263 -17290
rect 7303 -17324 7331 -17290
rect 7375 -17324 7399 -17290
rect 7433 -17324 7472 -17290
rect 7902 -17324 7941 -17290
rect 7975 -17324 7999 -17290
rect 8043 -17324 8071 -17290
rect 8111 -17324 8143 -17290
rect 8179 -17324 8213 -17290
rect 8249 -17324 8281 -17290
rect 8321 -17324 8349 -17290
rect 8393 -17324 8417 -17290
rect 8451 -17324 8490 -17290
rect 8920 -17324 8959 -17290
rect 8993 -17324 9017 -17290
rect 9061 -17324 9089 -17290
rect 9129 -17324 9161 -17290
rect 9197 -17324 9231 -17290
rect 9267 -17324 9299 -17290
rect 9339 -17324 9367 -17290
rect 9411 -17324 9435 -17290
rect 9469 -17324 9508 -17290
rect 9938 -17324 9977 -17290
rect 10011 -17324 10035 -17290
rect 10079 -17324 10107 -17290
rect 10147 -17324 10179 -17290
rect 10215 -17324 10249 -17290
rect 10285 -17324 10317 -17290
rect 10357 -17324 10385 -17290
rect 10429 -17324 10453 -17290
rect 10487 -17324 10526 -17290
rect 10956 -17324 10995 -17290
rect 11029 -17324 11053 -17290
rect 11097 -17324 11125 -17290
rect 11165 -17324 11197 -17290
rect 11233 -17324 11267 -17290
rect 11303 -17324 11335 -17290
rect 11375 -17324 11403 -17290
rect 11447 -17324 11471 -17290
rect 11505 -17324 11544 -17290
rect 11974 -17324 12013 -17290
rect 12047 -17324 12071 -17290
rect 12115 -17324 12143 -17290
rect 12183 -17324 12215 -17290
rect 12251 -17324 12285 -17290
rect 12321 -17324 12353 -17290
rect 12393 -17324 12421 -17290
rect 12465 -17324 12489 -17290
rect 12523 -17324 12562 -17290
rect 12992 -17324 13031 -17290
rect 13065 -17324 13089 -17290
rect 13133 -17324 13161 -17290
rect 13201 -17324 13233 -17290
rect 13269 -17324 13303 -17290
rect 13339 -17324 13371 -17290
rect 13411 -17324 13439 -17290
rect 13483 -17324 13507 -17290
rect 13541 -17324 13580 -17290
rect 14010 -17324 14049 -17290
rect 14083 -17324 14107 -17290
rect 14151 -17324 14179 -17290
rect 14219 -17324 14251 -17290
rect 14287 -17324 14321 -17290
rect 14357 -17324 14389 -17290
rect 14429 -17324 14457 -17290
rect 14501 -17324 14525 -17290
rect 14559 -17324 14598 -17290
rect 15028 -17324 15067 -17290
rect 15101 -17324 15125 -17290
rect 15169 -17324 15197 -17290
rect 15237 -17324 15269 -17290
rect 15305 -17324 15339 -17290
rect 15375 -17324 15407 -17290
rect 15447 -17324 15475 -17290
rect 15519 -17324 15543 -17290
rect 15577 -17324 15616 -17290
rect 16046 -17324 16085 -17290
rect 16119 -17324 16143 -17290
rect 16187 -17324 16215 -17290
rect 16255 -17324 16287 -17290
rect 16323 -17324 16357 -17290
rect 16393 -17324 16425 -17290
rect 16465 -17324 16493 -17290
rect 16537 -17324 16561 -17290
rect 16595 -17324 16634 -17290
rect 17064 -17324 17103 -17290
rect 17137 -17324 17161 -17290
rect 17205 -17324 17233 -17290
rect 17273 -17324 17305 -17290
rect 17341 -17324 17375 -17290
rect 17411 -17324 17443 -17290
rect 17483 -17324 17511 -17290
rect 17555 -17324 17579 -17290
rect 17613 -17324 17652 -17290
rect 18082 -17324 18121 -17290
rect 18155 -17324 18179 -17290
rect 18223 -17324 18251 -17290
rect 18291 -17324 18323 -17290
rect 18359 -17324 18393 -17290
rect 18429 -17324 18461 -17290
rect 18501 -17324 18529 -17290
rect 18573 -17324 18597 -17290
rect 18631 -17324 18670 -17290
rect 19100 -17324 19139 -17290
rect 19173 -17324 19197 -17290
rect 19241 -17324 19269 -17290
rect 19309 -17324 19341 -17290
rect 19377 -17324 19411 -17290
rect 19447 -17324 19479 -17290
rect 19519 -17324 19547 -17290
rect 19591 -17324 19615 -17290
rect 19649 -17324 19688 -17290
rect 20118 -17324 20157 -17290
rect 20191 -17324 20215 -17290
rect 20259 -17324 20287 -17290
rect 20327 -17324 20359 -17290
rect 20395 -17324 20429 -17290
rect 20465 -17324 20497 -17290
rect 20537 -17324 20565 -17290
rect 20609 -17324 20633 -17290
rect 20667 -17324 20706 -17290
rect 21136 -17324 21175 -17290
rect 21209 -17324 21233 -17290
rect 21277 -17324 21305 -17290
rect 21345 -17324 21379 -17290
rect 21413 -17324 21447 -17290
rect 21481 -17324 21515 -17290
rect 21555 -17324 21583 -17290
rect 21627 -17324 21651 -17290
rect 21685 -17324 21724 -17290
rect 22154 -17324 22193 -17290
rect 22227 -17324 22251 -17290
rect 22295 -17324 22323 -17290
rect 22363 -17324 22395 -17290
rect 22431 -17324 22465 -17290
rect 22501 -17324 22533 -17290
rect 22573 -17324 22601 -17290
rect 22645 -17324 22669 -17290
rect 22703 -17324 22742 -17290
rect 24822 -17313 24855 -17275
rect 24889 -17313 24922 -17275
rect -12322 -17381 -12289 -17347
rect -12255 -17381 -12222 -17347
rect 24822 -17347 24922 -17313
rect -12322 -17415 -12222 -17381
rect -8952 -17382 -8913 -17348
rect -8879 -17382 -8855 -17348
rect -8811 -17382 -8783 -17348
rect -8743 -17382 -8711 -17348
rect -8675 -17382 -8641 -17348
rect -8605 -17382 -8573 -17348
rect -8533 -17382 -8505 -17348
rect -8461 -17382 -8437 -17348
rect -8403 -17382 -8364 -17348
rect -7934 -17382 -7895 -17348
rect -7861 -17382 -7837 -17348
rect -7793 -17382 -7765 -17348
rect -7725 -17382 -7693 -17348
rect -7657 -17382 -7623 -17348
rect -7587 -17382 -7555 -17348
rect -7515 -17382 -7487 -17348
rect -7443 -17382 -7419 -17348
rect -7385 -17382 -7346 -17348
rect -6916 -17382 -6877 -17348
rect -6843 -17382 -6819 -17348
rect -6775 -17382 -6747 -17348
rect -6707 -17382 -6675 -17348
rect -6639 -17382 -6605 -17348
rect -6569 -17382 -6537 -17348
rect -6497 -17382 -6469 -17348
rect -6425 -17382 -6401 -17348
rect -6367 -17382 -6328 -17348
rect -5898 -17382 -5859 -17348
rect -5825 -17382 -5801 -17348
rect -5757 -17382 -5729 -17348
rect -5689 -17382 -5657 -17348
rect -5621 -17382 -5587 -17348
rect -5551 -17382 -5519 -17348
rect -5479 -17382 -5451 -17348
rect -5407 -17382 -5383 -17348
rect -5349 -17382 -5310 -17348
rect -4880 -17382 -4841 -17348
rect -4807 -17382 -4783 -17348
rect -4739 -17382 -4711 -17348
rect -4671 -17382 -4639 -17348
rect -4603 -17382 -4569 -17348
rect -4533 -17382 -4501 -17348
rect -4461 -17382 -4433 -17348
rect -4389 -17382 -4365 -17348
rect -4331 -17382 -4292 -17348
rect -3862 -17382 -3823 -17348
rect -3789 -17382 -3765 -17348
rect -3721 -17382 -3693 -17348
rect -3653 -17382 -3621 -17348
rect -3585 -17382 -3551 -17348
rect -3515 -17382 -3483 -17348
rect -3443 -17382 -3415 -17348
rect -3371 -17382 -3347 -17348
rect -3313 -17382 -3274 -17348
rect -2844 -17382 -2805 -17348
rect -2771 -17382 -2747 -17348
rect -2703 -17382 -2675 -17348
rect -2635 -17382 -2603 -17348
rect -2567 -17382 -2533 -17348
rect -2497 -17382 -2465 -17348
rect -2425 -17382 -2397 -17348
rect -2353 -17382 -2329 -17348
rect -2295 -17382 -2256 -17348
rect -1826 -17382 -1787 -17348
rect -1753 -17382 -1729 -17348
rect -1685 -17382 -1657 -17348
rect -1617 -17382 -1585 -17348
rect -1549 -17382 -1515 -17348
rect -1479 -17382 -1447 -17348
rect -1407 -17382 -1379 -17348
rect -1335 -17382 -1311 -17348
rect -1277 -17382 -1238 -17348
rect -808 -17382 -769 -17348
rect -735 -17382 -711 -17348
rect -667 -17382 -639 -17348
rect -599 -17382 -567 -17348
rect -531 -17382 -497 -17348
rect -461 -17382 -429 -17348
rect -389 -17382 -361 -17348
rect -317 -17382 -293 -17348
rect -259 -17382 -220 -17348
rect 24822 -17381 24855 -17347
rect 24889 -17381 24922 -17347
rect -12322 -17453 -12289 -17415
rect -12255 -17453 -12222 -17415
rect 24822 -17415 24922 -17381
rect -12322 -17483 -12222 -17453
rect -12322 -17525 -12289 -17483
rect -12255 -17525 -12222 -17483
rect -12322 -17551 -12222 -17525
rect -12322 -17597 -12289 -17551
rect -12255 -17597 -12222 -17551
rect -12322 -17619 -12222 -17597
rect -12322 -17669 -12289 -17619
rect -12255 -17669 -12222 -17619
rect -12322 -17687 -12222 -17669
rect -12322 -17741 -12289 -17687
rect -12255 -17741 -12222 -17687
rect -12322 -17755 -12222 -17741
rect -12322 -17813 -12289 -17755
rect -12255 -17813 -12222 -17755
rect -12322 -17823 -12222 -17813
rect -12322 -17885 -12289 -17823
rect -12255 -17885 -12222 -17823
rect -12322 -17891 -12222 -17885
rect -12322 -17957 -12289 -17891
rect -12255 -17957 -12222 -17891
rect -12322 -17959 -12222 -17957
rect -12322 -17993 -12289 -17959
rect -12255 -17993 -12222 -17959
rect -12322 -17995 -12222 -17993
rect -12322 -18061 -12289 -17995
rect -12255 -18061 -12222 -17995
rect -9184 -17451 -9150 -17416
rect -9184 -17523 -9150 -17499
rect -9184 -17595 -9150 -17567
rect -9184 -17667 -9150 -17635
rect -9184 -17737 -9150 -17703
rect -9184 -17805 -9150 -17773
rect -9184 -17873 -9150 -17845
rect -9184 -17941 -9150 -17917
rect -9184 -18024 -9150 -17989
rect -8166 -17451 -8132 -17416
rect -8166 -17523 -8132 -17499
rect -8166 -17595 -8132 -17567
rect -8166 -17667 -8132 -17635
rect -8166 -17737 -8132 -17703
rect -8166 -17805 -8132 -17773
rect -8166 -17873 -8132 -17845
rect -8166 -17941 -8132 -17917
rect -8166 -18024 -8132 -17989
rect -7148 -17451 -7114 -17416
rect -7148 -17523 -7114 -17499
rect -7148 -17595 -7114 -17567
rect -7148 -17667 -7114 -17635
rect -7148 -17737 -7114 -17703
rect -7148 -17805 -7114 -17773
rect -7148 -17873 -7114 -17845
rect -7148 -17941 -7114 -17917
rect -7148 -18024 -7114 -17989
rect -6130 -17451 -6096 -17416
rect -6130 -17523 -6096 -17499
rect -6130 -17595 -6096 -17567
rect -6130 -17667 -6096 -17635
rect -6130 -17737 -6096 -17703
rect -6130 -17805 -6096 -17773
rect -6130 -17873 -6096 -17845
rect -6130 -17941 -6096 -17917
rect -6130 -18024 -6096 -17989
rect -5112 -17451 -5078 -17416
rect -5112 -17523 -5078 -17499
rect -5112 -17595 -5078 -17567
rect -5112 -17667 -5078 -17635
rect -5112 -17737 -5078 -17703
rect -5112 -17805 -5078 -17773
rect -5112 -17873 -5078 -17845
rect -5112 -17941 -5078 -17917
rect -5112 -18024 -5078 -17989
rect -4094 -17451 -4060 -17416
rect -4094 -17523 -4060 -17499
rect -4094 -17595 -4060 -17567
rect -4094 -17667 -4060 -17635
rect -4094 -17737 -4060 -17703
rect -4094 -17805 -4060 -17773
rect -4094 -17873 -4060 -17845
rect -4094 -17941 -4060 -17917
rect -4094 -18024 -4060 -17989
rect -3076 -17451 -3042 -17416
rect -3076 -17523 -3042 -17499
rect -3076 -17595 -3042 -17567
rect -3076 -17667 -3042 -17635
rect -3076 -17737 -3042 -17703
rect -3076 -17805 -3042 -17773
rect -3076 -17873 -3042 -17845
rect -3076 -17941 -3042 -17917
rect -3076 -18024 -3042 -17989
rect -2058 -17451 -2024 -17416
rect -2058 -17523 -2024 -17499
rect -2058 -17595 -2024 -17567
rect -2058 -17667 -2024 -17635
rect -2058 -17737 -2024 -17703
rect -2058 -17805 -2024 -17773
rect -2058 -17873 -2024 -17845
rect -2058 -17941 -2024 -17917
rect -2058 -18024 -2024 -17989
rect -1040 -17451 -1006 -17416
rect -1040 -17523 -1006 -17499
rect -1040 -17595 -1006 -17567
rect -1040 -17667 -1006 -17635
rect -1040 -17737 -1006 -17703
rect -1040 -17805 -1006 -17773
rect -1040 -17873 -1006 -17845
rect -1040 -17941 -1006 -17917
rect -1040 -18024 -1006 -17989
rect -22 -17451 12 -17416
rect -22 -17523 12 -17499
rect -22 -17595 12 -17567
rect -22 -17667 12 -17635
rect -22 -17737 12 -17703
rect -22 -17805 12 -17773
rect 24822 -17453 24855 -17415
rect 24889 -17453 24922 -17415
rect 24822 -17483 24922 -17453
rect 24822 -17525 24855 -17483
rect 24889 -17525 24922 -17483
rect 24822 -17551 24922 -17525
rect 24822 -17597 24855 -17551
rect 24889 -17597 24922 -17551
rect 24822 -17619 24922 -17597
rect 24822 -17669 24855 -17619
rect 24889 -17669 24922 -17619
rect 24822 -17687 24922 -17669
rect 24822 -17741 24855 -17687
rect 24889 -17741 24922 -17687
rect 24822 -17755 24922 -17741
rect -22 -17873 12 -17845
rect 2812 -17846 2851 -17812
rect 2885 -17846 2909 -17812
rect 2953 -17846 2981 -17812
rect 3021 -17846 3053 -17812
rect 3089 -17846 3123 -17812
rect 3159 -17846 3191 -17812
rect 3231 -17846 3259 -17812
rect 3303 -17846 3327 -17812
rect 3361 -17846 3400 -17812
rect 3830 -17846 3869 -17812
rect 3903 -17846 3927 -17812
rect 3971 -17846 3999 -17812
rect 4039 -17846 4071 -17812
rect 4107 -17846 4141 -17812
rect 4177 -17846 4209 -17812
rect 4249 -17846 4277 -17812
rect 4321 -17846 4345 -17812
rect 4379 -17846 4418 -17812
rect 4848 -17846 4887 -17812
rect 4921 -17846 4945 -17812
rect 4989 -17846 5017 -17812
rect 5057 -17846 5089 -17812
rect 5125 -17846 5159 -17812
rect 5195 -17846 5227 -17812
rect 5267 -17846 5295 -17812
rect 5339 -17846 5363 -17812
rect 5397 -17846 5436 -17812
rect 5866 -17846 5905 -17812
rect 5939 -17846 5963 -17812
rect 6007 -17846 6035 -17812
rect 6075 -17846 6107 -17812
rect 6143 -17846 6177 -17812
rect 6213 -17846 6245 -17812
rect 6285 -17846 6313 -17812
rect 6357 -17846 6381 -17812
rect 6415 -17846 6454 -17812
rect 6884 -17846 6923 -17812
rect 6957 -17846 6981 -17812
rect 7025 -17846 7053 -17812
rect 7093 -17846 7125 -17812
rect 7161 -17846 7195 -17812
rect 7231 -17846 7263 -17812
rect 7303 -17846 7331 -17812
rect 7375 -17846 7399 -17812
rect 7433 -17846 7472 -17812
rect 7902 -17846 7941 -17812
rect 7975 -17846 7999 -17812
rect 8043 -17846 8071 -17812
rect 8111 -17846 8143 -17812
rect 8179 -17846 8213 -17812
rect 8249 -17846 8281 -17812
rect 8321 -17846 8349 -17812
rect 8393 -17846 8417 -17812
rect 8451 -17846 8490 -17812
rect 8920 -17846 8959 -17812
rect 8993 -17846 9017 -17812
rect 9061 -17846 9089 -17812
rect 9129 -17846 9161 -17812
rect 9197 -17846 9231 -17812
rect 9267 -17846 9299 -17812
rect 9339 -17846 9367 -17812
rect 9411 -17846 9435 -17812
rect 9469 -17846 9508 -17812
rect 9938 -17846 9977 -17812
rect 10011 -17846 10035 -17812
rect 10079 -17846 10107 -17812
rect 10147 -17846 10179 -17812
rect 10215 -17846 10249 -17812
rect 10285 -17846 10317 -17812
rect 10357 -17846 10385 -17812
rect 10429 -17846 10453 -17812
rect 10487 -17846 10526 -17812
rect 10956 -17846 10995 -17812
rect 11029 -17846 11053 -17812
rect 11097 -17846 11125 -17812
rect 11165 -17846 11197 -17812
rect 11233 -17846 11267 -17812
rect 11303 -17846 11335 -17812
rect 11375 -17846 11403 -17812
rect 11447 -17846 11471 -17812
rect 11505 -17846 11544 -17812
rect 11974 -17846 12013 -17812
rect 12047 -17846 12071 -17812
rect 12115 -17846 12143 -17812
rect 12183 -17846 12215 -17812
rect 12251 -17846 12285 -17812
rect 12321 -17846 12353 -17812
rect 12393 -17846 12421 -17812
rect 12465 -17846 12489 -17812
rect 12523 -17846 12562 -17812
rect 12992 -17846 13031 -17812
rect 13065 -17846 13089 -17812
rect 13133 -17846 13161 -17812
rect 13201 -17846 13233 -17812
rect 13269 -17846 13303 -17812
rect 13339 -17846 13371 -17812
rect 13411 -17846 13439 -17812
rect 13483 -17846 13507 -17812
rect 13541 -17846 13580 -17812
rect 14010 -17846 14049 -17812
rect 14083 -17846 14107 -17812
rect 14151 -17846 14179 -17812
rect 14219 -17846 14251 -17812
rect 14287 -17846 14321 -17812
rect 14357 -17846 14389 -17812
rect 14429 -17846 14457 -17812
rect 14501 -17846 14525 -17812
rect 14559 -17846 14598 -17812
rect 15028 -17846 15067 -17812
rect 15101 -17846 15125 -17812
rect 15169 -17846 15197 -17812
rect 15237 -17846 15269 -17812
rect 15305 -17846 15339 -17812
rect 15375 -17846 15407 -17812
rect 15447 -17846 15475 -17812
rect 15519 -17846 15543 -17812
rect 15577 -17846 15616 -17812
rect 16046 -17846 16085 -17812
rect 16119 -17846 16143 -17812
rect 16187 -17846 16215 -17812
rect 16255 -17846 16287 -17812
rect 16323 -17846 16357 -17812
rect 16393 -17846 16425 -17812
rect 16465 -17846 16493 -17812
rect 16537 -17846 16561 -17812
rect 16595 -17846 16634 -17812
rect 17064 -17846 17103 -17812
rect 17137 -17846 17161 -17812
rect 17205 -17846 17233 -17812
rect 17273 -17846 17305 -17812
rect 17341 -17846 17375 -17812
rect 17411 -17846 17443 -17812
rect 17483 -17846 17511 -17812
rect 17555 -17846 17579 -17812
rect 17613 -17846 17652 -17812
rect 18082 -17846 18121 -17812
rect 18155 -17846 18179 -17812
rect 18223 -17846 18251 -17812
rect 18291 -17846 18323 -17812
rect 18359 -17846 18393 -17812
rect 18429 -17846 18461 -17812
rect 18501 -17846 18529 -17812
rect 18573 -17846 18597 -17812
rect 18631 -17846 18670 -17812
rect 19100 -17846 19139 -17812
rect 19173 -17846 19197 -17812
rect 19241 -17846 19269 -17812
rect 19309 -17846 19341 -17812
rect 19377 -17846 19411 -17812
rect 19447 -17846 19479 -17812
rect 19519 -17846 19547 -17812
rect 19591 -17846 19615 -17812
rect 19649 -17846 19688 -17812
rect 20118 -17846 20157 -17812
rect 20191 -17846 20215 -17812
rect 20259 -17846 20287 -17812
rect 20327 -17846 20359 -17812
rect 20395 -17846 20429 -17812
rect 20465 -17846 20497 -17812
rect 20537 -17846 20565 -17812
rect 20609 -17846 20633 -17812
rect 20667 -17846 20706 -17812
rect 21136 -17846 21175 -17812
rect 21209 -17846 21233 -17812
rect 21277 -17846 21305 -17812
rect 21345 -17846 21377 -17812
rect 21413 -17846 21447 -17812
rect 21483 -17846 21515 -17812
rect 21555 -17846 21583 -17812
rect 21627 -17846 21651 -17812
rect 21685 -17846 21724 -17812
rect 22154 -17846 22193 -17812
rect 22227 -17846 22251 -17812
rect 22295 -17846 22323 -17812
rect 22363 -17846 22395 -17812
rect 22431 -17846 22465 -17812
rect 22501 -17846 22533 -17812
rect 22573 -17846 22601 -17812
rect 22645 -17846 22669 -17812
rect 22703 -17846 22742 -17812
rect 24822 -17813 24855 -17755
rect 24889 -17813 24922 -17755
rect 24822 -17823 24922 -17813
rect -22 -17941 12 -17917
rect -22 -18024 12 -17989
rect 2580 -17915 2614 -17880
rect 2580 -17987 2614 -17963
rect -8692 -18058 -8632 -18056
rect -7666 -18058 -7606 -18054
rect -6652 -18058 -6592 -18054
rect -5632 -18058 -5572 -18056
rect -4610 -18058 -4550 -18056
rect -2578 -18058 -2518 -18054
rect -1562 -18058 -1502 -18054
rect -542 -18058 -482 -18056
rect -12322 -18067 -12222 -18061
rect -12322 -18129 -12289 -18067
rect -12255 -18129 -12222 -18067
rect -8952 -18092 -8913 -18058
rect -8879 -18092 -8855 -18058
rect -8811 -18092 -8783 -18058
rect -8743 -18092 -8711 -18058
rect -8675 -18092 -8641 -18058
rect -8605 -18092 -8573 -18058
rect -8533 -18092 -8505 -18058
rect -8461 -18092 -8437 -18058
rect -8403 -18092 -8364 -18058
rect -7934 -18092 -7895 -18058
rect -7861 -18092 -7837 -18058
rect -7793 -18092 -7765 -18058
rect -7725 -18092 -7693 -18058
rect -7657 -18092 -7623 -18058
rect -7587 -18092 -7555 -18058
rect -7515 -18092 -7487 -18058
rect -7443 -18092 -7419 -18058
rect -7385 -18092 -7346 -18058
rect -6916 -18092 -6877 -18058
rect -6843 -18092 -6819 -18058
rect -6775 -18092 -6747 -18058
rect -6707 -18092 -6675 -18058
rect -6639 -18092 -6605 -18058
rect -6569 -18092 -6537 -18058
rect -6497 -18092 -6469 -18058
rect -6425 -18092 -6401 -18058
rect -6367 -18092 -6328 -18058
rect -5898 -18092 -5859 -18058
rect -5825 -18092 -5801 -18058
rect -5757 -18092 -5729 -18058
rect -5689 -18092 -5657 -18058
rect -5621 -18092 -5587 -18058
rect -5551 -18092 -5519 -18058
rect -5479 -18092 -5451 -18058
rect -5407 -18092 -5383 -18058
rect -5349 -18092 -5310 -18058
rect -4880 -18092 -4841 -18058
rect -4807 -18092 -4783 -18058
rect -4739 -18092 -4711 -18058
rect -4671 -18092 -4639 -18058
rect -4603 -18092 -4569 -18058
rect -4533 -18092 -4501 -18058
rect -4461 -18092 -4433 -18058
rect -4389 -18092 -4365 -18058
rect -4331 -18092 -4292 -18058
rect -3862 -18092 -3823 -18058
rect -3789 -18092 -3765 -18058
rect -3721 -18092 -3693 -18058
rect -3653 -18092 -3621 -18058
rect -3585 -18092 -3551 -18058
rect -3515 -18092 -3483 -18058
rect -3443 -18092 -3415 -18058
rect -3371 -18092 -3347 -18058
rect -3313 -18092 -3274 -18058
rect -2844 -18092 -2805 -18058
rect -2771 -18092 -2747 -18058
rect -2703 -18092 -2675 -18058
rect -2635 -18092 -2603 -18058
rect -2567 -18092 -2533 -18058
rect -2497 -18092 -2465 -18058
rect -2425 -18092 -2397 -18058
rect -2353 -18092 -2329 -18058
rect -2295 -18092 -2256 -18058
rect -1826 -18092 -1787 -18058
rect -1753 -18092 -1729 -18058
rect -1685 -18092 -1657 -18058
rect -1617 -18092 -1585 -18058
rect -1549 -18092 -1515 -18058
rect -1479 -18092 -1447 -18058
rect -1407 -18092 -1379 -18058
rect -1335 -18092 -1311 -18058
rect -1277 -18092 -1238 -18058
rect -808 -18092 -769 -18058
rect -735 -18092 -711 -18058
rect -667 -18092 -639 -18058
rect -599 -18092 -567 -18058
rect -531 -18092 -497 -18058
rect -461 -18092 -429 -18058
rect -389 -18092 -361 -18058
rect -317 -18092 -293 -18058
rect -259 -18092 -220 -18058
rect 2580 -18059 2614 -18031
rect -12322 -18139 -12222 -18129
rect -12322 -18197 -12289 -18139
rect -12255 -18197 -12222 -18139
rect 2580 -18131 2614 -18099
rect -12322 -18211 -12222 -18197
rect -8952 -18200 -8913 -18166
rect -8879 -18200 -8855 -18166
rect -8811 -18200 -8783 -18166
rect -8743 -18200 -8711 -18166
rect -8675 -18200 -8641 -18166
rect -8605 -18200 -8573 -18166
rect -8533 -18200 -8505 -18166
rect -8461 -18200 -8437 -18166
rect -8403 -18200 -8364 -18166
rect -7934 -18200 -7895 -18166
rect -7861 -18200 -7837 -18166
rect -7793 -18200 -7765 -18166
rect -7725 -18200 -7693 -18166
rect -7657 -18200 -7623 -18166
rect -7587 -18200 -7555 -18166
rect -7515 -18200 -7487 -18166
rect -7443 -18200 -7419 -18166
rect -7385 -18200 -7346 -18166
rect -6916 -18200 -6877 -18166
rect -6843 -18200 -6819 -18166
rect -6775 -18200 -6747 -18166
rect -6707 -18200 -6675 -18166
rect -6639 -18200 -6605 -18166
rect -6569 -18200 -6537 -18166
rect -6497 -18200 -6469 -18166
rect -6425 -18200 -6401 -18166
rect -6367 -18200 -6328 -18166
rect -5898 -18200 -5859 -18166
rect -5825 -18200 -5801 -18166
rect -5757 -18200 -5729 -18166
rect -5689 -18200 -5657 -18166
rect -5621 -18200 -5587 -18166
rect -5551 -18200 -5519 -18166
rect -5479 -18200 -5451 -18166
rect -5407 -18200 -5383 -18166
rect -5349 -18200 -5310 -18166
rect -4880 -18200 -4841 -18166
rect -4807 -18200 -4783 -18166
rect -4739 -18200 -4711 -18166
rect -4671 -18200 -4639 -18166
rect -4603 -18200 -4569 -18166
rect -4533 -18200 -4501 -18166
rect -4461 -18200 -4433 -18166
rect -4389 -18200 -4365 -18166
rect -4331 -18200 -4292 -18166
rect -3862 -18200 -3823 -18166
rect -3789 -18200 -3765 -18166
rect -3721 -18200 -3693 -18166
rect -3653 -18200 -3621 -18166
rect -3585 -18200 -3551 -18166
rect -3515 -18200 -3483 -18166
rect -3443 -18200 -3415 -18166
rect -3371 -18200 -3347 -18166
rect -3313 -18200 -3274 -18166
rect -2844 -18200 -2805 -18166
rect -2771 -18200 -2747 -18166
rect -2703 -18200 -2675 -18166
rect -2635 -18200 -2603 -18166
rect -2567 -18200 -2533 -18166
rect -2497 -18200 -2465 -18166
rect -2425 -18200 -2397 -18166
rect -2353 -18200 -2329 -18166
rect -2295 -18200 -2256 -18166
rect -1826 -18200 -1787 -18166
rect -1753 -18200 -1729 -18166
rect -1685 -18200 -1657 -18166
rect -1617 -18200 -1585 -18166
rect -1549 -18200 -1515 -18166
rect -1479 -18200 -1447 -18166
rect -1407 -18200 -1379 -18166
rect -1335 -18200 -1311 -18166
rect -1277 -18200 -1238 -18166
rect -808 -18200 -769 -18166
rect -735 -18200 -711 -18166
rect -667 -18200 -639 -18166
rect -599 -18200 -567 -18166
rect -531 -18200 -497 -18166
rect -461 -18200 -429 -18166
rect -389 -18200 -361 -18166
rect -317 -18200 -293 -18166
rect -259 -18200 -220 -18166
rect -12322 -18265 -12289 -18211
rect -12255 -18265 -12222 -18211
rect 2580 -18201 2614 -18167
rect -12322 -18283 -12222 -18265
rect -12322 -18333 -12289 -18283
rect -12255 -18333 -12222 -18283
rect -12322 -18355 -12222 -18333
rect -12322 -18401 -12289 -18355
rect -12255 -18401 -12222 -18355
rect -12322 -18427 -12222 -18401
rect -12322 -18469 -12289 -18427
rect -12255 -18469 -12222 -18427
rect -12322 -18499 -12222 -18469
rect -12322 -18537 -12289 -18499
rect -12255 -18537 -12222 -18499
rect -12322 -18571 -12222 -18537
rect -12322 -18605 -12289 -18571
rect -12255 -18605 -12222 -18571
rect -12322 -18639 -12222 -18605
rect -12322 -18677 -12289 -18639
rect -12255 -18677 -12222 -18639
rect -12322 -18707 -12222 -18677
rect -12322 -18749 -12289 -18707
rect -12255 -18749 -12222 -18707
rect -12322 -18775 -12222 -18749
rect -12322 -18821 -12289 -18775
rect -12255 -18821 -12222 -18775
rect -12322 -18843 -12222 -18821
rect -9184 -18269 -9150 -18234
rect -9184 -18341 -9150 -18317
rect -9184 -18413 -9150 -18385
rect -9184 -18485 -9150 -18453
rect -9184 -18555 -9150 -18521
rect -9184 -18623 -9150 -18591
rect -9184 -18691 -9150 -18663
rect -9184 -18759 -9150 -18735
rect -9184 -18842 -9150 -18807
rect -8166 -18269 -8132 -18234
rect -8166 -18341 -8132 -18317
rect -8166 -18413 -8132 -18385
rect -8166 -18485 -8132 -18453
rect -8166 -18555 -8132 -18521
rect -8166 -18623 -8132 -18591
rect -8166 -18691 -8132 -18663
rect -8166 -18759 -8132 -18735
rect -8166 -18842 -8132 -18807
rect -7148 -18269 -7114 -18234
rect -7148 -18341 -7114 -18317
rect -7148 -18413 -7114 -18385
rect -7148 -18485 -7114 -18453
rect -7148 -18555 -7114 -18521
rect -7148 -18623 -7114 -18591
rect -7148 -18691 -7114 -18663
rect -7148 -18759 -7114 -18735
rect -7148 -18842 -7114 -18807
rect -6130 -18269 -6096 -18234
rect -6130 -18341 -6096 -18317
rect -6130 -18413 -6096 -18385
rect -6130 -18485 -6096 -18453
rect -6130 -18555 -6096 -18521
rect -6130 -18623 -6096 -18591
rect -6130 -18691 -6096 -18663
rect -6130 -18759 -6096 -18735
rect -6130 -18842 -6096 -18807
rect -5112 -18269 -5078 -18234
rect -5112 -18341 -5078 -18317
rect -5112 -18413 -5078 -18385
rect -5112 -18485 -5078 -18453
rect -5112 -18555 -5078 -18521
rect -5112 -18623 -5078 -18591
rect -5112 -18691 -5078 -18663
rect -5112 -18759 -5078 -18735
rect -5112 -18842 -5078 -18807
rect -4094 -18269 -4060 -18234
rect -4094 -18341 -4060 -18317
rect -4094 -18413 -4060 -18385
rect -4094 -18485 -4060 -18453
rect -4094 -18555 -4060 -18521
rect -4094 -18623 -4060 -18591
rect -4094 -18691 -4060 -18663
rect -4094 -18759 -4060 -18735
rect -4094 -18842 -4060 -18807
rect -3076 -18269 -3042 -18234
rect -3076 -18341 -3042 -18317
rect -3076 -18413 -3042 -18385
rect -3076 -18485 -3042 -18453
rect -3076 -18555 -3042 -18521
rect -3076 -18623 -3042 -18591
rect -3076 -18691 -3042 -18663
rect -3076 -18759 -3042 -18735
rect -3076 -18842 -3042 -18807
rect -2058 -18269 -2024 -18234
rect -2058 -18341 -2024 -18317
rect -2058 -18413 -2024 -18385
rect -2058 -18485 -2024 -18453
rect -2058 -18555 -2024 -18521
rect -2058 -18623 -2024 -18591
rect -2058 -18691 -2024 -18663
rect -2058 -18759 -2024 -18735
rect -2058 -18842 -2024 -18807
rect -1040 -18269 -1006 -18234
rect -1040 -18341 -1006 -18317
rect -1040 -18413 -1006 -18385
rect -1040 -18485 -1006 -18453
rect -1040 -18555 -1006 -18521
rect -1040 -18623 -1006 -18591
rect -1040 -18691 -1006 -18663
rect -1040 -18759 -1006 -18735
rect -1040 -18842 -1006 -18807
rect -22 -18269 12 -18234
rect -22 -18341 12 -18317
rect -22 -18413 12 -18385
rect -22 -18485 12 -18453
rect 2580 -18269 2614 -18237
rect 2580 -18337 2614 -18309
rect 2580 -18405 2614 -18381
rect 2580 -18488 2614 -18453
rect 3598 -17915 3632 -17880
rect 3598 -17987 3632 -17963
rect 3598 -18059 3632 -18031
rect 3598 -18131 3632 -18099
rect 3598 -18201 3632 -18167
rect 3598 -18269 3632 -18237
rect 3598 -18337 3632 -18309
rect 3598 -18405 3632 -18381
rect 3598 -18488 3632 -18453
rect 4616 -17915 4650 -17880
rect 4616 -17987 4650 -17963
rect 4616 -18059 4650 -18031
rect 4616 -18131 4650 -18099
rect 4616 -18201 4650 -18167
rect 4616 -18269 4650 -18237
rect 4616 -18337 4650 -18309
rect 4616 -18405 4650 -18381
rect 4616 -18488 4650 -18453
rect 5634 -17915 5668 -17880
rect 5634 -17987 5668 -17963
rect 5634 -18059 5668 -18031
rect 5634 -18131 5668 -18099
rect 5634 -18201 5668 -18167
rect 5634 -18269 5668 -18237
rect 5634 -18337 5668 -18309
rect 5634 -18405 5668 -18381
rect 5634 -18488 5668 -18453
rect 6652 -17915 6686 -17880
rect 6652 -17987 6686 -17963
rect 6652 -18059 6686 -18031
rect 6652 -18131 6686 -18099
rect 6652 -18201 6686 -18167
rect 6652 -18269 6686 -18237
rect 6652 -18337 6686 -18309
rect 6652 -18405 6686 -18381
rect 6652 -18488 6686 -18453
rect 7670 -17915 7704 -17880
rect 7670 -17987 7704 -17963
rect 7670 -18059 7704 -18031
rect 7670 -18131 7704 -18099
rect 7670 -18201 7704 -18167
rect 7670 -18269 7704 -18237
rect 7670 -18337 7704 -18309
rect 7670 -18405 7704 -18381
rect 7670 -18488 7704 -18453
rect 8688 -17915 8722 -17880
rect 8688 -17987 8722 -17963
rect 8688 -18059 8722 -18031
rect 8688 -18131 8722 -18099
rect 8688 -18201 8722 -18167
rect 8688 -18269 8722 -18237
rect 8688 -18337 8722 -18309
rect 8688 -18405 8722 -18381
rect 8688 -18488 8722 -18453
rect 9706 -17915 9740 -17880
rect 9706 -17987 9740 -17963
rect 9706 -18059 9740 -18031
rect 9706 -18131 9740 -18099
rect 9706 -18201 9740 -18167
rect 9706 -18269 9740 -18237
rect 9706 -18337 9740 -18309
rect 9706 -18405 9740 -18381
rect 9706 -18488 9740 -18453
rect 10724 -17915 10758 -17880
rect 10724 -17987 10758 -17963
rect 10724 -18059 10758 -18031
rect 10724 -18131 10758 -18099
rect 10724 -18201 10758 -18167
rect 10724 -18269 10758 -18237
rect 10724 -18337 10758 -18309
rect 10724 -18405 10758 -18381
rect 10724 -18488 10758 -18453
rect 11742 -17915 11776 -17880
rect 11742 -17987 11776 -17963
rect 11742 -18059 11776 -18031
rect 11742 -18131 11776 -18099
rect 11742 -18201 11776 -18167
rect 11742 -18269 11776 -18237
rect 11742 -18337 11776 -18309
rect 11742 -18405 11776 -18381
rect 11742 -18488 11776 -18453
rect 12760 -17915 12794 -17880
rect 12760 -17987 12794 -17963
rect 12760 -18059 12794 -18031
rect 12760 -18131 12794 -18099
rect 12760 -18201 12794 -18167
rect 12760 -18269 12794 -18237
rect 12760 -18337 12794 -18309
rect 12760 -18405 12794 -18381
rect 12760 -18488 12794 -18453
rect 13778 -17915 13812 -17880
rect 13778 -17987 13812 -17963
rect 13778 -18059 13812 -18031
rect 13778 -18131 13812 -18099
rect 13778 -18201 13812 -18167
rect 13778 -18269 13812 -18237
rect 13778 -18337 13812 -18309
rect 13778 -18405 13812 -18381
rect 13778 -18488 13812 -18453
rect 14796 -17915 14830 -17880
rect 14796 -17987 14830 -17963
rect 14796 -18059 14830 -18031
rect 14796 -18131 14830 -18099
rect 14796 -18201 14830 -18167
rect 14796 -18269 14830 -18237
rect 14796 -18337 14830 -18309
rect 14796 -18405 14830 -18381
rect 14796 -18488 14830 -18453
rect 15814 -17915 15848 -17880
rect 15814 -17987 15848 -17963
rect 15814 -18059 15848 -18031
rect 15814 -18131 15848 -18099
rect 15814 -18201 15848 -18167
rect 15814 -18269 15848 -18237
rect 15814 -18337 15848 -18309
rect 15814 -18405 15848 -18381
rect 15814 -18488 15848 -18453
rect 16832 -17915 16866 -17880
rect 16832 -17987 16866 -17963
rect 16832 -18059 16866 -18031
rect 16832 -18131 16866 -18099
rect 16832 -18201 16866 -18167
rect 16832 -18269 16866 -18237
rect 16832 -18337 16866 -18309
rect 16832 -18405 16866 -18381
rect 16832 -18488 16866 -18453
rect 17850 -17915 17884 -17880
rect 17850 -17987 17884 -17963
rect 17850 -18059 17884 -18031
rect 17850 -18131 17884 -18099
rect 17850 -18201 17884 -18167
rect 17850 -18269 17884 -18237
rect 17850 -18337 17884 -18309
rect 17850 -18405 17884 -18381
rect 17850 -18488 17884 -18453
rect 18868 -17915 18902 -17880
rect 18868 -17987 18902 -17963
rect 18868 -18059 18902 -18031
rect 18868 -18131 18902 -18099
rect 18868 -18201 18902 -18167
rect 18868 -18269 18902 -18237
rect 18868 -18337 18902 -18309
rect 18868 -18405 18902 -18381
rect 18868 -18488 18902 -18453
rect 19886 -17915 19920 -17880
rect 19886 -17987 19920 -17963
rect 19886 -18059 19920 -18031
rect 19886 -18131 19920 -18099
rect 19886 -18201 19920 -18167
rect 19886 -18269 19920 -18237
rect 19886 -18337 19920 -18309
rect 19886 -18405 19920 -18381
rect 19886 -18488 19920 -18453
rect 20904 -17915 20938 -17880
rect 20904 -17987 20938 -17963
rect 20904 -18059 20938 -18031
rect 20904 -18131 20938 -18099
rect 20904 -18201 20938 -18167
rect 20904 -18269 20938 -18237
rect 20904 -18337 20938 -18309
rect 20904 -18405 20938 -18381
rect 20904 -18488 20938 -18453
rect 21922 -17915 21956 -17880
rect 21922 -17987 21956 -17963
rect 21922 -18059 21956 -18031
rect 21922 -18131 21956 -18099
rect 21922 -18201 21956 -18167
rect 21922 -18269 21956 -18237
rect 21922 -18337 21956 -18309
rect 21922 -18405 21956 -18381
rect 21922 -18488 21956 -18453
rect 22940 -17915 22974 -17880
rect 22940 -17987 22974 -17963
rect 22940 -18059 22974 -18031
rect 22940 -18131 22974 -18099
rect 22940 -18201 22974 -18167
rect 22940 -18269 22974 -18237
rect 22940 -18337 22974 -18309
rect 22940 -18405 22974 -18381
rect 22940 -18488 22974 -18453
rect 24822 -17885 24855 -17823
rect 24889 -17885 24922 -17823
rect 24822 -17891 24922 -17885
rect 24822 -17957 24855 -17891
rect 24889 -17957 24922 -17891
rect 24822 -17959 24922 -17957
rect 24822 -17993 24855 -17959
rect 24889 -17993 24922 -17959
rect 24822 -17995 24922 -17993
rect 24822 -18061 24855 -17995
rect 24889 -18061 24922 -17995
rect 24822 -18067 24922 -18061
rect 24822 -18129 24855 -18067
rect 24889 -18129 24922 -18067
rect 24822 -18139 24922 -18129
rect 24822 -18197 24855 -18139
rect 24889 -18197 24922 -18139
rect 24822 -18211 24922 -18197
rect 24822 -18265 24855 -18211
rect 24889 -18265 24922 -18211
rect 24822 -18283 24922 -18265
rect 24822 -18333 24855 -18283
rect 24889 -18333 24922 -18283
rect 24822 -18355 24922 -18333
rect 24822 -18401 24855 -18355
rect 24889 -18401 24922 -18355
rect 24822 -18427 24922 -18401
rect 24822 -18469 24855 -18427
rect 24889 -18469 24922 -18427
rect 24822 -18499 24922 -18469
rect -22 -18555 12 -18521
rect 11230 -18522 11290 -18520
rect 13274 -18522 13334 -18518
rect 21408 -18522 21468 -18520
rect 2812 -18556 2851 -18522
rect 2885 -18556 2909 -18522
rect 2953 -18556 2981 -18522
rect 3021 -18556 3053 -18522
rect 3089 -18556 3123 -18522
rect 3159 -18556 3191 -18522
rect 3231 -18556 3259 -18522
rect 3303 -18556 3327 -18522
rect 3361 -18556 3400 -18522
rect 3830 -18556 3869 -18522
rect 3903 -18556 3927 -18522
rect 3971 -18556 3999 -18522
rect 4039 -18556 4071 -18522
rect 4107 -18556 4141 -18522
rect 4177 -18556 4209 -18522
rect 4249 -18556 4277 -18522
rect 4321 -18556 4345 -18522
rect 4379 -18556 4418 -18522
rect 4848 -18556 4887 -18522
rect 4921 -18556 4945 -18522
rect 4989 -18556 5017 -18522
rect 5057 -18556 5089 -18522
rect 5125 -18556 5159 -18522
rect 5195 -18556 5227 -18522
rect 5267 -18556 5295 -18522
rect 5339 -18556 5363 -18522
rect 5397 -18556 5436 -18522
rect 5866 -18556 5905 -18522
rect 5939 -18556 5963 -18522
rect 6007 -18556 6035 -18522
rect 6075 -18556 6107 -18522
rect 6143 -18556 6177 -18522
rect 6213 -18556 6245 -18522
rect 6285 -18556 6313 -18522
rect 6357 -18556 6381 -18522
rect 6415 -18556 6454 -18522
rect 6884 -18556 6923 -18522
rect 6957 -18556 6981 -18522
rect 7025 -18556 7053 -18522
rect 7093 -18556 7125 -18522
rect 7161 -18556 7195 -18522
rect 7231 -18556 7263 -18522
rect 7303 -18556 7331 -18522
rect 7375 -18556 7399 -18522
rect 7433 -18556 7472 -18522
rect 7902 -18556 7941 -18522
rect 7975 -18556 7999 -18522
rect 8043 -18556 8071 -18522
rect 8111 -18556 8143 -18522
rect 8179 -18556 8213 -18522
rect 8249 -18556 8281 -18522
rect 8321 -18556 8349 -18522
rect 8393 -18556 8417 -18522
rect 8451 -18556 8490 -18522
rect 8920 -18556 8959 -18522
rect 8993 -18556 9017 -18522
rect 9061 -18556 9089 -18522
rect 9129 -18556 9161 -18522
rect 9197 -18556 9231 -18522
rect 9267 -18556 9299 -18522
rect 9339 -18556 9367 -18522
rect 9411 -18556 9435 -18522
rect 9469 -18556 9508 -18522
rect 9938 -18556 9977 -18522
rect 10011 -18556 10035 -18522
rect 10079 -18556 10107 -18522
rect 10147 -18556 10179 -18522
rect 10215 -18556 10249 -18522
rect 10285 -18556 10317 -18522
rect 10357 -18556 10385 -18522
rect 10429 -18556 10453 -18522
rect 10487 -18556 10526 -18522
rect 10956 -18556 10995 -18522
rect 11029 -18556 11053 -18522
rect 11097 -18556 11125 -18522
rect 11165 -18556 11197 -18522
rect 11233 -18556 11267 -18522
rect 11303 -18556 11335 -18522
rect 11375 -18556 11403 -18522
rect 11447 -18556 11471 -18522
rect 11505 -18556 11544 -18522
rect 11974 -18556 12013 -18522
rect 12047 -18556 12071 -18522
rect 12115 -18556 12143 -18522
rect 12183 -18556 12215 -18522
rect 12251 -18556 12285 -18522
rect 12321 -18556 12353 -18522
rect 12393 -18556 12421 -18522
rect 12465 -18556 12489 -18522
rect 12523 -18556 12562 -18522
rect 12992 -18556 13031 -18522
rect 13065 -18556 13089 -18522
rect 13133 -18556 13161 -18522
rect 13201 -18556 13233 -18522
rect 13269 -18556 13303 -18522
rect 13339 -18556 13371 -18522
rect 13411 -18556 13439 -18522
rect 13483 -18556 13507 -18522
rect 13541 -18556 13580 -18522
rect 14010 -18556 14049 -18522
rect 14083 -18556 14107 -18522
rect 14151 -18556 14179 -18522
rect 14219 -18556 14251 -18522
rect 14287 -18556 14321 -18522
rect 14357 -18556 14389 -18522
rect 14429 -18556 14457 -18522
rect 14501 -18556 14525 -18522
rect 14559 -18556 14598 -18522
rect 15028 -18556 15067 -18522
rect 15101 -18556 15125 -18522
rect 15169 -18556 15197 -18522
rect 15237 -18556 15269 -18522
rect 15305 -18556 15339 -18522
rect 15375 -18556 15407 -18522
rect 15447 -18556 15475 -18522
rect 15519 -18556 15543 -18522
rect 15577 -18556 15616 -18522
rect 16046 -18556 16085 -18522
rect 16119 -18556 16143 -18522
rect 16187 -18556 16215 -18522
rect 16255 -18556 16287 -18522
rect 16323 -18556 16357 -18522
rect 16393 -18556 16425 -18522
rect 16465 -18556 16493 -18522
rect 16537 -18556 16561 -18522
rect 16595 -18556 16634 -18522
rect 17064 -18556 17103 -18522
rect 17137 -18556 17161 -18522
rect 17205 -18556 17233 -18522
rect 17273 -18556 17305 -18522
rect 17341 -18556 17375 -18522
rect 17411 -18556 17443 -18522
rect 17483 -18556 17511 -18522
rect 17555 -18556 17579 -18522
rect 17613 -18556 17652 -18522
rect 18082 -18556 18121 -18522
rect 18155 -18556 18179 -18522
rect 18223 -18556 18251 -18522
rect 18291 -18556 18323 -18522
rect 18359 -18556 18393 -18522
rect 18429 -18556 18461 -18522
rect 18501 -18556 18529 -18522
rect 18573 -18556 18597 -18522
rect 18631 -18556 18670 -18522
rect 19100 -18556 19139 -18522
rect 19173 -18556 19197 -18522
rect 19241 -18556 19269 -18522
rect 19309 -18556 19341 -18522
rect 19377 -18556 19411 -18522
rect 19447 -18556 19479 -18522
rect 19519 -18556 19547 -18522
rect 19591 -18556 19615 -18522
rect 19649 -18556 19688 -18522
rect 20118 -18556 20157 -18522
rect 20191 -18556 20215 -18522
rect 20259 -18556 20287 -18522
rect 20327 -18556 20359 -18522
rect 20395 -18556 20429 -18522
rect 20465 -18556 20497 -18522
rect 20537 -18556 20565 -18522
rect 20609 -18556 20633 -18522
rect 20667 -18556 20706 -18522
rect 21136 -18556 21175 -18522
rect 21209 -18556 21233 -18522
rect 21277 -18556 21305 -18522
rect 21345 -18556 21377 -18522
rect 21413 -18556 21447 -18522
rect 21483 -18556 21515 -18522
rect 21555 -18556 21583 -18522
rect 21627 -18556 21651 -18522
rect 21685 -18556 21724 -18522
rect 22154 -18556 22193 -18522
rect 22227 -18556 22251 -18522
rect 22295 -18556 22323 -18522
rect 22363 -18556 22395 -18522
rect 22431 -18556 22465 -18522
rect 22501 -18556 22533 -18522
rect 22573 -18556 22601 -18522
rect 22645 -18556 22669 -18522
rect 22703 -18556 22742 -18522
rect 24822 -18537 24855 -18499
rect 24889 -18537 24922 -18499
rect -22 -18623 12 -18591
rect -22 -18691 12 -18663
rect -22 -18759 12 -18735
rect -22 -18842 12 -18807
rect 24822 -18571 24922 -18537
rect 24822 -18605 24855 -18571
rect 24889 -18605 24922 -18571
rect 24822 -18639 24922 -18605
rect 24822 -18677 24855 -18639
rect 24889 -18677 24922 -18639
rect 24822 -18707 24922 -18677
rect 24822 -18749 24855 -18707
rect 24889 -18749 24922 -18707
rect 24822 -18775 24922 -18749
rect 24822 -18821 24855 -18775
rect 24889 -18821 24922 -18775
rect -12322 -18893 -12289 -18843
rect -12255 -18893 -12222 -18843
rect 24822 -18843 24922 -18821
rect -12322 -18911 -12222 -18893
rect -8952 -18910 -8913 -18876
rect -8879 -18910 -8855 -18876
rect -8811 -18910 -8783 -18876
rect -8743 -18910 -8711 -18876
rect -8675 -18910 -8641 -18876
rect -8605 -18910 -8573 -18876
rect -8533 -18910 -8505 -18876
rect -8461 -18910 -8437 -18876
rect -8403 -18910 -8364 -18876
rect -7934 -18910 -7895 -18876
rect -7861 -18910 -7837 -18876
rect -7793 -18910 -7765 -18876
rect -7725 -18910 -7693 -18876
rect -7657 -18910 -7623 -18876
rect -7587 -18910 -7555 -18876
rect -7515 -18910 -7487 -18876
rect -7443 -18910 -7419 -18876
rect -7385 -18910 -7346 -18876
rect -6916 -18910 -6877 -18876
rect -6843 -18910 -6819 -18876
rect -6775 -18910 -6747 -18876
rect -6707 -18910 -6675 -18876
rect -6639 -18910 -6605 -18876
rect -6569 -18910 -6537 -18876
rect -6497 -18910 -6469 -18876
rect -6425 -18910 -6401 -18876
rect -6367 -18910 -6328 -18876
rect -5898 -18910 -5859 -18876
rect -5825 -18910 -5801 -18876
rect -5757 -18910 -5729 -18876
rect -5689 -18910 -5657 -18876
rect -5621 -18910 -5587 -18876
rect -5551 -18910 -5519 -18876
rect -5479 -18910 -5451 -18876
rect -5407 -18910 -5383 -18876
rect -5349 -18910 -5310 -18876
rect -4880 -18910 -4841 -18876
rect -4807 -18910 -4783 -18876
rect -4739 -18910 -4711 -18876
rect -4671 -18910 -4639 -18876
rect -4603 -18910 -4569 -18876
rect -4533 -18910 -4501 -18876
rect -4461 -18910 -4433 -18876
rect -4389 -18910 -4365 -18876
rect -4331 -18910 -4292 -18876
rect -3862 -18910 -3823 -18876
rect -3789 -18910 -3765 -18876
rect -3721 -18910 -3693 -18876
rect -3653 -18910 -3621 -18876
rect -3585 -18910 -3551 -18876
rect -3515 -18910 -3483 -18876
rect -3443 -18910 -3415 -18876
rect -3371 -18910 -3347 -18876
rect -3313 -18910 -3274 -18876
rect -2844 -18910 -2805 -18876
rect -2771 -18910 -2747 -18876
rect -2703 -18910 -2675 -18876
rect -2635 -18910 -2603 -18876
rect -2567 -18910 -2533 -18876
rect -2497 -18910 -2465 -18876
rect -2425 -18910 -2397 -18876
rect -2353 -18910 -2329 -18876
rect -2295 -18910 -2256 -18876
rect -1826 -18910 -1787 -18876
rect -1753 -18910 -1729 -18876
rect -1685 -18910 -1657 -18876
rect -1617 -18910 -1585 -18876
rect -1549 -18910 -1515 -18876
rect -1479 -18910 -1447 -18876
rect -1407 -18910 -1379 -18876
rect -1335 -18910 -1311 -18876
rect -1277 -18910 -1238 -18876
rect -808 -18910 -769 -18876
rect -735 -18910 -711 -18876
rect -667 -18910 -639 -18876
rect -599 -18910 -567 -18876
rect -531 -18910 -497 -18876
rect -461 -18910 -429 -18876
rect -389 -18910 -361 -18876
rect -317 -18910 -293 -18876
rect -259 -18910 -220 -18876
rect 24822 -18893 24855 -18843
rect 24889 -18893 24922 -18843
rect -12322 -18965 -12289 -18911
rect -12255 -18965 -12222 -18911
rect -12322 -18979 -12222 -18965
rect -12322 -19037 -12289 -18979
rect -12255 -19037 -12222 -18979
rect -12322 -19047 -12222 -19037
rect 24822 -18911 24922 -18893
rect 24822 -18965 24855 -18911
rect 24889 -18965 24922 -18911
rect 24822 -18979 24922 -18965
rect 24822 -19037 24855 -18979
rect 24889 -19037 24922 -18979
rect -12322 -19109 -12289 -19047
rect -12255 -19109 -12222 -19047
rect 2812 -19080 2851 -19046
rect 2885 -19080 2909 -19046
rect 2953 -19080 2981 -19046
rect 3021 -19080 3053 -19046
rect 3089 -19080 3123 -19046
rect 3159 -19080 3191 -19046
rect 3231 -19080 3259 -19046
rect 3303 -19080 3327 -19046
rect 3361 -19080 3400 -19046
rect 3830 -19080 3869 -19046
rect 3903 -19080 3927 -19046
rect 3971 -19080 3999 -19046
rect 4039 -19080 4071 -19046
rect 4107 -19080 4141 -19046
rect 4177 -19080 4209 -19046
rect 4249 -19080 4277 -19046
rect 4321 -19080 4345 -19046
rect 4379 -19080 4418 -19046
rect 4848 -19080 4887 -19046
rect 4921 -19080 4945 -19046
rect 4989 -19080 5017 -19046
rect 5057 -19080 5089 -19046
rect 5125 -19080 5159 -19046
rect 5195 -19080 5227 -19046
rect 5267 -19080 5295 -19046
rect 5339 -19080 5363 -19046
rect 5397 -19080 5436 -19046
rect 5866 -19080 5905 -19046
rect 5939 -19080 5963 -19046
rect 6007 -19080 6035 -19046
rect 6075 -19080 6107 -19046
rect 6143 -19080 6177 -19046
rect 6213 -19080 6245 -19046
rect 6285 -19080 6313 -19046
rect 6357 -19080 6381 -19046
rect 6415 -19080 6454 -19046
rect 6884 -19080 6923 -19046
rect 6957 -19080 6981 -19046
rect 7025 -19080 7053 -19046
rect 7093 -19080 7125 -19046
rect 7161 -19080 7195 -19046
rect 7231 -19080 7263 -19046
rect 7303 -19080 7331 -19046
rect 7375 -19080 7399 -19046
rect 7433 -19080 7472 -19046
rect 7902 -19080 7941 -19046
rect 7975 -19080 7999 -19046
rect 8043 -19080 8071 -19046
rect 8111 -19080 8143 -19046
rect 8179 -19080 8213 -19046
rect 8249 -19080 8281 -19046
rect 8321 -19080 8349 -19046
rect 8393 -19080 8417 -19046
rect 8451 -19080 8490 -19046
rect 8920 -19080 8959 -19046
rect 8993 -19080 9017 -19046
rect 9061 -19080 9089 -19046
rect 9129 -19080 9161 -19046
rect 9197 -19080 9231 -19046
rect 9267 -19080 9299 -19046
rect 9339 -19080 9367 -19046
rect 9411 -19080 9435 -19046
rect 9469 -19080 9508 -19046
rect 9938 -19080 9977 -19046
rect 10011 -19080 10035 -19046
rect 10079 -19080 10107 -19046
rect 10147 -19080 10179 -19046
rect 10215 -19080 10249 -19046
rect 10285 -19080 10317 -19046
rect 10357 -19080 10385 -19046
rect 10429 -19080 10453 -19046
rect 10487 -19080 10526 -19046
rect 10956 -19080 10995 -19046
rect 11029 -19080 11053 -19046
rect 11097 -19080 11125 -19046
rect 11165 -19080 11197 -19046
rect 11233 -19080 11267 -19046
rect 11303 -19080 11335 -19046
rect 11375 -19080 11403 -19046
rect 11447 -19080 11471 -19046
rect 11505 -19080 11544 -19046
rect 11974 -19080 12013 -19046
rect 12047 -19080 12071 -19046
rect 12115 -19080 12143 -19046
rect 12183 -19080 12215 -19046
rect 12251 -19080 12285 -19046
rect 12321 -19080 12353 -19046
rect 12393 -19080 12421 -19046
rect 12465 -19080 12489 -19046
rect 12523 -19080 12562 -19046
rect 12992 -19080 13031 -19046
rect 13065 -19080 13089 -19046
rect 13133 -19080 13161 -19046
rect 13201 -19080 13233 -19046
rect 13269 -19080 13303 -19046
rect 13339 -19080 13371 -19046
rect 13411 -19080 13439 -19046
rect 13483 -19080 13507 -19046
rect 13541 -19080 13580 -19046
rect 14010 -19080 14049 -19046
rect 14083 -19080 14107 -19046
rect 14151 -19080 14179 -19046
rect 14219 -19080 14251 -19046
rect 14287 -19080 14321 -19046
rect 14357 -19080 14389 -19046
rect 14429 -19080 14457 -19046
rect 14501 -19080 14525 -19046
rect 14559 -19080 14598 -19046
rect 15028 -19080 15067 -19046
rect 15101 -19080 15125 -19046
rect 15169 -19080 15197 -19046
rect 15237 -19080 15269 -19046
rect 15305 -19080 15339 -19046
rect 15375 -19080 15407 -19046
rect 15447 -19080 15475 -19046
rect 15519 -19080 15543 -19046
rect 15577 -19080 15616 -19046
rect 16046 -19080 16085 -19046
rect 16119 -19080 16143 -19046
rect 16187 -19080 16215 -19046
rect 16255 -19080 16287 -19046
rect 16323 -19080 16357 -19046
rect 16393 -19080 16425 -19046
rect 16465 -19080 16493 -19046
rect 16537 -19080 16561 -19046
rect 16595 -19080 16634 -19046
rect 17064 -19080 17103 -19046
rect 17137 -19080 17161 -19046
rect 17205 -19080 17233 -19046
rect 17273 -19080 17305 -19046
rect 17341 -19080 17375 -19046
rect 17411 -19080 17443 -19046
rect 17483 -19080 17511 -19046
rect 17555 -19080 17579 -19046
rect 17613 -19080 17652 -19046
rect 18082 -19080 18121 -19046
rect 18155 -19080 18179 -19046
rect 18223 -19080 18251 -19046
rect 18291 -19080 18323 -19046
rect 18359 -19080 18393 -19046
rect 18429 -19080 18461 -19046
rect 18501 -19080 18529 -19046
rect 18573 -19080 18597 -19046
rect 18631 -19080 18670 -19046
rect 19100 -19080 19139 -19046
rect 19173 -19080 19197 -19046
rect 19241 -19080 19269 -19046
rect 19309 -19080 19341 -19046
rect 19377 -19080 19411 -19046
rect 19447 -19080 19479 -19046
rect 19519 -19080 19547 -19046
rect 19591 -19080 19615 -19046
rect 19649 -19080 19688 -19046
rect 20118 -19080 20157 -19046
rect 20191 -19080 20215 -19046
rect 20259 -19080 20287 -19046
rect 20327 -19080 20359 -19046
rect 20395 -19080 20429 -19046
rect 20465 -19080 20497 -19046
rect 20537 -19080 20565 -19046
rect 20609 -19080 20633 -19046
rect 20667 -19080 20706 -19046
rect 21136 -19080 21175 -19046
rect 21209 -19080 21233 -19046
rect 21277 -19080 21305 -19046
rect 21345 -19080 21377 -19046
rect 21413 -19080 21447 -19046
rect 21483 -19080 21515 -19046
rect 21555 -19080 21583 -19046
rect 21627 -19080 21651 -19046
rect 21685 -19080 21724 -19046
rect 22154 -19080 22193 -19046
rect 22227 -19080 22251 -19046
rect 22295 -19080 22323 -19046
rect 22363 -19080 22395 -19046
rect 22431 -19080 22465 -19046
rect 22501 -19080 22533 -19046
rect 22573 -19080 22601 -19046
rect 22645 -19080 22669 -19046
rect 22703 -19080 22742 -19046
rect 24822 -19047 24922 -19037
rect -12322 -19115 -12222 -19109
rect 24822 -19109 24855 -19047
rect 24889 -19109 24922 -19047
rect -12322 -19181 -12289 -19115
rect -12255 -19181 -12222 -19115
rect -12322 -19183 -12222 -19181
rect -12322 -19217 -12289 -19183
rect -12255 -19217 -12222 -19183
rect -12322 -19219 -12222 -19217
rect -12322 -19285 -12289 -19219
rect -12255 -19285 -12222 -19219
rect -12322 -19291 -12222 -19285
rect -12322 -19353 -12289 -19291
rect -12255 -19353 -12222 -19291
rect -12322 -19363 -12222 -19353
rect -12322 -19421 -12289 -19363
rect -12255 -19421 -12222 -19363
rect -12322 -19435 -12222 -19421
rect -12322 -19489 -12289 -19435
rect -12255 -19489 -12222 -19435
rect -12322 -19507 -12222 -19489
rect -12322 -19557 -12289 -19507
rect -12255 -19557 -12222 -19507
rect 2580 -19149 2614 -19114
rect 2580 -19221 2614 -19197
rect 2580 -19293 2614 -19265
rect 2580 -19365 2614 -19333
rect 2580 -19435 2614 -19401
rect 2580 -19503 2614 -19471
rect -12322 -19579 -12222 -19557
rect -12322 -19625 -12289 -19579
rect -12255 -19625 -12222 -19579
rect -2252 -19584 -2215 -19550
rect -2181 -19584 -2144 -19550
rect -2034 -19584 -1997 -19550
rect -1963 -19584 -1926 -19550
rect -1816 -19584 -1779 -19550
rect -1745 -19584 -1708 -19550
rect -1598 -19584 -1561 -19550
rect -1527 -19584 -1490 -19550
rect -1380 -19584 -1343 -19550
rect -1309 -19584 -1272 -19550
rect -1162 -19584 -1125 -19550
rect -1091 -19584 -1054 -19550
rect -944 -19584 -907 -19550
rect -873 -19584 -836 -19550
rect -726 -19584 -689 -19550
rect -655 -19584 -618 -19550
rect -508 -19584 -471 -19550
rect -437 -19584 -400 -19550
rect -290 -19584 -253 -19550
rect -219 -19584 -182 -19550
rect 2580 -19571 2614 -19543
rect -12322 -19651 -12222 -19625
rect -12322 -19693 -12289 -19651
rect -12255 -19693 -12222 -19651
rect -12322 -19723 -12222 -19693
rect -12322 -19761 -12289 -19723
rect -12255 -19761 -12222 -19723
rect -12322 -19795 -12222 -19761
rect -12322 -19829 -12289 -19795
rect -12255 -19829 -12222 -19795
rect -2324 -19637 -2290 -19618
rect -2324 -19705 -2290 -19703
rect -2324 -19741 -2290 -19739
rect -2324 -19826 -2290 -19807
rect -2106 -19637 -2072 -19618
rect -2106 -19705 -2072 -19703
rect -2106 -19741 -2072 -19739
rect -2106 -19826 -2072 -19807
rect -1888 -19637 -1854 -19618
rect -1888 -19705 -1854 -19703
rect -1888 -19741 -1854 -19739
rect -1888 -19826 -1854 -19807
rect -1670 -19637 -1636 -19618
rect -1670 -19705 -1636 -19703
rect -1670 -19741 -1636 -19739
rect -1670 -19826 -1636 -19807
rect -1452 -19637 -1418 -19618
rect -1452 -19705 -1418 -19703
rect -1452 -19741 -1418 -19739
rect -1452 -19826 -1418 -19807
rect -1234 -19637 -1200 -19618
rect -1234 -19705 -1200 -19703
rect -1234 -19741 -1200 -19739
rect -1234 -19826 -1200 -19807
rect -1016 -19637 -982 -19618
rect -1016 -19705 -982 -19703
rect -1016 -19741 -982 -19739
rect -1016 -19826 -982 -19807
rect -798 -19637 -764 -19618
rect -798 -19705 -764 -19703
rect -798 -19741 -764 -19739
rect -798 -19826 -764 -19807
rect -580 -19637 -546 -19618
rect -580 -19705 -546 -19703
rect -580 -19741 -546 -19739
rect -580 -19826 -546 -19807
rect -362 -19637 -328 -19618
rect -362 -19705 -328 -19703
rect -362 -19741 -328 -19739
rect -362 -19826 -328 -19807
rect -144 -19637 -110 -19618
rect -144 -19705 -110 -19703
rect 2580 -19639 2614 -19615
rect 2580 -19722 2614 -19687
rect 3598 -19149 3632 -19114
rect 3598 -19221 3632 -19197
rect 3598 -19293 3632 -19265
rect 3598 -19365 3632 -19333
rect 3598 -19435 3632 -19401
rect 3598 -19503 3632 -19471
rect 3598 -19571 3632 -19543
rect 3598 -19639 3632 -19615
rect 3598 -19722 3632 -19687
rect 4616 -19149 4650 -19114
rect 4616 -19221 4650 -19197
rect 4616 -19293 4650 -19265
rect 4616 -19365 4650 -19333
rect 4616 -19435 4650 -19401
rect 4616 -19503 4650 -19471
rect 4616 -19571 4650 -19543
rect 4616 -19639 4650 -19615
rect 4616 -19722 4650 -19687
rect 5634 -19149 5668 -19114
rect 5634 -19221 5668 -19197
rect 5634 -19293 5668 -19265
rect 5634 -19365 5668 -19333
rect 5634 -19435 5668 -19401
rect 5634 -19503 5668 -19471
rect 5634 -19571 5668 -19543
rect 5634 -19639 5668 -19615
rect 5634 -19722 5668 -19687
rect 6652 -19149 6686 -19114
rect 6652 -19221 6686 -19197
rect 6652 -19293 6686 -19265
rect 6652 -19365 6686 -19333
rect 6652 -19435 6686 -19401
rect 6652 -19503 6686 -19471
rect 6652 -19571 6686 -19543
rect 6652 -19639 6686 -19615
rect 6652 -19722 6686 -19687
rect 7670 -19149 7704 -19114
rect 7670 -19221 7704 -19197
rect 7670 -19293 7704 -19265
rect 7670 -19365 7704 -19333
rect 7670 -19435 7704 -19401
rect 7670 -19503 7704 -19471
rect 7670 -19571 7704 -19543
rect 7670 -19639 7704 -19615
rect 7670 -19722 7704 -19687
rect 8688 -19149 8722 -19114
rect 8688 -19221 8722 -19197
rect 8688 -19293 8722 -19265
rect 8688 -19365 8722 -19333
rect 8688 -19435 8722 -19401
rect 8688 -19503 8722 -19471
rect 8688 -19571 8722 -19543
rect 8688 -19639 8722 -19615
rect 8688 -19722 8722 -19687
rect 9706 -19149 9740 -19114
rect 9706 -19221 9740 -19197
rect 9706 -19293 9740 -19265
rect 9706 -19365 9740 -19333
rect 9706 -19435 9740 -19401
rect 9706 -19503 9740 -19471
rect 9706 -19571 9740 -19543
rect 9706 -19639 9740 -19615
rect 9706 -19722 9740 -19687
rect 10724 -19149 10758 -19114
rect 10724 -19221 10758 -19197
rect 10724 -19293 10758 -19265
rect 10724 -19365 10758 -19333
rect 10724 -19435 10758 -19401
rect 10724 -19503 10758 -19471
rect 10724 -19571 10758 -19543
rect 10724 -19639 10758 -19615
rect 10724 -19722 10758 -19687
rect 11742 -19149 11776 -19114
rect 11742 -19221 11776 -19197
rect 11742 -19293 11776 -19265
rect 11742 -19365 11776 -19333
rect 11742 -19435 11776 -19401
rect 11742 -19503 11776 -19471
rect 11742 -19571 11776 -19543
rect 11742 -19639 11776 -19615
rect 11742 -19722 11776 -19687
rect 12760 -19149 12794 -19114
rect 12760 -19221 12794 -19197
rect 12760 -19293 12794 -19265
rect 12760 -19365 12794 -19333
rect 12760 -19435 12794 -19401
rect 12760 -19503 12794 -19471
rect 12760 -19571 12794 -19543
rect 12760 -19639 12794 -19615
rect 12760 -19722 12794 -19687
rect 13778 -19149 13812 -19114
rect 13778 -19221 13812 -19197
rect 13778 -19293 13812 -19265
rect 13778 -19365 13812 -19333
rect 13778 -19435 13812 -19401
rect 13778 -19503 13812 -19471
rect 13778 -19571 13812 -19543
rect 13778 -19639 13812 -19615
rect 13778 -19722 13812 -19687
rect 14796 -19149 14830 -19114
rect 14796 -19221 14830 -19197
rect 14796 -19293 14830 -19265
rect 14796 -19365 14830 -19333
rect 14796 -19435 14830 -19401
rect 14796 -19503 14830 -19471
rect 14796 -19571 14830 -19543
rect 14796 -19639 14830 -19615
rect 14796 -19722 14830 -19687
rect 15814 -19149 15848 -19114
rect 15814 -19221 15848 -19197
rect 15814 -19293 15848 -19265
rect 15814 -19365 15848 -19333
rect 15814 -19435 15848 -19401
rect 15814 -19503 15848 -19471
rect 15814 -19571 15848 -19543
rect 15814 -19639 15848 -19615
rect 15814 -19722 15848 -19687
rect 16832 -19149 16866 -19114
rect 16832 -19221 16866 -19197
rect 16832 -19293 16866 -19265
rect 16832 -19365 16866 -19333
rect 16832 -19435 16866 -19401
rect 16832 -19503 16866 -19471
rect 16832 -19571 16866 -19543
rect 16832 -19639 16866 -19615
rect 16832 -19722 16866 -19687
rect 17850 -19149 17884 -19114
rect 17850 -19221 17884 -19197
rect 17850 -19293 17884 -19265
rect 17850 -19365 17884 -19333
rect 17850 -19435 17884 -19401
rect 17850 -19503 17884 -19471
rect 17850 -19571 17884 -19543
rect 17850 -19639 17884 -19615
rect 17850 -19722 17884 -19687
rect 18868 -19149 18902 -19114
rect 18868 -19221 18902 -19197
rect 18868 -19293 18902 -19265
rect 18868 -19365 18902 -19333
rect 18868 -19435 18902 -19401
rect 18868 -19503 18902 -19471
rect 18868 -19571 18902 -19543
rect 18868 -19639 18902 -19615
rect 18868 -19722 18902 -19687
rect 19886 -19149 19920 -19114
rect 19886 -19221 19920 -19197
rect 19886 -19293 19920 -19265
rect 19886 -19365 19920 -19333
rect 19886 -19435 19920 -19401
rect 19886 -19503 19920 -19471
rect 19886 -19571 19920 -19543
rect 19886 -19639 19920 -19615
rect 19886 -19722 19920 -19687
rect 20904 -19149 20938 -19114
rect 20904 -19221 20938 -19197
rect 20904 -19293 20938 -19265
rect 20904 -19365 20938 -19333
rect 20904 -19435 20938 -19401
rect 20904 -19503 20938 -19471
rect 20904 -19571 20938 -19543
rect 20904 -19639 20938 -19615
rect 20904 -19722 20938 -19687
rect 21922 -19149 21956 -19114
rect 21922 -19221 21956 -19197
rect 21922 -19293 21956 -19265
rect 21922 -19365 21956 -19333
rect 21922 -19435 21956 -19401
rect 21922 -19503 21956 -19471
rect 21922 -19571 21956 -19543
rect 21922 -19639 21956 -19615
rect 21922 -19722 21956 -19687
rect 22940 -19149 22974 -19114
rect 22940 -19221 22974 -19197
rect 22940 -19293 22974 -19265
rect 22940 -19365 22974 -19333
rect 22940 -19435 22974 -19401
rect 22940 -19503 22974 -19471
rect 22940 -19571 22974 -19543
rect 22940 -19639 22974 -19615
rect 22940 -19722 22974 -19687
rect 24822 -19115 24922 -19109
rect 24822 -19181 24855 -19115
rect 24889 -19181 24922 -19115
rect 24822 -19183 24922 -19181
rect 24822 -19217 24855 -19183
rect 24889 -19217 24922 -19183
rect 24822 -19219 24922 -19217
rect 24822 -19285 24855 -19219
rect 24889 -19285 24922 -19219
rect 24822 -19291 24922 -19285
rect 24822 -19353 24855 -19291
rect 24889 -19353 24922 -19291
rect 24822 -19363 24922 -19353
rect 24822 -19421 24855 -19363
rect 24889 -19421 24922 -19363
rect 24822 -19435 24922 -19421
rect 24822 -19489 24855 -19435
rect 24889 -19489 24922 -19435
rect 24822 -19507 24922 -19489
rect 24822 -19557 24855 -19507
rect 24889 -19557 24922 -19507
rect 24822 -19579 24922 -19557
rect 24822 -19625 24855 -19579
rect 24889 -19625 24922 -19579
rect 24822 -19651 24922 -19625
rect 24822 -19693 24855 -19651
rect 24889 -19693 24922 -19651
rect -144 -19741 -110 -19739
rect 24822 -19723 24922 -19693
rect 5106 -19756 5166 -19752
rect 2812 -19790 2851 -19756
rect 2885 -19790 2909 -19756
rect 2953 -19790 2981 -19756
rect 3021 -19790 3053 -19756
rect 3089 -19790 3123 -19756
rect 3159 -19790 3191 -19756
rect 3231 -19790 3259 -19756
rect 3303 -19790 3327 -19756
rect 3361 -19790 3400 -19756
rect 3830 -19790 3869 -19756
rect 3903 -19790 3927 -19756
rect 3971 -19790 3999 -19756
rect 4039 -19790 4071 -19756
rect 4107 -19790 4141 -19756
rect 4177 -19790 4209 -19756
rect 4249 -19790 4277 -19756
rect 4321 -19790 4345 -19756
rect 4379 -19790 4418 -19756
rect 4848 -19790 4887 -19756
rect 4921 -19790 4945 -19756
rect 4989 -19790 5017 -19756
rect 5057 -19790 5089 -19756
rect 5125 -19790 5159 -19756
rect 5195 -19790 5227 -19756
rect 5267 -19790 5295 -19756
rect 5339 -19790 5363 -19756
rect 5397 -19790 5436 -19756
rect 5866 -19790 5905 -19756
rect 5939 -19790 5963 -19756
rect 6007 -19790 6035 -19756
rect 6075 -19790 6107 -19756
rect 6143 -19790 6177 -19756
rect 6213 -19790 6245 -19756
rect 6285 -19790 6313 -19756
rect 6357 -19790 6381 -19756
rect 6415 -19790 6454 -19756
rect 6884 -19790 6923 -19756
rect 6957 -19790 6981 -19756
rect 7025 -19790 7053 -19756
rect 7093 -19790 7125 -19756
rect 7161 -19790 7195 -19756
rect 7231 -19790 7263 -19756
rect 7303 -19790 7331 -19756
rect 7375 -19790 7399 -19756
rect 7433 -19790 7472 -19756
rect 7902 -19790 7941 -19756
rect 7975 -19790 7999 -19756
rect 8043 -19790 8071 -19756
rect 8111 -19790 8143 -19756
rect 8179 -19790 8213 -19756
rect 8249 -19790 8281 -19756
rect 8321 -19790 8349 -19756
rect 8393 -19790 8417 -19756
rect 8451 -19790 8490 -19756
rect 8920 -19790 8959 -19756
rect 8993 -19790 9017 -19756
rect 9061 -19790 9089 -19756
rect 9129 -19790 9161 -19756
rect 9197 -19790 9231 -19756
rect 9267 -19790 9299 -19756
rect 9339 -19790 9367 -19756
rect 9411 -19790 9435 -19756
rect 9469 -19790 9508 -19756
rect 9938 -19790 9977 -19756
rect 10011 -19790 10035 -19756
rect 10079 -19790 10107 -19756
rect 10147 -19790 10179 -19756
rect 10215 -19790 10249 -19756
rect 10285 -19790 10317 -19756
rect 10357 -19790 10385 -19756
rect 10429 -19790 10453 -19756
rect 10487 -19790 10526 -19756
rect 10956 -19790 10995 -19756
rect 11029 -19790 11053 -19756
rect 11097 -19790 11125 -19756
rect 11165 -19790 11197 -19756
rect 11233 -19790 11267 -19756
rect 11303 -19790 11335 -19756
rect 11375 -19790 11403 -19756
rect 11447 -19790 11471 -19756
rect 11505 -19790 11544 -19756
rect 11974 -19790 12013 -19756
rect 12047 -19790 12071 -19756
rect 12115 -19790 12143 -19756
rect 12183 -19790 12215 -19756
rect 12251 -19790 12285 -19756
rect 12321 -19790 12353 -19756
rect 12393 -19790 12421 -19756
rect 12465 -19790 12489 -19756
rect 12523 -19790 12562 -19756
rect 12992 -19790 13031 -19756
rect 13065 -19790 13089 -19756
rect 13133 -19790 13161 -19756
rect 13201 -19790 13233 -19756
rect 13269 -19790 13303 -19756
rect 13339 -19790 13371 -19756
rect 13411 -19790 13439 -19756
rect 13483 -19790 13507 -19756
rect 13541 -19790 13580 -19756
rect 14010 -19790 14049 -19756
rect 14083 -19790 14107 -19756
rect 14151 -19790 14179 -19756
rect 14219 -19790 14251 -19756
rect 14287 -19790 14321 -19756
rect 14357 -19790 14389 -19756
rect 14429 -19790 14457 -19756
rect 14501 -19790 14525 -19756
rect 14559 -19790 14598 -19756
rect 15028 -19790 15067 -19756
rect 15101 -19790 15125 -19756
rect 15169 -19790 15197 -19756
rect 15237 -19790 15269 -19756
rect 15305 -19790 15339 -19756
rect 15375 -19790 15407 -19756
rect 15447 -19790 15475 -19756
rect 15519 -19790 15543 -19756
rect 15577 -19790 15616 -19756
rect 16046 -19790 16085 -19756
rect 16119 -19790 16143 -19756
rect 16187 -19790 16215 -19756
rect 16255 -19790 16287 -19756
rect 16323 -19790 16357 -19756
rect 16393 -19790 16425 -19756
rect 16465 -19790 16493 -19756
rect 16537 -19790 16561 -19756
rect 16595 -19790 16634 -19756
rect 17064 -19790 17103 -19756
rect 17137 -19790 17161 -19756
rect 17205 -19790 17233 -19756
rect 17273 -19790 17305 -19756
rect 17341 -19790 17375 -19756
rect 17411 -19790 17443 -19756
rect 17483 -19790 17511 -19756
rect 17555 -19790 17579 -19756
rect 17613 -19790 17652 -19756
rect 18082 -19790 18121 -19756
rect 18155 -19790 18179 -19756
rect 18223 -19790 18251 -19756
rect 18291 -19790 18323 -19756
rect 18359 -19790 18393 -19756
rect 18429 -19790 18461 -19756
rect 18501 -19790 18529 -19756
rect 18573 -19790 18597 -19756
rect 18631 -19790 18670 -19756
rect 19100 -19790 19139 -19756
rect 19173 -19790 19197 -19756
rect 19241 -19790 19269 -19756
rect 19309 -19790 19341 -19756
rect 19377 -19790 19411 -19756
rect 19447 -19790 19479 -19756
rect 19519 -19790 19547 -19756
rect 19591 -19790 19615 -19756
rect 19649 -19790 19688 -19756
rect 20118 -19790 20157 -19756
rect 20191 -19790 20215 -19756
rect 20259 -19790 20287 -19756
rect 20327 -19790 20359 -19756
rect 20395 -19790 20429 -19756
rect 20465 -19790 20497 -19756
rect 20537 -19790 20565 -19756
rect 20609 -19790 20633 -19756
rect 20667 -19790 20706 -19756
rect 21136 -19790 21175 -19756
rect 21209 -19790 21233 -19756
rect 21277 -19790 21305 -19756
rect 21345 -19790 21377 -19756
rect 21413 -19790 21447 -19756
rect 21483 -19790 21515 -19756
rect 21555 -19790 21583 -19756
rect 21627 -19790 21651 -19756
rect 21685 -19790 21724 -19756
rect 22154 -19790 22193 -19756
rect 22227 -19790 22251 -19756
rect 22295 -19790 22323 -19756
rect 22363 -19790 22395 -19756
rect 22431 -19790 22465 -19756
rect 22501 -19790 22533 -19756
rect 22573 -19790 22601 -19756
rect 22645 -19790 22669 -19756
rect 22703 -19790 22742 -19756
rect 24822 -19761 24855 -19723
rect 24889 -19761 24922 -19723
rect -144 -19826 -110 -19807
rect 24822 -19795 24922 -19761
rect -12322 -19863 -12222 -19829
rect 24822 -19829 24855 -19795
rect 24889 -19829 24922 -19795
rect -12322 -19901 -12289 -19863
rect -12255 -19901 -12222 -19863
rect -2252 -19894 -2215 -19860
rect -2181 -19894 -2144 -19860
rect -2034 -19894 -1997 -19860
rect -1963 -19894 -1926 -19860
rect -1816 -19894 -1779 -19860
rect -1745 -19894 -1708 -19860
rect -1598 -19894 -1561 -19860
rect -1527 -19894 -1490 -19860
rect -1380 -19894 -1343 -19860
rect -1309 -19894 -1272 -19860
rect -1162 -19894 -1125 -19860
rect -1091 -19894 -1054 -19860
rect -944 -19894 -907 -19860
rect -873 -19894 -836 -19860
rect -726 -19894 -689 -19860
rect -655 -19894 -618 -19860
rect -508 -19894 -471 -19860
rect -437 -19894 -400 -19860
rect -290 -19894 -253 -19860
rect -219 -19894 -182 -19860
rect 24822 -19863 24922 -19829
rect -12322 -19931 -12222 -19901
rect -12322 -19973 -12289 -19931
rect -12255 -19973 -12222 -19931
rect -12322 -19999 -12222 -19973
rect -12322 -20045 -12289 -19999
rect -12255 -20045 -12222 -19999
rect -12322 -20067 -12222 -20045
rect -12322 -20117 -12289 -20067
rect -12255 -20117 -12222 -20067
rect -12322 -20135 -12222 -20117
rect -12322 -20189 -12289 -20135
rect -12255 -20189 -12222 -20135
rect -12322 -20203 -12222 -20189
rect -12322 -20261 -12289 -20203
rect -12255 -20261 -12222 -20203
rect -12322 -20271 -12222 -20261
rect -12322 -20333 -12289 -20271
rect -12255 -20333 -12222 -20271
rect 24822 -19901 24855 -19863
rect 24889 -19901 24922 -19863
rect 24822 -19931 24922 -19901
rect 24822 -19973 24855 -19931
rect 24889 -19973 24922 -19931
rect 24822 -19999 24922 -19973
rect 24822 -20045 24855 -19999
rect 24889 -20045 24922 -19999
rect 24822 -20067 24922 -20045
rect 24822 -20117 24855 -20067
rect 24889 -20117 24922 -20067
rect 24822 -20135 24922 -20117
rect 24822 -20189 24855 -20135
rect 24889 -20189 24922 -20135
rect 24822 -20203 24922 -20189
rect 24822 -20261 24855 -20203
rect 24889 -20261 24922 -20203
rect 24822 -20271 24922 -20261
rect 2812 -20314 2851 -20280
rect 2885 -20314 2909 -20280
rect 2953 -20314 2981 -20280
rect 3021 -20314 3053 -20280
rect 3089 -20314 3123 -20280
rect 3159 -20314 3191 -20280
rect 3231 -20314 3259 -20280
rect 3303 -20314 3327 -20280
rect 3361 -20314 3400 -20280
rect 3830 -20314 3869 -20280
rect 3903 -20314 3927 -20280
rect 3971 -20314 3999 -20280
rect 4039 -20314 4071 -20280
rect 4107 -20314 4141 -20280
rect 4177 -20314 4209 -20280
rect 4249 -20314 4277 -20280
rect 4321 -20314 4345 -20280
rect 4379 -20314 4418 -20280
rect 4848 -20314 4887 -20280
rect 4921 -20314 4945 -20280
rect 4989 -20314 5017 -20280
rect 5057 -20314 5089 -20280
rect 5125 -20314 5159 -20280
rect 5195 -20314 5227 -20280
rect 5267 -20314 5295 -20280
rect 5339 -20314 5363 -20280
rect 5397 -20314 5436 -20280
rect 5866 -20314 5905 -20280
rect 5939 -20314 5963 -20280
rect 6007 -20314 6035 -20280
rect 6075 -20314 6107 -20280
rect 6143 -20314 6177 -20280
rect 6213 -20314 6245 -20280
rect 6285 -20314 6313 -20280
rect 6357 -20314 6381 -20280
rect 6415 -20314 6454 -20280
rect 6884 -20314 6923 -20280
rect 6957 -20314 6981 -20280
rect 7025 -20314 7053 -20280
rect 7093 -20314 7125 -20280
rect 7161 -20314 7195 -20280
rect 7231 -20314 7263 -20280
rect 7303 -20314 7331 -20280
rect 7375 -20314 7399 -20280
rect 7433 -20314 7472 -20280
rect 7902 -20314 7941 -20280
rect 7975 -20314 7999 -20280
rect 8043 -20314 8071 -20280
rect 8111 -20314 8143 -20280
rect 8179 -20314 8213 -20280
rect 8249 -20314 8281 -20280
rect 8321 -20314 8349 -20280
rect 8393 -20314 8417 -20280
rect 8451 -20314 8490 -20280
rect 8920 -20314 8959 -20280
rect 8993 -20314 9017 -20280
rect 9061 -20314 9089 -20280
rect 9129 -20314 9161 -20280
rect 9197 -20314 9231 -20280
rect 9267 -20314 9299 -20280
rect 9339 -20314 9367 -20280
rect 9411 -20314 9435 -20280
rect 9469 -20314 9508 -20280
rect 9938 -20314 9977 -20280
rect 10011 -20314 10035 -20280
rect 10079 -20314 10107 -20280
rect 10147 -20314 10179 -20280
rect 10215 -20314 10249 -20280
rect 10285 -20314 10317 -20280
rect 10357 -20314 10385 -20280
rect 10429 -20314 10453 -20280
rect 10487 -20314 10526 -20280
rect 10956 -20314 10995 -20280
rect 11029 -20314 11053 -20280
rect 11097 -20314 11125 -20280
rect 11165 -20314 11197 -20280
rect 11233 -20314 11267 -20280
rect 11303 -20314 11335 -20280
rect 11375 -20314 11403 -20280
rect 11447 -20314 11471 -20280
rect 11505 -20314 11544 -20280
rect 11974 -20314 12013 -20280
rect 12047 -20314 12071 -20280
rect 12115 -20314 12143 -20280
rect 12183 -20314 12215 -20280
rect 12251 -20314 12285 -20280
rect 12321 -20314 12353 -20280
rect 12393 -20314 12421 -20280
rect 12465 -20314 12489 -20280
rect 12523 -20314 12562 -20280
rect 12992 -20314 13031 -20280
rect 13065 -20314 13089 -20280
rect 13133 -20314 13161 -20280
rect 13201 -20314 13233 -20280
rect 13269 -20314 13303 -20280
rect 13339 -20314 13371 -20280
rect 13411 -20314 13439 -20280
rect 13483 -20314 13507 -20280
rect 13541 -20314 13580 -20280
rect 14010 -20314 14049 -20280
rect 14083 -20314 14107 -20280
rect 14151 -20314 14179 -20280
rect 14219 -20314 14251 -20280
rect 14287 -20314 14321 -20280
rect 14357 -20314 14389 -20280
rect 14429 -20314 14457 -20280
rect 14501 -20314 14525 -20280
rect 14559 -20314 14598 -20280
rect 15028 -20314 15067 -20280
rect 15101 -20314 15125 -20280
rect 15169 -20314 15197 -20280
rect 15237 -20314 15269 -20280
rect 15305 -20314 15339 -20280
rect 15375 -20314 15407 -20280
rect 15447 -20314 15475 -20280
rect 15519 -20314 15543 -20280
rect 15577 -20314 15616 -20280
rect 16046 -20314 16085 -20280
rect 16119 -20314 16143 -20280
rect 16187 -20314 16215 -20280
rect 16255 -20314 16287 -20280
rect 16323 -20314 16357 -20280
rect 16393 -20314 16425 -20280
rect 16465 -20314 16493 -20280
rect 16537 -20314 16561 -20280
rect 16595 -20314 16634 -20280
rect 17064 -20314 17103 -20280
rect 17137 -20314 17161 -20280
rect 17205 -20314 17233 -20280
rect 17273 -20314 17305 -20280
rect 17341 -20314 17375 -20280
rect 17411 -20314 17443 -20280
rect 17483 -20314 17511 -20280
rect 17555 -20314 17579 -20280
rect 17613 -20314 17652 -20280
rect 18082 -20314 18121 -20280
rect 18155 -20314 18179 -20280
rect 18223 -20314 18251 -20280
rect 18291 -20314 18323 -20280
rect 18359 -20314 18393 -20280
rect 18429 -20314 18461 -20280
rect 18501 -20314 18529 -20280
rect 18573 -20314 18597 -20280
rect 18631 -20314 18670 -20280
rect 19100 -20314 19139 -20280
rect 19173 -20314 19197 -20280
rect 19241 -20314 19269 -20280
rect 19309 -20314 19341 -20280
rect 19377 -20314 19411 -20280
rect 19447 -20314 19479 -20280
rect 19519 -20314 19547 -20280
rect 19591 -20314 19615 -20280
rect 19649 -20314 19688 -20280
rect 20118 -20314 20157 -20280
rect 20191 -20314 20215 -20280
rect 20259 -20314 20287 -20280
rect 20327 -20314 20359 -20280
rect 20395 -20314 20429 -20280
rect 20465 -20314 20497 -20280
rect 20537 -20314 20565 -20280
rect 20609 -20314 20633 -20280
rect 20667 -20314 20706 -20280
rect 21136 -20314 21175 -20280
rect 21209 -20314 21233 -20280
rect 21277 -20314 21305 -20280
rect 21345 -20314 21377 -20280
rect 21413 -20314 21447 -20280
rect 21483 -20314 21515 -20280
rect 21555 -20314 21583 -20280
rect 21627 -20314 21651 -20280
rect 21685 -20314 21724 -20280
rect 22154 -20314 22193 -20280
rect 22227 -20314 22251 -20280
rect 22295 -20314 22323 -20280
rect 22363 -20314 22395 -20280
rect 22431 -20314 22465 -20280
rect 22501 -20314 22533 -20280
rect 22573 -20314 22601 -20280
rect 22645 -20314 22669 -20280
rect 22703 -20314 22742 -20280
rect -12322 -20339 -12222 -20333
rect -12322 -20405 -12289 -20339
rect -12255 -20405 -12222 -20339
rect 24822 -20333 24855 -20271
rect 24889 -20333 24922 -20271
rect 24822 -20339 24922 -20333
rect -12322 -20407 -12222 -20405
rect -12322 -20441 -12289 -20407
rect -12255 -20441 -12222 -20407
rect -2252 -20416 -2215 -20382
rect -2181 -20416 -2144 -20382
rect -2034 -20416 -1997 -20382
rect -1963 -20416 -1926 -20382
rect -1816 -20416 -1779 -20382
rect -1745 -20416 -1708 -20382
rect -1598 -20416 -1561 -20382
rect -1527 -20416 -1490 -20382
rect -1380 -20416 -1343 -20382
rect -1309 -20416 -1272 -20382
rect -1162 -20416 -1125 -20382
rect -1091 -20416 -1054 -20382
rect -944 -20416 -907 -20382
rect -873 -20416 -836 -20382
rect -726 -20416 -689 -20382
rect -655 -20416 -618 -20382
rect -508 -20416 -471 -20382
rect -437 -20416 -400 -20382
rect -290 -20416 -253 -20382
rect -219 -20416 -182 -20382
rect 2580 -20383 2614 -20348
rect -12322 -20443 -12222 -20441
rect -12322 -20509 -12289 -20443
rect -12255 -20509 -12222 -20443
rect -12322 -20515 -12222 -20509
rect -12322 -20577 -12289 -20515
rect -12255 -20577 -12222 -20515
rect -12322 -20587 -12222 -20577
rect -12322 -20645 -12289 -20587
rect -12255 -20645 -12222 -20587
rect -12322 -20659 -12222 -20645
rect -2324 -20469 -2290 -20450
rect -2324 -20537 -2290 -20535
rect -2324 -20573 -2290 -20571
rect -2324 -20658 -2290 -20639
rect -2106 -20469 -2072 -20450
rect -2106 -20537 -2072 -20535
rect -2106 -20573 -2072 -20571
rect -2106 -20658 -2072 -20639
rect -1888 -20469 -1854 -20450
rect -1888 -20537 -1854 -20535
rect -1888 -20573 -1854 -20571
rect -1888 -20658 -1854 -20639
rect -1670 -20469 -1636 -20450
rect -1670 -20537 -1636 -20535
rect -1670 -20573 -1636 -20571
rect -1670 -20658 -1636 -20639
rect -1452 -20469 -1418 -20450
rect -1452 -20537 -1418 -20535
rect -1452 -20573 -1418 -20571
rect -1452 -20658 -1418 -20639
rect -1234 -20469 -1200 -20450
rect -1234 -20537 -1200 -20535
rect -1234 -20573 -1200 -20571
rect -1234 -20658 -1200 -20639
rect -1016 -20469 -982 -20450
rect -1016 -20537 -982 -20535
rect -1016 -20573 -982 -20571
rect -1016 -20658 -982 -20639
rect -798 -20469 -764 -20450
rect -798 -20537 -764 -20535
rect -798 -20573 -764 -20571
rect -798 -20658 -764 -20639
rect -580 -20469 -546 -20450
rect -580 -20537 -546 -20535
rect -580 -20573 -546 -20571
rect -580 -20658 -546 -20639
rect -362 -20469 -328 -20450
rect -362 -20537 -328 -20535
rect -362 -20573 -328 -20571
rect -362 -20658 -328 -20639
rect -144 -20469 -110 -20450
rect -144 -20537 -110 -20535
rect -144 -20573 -110 -20571
rect -144 -20658 -110 -20639
rect 2580 -20455 2614 -20431
rect 2580 -20527 2614 -20499
rect 2580 -20599 2614 -20567
rect -12322 -20713 -12289 -20659
rect -12255 -20713 -12222 -20659
rect 2580 -20669 2614 -20635
rect -12322 -20731 -12222 -20713
rect -2252 -20726 -2215 -20692
rect -2181 -20726 -2144 -20692
rect -2034 -20726 -1997 -20692
rect -1963 -20726 -1926 -20692
rect -1816 -20726 -1779 -20692
rect -1745 -20726 -1708 -20692
rect -1598 -20726 -1561 -20692
rect -1527 -20726 -1490 -20692
rect -1380 -20726 -1343 -20692
rect -1309 -20726 -1272 -20692
rect -1162 -20726 -1125 -20692
rect -1091 -20726 -1054 -20692
rect -944 -20726 -907 -20692
rect -873 -20726 -836 -20692
rect -726 -20726 -689 -20692
rect -655 -20726 -618 -20692
rect -508 -20726 -471 -20692
rect -437 -20726 -400 -20692
rect -290 -20726 -253 -20692
rect -219 -20726 -182 -20692
rect -12322 -20781 -12289 -20731
rect -12255 -20781 -12222 -20731
rect -12322 -20803 -12222 -20781
rect -12322 -20849 -12289 -20803
rect -12255 -20849 -12222 -20803
rect -12322 -20875 -12222 -20849
rect -12322 -20917 -12289 -20875
rect -12255 -20917 -12222 -20875
rect -12322 -20947 -12222 -20917
rect -12322 -20985 -12289 -20947
rect -12255 -20985 -12222 -20947
rect 2580 -20737 2614 -20705
rect 2580 -20805 2614 -20777
rect 2580 -20873 2614 -20849
rect 2580 -20956 2614 -20921
rect 3598 -20383 3632 -20348
rect 3598 -20455 3632 -20431
rect 3598 -20527 3632 -20499
rect 3598 -20599 3632 -20567
rect 3598 -20669 3632 -20635
rect 3598 -20737 3632 -20705
rect 3598 -20805 3632 -20777
rect 3598 -20873 3632 -20849
rect 3598 -20956 3632 -20921
rect 4616 -20383 4650 -20348
rect 4616 -20455 4650 -20431
rect 4616 -20527 4650 -20499
rect 4616 -20599 4650 -20567
rect 4616 -20669 4650 -20635
rect 4616 -20737 4650 -20705
rect 4616 -20805 4650 -20777
rect 4616 -20873 4650 -20849
rect 4616 -20956 4650 -20921
rect 5634 -20383 5668 -20348
rect 5634 -20455 5668 -20431
rect 5634 -20527 5668 -20499
rect 5634 -20599 5668 -20567
rect 5634 -20669 5668 -20635
rect 5634 -20737 5668 -20705
rect 5634 -20805 5668 -20777
rect 5634 -20873 5668 -20849
rect 5634 -20956 5668 -20921
rect 6652 -20383 6686 -20348
rect 6652 -20455 6686 -20431
rect 6652 -20527 6686 -20499
rect 6652 -20599 6686 -20567
rect 6652 -20669 6686 -20635
rect 6652 -20737 6686 -20705
rect 6652 -20805 6686 -20777
rect 6652 -20873 6686 -20849
rect 6652 -20956 6686 -20921
rect 7670 -20383 7704 -20348
rect 7670 -20455 7704 -20431
rect 7670 -20527 7704 -20499
rect 7670 -20599 7704 -20567
rect 7670 -20669 7704 -20635
rect 7670 -20737 7704 -20705
rect 7670 -20805 7704 -20777
rect 7670 -20873 7704 -20849
rect 7670 -20956 7704 -20921
rect 8688 -20383 8722 -20348
rect 8688 -20455 8722 -20431
rect 8688 -20527 8722 -20499
rect 8688 -20599 8722 -20567
rect 8688 -20669 8722 -20635
rect 8688 -20737 8722 -20705
rect 8688 -20805 8722 -20777
rect 8688 -20873 8722 -20849
rect 8688 -20956 8722 -20921
rect 9706 -20383 9740 -20348
rect 9706 -20455 9740 -20431
rect 9706 -20527 9740 -20499
rect 9706 -20599 9740 -20567
rect 9706 -20669 9740 -20635
rect 9706 -20737 9740 -20705
rect 9706 -20805 9740 -20777
rect 9706 -20873 9740 -20849
rect 9706 -20956 9740 -20921
rect 10724 -20383 10758 -20348
rect 10724 -20455 10758 -20431
rect 10724 -20527 10758 -20499
rect 10724 -20599 10758 -20567
rect 10724 -20669 10758 -20635
rect 10724 -20737 10758 -20705
rect 10724 -20805 10758 -20777
rect 10724 -20873 10758 -20849
rect 10724 -20956 10758 -20921
rect 11742 -20383 11776 -20348
rect 11742 -20455 11776 -20431
rect 11742 -20527 11776 -20499
rect 11742 -20599 11776 -20567
rect 11742 -20669 11776 -20635
rect 11742 -20737 11776 -20705
rect 11742 -20805 11776 -20777
rect 11742 -20873 11776 -20849
rect 11742 -20956 11776 -20921
rect 12760 -20383 12794 -20348
rect 12760 -20455 12794 -20431
rect 12760 -20527 12794 -20499
rect 12760 -20599 12794 -20567
rect 12760 -20669 12794 -20635
rect 12760 -20737 12794 -20705
rect 12760 -20805 12794 -20777
rect 12760 -20873 12794 -20849
rect 12760 -20956 12794 -20921
rect 13778 -20383 13812 -20348
rect 13778 -20455 13812 -20431
rect 13778 -20527 13812 -20499
rect 13778 -20599 13812 -20567
rect 13778 -20669 13812 -20635
rect 13778 -20737 13812 -20705
rect 13778 -20805 13812 -20777
rect 13778 -20873 13812 -20849
rect 13778 -20956 13812 -20921
rect 14796 -20383 14830 -20348
rect 14796 -20455 14830 -20431
rect 14796 -20527 14830 -20499
rect 14796 -20599 14830 -20567
rect 14796 -20669 14830 -20635
rect 14796 -20737 14830 -20705
rect 14796 -20805 14830 -20777
rect 14796 -20873 14830 -20849
rect 14796 -20956 14830 -20921
rect 15814 -20383 15848 -20348
rect 15814 -20455 15848 -20431
rect 15814 -20527 15848 -20499
rect 15814 -20599 15848 -20567
rect 15814 -20669 15848 -20635
rect 15814 -20737 15848 -20705
rect 15814 -20805 15848 -20777
rect 15814 -20873 15848 -20849
rect 15814 -20956 15848 -20921
rect 16832 -20383 16866 -20348
rect 16832 -20455 16866 -20431
rect 16832 -20527 16866 -20499
rect 16832 -20599 16866 -20567
rect 16832 -20669 16866 -20635
rect 16832 -20737 16866 -20705
rect 16832 -20805 16866 -20777
rect 16832 -20873 16866 -20849
rect 16832 -20956 16866 -20921
rect 17850 -20383 17884 -20348
rect 17850 -20455 17884 -20431
rect 17850 -20527 17884 -20499
rect 17850 -20599 17884 -20567
rect 17850 -20669 17884 -20635
rect 17850 -20737 17884 -20705
rect 17850 -20805 17884 -20777
rect 17850 -20873 17884 -20849
rect 17850 -20956 17884 -20921
rect 18868 -20383 18902 -20348
rect 18868 -20455 18902 -20431
rect 18868 -20527 18902 -20499
rect 18868 -20599 18902 -20567
rect 18868 -20669 18902 -20635
rect 18868 -20737 18902 -20705
rect 18868 -20805 18902 -20777
rect 18868 -20873 18902 -20849
rect 18868 -20956 18902 -20921
rect 19886 -20383 19920 -20348
rect 19886 -20455 19920 -20431
rect 19886 -20527 19920 -20499
rect 19886 -20599 19920 -20567
rect 19886 -20669 19920 -20635
rect 19886 -20737 19920 -20705
rect 19886 -20805 19920 -20777
rect 19886 -20873 19920 -20849
rect 19886 -20956 19920 -20921
rect 20904 -20383 20938 -20348
rect 20904 -20455 20938 -20431
rect 20904 -20527 20938 -20499
rect 20904 -20599 20938 -20567
rect 20904 -20669 20938 -20635
rect 20904 -20737 20938 -20705
rect 20904 -20805 20938 -20777
rect 20904 -20873 20938 -20849
rect 20904 -20956 20938 -20921
rect 21922 -20383 21956 -20348
rect 21922 -20455 21956 -20431
rect 21922 -20527 21956 -20499
rect 21922 -20599 21956 -20567
rect 21922 -20669 21956 -20635
rect 21922 -20737 21956 -20705
rect 21922 -20805 21956 -20777
rect 21922 -20873 21956 -20849
rect 21922 -20956 21956 -20921
rect 22940 -20383 22974 -20348
rect 22940 -20455 22974 -20431
rect 22940 -20527 22974 -20499
rect 22940 -20599 22974 -20567
rect 22940 -20669 22974 -20635
rect 22940 -20737 22974 -20705
rect 22940 -20805 22974 -20777
rect 22940 -20873 22974 -20849
rect 22940 -20956 22974 -20921
rect 24822 -20405 24855 -20339
rect 24889 -20405 24922 -20339
rect 24822 -20407 24922 -20405
rect 24822 -20441 24855 -20407
rect 24889 -20441 24922 -20407
rect 24822 -20443 24922 -20441
rect 24822 -20509 24855 -20443
rect 24889 -20509 24922 -20443
rect 24822 -20515 24922 -20509
rect 24822 -20577 24855 -20515
rect 24889 -20577 24922 -20515
rect 24822 -20587 24922 -20577
rect 24822 -20645 24855 -20587
rect 24889 -20645 24922 -20587
rect 24822 -20659 24922 -20645
rect 24822 -20713 24855 -20659
rect 24889 -20713 24922 -20659
rect 24822 -20731 24922 -20713
rect 24822 -20781 24855 -20731
rect 24889 -20781 24922 -20731
rect 24822 -20803 24922 -20781
rect 24822 -20849 24855 -20803
rect 24889 -20849 24922 -20803
rect 24822 -20875 24922 -20849
rect 24822 -20917 24855 -20875
rect 24889 -20917 24922 -20875
rect 24822 -20947 24922 -20917
rect -12322 -21019 -12222 -20985
rect 24822 -20985 24855 -20947
rect 24889 -20985 24922 -20947
rect 11230 -20990 11290 -20988
rect 13274 -20990 13334 -20986
rect 16312 -20990 16372 -20986
rect -12322 -21053 -12289 -21019
rect -12255 -21053 -12222 -21019
rect 2812 -21024 2851 -20990
rect 2885 -21024 2909 -20990
rect 2953 -21024 2981 -20990
rect 3021 -21024 3053 -20990
rect 3089 -21024 3123 -20990
rect 3159 -21024 3191 -20990
rect 3231 -21024 3259 -20990
rect 3303 -21024 3327 -20990
rect 3361 -21024 3400 -20990
rect 3830 -21024 3869 -20990
rect 3903 -21024 3927 -20990
rect 3971 -21024 3999 -20990
rect 4039 -21024 4071 -20990
rect 4107 -21024 4141 -20990
rect 4177 -21024 4209 -20990
rect 4249 -21024 4277 -20990
rect 4321 -21024 4345 -20990
rect 4379 -21024 4418 -20990
rect 4848 -21024 4887 -20990
rect 4921 -21024 4945 -20990
rect 4989 -21024 5017 -20990
rect 5057 -21024 5089 -20990
rect 5125 -21024 5159 -20990
rect 5195 -21024 5227 -20990
rect 5267 -21024 5295 -20990
rect 5339 -21024 5363 -20990
rect 5397 -21024 5436 -20990
rect 5866 -21024 5905 -20990
rect 5939 -21024 5963 -20990
rect 6007 -21024 6035 -20990
rect 6075 -21024 6107 -20990
rect 6143 -21024 6177 -20990
rect 6213 -21024 6245 -20990
rect 6285 -21024 6313 -20990
rect 6357 -21024 6381 -20990
rect 6415 -21024 6454 -20990
rect 6884 -21024 6923 -20990
rect 6957 -21024 6981 -20990
rect 7025 -21024 7053 -20990
rect 7093 -21024 7125 -20990
rect 7161 -21024 7195 -20990
rect 7231 -21024 7263 -20990
rect 7303 -21024 7331 -20990
rect 7375 -21024 7399 -20990
rect 7433 -21024 7472 -20990
rect 7902 -21024 7941 -20990
rect 7975 -21024 7999 -20990
rect 8043 -21024 8071 -20990
rect 8111 -21024 8143 -20990
rect 8179 -21024 8213 -20990
rect 8249 -21024 8281 -20990
rect 8321 -21024 8349 -20990
rect 8393 -21024 8417 -20990
rect 8451 -21024 8490 -20990
rect 8920 -21024 8959 -20990
rect 8993 -21024 9017 -20990
rect 9061 -21024 9089 -20990
rect 9129 -21024 9161 -20990
rect 9197 -21024 9231 -20990
rect 9267 -21024 9299 -20990
rect 9339 -21024 9367 -20990
rect 9411 -21024 9435 -20990
rect 9469 -21024 9508 -20990
rect 9938 -21024 9977 -20990
rect 10011 -21024 10035 -20990
rect 10079 -21024 10107 -20990
rect 10147 -21024 10179 -20990
rect 10215 -21024 10249 -20990
rect 10285 -21024 10317 -20990
rect 10357 -21024 10385 -20990
rect 10429 -21024 10453 -20990
rect 10487 -21024 10526 -20990
rect 10956 -21024 10995 -20990
rect 11029 -21024 11053 -20990
rect 11097 -21024 11125 -20990
rect 11165 -21024 11197 -20990
rect 11233 -21024 11267 -20990
rect 11303 -21024 11335 -20990
rect 11375 -21024 11403 -20990
rect 11447 -21024 11471 -20990
rect 11505 -21024 11544 -20990
rect 11974 -21024 12013 -20990
rect 12047 -21024 12071 -20990
rect 12115 -21024 12143 -20990
rect 12183 -21024 12215 -20990
rect 12251 -21024 12285 -20990
rect 12321 -21024 12353 -20990
rect 12393 -21024 12421 -20990
rect 12465 -21024 12489 -20990
rect 12523 -21024 12562 -20990
rect 12992 -21024 13031 -20990
rect 13065 -21024 13089 -20990
rect 13133 -21024 13161 -20990
rect 13201 -21024 13233 -20990
rect 13269 -21024 13303 -20990
rect 13339 -21024 13371 -20990
rect 13411 -21024 13439 -20990
rect 13483 -21024 13507 -20990
rect 13541 -21024 13580 -20990
rect 14010 -21024 14049 -20990
rect 14083 -21024 14107 -20990
rect 14151 -21024 14179 -20990
rect 14219 -21024 14251 -20990
rect 14287 -21024 14321 -20990
rect 14357 -21024 14389 -20990
rect 14429 -21024 14457 -20990
rect 14501 -21024 14525 -20990
rect 14559 -21024 14598 -20990
rect 15028 -21024 15067 -20990
rect 15101 -21024 15125 -20990
rect 15169 -21024 15197 -20990
rect 15237 -21024 15269 -20990
rect 15305 -21024 15339 -20990
rect 15375 -21024 15407 -20990
rect 15447 -21024 15475 -20990
rect 15519 -21024 15543 -20990
rect 15577 -21024 15616 -20990
rect 16046 -21024 16085 -20990
rect 16119 -21024 16143 -20990
rect 16187 -21024 16215 -20990
rect 16255 -21024 16287 -20990
rect 16323 -21024 16357 -20990
rect 16393 -21024 16425 -20990
rect 16465 -21024 16493 -20990
rect 16537 -21024 16561 -20990
rect 16595 -21024 16634 -20990
rect 17064 -21024 17103 -20990
rect 17137 -21024 17161 -20990
rect 17205 -21024 17233 -20990
rect 17273 -21024 17305 -20990
rect 17341 -21024 17375 -20990
rect 17411 -21024 17443 -20990
rect 17483 -21024 17511 -20990
rect 17555 -21024 17579 -20990
rect 17613 -21024 17652 -20990
rect 18082 -21024 18121 -20990
rect 18155 -21024 18179 -20990
rect 18223 -21024 18251 -20990
rect 18291 -21024 18323 -20990
rect 18359 -21024 18393 -20990
rect 18429 -21024 18461 -20990
rect 18501 -21024 18529 -20990
rect 18573 -21024 18597 -20990
rect 18631 -21024 18670 -20990
rect 19100 -21024 19139 -20990
rect 19173 -21024 19197 -20990
rect 19241 -21024 19269 -20990
rect 19309 -21024 19341 -20990
rect 19377 -21024 19411 -20990
rect 19447 -21024 19479 -20990
rect 19519 -21024 19547 -20990
rect 19591 -21024 19615 -20990
rect 19649 -21024 19688 -20990
rect 20118 -21024 20157 -20990
rect 20191 -21024 20215 -20990
rect 20259 -21024 20287 -20990
rect 20327 -21024 20359 -20990
rect 20395 -21024 20429 -20990
rect 20465 -21024 20497 -20990
rect 20537 -21024 20565 -20990
rect 20609 -21024 20633 -20990
rect 20667 -21024 20706 -20990
rect 21136 -21024 21175 -20990
rect 21209 -21024 21233 -20990
rect 21277 -21024 21305 -20990
rect 21345 -21024 21377 -20990
rect 21413 -21024 21447 -20990
rect 21483 -21024 21515 -20990
rect 21555 -21024 21583 -20990
rect 21627 -21024 21651 -20990
rect 21685 -21024 21724 -20990
rect 22154 -21024 22193 -20990
rect 22227 -21024 22251 -20990
rect 22295 -21024 22323 -20990
rect 22363 -21024 22395 -20990
rect 22431 -21024 22465 -20990
rect 22501 -21024 22533 -20990
rect 22573 -21024 22601 -20990
rect 22645 -21024 22669 -20990
rect 22703 -21024 22742 -20990
rect 24822 -21019 24922 -20985
rect -12322 -21087 -12222 -21053
rect -12322 -21125 -12289 -21087
rect -12255 -21125 -12222 -21087
rect -12322 -21155 -12222 -21125
rect -12322 -21197 -12289 -21155
rect -12255 -21197 -12222 -21155
rect -12322 -21223 -12222 -21197
rect -12322 -21269 -12289 -21223
rect -12255 -21269 -12222 -21223
rect -12322 -21291 -12222 -21269
rect -12322 -21341 -12289 -21291
rect -12255 -21341 -12222 -21291
rect -12322 -21359 -12222 -21341
rect -12322 -21413 -12289 -21359
rect -12255 -21413 -12222 -21359
rect -12322 -21427 -12222 -21413
rect -12322 -21485 -12289 -21427
rect -12255 -21485 -12222 -21427
rect -12322 -21495 -12222 -21485
rect -12322 -21557 -12289 -21495
rect -12255 -21557 -12222 -21495
rect 24822 -21053 24855 -21019
rect 24889 -21053 24922 -21019
rect 24822 -21087 24922 -21053
rect 24822 -21125 24855 -21087
rect 24889 -21125 24922 -21087
rect 24822 -21155 24922 -21125
rect 24822 -21197 24855 -21155
rect 24889 -21197 24922 -21155
rect 24822 -21223 24922 -21197
rect 24822 -21269 24855 -21223
rect 24889 -21269 24922 -21223
rect 24822 -21291 24922 -21269
rect 24822 -21341 24855 -21291
rect 24889 -21341 24922 -21291
rect 24822 -21359 24922 -21341
rect 24822 -21413 24855 -21359
rect 24889 -21413 24922 -21359
rect 24822 -21427 24922 -21413
rect 24822 -21485 24855 -21427
rect 24889 -21485 24922 -21427
rect 24822 -21495 24922 -21485
rect 2812 -21546 2851 -21512
rect 2885 -21546 2909 -21512
rect 2953 -21546 2981 -21512
rect 3021 -21546 3053 -21512
rect 3089 -21546 3123 -21512
rect 3159 -21546 3191 -21512
rect 3231 -21546 3259 -21512
rect 3303 -21546 3327 -21512
rect 3361 -21546 3400 -21512
rect 3830 -21546 3869 -21512
rect 3903 -21546 3927 -21512
rect 3971 -21546 3999 -21512
rect 4039 -21546 4071 -21512
rect 4107 -21546 4141 -21512
rect 4177 -21546 4209 -21512
rect 4249 -21546 4277 -21512
rect 4321 -21546 4345 -21512
rect 4379 -21546 4418 -21512
rect 4848 -21546 4887 -21512
rect 4921 -21546 4945 -21512
rect 4989 -21546 5017 -21512
rect 5057 -21546 5089 -21512
rect 5125 -21546 5159 -21512
rect 5195 -21546 5227 -21512
rect 5267 -21546 5295 -21512
rect 5339 -21546 5363 -21512
rect 5397 -21546 5436 -21512
rect 5866 -21546 5905 -21512
rect 5939 -21546 5963 -21512
rect 6007 -21546 6035 -21512
rect 6075 -21546 6107 -21512
rect 6143 -21546 6177 -21512
rect 6213 -21546 6245 -21512
rect 6285 -21546 6313 -21512
rect 6357 -21546 6381 -21512
rect 6415 -21546 6454 -21512
rect 6884 -21546 6923 -21512
rect 6957 -21546 6981 -21512
rect 7025 -21546 7053 -21512
rect 7093 -21546 7125 -21512
rect 7161 -21546 7195 -21512
rect 7231 -21546 7263 -21512
rect 7303 -21546 7331 -21512
rect 7375 -21546 7399 -21512
rect 7433 -21546 7472 -21512
rect 7902 -21546 7941 -21512
rect 7975 -21546 7999 -21512
rect 8043 -21546 8071 -21512
rect 8111 -21546 8143 -21512
rect 8179 -21546 8213 -21512
rect 8249 -21546 8281 -21512
rect 8321 -21546 8349 -21512
rect 8393 -21546 8417 -21512
rect 8451 -21546 8490 -21512
rect 8920 -21546 8959 -21512
rect 8993 -21546 9017 -21512
rect 9061 -21546 9089 -21512
rect 9129 -21546 9161 -21512
rect 9197 -21546 9231 -21512
rect 9267 -21546 9299 -21512
rect 9339 -21546 9367 -21512
rect 9411 -21546 9435 -21512
rect 9469 -21546 9508 -21512
rect 9938 -21546 9977 -21512
rect 10011 -21546 10035 -21512
rect 10079 -21546 10107 -21512
rect 10147 -21546 10179 -21512
rect 10215 -21546 10249 -21512
rect 10285 -21546 10317 -21512
rect 10357 -21546 10385 -21512
rect 10429 -21546 10453 -21512
rect 10487 -21546 10526 -21512
rect 10956 -21546 10995 -21512
rect 11029 -21546 11053 -21512
rect 11097 -21546 11125 -21512
rect 11165 -21546 11197 -21512
rect 11233 -21546 11267 -21512
rect 11303 -21546 11335 -21512
rect 11375 -21546 11403 -21512
rect 11447 -21546 11471 -21512
rect 11505 -21546 11544 -21512
rect 11974 -21546 12013 -21512
rect 12047 -21546 12071 -21512
rect 12115 -21546 12143 -21512
rect 12183 -21546 12215 -21512
rect 12251 -21546 12285 -21512
rect 12321 -21546 12353 -21512
rect 12393 -21546 12421 -21512
rect 12465 -21546 12489 -21512
rect 12523 -21546 12562 -21512
rect 12992 -21546 13031 -21512
rect 13065 -21546 13089 -21512
rect 13133 -21546 13161 -21512
rect 13201 -21546 13233 -21512
rect 13269 -21546 13303 -21512
rect 13339 -21546 13371 -21512
rect 13411 -21546 13439 -21512
rect 13483 -21546 13507 -21512
rect 13541 -21546 13580 -21512
rect 14010 -21546 14049 -21512
rect 14083 -21546 14107 -21512
rect 14151 -21546 14179 -21512
rect 14219 -21546 14251 -21512
rect 14287 -21546 14321 -21512
rect 14357 -21546 14389 -21512
rect 14429 -21546 14457 -21512
rect 14501 -21546 14525 -21512
rect 14559 -21546 14598 -21512
rect 15028 -21546 15067 -21512
rect 15101 -21546 15125 -21512
rect 15169 -21546 15197 -21512
rect 15237 -21546 15269 -21512
rect 15305 -21546 15339 -21512
rect 15375 -21546 15407 -21512
rect 15447 -21546 15475 -21512
rect 15519 -21546 15543 -21512
rect 15577 -21546 15616 -21512
rect 16046 -21546 16085 -21512
rect 16119 -21546 16143 -21512
rect 16187 -21546 16215 -21512
rect 16255 -21546 16287 -21512
rect 16323 -21546 16357 -21512
rect 16393 -21546 16425 -21512
rect 16465 -21546 16493 -21512
rect 16537 -21546 16561 -21512
rect 16595 -21546 16634 -21512
rect 17064 -21546 17103 -21512
rect 17137 -21546 17161 -21512
rect 17205 -21546 17233 -21512
rect 17273 -21546 17305 -21512
rect 17341 -21546 17375 -21512
rect 17411 -21546 17443 -21512
rect 17483 -21546 17511 -21512
rect 17555 -21546 17579 -21512
rect 17613 -21546 17652 -21512
rect 18082 -21546 18121 -21512
rect 18155 -21546 18179 -21512
rect 18223 -21546 18251 -21512
rect 18291 -21546 18323 -21512
rect 18359 -21546 18393 -21512
rect 18429 -21546 18461 -21512
rect 18501 -21546 18529 -21512
rect 18573 -21546 18597 -21512
rect 18631 -21546 18670 -21512
rect 19100 -21546 19139 -21512
rect 19173 -21546 19197 -21512
rect 19241 -21546 19269 -21512
rect 19309 -21546 19341 -21512
rect 19377 -21546 19411 -21512
rect 19447 -21546 19479 -21512
rect 19519 -21546 19547 -21512
rect 19591 -21546 19615 -21512
rect 19649 -21546 19688 -21512
rect 20118 -21546 20157 -21512
rect 20191 -21546 20215 -21512
rect 20259 -21546 20287 -21512
rect 20327 -21546 20359 -21512
rect 20395 -21546 20429 -21512
rect 20465 -21546 20497 -21512
rect 20537 -21546 20565 -21512
rect 20609 -21546 20633 -21512
rect 20667 -21546 20706 -21512
rect 21136 -21546 21175 -21512
rect 21209 -21546 21233 -21512
rect 21277 -21546 21305 -21512
rect 21345 -21546 21377 -21512
rect 21413 -21546 21447 -21512
rect 21483 -21546 21515 -21512
rect 21555 -21546 21583 -21512
rect 21627 -21546 21651 -21512
rect 21685 -21546 21724 -21512
rect 22154 -21546 22193 -21512
rect 22227 -21546 22251 -21512
rect 22295 -21546 22323 -21512
rect 22363 -21546 22395 -21512
rect 22431 -21546 22465 -21512
rect 22501 -21546 22533 -21512
rect 22573 -21546 22601 -21512
rect 22645 -21546 22669 -21512
rect 22703 -21546 22742 -21512
rect 6134 -21548 6194 -21546
rect -12322 -21563 -12222 -21557
rect -12322 -21629 -12289 -21563
rect -12255 -21629 -12222 -21563
rect 24822 -21557 24855 -21495
rect 24889 -21557 24922 -21495
rect 24822 -21563 24922 -21557
rect -12322 -21631 -12222 -21629
rect -12322 -21665 -12289 -21631
rect -12255 -21665 -12222 -21631
rect -12322 -21667 -12222 -21665
rect -12322 -21733 -12289 -21667
rect -12255 -21733 -12222 -21667
rect 2580 -21615 2614 -21580
rect 2580 -21687 2614 -21663
rect -12322 -21739 -12222 -21733
rect -12322 -21801 -12289 -21739
rect -12255 -21801 -12222 -21739
rect -9173 -21743 -9134 -21709
rect -9100 -21743 -9076 -21709
rect -9032 -21743 -9004 -21709
rect -8964 -21743 -8932 -21709
rect -8896 -21743 -8862 -21709
rect -8826 -21743 -8794 -21709
rect -8754 -21743 -8726 -21709
rect -8682 -21743 -8658 -21709
rect -8624 -21743 -8585 -21709
rect -8155 -21743 -8116 -21709
rect -8082 -21743 -8058 -21709
rect -8014 -21743 -7986 -21709
rect -7946 -21743 -7914 -21709
rect -7878 -21743 -7844 -21709
rect -7808 -21743 -7776 -21709
rect -7736 -21743 -7708 -21709
rect -7664 -21743 -7640 -21709
rect -7606 -21743 -7567 -21709
rect -7137 -21743 -7098 -21709
rect -7064 -21743 -7040 -21709
rect -6996 -21743 -6968 -21709
rect -6928 -21743 -6896 -21709
rect -6860 -21743 -6826 -21709
rect -6790 -21743 -6758 -21709
rect -6718 -21743 -6690 -21709
rect -6646 -21743 -6622 -21709
rect -6588 -21743 -6549 -21709
rect -6119 -21743 -6080 -21709
rect -6046 -21743 -6022 -21709
rect -5978 -21743 -5950 -21709
rect -5910 -21743 -5878 -21709
rect -5842 -21743 -5808 -21709
rect -5772 -21743 -5740 -21709
rect -5700 -21743 -5672 -21709
rect -5628 -21743 -5604 -21709
rect -5570 -21743 -5531 -21709
rect -5101 -21743 -5062 -21709
rect -5028 -21743 -5004 -21709
rect -4960 -21743 -4932 -21709
rect -4892 -21743 -4860 -21709
rect -4824 -21743 -4790 -21709
rect -4754 -21743 -4722 -21709
rect -4682 -21743 -4654 -21709
rect -4610 -21743 -4586 -21709
rect -4552 -21743 -4513 -21709
rect -4083 -21743 -4044 -21709
rect -4010 -21743 -3986 -21709
rect -3942 -21743 -3914 -21709
rect -3874 -21743 -3842 -21709
rect -3806 -21743 -3772 -21709
rect -3736 -21743 -3704 -21709
rect -3664 -21743 -3636 -21709
rect -3592 -21743 -3568 -21709
rect -3534 -21743 -3495 -21709
rect -2322 -21742 -2295 -21708
rect -2193 -21742 -2166 -21708
rect -2024 -21742 -1997 -21708
rect -1895 -21742 -1868 -21708
rect -1726 -21742 -1699 -21708
rect -1597 -21742 -1570 -21708
rect -1428 -21742 -1401 -21708
rect -1299 -21742 -1272 -21708
rect -1130 -21742 -1103 -21708
rect -1001 -21742 -974 -21708
rect -832 -21742 -805 -21708
rect -703 -21742 -676 -21708
rect -534 -21742 -507 -21708
rect -405 -21742 -378 -21708
rect -236 -21742 -209 -21708
rect -107 -21742 -80 -21708
rect 62 -21742 89 -21708
rect 191 -21742 218 -21708
rect 360 -21742 387 -21708
rect 489 -21742 516 -21708
rect 658 -21742 685 -21708
rect 787 -21742 814 -21708
rect 2580 -21759 2614 -21731
rect -12322 -21811 -12222 -21801
rect -12322 -21869 -12289 -21811
rect -12255 -21869 -12222 -21811
rect -12322 -21883 -12222 -21869
rect -12322 -21937 -12289 -21883
rect -12255 -21937 -12222 -21883
rect -12322 -21955 -12222 -21937
rect -12322 -22005 -12289 -21955
rect -12255 -22005 -12222 -21955
rect -12322 -22027 -12222 -22005
rect -12322 -22073 -12289 -22027
rect -12255 -22073 -12222 -22027
rect -12322 -22099 -12222 -22073
rect -12322 -22141 -12289 -22099
rect -12255 -22141 -12222 -22099
rect -12322 -22171 -12222 -22141
rect -12322 -22209 -12289 -22171
rect -12255 -22209 -12222 -22171
rect -12322 -22243 -12222 -22209
rect -12322 -22277 -12289 -22243
rect -12255 -22277 -12222 -22243
rect -12322 -22311 -12222 -22277
rect -12322 -22349 -12289 -22311
rect -12255 -22349 -12222 -22311
rect -12322 -22379 -12222 -22349
rect -12322 -22421 -12289 -22379
rect -12255 -22421 -12222 -22379
rect -9405 -21812 -9371 -21777
rect -9405 -21884 -9371 -21860
rect -9405 -21956 -9371 -21928
rect -9405 -22028 -9371 -21996
rect -9405 -22098 -9371 -22064
rect -9405 -22166 -9371 -22134
rect -9405 -22234 -9371 -22206
rect -9405 -22302 -9371 -22278
rect -9405 -22385 -9371 -22350
rect -8387 -21812 -8353 -21777
rect -8387 -21884 -8353 -21860
rect -8387 -21956 -8353 -21928
rect -8387 -22028 -8353 -21996
rect -8387 -22098 -8353 -22064
rect -8387 -22166 -8353 -22134
rect -8387 -22234 -8353 -22206
rect -8387 -22302 -8353 -22278
rect -8387 -22385 -8353 -22350
rect -7369 -21812 -7335 -21777
rect -7369 -21884 -7335 -21860
rect -7369 -21956 -7335 -21928
rect -7369 -22028 -7335 -21996
rect -7369 -22098 -7335 -22064
rect -7369 -22166 -7335 -22134
rect -7369 -22234 -7335 -22206
rect -7369 -22302 -7335 -22278
rect -7369 -22385 -7335 -22350
rect -6351 -21812 -6317 -21777
rect -6351 -21884 -6317 -21860
rect -6351 -21956 -6317 -21928
rect -6351 -22028 -6317 -21996
rect -6351 -22098 -6317 -22064
rect -6351 -22166 -6317 -22134
rect -6351 -22234 -6317 -22206
rect -6351 -22302 -6317 -22278
rect -6351 -22385 -6317 -22350
rect -5333 -21812 -5299 -21777
rect -5333 -21884 -5299 -21860
rect -5333 -21956 -5299 -21928
rect -5333 -22028 -5299 -21996
rect -5333 -22098 -5299 -22064
rect -5333 -22166 -5299 -22134
rect -5333 -22234 -5299 -22206
rect -5333 -22302 -5299 -22278
rect -5333 -22385 -5299 -22350
rect -4315 -21812 -4281 -21777
rect -4315 -21884 -4281 -21860
rect -4315 -21956 -4281 -21928
rect -4315 -22028 -4281 -21996
rect -4315 -22098 -4281 -22064
rect -4315 -22166 -4281 -22134
rect -4315 -22234 -4281 -22206
rect -4315 -22302 -4281 -22278
rect -4315 -22385 -4281 -22350
rect -3297 -21812 -3263 -21777
rect -3297 -21884 -3263 -21860
rect -3297 -21956 -3263 -21928
rect -3297 -22028 -3263 -21996
rect -3297 -22098 -3263 -22064
rect -3297 -22166 -3263 -22134
rect -3297 -22234 -3263 -22206
rect -3297 -22302 -3263 -22278
rect -3297 -22385 -3263 -22350
rect -2410 -21811 -2376 -21776
rect -2410 -21883 -2376 -21859
rect -2410 -21955 -2376 -21927
rect -2410 -22027 -2376 -21995
rect -2410 -22097 -2376 -22063
rect -2410 -22165 -2376 -22133
rect -2410 -22233 -2376 -22205
rect -2410 -22301 -2376 -22277
rect -2410 -22384 -2376 -22349
rect -2112 -21811 -2078 -21776
rect -2112 -21883 -2078 -21859
rect -2112 -21955 -2078 -21927
rect -2112 -22027 -2078 -21995
rect -2112 -22097 -2078 -22063
rect -2112 -22165 -2078 -22133
rect -2112 -22233 -2078 -22205
rect -2112 -22301 -2078 -22277
rect -2112 -22384 -2078 -22349
rect -1814 -21811 -1780 -21776
rect -1814 -21883 -1780 -21859
rect -1814 -21955 -1780 -21927
rect -1814 -22027 -1780 -21995
rect -1814 -22097 -1780 -22063
rect -1814 -22165 -1780 -22133
rect -1814 -22233 -1780 -22205
rect -1814 -22301 -1780 -22277
rect -1814 -22384 -1780 -22349
rect -1516 -21811 -1482 -21776
rect -1516 -21883 -1482 -21859
rect -1516 -21955 -1482 -21927
rect -1516 -22027 -1482 -21995
rect -1516 -22097 -1482 -22063
rect -1516 -22165 -1482 -22133
rect -1516 -22233 -1482 -22205
rect -1516 -22301 -1482 -22277
rect -1516 -22384 -1482 -22349
rect -1218 -21811 -1184 -21776
rect -1218 -21883 -1184 -21859
rect -1218 -21955 -1184 -21927
rect -1218 -22027 -1184 -21995
rect -1218 -22097 -1184 -22063
rect -1218 -22165 -1184 -22133
rect -1218 -22233 -1184 -22205
rect -1218 -22301 -1184 -22277
rect -1218 -22384 -1184 -22349
rect -920 -21811 -886 -21776
rect -920 -21883 -886 -21859
rect -920 -21955 -886 -21927
rect -920 -22027 -886 -21995
rect -920 -22097 -886 -22063
rect -920 -22165 -886 -22133
rect -920 -22233 -886 -22205
rect -920 -22301 -886 -22277
rect -920 -22384 -886 -22349
rect -622 -21811 -588 -21776
rect -622 -21883 -588 -21859
rect -622 -21955 -588 -21927
rect -622 -22027 -588 -21995
rect -622 -22097 -588 -22063
rect -622 -22165 -588 -22133
rect -622 -22233 -588 -22205
rect -622 -22301 -588 -22277
rect -622 -22384 -588 -22349
rect -324 -21811 -290 -21776
rect -324 -21883 -290 -21859
rect -324 -21955 -290 -21927
rect -324 -22027 -290 -21995
rect -324 -22097 -290 -22063
rect -324 -22165 -290 -22133
rect -324 -22233 -290 -22205
rect -324 -22301 -290 -22277
rect -324 -22384 -290 -22349
rect -26 -21811 8 -21776
rect -26 -21883 8 -21859
rect -26 -21955 8 -21927
rect -26 -22027 8 -21995
rect -26 -22097 8 -22063
rect -26 -22165 8 -22133
rect -26 -22233 8 -22205
rect -26 -22301 8 -22277
rect -26 -22384 8 -22349
rect 272 -21811 306 -21776
rect 272 -21883 306 -21859
rect 272 -21955 306 -21927
rect 272 -22027 306 -21995
rect 272 -22097 306 -22063
rect 272 -22165 306 -22133
rect 272 -22233 306 -22205
rect 272 -22301 306 -22277
rect 272 -22384 306 -22349
rect 570 -21811 604 -21776
rect 570 -21883 604 -21859
rect 570 -21955 604 -21927
rect 570 -22027 604 -21995
rect 570 -22097 604 -22063
rect 570 -22165 604 -22133
rect 570 -22233 604 -22205
rect 570 -22301 604 -22277
rect 570 -22384 604 -22349
rect 868 -21811 902 -21776
rect 868 -21883 902 -21859
rect 868 -21955 902 -21927
rect 868 -22027 902 -21995
rect 868 -22097 902 -22063
rect 868 -22165 902 -22133
rect 2580 -21831 2614 -21799
rect 2580 -21901 2614 -21867
rect 2580 -21969 2614 -21937
rect 2580 -22037 2614 -22009
rect 2580 -22105 2614 -22081
rect 2580 -22188 2614 -22153
rect 3598 -21615 3632 -21580
rect 3598 -21687 3632 -21663
rect 3598 -21759 3632 -21731
rect 3598 -21831 3632 -21799
rect 3598 -21901 3632 -21867
rect 3598 -21969 3632 -21937
rect 3598 -22037 3632 -22009
rect 3598 -22105 3632 -22081
rect 3598 -22188 3632 -22153
rect 4616 -21615 4650 -21580
rect 4616 -21687 4650 -21663
rect 4616 -21759 4650 -21731
rect 4616 -21831 4650 -21799
rect 4616 -21901 4650 -21867
rect 4616 -21969 4650 -21937
rect 4616 -22037 4650 -22009
rect 4616 -22105 4650 -22081
rect 4616 -22188 4650 -22153
rect 5634 -21615 5668 -21580
rect 5634 -21687 5668 -21663
rect 5634 -21759 5668 -21731
rect 5634 -21831 5668 -21799
rect 5634 -21901 5668 -21867
rect 5634 -21969 5668 -21937
rect 5634 -22037 5668 -22009
rect 5634 -22105 5668 -22081
rect 5634 -22188 5668 -22153
rect 6652 -21615 6686 -21580
rect 6652 -21687 6686 -21663
rect 6652 -21759 6686 -21731
rect 6652 -21831 6686 -21799
rect 6652 -21901 6686 -21867
rect 6652 -21969 6686 -21937
rect 6652 -22037 6686 -22009
rect 6652 -22105 6686 -22081
rect 6652 -22188 6686 -22153
rect 7670 -21615 7704 -21580
rect 7670 -21687 7704 -21663
rect 7670 -21759 7704 -21731
rect 7670 -21831 7704 -21799
rect 7670 -21901 7704 -21867
rect 7670 -21969 7704 -21937
rect 7670 -22037 7704 -22009
rect 7670 -22105 7704 -22081
rect 7670 -22188 7704 -22153
rect 8688 -21615 8722 -21580
rect 8688 -21687 8722 -21663
rect 8688 -21759 8722 -21731
rect 8688 -21831 8722 -21799
rect 8688 -21901 8722 -21867
rect 8688 -21969 8722 -21937
rect 8688 -22037 8722 -22009
rect 8688 -22105 8722 -22081
rect 8688 -22188 8722 -22153
rect 9706 -21615 9740 -21580
rect 9706 -21687 9740 -21663
rect 9706 -21759 9740 -21731
rect 9706 -21831 9740 -21799
rect 9706 -21901 9740 -21867
rect 9706 -21969 9740 -21937
rect 9706 -22037 9740 -22009
rect 9706 -22105 9740 -22081
rect 9706 -22188 9740 -22153
rect 10724 -21615 10758 -21580
rect 10724 -21687 10758 -21663
rect 10724 -21759 10758 -21731
rect 10724 -21831 10758 -21799
rect 10724 -21901 10758 -21867
rect 10724 -21969 10758 -21937
rect 10724 -22037 10758 -22009
rect 10724 -22105 10758 -22081
rect 10724 -22188 10758 -22153
rect 11742 -21615 11776 -21580
rect 11742 -21687 11776 -21663
rect 11742 -21759 11776 -21731
rect 11742 -21831 11776 -21799
rect 11742 -21901 11776 -21867
rect 11742 -21969 11776 -21937
rect 11742 -22037 11776 -22009
rect 11742 -22105 11776 -22081
rect 11742 -22188 11776 -22153
rect 12760 -21615 12794 -21580
rect 12760 -21687 12794 -21663
rect 12760 -21759 12794 -21731
rect 12760 -21831 12794 -21799
rect 12760 -21901 12794 -21867
rect 12760 -21969 12794 -21937
rect 12760 -22037 12794 -22009
rect 12760 -22105 12794 -22081
rect 12760 -22188 12794 -22153
rect 13778 -21615 13812 -21580
rect 13778 -21687 13812 -21663
rect 13778 -21759 13812 -21731
rect 13778 -21831 13812 -21799
rect 13778 -21901 13812 -21867
rect 13778 -21969 13812 -21937
rect 13778 -22037 13812 -22009
rect 13778 -22105 13812 -22081
rect 13778 -22188 13812 -22153
rect 14796 -21615 14830 -21580
rect 14796 -21687 14830 -21663
rect 14796 -21759 14830 -21731
rect 14796 -21831 14830 -21799
rect 14796 -21901 14830 -21867
rect 14796 -21969 14830 -21937
rect 14796 -22037 14830 -22009
rect 14796 -22105 14830 -22081
rect 14796 -22188 14830 -22153
rect 15814 -21615 15848 -21580
rect 15814 -21687 15848 -21663
rect 15814 -21759 15848 -21731
rect 15814 -21831 15848 -21799
rect 15814 -21901 15848 -21867
rect 15814 -21969 15848 -21937
rect 15814 -22037 15848 -22009
rect 15814 -22105 15848 -22081
rect 15814 -22188 15848 -22153
rect 16832 -21615 16866 -21580
rect 16832 -21687 16866 -21663
rect 16832 -21759 16866 -21731
rect 16832 -21831 16866 -21799
rect 16832 -21901 16866 -21867
rect 16832 -21969 16866 -21937
rect 16832 -22037 16866 -22009
rect 16832 -22105 16866 -22081
rect 16832 -22188 16866 -22153
rect 17850 -21615 17884 -21580
rect 17850 -21687 17884 -21663
rect 17850 -21759 17884 -21731
rect 17850 -21831 17884 -21799
rect 17850 -21901 17884 -21867
rect 17850 -21969 17884 -21937
rect 17850 -22037 17884 -22009
rect 17850 -22105 17884 -22081
rect 17850 -22188 17884 -22153
rect 18868 -21615 18902 -21580
rect 18868 -21687 18902 -21663
rect 18868 -21759 18902 -21731
rect 18868 -21831 18902 -21799
rect 18868 -21901 18902 -21867
rect 18868 -21969 18902 -21937
rect 18868 -22037 18902 -22009
rect 18868 -22105 18902 -22081
rect 18868 -22188 18902 -22153
rect 19886 -21615 19920 -21580
rect 19886 -21687 19920 -21663
rect 19886 -21759 19920 -21731
rect 19886 -21831 19920 -21799
rect 19886 -21901 19920 -21867
rect 19886 -21969 19920 -21937
rect 19886 -22037 19920 -22009
rect 19886 -22105 19920 -22081
rect 19886 -22188 19920 -22153
rect 20904 -21615 20938 -21580
rect 20904 -21687 20938 -21663
rect 20904 -21759 20938 -21731
rect 20904 -21831 20938 -21799
rect 20904 -21901 20938 -21867
rect 20904 -21969 20938 -21937
rect 20904 -22037 20938 -22009
rect 20904 -22105 20938 -22081
rect 20904 -22188 20938 -22153
rect 21922 -21615 21956 -21580
rect 21922 -21687 21956 -21663
rect 21922 -21759 21956 -21731
rect 21922 -21831 21956 -21799
rect 21922 -21901 21956 -21867
rect 21922 -21969 21956 -21937
rect 21922 -22037 21956 -22009
rect 21922 -22105 21956 -22081
rect 21922 -22172 21956 -22153
rect 22940 -21615 22974 -21580
rect 22940 -21687 22974 -21663
rect 22940 -21759 22974 -21731
rect 22940 -21831 22974 -21799
rect 22940 -21901 22974 -21867
rect 22940 -21969 22974 -21937
rect 22940 -22037 22974 -22009
rect 22940 -22105 22974 -22081
rect 22940 -22188 22974 -22153
rect 24822 -21629 24855 -21563
rect 24889 -21629 24922 -21563
rect 24822 -21631 24922 -21629
rect 24822 -21665 24855 -21631
rect 24889 -21665 24922 -21631
rect 24822 -21667 24922 -21665
rect 24822 -21733 24855 -21667
rect 24889 -21733 24922 -21667
rect 24822 -21739 24922 -21733
rect 24822 -21801 24855 -21739
rect 24889 -21801 24922 -21739
rect 24822 -21811 24922 -21801
rect 24822 -21869 24855 -21811
rect 24889 -21869 24922 -21811
rect 24822 -21883 24922 -21869
rect 24822 -21937 24855 -21883
rect 24889 -21937 24922 -21883
rect 24822 -21955 24922 -21937
rect 24822 -22005 24855 -21955
rect 24889 -22005 24922 -21955
rect 24822 -22027 24922 -22005
rect 24822 -22073 24855 -22027
rect 24889 -22073 24922 -22027
rect 24822 -22099 24922 -22073
rect 24822 -22141 24855 -22099
rect 24889 -22141 24922 -22099
rect 24822 -22171 24922 -22141
rect 868 -22233 902 -22205
rect 24822 -22209 24855 -22171
rect 24889 -22209 24922 -22171
rect 10206 -22222 10266 -22212
rect 2812 -22256 2851 -22222
rect 2885 -22256 2909 -22222
rect 2953 -22256 2981 -22222
rect 3021 -22256 3053 -22222
rect 3089 -22256 3123 -22222
rect 3159 -22256 3191 -22222
rect 3231 -22256 3259 -22222
rect 3303 -22256 3327 -22222
rect 3361 -22256 3400 -22222
rect 3830 -22256 3869 -22222
rect 3903 -22256 3927 -22222
rect 3971 -22256 3999 -22222
rect 4039 -22256 4071 -22222
rect 4107 -22256 4141 -22222
rect 4177 -22256 4209 -22222
rect 4249 -22256 4277 -22222
rect 4321 -22256 4345 -22222
rect 4379 -22256 4418 -22222
rect 4848 -22256 4887 -22222
rect 4921 -22256 4945 -22222
rect 4989 -22256 5017 -22222
rect 5057 -22256 5089 -22222
rect 5125 -22256 5159 -22222
rect 5195 -22256 5227 -22222
rect 5267 -22256 5295 -22222
rect 5339 -22256 5363 -22222
rect 5397 -22256 5436 -22222
rect 5866 -22256 5905 -22222
rect 5939 -22256 5963 -22222
rect 6007 -22256 6035 -22222
rect 6075 -22256 6107 -22222
rect 6143 -22256 6177 -22222
rect 6213 -22256 6245 -22222
rect 6285 -22256 6313 -22222
rect 6357 -22256 6381 -22222
rect 6415 -22256 6454 -22222
rect 6884 -22256 6923 -22222
rect 6957 -22256 6981 -22222
rect 7025 -22256 7053 -22222
rect 7093 -22256 7125 -22222
rect 7161 -22256 7195 -22222
rect 7231 -22256 7263 -22222
rect 7303 -22256 7331 -22222
rect 7375 -22256 7399 -22222
rect 7433 -22256 7472 -22222
rect 7902 -22256 7941 -22222
rect 7975 -22256 7999 -22222
rect 8043 -22256 8071 -22222
rect 8111 -22256 8143 -22222
rect 8179 -22256 8213 -22222
rect 8249 -22256 8281 -22222
rect 8321 -22256 8349 -22222
rect 8393 -22256 8417 -22222
rect 8451 -22256 8490 -22222
rect 8920 -22256 8959 -22222
rect 8993 -22256 9017 -22222
rect 9061 -22256 9089 -22222
rect 9129 -22256 9161 -22222
rect 9197 -22256 9231 -22222
rect 9267 -22256 9299 -22222
rect 9339 -22256 9367 -22222
rect 9411 -22256 9435 -22222
rect 9469 -22256 9508 -22222
rect 9938 -22256 9977 -22222
rect 10011 -22256 10035 -22222
rect 10079 -22256 10107 -22222
rect 10147 -22256 10179 -22222
rect 10215 -22256 10249 -22222
rect 10285 -22256 10317 -22222
rect 10357 -22256 10385 -22222
rect 10429 -22256 10453 -22222
rect 10487 -22256 10526 -22222
rect 10956 -22256 10995 -22222
rect 11029 -22256 11053 -22222
rect 11097 -22256 11125 -22222
rect 11165 -22256 11197 -22222
rect 11233 -22256 11267 -22222
rect 11303 -22256 11335 -22222
rect 11375 -22256 11403 -22222
rect 11447 -22256 11471 -22222
rect 11505 -22256 11544 -22222
rect 11974 -22256 12013 -22222
rect 12047 -22256 12071 -22222
rect 12115 -22256 12143 -22222
rect 12183 -22256 12215 -22222
rect 12251 -22256 12285 -22222
rect 12321 -22256 12353 -22222
rect 12393 -22256 12421 -22222
rect 12465 -22256 12489 -22222
rect 12523 -22256 12562 -22222
rect 12992 -22256 13031 -22222
rect 13065 -22256 13089 -22222
rect 13133 -22256 13161 -22222
rect 13201 -22256 13233 -22222
rect 13269 -22256 13303 -22222
rect 13339 -22256 13371 -22222
rect 13411 -22256 13439 -22222
rect 13483 -22256 13507 -22222
rect 13541 -22256 13580 -22222
rect 14010 -22256 14049 -22222
rect 14083 -22256 14107 -22222
rect 14151 -22256 14179 -22222
rect 14219 -22256 14251 -22222
rect 14287 -22256 14321 -22222
rect 14357 -22256 14389 -22222
rect 14429 -22256 14457 -22222
rect 14501 -22256 14525 -22222
rect 14559 -22256 14598 -22222
rect 15028 -22256 15067 -22222
rect 15101 -22256 15125 -22222
rect 15169 -22256 15197 -22222
rect 15237 -22256 15269 -22222
rect 15305 -22256 15339 -22222
rect 15375 -22256 15407 -22222
rect 15447 -22256 15475 -22222
rect 15519 -22256 15543 -22222
rect 15577 -22256 15616 -22222
rect 16046 -22256 16085 -22222
rect 16119 -22256 16143 -22222
rect 16187 -22256 16215 -22222
rect 16255 -22256 16287 -22222
rect 16323 -22256 16357 -22222
rect 16393 -22256 16425 -22222
rect 16465 -22256 16493 -22222
rect 16537 -22256 16561 -22222
rect 16595 -22256 16634 -22222
rect 17064 -22256 17103 -22222
rect 17137 -22256 17161 -22222
rect 17205 -22256 17233 -22222
rect 17273 -22256 17305 -22222
rect 17341 -22256 17375 -22222
rect 17411 -22256 17443 -22222
rect 17483 -22256 17511 -22222
rect 17555 -22256 17579 -22222
rect 17613 -22256 17652 -22222
rect 18082 -22256 18121 -22222
rect 18155 -22256 18179 -22222
rect 18223 -22256 18251 -22222
rect 18291 -22256 18323 -22222
rect 18359 -22256 18393 -22222
rect 18429 -22256 18461 -22222
rect 18501 -22256 18529 -22222
rect 18573 -22256 18597 -22222
rect 18631 -22256 18670 -22222
rect 19100 -22256 19139 -22222
rect 19173 -22256 19197 -22222
rect 19241 -22256 19269 -22222
rect 19309 -22256 19341 -22222
rect 19377 -22256 19411 -22222
rect 19447 -22256 19479 -22222
rect 19519 -22256 19547 -22222
rect 19591 -22256 19615 -22222
rect 19649 -22256 19688 -22222
rect 20118 -22256 20157 -22222
rect 20191 -22256 20215 -22222
rect 20259 -22256 20287 -22222
rect 20327 -22256 20359 -22222
rect 20395 -22256 20429 -22222
rect 20465 -22256 20497 -22222
rect 20537 -22256 20565 -22222
rect 20609 -22256 20633 -22222
rect 20667 -22256 20706 -22222
rect 21136 -22256 21175 -22222
rect 21209 -22256 21233 -22222
rect 21277 -22256 21305 -22222
rect 21345 -22256 21379 -22222
rect 21413 -22256 21447 -22222
rect 21481 -22256 21515 -22222
rect 21555 -22256 21583 -22222
rect 21627 -22256 21651 -22222
rect 21685 -22256 21724 -22222
rect 22154 -22256 22193 -22222
rect 22227 -22256 22251 -22222
rect 22295 -22256 22323 -22222
rect 22363 -22256 22395 -22222
rect 22431 -22256 22465 -22222
rect 22501 -22256 22533 -22222
rect 22573 -22256 22601 -22222
rect 22645 -22256 22669 -22222
rect 22703 -22256 22742 -22222
rect 24822 -22243 24922 -22209
rect 868 -22301 902 -22277
rect 868 -22384 902 -22349
rect 24822 -22277 24855 -22243
rect 24889 -22277 24922 -22243
rect 24822 -22311 24922 -22277
rect 24822 -22349 24855 -22311
rect 24889 -22349 24922 -22311
rect 24822 -22379 24922 -22349
rect -7892 -22419 -7832 -22418
rect -6882 -22419 -6822 -22418
rect -4834 -22419 -4774 -22418
rect -12322 -22447 -12222 -22421
rect -12322 -22493 -12289 -22447
rect -12255 -22493 -12222 -22447
rect -9173 -22453 -9134 -22419
rect -9100 -22453 -9076 -22419
rect -9032 -22453 -9004 -22419
rect -8964 -22453 -8932 -22419
rect -8896 -22453 -8862 -22419
rect -8826 -22453 -8794 -22419
rect -8754 -22453 -8726 -22419
rect -8682 -22453 -8658 -22419
rect -8624 -22453 -8585 -22419
rect -8155 -22453 -8116 -22419
rect -8082 -22453 -8058 -22419
rect -8014 -22453 -7986 -22419
rect -7946 -22453 -7914 -22419
rect -7878 -22453 -7844 -22419
rect -7808 -22453 -7776 -22419
rect -7736 -22453 -7708 -22419
rect -7664 -22453 -7640 -22419
rect -7606 -22453 -7567 -22419
rect -7137 -22453 -7098 -22419
rect -7064 -22453 -7040 -22419
rect -6996 -22453 -6968 -22419
rect -6928 -22453 -6896 -22419
rect -6860 -22453 -6826 -22419
rect -6790 -22453 -6758 -22419
rect -6718 -22453 -6690 -22419
rect -6646 -22453 -6622 -22419
rect -6588 -22453 -6549 -22419
rect -6119 -22453 -6080 -22419
rect -6046 -22453 -6022 -22419
rect -5978 -22453 -5950 -22419
rect -5910 -22453 -5878 -22419
rect -5842 -22453 -5808 -22419
rect -5772 -22453 -5740 -22419
rect -5700 -22453 -5672 -22419
rect -5628 -22453 -5604 -22419
rect -5570 -22453 -5531 -22419
rect -5101 -22453 -5062 -22419
rect -5028 -22453 -5004 -22419
rect -4960 -22453 -4932 -22419
rect -4892 -22453 -4860 -22419
rect -4824 -22453 -4790 -22419
rect -4754 -22453 -4722 -22419
rect -4682 -22453 -4654 -22419
rect -4610 -22453 -4586 -22419
rect -4552 -22453 -4513 -22419
rect -4083 -22453 -4044 -22419
rect -4010 -22453 -3986 -22419
rect -3942 -22453 -3914 -22419
rect -3874 -22453 -3842 -22419
rect -3806 -22453 -3772 -22419
rect -3736 -22453 -3704 -22419
rect -3664 -22453 -3636 -22419
rect -3592 -22453 -3568 -22419
rect -3534 -22453 -3495 -22419
rect -2322 -22452 -2295 -22418
rect -2193 -22452 -2166 -22418
rect -2024 -22452 -1997 -22418
rect -1895 -22452 -1868 -22418
rect -1726 -22452 -1699 -22418
rect -1597 -22452 -1570 -22418
rect -1428 -22452 -1401 -22418
rect -1299 -22452 -1272 -22418
rect -1130 -22452 -1103 -22418
rect -1001 -22452 -974 -22418
rect -832 -22452 -805 -22418
rect -703 -22452 -676 -22418
rect -534 -22452 -507 -22418
rect -405 -22452 -378 -22418
rect -236 -22452 -209 -22418
rect -107 -22452 -80 -22418
rect 62 -22452 89 -22418
rect 191 -22452 218 -22418
rect 360 -22452 387 -22418
rect 489 -22452 516 -22418
rect 658 -22452 685 -22418
rect 787 -22452 814 -22418
rect 24822 -22421 24855 -22379
rect 24889 -22421 24922 -22379
rect 24822 -22447 24922 -22421
rect -1974 -22472 -1914 -22452
rect -12322 -22515 -12222 -22493
rect -12322 -22565 -12289 -22515
rect -12255 -22565 -12222 -22515
rect -12322 -22583 -12222 -22565
rect -12322 -22637 -12289 -22583
rect -12255 -22637 -12222 -22583
rect -12322 -22651 -12222 -22637
rect -12322 -22709 -12289 -22651
rect -12255 -22709 -12222 -22651
rect -12322 -22719 -12222 -22709
rect -12322 -22781 -12289 -22719
rect -12255 -22781 -12222 -22719
rect 24822 -22493 24855 -22447
rect 24889 -22493 24922 -22447
rect 24822 -22515 24922 -22493
rect 24822 -22565 24855 -22515
rect 24889 -22565 24922 -22515
rect 24822 -22583 24922 -22565
rect 24822 -22637 24855 -22583
rect 24889 -22637 24922 -22583
rect 24822 -22651 24922 -22637
rect 24822 -22709 24855 -22651
rect 24889 -22709 24922 -22651
rect 24822 -22719 24922 -22709
rect 2812 -22780 2851 -22746
rect 2885 -22780 2909 -22746
rect 2953 -22780 2981 -22746
rect 3021 -22780 3053 -22746
rect 3089 -22780 3123 -22746
rect 3159 -22780 3191 -22746
rect 3231 -22780 3259 -22746
rect 3303 -22780 3327 -22746
rect 3361 -22780 3400 -22746
rect 3830 -22780 3869 -22746
rect 3903 -22780 3927 -22746
rect 3971 -22780 3999 -22746
rect 4039 -22780 4071 -22746
rect 4107 -22780 4141 -22746
rect 4177 -22780 4209 -22746
rect 4249 -22780 4277 -22746
rect 4321 -22780 4345 -22746
rect 4379 -22780 4418 -22746
rect 4848 -22780 4887 -22746
rect 4921 -22780 4945 -22746
rect 4989 -22780 5017 -22746
rect 5057 -22780 5089 -22746
rect 5125 -22780 5159 -22746
rect 5195 -22780 5227 -22746
rect 5267 -22780 5295 -22746
rect 5339 -22780 5363 -22746
rect 5397 -22780 5436 -22746
rect 5866 -22780 5905 -22746
rect 5939 -22780 5963 -22746
rect 6007 -22780 6035 -22746
rect 6075 -22780 6107 -22746
rect 6143 -22780 6177 -22746
rect 6213 -22780 6245 -22746
rect 6285 -22780 6313 -22746
rect 6357 -22780 6381 -22746
rect 6415 -22780 6454 -22746
rect 6884 -22780 6923 -22746
rect 6957 -22780 6981 -22746
rect 7025 -22780 7053 -22746
rect 7093 -22780 7125 -22746
rect 7161 -22780 7195 -22746
rect 7231 -22780 7263 -22746
rect 7303 -22780 7331 -22746
rect 7375 -22780 7399 -22746
rect 7433 -22780 7472 -22746
rect 7902 -22780 7941 -22746
rect 7975 -22780 7999 -22746
rect 8043 -22780 8071 -22746
rect 8111 -22780 8143 -22746
rect 8179 -22780 8213 -22746
rect 8249 -22780 8281 -22746
rect 8321 -22780 8349 -22746
rect 8393 -22780 8417 -22746
rect 8451 -22780 8490 -22746
rect 8920 -22780 8959 -22746
rect 8993 -22780 9017 -22746
rect 9061 -22780 9089 -22746
rect 9129 -22780 9161 -22746
rect 9197 -22780 9231 -22746
rect 9267 -22780 9299 -22746
rect 9339 -22780 9367 -22746
rect 9411 -22780 9435 -22746
rect 9469 -22780 9508 -22746
rect 9938 -22780 9977 -22746
rect 10011 -22780 10035 -22746
rect 10079 -22780 10107 -22746
rect 10147 -22780 10179 -22746
rect 10215 -22780 10249 -22746
rect 10285 -22780 10317 -22746
rect 10357 -22780 10385 -22746
rect 10429 -22780 10453 -22746
rect 10487 -22780 10526 -22746
rect 10956 -22780 10995 -22746
rect 11029 -22780 11053 -22746
rect 11097 -22780 11125 -22746
rect 11165 -22780 11197 -22746
rect 11233 -22780 11267 -22746
rect 11303 -22780 11335 -22746
rect 11375 -22780 11403 -22746
rect 11447 -22780 11471 -22746
rect 11505 -22780 11544 -22746
rect 11974 -22780 12013 -22746
rect 12047 -22780 12071 -22746
rect 12115 -22780 12143 -22746
rect 12183 -22780 12215 -22746
rect 12251 -22780 12285 -22746
rect 12321 -22780 12353 -22746
rect 12393 -22780 12421 -22746
rect 12465 -22780 12489 -22746
rect 12523 -22780 12562 -22746
rect 12992 -22780 13031 -22746
rect 13065 -22780 13089 -22746
rect 13133 -22780 13161 -22746
rect 13201 -22780 13233 -22746
rect 13269 -22780 13303 -22746
rect 13339 -22780 13371 -22746
rect 13411 -22780 13439 -22746
rect 13483 -22780 13507 -22746
rect 13541 -22780 13580 -22746
rect 14010 -22780 14049 -22746
rect 14083 -22780 14107 -22746
rect 14151 -22780 14179 -22746
rect 14219 -22780 14251 -22746
rect 14287 -22780 14321 -22746
rect 14357 -22780 14389 -22746
rect 14429 -22780 14457 -22746
rect 14501 -22780 14525 -22746
rect 14559 -22780 14598 -22746
rect 15028 -22780 15067 -22746
rect 15101 -22780 15125 -22746
rect 15169 -22780 15197 -22746
rect 15237 -22780 15269 -22746
rect 15305 -22780 15339 -22746
rect 15375 -22780 15407 -22746
rect 15447 -22780 15475 -22746
rect 15519 -22780 15543 -22746
rect 15577 -22780 15616 -22746
rect 16046 -22780 16085 -22746
rect 16119 -22780 16143 -22746
rect 16187 -22780 16215 -22746
rect 16255 -22780 16287 -22746
rect 16323 -22780 16357 -22746
rect 16393 -22780 16425 -22746
rect 16465 -22780 16493 -22746
rect 16537 -22780 16561 -22746
rect 16595 -22780 16634 -22746
rect 17064 -22780 17103 -22746
rect 17137 -22780 17161 -22746
rect 17205 -22780 17233 -22746
rect 17273 -22780 17305 -22746
rect 17341 -22780 17375 -22746
rect 17411 -22780 17443 -22746
rect 17483 -22780 17511 -22746
rect 17555 -22780 17579 -22746
rect 17613 -22780 17652 -22746
rect 18082 -22780 18121 -22746
rect 18155 -22780 18179 -22746
rect 18223 -22780 18251 -22746
rect 18291 -22780 18323 -22746
rect 18359 -22780 18393 -22746
rect 18429 -22780 18461 -22746
rect 18501 -22780 18529 -22746
rect 18573 -22780 18597 -22746
rect 18631 -22780 18670 -22746
rect 19100 -22780 19139 -22746
rect 19173 -22780 19197 -22746
rect 19241 -22780 19269 -22746
rect 19309 -22780 19341 -22746
rect 19377 -22780 19411 -22746
rect 19447 -22780 19479 -22746
rect 19519 -22780 19547 -22746
rect 19591 -22780 19615 -22746
rect 19649 -22780 19688 -22746
rect 20118 -22780 20157 -22746
rect 20191 -22780 20215 -22746
rect 20259 -22780 20287 -22746
rect 20327 -22780 20359 -22746
rect 20395 -22780 20429 -22746
rect 20465 -22780 20497 -22746
rect 20537 -22780 20565 -22746
rect 20609 -22780 20633 -22746
rect 20667 -22780 20706 -22746
rect 21136 -22780 21175 -22746
rect 21209 -22780 21233 -22746
rect 21277 -22780 21305 -22746
rect 21345 -22780 21377 -22746
rect 21413 -22780 21447 -22746
rect 21483 -22780 21515 -22746
rect 21555 -22780 21583 -22746
rect 21627 -22780 21651 -22746
rect 21685 -22780 21724 -22746
rect 22154 -22780 22193 -22746
rect 22227 -22780 22251 -22746
rect 22295 -22780 22323 -22746
rect 22363 -22780 22395 -22746
rect 22431 -22780 22465 -22746
rect 22501 -22780 22533 -22746
rect 22573 -22780 22601 -22746
rect 22645 -22780 22669 -22746
rect 22703 -22780 22742 -22746
rect -12322 -22787 -12222 -22781
rect 6120 -22782 6180 -22780
rect 24822 -22781 24855 -22719
rect 24889 -22781 24922 -22719
rect -12322 -22853 -12289 -22787
rect -12255 -22853 -12222 -22787
rect 24822 -22787 24922 -22781
rect -12322 -22855 -12222 -22853
rect -12322 -22889 -12289 -22855
rect -12255 -22889 -12222 -22855
rect -9174 -22856 -9135 -22822
rect -9101 -22856 -9077 -22822
rect -9033 -22856 -9005 -22822
rect -8965 -22856 -8933 -22822
rect -8897 -22856 -8863 -22822
rect -8827 -22856 -8795 -22822
rect -8755 -22856 -8727 -22822
rect -8683 -22856 -8659 -22822
rect -8625 -22856 -8586 -22822
rect -8156 -22856 -8117 -22822
rect -8083 -22856 -8059 -22822
rect -8015 -22856 -7987 -22822
rect -7947 -22856 -7915 -22822
rect -7879 -22856 -7845 -22822
rect -7809 -22856 -7777 -22822
rect -7737 -22856 -7709 -22822
rect -7665 -22856 -7641 -22822
rect -7607 -22856 -7568 -22822
rect -7138 -22856 -7099 -22822
rect -7065 -22856 -7041 -22822
rect -6997 -22856 -6969 -22822
rect -6929 -22856 -6897 -22822
rect -6861 -22856 -6827 -22822
rect -6791 -22856 -6759 -22822
rect -6719 -22856 -6691 -22822
rect -6647 -22856 -6623 -22822
rect -6589 -22856 -6550 -22822
rect -6120 -22856 -6081 -22822
rect -6047 -22856 -6023 -22822
rect -5979 -22856 -5951 -22822
rect -5911 -22856 -5879 -22822
rect -5843 -22856 -5809 -22822
rect -5773 -22856 -5741 -22822
rect -5701 -22856 -5673 -22822
rect -5629 -22856 -5605 -22822
rect -5571 -22856 -5532 -22822
rect -5102 -22856 -5063 -22822
rect -5029 -22856 -5005 -22822
rect -4961 -22856 -4933 -22822
rect -4893 -22856 -4861 -22822
rect -4825 -22856 -4791 -22822
rect -4755 -22856 -4723 -22822
rect -4683 -22856 -4655 -22822
rect -4611 -22856 -4587 -22822
rect -4553 -22856 -4514 -22822
rect -4084 -22856 -4045 -22822
rect -4011 -22856 -3987 -22822
rect -3943 -22856 -3915 -22822
rect -3875 -22856 -3843 -22822
rect -3807 -22856 -3773 -22822
rect -3737 -22856 -3705 -22822
rect -3665 -22856 -3637 -22822
rect -3593 -22856 -3569 -22822
rect -3535 -22856 -3496 -22822
rect -2322 -22854 -2295 -22820
rect -2193 -22854 -2166 -22820
rect -2024 -22854 -1997 -22820
rect -1895 -22854 -1868 -22820
rect -1726 -22854 -1699 -22820
rect -1597 -22854 -1570 -22820
rect -1428 -22854 -1401 -22820
rect -1299 -22854 -1272 -22820
rect -1130 -22854 -1103 -22820
rect -1001 -22854 -974 -22820
rect -832 -22854 -805 -22820
rect -703 -22854 -676 -22820
rect -534 -22854 -507 -22820
rect -405 -22854 -378 -22820
rect -236 -22854 -209 -22820
rect -107 -22854 -80 -22820
rect 62 -22854 89 -22820
rect 191 -22854 218 -22820
rect 360 -22854 387 -22820
rect 489 -22854 516 -22820
rect 658 -22854 685 -22820
rect 787 -22854 814 -22820
rect 2580 -22849 2614 -22814
rect -7892 -22858 -7832 -22856
rect -5856 -22858 -5796 -22856
rect -4834 -22858 -4774 -22856
rect -12322 -22891 -12222 -22889
rect -12322 -22957 -12289 -22891
rect -12255 -22957 -12222 -22891
rect -12322 -22963 -12222 -22957
rect -12322 -23025 -12289 -22963
rect -12255 -23025 -12222 -22963
rect -12322 -23035 -12222 -23025
rect -12322 -23093 -12289 -23035
rect -12255 -23093 -12222 -23035
rect -12322 -23107 -12222 -23093
rect -12322 -23161 -12289 -23107
rect -12255 -23161 -12222 -23107
rect -12322 -23179 -12222 -23161
rect -12322 -23229 -12289 -23179
rect -12255 -23229 -12222 -23179
rect -12322 -23251 -12222 -23229
rect -12322 -23297 -12289 -23251
rect -12255 -23297 -12222 -23251
rect -12322 -23323 -12222 -23297
rect -12322 -23365 -12289 -23323
rect -12255 -23365 -12222 -23323
rect -12322 -23395 -12222 -23365
rect -12322 -23433 -12289 -23395
rect -12255 -23433 -12222 -23395
rect -12322 -23467 -12222 -23433
rect -12322 -23501 -12289 -23467
rect -12255 -23501 -12222 -23467
rect -9406 -22925 -9372 -22890
rect -9406 -22997 -9372 -22973
rect -9406 -23069 -9372 -23041
rect -9406 -23141 -9372 -23109
rect -9406 -23211 -9372 -23177
rect -9406 -23279 -9372 -23247
rect -9406 -23347 -9372 -23319
rect -9406 -23415 -9372 -23391
rect -9406 -23498 -9372 -23463
rect -8388 -22925 -8354 -22890
rect -8388 -22997 -8354 -22973
rect -8388 -23069 -8354 -23041
rect -8388 -23141 -8354 -23109
rect -8388 -23211 -8354 -23177
rect -8388 -23279 -8354 -23247
rect -8388 -23347 -8354 -23319
rect -8388 -23415 -8354 -23391
rect -8388 -23498 -8354 -23463
rect -7370 -22925 -7336 -22890
rect -7370 -22997 -7336 -22973
rect -7370 -23069 -7336 -23041
rect -7370 -23141 -7336 -23109
rect -7370 -23211 -7336 -23177
rect -7370 -23279 -7336 -23247
rect -7370 -23347 -7336 -23319
rect -7370 -23415 -7336 -23391
rect -7370 -23498 -7336 -23463
rect -6352 -22925 -6318 -22890
rect -6352 -22997 -6318 -22973
rect -6352 -23069 -6318 -23041
rect -6352 -23141 -6318 -23109
rect -6352 -23211 -6318 -23177
rect -6352 -23279 -6318 -23247
rect -6352 -23347 -6318 -23319
rect -6352 -23415 -6318 -23391
rect -6352 -23498 -6318 -23463
rect -5334 -22925 -5300 -22890
rect -5334 -22997 -5300 -22973
rect -5334 -23069 -5300 -23041
rect -5334 -23141 -5300 -23109
rect -5334 -23211 -5300 -23177
rect -5334 -23279 -5300 -23247
rect -5334 -23347 -5300 -23319
rect -5334 -23415 -5300 -23391
rect -5334 -23498 -5300 -23463
rect -4316 -22925 -4282 -22890
rect -4316 -22997 -4282 -22973
rect -4316 -23069 -4282 -23041
rect -4316 -23141 -4282 -23109
rect -4316 -23211 -4282 -23177
rect -4316 -23279 -4282 -23247
rect -4316 -23347 -4282 -23319
rect -4316 -23415 -4282 -23391
rect -4316 -23498 -4282 -23463
rect -3298 -22925 -3264 -22890
rect -3298 -22997 -3264 -22973
rect -3298 -23069 -3264 -23041
rect -3298 -23141 -3264 -23109
rect -3298 -23211 -3264 -23177
rect -3298 -23279 -3264 -23247
rect -3298 -23347 -3264 -23319
rect -3298 -23415 -3264 -23391
rect -3298 -23498 -3264 -23463
rect -2410 -22923 -2376 -22888
rect -2410 -22995 -2376 -22971
rect -2410 -23067 -2376 -23039
rect -2410 -23139 -2376 -23107
rect -2410 -23209 -2376 -23175
rect -2410 -23277 -2376 -23245
rect -2410 -23345 -2376 -23317
rect -2410 -23413 -2376 -23389
rect -2410 -23496 -2376 -23461
rect -2112 -22923 -2078 -22888
rect -2112 -22995 -2078 -22971
rect -2112 -23067 -2078 -23039
rect -2112 -23139 -2078 -23107
rect -2112 -23209 -2078 -23175
rect -2112 -23277 -2078 -23245
rect -2112 -23345 -2078 -23317
rect -2112 -23413 -2078 -23389
rect -2112 -23496 -2078 -23461
rect -1814 -22923 -1780 -22888
rect -1814 -22995 -1780 -22971
rect -1814 -23067 -1780 -23039
rect -1814 -23139 -1780 -23107
rect -1814 -23209 -1780 -23175
rect -1814 -23277 -1780 -23245
rect -1814 -23345 -1780 -23317
rect -1814 -23413 -1780 -23389
rect -1814 -23496 -1780 -23461
rect -1516 -22923 -1482 -22888
rect -1516 -22995 -1482 -22971
rect -1516 -23067 -1482 -23039
rect -1516 -23139 -1482 -23107
rect -1516 -23209 -1482 -23175
rect -1516 -23277 -1482 -23245
rect -1516 -23345 -1482 -23317
rect -1516 -23413 -1482 -23389
rect -1516 -23496 -1482 -23461
rect -1218 -22923 -1184 -22888
rect -1218 -22995 -1184 -22971
rect -1218 -23067 -1184 -23039
rect -1218 -23139 -1184 -23107
rect -1218 -23209 -1184 -23175
rect -1218 -23277 -1184 -23245
rect -1218 -23345 -1184 -23317
rect -1218 -23413 -1184 -23389
rect -1218 -23496 -1184 -23461
rect -920 -22923 -886 -22888
rect -920 -22995 -886 -22971
rect -920 -23067 -886 -23039
rect -920 -23139 -886 -23107
rect -920 -23209 -886 -23175
rect -920 -23277 -886 -23245
rect -920 -23345 -886 -23317
rect -920 -23413 -886 -23389
rect -920 -23496 -886 -23461
rect -622 -22923 -588 -22888
rect -622 -22995 -588 -22971
rect -622 -23067 -588 -23039
rect -622 -23139 -588 -23107
rect -622 -23209 -588 -23175
rect -622 -23277 -588 -23245
rect -622 -23345 -588 -23317
rect -622 -23413 -588 -23389
rect -622 -23496 -588 -23461
rect -324 -22923 -290 -22888
rect -324 -22995 -290 -22971
rect -324 -23067 -290 -23039
rect -324 -23139 -290 -23107
rect -324 -23209 -290 -23175
rect -324 -23277 -290 -23245
rect -324 -23345 -290 -23317
rect -324 -23413 -290 -23389
rect -324 -23496 -290 -23461
rect -26 -22923 8 -22888
rect -26 -22995 8 -22971
rect -26 -23067 8 -23039
rect -26 -23139 8 -23107
rect -26 -23209 8 -23175
rect -26 -23277 8 -23245
rect -26 -23345 8 -23317
rect -26 -23413 8 -23389
rect -26 -23496 8 -23461
rect 272 -22923 306 -22888
rect 272 -22995 306 -22971
rect 272 -23067 306 -23039
rect 272 -23139 306 -23107
rect 272 -23209 306 -23175
rect 272 -23277 306 -23245
rect 272 -23345 306 -23317
rect 272 -23413 306 -23389
rect 272 -23496 306 -23461
rect 570 -22923 604 -22888
rect 570 -22995 604 -22971
rect 570 -23067 604 -23039
rect 570 -23139 604 -23107
rect 570 -23209 604 -23175
rect 570 -23277 604 -23245
rect 570 -23345 604 -23317
rect 570 -23413 604 -23389
rect 570 -23496 604 -23461
rect 868 -22923 902 -22888
rect 868 -22995 902 -22971
rect 868 -23067 902 -23039
rect 868 -23139 902 -23107
rect 868 -23209 902 -23175
rect 868 -23277 902 -23245
rect 868 -23345 902 -23317
rect 868 -23413 902 -23389
rect 2580 -22921 2614 -22897
rect 2580 -22993 2614 -22965
rect 2580 -23065 2614 -23033
rect 2580 -23135 2614 -23101
rect 2580 -23203 2614 -23171
rect 2580 -23271 2614 -23243
rect 2580 -23339 2614 -23315
rect 2580 -23422 2614 -23387
rect 3598 -22849 3632 -22814
rect 3598 -22921 3632 -22897
rect 3598 -22993 3632 -22965
rect 3598 -23065 3632 -23033
rect 3598 -23135 3632 -23101
rect 3598 -23203 3632 -23171
rect 3598 -23271 3632 -23243
rect 3598 -23339 3632 -23315
rect 3598 -23422 3632 -23387
rect 4616 -22849 4650 -22814
rect 4616 -22921 4650 -22897
rect 4616 -22993 4650 -22965
rect 4616 -23065 4650 -23033
rect 4616 -23135 4650 -23101
rect 4616 -23203 4650 -23171
rect 4616 -23271 4650 -23243
rect 4616 -23339 4650 -23315
rect 4616 -23422 4650 -23387
rect 5634 -22849 5668 -22814
rect 5634 -22921 5668 -22897
rect 5634 -22993 5668 -22965
rect 5634 -23065 5668 -23033
rect 5634 -23135 5668 -23101
rect 5634 -23203 5668 -23171
rect 5634 -23271 5668 -23243
rect 5634 -23339 5668 -23315
rect 5634 -23422 5668 -23387
rect 6652 -22849 6686 -22814
rect 6652 -22921 6686 -22897
rect 6652 -22993 6686 -22965
rect 6652 -23065 6686 -23033
rect 6652 -23135 6686 -23101
rect 6652 -23203 6686 -23171
rect 6652 -23271 6686 -23243
rect 6652 -23339 6686 -23315
rect 6652 -23422 6686 -23387
rect 7670 -22849 7704 -22814
rect 7670 -22921 7704 -22897
rect 7670 -22993 7704 -22965
rect 7670 -23065 7704 -23033
rect 7670 -23135 7704 -23101
rect 7670 -23203 7704 -23171
rect 7670 -23271 7704 -23243
rect 7670 -23339 7704 -23315
rect 7670 -23422 7704 -23387
rect 8688 -22849 8722 -22814
rect 8688 -22921 8722 -22897
rect 8688 -22993 8722 -22965
rect 8688 -23065 8722 -23033
rect 8688 -23135 8722 -23101
rect 8688 -23203 8722 -23171
rect 8688 -23271 8722 -23243
rect 8688 -23339 8722 -23315
rect 8688 -23422 8722 -23387
rect 9706 -22849 9740 -22814
rect 9706 -22921 9740 -22897
rect 9706 -22993 9740 -22965
rect 9706 -23065 9740 -23033
rect 9706 -23135 9740 -23101
rect 9706 -23203 9740 -23171
rect 9706 -23271 9740 -23243
rect 9706 -23339 9740 -23315
rect 9706 -23422 9740 -23387
rect 10724 -22849 10758 -22814
rect 10724 -22921 10758 -22897
rect 10724 -22993 10758 -22965
rect 10724 -23065 10758 -23033
rect 10724 -23135 10758 -23101
rect 10724 -23203 10758 -23171
rect 10724 -23271 10758 -23243
rect 10724 -23339 10758 -23315
rect 10724 -23422 10758 -23387
rect 11742 -22849 11776 -22814
rect 11742 -22921 11776 -22897
rect 11742 -22993 11776 -22965
rect 11742 -23065 11776 -23033
rect 11742 -23135 11776 -23101
rect 11742 -23203 11776 -23171
rect 11742 -23271 11776 -23243
rect 11742 -23339 11776 -23315
rect 11742 -23422 11776 -23387
rect 12760 -22849 12794 -22814
rect 12760 -22921 12794 -22897
rect 12760 -22993 12794 -22965
rect 12760 -23065 12794 -23033
rect 12760 -23135 12794 -23101
rect 12760 -23203 12794 -23171
rect 12760 -23271 12794 -23243
rect 12760 -23339 12794 -23315
rect 12760 -23422 12794 -23387
rect 13778 -22849 13812 -22814
rect 13778 -22921 13812 -22897
rect 13778 -22993 13812 -22965
rect 13778 -23065 13812 -23033
rect 13778 -23135 13812 -23101
rect 13778 -23203 13812 -23171
rect 13778 -23271 13812 -23243
rect 13778 -23339 13812 -23315
rect 13778 -23422 13812 -23387
rect 14796 -22849 14830 -22814
rect 14796 -22921 14830 -22897
rect 14796 -22993 14830 -22965
rect 14796 -23065 14830 -23033
rect 14796 -23135 14830 -23101
rect 14796 -23203 14830 -23171
rect 14796 -23271 14830 -23243
rect 14796 -23339 14830 -23315
rect 14796 -23422 14830 -23387
rect 15814 -22849 15848 -22814
rect 15814 -22921 15848 -22897
rect 15814 -22993 15848 -22965
rect 15814 -23065 15848 -23033
rect 15814 -23135 15848 -23101
rect 15814 -23203 15848 -23171
rect 15814 -23271 15848 -23243
rect 15814 -23339 15848 -23315
rect 15814 -23422 15848 -23387
rect 16832 -22849 16866 -22814
rect 16832 -22921 16866 -22897
rect 16832 -22993 16866 -22965
rect 16832 -23065 16866 -23033
rect 16832 -23135 16866 -23101
rect 16832 -23203 16866 -23171
rect 16832 -23271 16866 -23243
rect 16832 -23339 16866 -23315
rect 16832 -23422 16866 -23387
rect 17850 -22849 17884 -22814
rect 17850 -22921 17884 -22897
rect 17850 -22993 17884 -22965
rect 17850 -23065 17884 -23033
rect 17850 -23135 17884 -23101
rect 17850 -23203 17884 -23171
rect 17850 -23271 17884 -23243
rect 17850 -23339 17884 -23315
rect 17850 -23422 17884 -23387
rect 18868 -22849 18902 -22814
rect 18868 -22921 18902 -22897
rect 18868 -22993 18902 -22965
rect 18868 -23065 18902 -23033
rect 18868 -23135 18902 -23101
rect 18868 -23203 18902 -23171
rect 18868 -23271 18902 -23243
rect 18868 -23339 18902 -23315
rect 18868 -23422 18902 -23387
rect 19886 -22849 19920 -22814
rect 19886 -22921 19920 -22897
rect 19886 -22993 19920 -22965
rect 19886 -23065 19920 -23033
rect 19886 -23135 19920 -23101
rect 19886 -23203 19920 -23171
rect 19886 -23271 19920 -23243
rect 19886 -23339 19920 -23315
rect 19886 -23422 19920 -23387
rect 20904 -22849 20938 -22814
rect 20904 -22921 20938 -22897
rect 20904 -22993 20938 -22965
rect 20904 -23065 20938 -23033
rect 20904 -23135 20938 -23101
rect 20904 -23203 20938 -23171
rect 20904 -23271 20938 -23243
rect 20904 -23339 20938 -23315
rect 20904 -23422 20938 -23387
rect 21922 -22849 21956 -22814
rect 21922 -22921 21956 -22897
rect 21922 -22993 21956 -22965
rect 21922 -23065 21956 -23033
rect 21922 -23135 21956 -23101
rect 21922 -23203 21956 -23171
rect 21922 -23271 21956 -23243
rect 21922 -23339 21956 -23315
rect 21922 -23422 21956 -23387
rect 22940 -22849 22974 -22814
rect 22940 -22921 22974 -22897
rect 22940 -22993 22974 -22965
rect 22940 -23065 22974 -23033
rect 22940 -23135 22974 -23101
rect 22940 -23203 22974 -23171
rect 22940 -23271 22974 -23243
rect 22940 -23339 22974 -23315
rect 22940 -23422 22974 -23387
rect 24822 -22853 24855 -22787
rect 24889 -22853 24922 -22787
rect 24822 -22855 24922 -22853
rect 24822 -22889 24855 -22855
rect 24889 -22889 24922 -22855
rect 24822 -22891 24922 -22889
rect 24822 -22957 24855 -22891
rect 24889 -22957 24922 -22891
rect 24822 -22963 24922 -22957
rect 24822 -23025 24855 -22963
rect 24889 -23025 24922 -22963
rect 24822 -23035 24922 -23025
rect 24822 -23093 24855 -23035
rect 24889 -23093 24922 -23035
rect 24822 -23107 24922 -23093
rect 24822 -23161 24855 -23107
rect 24889 -23161 24922 -23107
rect 24822 -23179 24922 -23161
rect 24822 -23229 24855 -23179
rect 24889 -23229 24922 -23179
rect 24822 -23251 24922 -23229
rect 24822 -23297 24855 -23251
rect 24889 -23297 24922 -23251
rect 24822 -23323 24922 -23297
rect 24822 -23365 24855 -23323
rect 24889 -23365 24922 -23323
rect 24822 -23395 24922 -23365
rect 24822 -23433 24855 -23395
rect 24889 -23433 24922 -23395
rect 4088 -23456 4148 -23454
rect 10200 -23456 10260 -23454
rect 12234 -23456 12294 -23454
rect 16300 -23456 16360 -23450
rect 20376 -23456 20436 -23454
rect 21392 -23456 21452 -23454
rect 868 -23496 902 -23461
rect 2812 -23490 2851 -23456
rect 2885 -23490 2909 -23456
rect 2953 -23490 2981 -23456
rect 3021 -23490 3053 -23456
rect 3089 -23490 3123 -23456
rect 3159 -23490 3191 -23456
rect 3231 -23490 3259 -23456
rect 3303 -23490 3327 -23456
rect 3361 -23490 3400 -23456
rect 3830 -23490 3869 -23456
rect 3903 -23490 3927 -23456
rect 3971 -23490 3999 -23456
rect 4039 -23490 4071 -23456
rect 4107 -23490 4141 -23456
rect 4177 -23490 4209 -23456
rect 4249 -23490 4277 -23456
rect 4321 -23490 4345 -23456
rect 4379 -23490 4418 -23456
rect 4848 -23490 4887 -23456
rect 4921 -23490 4945 -23456
rect 4989 -23490 5017 -23456
rect 5057 -23490 5089 -23456
rect 5125 -23490 5159 -23456
rect 5195 -23490 5227 -23456
rect 5267 -23490 5295 -23456
rect 5339 -23490 5363 -23456
rect 5397 -23490 5436 -23456
rect 5866 -23490 5905 -23456
rect 5939 -23490 5963 -23456
rect 6007 -23490 6035 -23456
rect 6075 -23490 6107 -23456
rect 6143 -23490 6177 -23456
rect 6213 -23490 6245 -23456
rect 6285 -23490 6313 -23456
rect 6357 -23490 6381 -23456
rect 6415 -23490 6454 -23456
rect 6884 -23490 6923 -23456
rect 6957 -23490 6981 -23456
rect 7025 -23490 7053 -23456
rect 7093 -23490 7125 -23456
rect 7161 -23490 7195 -23456
rect 7231 -23490 7263 -23456
rect 7303 -23490 7331 -23456
rect 7375 -23490 7399 -23456
rect 7433 -23490 7472 -23456
rect 7902 -23490 7941 -23456
rect 7975 -23490 7999 -23456
rect 8043 -23490 8071 -23456
rect 8111 -23490 8143 -23456
rect 8179 -23490 8213 -23456
rect 8249 -23490 8281 -23456
rect 8321 -23490 8349 -23456
rect 8393 -23490 8417 -23456
rect 8451 -23490 8490 -23456
rect 8920 -23490 8959 -23456
rect 8993 -23490 9017 -23456
rect 9061 -23490 9089 -23456
rect 9129 -23490 9161 -23456
rect 9197 -23490 9231 -23456
rect 9267 -23490 9299 -23456
rect 9339 -23490 9367 -23456
rect 9411 -23490 9435 -23456
rect 9469 -23490 9508 -23456
rect 9938 -23490 9977 -23456
rect 10011 -23490 10035 -23456
rect 10079 -23490 10107 -23456
rect 10147 -23490 10179 -23456
rect 10215 -23490 10249 -23456
rect 10285 -23490 10317 -23456
rect 10357 -23490 10385 -23456
rect 10429 -23490 10453 -23456
rect 10487 -23490 10526 -23456
rect 10956 -23490 10995 -23456
rect 11029 -23490 11053 -23456
rect 11097 -23490 11125 -23456
rect 11165 -23490 11197 -23456
rect 11233 -23490 11267 -23456
rect 11303 -23490 11335 -23456
rect 11375 -23490 11403 -23456
rect 11447 -23490 11471 -23456
rect 11505 -23490 11544 -23456
rect 11974 -23490 12013 -23456
rect 12047 -23490 12071 -23456
rect 12115 -23490 12143 -23456
rect 12183 -23490 12215 -23456
rect 12251 -23490 12285 -23456
rect 12321 -23490 12353 -23456
rect 12393 -23490 12421 -23456
rect 12465 -23490 12489 -23456
rect 12523 -23490 12562 -23456
rect 12992 -23490 13031 -23456
rect 13065 -23490 13089 -23456
rect 13133 -23490 13161 -23456
rect 13201 -23490 13233 -23456
rect 13269 -23490 13303 -23456
rect 13339 -23490 13371 -23456
rect 13411 -23490 13439 -23456
rect 13483 -23490 13507 -23456
rect 13541 -23490 13580 -23456
rect 14010 -23490 14049 -23456
rect 14083 -23490 14107 -23456
rect 14151 -23490 14179 -23456
rect 14219 -23490 14251 -23456
rect 14287 -23490 14321 -23456
rect 14357 -23490 14389 -23456
rect 14429 -23490 14457 -23456
rect 14501 -23490 14525 -23456
rect 14559 -23490 14598 -23456
rect 15028 -23490 15067 -23456
rect 15101 -23490 15125 -23456
rect 15169 -23490 15197 -23456
rect 15237 -23490 15269 -23456
rect 15305 -23490 15339 -23456
rect 15375 -23490 15407 -23456
rect 15447 -23490 15475 -23456
rect 15519 -23490 15543 -23456
rect 15577 -23490 15616 -23456
rect 16046 -23490 16085 -23456
rect 16119 -23490 16143 -23456
rect 16187 -23490 16215 -23456
rect 16255 -23490 16287 -23456
rect 16323 -23490 16357 -23456
rect 16393 -23490 16425 -23456
rect 16465 -23490 16493 -23456
rect 16537 -23490 16561 -23456
rect 16595 -23490 16634 -23456
rect 17064 -23490 17103 -23456
rect 17137 -23490 17161 -23456
rect 17205 -23490 17233 -23456
rect 17273 -23490 17305 -23456
rect 17341 -23490 17375 -23456
rect 17411 -23490 17443 -23456
rect 17483 -23490 17511 -23456
rect 17555 -23490 17579 -23456
rect 17613 -23490 17652 -23456
rect 18082 -23490 18121 -23456
rect 18155 -23490 18179 -23456
rect 18223 -23490 18251 -23456
rect 18291 -23490 18323 -23456
rect 18359 -23490 18393 -23456
rect 18429 -23490 18461 -23456
rect 18501 -23490 18529 -23456
rect 18573 -23490 18597 -23456
rect 18631 -23490 18670 -23456
rect 19100 -23490 19139 -23456
rect 19173 -23490 19197 -23456
rect 19241 -23490 19269 -23456
rect 19309 -23490 19341 -23456
rect 19377 -23490 19411 -23456
rect 19447 -23490 19479 -23456
rect 19519 -23490 19547 -23456
rect 19591 -23490 19615 -23456
rect 19649 -23490 19688 -23456
rect 20118 -23490 20157 -23456
rect 20191 -23490 20215 -23456
rect 20259 -23490 20287 -23456
rect 20327 -23490 20359 -23456
rect 20395 -23490 20429 -23456
rect 20465 -23490 20497 -23456
rect 20537 -23490 20565 -23456
rect 20609 -23490 20633 -23456
rect 20667 -23490 20706 -23456
rect 21136 -23490 21175 -23456
rect 21209 -23490 21233 -23456
rect 21277 -23490 21305 -23456
rect 21345 -23490 21377 -23456
rect 21413 -23490 21447 -23456
rect 21483 -23490 21515 -23456
rect 21555 -23490 21583 -23456
rect 21627 -23490 21651 -23456
rect 21685 -23490 21724 -23456
rect 22154 -23490 22193 -23456
rect 22227 -23490 22251 -23456
rect 22295 -23490 22323 -23456
rect 22363 -23490 22395 -23456
rect 22431 -23490 22465 -23456
rect 22501 -23490 22533 -23456
rect 22573 -23490 22601 -23456
rect 22645 -23490 22669 -23456
rect 22703 -23490 22742 -23456
rect 24822 -23467 24922 -23433
rect -12322 -23535 -12222 -23501
rect 24822 -23501 24855 -23467
rect 24889 -23501 24922 -23467
rect -7890 -23532 -7830 -23528
rect -6880 -23532 -6820 -23528
rect -4832 -23532 -4772 -23528
rect -12322 -23573 -12289 -23535
rect -12255 -23573 -12222 -23535
rect -9174 -23566 -9135 -23532
rect -9101 -23566 -9077 -23532
rect -9033 -23566 -9005 -23532
rect -8965 -23566 -8933 -23532
rect -8897 -23566 -8863 -23532
rect -8827 -23566 -8795 -23532
rect -8755 -23566 -8727 -23532
rect -8683 -23566 -8659 -23532
rect -8625 -23566 -8586 -23532
rect -8156 -23566 -8117 -23532
rect -8083 -23566 -8059 -23532
rect -8015 -23566 -7987 -23532
rect -7947 -23566 -7915 -23532
rect -7879 -23566 -7845 -23532
rect -7809 -23566 -7777 -23532
rect -7737 -23566 -7709 -23532
rect -7665 -23566 -7641 -23532
rect -7607 -23566 -7568 -23532
rect -7138 -23566 -7099 -23532
rect -7065 -23566 -7041 -23532
rect -6997 -23566 -6969 -23532
rect -6929 -23566 -6897 -23532
rect -6861 -23566 -6827 -23532
rect -6791 -23566 -6759 -23532
rect -6719 -23566 -6691 -23532
rect -6647 -23566 -6623 -23532
rect -6589 -23566 -6550 -23532
rect -6120 -23566 -6081 -23532
rect -6047 -23566 -6023 -23532
rect -5979 -23566 -5951 -23532
rect -5911 -23566 -5879 -23532
rect -5843 -23566 -5809 -23532
rect -5773 -23566 -5741 -23532
rect -5701 -23566 -5673 -23532
rect -5629 -23566 -5605 -23532
rect -5571 -23566 -5532 -23532
rect -5102 -23566 -5063 -23532
rect -5029 -23566 -5005 -23532
rect -4961 -23566 -4933 -23532
rect -4893 -23566 -4861 -23532
rect -4825 -23566 -4791 -23532
rect -4755 -23566 -4723 -23532
rect -4683 -23566 -4655 -23532
rect -4611 -23566 -4587 -23532
rect -4553 -23566 -4514 -23532
rect -4084 -23566 -4045 -23532
rect -4011 -23566 -3987 -23532
rect -3943 -23566 -3915 -23532
rect -3875 -23566 -3843 -23532
rect -3807 -23566 -3773 -23532
rect -3737 -23566 -3705 -23532
rect -3665 -23566 -3637 -23532
rect -3593 -23566 -3569 -23532
rect -3535 -23566 -3496 -23532
rect -2322 -23564 -2295 -23530
rect -2193 -23564 -2166 -23530
rect -2024 -23564 -1997 -23530
rect -1895 -23564 -1868 -23530
rect -1726 -23564 -1699 -23530
rect -1597 -23564 -1570 -23530
rect -1428 -23564 -1401 -23530
rect -1299 -23564 -1272 -23530
rect -1130 -23564 -1103 -23530
rect -1001 -23564 -974 -23530
rect -832 -23564 -805 -23530
rect -703 -23564 -676 -23530
rect -534 -23564 -507 -23530
rect -405 -23564 -378 -23530
rect -236 -23564 -209 -23530
rect -107 -23564 -80 -23530
rect 62 -23564 89 -23530
rect 191 -23564 218 -23530
rect 360 -23564 387 -23530
rect 489 -23564 516 -23530
rect 658 -23564 685 -23530
rect 787 -23564 814 -23530
rect 24822 -23535 24922 -23501
rect -12322 -23603 -12222 -23573
rect -12322 -23645 -12289 -23603
rect -12255 -23645 -12222 -23603
rect -12322 -23671 -12222 -23645
rect -12322 -23717 -12289 -23671
rect -12255 -23717 -12222 -23671
rect -12322 -23739 -12222 -23717
rect -12322 -23789 -12289 -23739
rect -12255 -23789 -12222 -23739
rect -12322 -23807 -12222 -23789
rect -12322 -23861 -12289 -23807
rect -12255 -23861 -12222 -23807
rect -12322 -23875 -12222 -23861
rect -12322 -23933 -12289 -23875
rect -12255 -23933 -12222 -23875
rect 24822 -23573 24855 -23535
rect 24889 -23573 24922 -23535
rect 24822 -23603 24922 -23573
rect 24822 -23645 24855 -23603
rect 24889 -23645 24922 -23603
rect 24822 -23671 24922 -23645
rect 24822 -23717 24855 -23671
rect 24889 -23717 24922 -23671
rect 24822 -23739 24922 -23717
rect 24822 -23789 24855 -23739
rect 24889 -23789 24922 -23739
rect 24822 -23807 24922 -23789
rect 24822 -23861 24855 -23807
rect 24889 -23861 24922 -23807
rect 24822 -23875 24922 -23861
rect -12322 -23943 -12222 -23933
rect -12322 -24005 -12289 -23943
rect -12255 -24005 -12222 -23943
rect -9173 -23967 -9134 -23933
rect -9100 -23967 -9076 -23933
rect -9032 -23967 -9004 -23933
rect -8964 -23967 -8932 -23933
rect -8896 -23967 -8862 -23933
rect -8826 -23967 -8794 -23933
rect -8754 -23967 -8726 -23933
rect -8682 -23967 -8658 -23933
rect -8624 -23967 -8585 -23933
rect -8155 -23967 -8116 -23933
rect -8082 -23967 -8058 -23933
rect -8014 -23967 -7986 -23933
rect -7946 -23967 -7914 -23933
rect -7878 -23967 -7844 -23933
rect -7808 -23967 -7776 -23933
rect -7736 -23967 -7708 -23933
rect -7664 -23967 -7640 -23933
rect -7606 -23967 -7567 -23933
rect -7137 -23967 -7098 -23933
rect -7064 -23967 -7040 -23933
rect -6996 -23967 -6968 -23933
rect -6928 -23967 -6896 -23933
rect -6860 -23967 -6826 -23933
rect -6790 -23967 -6758 -23933
rect -6718 -23967 -6690 -23933
rect -6646 -23967 -6622 -23933
rect -6588 -23967 -6549 -23933
rect -6119 -23967 -6080 -23933
rect -6046 -23967 -6022 -23933
rect -5978 -23967 -5950 -23933
rect -5910 -23967 -5878 -23933
rect -5842 -23967 -5808 -23933
rect -5772 -23967 -5740 -23933
rect -5700 -23967 -5672 -23933
rect -5628 -23967 -5604 -23933
rect -5570 -23967 -5531 -23933
rect -5101 -23967 -5062 -23933
rect -5028 -23967 -5004 -23933
rect -4960 -23967 -4932 -23933
rect -4892 -23967 -4860 -23933
rect -4824 -23967 -4790 -23933
rect -4754 -23967 -4722 -23933
rect -4682 -23967 -4654 -23933
rect -4610 -23967 -4586 -23933
rect -4552 -23967 -4513 -23933
rect -4083 -23967 -4044 -23933
rect -4010 -23967 -3986 -23933
rect -3942 -23967 -3914 -23933
rect -3874 -23967 -3842 -23933
rect -3806 -23967 -3772 -23933
rect -3736 -23967 -3704 -23933
rect -3664 -23967 -3636 -23933
rect -3592 -23967 -3568 -23933
rect -3534 -23967 -3495 -23933
rect -2324 -23966 -2297 -23932
rect -2195 -23966 -2168 -23932
rect -2026 -23966 -1999 -23932
rect -1897 -23966 -1870 -23932
rect -1728 -23966 -1701 -23932
rect -1599 -23966 -1572 -23932
rect -1430 -23966 -1403 -23932
rect -1301 -23966 -1274 -23932
rect -1132 -23966 -1105 -23932
rect -1003 -23966 -976 -23932
rect -834 -23966 -807 -23932
rect -705 -23966 -678 -23932
rect -536 -23966 -509 -23932
rect -407 -23966 -380 -23932
rect -238 -23966 -211 -23932
rect -109 -23966 -82 -23932
rect 60 -23966 87 -23932
rect 189 -23966 216 -23932
rect 358 -23966 385 -23932
rect 487 -23966 514 -23932
rect 656 -23966 683 -23932
rect 785 -23966 812 -23932
rect 24822 -23933 24855 -23875
rect 24889 -23933 24922 -23875
rect 24822 -23943 24922 -23933
rect -7890 -23968 -7830 -23967
rect -5854 -23968 -5794 -23967
rect -4832 -23968 -4772 -23967
rect -12322 -24011 -12222 -24005
rect -12322 -24077 -12289 -24011
rect -12255 -24077 -12222 -24011
rect -12322 -24079 -12222 -24077
rect -12322 -24113 -12289 -24079
rect -12255 -24113 -12222 -24079
rect -12322 -24115 -12222 -24113
rect -12322 -24181 -12289 -24115
rect -12255 -24181 -12222 -24115
rect -12322 -24187 -12222 -24181
rect -12322 -24249 -12289 -24187
rect -12255 -24249 -12222 -24187
rect -12322 -24259 -12222 -24249
rect -12322 -24317 -12289 -24259
rect -12255 -24317 -12222 -24259
rect -12322 -24331 -12222 -24317
rect -12322 -24385 -12289 -24331
rect -12255 -24385 -12222 -24331
rect -12322 -24403 -12222 -24385
rect -12322 -24453 -12289 -24403
rect -12255 -24453 -12222 -24403
rect -12322 -24475 -12222 -24453
rect -12322 -24521 -12289 -24475
rect -12255 -24521 -12222 -24475
rect -12322 -24547 -12222 -24521
rect -12322 -24589 -12289 -24547
rect -12255 -24589 -12222 -24547
rect -12322 -24619 -12222 -24589
rect -9405 -24036 -9371 -24001
rect -9405 -24108 -9371 -24084
rect -9405 -24180 -9371 -24152
rect -9405 -24252 -9371 -24220
rect -9405 -24322 -9371 -24288
rect -9405 -24390 -9371 -24358
rect -9405 -24458 -9371 -24430
rect -9405 -24526 -9371 -24502
rect -9405 -24609 -9371 -24574
rect -8387 -24036 -8353 -24001
rect -8387 -24108 -8353 -24084
rect -8387 -24180 -8353 -24152
rect -8387 -24252 -8353 -24220
rect -8387 -24322 -8353 -24288
rect -8387 -24390 -8353 -24358
rect -8387 -24458 -8353 -24430
rect -8387 -24526 -8353 -24502
rect -8387 -24609 -8353 -24574
rect -7369 -24036 -7335 -24001
rect -7369 -24108 -7335 -24084
rect -7369 -24180 -7335 -24152
rect -7369 -24252 -7335 -24220
rect -7369 -24322 -7335 -24288
rect -7369 -24390 -7335 -24358
rect -7369 -24458 -7335 -24430
rect -7369 -24526 -7335 -24502
rect -7369 -24609 -7335 -24574
rect -6351 -24036 -6317 -24001
rect -6351 -24108 -6317 -24084
rect -6351 -24180 -6317 -24152
rect -6351 -24252 -6317 -24220
rect -6351 -24322 -6317 -24288
rect -6351 -24390 -6317 -24358
rect -6351 -24458 -6317 -24430
rect -6351 -24526 -6317 -24502
rect -6351 -24609 -6317 -24574
rect -5333 -24036 -5299 -24001
rect -5333 -24108 -5299 -24084
rect -5333 -24180 -5299 -24152
rect -5333 -24252 -5299 -24220
rect -5333 -24322 -5299 -24288
rect -5333 -24390 -5299 -24358
rect -5333 -24458 -5299 -24430
rect -5333 -24526 -5299 -24502
rect -5333 -24609 -5299 -24574
rect -4315 -24036 -4281 -24001
rect -4315 -24108 -4281 -24084
rect -4315 -24180 -4281 -24152
rect -4315 -24252 -4281 -24220
rect -4315 -24322 -4281 -24288
rect -4315 -24390 -4281 -24358
rect -4315 -24458 -4281 -24430
rect -4315 -24526 -4281 -24502
rect -4315 -24609 -4281 -24574
rect -3297 -24036 -3263 -24001
rect -3297 -24108 -3263 -24084
rect -3297 -24180 -3263 -24152
rect -3297 -24252 -3263 -24220
rect -3297 -24322 -3263 -24288
rect -3297 -24390 -3263 -24358
rect -3297 -24458 -3263 -24430
rect -3297 -24526 -3263 -24502
rect -3297 -24609 -3263 -24574
rect -2412 -24035 -2378 -24000
rect -2412 -24107 -2378 -24083
rect -2412 -24179 -2378 -24151
rect -2412 -24251 -2378 -24219
rect -2412 -24321 -2378 -24287
rect -2412 -24389 -2378 -24357
rect -2412 -24457 -2378 -24429
rect -2412 -24525 -2378 -24501
rect -2412 -24608 -2378 -24573
rect -2114 -24035 -2080 -24000
rect -2114 -24107 -2080 -24083
rect -2114 -24179 -2080 -24151
rect -2114 -24251 -2080 -24219
rect -2114 -24321 -2080 -24287
rect -2114 -24389 -2080 -24357
rect -2114 -24457 -2080 -24429
rect -2114 -24525 -2080 -24501
rect -2114 -24608 -2080 -24573
rect -1816 -24035 -1782 -24000
rect -1816 -24107 -1782 -24083
rect -1816 -24179 -1782 -24151
rect -1816 -24251 -1782 -24219
rect -1816 -24321 -1782 -24287
rect -1816 -24389 -1782 -24357
rect -1816 -24457 -1782 -24429
rect -1816 -24525 -1782 -24501
rect -1816 -24608 -1782 -24573
rect -1518 -24035 -1484 -24000
rect -1518 -24107 -1484 -24083
rect -1518 -24179 -1484 -24151
rect -1518 -24251 -1484 -24219
rect -1518 -24321 -1484 -24287
rect -1518 -24389 -1484 -24357
rect -1518 -24457 -1484 -24429
rect -1518 -24525 -1484 -24501
rect -1518 -24608 -1484 -24573
rect -1220 -24035 -1186 -24000
rect -1220 -24107 -1186 -24083
rect -1220 -24179 -1186 -24151
rect -1220 -24251 -1186 -24219
rect -1220 -24321 -1186 -24287
rect -1220 -24389 -1186 -24357
rect -1220 -24457 -1186 -24429
rect -1220 -24525 -1186 -24501
rect -1220 -24608 -1186 -24573
rect -922 -24035 -888 -24000
rect -922 -24107 -888 -24083
rect -922 -24179 -888 -24151
rect -922 -24251 -888 -24219
rect -922 -24321 -888 -24287
rect -922 -24389 -888 -24357
rect -922 -24457 -888 -24429
rect -922 -24525 -888 -24501
rect -922 -24608 -888 -24573
rect -624 -24035 -590 -24000
rect -624 -24107 -590 -24083
rect -624 -24179 -590 -24151
rect -624 -24251 -590 -24219
rect -624 -24321 -590 -24287
rect -624 -24389 -590 -24357
rect -624 -24457 -590 -24429
rect -624 -24525 -590 -24501
rect -624 -24608 -590 -24573
rect -326 -24035 -292 -24000
rect -326 -24107 -292 -24083
rect -326 -24179 -292 -24151
rect -326 -24251 -292 -24219
rect -326 -24321 -292 -24287
rect -326 -24389 -292 -24357
rect -326 -24457 -292 -24429
rect -326 -24525 -292 -24501
rect -326 -24608 -292 -24573
rect -28 -24035 6 -24000
rect -28 -24107 6 -24083
rect -28 -24179 6 -24151
rect -28 -24251 6 -24219
rect -28 -24321 6 -24287
rect -28 -24389 6 -24357
rect -28 -24457 6 -24429
rect -28 -24525 6 -24501
rect -28 -24608 6 -24573
rect 270 -24035 304 -24000
rect 270 -24107 304 -24083
rect 270 -24179 304 -24151
rect 270 -24251 304 -24219
rect 270 -24321 304 -24287
rect 270 -24389 304 -24357
rect 270 -24457 304 -24429
rect 270 -24525 304 -24501
rect 270 -24608 304 -24573
rect 568 -24035 602 -24000
rect 568 -24107 602 -24083
rect 568 -24179 602 -24151
rect 568 -24251 602 -24219
rect 568 -24321 602 -24287
rect 568 -24389 602 -24357
rect 568 -24457 602 -24429
rect 568 -24525 602 -24501
rect 568 -24608 602 -24573
rect 866 -24035 900 -24000
rect 2812 -24014 2851 -23980
rect 2885 -24014 2909 -23980
rect 2953 -24014 2981 -23980
rect 3021 -24014 3053 -23980
rect 3089 -24014 3123 -23980
rect 3159 -24014 3191 -23980
rect 3231 -24014 3259 -23980
rect 3303 -24014 3327 -23980
rect 3361 -24014 3400 -23980
rect 3830 -24014 3869 -23980
rect 3903 -24014 3927 -23980
rect 3971 -24014 3999 -23980
rect 4039 -24014 4071 -23980
rect 4107 -24014 4141 -23980
rect 4177 -24014 4209 -23980
rect 4249 -24014 4277 -23980
rect 4321 -24014 4345 -23980
rect 4379 -24014 4418 -23980
rect 4848 -24014 4887 -23980
rect 4921 -24014 4945 -23980
rect 4989 -24014 5017 -23980
rect 5057 -24014 5089 -23980
rect 5125 -24014 5159 -23980
rect 5195 -24014 5227 -23980
rect 5267 -24014 5295 -23980
rect 5339 -24014 5363 -23980
rect 5397 -24014 5436 -23980
rect 5866 -24014 5905 -23980
rect 5939 -24014 5963 -23980
rect 6007 -24014 6035 -23980
rect 6075 -24014 6107 -23980
rect 6143 -24014 6177 -23980
rect 6213 -24014 6245 -23980
rect 6285 -24014 6313 -23980
rect 6357 -24014 6381 -23980
rect 6415 -24014 6454 -23980
rect 6884 -24014 6923 -23980
rect 6957 -24014 6981 -23980
rect 7025 -24014 7053 -23980
rect 7093 -24014 7125 -23980
rect 7161 -24014 7195 -23980
rect 7231 -24014 7263 -23980
rect 7303 -24014 7331 -23980
rect 7375 -24014 7399 -23980
rect 7433 -24014 7472 -23980
rect 7902 -24014 7941 -23980
rect 7975 -24014 7999 -23980
rect 8043 -24014 8071 -23980
rect 8111 -24014 8143 -23980
rect 8179 -24014 8213 -23980
rect 8249 -24014 8281 -23980
rect 8321 -24014 8349 -23980
rect 8393 -24014 8417 -23980
rect 8451 -24014 8490 -23980
rect 8920 -24014 8959 -23980
rect 8993 -24014 9017 -23980
rect 9061 -24014 9089 -23980
rect 9129 -24014 9161 -23980
rect 9197 -24014 9231 -23980
rect 9267 -24014 9299 -23980
rect 9339 -24014 9367 -23980
rect 9411 -24014 9435 -23980
rect 9469 -24014 9508 -23980
rect 9938 -24014 9977 -23980
rect 10011 -24014 10035 -23980
rect 10079 -24014 10107 -23980
rect 10147 -24014 10179 -23980
rect 10215 -24014 10249 -23980
rect 10285 -24014 10317 -23980
rect 10357 -24014 10385 -23980
rect 10429 -24014 10453 -23980
rect 10487 -24014 10526 -23980
rect 10956 -24014 10995 -23980
rect 11029 -24014 11053 -23980
rect 11097 -24014 11125 -23980
rect 11165 -24014 11197 -23980
rect 11233 -24014 11267 -23980
rect 11303 -24014 11335 -23980
rect 11375 -24014 11403 -23980
rect 11447 -24014 11471 -23980
rect 11505 -24014 11544 -23980
rect 11974 -24014 12013 -23980
rect 12047 -24014 12071 -23980
rect 12115 -24014 12143 -23980
rect 12183 -24014 12215 -23980
rect 12251 -24014 12285 -23980
rect 12321 -24014 12353 -23980
rect 12393 -24014 12421 -23980
rect 12465 -24014 12489 -23980
rect 12523 -24014 12562 -23980
rect 12992 -24014 13031 -23980
rect 13065 -24014 13089 -23980
rect 13133 -24014 13161 -23980
rect 13201 -24014 13233 -23980
rect 13269 -24014 13303 -23980
rect 13339 -24014 13371 -23980
rect 13411 -24014 13439 -23980
rect 13483 -24014 13507 -23980
rect 13541 -24014 13580 -23980
rect 14010 -24014 14049 -23980
rect 14083 -24014 14107 -23980
rect 14151 -24014 14179 -23980
rect 14219 -24014 14251 -23980
rect 14287 -24014 14321 -23980
rect 14357 -24014 14389 -23980
rect 14429 -24014 14457 -23980
rect 14501 -24014 14525 -23980
rect 14559 -24014 14598 -23980
rect 15028 -24014 15067 -23980
rect 15101 -24014 15125 -23980
rect 15169 -24014 15197 -23980
rect 15237 -24014 15269 -23980
rect 15305 -24014 15339 -23980
rect 15375 -24014 15407 -23980
rect 15447 -24014 15475 -23980
rect 15519 -24014 15543 -23980
rect 15577 -24014 15616 -23980
rect 16046 -24014 16085 -23980
rect 16119 -24014 16143 -23980
rect 16187 -24014 16215 -23980
rect 16255 -24014 16287 -23980
rect 16323 -24014 16357 -23980
rect 16393 -24014 16425 -23980
rect 16465 -24014 16493 -23980
rect 16537 -24014 16561 -23980
rect 16595 -24014 16634 -23980
rect 17064 -24014 17103 -23980
rect 17137 -24014 17161 -23980
rect 17205 -24014 17233 -23980
rect 17273 -24014 17305 -23980
rect 17341 -24014 17375 -23980
rect 17411 -24014 17443 -23980
rect 17483 -24014 17511 -23980
rect 17555 -24014 17579 -23980
rect 17613 -24014 17652 -23980
rect 18082 -24014 18121 -23980
rect 18155 -24014 18179 -23980
rect 18223 -24014 18251 -23980
rect 18291 -24014 18323 -23980
rect 18359 -24014 18393 -23980
rect 18429 -24014 18461 -23980
rect 18501 -24014 18529 -23980
rect 18573 -24014 18597 -23980
rect 18631 -24014 18670 -23980
rect 19100 -24014 19139 -23980
rect 19173 -24014 19197 -23980
rect 19241 -24014 19269 -23980
rect 19309 -24014 19341 -23980
rect 19377 -24014 19411 -23980
rect 19447 -24014 19479 -23980
rect 19519 -24014 19547 -23980
rect 19591 -24014 19615 -23980
rect 19649 -24014 19688 -23980
rect 20118 -24014 20157 -23980
rect 20191 -24014 20215 -23980
rect 20259 -24014 20287 -23980
rect 20327 -24014 20359 -23980
rect 20395 -24014 20429 -23980
rect 20465 -24014 20497 -23980
rect 20537 -24014 20565 -23980
rect 20609 -24014 20633 -23980
rect 20667 -24014 20706 -23980
rect 21136 -24014 21175 -23980
rect 21209 -24014 21233 -23980
rect 21277 -24014 21305 -23980
rect 21345 -24014 21377 -23980
rect 21413 -24014 21447 -23980
rect 21483 -24014 21515 -23980
rect 21555 -24014 21583 -23980
rect 21627 -24014 21651 -23980
rect 21685 -24014 21724 -23980
rect 22154 -24014 22193 -23980
rect 22227 -24014 22251 -23980
rect 22295 -24014 22323 -23980
rect 22363 -24014 22395 -23980
rect 22431 -24014 22465 -23980
rect 22501 -24014 22533 -23980
rect 22573 -24014 22601 -23980
rect 22645 -24014 22669 -23980
rect 22703 -24014 22742 -23980
rect 24822 -24005 24855 -23943
rect 24889 -24005 24922 -23943
rect 24822 -24011 24922 -24005
rect 9198 -24020 9258 -24014
rect 14270 -24020 14330 -24014
rect 15290 -24020 15350 -24014
rect 17326 -24020 17386 -24014
rect 866 -24107 900 -24083
rect 866 -24179 900 -24151
rect 866 -24251 900 -24219
rect 866 -24321 900 -24287
rect 866 -24389 900 -24357
rect 866 -24457 900 -24429
rect 866 -24525 900 -24501
rect 866 -24608 900 -24573
rect 2580 -24083 2614 -24048
rect 2580 -24155 2614 -24131
rect 2580 -24227 2614 -24199
rect 2580 -24299 2614 -24267
rect 2580 -24369 2614 -24335
rect 2580 -24437 2614 -24405
rect 2580 -24505 2614 -24477
rect 2580 -24573 2614 -24549
rect -12322 -24657 -12289 -24619
rect -12255 -24657 -12222 -24619
rect -7888 -24643 -7828 -24638
rect -6878 -24643 -6818 -24638
rect -5852 -24643 -5792 -24642
rect -4830 -24643 -4770 -24638
rect -12322 -24691 -12222 -24657
rect -9173 -24677 -9134 -24643
rect -9100 -24677 -9076 -24643
rect -9032 -24677 -9004 -24643
rect -8964 -24677 -8932 -24643
rect -8896 -24677 -8862 -24643
rect -8826 -24677 -8794 -24643
rect -8754 -24677 -8726 -24643
rect -8682 -24677 -8658 -24643
rect -8624 -24677 -8585 -24643
rect -8155 -24677 -8116 -24643
rect -8082 -24677 -8058 -24643
rect -8014 -24677 -7986 -24643
rect -7946 -24677 -7914 -24643
rect -7878 -24677 -7844 -24643
rect -7808 -24677 -7776 -24643
rect -7736 -24677 -7708 -24643
rect -7664 -24677 -7640 -24643
rect -7606 -24677 -7567 -24643
rect -7137 -24677 -7098 -24643
rect -7064 -24677 -7040 -24643
rect -6996 -24677 -6968 -24643
rect -6928 -24677 -6896 -24643
rect -6860 -24677 -6826 -24643
rect -6790 -24677 -6758 -24643
rect -6718 -24677 -6690 -24643
rect -6646 -24677 -6622 -24643
rect -6588 -24677 -6549 -24643
rect -6119 -24677 -6080 -24643
rect -6046 -24677 -6022 -24643
rect -5978 -24677 -5950 -24643
rect -5910 -24677 -5878 -24643
rect -5842 -24677 -5808 -24643
rect -5772 -24677 -5740 -24643
rect -5700 -24677 -5672 -24643
rect -5628 -24677 -5604 -24643
rect -5570 -24677 -5531 -24643
rect -5101 -24677 -5062 -24643
rect -5028 -24677 -5004 -24643
rect -4960 -24677 -4932 -24643
rect -4892 -24677 -4860 -24643
rect -4824 -24677 -4790 -24643
rect -4754 -24677 -4722 -24643
rect -4682 -24677 -4654 -24643
rect -4610 -24677 -4586 -24643
rect -4552 -24677 -4513 -24643
rect -4083 -24677 -4044 -24643
rect -4010 -24677 -3986 -24643
rect -3942 -24677 -3914 -24643
rect -3874 -24677 -3842 -24643
rect -3806 -24677 -3772 -24643
rect -3736 -24677 -3704 -24643
rect -3664 -24677 -3636 -24643
rect -3592 -24677 -3568 -24643
rect -3534 -24677 -3495 -24643
rect -2324 -24676 -2297 -24642
rect -2195 -24676 -2168 -24642
rect -2026 -24676 -1999 -24642
rect -1897 -24676 -1870 -24642
rect -1728 -24676 -1701 -24642
rect -1599 -24676 -1572 -24642
rect -1430 -24676 -1403 -24642
rect -1301 -24676 -1274 -24642
rect -1132 -24676 -1105 -24642
rect -1003 -24676 -976 -24642
rect -834 -24676 -807 -24642
rect -705 -24676 -678 -24642
rect -536 -24676 -509 -24642
rect -407 -24676 -380 -24642
rect -238 -24676 -211 -24642
rect -109 -24676 -82 -24642
rect 60 -24676 87 -24642
rect 189 -24676 216 -24642
rect 358 -24676 385 -24642
rect 487 -24676 514 -24642
rect 656 -24676 683 -24642
rect 785 -24676 812 -24642
rect 2580 -24656 2614 -24621
rect 3598 -24083 3632 -24048
rect 3598 -24155 3632 -24131
rect 3598 -24227 3632 -24199
rect 3598 -24299 3632 -24267
rect 3598 -24369 3632 -24335
rect 3598 -24437 3632 -24405
rect 3598 -24505 3632 -24477
rect 3598 -24573 3632 -24549
rect 3598 -24656 3632 -24621
rect 4616 -24083 4650 -24048
rect 4616 -24155 4650 -24131
rect 4616 -24227 4650 -24199
rect 4616 -24299 4650 -24267
rect 4616 -24369 4650 -24335
rect 4616 -24437 4650 -24405
rect 4616 -24505 4650 -24477
rect 4616 -24573 4650 -24549
rect 4616 -24656 4650 -24621
rect 5634 -24083 5668 -24048
rect 5634 -24155 5668 -24131
rect 5634 -24227 5668 -24199
rect 5634 -24299 5668 -24267
rect 5634 -24369 5668 -24335
rect 5634 -24437 5668 -24405
rect 5634 -24505 5668 -24477
rect 5634 -24573 5668 -24549
rect 5634 -24656 5668 -24621
rect 6652 -24083 6686 -24048
rect 6652 -24155 6686 -24131
rect 6652 -24227 6686 -24199
rect 6652 -24299 6686 -24267
rect 6652 -24369 6686 -24335
rect 6652 -24437 6686 -24405
rect 6652 -24505 6686 -24477
rect 6652 -24573 6686 -24549
rect 6652 -24656 6686 -24621
rect 7670 -24083 7704 -24048
rect 7670 -24155 7704 -24131
rect 7670 -24227 7704 -24199
rect 7670 -24299 7704 -24267
rect 7670 -24369 7704 -24335
rect 7670 -24437 7704 -24405
rect 7670 -24505 7704 -24477
rect 7670 -24573 7704 -24549
rect 7670 -24656 7704 -24621
rect 8688 -24083 8722 -24048
rect 8688 -24155 8722 -24131
rect 8688 -24227 8722 -24199
rect 8688 -24299 8722 -24267
rect 8688 -24369 8722 -24335
rect 8688 -24437 8722 -24405
rect 8688 -24505 8722 -24477
rect 8688 -24573 8722 -24549
rect 8688 -24656 8722 -24621
rect 9706 -24083 9740 -24048
rect 9706 -24155 9740 -24131
rect 9706 -24227 9740 -24199
rect 9706 -24299 9740 -24267
rect 9706 -24369 9740 -24335
rect 9706 -24437 9740 -24405
rect 9706 -24505 9740 -24477
rect 9706 -24573 9740 -24549
rect 9706 -24656 9740 -24621
rect 10724 -24083 10758 -24048
rect 10724 -24155 10758 -24131
rect 10724 -24227 10758 -24199
rect 10724 -24299 10758 -24267
rect 10724 -24369 10758 -24335
rect 10724 -24437 10758 -24405
rect 10724 -24505 10758 -24477
rect 10724 -24573 10758 -24549
rect 10724 -24656 10758 -24621
rect 11742 -24083 11776 -24048
rect 11742 -24155 11776 -24131
rect 11742 -24227 11776 -24199
rect 11742 -24299 11776 -24267
rect 11742 -24369 11776 -24335
rect 11742 -24437 11776 -24405
rect 11742 -24505 11776 -24477
rect 11742 -24573 11776 -24549
rect 11742 -24656 11776 -24621
rect 12760 -24083 12794 -24048
rect 12760 -24155 12794 -24131
rect 12760 -24227 12794 -24199
rect 12760 -24299 12794 -24267
rect 12760 -24369 12794 -24335
rect 12760 -24437 12794 -24405
rect 12760 -24505 12794 -24477
rect 12760 -24573 12794 -24549
rect 12760 -24656 12794 -24621
rect 13778 -24083 13812 -24048
rect 13778 -24155 13812 -24131
rect 13778 -24227 13812 -24199
rect 13778 -24299 13812 -24267
rect 13778 -24369 13812 -24335
rect 13778 -24437 13812 -24405
rect 13778 -24505 13812 -24477
rect 13778 -24573 13812 -24549
rect 13778 -24656 13812 -24621
rect 14796 -24083 14830 -24048
rect 14796 -24155 14830 -24131
rect 14796 -24227 14830 -24199
rect 14796 -24299 14830 -24267
rect 14796 -24369 14830 -24335
rect 14796 -24437 14830 -24405
rect 14796 -24505 14830 -24477
rect 14796 -24573 14830 -24549
rect 14796 -24656 14830 -24621
rect 15814 -24083 15848 -24048
rect 15814 -24155 15848 -24131
rect 15814 -24227 15848 -24199
rect 15814 -24299 15848 -24267
rect 15814 -24369 15848 -24335
rect 15814 -24437 15848 -24405
rect 15814 -24505 15848 -24477
rect 15814 -24573 15848 -24549
rect 15814 -24656 15848 -24621
rect 16832 -24083 16866 -24048
rect 16832 -24155 16866 -24131
rect 16832 -24227 16866 -24199
rect 16832 -24299 16866 -24267
rect 16832 -24369 16866 -24335
rect 16832 -24437 16866 -24405
rect 16832 -24505 16866 -24477
rect 16832 -24573 16866 -24549
rect 16832 -24656 16866 -24621
rect 17850 -24083 17884 -24048
rect 17850 -24155 17884 -24131
rect 17850 -24227 17884 -24199
rect 17850 -24299 17884 -24267
rect 17850 -24369 17884 -24335
rect 17850 -24437 17884 -24405
rect 17850 -24505 17884 -24477
rect 17850 -24573 17884 -24549
rect 17850 -24656 17884 -24621
rect 18868 -24083 18902 -24048
rect 18868 -24155 18902 -24131
rect 18868 -24227 18902 -24199
rect 18868 -24299 18902 -24267
rect 18868 -24369 18902 -24335
rect 18868 -24437 18902 -24405
rect 18868 -24505 18902 -24477
rect 18868 -24573 18902 -24549
rect 18868 -24656 18902 -24621
rect 19886 -24083 19920 -24048
rect 19886 -24155 19920 -24131
rect 19886 -24227 19920 -24199
rect 19886 -24299 19920 -24267
rect 19886 -24369 19920 -24335
rect 19886 -24437 19920 -24405
rect 19886 -24505 19920 -24477
rect 19886 -24573 19920 -24549
rect 19886 -24656 19920 -24621
rect 20904 -24083 20938 -24048
rect 20904 -24155 20938 -24131
rect 20904 -24227 20938 -24199
rect 20904 -24299 20938 -24267
rect 20904 -24369 20938 -24335
rect 20904 -24437 20938 -24405
rect 20904 -24505 20938 -24477
rect 20904 -24573 20938 -24549
rect 20904 -24656 20938 -24621
rect 21922 -24083 21956 -24048
rect 21922 -24155 21956 -24131
rect 21922 -24227 21956 -24199
rect 21922 -24299 21956 -24267
rect 21922 -24369 21956 -24335
rect 21922 -24437 21956 -24405
rect 21922 -24505 21956 -24477
rect 21922 -24573 21956 -24549
rect 21922 -24656 21956 -24621
rect 22940 -24083 22974 -24048
rect 22940 -24155 22974 -24131
rect 22940 -24227 22974 -24199
rect 22940 -24299 22974 -24267
rect 22940 -24369 22974 -24335
rect 22940 -24437 22974 -24405
rect 22940 -24505 22974 -24477
rect 22940 -24573 22974 -24549
rect 22940 -24656 22974 -24621
rect 24822 -24077 24855 -24011
rect 24889 -24077 24922 -24011
rect 24822 -24079 24922 -24077
rect 24822 -24113 24855 -24079
rect 24889 -24113 24922 -24079
rect 24822 -24115 24922 -24113
rect 24822 -24181 24855 -24115
rect 24889 -24181 24922 -24115
rect 24822 -24187 24922 -24181
rect 24822 -24249 24855 -24187
rect 24889 -24249 24922 -24187
rect 24822 -24259 24922 -24249
rect 24822 -24317 24855 -24259
rect 24889 -24317 24922 -24259
rect 24822 -24331 24922 -24317
rect 24822 -24385 24855 -24331
rect 24889 -24385 24922 -24331
rect 24822 -24403 24922 -24385
rect 24822 -24453 24855 -24403
rect 24889 -24453 24922 -24403
rect 24822 -24475 24922 -24453
rect 24822 -24521 24855 -24475
rect 24889 -24521 24922 -24475
rect 24822 -24547 24922 -24521
rect 24822 -24589 24855 -24547
rect 24889 -24589 24922 -24547
rect 24822 -24619 24922 -24589
rect 24822 -24657 24855 -24619
rect 24889 -24657 24922 -24619
rect 13254 -24690 13314 -24684
rect -12322 -24725 -12289 -24691
rect -12255 -24725 -12222 -24691
rect 2812 -24724 2851 -24690
rect 2885 -24724 2909 -24690
rect 2953 -24724 2981 -24690
rect 3021 -24724 3053 -24690
rect 3089 -24724 3123 -24690
rect 3159 -24724 3191 -24690
rect 3231 -24724 3259 -24690
rect 3303 -24724 3327 -24690
rect 3361 -24724 3400 -24690
rect 3830 -24724 3869 -24690
rect 3903 -24724 3927 -24690
rect 3971 -24724 3999 -24690
rect 4039 -24724 4071 -24690
rect 4107 -24724 4141 -24690
rect 4177 -24724 4209 -24690
rect 4249 -24724 4277 -24690
rect 4321 -24724 4345 -24690
rect 4379 -24724 4418 -24690
rect 4848 -24724 4887 -24690
rect 4921 -24724 4945 -24690
rect 4989 -24724 5017 -24690
rect 5057 -24724 5089 -24690
rect 5125 -24724 5159 -24690
rect 5195 -24724 5227 -24690
rect 5267 -24724 5295 -24690
rect 5339 -24724 5363 -24690
rect 5397 -24724 5436 -24690
rect 5866 -24724 5905 -24690
rect 5939 -24724 5963 -24690
rect 6007 -24724 6035 -24690
rect 6075 -24724 6107 -24690
rect 6143 -24724 6177 -24690
rect 6213 -24724 6245 -24690
rect 6285 -24724 6313 -24690
rect 6357 -24724 6381 -24690
rect 6415 -24724 6454 -24690
rect 6884 -24724 6923 -24690
rect 6957 -24724 6981 -24690
rect 7025 -24724 7053 -24690
rect 7093 -24724 7125 -24690
rect 7161 -24724 7195 -24690
rect 7231 -24724 7263 -24690
rect 7303 -24724 7331 -24690
rect 7375 -24724 7399 -24690
rect 7433 -24724 7472 -24690
rect 7902 -24724 7941 -24690
rect 7975 -24724 7999 -24690
rect 8043 -24724 8071 -24690
rect 8111 -24724 8143 -24690
rect 8179 -24724 8213 -24690
rect 8249 -24724 8281 -24690
rect 8321 -24724 8349 -24690
rect 8393 -24724 8417 -24690
rect 8451 -24724 8490 -24690
rect 8920 -24724 8959 -24690
rect 8993 -24724 9017 -24690
rect 9061 -24724 9089 -24690
rect 9129 -24724 9161 -24690
rect 9197 -24724 9231 -24690
rect 9267 -24724 9299 -24690
rect 9339 -24724 9367 -24690
rect 9411 -24724 9435 -24690
rect 9469 -24724 9508 -24690
rect 9938 -24724 9977 -24690
rect 10011 -24724 10035 -24690
rect 10079 -24724 10107 -24690
rect 10147 -24724 10179 -24690
rect 10215 -24724 10249 -24690
rect 10285 -24724 10317 -24690
rect 10357 -24724 10385 -24690
rect 10429 -24724 10453 -24690
rect 10487 -24724 10526 -24690
rect 10956 -24724 10995 -24690
rect 11029 -24724 11053 -24690
rect 11097 -24724 11125 -24690
rect 11165 -24724 11197 -24690
rect 11233 -24724 11267 -24690
rect 11303 -24724 11335 -24690
rect 11375 -24724 11403 -24690
rect 11447 -24724 11471 -24690
rect 11505 -24724 11544 -24690
rect 11974 -24724 12013 -24690
rect 12047 -24724 12071 -24690
rect 12115 -24724 12143 -24690
rect 12183 -24724 12215 -24690
rect 12251 -24724 12285 -24690
rect 12321 -24724 12353 -24690
rect 12393 -24724 12421 -24690
rect 12465 -24724 12489 -24690
rect 12523 -24724 12562 -24690
rect 12992 -24724 13031 -24690
rect 13065 -24724 13089 -24690
rect 13133 -24724 13161 -24690
rect 13201 -24724 13233 -24690
rect 13269 -24724 13303 -24690
rect 13339 -24724 13371 -24690
rect 13411 -24724 13439 -24690
rect 13483 -24724 13507 -24690
rect 13541 -24724 13580 -24690
rect 14010 -24724 14049 -24690
rect 14083 -24724 14107 -24690
rect 14151 -24724 14179 -24690
rect 14219 -24724 14251 -24690
rect 14287 -24724 14321 -24690
rect 14357 -24724 14389 -24690
rect 14429 -24724 14457 -24690
rect 14501 -24724 14525 -24690
rect 14559 -24724 14598 -24690
rect 15028 -24724 15067 -24690
rect 15101 -24724 15125 -24690
rect 15169 -24724 15197 -24690
rect 15237 -24724 15269 -24690
rect 15305 -24724 15339 -24690
rect 15375 -24724 15407 -24690
rect 15447 -24724 15475 -24690
rect 15519 -24724 15543 -24690
rect 15577 -24724 15616 -24690
rect 16046 -24724 16085 -24690
rect 16119 -24724 16143 -24690
rect 16187 -24724 16215 -24690
rect 16255 -24724 16287 -24690
rect 16323 -24724 16357 -24690
rect 16393 -24724 16425 -24690
rect 16465 -24724 16493 -24690
rect 16537 -24724 16561 -24690
rect 16595 -24724 16634 -24690
rect 17064 -24724 17103 -24690
rect 17137 -24724 17161 -24690
rect 17205 -24724 17233 -24690
rect 17273 -24724 17305 -24690
rect 17341 -24724 17375 -24690
rect 17411 -24724 17443 -24690
rect 17483 -24724 17511 -24690
rect 17555 -24724 17579 -24690
rect 17613 -24724 17652 -24690
rect 18082 -24724 18121 -24690
rect 18155 -24724 18179 -24690
rect 18223 -24724 18251 -24690
rect 18291 -24724 18323 -24690
rect 18359 -24724 18393 -24690
rect 18429 -24724 18461 -24690
rect 18501 -24724 18529 -24690
rect 18573 -24724 18597 -24690
rect 18631 -24724 18670 -24690
rect 19100 -24724 19139 -24690
rect 19173 -24724 19197 -24690
rect 19241 -24724 19269 -24690
rect 19309 -24724 19341 -24690
rect 19377 -24724 19411 -24690
rect 19447 -24724 19479 -24690
rect 19519 -24724 19547 -24690
rect 19591 -24724 19615 -24690
rect 19649 -24724 19688 -24690
rect 20118 -24724 20157 -24690
rect 20191 -24724 20215 -24690
rect 20259 -24724 20287 -24690
rect 20327 -24724 20359 -24690
rect 20395 -24724 20429 -24690
rect 20465 -24724 20497 -24690
rect 20537 -24724 20565 -24690
rect 20609 -24724 20633 -24690
rect 20667 -24724 20706 -24690
rect 21136 -24724 21175 -24690
rect 21209 -24724 21233 -24690
rect 21277 -24724 21305 -24690
rect 21345 -24724 21377 -24690
rect 21413 -24724 21447 -24690
rect 21483 -24724 21515 -24690
rect 21555 -24724 21583 -24690
rect 21627 -24724 21651 -24690
rect 21685 -24724 21724 -24690
rect 22154 -24724 22193 -24690
rect 22227 -24724 22251 -24690
rect 22295 -24724 22323 -24690
rect 22363 -24724 22395 -24690
rect 22431 -24724 22465 -24690
rect 22501 -24724 22533 -24690
rect 22573 -24724 22601 -24690
rect 22645 -24724 22669 -24690
rect 22703 -24724 22742 -24690
rect 24822 -24691 24922 -24657
rect -12322 -24759 -12222 -24725
rect -12322 -24797 -12289 -24759
rect -12255 -24797 -12222 -24759
rect -12322 -24827 -12222 -24797
rect -12322 -24869 -12289 -24827
rect -12255 -24869 -12222 -24827
rect -12322 -24895 -12222 -24869
rect -12322 -24941 -12289 -24895
rect -12255 -24941 -12222 -24895
rect -12322 -24963 -12222 -24941
rect -12322 -25013 -12289 -24963
rect -12255 -25013 -12222 -24963
rect -12322 -25031 -12222 -25013
rect -12322 -25085 -12289 -25031
rect -12255 -25085 -12222 -25031
rect 24822 -24725 24855 -24691
rect 24889 -24725 24922 -24691
rect 24822 -24759 24922 -24725
rect 24822 -24797 24855 -24759
rect 24889 -24797 24922 -24759
rect 24822 -24827 24922 -24797
rect 24822 -24869 24855 -24827
rect 24889 -24869 24922 -24827
rect 24822 -24895 24922 -24869
rect 24822 -24941 24855 -24895
rect 24889 -24941 24922 -24895
rect 24822 -24963 24922 -24941
rect 24822 -25013 24855 -24963
rect 24889 -25013 24922 -24963
rect 24822 -25031 24922 -25013
rect -9174 -25080 -9135 -25046
rect -9101 -25080 -9077 -25046
rect -9033 -25080 -9005 -25046
rect -8965 -25080 -8933 -25046
rect -8897 -25080 -8863 -25046
rect -8827 -25080 -8795 -25046
rect -8755 -25080 -8727 -25046
rect -8683 -25080 -8659 -25046
rect -8625 -25080 -8586 -25046
rect -8156 -25080 -8117 -25046
rect -8083 -25080 -8059 -25046
rect -8015 -25080 -7987 -25046
rect -7947 -25080 -7915 -25046
rect -7879 -25080 -7845 -25046
rect -7809 -25080 -7777 -25046
rect -7737 -25080 -7709 -25046
rect -7665 -25080 -7641 -25046
rect -7607 -25080 -7568 -25046
rect -7138 -25080 -7099 -25046
rect -7065 -25080 -7041 -25046
rect -6997 -25080 -6969 -25046
rect -6929 -25080 -6897 -25046
rect -6861 -25080 -6827 -25046
rect -6791 -25080 -6759 -25046
rect -6719 -25080 -6691 -25046
rect -6647 -25080 -6623 -25046
rect -6589 -25080 -6550 -25046
rect -6120 -25080 -6081 -25046
rect -6047 -25080 -6023 -25046
rect -5979 -25080 -5951 -25046
rect -5911 -25080 -5879 -25046
rect -5843 -25080 -5809 -25046
rect -5773 -25080 -5741 -25046
rect -5701 -25080 -5673 -25046
rect -5629 -25080 -5605 -25046
rect -5571 -25080 -5532 -25046
rect -5102 -25080 -5063 -25046
rect -5029 -25080 -5005 -25046
rect -4961 -25080 -4933 -25046
rect -4893 -25080 -4861 -25046
rect -4825 -25080 -4791 -25046
rect -4755 -25080 -4723 -25046
rect -4683 -25080 -4655 -25046
rect -4611 -25080 -4587 -25046
rect -4553 -25080 -4514 -25046
rect -4084 -25080 -4045 -25046
rect -4011 -25080 -3987 -25046
rect -3943 -25080 -3915 -25046
rect -3875 -25080 -3843 -25046
rect -3807 -25080 -3773 -25046
rect -3737 -25080 -3705 -25046
rect -3665 -25080 -3637 -25046
rect -3593 -25080 -3569 -25046
rect -3535 -25080 -3496 -25046
rect -2324 -25076 -2297 -25042
rect -2195 -25076 -2168 -25042
rect -2026 -25076 -1999 -25042
rect -1897 -25076 -1870 -25042
rect -1728 -25076 -1701 -25042
rect -1599 -25076 -1572 -25042
rect -1430 -25076 -1403 -25042
rect -1301 -25076 -1274 -25042
rect -1132 -25076 -1105 -25042
rect -1003 -25076 -976 -25042
rect -834 -25076 -807 -25042
rect -705 -25076 -678 -25042
rect -536 -25076 -509 -25042
rect -407 -25076 -380 -25042
rect -238 -25076 -211 -25042
rect -109 -25076 -82 -25042
rect 60 -25076 87 -25042
rect 189 -25076 216 -25042
rect 358 -25076 385 -25042
rect 487 -25076 514 -25042
rect 656 -25076 683 -25042
rect 785 -25076 812 -25042
rect -12322 -25099 -12222 -25085
rect -12322 -25157 -12289 -25099
rect -12255 -25157 -12222 -25099
rect 24822 -25085 24855 -25031
rect 24889 -25085 24922 -25031
rect 24822 -25099 24922 -25085
rect -12322 -25167 -12222 -25157
rect -12322 -25229 -12289 -25167
rect -12255 -25229 -12222 -25167
rect -12322 -25235 -12222 -25229
rect -12322 -25301 -12289 -25235
rect -12255 -25301 -12222 -25235
rect -12322 -25303 -12222 -25301
rect -12322 -25337 -12289 -25303
rect -12255 -25337 -12222 -25303
rect -12322 -25339 -12222 -25337
rect -12322 -25405 -12289 -25339
rect -12255 -25405 -12222 -25339
rect -12322 -25411 -12222 -25405
rect -12322 -25473 -12289 -25411
rect -12255 -25473 -12222 -25411
rect -12322 -25483 -12222 -25473
rect -12322 -25541 -12289 -25483
rect -12255 -25541 -12222 -25483
rect -12322 -25555 -12222 -25541
rect -12322 -25609 -12289 -25555
rect -12255 -25609 -12222 -25555
rect -12322 -25627 -12222 -25609
rect -12322 -25677 -12289 -25627
rect -12255 -25677 -12222 -25627
rect -12322 -25699 -12222 -25677
rect -12322 -25745 -12289 -25699
rect -12255 -25745 -12222 -25699
rect -9406 -25149 -9372 -25114
rect -9406 -25221 -9372 -25197
rect -9406 -25293 -9372 -25265
rect -9406 -25365 -9372 -25333
rect -9406 -25435 -9372 -25401
rect -9406 -25503 -9372 -25471
rect -9406 -25571 -9372 -25543
rect -9406 -25639 -9372 -25615
rect -9406 -25722 -9372 -25687
rect -8388 -25149 -8354 -25114
rect -8388 -25221 -8354 -25197
rect -8388 -25293 -8354 -25265
rect -8388 -25365 -8354 -25333
rect -8388 -25435 -8354 -25401
rect -8388 -25503 -8354 -25471
rect -8388 -25571 -8354 -25543
rect -8388 -25639 -8354 -25615
rect -8388 -25722 -8354 -25687
rect -7370 -25149 -7336 -25114
rect -7370 -25221 -7336 -25197
rect -7370 -25293 -7336 -25265
rect -7370 -25365 -7336 -25333
rect -7370 -25435 -7336 -25401
rect -7370 -25503 -7336 -25471
rect -7370 -25571 -7336 -25543
rect -7370 -25639 -7336 -25615
rect -7370 -25722 -7336 -25687
rect -6352 -25149 -6318 -25114
rect -6352 -25221 -6318 -25197
rect -6352 -25293 -6318 -25265
rect -6352 -25365 -6318 -25333
rect -6352 -25435 -6318 -25401
rect -6352 -25503 -6318 -25471
rect -6352 -25571 -6318 -25543
rect -6352 -25639 -6318 -25615
rect -6352 -25722 -6318 -25687
rect -5334 -25149 -5300 -25114
rect -5334 -25221 -5300 -25197
rect -5334 -25293 -5300 -25265
rect -5334 -25365 -5300 -25333
rect -5334 -25435 -5300 -25401
rect -5334 -25503 -5300 -25471
rect -5334 -25571 -5300 -25543
rect -5334 -25639 -5300 -25615
rect -5334 -25722 -5300 -25687
rect -4316 -25149 -4282 -25114
rect -4316 -25221 -4282 -25197
rect -4316 -25293 -4282 -25265
rect -4316 -25365 -4282 -25333
rect -4316 -25435 -4282 -25401
rect -4316 -25503 -4282 -25471
rect -4316 -25571 -4282 -25543
rect -4316 -25639 -4282 -25615
rect -4316 -25722 -4282 -25687
rect -3298 -25149 -3264 -25114
rect -3298 -25221 -3264 -25197
rect -3298 -25293 -3264 -25265
rect -3298 -25365 -3264 -25333
rect -3298 -25435 -3264 -25401
rect -3298 -25503 -3264 -25471
rect -3298 -25571 -3264 -25543
rect -3298 -25639 -3264 -25615
rect -3298 -25722 -3264 -25687
rect -2412 -25145 -2378 -25110
rect -2412 -25217 -2378 -25193
rect -2412 -25289 -2378 -25261
rect -2412 -25361 -2378 -25329
rect -2412 -25431 -2378 -25397
rect -2412 -25499 -2378 -25467
rect -2412 -25567 -2378 -25539
rect -2412 -25635 -2378 -25611
rect -2412 -25718 -2378 -25683
rect -2114 -25145 -2080 -25110
rect -2114 -25217 -2080 -25193
rect -2114 -25289 -2080 -25261
rect -2114 -25361 -2080 -25329
rect -2114 -25431 -2080 -25397
rect -2114 -25499 -2080 -25467
rect -2114 -25567 -2080 -25539
rect -2114 -25635 -2080 -25611
rect -2114 -25718 -2080 -25683
rect -1816 -25145 -1782 -25110
rect -1816 -25217 -1782 -25193
rect -1816 -25289 -1782 -25261
rect -1816 -25361 -1782 -25329
rect -1816 -25431 -1782 -25397
rect -1816 -25499 -1782 -25467
rect -1816 -25567 -1782 -25539
rect -1816 -25635 -1782 -25611
rect -1816 -25718 -1782 -25683
rect -1518 -25145 -1484 -25110
rect -1518 -25217 -1484 -25193
rect -1518 -25289 -1484 -25261
rect -1518 -25361 -1484 -25329
rect -1518 -25431 -1484 -25397
rect -1518 -25499 -1484 -25467
rect -1518 -25567 -1484 -25539
rect -1518 -25635 -1484 -25611
rect -1518 -25718 -1484 -25683
rect -1220 -25145 -1186 -25110
rect -1220 -25217 -1186 -25193
rect -1220 -25289 -1186 -25261
rect -1220 -25361 -1186 -25329
rect -1220 -25431 -1186 -25397
rect -1220 -25499 -1186 -25467
rect -1220 -25567 -1186 -25539
rect -1220 -25635 -1186 -25611
rect -1220 -25718 -1186 -25683
rect -922 -25145 -888 -25110
rect -922 -25217 -888 -25193
rect -922 -25289 -888 -25261
rect -922 -25361 -888 -25329
rect -922 -25431 -888 -25397
rect -922 -25499 -888 -25467
rect -922 -25567 -888 -25539
rect -922 -25635 -888 -25611
rect -922 -25718 -888 -25683
rect -624 -25145 -590 -25110
rect -624 -25217 -590 -25193
rect -624 -25289 -590 -25261
rect -624 -25361 -590 -25329
rect -624 -25431 -590 -25397
rect -624 -25499 -590 -25467
rect -624 -25567 -590 -25539
rect -624 -25635 -590 -25611
rect -624 -25718 -590 -25683
rect -326 -25145 -292 -25110
rect -326 -25217 -292 -25193
rect -326 -25289 -292 -25261
rect -326 -25361 -292 -25329
rect -326 -25431 -292 -25397
rect -326 -25499 -292 -25467
rect -326 -25567 -292 -25539
rect -326 -25635 -292 -25611
rect -326 -25718 -292 -25683
rect -28 -25145 6 -25110
rect -28 -25217 6 -25193
rect -28 -25289 6 -25261
rect -28 -25361 6 -25329
rect -28 -25431 6 -25397
rect -28 -25499 6 -25467
rect -28 -25567 6 -25539
rect -28 -25635 6 -25611
rect -28 -25718 6 -25683
rect 270 -25145 304 -25110
rect 270 -25217 304 -25193
rect 270 -25289 304 -25261
rect 270 -25361 304 -25329
rect 270 -25431 304 -25397
rect 270 -25499 304 -25467
rect 270 -25567 304 -25539
rect 270 -25635 304 -25611
rect 270 -25718 304 -25683
rect 568 -25145 602 -25110
rect 568 -25217 602 -25193
rect 568 -25289 602 -25261
rect 568 -25361 602 -25329
rect 568 -25431 602 -25397
rect 568 -25499 602 -25467
rect 568 -25567 602 -25539
rect 568 -25635 602 -25611
rect 568 -25718 602 -25683
rect 866 -25145 900 -25110
rect 866 -25217 900 -25193
rect 24822 -25157 24855 -25099
rect 24889 -25157 24922 -25099
rect 24822 -25167 24922 -25157
rect 2812 -25246 2851 -25212
rect 2885 -25246 2909 -25212
rect 2953 -25246 2981 -25212
rect 3021 -25246 3053 -25212
rect 3089 -25246 3123 -25212
rect 3159 -25246 3191 -25212
rect 3231 -25246 3259 -25212
rect 3303 -25246 3327 -25212
rect 3361 -25246 3400 -25212
rect 3830 -25246 3869 -25212
rect 3903 -25246 3927 -25212
rect 3971 -25246 3999 -25212
rect 4039 -25246 4071 -25212
rect 4107 -25246 4141 -25212
rect 4177 -25246 4209 -25212
rect 4249 -25246 4277 -25212
rect 4321 -25246 4345 -25212
rect 4379 -25246 4418 -25212
rect 4848 -25246 4887 -25212
rect 4921 -25246 4945 -25212
rect 4989 -25246 5017 -25212
rect 5057 -25246 5089 -25212
rect 5125 -25246 5159 -25212
rect 5195 -25246 5227 -25212
rect 5267 -25246 5295 -25212
rect 5339 -25246 5363 -25212
rect 5397 -25246 5436 -25212
rect 5866 -25246 5905 -25212
rect 5939 -25246 5963 -25212
rect 6007 -25246 6035 -25212
rect 6075 -25246 6107 -25212
rect 6143 -25246 6177 -25212
rect 6213 -25246 6245 -25212
rect 6285 -25246 6313 -25212
rect 6357 -25246 6381 -25212
rect 6415 -25246 6454 -25212
rect 6884 -25246 6923 -25212
rect 6957 -25246 6981 -25212
rect 7025 -25246 7053 -25212
rect 7093 -25246 7125 -25212
rect 7161 -25246 7195 -25212
rect 7231 -25246 7263 -25212
rect 7303 -25246 7331 -25212
rect 7375 -25246 7399 -25212
rect 7433 -25246 7472 -25212
rect 7902 -25246 7941 -25212
rect 7975 -25246 7999 -25212
rect 8043 -25246 8071 -25212
rect 8111 -25246 8143 -25212
rect 8179 -25246 8213 -25212
rect 8249 -25246 8281 -25212
rect 8321 -25246 8349 -25212
rect 8393 -25246 8417 -25212
rect 8451 -25246 8490 -25212
rect 8920 -25246 8959 -25212
rect 8993 -25246 9017 -25212
rect 9061 -25246 9089 -25212
rect 9129 -25246 9161 -25212
rect 9197 -25246 9231 -25212
rect 9267 -25246 9299 -25212
rect 9339 -25246 9367 -25212
rect 9411 -25246 9435 -25212
rect 9469 -25246 9508 -25212
rect 9938 -25246 9977 -25212
rect 10011 -25246 10035 -25212
rect 10079 -25246 10107 -25212
rect 10147 -25246 10179 -25212
rect 10215 -25246 10249 -25212
rect 10285 -25246 10317 -25212
rect 10357 -25246 10385 -25212
rect 10429 -25246 10453 -25212
rect 10487 -25246 10526 -25212
rect 10956 -25246 10995 -25212
rect 11029 -25246 11053 -25212
rect 11097 -25246 11125 -25212
rect 11165 -25246 11197 -25212
rect 11233 -25246 11267 -25212
rect 11303 -25246 11335 -25212
rect 11375 -25246 11403 -25212
rect 11447 -25246 11471 -25212
rect 11505 -25246 11544 -25212
rect 11974 -25246 12013 -25212
rect 12047 -25246 12071 -25212
rect 12115 -25246 12143 -25212
rect 12183 -25246 12215 -25212
rect 12251 -25246 12285 -25212
rect 12321 -25246 12353 -25212
rect 12393 -25246 12421 -25212
rect 12465 -25246 12489 -25212
rect 12523 -25246 12562 -25212
rect 12992 -25246 13031 -25212
rect 13065 -25246 13089 -25212
rect 13133 -25246 13161 -25212
rect 13201 -25246 13233 -25212
rect 13269 -25246 13303 -25212
rect 13339 -25246 13371 -25212
rect 13411 -25246 13439 -25212
rect 13483 -25246 13507 -25212
rect 13541 -25246 13580 -25212
rect 14010 -25246 14049 -25212
rect 14083 -25246 14107 -25212
rect 14151 -25246 14179 -25212
rect 14219 -25246 14251 -25212
rect 14287 -25246 14321 -25212
rect 14357 -25246 14389 -25212
rect 14429 -25246 14457 -25212
rect 14501 -25246 14525 -25212
rect 14559 -25246 14598 -25212
rect 15028 -25246 15067 -25212
rect 15101 -25246 15125 -25212
rect 15169 -25246 15197 -25212
rect 15237 -25246 15269 -25212
rect 15305 -25246 15339 -25212
rect 15375 -25246 15407 -25212
rect 15447 -25246 15475 -25212
rect 15519 -25246 15543 -25212
rect 15577 -25246 15616 -25212
rect 16046 -25246 16085 -25212
rect 16119 -25246 16143 -25212
rect 16187 -25246 16215 -25212
rect 16255 -25246 16287 -25212
rect 16323 -25246 16357 -25212
rect 16393 -25246 16425 -25212
rect 16465 -25246 16493 -25212
rect 16537 -25246 16561 -25212
rect 16595 -25246 16634 -25212
rect 17064 -25246 17103 -25212
rect 17137 -25246 17161 -25212
rect 17205 -25246 17233 -25212
rect 17273 -25246 17305 -25212
rect 17341 -25246 17375 -25212
rect 17411 -25246 17443 -25212
rect 17483 -25246 17511 -25212
rect 17555 -25246 17579 -25212
rect 17613 -25246 17652 -25212
rect 18082 -25246 18121 -25212
rect 18155 -25246 18179 -25212
rect 18223 -25246 18251 -25212
rect 18291 -25246 18323 -25212
rect 18359 -25246 18393 -25212
rect 18429 -25246 18461 -25212
rect 18501 -25246 18529 -25212
rect 18573 -25246 18597 -25212
rect 18631 -25246 18670 -25212
rect 19100 -25246 19139 -25212
rect 19173 -25246 19197 -25212
rect 19241 -25246 19269 -25212
rect 19309 -25246 19341 -25212
rect 19377 -25246 19411 -25212
rect 19447 -25246 19479 -25212
rect 19519 -25246 19547 -25212
rect 19591 -25246 19615 -25212
rect 19649 -25246 19688 -25212
rect 20118 -25246 20157 -25212
rect 20191 -25246 20215 -25212
rect 20259 -25246 20287 -25212
rect 20327 -25246 20359 -25212
rect 20395 -25246 20429 -25212
rect 20465 -25246 20497 -25212
rect 20537 -25246 20565 -25212
rect 20609 -25246 20633 -25212
rect 20667 -25246 20706 -25212
rect 21136 -25246 21175 -25212
rect 21209 -25246 21233 -25212
rect 21277 -25246 21305 -25212
rect 21345 -25246 21377 -25212
rect 21413 -25246 21447 -25212
rect 21483 -25246 21515 -25212
rect 21555 -25246 21583 -25212
rect 21627 -25246 21651 -25212
rect 21685 -25246 21724 -25212
rect 22154 -25246 22193 -25212
rect 22227 -25246 22251 -25212
rect 22295 -25246 22323 -25212
rect 22363 -25246 22395 -25212
rect 22431 -25246 22465 -25212
rect 22501 -25246 22533 -25212
rect 22573 -25246 22601 -25212
rect 22645 -25246 22669 -25212
rect 22703 -25246 22742 -25212
rect 24822 -25229 24855 -25167
rect 24889 -25229 24922 -25167
rect 24822 -25235 24922 -25229
rect 3066 -25250 3126 -25246
rect 4088 -25250 4148 -25246
rect 5114 -25250 5174 -25246
rect 6130 -25250 6190 -25246
rect 7144 -25250 7204 -25246
rect 8174 -25256 8234 -25246
rect 9190 -25256 9250 -25246
rect 10194 -25250 10254 -25246
rect 11224 -25256 11284 -25246
rect 12244 -25250 12304 -25246
rect 13254 -25250 13314 -25246
rect 14278 -25256 14338 -25246
rect 16304 -25250 16364 -25246
rect 17324 -25256 17384 -25246
rect 18348 -25250 18408 -25246
rect 21392 -25250 21452 -25246
rect 22414 -25248 22474 -25246
rect 866 -25289 900 -25261
rect 866 -25361 900 -25329
rect 866 -25431 900 -25397
rect 866 -25499 900 -25467
rect 866 -25567 900 -25539
rect 866 -25635 900 -25611
rect 866 -25718 900 -25683
rect 2580 -25315 2614 -25280
rect 2580 -25387 2614 -25363
rect 2580 -25459 2614 -25431
rect 2580 -25531 2614 -25499
rect 2580 -25601 2614 -25567
rect 2580 -25669 2614 -25637
rect -12322 -25771 -12222 -25745
rect 2580 -25737 2614 -25709
rect -12322 -25813 -12289 -25771
rect -12255 -25813 -12222 -25771
rect -9174 -25790 -9135 -25756
rect -9101 -25790 -9077 -25756
rect -9033 -25790 -9005 -25756
rect -8965 -25790 -8933 -25756
rect -8897 -25790 -8863 -25756
rect -8827 -25790 -8795 -25756
rect -8755 -25790 -8727 -25756
rect -8683 -25790 -8659 -25756
rect -8625 -25790 -8586 -25756
rect -8156 -25790 -8117 -25756
rect -8083 -25790 -8059 -25756
rect -8015 -25790 -7987 -25756
rect -7947 -25790 -7915 -25756
rect -7879 -25790 -7845 -25756
rect -7809 -25790 -7777 -25756
rect -7737 -25790 -7709 -25756
rect -7665 -25790 -7641 -25756
rect -7607 -25790 -7568 -25756
rect -7138 -25790 -7099 -25756
rect -7065 -25790 -7041 -25756
rect -6997 -25790 -6969 -25756
rect -6929 -25790 -6897 -25756
rect -6861 -25790 -6827 -25756
rect -6791 -25790 -6759 -25756
rect -6719 -25790 -6691 -25756
rect -6647 -25790 -6623 -25756
rect -6589 -25790 -6550 -25756
rect -6120 -25790 -6081 -25756
rect -6047 -25790 -6023 -25756
rect -5979 -25790 -5951 -25756
rect -5911 -25790 -5879 -25756
rect -5843 -25790 -5809 -25756
rect -5773 -25790 -5741 -25756
rect -5701 -25790 -5673 -25756
rect -5629 -25790 -5605 -25756
rect -5571 -25790 -5532 -25756
rect -5102 -25790 -5063 -25756
rect -5029 -25790 -5005 -25756
rect -4961 -25790 -4933 -25756
rect -4893 -25790 -4861 -25756
rect -4825 -25790 -4791 -25756
rect -4755 -25790 -4723 -25756
rect -4683 -25790 -4655 -25756
rect -4611 -25790 -4587 -25756
rect -4553 -25790 -4514 -25756
rect -4084 -25790 -4045 -25756
rect -4011 -25790 -3987 -25756
rect -3943 -25790 -3915 -25756
rect -3875 -25790 -3843 -25756
rect -3807 -25790 -3773 -25756
rect -3737 -25790 -3705 -25756
rect -3665 -25790 -3637 -25756
rect -3593 -25790 -3569 -25756
rect -3535 -25790 -3496 -25756
rect -2324 -25786 -2297 -25752
rect -2195 -25786 -2168 -25752
rect -2026 -25786 -1999 -25752
rect -1897 -25786 -1870 -25752
rect -1728 -25786 -1701 -25752
rect -1599 -25786 -1572 -25752
rect -1430 -25786 -1403 -25752
rect -1301 -25786 -1274 -25752
rect -1132 -25786 -1105 -25752
rect -1003 -25786 -976 -25752
rect -834 -25786 -807 -25752
rect -705 -25786 -678 -25752
rect -536 -25786 -509 -25752
rect -407 -25786 -380 -25752
rect -238 -25786 -211 -25752
rect -109 -25786 -82 -25752
rect 60 -25786 87 -25752
rect 189 -25786 216 -25752
rect 358 -25786 385 -25752
rect 487 -25786 514 -25752
rect 656 -25786 683 -25752
rect 785 -25786 812 -25752
rect -12322 -25843 -12222 -25813
rect -12322 -25881 -12289 -25843
rect -12255 -25881 -12222 -25843
rect -12322 -25915 -12222 -25881
rect 2580 -25805 2614 -25781
rect 3598 -25315 3632 -25280
rect 3598 -25387 3632 -25363
rect 3598 -25459 3632 -25431
rect 3598 -25531 3632 -25499
rect 3598 -25601 3632 -25567
rect 3598 -25669 3632 -25637
rect 3598 -25737 3632 -25709
rect 3598 -25805 3632 -25781
rect 2580 -25888 2614 -25853
rect 3582 -25853 3598 -25832
rect 4616 -25315 4650 -25280
rect 4616 -25387 4650 -25363
rect 4616 -25459 4650 -25431
rect 4616 -25531 4650 -25499
rect 4616 -25601 4650 -25567
rect 4616 -25669 4650 -25637
rect 4616 -25737 4650 -25709
rect 4616 -25805 4650 -25781
rect 3632 -25853 3642 -25832
rect 3582 -25872 3642 -25853
rect 4616 -25888 4650 -25853
rect 5634 -25315 5668 -25280
rect 5634 -25387 5668 -25363
rect 5634 -25459 5668 -25431
rect 5634 -25531 5668 -25499
rect 5634 -25601 5668 -25567
rect 5634 -25669 5668 -25637
rect 5634 -25737 5668 -25709
rect 5634 -25805 5668 -25781
rect 5634 -25872 5668 -25853
rect 6652 -25315 6686 -25280
rect 6652 -25387 6686 -25363
rect 6652 -25459 6686 -25431
rect 6652 -25531 6686 -25499
rect 6652 -25601 6686 -25567
rect 6652 -25669 6686 -25637
rect 6652 -25737 6686 -25709
rect 6652 -25805 6686 -25781
rect 7670 -25315 7704 -25280
rect 7670 -25387 7704 -25363
rect 7670 -25459 7704 -25431
rect 7670 -25531 7704 -25499
rect 7670 -25601 7704 -25567
rect 7670 -25669 7704 -25637
rect 7670 -25737 7704 -25709
rect 7670 -25805 7704 -25781
rect 6652 -25888 6686 -25853
rect 7656 -25853 7670 -25828
rect 8688 -25315 8722 -25280
rect 8688 -25387 8722 -25363
rect 8688 -25459 8722 -25431
rect 8688 -25531 8722 -25499
rect 8688 -25601 8722 -25567
rect 8688 -25669 8722 -25637
rect 8688 -25737 8722 -25709
rect 8688 -25805 8722 -25781
rect 7704 -25853 7716 -25828
rect 7656 -25872 7716 -25853
rect 8688 -25888 8722 -25853
rect 9706 -25315 9740 -25280
rect 9706 -25387 9740 -25363
rect 9706 -25459 9740 -25431
rect 9706 -25531 9740 -25499
rect 9706 -25601 9740 -25567
rect 9706 -25669 9740 -25637
rect 9706 -25737 9740 -25709
rect 9706 -25805 9740 -25781
rect 9706 -25872 9740 -25853
rect 10724 -25315 10758 -25280
rect 10724 -25387 10758 -25363
rect 10724 -25459 10758 -25431
rect 10724 -25531 10758 -25499
rect 10724 -25601 10758 -25567
rect 10724 -25669 10758 -25637
rect 10724 -25737 10758 -25709
rect 10724 -25805 10758 -25781
rect 10724 -25888 10758 -25853
rect 11742 -25315 11776 -25280
rect 11742 -25387 11776 -25363
rect 11742 -25459 11776 -25431
rect 11742 -25531 11776 -25499
rect 11742 -25601 11776 -25567
rect 11742 -25669 11776 -25637
rect 11742 -25737 11776 -25709
rect 11742 -25805 11776 -25781
rect 11742 -25872 11776 -25853
rect 12760 -25315 12794 -25280
rect 12760 -25387 12794 -25363
rect 12760 -25459 12794 -25431
rect 12760 -25531 12794 -25499
rect 12760 -25601 12794 -25567
rect 12760 -25669 12794 -25637
rect 12760 -25737 12794 -25709
rect 12760 -25805 12794 -25781
rect 13778 -25315 13812 -25280
rect 13778 -25387 13812 -25363
rect 13778 -25459 13812 -25431
rect 13778 -25531 13812 -25499
rect 13778 -25601 13812 -25567
rect 13778 -25669 13812 -25637
rect 13778 -25737 13812 -25709
rect 13778 -25805 13812 -25781
rect 12760 -25888 12794 -25853
rect 13764 -25853 13778 -25826
rect 14796 -25315 14830 -25280
rect 14796 -25387 14830 -25363
rect 14796 -25459 14830 -25431
rect 14796 -25531 14830 -25499
rect 14796 -25601 14830 -25567
rect 14796 -25669 14830 -25637
rect 14796 -25737 14830 -25709
rect 14796 -25805 14830 -25781
rect 13812 -25853 13824 -25826
rect 13764 -25872 13824 -25853
rect 14796 -25888 14830 -25853
rect 15814 -25315 15848 -25280
rect 15814 -25387 15848 -25363
rect 15814 -25459 15848 -25431
rect 15814 -25531 15848 -25499
rect 15814 -25601 15848 -25567
rect 15814 -25669 15848 -25637
rect 15814 -25737 15848 -25709
rect 15814 -25805 15848 -25781
rect 15814 -25872 15848 -25853
rect 16832 -25315 16866 -25280
rect 16832 -25387 16866 -25363
rect 16832 -25459 16866 -25431
rect 16832 -25531 16866 -25499
rect 16832 -25601 16866 -25567
rect 16832 -25669 16866 -25637
rect 16832 -25737 16866 -25709
rect 16832 -25805 16866 -25781
rect 17850 -25315 17884 -25280
rect 17850 -25387 17884 -25363
rect 17850 -25459 17884 -25431
rect 17850 -25531 17884 -25499
rect 17850 -25601 17884 -25567
rect 17850 -25669 17884 -25637
rect 17850 -25737 17884 -25709
rect 17850 -25805 17884 -25781
rect 16832 -25888 16866 -25853
rect 17836 -25853 17850 -25836
rect 18868 -25315 18902 -25280
rect 18868 -25387 18902 -25363
rect 18868 -25459 18902 -25431
rect 18868 -25531 18902 -25499
rect 18868 -25601 18902 -25567
rect 18868 -25669 18902 -25637
rect 18868 -25737 18902 -25709
rect 18868 -25805 18902 -25781
rect 17884 -25853 17896 -25836
rect 17836 -25872 17896 -25853
rect 18868 -25888 18902 -25853
rect 19886 -25315 19920 -25280
rect 19886 -25387 19920 -25363
rect 19886 -25459 19920 -25431
rect 19886 -25531 19920 -25499
rect 19886 -25601 19920 -25567
rect 19886 -25669 19920 -25637
rect 19886 -25737 19920 -25709
rect 19886 -25805 19920 -25781
rect 19886 -25872 19920 -25853
rect 20904 -25315 20938 -25280
rect 20904 -25387 20938 -25363
rect 20904 -25459 20938 -25431
rect 20904 -25531 20938 -25499
rect 20904 -25601 20938 -25567
rect 20904 -25669 20938 -25637
rect 20904 -25737 20938 -25709
rect 20904 -25805 20938 -25781
rect 21922 -25315 21956 -25280
rect 21922 -25387 21956 -25363
rect 21922 -25459 21956 -25431
rect 21922 -25531 21956 -25499
rect 21922 -25601 21956 -25567
rect 21922 -25669 21956 -25637
rect 21922 -25737 21956 -25709
rect 21922 -25805 21956 -25781
rect 20904 -25888 20938 -25853
rect 21906 -25853 21922 -25834
rect 22940 -25315 22974 -25280
rect 22940 -25387 22974 -25363
rect 22940 -25459 22974 -25431
rect 22940 -25531 22974 -25499
rect 22940 -25601 22974 -25567
rect 22940 -25669 22974 -25637
rect 22940 -25737 22974 -25709
rect 22940 -25805 22974 -25781
rect 21956 -25853 21966 -25834
rect 21906 -25872 21966 -25853
rect 22940 -25888 22974 -25853
rect 24822 -25301 24855 -25235
rect 24889 -25301 24922 -25235
rect 24822 -25303 24922 -25301
rect 24822 -25337 24855 -25303
rect 24889 -25337 24922 -25303
rect 24822 -25339 24922 -25337
rect 24822 -25405 24855 -25339
rect 24889 -25405 24922 -25339
rect 24822 -25411 24922 -25405
rect 24822 -25473 24855 -25411
rect 24889 -25473 24922 -25411
rect 24822 -25483 24922 -25473
rect 24822 -25541 24855 -25483
rect 24889 -25541 24922 -25483
rect 24822 -25555 24922 -25541
rect 24822 -25609 24855 -25555
rect 24889 -25609 24922 -25555
rect 24822 -25627 24922 -25609
rect 24822 -25677 24855 -25627
rect 24889 -25677 24922 -25627
rect 24822 -25699 24922 -25677
rect 24822 -25745 24855 -25699
rect 24889 -25745 24922 -25699
rect 24822 -25771 24922 -25745
rect 24822 -25813 24855 -25771
rect 24889 -25813 24922 -25771
rect 24822 -25843 24922 -25813
rect 24822 -25881 24855 -25843
rect 24889 -25881 24922 -25843
rect -12322 -25949 -12289 -25915
rect -12255 -25949 -12222 -25915
rect 24822 -25915 24922 -25881
rect 9186 -25922 9246 -25920
rect 15298 -25922 15358 -25920
rect 20384 -25922 20444 -25920
rect -12322 -25983 -12222 -25949
rect 2812 -25956 2851 -25922
rect 2885 -25956 2909 -25922
rect 2953 -25956 2981 -25922
rect 3021 -25956 3053 -25922
rect 3089 -25956 3123 -25922
rect 3159 -25956 3191 -25922
rect 3231 -25956 3259 -25922
rect 3303 -25956 3327 -25922
rect 3361 -25956 3400 -25922
rect 3830 -25956 3869 -25922
rect 3903 -25956 3927 -25922
rect 3971 -25956 3999 -25922
rect 4039 -25956 4071 -25922
rect 4107 -25956 4141 -25922
rect 4177 -25956 4209 -25922
rect 4249 -25956 4277 -25922
rect 4321 -25956 4345 -25922
rect 4379 -25956 4418 -25922
rect 4848 -25956 4887 -25922
rect 4921 -25956 4945 -25922
rect 4989 -25956 5017 -25922
rect 5057 -25956 5089 -25922
rect 5125 -25956 5159 -25922
rect 5195 -25956 5227 -25922
rect 5267 -25956 5295 -25922
rect 5339 -25956 5363 -25922
rect 5397 -25956 5436 -25922
rect 5866 -25956 5905 -25922
rect 5939 -25956 5963 -25922
rect 6007 -25956 6035 -25922
rect 6075 -25956 6107 -25922
rect 6143 -25956 6177 -25922
rect 6213 -25956 6245 -25922
rect 6285 -25956 6313 -25922
rect 6357 -25956 6381 -25922
rect 6415 -25956 6454 -25922
rect 6884 -25956 6923 -25922
rect 6957 -25956 6981 -25922
rect 7025 -25956 7053 -25922
rect 7093 -25956 7125 -25922
rect 7161 -25956 7195 -25922
rect 7231 -25956 7263 -25922
rect 7303 -25956 7331 -25922
rect 7375 -25956 7399 -25922
rect 7433 -25956 7472 -25922
rect 7902 -25956 7941 -25922
rect 7975 -25956 7999 -25922
rect 8043 -25956 8071 -25922
rect 8111 -25956 8143 -25922
rect 8179 -25956 8213 -25922
rect 8249 -25956 8281 -25922
rect 8321 -25956 8349 -25922
rect 8393 -25956 8417 -25922
rect 8451 -25956 8490 -25922
rect 8920 -25956 8959 -25922
rect 8993 -25956 9017 -25922
rect 9061 -25956 9089 -25922
rect 9129 -25956 9161 -25922
rect 9197 -25956 9231 -25922
rect 9267 -25956 9299 -25922
rect 9339 -25956 9367 -25922
rect 9411 -25956 9435 -25922
rect 9469 -25956 9508 -25922
rect 9938 -25956 9977 -25922
rect 10011 -25956 10035 -25922
rect 10079 -25956 10107 -25922
rect 10147 -25956 10179 -25922
rect 10215 -25956 10249 -25922
rect 10285 -25956 10317 -25922
rect 10357 -25956 10385 -25922
rect 10429 -25956 10453 -25922
rect 10487 -25956 10526 -25922
rect 10956 -25956 10995 -25922
rect 11029 -25956 11053 -25922
rect 11097 -25956 11125 -25922
rect 11165 -25956 11197 -25922
rect 11233 -25956 11267 -25922
rect 11303 -25956 11335 -25922
rect 11375 -25956 11403 -25922
rect 11447 -25956 11471 -25922
rect 11505 -25956 11544 -25922
rect 11974 -25956 12013 -25922
rect 12047 -25956 12071 -25922
rect 12115 -25956 12143 -25922
rect 12183 -25956 12215 -25922
rect 12251 -25956 12285 -25922
rect 12321 -25956 12353 -25922
rect 12393 -25956 12421 -25922
rect 12465 -25956 12489 -25922
rect 12523 -25956 12562 -25922
rect 12992 -25956 13031 -25922
rect 13065 -25956 13089 -25922
rect 13133 -25956 13161 -25922
rect 13201 -25956 13233 -25922
rect 13269 -25956 13303 -25922
rect 13339 -25956 13371 -25922
rect 13411 -25956 13439 -25922
rect 13483 -25956 13507 -25922
rect 13541 -25956 13580 -25922
rect 14010 -25956 14049 -25922
rect 14083 -25956 14107 -25922
rect 14151 -25956 14179 -25922
rect 14219 -25956 14251 -25922
rect 14287 -25956 14321 -25922
rect 14357 -25956 14389 -25922
rect 14429 -25956 14457 -25922
rect 14501 -25956 14525 -25922
rect 14559 -25956 14598 -25922
rect 15028 -25956 15067 -25922
rect 15101 -25956 15125 -25922
rect 15169 -25956 15197 -25922
rect 15237 -25956 15269 -25922
rect 15305 -25956 15339 -25922
rect 15375 -25956 15407 -25922
rect 15447 -25956 15475 -25922
rect 15519 -25956 15543 -25922
rect 15577 -25956 15616 -25922
rect 16046 -25956 16085 -25922
rect 16119 -25956 16143 -25922
rect 16187 -25956 16215 -25922
rect 16255 -25956 16287 -25922
rect 16323 -25956 16357 -25922
rect 16393 -25956 16425 -25922
rect 16465 -25956 16493 -25922
rect 16537 -25956 16561 -25922
rect 16595 -25956 16634 -25922
rect 17064 -25956 17103 -25922
rect 17137 -25956 17161 -25922
rect 17205 -25956 17233 -25922
rect 17273 -25956 17305 -25922
rect 17341 -25956 17375 -25922
rect 17411 -25956 17443 -25922
rect 17483 -25956 17511 -25922
rect 17555 -25956 17579 -25922
rect 17613 -25956 17652 -25922
rect 18082 -25956 18121 -25922
rect 18155 -25956 18179 -25922
rect 18223 -25956 18251 -25922
rect 18291 -25956 18323 -25922
rect 18359 -25956 18393 -25922
rect 18429 -25956 18461 -25922
rect 18501 -25956 18529 -25922
rect 18573 -25956 18597 -25922
rect 18631 -25956 18670 -25922
rect 19100 -25956 19139 -25922
rect 19173 -25956 19197 -25922
rect 19241 -25956 19269 -25922
rect 19309 -25956 19341 -25922
rect 19377 -25956 19411 -25922
rect 19447 -25956 19479 -25922
rect 19519 -25956 19547 -25922
rect 19591 -25956 19615 -25922
rect 19649 -25956 19688 -25922
rect 20118 -25956 20157 -25922
rect 20191 -25956 20215 -25922
rect 20259 -25956 20287 -25922
rect 20327 -25956 20359 -25922
rect 20395 -25956 20429 -25922
rect 20465 -25956 20497 -25922
rect 20537 -25956 20565 -25922
rect 20609 -25956 20633 -25922
rect 20667 -25956 20706 -25922
rect 21136 -25956 21175 -25922
rect 21209 -25956 21233 -25922
rect 21277 -25956 21305 -25922
rect 21345 -25956 21377 -25922
rect 21413 -25956 21447 -25922
rect 21483 -25956 21515 -25922
rect 21555 -25956 21583 -25922
rect 21627 -25956 21651 -25922
rect 21685 -25956 21724 -25922
rect 22154 -25956 22193 -25922
rect 22227 -25956 22251 -25922
rect 22295 -25956 22323 -25922
rect 22363 -25956 22395 -25922
rect 22431 -25956 22465 -25922
rect 22501 -25956 22533 -25922
rect 22573 -25956 22601 -25922
rect 22645 -25956 22669 -25922
rect 22703 -25956 22742 -25922
rect 24822 -25949 24855 -25915
rect 24889 -25949 24922 -25915
rect -12322 -26021 -12289 -25983
rect -12255 -26021 -12222 -25983
rect -12322 -26051 -12222 -26021
rect -12322 -26093 -12289 -26051
rect -12255 -26093 -12222 -26051
rect -12322 -26119 -12222 -26093
rect -12322 -26165 -12289 -26119
rect -12255 -26165 -12222 -26119
rect -12322 -26187 -12222 -26165
rect -12322 -26237 -12289 -26187
rect -12255 -26237 -12222 -26187
rect -12322 -26255 -12222 -26237
rect -12322 -26309 -12289 -26255
rect -12255 -26309 -12222 -26255
rect -12322 -26323 -12222 -26309
rect -12322 -26357 -12289 -26323
rect -12255 -26357 -12222 -26323
rect -12322 -26391 -12222 -26357
rect -12322 -26425 -12289 -26391
rect -12255 -26425 -12222 -26391
rect -12322 -26459 -12222 -26425
rect -12322 -26493 -12289 -26459
rect -12255 -26493 -12222 -26459
rect -12322 -26527 -12222 -26493
rect -12322 -26561 -12289 -26527
rect -12255 -26561 -12222 -26527
rect -12322 -26595 -12222 -26561
rect -12322 -26629 -12289 -26595
rect -12255 -26629 -12222 -26595
rect -12322 -26663 -12222 -26629
rect -12322 -26697 -12289 -26663
rect -12255 -26697 -12222 -26663
rect -12322 -26731 -12222 -26697
rect -12322 -26765 -12289 -26731
rect -12255 -26765 -12222 -26731
rect -12322 -26799 -12222 -26765
rect -12322 -26833 -12289 -26799
rect -12255 -26833 -12222 -26799
rect -12322 -26867 -12222 -26833
rect -12322 -26901 -12289 -26867
rect -12255 -26901 -12222 -26867
rect -12322 -26935 -12222 -26901
rect -12322 -26969 -12289 -26935
rect -12255 -26969 -12222 -26935
rect -12322 -27003 -12222 -26969
rect -12322 -27037 -12289 -27003
rect -12255 -27037 -12222 -27003
rect -12322 -27122 -12222 -27037
rect 24822 -25983 24922 -25949
rect 24822 -26021 24855 -25983
rect 24889 -26021 24922 -25983
rect 24822 -26051 24922 -26021
rect 24822 -26093 24855 -26051
rect 24889 -26093 24922 -26051
rect 24822 -26119 24922 -26093
rect 24822 -26165 24855 -26119
rect 24889 -26165 24922 -26119
rect 24822 -26187 24922 -26165
rect 24822 -26237 24855 -26187
rect 24889 -26237 24922 -26187
rect 24822 -26255 24922 -26237
rect 24822 -26309 24855 -26255
rect 24889 -26309 24922 -26255
rect 24822 -26323 24922 -26309
rect 24822 -26357 24855 -26323
rect 24889 -26357 24922 -26323
rect 24822 -26391 24922 -26357
rect 24822 -26425 24855 -26391
rect 24889 -26425 24922 -26391
rect 24822 -26459 24922 -26425
rect 24822 -26493 24855 -26459
rect 24889 -26493 24922 -26459
rect 24822 -26527 24922 -26493
rect 24822 -26561 24855 -26527
rect 24889 -26561 24922 -26527
rect 24822 -26595 24922 -26561
rect 24822 -26629 24855 -26595
rect 24889 -26629 24922 -26595
rect 24822 -26663 24922 -26629
rect 24822 -26697 24855 -26663
rect 24889 -26697 24922 -26663
rect 24822 -26731 24922 -26697
rect 24822 -26765 24855 -26731
rect 24889 -26765 24922 -26731
rect 24822 -26799 24922 -26765
rect 24822 -26833 24855 -26799
rect 24889 -26833 24922 -26799
rect 24822 -26867 24922 -26833
rect 24822 -26901 24855 -26867
rect 24889 -26901 24922 -26867
rect 24822 -26935 24922 -26901
rect 24822 -26969 24855 -26935
rect 24889 -26969 24922 -26935
rect 24822 -27003 24922 -26969
rect 24822 -27037 24855 -27003
rect 24889 -27037 24922 -27003
rect 24822 -27122 24922 -27037
rect -12322 -27155 24922 -27122
rect -12322 -27189 -12221 -27155
rect -12187 -27189 -12149 -27155
rect -12111 -27189 -12077 -27155
rect -12043 -27189 -12009 -27155
rect -11971 -27189 -11941 -27155
rect -11899 -27189 -11873 -27155
rect -11827 -27189 -11805 -27155
rect -11755 -27189 -11737 -27155
rect -11683 -27189 -11669 -27155
rect -11611 -27189 -11601 -27155
rect -11539 -27189 -11533 -27155
rect -11467 -27189 -11465 -27155
rect -11431 -27189 -11429 -27155
rect -11363 -27189 -11357 -27155
rect -11295 -27189 -11285 -27155
rect -11227 -27189 -11213 -27155
rect -11159 -27189 -11141 -27155
rect -11091 -27189 -11069 -27155
rect -11023 -27189 -10997 -27155
rect -10955 -27189 -10925 -27155
rect -10887 -27189 -10853 -27155
rect -10819 -27189 -10785 -27155
rect -10747 -27189 -10717 -27155
rect -10675 -27189 -10649 -27155
rect -10603 -27189 -10581 -27155
rect -10531 -27189 -10513 -27155
rect -10459 -27189 -10445 -27155
rect -10387 -27189 -10377 -27155
rect -10315 -27189 -10309 -27155
rect -10243 -27189 -10241 -27155
rect -10207 -27189 -10205 -27155
rect -10139 -27189 -10133 -27155
rect -10071 -27189 -10061 -27155
rect -10003 -27189 -9989 -27155
rect -9935 -27189 -9917 -27155
rect -9867 -27189 -9845 -27155
rect -9799 -27189 -9773 -27155
rect -9731 -27189 -9701 -27155
rect -9663 -27189 -9629 -27155
rect -9595 -27189 -9561 -27155
rect -9523 -27189 -9493 -27155
rect -9451 -27189 -9425 -27155
rect -9379 -27189 -9357 -27155
rect -9307 -27189 -9289 -27155
rect -9235 -27189 -9221 -27155
rect -9163 -27189 -9153 -27155
rect -9091 -27189 -9085 -27155
rect -9019 -27189 -9017 -27155
rect -8983 -27189 -8981 -27155
rect -8915 -27189 -8909 -27155
rect -8847 -27189 -8837 -27155
rect -8779 -27189 -8765 -27155
rect -8711 -27189 -8693 -27155
rect -8643 -27189 -8621 -27155
rect -8575 -27189 -8549 -27155
rect -8507 -27189 -8477 -27155
rect -8439 -27189 -8405 -27155
rect -8371 -27189 -8337 -27155
rect -8299 -27189 -8269 -27155
rect -8227 -27189 -8201 -27155
rect -8155 -27189 -8133 -27155
rect -8083 -27189 -8065 -27155
rect -8011 -27189 -7997 -27155
rect -7939 -27189 -7929 -27155
rect -7867 -27189 -7861 -27155
rect -7795 -27189 -7793 -27155
rect -7759 -27189 -7757 -27155
rect -7691 -27189 -7685 -27155
rect -7623 -27189 -7613 -27155
rect -7555 -27189 -7541 -27155
rect -7487 -27189 -7469 -27155
rect -7419 -27189 -7397 -27155
rect -7351 -27189 -7325 -27155
rect -7283 -27189 -7253 -27155
rect -7215 -27189 -7181 -27155
rect -7147 -27189 -7113 -27155
rect -7075 -27189 -7045 -27155
rect -7003 -27189 -6977 -27155
rect -6931 -27189 -6909 -27155
rect -6859 -27189 -6841 -27155
rect -6787 -27189 -6773 -27155
rect -6715 -27189 -6705 -27155
rect -6643 -27189 -6637 -27155
rect -6571 -27189 -6569 -27155
rect -6535 -27189 -6533 -27155
rect -6467 -27189 -6461 -27155
rect -6399 -27189 -6389 -27155
rect -6331 -27189 -6317 -27155
rect -6263 -27189 -6245 -27155
rect -6195 -27189 -6173 -27155
rect -6127 -27189 -6101 -27155
rect -6059 -27189 -6029 -27155
rect -5991 -27189 -5957 -27155
rect -5923 -27189 -5889 -27155
rect -5851 -27189 -5821 -27155
rect -5779 -27189 -5753 -27155
rect -5707 -27189 -5685 -27155
rect -5635 -27189 -5617 -27155
rect -5563 -27189 -5549 -27155
rect -5491 -27189 -5481 -27155
rect -5419 -27189 -5413 -27155
rect -5347 -27189 -5345 -27155
rect -5311 -27189 -5309 -27155
rect -5243 -27189 -5237 -27155
rect -5175 -27189 -5165 -27155
rect -5107 -27189 -5093 -27155
rect -5039 -27189 -5021 -27155
rect -4971 -27189 -4949 -27155
rect -4903 -27189 -4877 -27155
rect -4835 -27189 -4805 -27155
rect -4767 -27189 -4733 -27155
rect -4699 -27189 -4665 -27155
rect -4627 -27189 -4597 -27155
rect -4555 -27189 -4529 -27155
rect -4483 -27189 -4461 -27155
rect -4411 -27189 -4393 -27155
rect -4339 -27189 -4325 -27155
rect -4267 -27189 -4257 -27155
rect -4195 -27189 -4189 -27155
rect -4123 -27189 -4121 -27155
rect -4087 -27189 -4085 -27155
rect -4019 -27189 -4013 -27155
rect -3951 -27189 -3941 -27155
rect -3883 -27189 -3869 -27155
rect -3815 -27189 -3797 -27155
rect -3747 -27189 -3725 -27155
rect -3679 -27189 -3653 -27155
rect -3611 -27189 -3581 -27155
rect -3543 -27189 -3509 -27155
rect -3475 -27189 -3441 -27155
rect -3403 -27189 -3373 -27155
rect -3331 -27189 -3305 -27155
rect -3259 -27189 -3237 -27155
rect -3187 -27189 -3169 -27155
rect -3115 -27189 -3101 -27155
rect -3043 -27189 -3033 -27155
rect -2971 -27189 -2965 -27155
rect -2899 -27189 -2897 -27155
rect -2863 -27189 -2861 -27155
rect -2795 -27189 -2789 -27155
rect -2727 -27189 -2717 -27155
rect -2659 -27189 -2645 -27155
rect -2591 -27189 -2573 -27155
rect -2523 -27189 -2501 -27155
rect -2455 -27189 -2429 -27155
rect -2387 -27189 -2357 -27155
rect -2319 -27189 -2285 -27155
rect -2251 -27189 -2217 -27155
rect -2179 -27189 -2149 -27155
rect -2107 -27189 -2081 -27155
rect -2035 -27189 -2013 -27155
rect -1963 -27189 -1945 -27155
rect -1891 -27189 -1877 -27155
rect -1819 -27189 -1809 -27155
rect -1747 -27189 -1741 -27155
rect -1675 -27189 -1673 -27155
rect -1639 -27189 -1637 -27155
rect -1571 -27189 -1565 -27155
rect -1503 -27189 -1493 -27155
rect -1435 -27189 -1421 -27155
rect -1367 -27189 -1349 -27155
rect -1299 -27189 -1277 -27155
rect -1231 -27189 -1205 -27155
rect -1163 -27189 -1133 -27155
rect -1095 -27189 -1061 -27155
rect -1027 -27189 -993 -27155
rect -955 -27189 -925 -27155
rect -883 -27189 -857 -27155
rect -811 -27189 -789 -27155
rect -739 -27189 -721 -27155
rect -667 -27189 -653 -27155
rect -595 -27189 -585 -27155
rect -523 -27189 -517 -27155
rect -451 -27189 -449 -27155
rect -415 -27189 -413 -27155
rect -347 -27189 -341 -27155
rect -279 -27189 -269 -27155
rect -211 -27189 -197 -27155
rect -143 -27189 -125 -27155
rect -75 -27189 -53 -27155
rect -7 -27189 19 -27155
rect 61 -27189 91 -27155
rect 129 -27189 163 -27155
rect 197 -27189 231 -27155
rect 269 -27189 299 -27155
rect 341 -27189 367 -27155
rect 413 -27189 435 -27155
rect 485 -27189 503 -27155
rect 557 -27189 571 -27155
rect 629 -27189 639 -27155
rect 701 -27189 707 -27155
rect 773 -27189 775 -27155
rect 809 -27189 811 -27155
rect 877 -27189 883 -27155
rect 945 -27189 955 -27155
rect 1013 -27189 1027 -27155
rect 1081 -27189 1099 -27155
rect 1149 -27189 1171 -27155
rect 1217 -27189 1243 -27155
rect 1285 -27189 1315 -27155
rect 1353 -27189 1387 -27155
rect 1421 -27189 1455 -27155
rect 1493 -27189 1523 -27155
rect 1565 -27189 1591 -27155
rect 1637 -27189 1659 -27155
rect 1709 -27189 1727 -27155
rect 1781 -27189 1795 -27155
rect 1853 -27189 1863 -27155
rect 1925 -27189 1931 -27155
rect 1997 -27189 1999 -27155
rect 2033 -27189 2035 -27155
rect 2101 -27189 2107 -27155
rect 2169 -27189 2179 -27155
rect 2237 -27189 2251 -27155
rect 2305 -27189 2323 -27155
rect 2373 -27189 2395 -27155
rect 2441 -27189 2467 -27155
rect 2509 -27189 2539 -27155
rect 2577 -27189 2611 -27155
rect 2645 -27189 2679 -27155
rect 2717 -27189 2747 -27155
rect 2789 -27189 2815 -27155
rect 2861 -27189 2883 -27155
rect 2933 -27189 2951 -27155
rect 3005 -27189 3019 -27155
rect 3077 -27189 3087 -27155
rect 3149 -27189 3155 -27155
rect 3221 -27189 3223 -27155
rect 3257 -27189 3259 -27155
rect 3325 -27189 3331 -27155
rect 3393 -27189 3403 -27155
rect 3461 -27189 3475 -27155
rect 3529 -27189 3547 -27155
rect 3597 -27189 3619 -27155
rect 3665 -27189 3691 -27155
rect 3733 -27189 3763 -27155
rect 3801 -27189 3835 -27155
rect 3869 -27189 3903 -27155
rect 3941 -27189 3971 -27155
rect 4013 -27189 4039 -27155
rect 4085 -27189 4107 -27155
rect 4157 -27189 4175 -27155
rect 4229 -27189 4243 -27155
rect 4301 -27189 4311 -27155
rect 4373 -27189 4379 -27155
rect 4445 -27189 4447 -27155
rect 4481 -27189 4483 -27155
rect 4549 -27189 4555 -27155
rect 4617 -27189 4627 -27155
rect 4685 -27189 4699 -27155
rect 4753 -27189 4771 -27155
rect 4821 -27189 4843 -27155
rect 4889 -27189 4915 -27155
rect 4957 -27189 4987 -27155
rect 5025 -27189 5059 -27155
rect 5093 -27189 5127 -27155
rect 5165 -27189 5195 -27155
rect 5237 -27189 5263 -27155
rect 5309 -27189 5331 -27155
rect 5381 -27189 5399 -27155
rect 5453 -27189 5467 -27155
rect 5525 -27189 5535 -27155
rect 5597 -27189 5603 -27155
rect 5669 -27189 5671 -27155
rect 5705 -27189 5707 -27155
rect 5773 -27189 5779 -27155
rect 5841 -27189 5851 -27155
rect 5909 -27189 5923 -27155
rect 5977 -27189 5995 -27155
rect 6045 -27189 6067 -27155
rect 6113 -27189 6139 -27155
rect 6181 -27189 6211 -27155
rect 6249 -27189 6283 -27155
rect 6317 -27189 6351 -27155
rect 6389 -27189 6419 -27155
rect 6461 -27189 6487 -27155
rect 6533 -27189 6555 -27155
rect 6605 -27189 6623 -27155
rect 6677 -27189 6691 -27155
rect 6749 -27189 6759 -27155
rect 6821 -27189 6827 -27155
rect 6893 -27189 6895 -27155
rect 6929 -27189 6931 -27155
rect 6997 -27189 7003 -27155
rect 7065 -27189 7075 -27155
rect 7133 -27189 7147 -27155
rect 7201 -27189 7219 -27155
rect 7269 -27189 7291 -27155
rect 7337 -27189 7363 -27155
rect 7405 -27189 7435 -27155
rect 7473 -27189 7507 -27155
rect 7541 -27189 7575 -27155
rect 7613 -27189 7643 -27155
rect 7685 -27189 7711 -27155
rect 7757 -27189 7779 -27155
rect 7829 -27189 7847 -27155
rect 7901 -27189 7915 -27155
rect 7973 -27189 7983 -27155
rect 8045 -27189 8051 -27155
rect 8117 -27189 8119 -27155
rect 8153 -27189 8155 -27155
rect 8221 -27189 8227 -27155
rect 8289 -27189 8299 -27155
rect 8357 -27189 8371 -27155
rect 8425 -27189 8443 -27155
rect 8493 -27189 8515 -27155
rect 8561 -27189 8587 -27155
rect 8629 -27189 8659 -27155
rect 8697 -27189 8731 -27155
rect 8765 -27189 8799 -27155
rect 8837 -27189 8867 -27155
rect 8909 -27189 8935 -27155
rect 8981 -27189 9003 -27155
rect 9053 -27189 9071 -27155
rect 9125 -27189 9139 -27155
rect 9197 -27189 9207 -27155
rect 9269 -27189 9275 -27155
rect 9341 -27189 9343 -27155
rect 9377 -27189 9379 -27155
rect 9445 -27189 9451 -27155
rect 9513 -27189 9523 -27155
rect 9581 -27189 9595 -27155
rect 9649 -27189 9667 -27155
rect 9717 -27189 9739 -27155
rect 9785 -27189 9811 -27155
rect 9853 -27189 9883 -27155
rect 9921 -27189 9955 -27155
rect 9989 -27189 10023 -27155
rect 10061 -27189 10091 -27155
rect 10133 -27189 10159 -27155
rect 10205 -27189 10227 -27155
rect 10277 -27189 10295 -27155
rect 10349 -27189 10363 -27155
rect 10421 -27189 10431 -27155
rect 10493 -27189 10499 -27155
rect 10565 -27189 10567 -27155
rect 10601 -27189 10603 -27155
rect 10669 -27189 10675 -27155
rect 10737 -27189 10747 -27155
rect 10805 -27189 10819 -27155
rect 10873 -27189 10891 -27155
rect 10941 -27189 10963 -27155
rect 11009 -27189 11035 -27155
rect 11077 -27189 11107 -27155
rect 11145 -27189 11179 -27155
rect 11213 -27189 11247 -27155
rect 11285 -27189 11315 -27155
rect 11357 -27189 11383 -27155
rect 11429 -27189 11451 -27155
rect 11501 -27189 11519 -27155
rect 11573 -27189 11587 -27155
rect 11645 -27189 11655 -27155
rect 11717 -27189 11723 -27155
rect 11789 -27189 11791 -27155
rect 11825 -27189 11827 -27155
rect 11893 -27189 11899 -27155
rect 11961 -27189 11971 -27155
rect 12029 -27189 12043 -27155
rect 12097 -27189 12115 -27155
rect 12165 -27189 12187 -27155
rect 12233 -27189 12259 -27155
rect 12301 -27189 12331 -27155
rect 12369 -27189 12403 -27155
rect 12437 -27189 12471 -27155
rect 12509 -27189 12539 -27155
rect 12581 -27189 12607 -27155
rect 12653 -27189 12675 -27155
rect 12725 -27189 12743 -27155
rect 12797 -27189 12811 -27155
rect 12869 -27189 12879 -27155
rect 12941 -27189 12947 -27155
rect 13013 -27189 13015 -27155
rect 13049 -27189 13051 -27155
rect 13117 -27189 13123 -27155
rect 13185 -27189 13195 -27155
rect 13253 -27189 13267 -27155
rect 13321 -27189 13339 -27155
rect 13389 -27189 13411 -27155
rect 13457 -27189 13483 -27155
rect 13525 -27189 13555 -27155
rect 13593 -27189 13627 -27155
rect 13661 -27189 13695 -27155
rect 13733 -27189 13763 -27155
rect 13805 -27189 13831 -27155
rect 13877 -27189 13899 -27155
rect 13949 -27189 13967 -27155
rect 14021 -27189 14035 -27155
rect 14093 -27189 14103 -27155
rect 14165 -27189 14171 -27155
rect 14237 -27189 14239 -27155
rect 14273 -27189 14275 -27155
rect 14341 -27189 14347 -27155
rect 14409 -27189 14419 -27155
rect 14477 -27189 14491 -27155
rect 14545 -27189 14563 -27155
rect 14613 -27189 14635 -27155
rect 14681 -27189 14707 -27155
rect 14749 -27189 14779 -27155
rect 14817 -27189 14851 -27155
rect 14885 -27189 14919 -27155
rect 14957 -27189 14987 -27155
rect 15029 -27189 15055 -27155
rect 15101 -27189 15123 -27155
rect 15173 -27189 15191 -27155
rect 15245 -27189 15259 -27155
rect 15317 -27189 15327 -27155
rect 15389 -27189 15395 -27155
rect 15461 -27189 15463 -27155
rect 15497 -27189 15499 -27155
rect 15565 -27189 15571 -27155
rect 15633 -27189 15643 -27155
rect 15701 -27189 15715 -27155
rect 15769 -27189 15787 -27155
rect 15837 -27189 15859 -27155
rect 15905 -27189 15931 -27155
rect 15973 -27189 16003 -27155
rect 16041 -27189 16075 -27155
rect 16109 -27189 16143 -27155
rect 16181 -27189 16211 -27155
rect 16253 -27189 16279 -27155
rect 16325 -27189 16347 -27155
rect 16397 -27189 16415 -27155
rect 16469 -27189 16483 -27155
rect 16541 -27189 16551 -27155
rect 16613 -27189 16619 -27155
rect 16685 -27189 16687 -27155
rect 16721 -27189 16723 -27155
rect 16789 -27189 16795 -27155
rect 16857 -27189 16867 -27155
rect 16925 -27189 16939 -27155
rect 16993 -27189 17011 -27155
rect 17061 -27189 17083 -27155
rect 17129 -27189 17155 -27155
rect 17197 -27189 17227 -27155
rect 17265 -27189 17299 -27155
rect 17333 -27189 17367 -27155
rect 17405 -27189 17435 -27155
rect 17477 -27189 17503 -27155
rect 17549 -27189 17571 -27155
rect 17621 -27189 17639 -27155
rect 17693 -27189 17707 -27155
rect 17765 -27189 17775 -27155
rect 17837 -27189 17843 -27155
rect 17909 -27189 17911 -27155
rect 17945 -27189 17947 -27155
rect 18013 -27189 18019 -27155
rect 18081 -27189 18091 -27155
rect 18149 -27189 18163 -27155
rect 18217 -27189 18235 -27155
rect 18285 -27189 18307 -27155
rect 18353 -27189 18379 -27155
rect 18421 -27189 18451 -27155
rect 18489 -27189 18523 -27155
rect 18557 -27189 18591 -27155
rect 18629 -27189 18659 -27155
rect 18701 -27189 18727 -27155
rect 18773 -27189 18795 -27155
rect 18845 -27189 18863 -27155
rect 18917 -27189 18931 -27155
rect 18989 -27189 18999 -27155
rect 19061 -27189 19067 -27155
rect 19133 -27189 19135 -27155
rect 19169 -27189 19171 -27155
rect 19237 -27189 19243 -27155
rect 19305 -27189 19315 -27155
rect 19373 -27189 19387 -27155
rect 19441 -27189 19459 -27155
rect 19509 -27189 19531 -27155
rect 19577 -27189 19603 -27155
rect 19645 -27189 19675 -27155
rect 19713 -27189 19747 -27155
rect 19781 -27189 19815 -27155
rect 19853 -27189 19883 -27155
rect 19925 -27189 19951 -27155
rect 19997 -27189 20019 -27155
rect 20069 -27189 20087 -27155
rect 20141 -27189 20155 -27155
rect 20213 -27189 20223 -27155
rect 20285 -27189 20291 -27155
rect 20357 -27189 20359 -27155
rect 20393 -27189 20395 -27155
rect 20461 -27189 20467 -27155
rect 20529 -27189 20539 -27155
rect 20597 -27189 20611 -27155
rect 20665 -27189 20683 -27155
rect 20733 -27189 20755 -27155
rect 20801 -27189 20827 -27155
rect 20869 -27189 20899 -27155
rect 20937 -27189 20971 -27155
rect 21005 -27189 21039 -27155
rect 21077 -27189 21107 -27155
rect 21149 -27189 21175 -27155
rect 21221 -27189 21243 -27155
rect 21293 -27189 21311 -27155
rect 21365 -27189 21379 -27155
rect 21437 -27189 21447 -27155
rect 21509 -27189 21515 -27155
rect 21581 -27189 21583 -27155
rect 21617 -27189 21619 -27155
rect 21685 -27189 21691 -27155
rect 21753 -27189 21763 -27155
rect 21821 -27189 21835 -27155
rect 21889 -27189 21907 -27155
rect 21957 -27189 21979 -27155
rect 22025 -27189 22051 -27155
rect 22093 -27189 22123 -27155
rect 22161 -27189 22195 -27155
rect 22229 -27189 22263 -27155
rect 22301 -27189 22331 -27155
rect 22373 -27189 22399 -27155
rect 22445 -27189 22467 -27155
rect 22517 -27189 22535 -27155
rect 22589 -27189 22603 -27155
rect 22661 -27189 22671 -27155
rect 22733 -27189 22739 -27155
rect 22805 -27189 22807 -27155
rect 22841 -27189 22843 -27155
rect 22909 -27189 22915 -27155
rect 22977 -27189 22987 -27155
rect 23045 -27189 23059 -27155
rect 23113 -27189 23131 -27155
rect 23181 -27189 23203 -27155
rect 23249 -27189 23275 -27155
rect 23317 -27189 23347 -27155
rect 23385 -27189 23419 -27155
rect 23453 -27189 23487 -27155
rect 23525 -27189 23555 -27155
rect 23597 -27189 23623 -27155
rect 23669 -27189 23691 -27155
rect 23741 -27189 23759 -27155
rect 23813 -27189 23827 -27155
rect 23885 -27189 23895 -27155
rect 23957 -27189 23963 -27155
rect 24029 -27189 24031 -27155
rect 24065 -27189 24067 -27155
rect 24133 -27189 24139 -27155
rect 24201 -27189 24211 -27155
rect 24269 -27189 24283 -27155
rect 24337 -27189 24355 -27155
rect 24405 -27189 24427 -27155
rect 24473 -27189 24499 -27155
rect 24541 -27189 24571 -27155
rect 24609 -27189 24643 -27155
rect 24677 -27189 24711 -27155
rect 24749 -27189 24787 -27155
rect 24821 -27189 24922 -27155
rect -12322 -27222 24922 -27189
<< viali >>
rect 487 1655 521 1689
rect 559 1655 581 1689
rect 581 1655 593 1689
rect 631 1655 649 1689
rect 649 1655 665 1689
rect 703 1655 717 1689
rect 717 1655 737 1689
rect 775 1655 785 1689
rect 785 1655 809 1689
rect 847 1655 853 1689
rect 853 1655 881 1689
rect 919 1655 921 1689
rect 921 1655 953 1689
rect 991 1655 1023 1689
rect 1023 1655 1025 1689
rect 1063 1655 1091 1689
rect 1091 1655 1097 1689
rect 1135 1655 1159 1689
rect 1159 1655 1169 1689
rect 1207 1655 1227 1689
rect 1227 1655 1241 1689
rect 1279 1655 1295 1689
rect 1295 1655 1313 1689
rect 1351 1655 1363 1689
rect 1363 1655 1385 1689
rect 1423 1655 1431 1689
rect 1431 1655 1457 1689
rect 1495 1655 1499 1689
rect 1499 1655 1529 1689
rect 1567 1655 1601 1689
rect 1639 1655 1669 1689
rect 1669 1655 1673 1689
rect 1711 1655 1737 1689
rect 1737 1655 1745 1689
rect 1783 1655 1805 1689
rect 1805 1655 1817 1689
rect 1855 1655 1873 1689
rect 1873 1655 1889 1689
rect 1927 1655 1941 1689
rect 1941 1655 1961 1689
rect 1999 1655 2009 1689
rect 2009 1655 2033 1689
rect 2071 1655 2077 1689
rect 2077 1655 2105 1689
rect 2143 1655 2145 1689
rect 2145 1655 2177 1689
rect 2215 1655 2247 1689
rect 2247 1655 2249 1689
rect 2287 1655 2315 1689
rect 2315 1655 2321 1689
rect 2359 1655 2383 1689
rect 2383 1655 2393 1689
rect 2431 1655 2451 1689
rect 2451 1655 2465 1689
rect 2503 1655 2519 1689
rect 2519 1655 2537 1689
rect 2575 1655 2587 1689
rect 2587 1655 2609 1689
rect 2647 1655 2655 1689
rect 2655 1655 2681 1689
rect 2719 1655 2723 1689
rect 2723 1655 2753 1689
rect 2791 1655 2825 1689
rect 2863 1655 2893 1689
rect 2893 1655 2897 1689
rect 2935 1655 2961 1689
rect 2961 1655 2969 1689
rect 3007 1655 3029 1689
rect 3029 1655 3041 1689
rect 3079 1655 3097 1689
rect 3097 1655 3113 1689
rect 3151 1655 3165 1689
rect 3165 1655 3185 1689
rect 3223 1655 3233 1689
rect 3233 1655 3257 1689
rect 3295 1655 3301 1689
rect 3301 1655 3329 1689
rect 3367 1655 3369 1689
rect 3369 1655 3401 1689
rect 3439 1655 3471 1689
rect 3471 1655 3473 1689
rect 3511 1655 3539 1689
rect 3539 1655 3545 1689
rect 3583 1655 3607 1689
rect 3607 1655 3617 1689
rect 3655 1655 3675 1689
rect 3675 1655 3689 1689
rect 3727 1655 3743 1689
rect 3743 1655 3761 1689
rect 3799 1655 3811 1689
rect 3811 1655 3833 1689
rect 3871 1655 3879 1689
rect 3879 1655 3905 1689
rect 3943 1655 3947 1689
rect 3947 1655 3977 1689
rect 4015 1655 4049 1689
rect 4087 1655 4117 1689
rect 4117 1655 4121 1689
rect 4159 1655 4185 1689
rect 4185 1655 4193 1689
rect 4231 1655 4253 1689
rect 4253 1655 4265 1689
rect 4303 1655 4321 1689
rect 4321 1655 4337 1689
rect 4375 1655 4389 1689
rect 4389 1655 4409 1689
rect 4447 1655 4457 1689
rect 4457 1655 4481 1689
rect 4519 1655 4525 1689
rect 4525 1655 4553 1689
rect 4591 1655 4593 1689
rect 4593 1655 4625 1689
rect 4663 1655 4695 1689
rect 4695 1655 4697 1689
rect 4735 1655 4763 1689
rect 4763 1655 4769 1689
rect 4807 1655 4831 1689
rect 4831 1655 4841 1689
rect 4879 1655 4899 1689
rect 4899 1655 4913 1689
rect 4951 1655 4967 1689
rect 4967 1655 4985 1689
rect 5023 1655 5035 1689
rect 5035 1655 5057 1689
rect 5095 1655 5103 1689
rect 5103 1655 5129 1689
rect 5167 1655 5171 1689
rect 5171 1655 5201 1689
rect 5239 1655 5273 1689
rect 5311 1655 5341 1689
rect 5341 1655 5345 1689
rect 5383 1655 5409 1689
rect 5409 1655 5417 1689
rect 5455 1655 5477 1689
rect 5477 1655 5489 1689
rect 5527 1655 5545 1689
rect 5545 1655 5561 1689
rect 5599 1655 5613 1689
rect 5613 1655 5633 1689
rect 5671 1655 5681 1689
rect 5681 1655 5705 1689
rect 5743 1655 5749 1689
rect 5749 1655 5777 1689
rect 5815 1655 5817 1689
rect 5817 1655 5849 1689
rect 5887 1655 5919 1689
rect 5919 1655 5921 1689
rect 5959 1655 5987 1689
rect 5987 1655 5993 1689
rect 6031 1655 6055 1689
rect 6055 1655 6065 1689
rect 6103 1655 6123 1689
rect 6123 1655 6137 1689
rect 6175 1655 6191 1689
rect 6191 1655 6209 1689
rect 6247 1655 6259 1689
rect 6259 1655 6281 1689
rect 6319 1655 6327 1689
rect 6327 1655 6353 1689
rect 6391 1655 6395 1689
rect 6395 1655 6425 1689
rect 6463 1655 6497 1689
rect 6535 1655 6565 1689
rect 6565 1655 6569 1689
rect 6607 1655 6633 1689
rect 6633 1655 6641 1689
rect 6679 1655 6701 1689
rect 6701 1655 6713 1689
rect 6751 1655 6769 1689
rect 6769 1655 6785 1689
rect 6823 1655 6837 1689
rect 6837 1655 6857 1689
rect 6895 1655 6905 1689
rect 6905 1655 6929 1689
rect 6967 1655 6973 1689
rect 6973 1655 7001 1689
rect 7039 1655 7041 1689
rect 7041 1655 7073 1689
rect 7111 1655 7143 1689
rect 7143 1655 7145 1689
rect 7183 1655 7211 1689
rect 7211 1655 7217 1689
rect 7255 1655 7279 1689
rect 7279 1655 7289 1689
rect 7327 1655 7347 1689
rect 7347 1655 7361 1689
rect 7399 1655 7415 1689
rect 7415 1655 7433 1689
rect 7471 1655 7483 1689
rect 7483 1655 7505 1689
rect 7543 1655 7551 1689
rect 7551 1655 7577 1689
rect 7615 1655 7619 1689
rect 7619 1655 7649 1689
rect 7687 1655 7721 1689
rect 7759 1655 7789 1689
rect 7789 1655 7793 1689
rect 7831 1655 7857 1689
rect 7857 1655 7865 1689
rect 7903 1655 7925 1689
rect 7925 1655 7937 1689
rect 7975 1655 7993 1689
rect 7993 1655 8009 1689
rect 8047 1655 8061 1689
rect 8061 1655 8081 1689
rect 8119 1655 8129 1689
rect 8129 1655 8153 1689
rect 8191 1655 8197 1689
rect 8197 1655 8225 1689
rect 8263 1655 8265 1689
rect 8265 1655 8297 1689
rect 8335 1655 8367 1689
rect 8367 1655 8369 1689
rect 8407 1655 8435 1689
rect 8435 1655 8441 1689
rect 8479 1655 8503 1689
rect 8503 1655 8513 1689
rect 8551 1655 8571 1689
rect 8571 1655 8585 1689
rect 8623 1655 8639 1689
rect 8639 1655 8657 1689
rect 8695 1655 8707 1689
rect 8707 1655 8729 1689
rect 8767 1655 8775 1689
rect 8775 1655 8801 1689
rect 8839 1655 8843 1689
rect 8843 1655 8873 1689
rect 8911 1655 8945 1689
rect 8983 1655 9013 1689
rect 9013 1655 9017 1689
rect 9055 1655 9081 1689
rect 9081 1655 9089 1689
rect 9127 1655 9149 1689
rect 9149 1655 9161 1689
rect 9199 1655 9217 1689
rect 9217 1655 9233 1689
rect 9271 1655 9285 1689
rect 9285 1655 9305 1689
rect 9343 1655 9353 1689
rect 9353 1655 9377 1689
rect 9415 1655 9421 1689
rect 9421 1655 9449 1689
rect 9487 1655 9489 1689
rect 9489 1655 9521 1689
rect 9559 1655 9591 1689
rect 9591 1655 9593 1689
rect 9631 1655 9659 1689
rect 9659 1655 9665 1689
rect 9703 1655 9727 1689
rect 9727 1655 9737 1689
rect 9775 1655 9795 1689
rect 9795 1655 9809 1689
rect 9847 1655 9863 1689
rect 9863 1655 9881 1689
rect 9919 1655 9931 1689
rect 9931 1655 9953 1689
rect 9991 1655 9999 1689
rect 9999 1655 10025 1689
rect 10063 1655 10067 1689
rect 10067 1655 10097 1689
rect 10135 1655 10169 1689
rect 10207 1655 10237 1689
rect 10237 1655 10241 1689
rect 10279 1655 10305 1689
rect 10305 1655 10313 1689
rect 10351 1655 10373 1689
rect 10373 1655 10385 1689
rect 10423 1655 10441 1689
rect 10441 1655 10457 1689
rect 10495 1655 10509 1689
rect 10509 1655 10529 1689
rect 10567 1655 10577 1689
rect 10577 1655 10601 1689
rect 10639 1655 10645 1689
rect 10645 1655 10673 1689
rect 10711 1655 10713 1689
rect 10713 1655 10745 1689
rect 10783 1655 10815 1689
rect 10815 1655 10817 1689
rect 10855 1655 10883 1689
rect 10883 1655 10889 1689
rect 10927 1655 10951 1689
rect 10951 1655 10961 1689
rect 10999 1655 11019 1689
rect 11019 1655 11033 1689
rect 11071 1655 11087 1689
rect 11087 1655 11105 1689
rect 11143 1655 11155 1689
rect 11155 1655 11177 1689
rect 11215 1655 11223 1689
rect 11223 1655 11249 1689
rect 11287 1655 11291 1689
rect 11291 1655 11321 1689
rect 11359 1655 11393 1689
rect 11431 1655 11461 1689
rect 11461 1655 11465 1689
rect 11503 1655 11529 1689
rect 11529 1655 11537 1689
rect 11575 1655 11597 1689
rect 11597 1655 11609 1689
rect 11647 1655 11665 1689
rect 11665 1655 11681 1689
rect 11719 1655 11733 1689
rect 11733 1655 11753 1689
rect 11791 1655 11801 1689
rect 11801 1655 11825 1689
rect 11863 1655 11869 1689
rect 11869 1655 11897 1689
rect 11935 1655 11937 1689
rect 11937 1655 11969 1689
rect 12007 1655 12039 1689
rect 12039 1655 12041 1689
rect 12079 1655 12107 1689
rect 12107 1655 12113 1689
rect 12151 1655 12175 1689
rect 12175 1655 12185 1689
rect 12223 1655 12243 1689
rect 12243 1655 12257 1689
rect 12295 1655 12311 1689
rect 12311 1655 12329 1689
rect 12367 1655 12379 1689
rect 12379 1655 12401 1689
rect 12439 1655 12447 1689
rect 12447 1655 12473 1689
rect 12511 1655 12515 1689
rect 12515 1655 12545 1689
rect 12583 1655 12617 1689
rect 12655 1655 12685 1689
rect 12685 1655 12689 1689
rect 12727 1655 12753 1689
rect 12753 1655 12761 1689
rect 12799 1655 12821 1689
rect 12821 1655 12833 1689
rect 12871 1655 12889 1689
rect 12889 1655 12905 1689
rect 12943 1655 12957 1689
rect 12957 1655 12977 1689
rect 13015 1655 13025 1689
rect 13025 1655 13049 1689
rect 13087 1655 13093 1689
rect 13093 1655 13121 1689
rect 13159 1655 13161 1689
rect 13161 1655 13193 1689
rect 13231 1655 13263 1689
rect 13263 1655 13265 1689
rect 13303 1655 13331 1689
rect 13331 1655 13337 1689
rect 13375 1655 13399 1689
rect 13399 1655 13409 1689
rect 13447 1655 13467 1689
rect 13467 1655 13481 1689
rect 13519 1655 13535 1689
rect 13535 1655 13553 1689
rect 13591 1655 13603 1689
rect 13603 1655 13625 1689
rect 13663 1655 13671 1689
rect 13671 1655 13697 1689
rect 13735 1655 13739 1689
rect 13739 1655 13769 1689
rect 13807 1655 13841 1689
rect 13879 1655 13909 1689
rect 13909 1655 13913 1689
rect 13951 1655 13977 1689
rect 13977 1655 13985 1689
rect 14023 1655 14045 1689
rect 14045 1655 14057 1689
rect 14095 1655 14113 1689
rect 14113 1655 14129 1689
rect 14167 1655 14181 1689
rect 14181 1655 14201 1689
rect 14239 1655 14249 1689
rect 14249 1655 14273 1689
rect 14311 1655 14317 1689
rect 14317 1655 14345 1689
rect 14383 1655 14385 1689
rect 14385 1655 14417 1689
rect 14455 1655 14487 1689
rect 14487 1655 14489 1689
rect 14527 1655 14555 1689
rect 14555 1655 14561 1689
rect 14599 1655 14623 1689
rect 14623 1655 14633 1689
rect 14671 1655 14691 1689
rect 14691 1655 14705 1689
rect 14743 1655 14759 1689
rect 14759 1655 14777 1689
rect 14815 1655 14827 1689
rect 14827 1655 14849 1689
rect 14887 1655 14895 1689
rect 14895 1655 14921 1689
rect 14959 1655 14963 1689
rect 14963 1655 14993 1689
rect 15031 1655 15065 1689
rect 15103 1655 15133 1689
rect 15133 1655 15137 1689
rect 15175 1655 15201 1689
rect 15201 1655 15209 1689
rect 15247 1655 15269 1689
rect 15269 1655 15281 1689
rect 15319 1655 15337 1689
rect 15337 1655 15353 1689
rect 15391 1655 15405 1689
rect 15405 1655 15425 1689
rect 15463 1655 15473 1689
rect 15473 1655 15497 1689
rect 15535 1655 15541 1689
rect 15541 1655 15569 1689
rect 15607 1655 15609 1689
rect 15609 1655 15641 1689
rect 15679 1655 15711 1689
rect 15711 1655 15713 1689
rect 15751 1655 15779 1689
rect 15779 1655 15785 1689
rect 15823 1655 15847 1689
rect 15847 1655 15857 1689
rect 15895 1655 15915 1689
rect 15915 1655 15929 1689
rect 15967 1655 15983 1689
rect 15983 1655 16001 1689
rect 16039 1655 16051 1689
rect 16051 1655 16073 1689
rect 16111 1655 16119 1689
rect 16119 1655 16145 1689
rect 16183 1655 16187 1689
rect 16187 1655 16217 1689
rect 16255 1655 16289 1689
rect 16327 1655 16357 1689
rect 16357 1655 16361 1689
rect 16399 1655 16425 1689
rect 16425 1655 16433 1689
rect 16471 1655 16493 1689
rect 16493 1655 16505 1689
rect 16543 1655 16561 1689
rect 16561 1655 16577 1689
rect 16615 1655 16629 1689
rect 16629 1655 16649 1689
rect 16687 1655 16697 1689
rect 16697 1655 16721 1689
rect 16759 1655 16765 1689
rect 16765 1655 16793 1689
rect 16831 1655 16833 1689
rect 16833 1655 16865 1689
rect 16903 1655 16935 1689
rect 16935 1655 16937 1689
rect 16975 1655 17003 1689
rect 17003 1655 17009 1689
rect 17047 1655 17071 1689
rect 17071 1655 17081 1689
rect 17119 1655 17139 1689
rect 17139 1655 17153 1689
rect 17191 1655 17207 1689
rect 17207 1655 17225 1689
rect 17263 1655 17275 1689
rect 17275 1655 17297 1689
rect 17335 1655 17343 1689
rect 17343 1655 17369 1689
rect 17407 1655 17411 1689
rect 17411 1655 17441 1689
rect 17479 1655 17513 1689
rect 17551 1655 17581 1689
rect 17581 1655 17585 1689
rect 17623 1655 17649 1689
rect 17649 1655 17657 1689
rect 17695 1655 17717 1689
rect 17717 1655 17729 1689
rect 17767 1655 17785 1689
rect 17785 1655 17801 1689
rect 17839 1655 17853 1689
rect 17853 1655 17873 1689
rect 17911 1655 17921 1689
rect 17921 1655 17945 1689
rect 17983 1655 17989 1689
rect 17989 1655 18017 1689
rect 18055 1655 18057 1689
rect 18057 1655 18089 1689
rect 18127 1655 18159 1689
rect 18159 1655 18161 1689
rect 18199 1655 18227 1689
rect 18227 1655 18233 1689
rect 18271 1655 18295 1689
rect 18295 1655 18305 1689
rect 18343 1655 18363 1689
rect 18363 1655 18377 1689
rect 18415 1655 18431 1689
rect 18431 1655 18449 1689
rect 18487 1655 18499 1689
rect 18499 1655 18521 1689
rect 18559 1655 18567 1689
rect 18567 1655 18593 1689
rect 18631 1655 18635 1689
rect 18635 1655 18665 1689
rect 18703 1655 18737 1689
rect 18775 1655 18805 1689
rect 18805 1655 18809 1689
rect 18847 1655 18873 1689
rect 18873 1655 18881 1689
rect 18919 1655 18941 1689
rect 18941 1655 18953 1689
rect 18991 1655 19009 1689
rect 19009 1655 19025 1689
rect 19063 1655 19077 1689
rect 19077 1655 19097 1689
rect 19135 1655 19145 1689
rect 19145 1655 19169 1689
rect 19207 1655 19213 1689
rect 19213 1655 19241 1689
rect 19279 1655 19281 1689
rect 19281 1655 19313 1689
rect 19351 1655 19383 1689
rect 19383 1655 19385 1689
rect 19423 1655 19451 1689
rect 19451 1655 19457 1689
rect 19495 1655 19519 1689
rect 19519 1655 19529 1689
rect 19567 1655 19587 1689
rect 19587 1655 19601 1689
rect 19639 1655 19655 1689
rect 19655 1655 19673 1689
rect 19711 1655 19723 1689
rect 19723 1655 19745 1689
rect 19783 1655 19791 1689
rect 19791 1655 19817 1689
rect 19855 1655 19859 1689
rect 19859 1655 19889 1689
rect 19927 1655 19961 1689
rect 19999 1655 20029 1689
rect 20029 1655 20033 1689
rect 20071 1655 20097 1689
rect 20097 1655 20105 1689
rect 20143 1655 20165 1689
rect 20165 1655 20177 1689
rect 20215 1655 20233 1689
rect 20233 1655 20249 1689
rect 20287 1655 20301 1689
rect 20301 1655 20321 1689
rect 20359 1655 20369 1689
rect 20369 1655 20393 1689
rect 20431 1655 20437 1689
rect 20437 1655 20465 1689
rect 20503 1655 20505 1689
rect 20505 1655 20537 1689
rect 20575 1655 20607 1689
rect 20607 1655 20609 1689
rect 20647 1655 20675 1689
rect 20675 1655 20681 1689
rect 20719 1655 20743 1689
rect 20743 1655 20753 1689
rect 20791 1655 20811 1689
rect 20811 1655 20825 1689
rect 20863 1655 20879 1689
rect 20879 1655 20897 1689
rect 20935 1655 20947 1689
rect 20947 1655 20969 1689
rect 21007 1655 21015 1689
rect 21015 1655 21041 1689
rect 21079 1655 21083 1689
rect 21083 1655 21113 1689
rect 21151 1655 21185 1689
rect 21223 1655 21253 1689
rect 21253 1655 21257 1689
rect 21295 1655 21321 1689
rect 21321 1655 21329 1689
rect 21367 1655 21389 1689
rect 21389 1655 21401 1689
rect 21439 1655 21457 1689
rect 21457 1655 21473 1689
rect 21511 1655 21525 1689
rect 21525 1655 21545 1689
rect 21583 1655 21593 1689
rect 21593 1655 21617 1689
rect 21655 1655 21661 1689
rect 21661 1655 21689 1689
rect 21727 1655 21729 1689
rect 21729 1655 21761 1689
rect 21799 1655 21831 1689
rect 21831 1655 21833 1689
rect 21871 1655 21899 1689
rect 21899 1655 21905 1689
rect 21943 1655 21967 1689
rect 21967 1655 21977 1689
rect 22015 1655 22035 1689
rect 22035 1655 22049 1689
rect 22087 1655 22103 1689
rect 22103 1655 22121 1689
rect 22159 1655 22171 1689
rect 22171 1655 22193 1689
rect 22231 1655 22239 1689
rect 22239 1655 22265 1689
rect 22303 1655 22307 1689
rect 22307 1655 22337 1689
rect 22375 1655 22409 1689
rect 22447 1655 22477 1689
rect 22477 1655 22481 1689
rect 22519 1655 22545 1689
rect 22545 1655 22553 1689
rect 22591 1655 22613 1689
rect 22613 1655 22625 1689
rect 22663 1655 22681 1689
rect 22681 1655 22697 1689
rect 22735 1655 22749 1689
rect 22749 1655 22769 1689
rect 22807 1655 22817 1689
rect 22817 1655 22841 1689
rect 22879 1655 22885 1689
rect 22885 1655 22913 1689
rect 22951 1655 22953 1689
rect 22953 1655 22985 1689
rect 23023 1655 23055 1689
rect 23055 1655 23057 1689
rect 23095 1655 23123 1689
rect 23123 1655 23129 1689
rect 23167 1655 23191 1689
rect 23191 1655 23201 1689
rect 23239 1655 23259 1689
rect 23259 1655 23273 1689
rect 23311 1655 23327 1689
rect 23327 1655 23345 1689
rect 23383 1655 23395 1689
rect 23395 1655 23417 1689
rect 23455 1655 23463 1689
rect 23463 1655 23489 1689
rect 23527 1655 23531 1689
rect 23531 1655 23561 1689
rect 23599 1655 23633 1689
rect 23671 1655 23701 1689
rect 23701 1655 23705 1689
rect 23743 1655 23769 1689
rect 23769 1655 23777 1689
rect 23815 1655 23837 1689
rect 23837 1655 23849 1689
rect 23887 1655 23905 1689
rect 23905 1655 23921 1689
rect 23959 1655 23973 1689
rect 23973 1655 23993 1689
rect 24031 1655 24041 1689
rect 24041 1655 24065 1689
rect 24103 1655 24109 1689
rect 24109 1655 24137 1689
rect 24175 1655 24177 1689
rect 24177 1655 24209 1689
rect 24247 1655 24279 1689
rect 24279 1655 24281 1689
rect 24319 1655 24347 1689
rect 24347 1655 24353 1689
rect 24391 1655 24415 1689
rect 24415 1655 24425 1689
rect 24463 1655 24483 1689
rect 24483 1655 24497 1689
rect 24535 1655 24551 1689
rect 24551 1655 24569 1689
rect 24607 1655 24619 1689
rect 24619 1655 24641 1689
rect 24679 1655 24713 1689
rect 411 1061 445 1081
rect 411 1047 445 1061
rect 411 993 445 1009
rect 411 975 445 993
rect 411 925 445 937
rect 411 903 445 925
rect 411 857 445 865
rect 411 831 445 857
rect 411 789 445 793
rect 411 759 445 789
rect 411 687 445 721
rect 411 619 445 649
rect 411 615 445 619
rect 411 551 445 577
rect 411 543 445 551
rect 411 483 445 505
rect 411 471 445 483
rect 411 415 445 433
rect 411 399 445 415
rect 411 347 445 361
rect 411 327 445 347
rect 411 279 445 289
rect 411 255 445 279
rect 411 211 445 217
rect 411 183 445 211
rect 411 143 445 145
rect 411 111 445 143
rect 411 41 445 73
rect 411 39 445 41
rect 411 -27 445 1
rect 411 -33 445 -27
rect 411 -95 445 -71
rect 411 -105 445 -95
rect 411 -163 445 -143
rect 411 -177 445 -163
rect 411 -231 445 -215
rect 411 -249 445 -231
rect 411 -299 445 -287
rect 411 -321 445 -299
rect 411 -367 445 -359
rect 411 -393 445 -367
rect 411 -435 445 -431
rect 411 -465 445 -435
rect 411 -537 445 -503
rect 411 -605 445 -575
rect 411 -609 445 -605
rect 411 -673 445 -647
rect 411 -681 445 -673
rect 411 -741 445 -719
rect 411 -753 445 -741
rect 411 -809 445 -791
rect 411 -825 445 -809
rect 411 -877 445 -863
rect 411 -897 445 -877
rect 411 -945 445 -935
rect 411 -969 445 -945
rect 411 -1013 445 -1007
rect 411 -1041 445 -1013
rect 411 -1081 445 -1079
rect 411 -1113 445 -1081
rect 411 -1183 445 -1151
rect 411 -1185 445 -1183
rect 411 -1251 445 -1223
rect 411 -1257 445 -1251
rect 411 -1319 445 -1295
rect 411 -1329 445 -1319
rect 411 -1387 445 -1367
rect 411 -1401 445 -1387
rect 411 -1455 445 -1439
rect 411 -1473 445 -1455
rect 411 -1523 445 -1511
rect 411 -1545 445 -1523
rect 411 -1591 445 -1583
rect 411 -1617 445 -1591
rect 411 -1659 445 -1655
rect 411 -1689 445 -1659
rect 411 -1761 445 -1727
rect 411 -1829 445 -1799
rect 411 -1833 445 -1829
rect 411 -1897 445 -1871
rect 411 -1905 445 -1897
rect 411 -1965 445 -1943
rect 411 -1977 445 -1965
rect 411 -2033 445 -2015
rect 411 -2049 445 -2033
rect 411 -2101 445 -2087
rect 411 -2121 445 -2101
rect 411 -2169 445 -2159
rect 411 -2193 445 -2169
rect 411 -2237 445 -2231
rect 411 -2265 445 -2237
rect 411 -2305 445 -2303
rect 411 -2337 445 -2305
rect 411 -2407 445 -2375
rect 411 -2409 445 -2407
rect 411 -2475 445 -2447
rect 411 -2481 445 -2475
rect 411 -2543 445 -2519
rect 411 -2553 445 -2543
rect 411 -2611 445 -2591
rect 411 -2625 445 -2611
rect 411 -2679 445 -2663
rect 411 -2697 445 -2679
rect 411 -2747 445 -2735
rect 411 -2769 445 -2747
rect 411 -2815 445 -2807
rect 411 -2841 445 -2815
rect 411 -2883 445 -2879
rect 411 -2913 445 -2883
rect 411 -2985 445 -2951
rect 411 -3053 445 -3023
rect 411 -3057 445 -3053
rect 411 -3121 445 -3095
rect 411 -3129 445 -3121
rect 411 -3189 445 -3167
rect 411 -3201 445 -3189
rect 411 -3257 445 -3239
rect 411 -3273 445 -3257
rect 411 -3325 445 -3311
rect 411 -3345 445 -3325
rect 411 -3393 445 -3383
rect 411 -3417 445 -3393
rect 411 -3461 445 -3455
rect 411 -3489 445 -3461
rect 411 -3529 445 -3527
rect 411 -3561 445 -3529
rect 411 -3631 445 -3599
rect 411 -3633 445 -3631
rect 411 -3699 445 -3671
rect 411 -3705 445 -3699
rect 411 -3767 445 -3743
rect 411 -3777 445 -3767
rect 411 -3835 445 -3815
rect 411 -3849 445 -3835
rect 411 -3903 445 -3887
rect 411 -3921 445 -3903
rect 411 -3971 445 -3959
rect 411 -3993 445 -3971
rect 411 -4039 445 -4031
rect 411 -4065 445 -4039
rect 411 -4107 445 -4103
rect 411 -4137 445 -4107
rect 411 -4209 445 -4175
rect 411 -4277 445 -4247
rect 411 -4281 445 -4277
rect 411 -4345 445 -4319
rect 411 -4353 445 -4345
rect 411 -4413 445 -4391
rect 411 -4425 445 -4413
rect 411 -4481 445 -4463
rect 411 -4497 445 -4481
rect 411 -4549 445 -4535
rect 411 -4569 445 -4549
rect 411 -4617 445 -4607
rect 411 -4641 445 -4617
rect 24755 1061 24789 1081
rect 24755 1047 24789 1061
rect 24755 993 24789 1009
rect 24755 975 24789 993
rect 24755 925 24789 937
rect 24755 903 24789 925
rect 24755 857 24789 865
rect 24755 831 24789 857
rect 24755 789 24789 793
rect 24755 759 24789 789
rect 24755 687 24789 721
rect 24755 619 24789 649
rect 24755 615 24789 619
rect 24755 551 24789 577
rect 24755 543 24789 551
rect 24755 483 24789 505
rect 24755 471 24789 483
rect 24755 415 24789 433
rect 24755 399 24789 415
rect 24755 347 24789 361
rect 24755 327 24789 347
rect 24755 279 24789 289
rect 24755 255 24789 279
rect 24755 211 24789 217
rect 24755 183 24789 211
rect 24755 143 24789 145
rect 24755 111 24789 143
rect 24755 41 24789 73
rect 24755 39 24789 41
rect 24755 -27 24789 1
rect 24755 -33 24789 -27
rect 24755 -95 24789 -71
rect 24755 -105 24789 -95
rect 24755 -163 24789 -143
rect 24755 -177 24789 -163
rect 24755 -231 24789 -215
rect 24755 -249 24789 -231
rect 24755 -299 24789 -287
rect 24755 -321 24789 -299
rect 24755 -367 24789 -359
rect 24755 -393 24789 -367
rect 24755 -435 24789 -431
rect 24755 -465 24789 -435
rect 24755 -537 24789 -503
rect 24755 -605 24789 -575
rect 24755 -609 24789 -605
rect 24755 -673 24789 -647
rect 24755 -681 24789 -673
rect 24755 -741 24789 -719
rect 24755 -753 24789 -741
rect 24755 -809 24789 -791
rect 24755 -825 24789 -809
rect 24755 -877 24789 -863
rect 24755 -897 24789 -877
rect 24755 -945 24789 -935
rect 24755 -969 24789 -945
rect 24755 -1013 24789 -1007
rect 24755 -1041 24789 -1013
rect 24755 -1081 24789 -1079
rect 24755 -1113 24789 -1081
rect 24755 -1183 24789 -1151
rect 24755 -1185 24789 -1183
rect 24755 -1251 24789 -1223
rect 24755 -1257 24789 -1251
rect 24755 -1319 24789 -1295
rect 24755 -1329 24789 -1319
rect 24755 -1387 24789 -1367
rect 24755 -1401 24789 -1387
rect 24755 -1455 24789 -1439
rect 24755 -1473 24789 -1455
rect 24755 -1523 24789 -1511
rect 24755 -1545 24789 -1523
rect 24755 -1591 24789 -1583
rect 24755 -1617 24789 -1591
rect 24755 -1659 24789 -1655
rect 24755 -1689 24789 -1659
rect 24755 -1761 24789 -1727
rect 24755 -1829 24789 -1799
rect 24755 -1833 24789 -1829
rect 24755 -1897 24789 -1871
rect 24755 -1905 24789 -1897
rect 24755 -1965 24789 -1943
rect 24755 -1977 24789 -1965
rect 24755 -2033 24789 -2015
rect 24755 -2049 24789 -2033
rect 24755 -2101 24789 -2087
rect 24755 -2121 24789 -2101
rect 24755 -2169 24789 -2159
rect 24755 -2193 24789 -2169
rect 24755 -2237 24789 -2231
rect 24755 -2265 24789 -2237
rect 24755 -2305 24789 -2303
rect 24755 -2337 24789 -2305
rect 24755 -2407 24789 -2375
rect 24755 -2409 24789 -2407
rect 24755 -2475 24789 -2447
rect 24755 -2481 24789 -2475
rect 24755 -2543 24789 -2519
rect 24755 -2553 24789 -2543
rect 24755 -2611 24789 -2591
rect 24755 -2625 24789 -2611
rect 24755 -2679 24789 -2663
rect 24755 -2697 24789 -2679
rect 24755 -2747 24789 -2735
rect 24755 -2769 24789 -2747
rect 24755 -2815 24789 -2807
rect 24755 -2841 24789 -2815
rect 24755 -2883 24789 -2879
rect 24755 -2913 24789 -2883
rect 24755 -2985 24789 -2951
rect 24755 -3053 24789 -3023
rect 24755 -3057 24789 -3053
rect 24755 -3121 24789 -3095
rect 24755 -3129 24789 -3121
rect 24755 -3189 24789 -3167
rect 24755 -3201 24789 -3189
rect 24755 -3257 24789 -3239
rect 24755 -3273 24789 -3257
rect 24755 -3325 24789 -3311
rect 24755 -3345 24789 -3325
rect 24755 -3393 24789 -3383
rect 24755 -3417 24789 -3393
rect 24755 -3461 24789 -3455
rect 24755 -3489 24789 -3461
rect 24755 -3529 24789 -3527
rect 24755 -3561 24789 -3529
rect 24755 -3631 24789 -3599
rect 24755 -3633 24789 -3631
rect 24755 -3699 24789 -3671
rect 24755 -3705 24789 -3699
rect 24755 -3767 24789 -3743
rect 24755 -3777 24789 -3767
rect 24755 -3835 24789 -3815
rect 24755 -3849 24789 -3835
rect 24755 -3903 24789 -3887
rect 24755 -3921 24789 -3903
rect 24755 -3971 24789 -3959
rect 24755 -3993 24789 -3971
rect 24755 -4039 24789 -4031
rect 24755 -4065 24789 -4039
rect 24755 -4107 24789 -4103
rect 24755 -4137 24789 -4107
rect 24755 -4209 24789 -4175
rect 24755 -4277 24789 -4247
rect 24755 -4281 24789 -4277
rect 24755 -4345 24789 -4319
rect 24755 -4353 24789 -4345
rect 24755 -4413 24789 -4391
rect 24755 -4425 24789 -4413
rect 24755 -4481 24789 -4463
rect 24755 -4497 24789 -4481
rect 24755 -4549 24789 -4535
rect 24755 -4569 24789 -4549
rect 3735 -4643 3769 -4609
rect 3953 -4643 3987 -4609
rect 4171 -4643 4205 -4609
rect 4389 -4643 4423 -4609
rect 4607 -4643 4641 -4609
rect 4825 -4643 4859 -4609
rect 5043 -4643 5077 -4609
rect 5261 -4643 5295 -4609
rect 5479 -4643 5513 -4609
rect 5697 -4643 5731 -4609
rect 24755 -4617 24789 -4607
rect 24755 -4641 24789 -4617
rect 411 -4685 445 -4679
rect 411 -4713 445 -4685
rect 411 -4753 445 -4751
rect 411 -4785 445 -4753
rect 411 -4855 445 -4823
rect 411 -4857 445 -4855
rect 411 -4923 445 -4895
rect 411 -4929 445 -4923
rect 411 -4991 445 -4967
rect 411 -5001 445 -4991
rect 411 -5059 445 -5039
rect 411 -5073 445 -5059
rect 3626 -4737 3660 -4729
rect 3626 -4763 3660 -4737
rect 3626 -4805 3660 -4801
rect 3626 -4835 3660 -4805
rect 3626 -4907 3660 -4873
rect 3626 -4975 3660 -4945
rect 3626 -4979 3660 -4975
rect 3626 -5043 3660 -5017
rect 3626 -5051 3660 -5043
rect 3844 -4737 3878 -4729
rect 3844 -4763 3878 -4737
rect 3844 -4805 3878 -4801
rect 3844 -4835 3878 -4805
rect 3844 -4907 3878 -4873
rect 3844 -4975 3878 -4945
rect 3844 -4979 3878 -4975
rect 3844 -5043 3878 -5017
rect 3844 -5051 3878 -5043
rect 4062 -4737 4096 -4729
rect 4062 -4763 4096 -4737
rect 4062 -4805 4096 -4801
rect 4062 -4835 4096 -4805
rect 4062 -4907 4096 -4873
rect 4062 -4975 4096 -4945
rect 4062 -4979 4096 -4975
rect 4062 -5043 4096 -5017
rect 4062 -5051 4096 -5043
rect 4280 -4737 4314 -4729
rect 4280 -4763 4314 -4737
rect 4280 -4805 4314 -4801
rect 4280 -4835 4314 -4805
rect 4280 -4907 4314 -4873
rect 4280 -4975 4314 -4945
rect 4280 -4979 4314 -4975
rect 4280 -5043 4314 -5017
rect 4280 -5051 4314 -5043
rect 4498 -4737 4532 -4729
rect 4498 -4763 4532 -4737
rect 4498 -4805 4532 -4801
rect 4498 -4835 4532 -4805
rect 4498 -4907 4532 -4873
rect 4498 -4975 4532 -4945
rect 4498 -4979 4532 -4975
rect 4498 -5043 4532 -5017
rect 4498 -5051 4532 -5043
rect 4716 -4737 4750 -4729
rect 4716 -4763 4750 -4737
rect 4716 -4805 4750 -4801
rect 4716 -4835 4750 -4805
rect 4716 -4907 4750 -4873
rect 4716 -4975 4750 -4945
rect 4716 -4979 4750 -4975
rect 4716 -5043 4750 -5017
rect 4716 -5051 4750 -5043
rect 4934 -4737 4968 -4729
rect 4934 -4763 4968 -4737
rect 4934 -4805 4968 -4801
rect 4934 -4835 4968 -4805
rect 4934 -4907 4968 -4873
rect 4934 -4975 4968 -4945
rect 4934 -4979 4968 -4975
rect 4934 -5043 4968 -5017
rect 4934 -5051 4968 -5043
rect 5152 -4737 5186 -4729
rect 5152 -4763 5186 -4737
rect 5152 -4805 5186 -4801
rect 5152 -4835 5186 -4805
rect 5152 -4907 5186 -4873
rect 5152 -4975 5186 -4945
rect 5152 -4979 5186 -4975
rect 5152 -5043 5186 -5017
rect 5152 -5051 5186 -5043
rect 5370 -4737 5404 -4729
rect 5370 -4763 5404 -4737
rect 5370 -4805 5404 -4801
rect 5370 -4835 5404 -4805
rect 5370 -4907 5404 -4873
rect 5370 -4975 5404 -4945
rect 5370 -4979 5404 -4975
rect 5370 -5043 5404 -5017
rect 5370 -5051 5404 -5043
rect 5588 -4737 5622 -4729
rect 5588 -4763 5622 -4737
rect 5588 -4805 5622 -4801
rect 5588 -4835 5622 -4805
rect 5588 -4907 5622 -4873
rect 5588 -4975 5622 -4945
rect 5588 -4979 5622 -4975
rect 5588 -5043 5622 -5017
rect 5588 -5051 5622 -5043
rect 5806 -4737 5840 -4729
rect 5806 -4763 5840 -4737
rect 5806 -4805 5840 -4801
rect 5806 -4835 5840 -4805
rect 5806 -4907 5840 -4873
rect 5806 -4975 5840 -4945
rect 5806 -4979 5840 -4975
rect 5806 -5043 5840 -5017
rect 5806 -5051 5840 -5043
rect 24755 -4685 24789 -4679
rect 24755 -4713 24789 -4685
rect 24755 -4753 24789 -4751
rect 24755 -4785 24789 -4753
rect 24755 -4855 24789 -4823
rect 24755 -4857 24789 -4855
rect 24755 -4923 24789 -4895
rect 24755 -4929 24789 -4923
rect 24755 -4991 24789 -4967
rect 24755 -5001 24789 -4991
rect 24755 -5059 24789 -5039
rect 24755 -5073 24789 -5059
rect 411 -5127 445 -5111
rect 411 -5145 445 -5127
rect 3735 -5171 3769 -5137
rect 3953 -5171 3987 -5137
rect 4171 -5171 4205 -5137
rect 4389 -5171 4423 -5137
rect 4607 -5171 4641 -5137
rect 4825 -5171 4859 -5137
rect 5043 -5171 5077 -5137
rect 5261 -5171 5295 -5137
rect 5479 -5171 5513 -5137
rect 5697 -5171 5731 -5137
rect 24755 -5127 24789 -5111
rect 24755 -5145 24789 -5127
rect 411 -5195 445 -5183
rect 411 -5217 445 -5195
rect 411 -5263 445 -5255
rect 411 -5289 445 -5263
rect 411 -5331 445 -5327
rect 411 -5361 445 -5331
rect 411 -5433 445 -5399
rect 411 -5501 445 -5471
rect 411 -5505 445 -5501
rect 411 -5569 445 -5543
rect 411 -5577 445 -5569
rect 24755 -5195 24789 -5183
rect 24755 -5217 24789 -5195
rect 24755 -5263 24789 -5255
rect 24755 -5289 24789 -5263
rect 24755 -5331 24789 -5327
rect 24755 -5361 24789 -5331
rect 24755 -5433 24789 -5399
rect 24755 -5501 24789 -5471
rect 24755 -5505 24789 -5501
rect 3735 -5581 3769 -5547
rect 3953 -5581 3987 -5547
rect 4171 -5581 4205 -5547
rect 4389 -5581 4423 -5547
rect 4607 -5581 4641 -5547
rect 4825 -5581 4859 -5547
rect 5043 -5581 5077 -5547
rect 5261 -5581 5295 -5547
rect 5479 -5581 5513 -5547
rect 5697 -5581 5731 -5547
rect 24755 -5569 24789 -5543
rect 24755 -5577 24789 -5569
rect 411 -5637 445 -5615
rect 411 -5649 445 -5637
rect 411 -5705 445 -5687
rect 411 -5721 445 -5705
rect 411 -5773 445 -5759
rect 411 -5793 445 -5773
rect 411 -5841 445 -5831
rect 411 -5865 445 -5841
rect 411 -5909 445 -5903
rect 411 -5937 445 -5909
rect 411 -5977 445 -5975
rect 411 -6009 445 -5977
rect 3626 -5675 3660 -5667
rect 3626 -5701 3660 -5675
rect 3626 -5743 3660 -5739
rect 3626 -5773 3660 -5743
rect 3626 -5845 3660 -5811
rect 3626 -5913 3660 -5883
rect 3626 -5917 3660 -5913
rect 3626 -5981 3660 -5955
rect 3626 -5989 3660 -5981
rect 3844 -5675 3878 -5667
rect 3844 -5701 3878 -5675
rect 3844 -5743 3878 -5739
rect 3844 -5773 3878 -5743
rect 3844 -5845 3878 -5811
rect 3844 -5913 3878 -5883
rect 3844 -5917 3878 -5913
rect 3844 -5981 3878 -5955
rect 3844 -5989 3878 -5981
rect 4062 -5675 4096 -5667
rect 4062 -5701 4096 -5675
rect 4062 -5743 4096 -5739
rect 4062 -5773 4096 -5743
rect 4062 -5845 4096 -5811
rect 4062 -5913 4096 -5883
rect 4062 -5917 4096 -5913
rect 4062 -5981 4096 -5955
rect 4062 -5989 4096 -5981
rect 4280 -5675 4314 -5667
rect 4280 -5701 4314 -5675
rect 4280 -5743 4314 -5739
rect 4280 -5773 4314 -5743
rect 4280 -5845 4314 -5811
rect 4280 -5913 4314 -5883
rect 4280 -5917 4314 -5913
rect 4280 -5981 4314 -5955
rect 4280 -5989 4314 -5981
rect 4498 -5675 4532 -5667
rect 4498 -5701 4532 -5675
rect 4498 -5743 4532 -5739
rect 4498 -5773 4532 -5743
rect 4498 -5845 4532 -5811
rect 4498 -5913 4532 -5883
rect 4498 -5917 4532 -5913
rect 4498 -5981 4532 -5955
rect 4498 -5989 4532 -5981
rect 4716 -5675 4750 -5667
rect 4716 -5701 4750 -5675
rect 4716 -5743 4750 -5739
rect 4716 -5773 4750 -5743
rect 4716 -5845 4750 -5811
rect 4716 -5913 4750 -5883
rect 4716 -5917 4750 -5913
rect 4716 -5981 4750 -5955
rect 4716 -5989 4750 -5981
rect 4934 -5675 4968 -5667
rect 4934 -5701 4968 -5675
rect 4934 -5743 4968 -5739
rect 4934 -5773 4968 -5743
rect 4934 -5845 4968 -5811
rect 4934 -5913 4968 -5883
rect 4934 -5917 4968 -5913
rect 4934 -5981 4968 -5955
rect 4934 -5989 4968 -5981
rect 5152 -5675 5186 -5667
rect 5152 -5701 5186 -5675
rect 5152 -5743 5186 -5739
rect 5152 -5773 5186 -5743
rect 5152 -5845 5186 -5811
rect 5152 -5913 5186 -5883
rect 5152 -5917 5186 -5913
rect 5152 -5981 5186 -5955
rect 5152 -5989 5186 -5981
rect 5370 -5675 5404 -5667
rect 5370 -5701 5404 -5675
rect 5370 -5743 5404 -5739
rect 5370 -5773 5404 -5743
rect 5370 -5845 5404 -5811
rect 5370 -5913 5404 -5883
rect 5370 -5917 5404 -5913
rect 5370 -5981 5404 -5955
rect 5370 -5989 5404 -5981
rect 5588 -5675 5622 -5667
rect 5588 -5701 5622 -5675
rect 5588 -5743 5622 -5739
rect 5588 -5773 5622 -5743
rect 5588 -5845 5622 -5811
rect 5588 -5913 5622 -5883
rect 5588 -5917 5622 -5913
rect 5588 -5981 5622 -5955
rect 5588 -5989 5622 -5981
rect 5806 -5675 5840 -5667
rect 5806 -5701 5840 -5675
rect 5806 -5743 5840 -5739
rect 5806 -5773 5840 -5743
rect 5806 -5845 5840 -5811
rect 5806 -5913 5840 -5883
rect 5806 -5917 5840 -5913
rect 5806 -5981 5840 -5955
rect 5806 -5989 5840 -5981
rect 24755 -5637 24789 -5615
rect 24755 -5649 24789 -5637
rect 24755 -5705 24789 -5687
rect 24755 -5721 24789 -5705
rect 24755 -5773 24789 -5759
rect 24755 -5793 24789 -5773
rect 24755 -5841 24789 -5831
rect 24755 -5865 24789 -5841
rect 24755 -5909 24789 -5903
rect 24755 -5937 24789 -5909
rect 24755 -5977 24789 -5975
rect 24755 -6009 24789 -5977
rect 411 -6079 445 -6047
rect 411 -6081 445 -6079
rect 3735 -6109 3769 -6075
rect 3953 -6109 3987 -6075
rect 4171 -6109 4205 -6075
rect 4389 -6109 4423 -6075
rect 4607 -6109 4641 -6075
rect 4825 -6109 4859 -6075
rect 5043 -6109 5077 -6075
rect 5261 -6109 5295 -6075
rect 5479 -6109 5513 -6075
rect 5697 -6109 5731 -6075
rect 411 -6147 445 -6119
rect 411 -6153 445 -6147
rect 411 -6215 445 -6191
rect 411 -6225 445 -6215
rect 411 -6283 445 -6263
rect 411 -6297 445 -6283
rect 411 -6351 445 -6335
rect 411 -6369 445 -6351
rect 411 -6419 445 -6407
rect 411 -6441 445 -6419
rect 411 -6487 445 -6479
rect 411 -6513 445 -6487
rect 24755 -6079 24789 -6047
rect 24755 -6081 24789 -6079
rect 24755 -6147 24789 -6119
rect 24755 -6153 24789 -6147
rect 24755 -6215 24789 -6191
rect 24755 -6225 24789 -6215
rect 24755 -6283 24789 -6263
rect 24755 -6297 24789 -6283
rect 24755 -6351 24789 -6335
rect 24755 -6369 24789 -6351
rect 24755 -6419 24789 -6407
rect 24755 -6441 24789 -6419
rect 3735 -6519 3769 -6485
rect 3953 -6519 3987 -6485
rect 4171 -6519 4205 -6485
rect 4389 -6519 4423 -6485
rect 4607 -6519 4641 -6485
rect 4825 -6519 4859 -6485
rect 5043 -6519 5077 -6485
rect 5261 -6519 5295 -6485
rect 5479 -6519 5513 -6485
rect 5697 -6519 5731 -6485
rect 411 -6555 445 -6551
rect 411 -6585 445 -6555
rect 24755 -6487 24789 -6479
rect 24755 -6513 24789 -6487
rect 411 -6657 445 -6623
rect 411 -6725 445 -6695
rect 411 -6729 445 -6725
rect 411 -6793 445 -6767
rect 411 -6801 445 -6793
rect 411 -6861 445 -6839
rect 411 -6873 445 -6861
rect 411 -6929 445 -6911
rect 411 -6945 445 -6929
rect 411 -6997 445 -6983
rect 411 -7017 445 -6997
rect 3626 -6613 3660 -6605
rect 3626 -6639 3660 -6613
rect 3626 -6681 3660 -6677
rect 3626 -6711 3660 -6681
rect 3626 -6783 3660 -6749
rect 3626 -6851 3660 -6821
rect 3626 -6855 3660 -6851
rect 3626 -6919 3660 -6893
rect 3626 -6927 3660 -6919
rect 3844 -6613 3878 -6605
rect 3844 -6639 3878 -6613
rect 3844 -6681 3878 -6677
rect 3844 -6711 3878 -6681
rect 3844 -6783 3878 -6749
rect 3844 -6851 3878 -6821
rect 3844 -6855 3878 -6851
rect 3844 -6919 3878 -6893
rect 3844 -6927 3878 -6919
rect 4062 -6613 4096 -6605
rect 4062 -6639 4096 -6613
rect 4062 -6681 4096 -6677
rect 4062 -6711 4096 -6681
rect 4062 -6783 4096 -6749
rect 4062 -6851 4096 -6821
rect 4062 -6855 4096 -6851
rect 4062 -6919 4096 -6893
rect 4062 -6927 4096 -6919
rect 4280 -6613 4314 -6605
rect 4280 -6639 4314 -6613
rect 4280 -6681 4314 -6677
rect 4280 -6711 4314 -6681
rect 4280 -6783 4314 -6749
rect 4280 -6851 4314 -6821
rect 4280 -6855 4314 -6851
rect 4280 -6919 4314 -6893
rect 4280 -6927 4314 -6919
rect 4498 -6613 4532 -6605
rect 4498 -6639 4532 -6613
rect 4498 -6681 4532 -6677
rect 4498 -6711 4532 -6681
rect 4498 -6783 4532 -6749
rect 4498 -6851 4532 -6821
rect 4498 -6855 4532 -6851
rect 4498 -6919 4532 -6893
rect 4498 -6927 4532 -6919
rect 4716 -6613 4750 -6605
rect 4716 -6639 4750 -6613
rect 4716 -6681 4750 -6677
rect 4716 -6711 4750 -6681
rect 4716 -6783 4750 -6749
rect 4716 -6851 4750 -6821
rect 4716 -6855 4750 -6851
rect 4716 -6919 4750 -6893
rect 4716 -6927 4750 -6919
rect 4934 -6613 4968 -6605
rect 4934 -6639 4968 -6613
rect 4934 -6681 4968 -6677
rect 4934 -6711 4968 -6681
rect 4934 -6783 4968 -6749
rect 4934 -6851 4968 -6821
rect 4934 -6855 4968 -6851
rect 4934 -6919 4968 -6893
rect 4934 -6927 4968 -6919
rect 5152 -6613 5186 -6605
rect 5152 -6639 5186 -6613
rect 5152 -6681 5186 -6677
rect 5152 -6711 5186 -6681
rect 5152 -6783 5186 -6749
rect 5152 -6851 5186 -6821
rect 5152 -6855 5186 -6851
rect 5152 -6919 5186 -6893
rect 5152 -6927 5186 -6919
rect 5370 -6613 5404 -6605
rect 5370 -6639 5404 -6613
rect 5370 -6681 5404 -6677
rect 5370 -6711 5404 -6681
rect 5370 -6783 5404 -6749
rect 5370 -6851 5404 -6821
rect 5370 -6855 5404 -6851
rect 5370 -6919 5404 -6893
rect 5370 -6927 5404 -6919
rect 5588 -6613 5622 -6605
rect 5588 -6639 5622 -6613
rect 5588 -6681 5622 -6677
rect 5588 -6711 5622 -6681
rect 5588 -6783 5622 -6749
rect 5588 -6851 5622 -6821
rect 5588 -6855 5622 -6851
rect 5588 -6919 5622 -6893
rect 5588 -6927 5622 -6919
rect 5806 -6613 5840 -6605
rect 5806 -6639 5840 -6613
rect 5806 -6681 5840 -6677
rect 5806 -6711 5840 -6681
rect 5806 -6783 5840 -6749
rect 5806 -6851 5840 -6821
rect 5806 -6855 5840 -6851
rect 5806 -6919 5840 -6893
rect 5806 -6927 5840 -6919
rect 24755 -6555 24789 -6551
rect 24755 -6585 24789 -6555
rect 24755 -6657 24789 -6623
rect 24755 -6725 24789 -6695
rect 24755 -6729 24789 -6725
rect 24755 -6793 24789 -6767
rect 24755 -6801 24789 -6793
rect 24755 -6861 24789 -6839
rect 24755 -6873 24789 -6861
rect 24755 -6929 24789 -6911
rect 24755 -6945 24789 -6929
rect 411 -7065 445 -7055
rect 411 -7089 445 -7065
rect 3735 -7047 3769 -7013
rect 3953 -7047 3987 -7013
rect 4171 -7047 4205 -7013
rect 4389 -7047 4423 -7013
rect 4607 -7047 4641 -7013
rect 4825 -7047 4859 -7013
rect 5043 -7047 5077 -7013
rect 5261 -7047 5295 -7013
rect 5479 -7047 5513 -7013
rect 5697 -7047 5731 -7013
rect 24755 -6997 24789 -6983
rect 24755 -7017 24789 -6997
rect 411 -7133 445 -7127
rect 411 -7161 445 -7133
rect 411 -7201 445 -7199
rect 411 -7233 445 -7201
rect 411 -7303 445 -7271
rect 411 -7305 445 -7303
rect 411 -7371 445 -7343
rect 411 -7377 445 -7371
rect 411 -7439 445 -7415
rect 411 -7449 445 -7439
rect 24755 -7065 24789 -7055
rect 24755 -7089 24789 -7065
rect 24755 -7133 24789 -7127
rect 24755 -7161 24789 -7133
rect 24755 -7201 24789 -7199
rect 24755 -7233 24789 -7201
rect 24755 -7303 24789 -7271
rect 24755 -7305 24789 -7303
rect 24755 -7371 24789 -7343
rect 24755 -7377 24789 -7371
rect 3735 -7457 3769 -7423
rect 3953 -7457 3987 -7423
rect 4171 -7457 4205 -7423
rect 4389 -7457 4423 -7423
rect 4607 -7457 4641 -7423
rect 4825 -7457 4859 -7423
rect 5043 -7457 5077 -7423
rect 5261 -7457 5295 -7423
rect 5479 -7457 5513 -7423
rect 5697 -7457 5731 -7423
rect 411 -7507 445 -7487
rect 411 -7521 445 -7507
rect 24755 -7439 24789 -7415
rect 24755 -7449 24789 -7439
rect 411 -7575 445 -7559
rect 411 -7593 445 -7575
rect 411 -7643 445 -7631
rect 411 -7665 445 -7643
rect 411 -7711 445 -7703
rect 411 -7737 445 -7711
rect 411 -7779 445 -7775
rect 411 -7809 445 -7779
rect 411 -7881 445 -7847
rect 3626 -7551 3660 -7543
rect 3626 -7577 3660 -7551
rect 3626 -7619 3660 -7615
rect 3626 -7649 3660 -7619
rect 3626 -7721 3660 -7687
rect 3626 -7789 3660 -7759
rect 3626 -7793 3660 -7789
rect 3626 -7857 3660 -7831
rect 3626 -7865 3660 -7857
rect 3844 -7551 3878 -7543
rect 3844 -7577 3878 -7551
rect 3844 -7619 3878 -7615
rect 3844 -7649 3878 -7619
rect 3844 -7721 3878 -7687
rect 3844 -7789 3878 -7759
rect 3844 -7793 3878 -7789
rect 3844 -7857 3878 -7831
rect 3844 -7865 3878 -7857
rect 4062 -7551 4096 -7543
rect 4062 -7577 4096 -7551
rect 4062 -7619 4096 -7615
rect 4062 -7649 4096 -7619
rect 4062 -7721 4096 -7687
rect 4062 -7789 4096 -7759
rect 4062 -7793 4096 -7789
rect 4062 -7857 4096 -7831
rect 4062 -7865 4096 -7857
rect 4280 -7551 4314 -7543
rect 4280 -7577 4314 -7551
rect 4280 -7619 4314 -7615
rect 4280 -7649 4314 -7619
rect 4280 -7721 4314 -7687
rect 4280 -7789 4314 -7759
rect 4280 -7793 4314 -7789
rect 4280 -7857 4314 -7831
rect 4280 -7865 4314 -7857
rect 4498 -7551 4532 -7543
rect 4498 -7577 4532 -7551
rect 4498 -7619 4532 -7615
rect 4498 -7649 4532 -7619
rect 4498 -7721 4532 -7687
rect 4498 -7789 4532 -7759
rect 4498 -7793 4532 -7789
rect 4498 -7857 4532 -7831
rect 4498 -7865 4532 -7857
rect 4716 -7551 4750 -7543
rect 4716 -7577 4750 -7551
rect 4716 -7619 4750 -7615
rect 4716 -7649 4750 -7619
rect 4716 -7721 4750 -7687
rect 4716 -7789 4750 -7759
rect 4716 -7793 4750 -7789
rect 4716 -7857 4750 -7831
rect 4716 -7865 4750 -7857
rect 4934 -7551 4968 -7543
rect 4934 -7577 4968 -7551
rect 4934 -7619 4968 -7615
rect 4934 -7649 4968 -7619
rect 4934 -7721 4968 -7687
rect 4934 -7789 4968 -7759
rect 4934 -7793 4968 -7789
rect 4934 -7857 4968 -7831
rect 4934 -7865 4968 -7857
rect 5152 -7551 5186 -7543
rect 5152 -7577 5186 -7551
rect 5152 -7619 5186 -7615
rect 5152 -7649 5186 -7619
rect 5152 -7721 5186 -7687
rect 5152 -7789 5186 -7759
rect 5152 -7793 5186 -7789
rect 5152 -7857 5186 -7831
rect 5152 -7865 5186 -7857
rect 5370 -7551 5404 -7543
rect 5370 -7577 5404 -7551
rect 5370 -7619 5404 -7615
rect 5370 -7649 5404 -7619
rect 5370 -7721 5404 -7687
rect 5370 -7789 5404 -7759
rect 5370 -7793 5404 -7789
rect 5370 -7857 5404 -7831
rect 5370 -7865 5404 -7857
rect 5588 -7551 5622 -7543
rect 5588 -7577 5622 -7551
rect 5588 -7619 5622 -7615
rect 5588 -7649 5622 -7619
rect 5588 -7721 5622 -7687
rect 5588 -7789 5622 -7759
rect 5588 -7793 5622 -7789
rect 5588 -7857 5622 -7831
rect 5588 -7865 5622 -7857
rect 5806 -7551 5840 -7543
rect 5806 -7577 5840 -7551
rect 5806 -7619 5840 -7615
rect 5806 -7649 5840 -7619
rect 5806 -7721 5840 -7687
rect 5806 -7789 5840 -7759
rect 5806 -7793 5840 -7789
rect 5806 -7857 5840 -7831
rect 5806 -7865 5840 -7857
rect 24755 -7507 24789 -7487
rect 24755 -7521 24789 -7507
rect 24755 -7575 24789 -7559
rect 24755 -7593 24789 -7575
rect 24755 -7643 24789 -7631
rect 24755 -7665 24789 -7643
rect 24755 -7711 24789 -7703
rect 24755 -7737 24789 -7711
rect 24755 -7779 24789 -7775
rect 24755 -7809 24789 -7779
rect 24755 -7881 24789 -7847
rect 411 -7949 445 -7919
rect 411 -7953 445 -7949
rect 411 -8017 445 -7991
rect 411 -8025 445 -8017
rect 3735 -7985 3769 -7951
rect 3953 -7985 3987 -7951
rect 4171 -7985 4205 -7951
rect 4389 -7985 4423 -7951
rect 4607 -7985 4641 -7951
rect 4825 -7985 4859 -7951
rect 5043 -7985 5077 -7951
rect 5261 -7985 5295 -7951
rect 5479 -7985 5513 -7951
rect 5697 -7985 5731 -7951
rect 24755 -7949 24789 -7919
rect 24755 -7953 24789 -7949
rect 411 -8085 445 -8063
rect 411 -8097 445 -8085
rect 411 -8153 445 -8135
rect 411 -8169 445 -8153
rect 411 -8221 445 -8207
rect 411 -8241 445 -8221
rect 24755 -8017 24789 -7991
rect 24755 -8025 24789 -8017
rect 24755 -8085 24789 -8063
rect 24755 -8097 24789 -8085
rect 24755 -8153 24789 -8135
rect 24755 -8169 24789 -8153
rect 24755 -8221 24789 -8207
rect 24755 -8241 24789 -8221
rect 487 -8849 521 -8815
rect 559 -8849 581 -8815
rect 581 -8849 593 -8815
rect 631 -8849 649 -8815
rect 649 -8849 665 -8815
rect 703 -8849 717 -8815
rect 717 -8849 737 -8815
rect 775 -8849 785 -8815
rect 785 -8849 809 -8815
rect 847 -8849 853 -8815
rect 853 -8849 881 -8815
rect 919 -8849 921 -8815
rect 921 -8849 953 -8815
rect 991 -8849 1023 -8815
rect 1023 -8849 1025 -8815
rect 1063 -8849 1091 -8815
rect 1091 -8849 1097 -8815
rect 1135 -8849 1159 -8815
rect 1159 -8849 1169 -8815
rect 1207 -8849 1227 -8815
rect 1227 -8849 1241 -8815
rect 1279 -8849 1295 -8815
rect 1295 -8849 1313 -8815
rect 1351 -8849 1363 -8815
rect 1363 -8849 1385 -8815
rect 1423 -8849 1431 -8815
rect 1431 -8849 1457 -8815
rect 1495 -8849 1499 -8815
rect 1499 -8849 1529 -8815
rect 1567 -8849 1601 -8815
rect 1639 -8849 1669 -8815
rect 1669 -8849 1673 -8815
rect 1711 -8849 1737 -8815
rect 1737 -8849 1745 -8815
rect 1783 -8849 1805 -8815
rect 1805 -8849 1817 -8815
rect 1855 -8849 1873 -8815
rect 1873 -8849 1889 -8815
rect 1927 -8849 1941 -8815
rect 1941 -8849 1961 -8815
rect 1999 -8849 2009 -8815
rect 2009 -8849 2033 -8815
rect 2071 -8849 2077 -8815
rect 2077 -8849 2105 -8815
rect 2143 -8849 2145 -8815
rect 2145 -8849 2177 -8815
rect 2215 -8849 2247 -8815
rect 2247 -8849 2249 -8815
rect 2287 -8849 2315 -8815
rect 2315 -8849 2321 -8815
rect 2359 -8849 2383 -8815
rect 2383 -8849 2393 -8815
rect 2431 -8849 2451 -8815
rect 2451 -8849 2465 -8815
rect 2503 -8849 2519 -8815
rect 2519 -8849 2537 -8815
rect 2575 -8849 2587 -8815
rect 2587 -8849 2609 -8815
rect 2647 -8849 2655 -8815
rect 2655 -8849 2681 -8815
rect 2719 -8849 2723 -8815
rect 2723 -8849 2753 -8815
rect 2791 -8849 2825 -8815
rect 2863 -8849 2893 -8815
rect 2893 -8849 2897 -8815
rect 2935 -8849 2961 -8815
rect 2961 -8849 2969 -8815
rect 3007 -8849 3029 -8815
rect 3029 -8849 3041 -8815
rect 3079 -8849 3097 -8815
rect 3097 -8849 3113 -8815
rect 3151 -8849 3165 -8815
rect 3165 -8849 3185 -8815
rect 3223 -8849 3233 -8815
rect 3233 -8849 3257 -8815
rect 3295 -8849 3301 -8815
rect 3301 -8849 3329 -8815
rect 3367 -8849 3369 -8815
rect 3369 -8849 3401 -8815
rect 3439 -8849 3471 -8815
rect 3471 -8849 3473 -8815
rect 3511 -8849 3539 -8815
rect 3539 -8849 3545 -8815
rect 3583 -8849 3607 -8815
rect 3607 -8849 3617 -8815
rect 3655 -8849 3675 -8815
rect 3675 -8849 3689 -8815
rect 3727 -8849 3743 -8815
rect 3743 -8849 3761 -8815
rect 3799 -8849 3811 -8815
rect 3811 -8849 3833 -8815
rect 3871 -8849 3879 -8815
rect 3879 -8849 3905 -8815
rect 3943 -8849 3947 -8815
rect 3947 -8849 3977 -8815
rect 4015 -8849 4049 -8815
rect 4087 -8849 4117 -8815
rect 4117 -8849 4121 -8815
rect 4159 -8849 4185 -8815
rect 4185 -8849 4193 -8815
rect 4231 -8849 4253 -8815
rect 4253 -8849 4265 -8815
rect 4303 -8849 4321 -8815
rect 4321 -8849 4337 -8815
rect 4375 -8849 4389 -8815
rect 4389 -8849 4409 -8815
rect 4447 -8849 4457 -8815
rect 4457 -8849 4481 -8815
rect 4519 -8849 4525 -8815
rect 4525 -8849 4553 -8815
rect 4591 -8849 4593 -8815
rect 4593 -8849 4625 -8815
rect 4663 -8849 4695 -8815
rect 4695 -8849 4697 -8815
rect 4735 -8849 4763 -8815
rect 4763 -8849 4769 -8815
rect 4807 -8849 4831 -8815
rect 4831 -8849 4841 -8815
rect 4879 -8849 4899 -8815
rect 4899 -8849 4913 -8815
rect 4951 -8849 4967 -8815
rect 4967 -8849 4985 -8815
rect 5023 -8849 5035 -8815
rect 5035 -8849 5057 -8815
rect 5095 -8849 5103 -8815
rect 5103 -8849 5129 -8815
rect 5167 -8849 5171 -8815
rect 5171 -8849 5201 -8815
rect 5239 -8849 5273 -8815
rect 5311 -8849 5341 -8815
rect 5341 -8849 5345 -8815
rect 5383 -8849 5409 -8815
rect 5409 -8849 5417 -8815
rect 5455 -8849 5477 -8815
rect 5477 -8849 5489 -8815
rect 5527 -8849 5545 -8815
rect 5545 -8849 5561 -8815
rect 5599 -8849 5613 -8815
rect 5613 -8849 5633 -8815
rect 5671 -8849 5681 -8815
rect 5681 -8849 5705 -8815
rect 5743 -8849 5749 -8815
rect 5749 -8849 5777 -8815
rect 5815 -8849 5817 -8815
rect 5817 -8849 5849 -8815
rect 5887 -8849 5919 -8815
rect 5919 -8849 5921 -8815
rect 5959 -8849 5987 -8815
rect 5987 -8849 5993 -8815
rect 6031 -8849 6055 -8815
rect 6055 -8849 6065 -8815
rect 6103 -8849 6123 -8815
rect 6123 -8849 6137 -8815
rect 6175 -8849 6191 -8815
rect 6191 -8849 6209 -8815
rect 6247 -8849 6259 -8815
rect 6259 -8849 6281 -8815
rect 6319 -8849 6327 -8815
rect 6327 -8849 6353 -8815
rect 6391 -8849 6395 -8815
rect 6395 -8849 6425 -8815
rect 6463 -8849 6497 -8815
rect 6535 -8849 6565 -8815
rect 6565 -8849 6569 -8815
rect 6607 -8849 6633 -8815
rect 6633 -8849 6641 -8815
rect 6679 -8849 6701 -8815
rect 6701 -8849 6713 -8815
rect 6751 -8849 6769 -8815
rect 6769 -8849 6785 -8815
rect 6823 -8849 6837 -8815
rect 6837 -8849 6857 -8815
rect 6895 -8849 6905 -8815
rect 6905 -8849 6929 -8815
rect 6967 -8849 6973 -8815
rect 6973 -8849 7001 -8815
rect 7039 -8849 7041 -8815
rect 7041 -8849 7073 -8815
rect 7111 -8849 7143 -8815
rect 7143 -8849 7145 -8815
rect 7183 -8849 7211 -8815
rect 7211 -8849 7217 -8815
rect 7255 -8849 7279 -8815
rect 7279 -8849 7289 -8815
rect 7327 -8849 7347 -8815
rect 7347 -8849 7361 -8815
rect 7399 -8849 7415 -8815
rect 7415 -8849 7433 -8815
rect 7471 -8849 7483 -8815
rect 7483 -8849 7505 -8815
rect 7543 -8849 7551 -8815
rect 7551 -8849 7577 -8815
rect 7615 -8849 7619 -8815
rect 7619 -8849 7649 -8815
rect 7687 -8849 7721 -8815
rect 7759 -8849 7789 -8815
rect 7789 -8849 7793 -8815
rect 7831 -8849 7857 -8815
rect 7857 -8849 7865 -8815
rect 7903 -8849 7925 -8815
rect 7925 -8849 7937 -8815
rect 7975 -8849 7993 -8815
rect 7993 -8849 8009 -8815
rect 8047 -8849 8061 -8815
rect 8061 -8849 8081 -8815
rect 8119 -8849 8129 -8815
rect 8129 -8849 8153 -8815
rect 8191 -8849 8197 -8815
rect 8197 -8849 8225 -8815
rect 8263 -8849 8265 -8815
rect 8265 -8849 8297 -8815
rect 8335 -8849 8367 -8815
rect 8367 -8849 8369 -8815
rect 8407 -8849 8435 -8815
rect 8435 -8849 8441 -8815
rect 8479 -8849 8503 -8815
rect 8503 -8849 8513 -8815
rect 8551 -8849 8571 -8815
rect 8571 -8849 8585 -8815
rect 8623 -8849 8639 -8815
rect 8639 -8849 8657 -8815
rect 8695 -8849 8707 -8815
rect 8707 -8849 8729 -8815
rect 8767 -8849 8775 -8815
rect 8775 -8849 8801 -8815
rect 8839 -8849 8843 -8815
rect 8843 -8849 8873 -8815
rect 8911 -8849 8945 -8815
rect 8983 -8849 9013 -8815
rect 9013 -8849 9017 -8815
rect 9055 -8849 9081 -8815
rect 9081 -8849 9089 -8815
rect 9127 -8849 9149 -8815
rect 9149 -8849 9161 -8815
rect 9199 -8849 9217 -8815
rect 9217 -8849 9233 -8815
rect 9271 -8849 9285 -8815
rect 9285 -8849 9305 -8815
rect 9343 -8849 9353 -8815
rect 9353 -8849 9377 -8815
rect 9415 -8849 9421 -8815
rect 9421 -8849 9449 -8815
rect 9487 -8849 9489 -8815
rect 9489 -8849 9521 -8815
rect 9559 -8849 9591 -8815
rect 9591 -8849 9593 -8815
rect 9631 -8849 9659 -8815
rect 9659 -8849 9665 -8815
rect 9703 -8849 9727 -8815
rect 9727 -8849 9737 -8815
rect 9775 -8849 9795 -8815
rect 9795 -8849 9809 -8815
rect 9847 -8849 9863 -8815
rect 9863 -8849 9881 -8815
rect 9919 -8849 9931 -8815
rect 9931 -8849 9953 -8815
rect 9991 -8849 9999 -8815
rect 9999 -8849 10025 -8815
rect 10063 -8849 10067 -8815
rect 10067 -8849 10097 -8815
rect 10135 -8849 10169 -8815
rect 10207 -8849 10237 -8815
rect 10237 -8849 10241 -8815
rect 10279 -8849 10305 -8815
rect 10305 -8849 10313 -8815
rect 10351 -8849 10373 -8815
rect 10373 -8849 10385 -8815
rect 10423 -8849 10441 -8815
rect 10441 -8849 10457 -8815
rect 10495 -8849 10509 -8815
rect 10509 -8849 10529 -8815
rect 10567 -8849 10577 -8815
rect 10577 -8849 10601 -8815
rect 10639 -8849 10645 -8815
rect 10645 -8849 10673 -8815
rect 10711 -8849 10713 -8815
rect 10713 -8849 10745 -8815
rect 10783 -8849 10815 -8815
rect 10815 -8849 10817 -8815
rect 10855 -8849 10883 -8815
rect 10883 -8849 10889 -8815
rect 10927 -8849 10951 -8815
rect 10951 -8849 10961 -8815
rect 10999 -8849 11019 -8815
rect 11019 -8849 11033 -8815
rect 11071 -8849 11087 -8815
rect 11087 -8849 11105 -8815
rect 11143 -8849 11155 -8815
rect 11155 -8849 11177 -8815
rect 11215 -8849 11223 -8815
rect 11223 -8849 11249 -8815
rect 11287 -8849 11291 -8815
rect 11291 -8849 11321 -8815
rect 11359 -8849 11393 -8815
rect 11431 -8849 11461 -8815
rect 11461 -8849 11465 -8815
rect 11503 -8849 11529 -8815
rect 11529 -8849 11537 -8815
rect 11575 -8849 11597 -8815
rect 11597 -8849 11609 -8815
rect 11647 -8849 11665 -8815
rect 11665 -8849 11681 -8815
rect 11719 -8849 11733 -8815
rect 11733 -8849 11753 -8815
rect 11791 -8849 11801 -8815
rect 11801 -8849 11825 -8815
rect 11863 -8849 11869 -8815
rect 11869 -8849 11897 -8815
rect 11935 -8849 11937 -8815
rect 11937 -8849 11969 -8815
rect 12007 -8849 12039 -8815
rect 12039 -8849 12041 -8815
rect 12079 -8849 12107 -8815
rect 12107 -8849 12113 -8815
rect 12151 -8849 12175 -8815
rect 12175 -8849 12185 -8815
rect 12223 -8849 12243 -8815
rect 12243 -8849 12257 -8815
rect 12295 -8849 12311 -8815
rect 12311 -8849 12329 -8815
rect 12367 -8849 12379 -8815
rect 12379 -8849 12401 -8815
rect 12439 -8849 12447 -8815
rect 12447 -8849 12473 -8815
rect 12511 -8849 12515 -8815
rect 12515 -8849 12545 -8815
rect 12583 -8849 12617 -8815
rect 12655 -8849 12685 -8815
rect 12685 -8849 12689 -8815
rect 12727 -8849 12753 -8815
rect 12753 -8849 12761 -8815
rect 12799 -8849 12821 -8815
rect 12821 -8849 12833 -8815
rect 12871 -8849 12889 -8815
rect 12889 -8849 12905 -8815
rect 12943 -8849 12957 -8815
rect 12957 -8849 12977 -8815
rect 13015 -8849 13025 -8815
rect 13025 -8849 13049 -8815
rect 13087 -8849 13093 -8815
rect 13093 -8849 13121 -8815
rect 13159 -8849 13161 -8815
rect 13161 -8849 13193 -8815
rect 13231 -8849 13263 -8815
rect 13263 -8849 13265 -8815
rect 13303 -8849 13331 -8815
rect 13331 -8849 13337 -8815
rect 13375 -8849 13399 -8815
rect 13399 -8849 13409 -8815
rect 13447 -8849 13467 -8815
rect 13467 -8849 13481 -8815
rect 13519 -8849 13535 -8815
rect 13535 -8849 13553 -8815
rect 13591 -8849 13603 -8815
rect 13603 -8849 13625 -8815
rect 13663 -8849 13671 -8815
rect 13671 -8849 13697 -8815
rect 13735 -8849 13739 -8815
rect 13739 -8849 13769 -8815
rect 13807 -8849 13841 -8815
rect 13879 -8849 13909 -8815
rect 13909 -8849 13913 -8815
rect 13951 -8849 13977 -8815
rect 13977 -8849 13985 -8815
rect 14023 -8849 14045 -8815
rect 14045 -8849 14057 -8815
rect 14095 -8849 14113 -8815
rect 14113 -8849 14129 -8815
rect 14167 -8849 14181 -8815
rect 14181 -8849 14201 -8815
rect 14239 -8849 14249 -8815
rect 14249 -8849 14273 -8815
rect 14311 -8849 14317 -8815
rect 14317 -8849 14345 -8815
rect 14383 -8849 14385 -8815
rect 14385 -8849 14417 -8815
rect 14455 -8849 14487 -8815
rect 14487 -8849 14489 -8815
rect 14527 -8849 14555 -8815
rect 14555 -8849 14561 -8815
rect 14599 -8849 14623 -8815
rect 14623 -8849 14633 -8815
rect 14671 -8849 14691 -8815
rect 14691 -8849 14705 -8815
rect 14743 -8849 14759 -8815
rect 14759 -8849 14777 -8815
rect 14815 -8849 14827 -8815
rect 14827 -8849 14849 -8815
rect 14887 -8849 14895 -8815
rect 14895 -8849 14921 -8815
rect 14959 -8849 14963 -8815
rect 14963 -8849 14993 -8815
rect 15031 -8849 15065 -8815
rect 15103 -8849 15133 -8815
rect 15133 -8849 15137 -8815
rect 15175 -8849 15201 -8815
rect 15201 -8849 15209 -8815
rect 15247 -8849 15269 -8815
rect 15269 -8849 15281 -8815
rect 15319 -8849 15337 -8815
rect 15337 -8849 15353 -8815
rect 15391 -8849 15405 -8815
rect 15405 -8849 15425 -8815
rect 15463 -8849 15473 -8815
rect 15473 -8849 15497 -8815
rect 15535 -8849 15541 -8815
rect 15541 -8849 15569 -8815
rect 15607 -8849 15609 -8815
rect 15609 -8849 15641 -8815
rect 15679 -8849 15711 -8815
rect 15711 -8849 15713 -8815
rect 15751 -8849 15779 -8815
rect 15779 -8849 15785 -8815
rect 15823 -8849 15847 -8815
rect 15847 -8849 15857 -8815
rect 15895 -8849 15915 -8815
rect 15915 -8849 15929 -8815
rect 15967 -8849 15983 -8815
rect 15983 -8849 16001 -8815
rect 16039 -8849 16051 -8815
rect 16051 -8849 16073 -8815
rect 16111 -8849 16119 -8815
rect 16119 -8849 16145 -8815
rect 16183 -8849 16187 -8815
rect 16187 -8849 16217 -8815
rect 16255 -8849 16289 -8815
rect 16327 -8849 16357 -8815
rect 16357 -8849 16361 -8815
rect 16399 -8849 16425 -8815
rect 16425 -8849 16433 -8815
rect 16471 -8849 16493 -8815
rect 16493 -8849 16505 -8815
rect 16543 -8849 16561 -8815
rect 16561 -8849 16577 -8815
rect 16615 -8849 16629 -8815
rect 16629 -8849 16649 -8815
rect 16687 -8849 16697 -8815
rect 16697 -8849 16721 -8815
rect 16759 -8849 16765 -8815
rect 16765 -8849 16793 -8815
rect 16831 -8849 16833 -8815
rect 16833 -8849 16865 -8815
rect 16903 -8849 16935 -8815
rect 16935 -8849 16937 -8815
rect 16975 -8849 17003 -8815
rect 17003 -8849 17009 -8815
rect 17047 -8849 17071 -8815
rect 17071 -8849 17081 -8815
rect 17119 -8849 17139 -8815
rect 17139 -8849 17153 -8815
rect 17191 -8849 17207 -8815
rect 17207 -8849 17225 -8815
rect 17263 -8849 17275 -8815
rect 17275 -8849 17297 -8815
rect 17335 -8849 17343 -8815
rect 17343 -8849 17369 -8815
rect 17407 -8849 17411 -8815
rect 17411 -8849 17441 -8815
rect 17479 -8849 17513 -8815
rect 17551 -8849 17581 -8815
rect 17581 -8849 17585 -8815
rect 17623 -8849 17649 -8815
rect 17649 -8849 17657 -8815
rect 17695 -8849 17717 -8815
rect 17717 -8849 17729 -8815
rect 17767 -8849 17785 -8815
rect 17785 -8849 17801 -8815
rect 17839 -8849 17853 -8815
rect 17853 -8849 17873 -8815
rect 17911 -8849 17921 -8815
rect 17921 -8849 17945 -8815
rect 17983 -8849 17989 -8815
rect 17989 -8849 18017 -8815
rect 18055 -8849 18057 -8815
rect 18057 -8849 18089 -8815
rect 18127 -8849 18159 -8815
rect 18159 -8849 18161 -8815
rect 18199 -8849 18227 -8815
rect 18227 -8849 18233 -8815
rect 18271 -8849 18295 -8815
rect 18295 -8849 18305 -8815
rect 18343 -8849 18363 -8815
rect 18363 -8849 18377 -8815
rect 18415 -8849 18431 -8815
rect 18431 -8849 18449 -8815
rect 18487 -8849 18499 -8815
rect 18499 -8849 18521 -8815
rect 18559 -8849 18567 -8815
rect 18567 -8849 18593 -8815
rect 18631 -8849 18635 -8815
rect 18635 -8849 18665 -8815
rect 18703 -8849 18737 -8815
rect 18775 -8849 18805 -8815
rect 18805 -8849 18809 -8815
rect 18847 -8849 18873 -8815
rect 18873 -8849 18881 -8815
rect 18919 -8849 18941 -8815
rect 18941 -8849 18953 -8815
rect 18991 -8849 19009 -8815
rect 19009 -8849 19025 -8815
rect 19063 -8849 19077 -8815
rect 19077 -8849 19097 -8815
rect 19135 -8849 19145 -8815
rect 19145 -8849 19169 -8815
rect 19207 -8849 19213 -8815
rect 19213 -8849 19241 -8815
rect 19279 -8849 19281 -8815
rect 19281 -8849 19313 -8815
rect 19351 -8849 19383 -8815
rect 19383 -8849 19385 -8815
rect 19423 -8849 19451 -8815
rect 19451 -8849 19457 -8815
rect 19495 -8849 19519 -8815
rect 19519 -8849 19529 -8815
rect 19567 -8849 19587 -8815
rect 19587 -8849 19601 -8815
rect 19639 -8849 19655 -8815
rect 19655 -8849 19673 -8815
rect 19711 -8849 19723 -8815
rect 19723 -8849 19745 -8815
rect 19783 -8849 19791 -8815
rect 19791 -8849 19817 -8815
rect 19855 -8849 19859 -8815
rect 19859 -8849 19889 -8815
rect 19927 -8849 19961 -8815
rect 19999 -8849 20029 -8815
rect 20029 -8849 20033 -8815
rect 20071 -8849 20097 -8815
rect 20097 -8849 20105 -8815
rect 20143 -8849 20165 -8815
rect 20165 -8849 20177 -8815
rect 20215 -8849 20233 -8815
rect 20233 -8849 20249 -8815
rect 20287 -8849 20301 -8815
rect 20301 -8849 20321 -8815
rect 20359 -8849 20369 -8815
rect 20369 -8849 20393 -8815
rect 20431 -8849 20437 -8815
rect 20437 -8849 20465 -8815
rect 20503 -8849 20505 -8815
rect 20505 -8849 20537 -8815
rect 20575 -8849 20607 -8815
rect 20607 -8849 20609 -8815
rect 20647 -8849 20675 -8815
rect 20675 -8849 20681 -8815
rect 20719 -8849 20743 -8815
rect 20743 -8849 20753 -8815
rect 20791 -8849 20811 -8815
rect 20811 -8849 20825 -8815
rect 20863 -8849 20879 -8815
rect 20879 -8849 20897 -8815
rect 20935 -8849 20947 -8815
rect 20947 -8849 20969 -8815
rect 21007 -8849 21015 -8815
rect 21015 -8849 21041 -8815
rect 21079 -8849 21083 -8815
rect 21083 -8849 21113 -8815
rect 21151 -8849 21185 -8815
rect 21223 -8849 21253 -8815
rect 21253 -8849 21257 -8815
rect 21295 -8849 21321 -8815
rect 21321 -8849 21329 -8815
rect 21367 -8849 21389 -8815
rect 21389 -8849 21401 -8815
rect 21439 -8849 21457 -8815
rect 21457 -8849 21473 -8815
rect 21511 -8849 21525 -8815
rect 21525 -8849 21545 -8815
rect 21583 -8849 21593 -8815
rect 21593 -8849 21617 -8815
rect 21655 -8849 21661 -8815
rect 21661 -8849 21689 -8815
rect 21727 -8849 21729 -8815
rect 21729 -8849 21761 -8815
rect 21799 -8849 21831 -8815
rect 21831 -8849 21833 -8815
rect 21871 -8849 21899 -8815
rect 21899 -8849 21905 -8815
rect 21943 -8849 21967 -8815
rect 21967 -8849 21977 -8815
rect 22015 -8849 22035 -8815
rect 22035 -8849 22049 -8815
rect 22087 -8849 22103 -8815
rect 22103 -8849 22121 -8815
rect 22159 -8849 22171 -8815
rect 22171 -8849 22193 -8815
rect 22231 -8849 22239 -8815
rect 22239 -8849 22265 -8815
rect 22303 -8849 22307 -8815
rect 22307 -8849 22337 -8815
rect 22375 -8849 22409 -8815
rect 22447 -8849 22477 -8815
rect 22477 -8849 22481 -8815
rect 22519 -8849 22545 -8815
rect 22545 -8849 22553 -8815
rect 22591 -8849 22613 -8815
rect 22613 -8849 22625 -8815
rect 22663 -8849 22681 -8815
rect 22681 -8849 22697 -8815
rect 22735 -8849 22749 -8815
rect 22749 -8849 22769 -8815
rect 22807 -8849 22817 -8815
rect 22817 -8849 22841 -8815
rect 22879 -8849 22885 -8815
rect 22885 -8849 22913 -8815
rect 22951 -8849 22953 -8815
rect 22953 -8849 22985 -8815
rect 23023 -8849 23055 -8815
rect 23055 -8849 23057 -8815
rect 23095 -8849 23123 -8815
rect 23123 -8849 23129 -8815
rect 23167 -8849 23191 -8815
rect 23191 -8849 23201 -8815
rect 23239 -8849 23259 -8815
rect 23259 -8849 23273 -8815
rect 23311 -8849 23327 -8815
rect 23327 -8849 23345 -8815
rect 23383 -8849 23395 -8815
rect 23395 -8849 23417 -8815
rect 23455 -8849 23463 -8815
rect 23463 -8849 23489 -8815
rect 23527 -8849 23531 -8815
rect 23531 -8849 23561 -8815
rect 23599 -8849 23633 -8815
rect 23671 -8849 23701 -8815
rect 23701 -8849 23705 -8815
rect 23743 -8849 23769 -8815
rect 23769 -8849 23777 -8815
rect 23815 -8849 23837 -8815
rect 23837 -8849 23849 -8815
rect 23887 -8849 23905 -8815
rect 23905 -8849 23921 -8815
rect 23959 -8849 23973 -8815
rect 23973 -8849 23993 -8815
rect 24031 -8849 24041 -8815
rect 24041 -8849 24065 -8815
rect 24103 -8849 24109 -8815
rect 24109 -8849 24137 -8815
rect 24175 -8849 24177 -8815
rect 24177 -8849 24209 -8815
rect 24247 -8849 24279 -8815
rect 24279 -8849 24281 -8815
rect 24319 -8849 24347 -8815
rect 24347 -8849 24353 -8815
rect 24391 -8849 24415 -8815
rect 24415 -8849 24425 -8815
rect 24463 -8849 24483 -8815
rect 24483 -8849 24497 -8815
rect 24535 -8849 24551 -8815
rect 24551 -8849 24569 -8815
rect 24607 -8849 24619 -8815
rect 24619 -8849 24641 -8815
rect 24679 -8849 24713 -8815
rect -12221 -11245 -12187 -11211
rect -12149 -11245 -12145 -11211
rect -12145 -11245 -12115 -11211
rect -12077 -11245 -12043 -11211
rect -12005 -11245 -11975 -11211
rect -11975 -11245 -11971 -11211
rect -11933 -11245 -11907 -11211
rect -11907 -11245 -11899 -11211
rect -11861 -11245 -11839 -11211
rect -11839 -11245 -11827 -11211
rect -11789 -11245 -11771 -11211
rect -11771 -11245 -11755 -11211
rect -11717 -11245 -11703 -11211
rect -11703 -11245 -11683 -11211
rect -11645 -11245 -11635 -11211
rect -11635 -11245 -11611 -11211
rect -11573 -11245 -11567 -11211
rect -11567 -11245 -11539 -11211
rect -11501 -11245 -11499 -11211
rect -11499 -11245 -11467 -11211
rect -11429 -11245 -11397 -11211
rect -11397 -11245 -11395 -11211
rect -11357 -11245 -11329 -11211
rect -11329 -11245 -11323 -11211
rect -11285 -11245 -11261 -11211
rect -11261 -11245 -11251 -11211
rect -11213 -11245 -11193 -11211
rect -11193 -11245 -11179 -11211
rect -11141 -11245 -11125 -11211
rect -11125 -11245 -11107 -11211
rect -11069 -11245 -11057 -11211
rect -11057 -11245 -11035 -11211
rect -10997 -11245 -10989 -11211
rect -10989 -11245 -10963 -11211
rect -10925 -11245 -10921 -11211
rect -10921 -11245 -10891 -11211
rect -10853 -11245 -10819 -11211
rect -10781 -11245 -10751 -11211
rect -10751 -11245 -10747 -11211
rect -10709 -11245 -10683 -11211
rect -10683 -11245 -10675 -11211
rect -10637 -11245 -10615 -11211
rect -10615 -11245 -10603 -11211
rect -10565 -11245 -10547 -11211
rect -10547 -11245 -10531 -11211
rect -10493 -11245 -10479 -11211
rect -10479 -11245 -10459 -11211
rect -10421 -11245 -10411 -11211
rect -10411 -11245 -10387 -11211
rect -10349 -11245 -10343 -11211
rect -10343 -11245 -10315 -11211
rect -10277 -11245 -10275 -11211
rect -10275 -11245 -10243 -11211
rect -10205 -11245 -10173 -11211
rect -10173 -11245 -10171 -11211
rect -10133 -11245 -10105 -11211
rect -10105 -11245 -10099 -11211
rect -10061 -11245 -10037 -11211
rect -10037 -11245 -10027 -11211
rect -9989 -11245 -9969 -11211
rect -9969 -11245 -9955 -11211
rect -9917 -11245 -9901 -11211
rect -9901 -11245 -9883 -11211
rect -9845 -11245 -9833 -11211
rect -9833 -11245 -9811 -11211
rect -9773 -11245 -9765 -11211
rect -9765 -11245 -9739 -11211
rect -9701 -11245 -9697 -11211
rect -9697 -11245 -9667 -11211
rect -9629 -11245 -9595 -11211
rect -9557 -11245 -9527 -11211
rect -9527 -11245 -9523 -11211
rect -9485 -11245 -9459 -11211
rect -9459 -11245 -9451 -11211
rect -9413 -11245 -9391 -11211
rect -9391 -11245 -9379 -11211
rect -9341 -11245 -9323 -11211
rect -9323 -11245 -9307 -11211
rect -9269 -11245 -9255 -11211
rect -9255 -11245 -9235 -11211
rect -9197 -11245 -9187 -11211
rect -9187 -11245 -9163 -11211
rect -9125 -11245 -9119 -11211
rect -9119 -11245 -9091 -11211
rect -9053 -11245 -9051 -11211
rect -9051 -11245 -9019 -11211
rect -8981 -11245 -8949 -11211
rect -8949 -11245 -8947 -11211
rect -8909 -11245 -8881 -11211
rect -8881 -11245 -8875 -11211
rect -8837 -11245 -8813 -11211
rect -8813 -11245 -8803 -11211
rect -8765 -11245 -8745 -11211
rect -8745 -11245 -8731 -11211
rect -8693 -11245 -8677 -11211
rect -8677 -11245 -8659 -11211
rect -8621 -11245 -8609 -11211
rect -8609 -11245 -8587 -11211
rect -8549 -11245 -8541 -11211
rect -8541 -11245 -8515 -11211
rect -8477 -11245 -8473 -11211
rect -8473 -11245 -8443 -11211
rect -8405 -11245 -8371 -11211
rect -8333 -11245 -8303 -11211
rect -8303 -11245 -8299 -11211
rect -8261 -11245 -8235 -11211
rect -8235 -11245 -8227 -11211
rect -8189 -11245 -8167 -11211
rect -8167 -11245 -8155 -11211
rect -8117 -11245 -8099 -11211
rect -8099 -11245 -8083 -11211
rect -8045 -11245 -8031 -11211
rect -8031 -11245 -8011 -11211
rect -7973 -11245 -7963 -11211
rect -7963 -11245 -7939 -11211
rect -7901 -11245 -7895 -11211
rect -7895 -11245 -7867 -11211
rect -7829 -11245 -7827 -11211
rect -7827 -11245 -7795 -11211
rect -7757 -11245 -7725 -11211
rect -7725 -11245 -7723 -11211
rect -7685 -11245 -7657 -11211
rect -7657 -11245 -7651 -11211
rect -7613 -11245 -7589 -11211
rect -7589 -11245 -7579 -11211
rect -7541 -11245 -7521 -11211
rect -7521 -11245 -7507 -11211
rect -7469 -11245 -7453 -11211
rect -7453 -11245 -7435 -11211
rect -7397 -11245 -7385 -11211
rect -7385 -11245 -7363 -11211
rect -7325 -11245 -7317 -11211
rect -7317 -11245 -7291 -11211
rect -7253 -11245 -7249 -11211
rect -7249 -11245 -7219 -11211
rect -7181 -11245 -7147 -11211
rect -7109 -11245 -7079 -11211
rect -7079 -11245 -7075 -11211
rect -7037 -11245 -7011 -11211
rect -7011 -11245 -7003 -11211
rect -6965 -11245 -6943 -11211
rect -6943 -11245 -6931 -11211
rect -6893 -11245 -6875 -11211
rect -6875 -11245 -6859 -11211
rect -6821 -11245 -6807 -11211
rect -6807 -11245 -6787 -11211
rect -6749 -11245 -6739 -11211
rect -6739 -11245 -6715 -11211
rect -6677 -11245 -6671 -11211
rect -6671 -11245 -6643 -11211
rect -6605 -11245 -6603 -11211
rect -6603 -11245 -6571 -11211
rect -6533 -11245 -6501 -11211
rect -6501 -11245 -6499 -11211
rect -6461 -11245 -6433 -11211
rect -6433 -11245 -6427 -11211
rect -6389 -11245 -6365 -11211
rect -6365 -11245 -6355 -11211
rect -6317 -11245 -6297 -11211
rect -6297 -11245 -6283 -11211
rect -6245 -11245 -6229 -11211
rect -6229 -11245 -6211 -11211
rect -6173 -11245 -6161 -11211
rect -6161 -11245 -6139 -11211
rect -6101 -11245 -6093 -11211
rect -6093 -11245 -6067 -11211
rect -6029 -11245 -6025 -11211
rect -6025 -11245 -5995 -11211
rect -5957 -11245 -5923 -11211
rect -5885 -11245 -5855 -11211
rect -5855 -11245 -5851 -11211
rect -5813 -11245 -5787 -11211
rect -5787 -11245 -5779 -11211
rect -5741 -11245 -5719 -11211
rect -5719 -11245 -5707 -11211
rect -5669 -11245 -5651 -11211
rect -5651 -11245 -5635 -11211
rect -5597 -11245 -5583 -11211
rect -5583 -11245 -5563 -11211
rect -5525 -11245 -5515 -11211
rect -5515 -11245 -5491 -11211
rect -5453 -11245 -5447 -11211
rect -5447 -11245 -5419 -11211
rect -5381 -11245 -5379 -11211
rect -5379 -11245 -5347 -11211
rect -5309 -11245 -5277 -11211
rect -5277 -11245 -5275 -11211
rect -5237 -11245 -5209 -11211
rect -5209 -11245 -5203 -11211
rect -5165 -11245 -5141 -11211
rect -5141 -11245 -5131 -11211
rect -5093 -11245 -5073 -11211
rect -5073 -11245 -5059 -11211
rect -5021 -11245 -5005 -11211
rect -5005 -11245 -4987 -11211
rect -4949 -11245 -4937 -11211
rect -4937 -11245 -4915 -11211
rect -4877 -11245 -4869 -11211
rect -4869 -11245 -4843 -11211
rect -4805 -11245 -4801 -11211
rect -4801 -11245 -4771 -11211
rect -4733 -11245 -4699 -11211
rect -4661 -11245 -4631 -11211
rect -4631 -11245 -4627 -11211
rect -4589 -11245 -4563 -11211
rect -4563 -11245 -4555 -11211
rect -4517 -11245 -4495 -11211
rect -4495 -11245 -4483 -11211
rect -4445 -11245 -4427 -11211
rect -4427 -11245 -4411 -11211
rect -4373 -11245 -4359 -11211
rect -4359 -11245 -4339 -11211
rect -4301 -11245 -4291 -11211
rect -4291 -11245 -4267 -11211
rect -4229 -11245 -4223 -11211
rect -4223 -11245 -4195 -11211
rect -4157 -11245 -4155 -11211
rect -4155 -11245 -4123 -11211
rect -4085 -11245 -4053 -11211
rect -4053 -11245 -4051 -11211
rect -4013 -11245 -3985 -11211
rect -3985 -11245 -3979 -11211
rect -3941 -11245 -3917 -11211
rect -3917 -11245 -3907 -11211
rect -3869 -11245 -3849 -11211
rect -3849 -11245 -3835 -11211
rect -3797 -11245 -3781 -11211
rect -3781 -11245 -3763 -11211
rect -3725 -11245 -3713 -11211
rect -3713 -11245 -3691 -11211
rect -3653 -11245 -3645 -11211
rect -3645 -11245 -3619 -11211
rect -3581 -11245 -3577 -11211
rect -3577 -11245 -3547 -11211
rect -3509 -11245 -3475 -11211
rect -3437 -11245 -3407 -11211
rect -3407 -11245 -3403 -11211
rect -3365 -11245 -3339 -11211
rect -3339 -11245 -3331 -11211
rect -3293 -11245 -3271 -11211
rect -3271 -11245 -3259 -11211
rect -3221 -11245 -3203 -11211
rect -3203 -11245 -3187 -11211
rect -3149 -11245 -3135 -11211
rect -3135 -11245 -3115 -11211
rect -3077 -11245 -3067 -11211
rect -3067 -11245 -3043 -11211
rect -3005 -11245 -2999 -11211
rect -2999 -11245 -2971 -11211
rect -2933 -11245 -2931 -11211
rect -2931 -11245 -2899 -11211
rect -2861 -11245 -2829 -11211
rect -2829 -11245 -2827 -11211
rect -2789 -11245 -2761 -11211
rect -2761 -11245 -2755 -11211
rect -2717 -11245 -2693 -11211
rect -2693 -11245 -2683 -11211
rect -2645 -11245 -2625 -11211
rect -2625 -11245 -2611 -11211
rect -2573 -11245 -2557 -11211
rect -2557 -11245 -2539 -11211
rect -2501 -11245 -2489 -11211
rect -2489 -11245 -2467 -11211
rect -2429 -11245 -2421 -11211
rect -2421 -11245 -2395 -11211
rect -2357 -11245 -2353 -11211
rect -2353 -11245 -2323 -11211
rect -2285 -11245 -2251 -11211
rect -2213 -11245 -2183 -11211
rect -2183 -11245 -2179 -11211
rect -2141 -11245 -2115 -11211
rect -2115 -11245 -2107 -11211
rect -2069 -11245 -2047 -11211
rect -2047 -11245 -2035 -11211
rect -1997 -11245 -1979 -11211
rect -1979 -11245 -1963 -11211
rect -1925 -11245 -1911 -11211
rect -1911 -11245 -1891 -11211
rect -1853 -11245 -1843 -11211
rect -1843 -11245 -1819 -11211
rect -1781 -11245 -1775 -11211
rect -1775 -11245 -1747 -11211
rect -1709 -11245 -1707 -11211
rect -1707 -11245 -1675 -11211
rect -1637 -11245 -1605 -11211
rect -1605 -11245 -1603 -11211
rect -1565 -11245 -1537 -11211
rect -1537 -11245 -1531 -11211
rect -1493 -11245 -1469 -11211
rect -1469 -11245 -1459 -11211
rect -1421 -11245 -1401 -11211
rect -1401 -11245 -1387 -11211
rect -1349 -11245 -1333 -11211
rect -1333 -11245 -1315 -11211
rect -1277 -11245 -1265 -11211
rect -1265 -11245 -1243 -11211
rect -1205 -11245 -1197 -11211
rect -1197 -11245 -1171 -11211
rect -1133 -11245 -1129 -11211
rect -1129 -11245 -1099 -11211
rect -1061 -11245 -1027 -11211
rect -989 -11245 -959 -11211
rect -959 -11245 -955 -11211
rect -917 -11245 -891 -11211
rect -891 -11245 -883 -11211
rect -845 -11245 -823 -11211
rect -823 -11245 -811 -11211
rect -773 -11245 -755 -11211
rect -755 -11245 -739 -11211
rect -701 -11245 -687 -11211
rect -687 -11245 -667 -11211
rect -629 -11245 -619 -11211
rect -619 -11245 -595 -11211
rect -557 -11245 -551 -11211
rect -551 -11245 -523 -11211
rect -485 -11245 -483 -11211
rect -483 -11245 -451 -11211
rect -413 -11245 -381 -11211
rect -381 -11245 -379 -11211
rect -341 -11245 -313 -11211
rect -313 -11245 -307 -11211
rect -269 -11245 -245 -11211
rect -245 -11245 -235 -11211
rect -197 -11245 -177 -11211
rect -177 -11245 -163 -11211
rect -125 -11245 -109 -11211
rect -109 -11245 -91 -11211
rect -53 -11245 -41 -11211
rect -41 -11245 -19 -11211
rect 19 -11245 27 -11211
rect 27 -11245 53 -11211
rect 91 -11245 95 -11211
rect 95 -11245 125 -11211
rect 163 -11245 197 -11211
rect 235 -11245 265 -11211
rect 265 -11245 269 -11211
rect 307 -11245 333 -11211
rect 333 -11245 341 -11211
rect 379 -11245 401 -11211
rect 401 -11245 413 -11211
rect 451 -11245 469 -11211
rect 469 -11245 485 -11211
rect 523 -11245 537 -11211
rect 537 -11245 557 -11211
rect 595 -11245 605 -11211
rect 605 -11245 629 -11211
rect 667 -11245 673 -11211
rect 673 -11245 701 -11211
rect 739 -11245 741 -11211
rect 741 -11245 773 -11211
rect 811 -11245 843 -11211
rect 843 -11245 845 -11211
rect 883 -11245 911 -11211
rect 911 -11245 917 -11211
rect 955 -11245 979 -11211
rect 979 -11245 989 -11211
rect 1027 -11245 1047 -11211
rect 1047 -11245 1061 -11211
rect 1099 -11245 1115 -11211
rect 1115 -11245 1133 -11211
rect 1171 -11245 1183 -11211
rect 1183 -11245 1205 -11211
rect 1243 -11245 1251 -11211
rect 1251 -11245 1277 -11211
rect 1315 -11245 1319 -11211
rect 1319 -11245 1349 -11211
rect 1387 -11245 1421 -11211
rect 1459 -11245 1489 -11211
rect 1489 -11245 1493 -11211
rect 1531 -11245 1557 -11211
rect 1557 -11245 1565 -11211
rect 1603 -11245 1625 -11211
rect 1625 -11245 1637 -11211
rect 1675 -11245 1693 -11211
rect 1693 -11245 1709 -11211
rect 1747 -11245 1761 -11211
rect 1761 -11245 1781 -11211
rect 1819 -11245 1829 -11211
rect 1829 -11245 1853 -11211
rect 1891 -11245 1897 -11211
rect 1897 -11245 1925 -11211
rect 1963 -11245 1965 -11211
rect 1965 -11245 1997 -11211
rect 2035 -11245 2067 -11211
rect 2067 -11245 2069 -11211
rect 2107 -11245 2135 -11211
rect 2135 -11245 2141 -11211
rect 2179 -11245 2203 -11211
rect 2203 -11245 2213 -11211
rect 2251 -11245 2271 -11211
rect 2271 -11245 2285 -11211
rect 2323 -11245 2339 -11211
rect 2339 -11245 2357 -11211
rect 2395 -11245 2407 -11211
rect 2407 -11245 2429 -11211
rect 2467 -11245 2475 -11211
rect 2475 -11245 2501 -11211
rect 2539 -11245 2543 -11211
rect 2543 -11245 2573 -11211
rect 2611 -11245 2645 -11211
rect 2683 -11245 2713 -11211
rect 2713 -11245 2717 -11211
rect 2755 -11245 2781 -11211
rect 2781 -11245 2789 -11211
rect 2827 -11245 2849 -11211
rect 2849 -11245 2861 -11211
rect 2899 -11245 2917 -11211
rect 2917 -11245 2933 -11211
rect 2971 -11245 2985 -11211
rect 2985 -11245 3005 -11211
rect 3043 -11245 3053 -11211
rect 3053 -11245 3077 -11211
rect 3115 -11245 3121 -11211
rect 3121 -11245 3149 -11211
rect 3187 -11245 3189 -11211
rect 3189 -11245 3221 -11211
rect 3259 -11245 3291 -11211
rect 3291 -11245 3293 -11211
rect 3331 -11245 3359 -11211
rect 3359 -11245 3365 -11211
rect 3403 -11245 3427 -11211
rect 3427 -11245 3437 -11211
rect 3475 -11245 3495 -11211
rect 3495 -11245 3509 -11211
rect 3547 -11245 3563 -11211
rect 3563 -11245 3581 -11211
rect 3619 -11245 3631 -11211
rect 3631 -11245 3653 -11211
rect 3691 -11245 3699 -11211
rect 3699 -11245 3725 -11211
rect 3763 -11245 3767 -11211
rect 3767 -11245 3797 -11211
rect 3835 -11245 3869 -11211
rect 3907 -11245 3937 -11211
rect 3937 -11245 3941 -11211
rect 3979 -11245 4005 -11211
rect 4005 -11245 4013 -11211
rect 4051 -11245 4073 -11211
rect 4073 -11245 4085 -11211
rect 4123 -11245 4141 -11211
rect 4141 -11245 4157 -11211
rect 4195 -11245 4209 -11211
rect 4209 -11245 4229 -11211
rect 4267 -11245 4277 -11211
rect 4277 -11245 4301 -11211
rect 4339 -11245 4345 -11211
rect 4345 -11245 4373 -11211
rect 4411 -11245 4413 -11211
rect 4413 -11245 4445 -11211
rect 4483 -11245 4515 -11211
rect 4515 -11245 4517 -11211
rect 4555 -11245 4583 -11211
rect 4583 -11245 4589 -11211
rect 4627 -11245 4651 -11211
rect 4651 -11245 4661 -11211
rect 4699 -11245 4719 -11211
rect 4719 -11245 4733 -11211
rect 4771 -11245 4787 -11211
rect 4787 -11245 4805 -11211
rect 4843 -11245 4855 -11211
rect 4855 -11245 4877 -11211
rect 4915 -11245 4923 -11211
rect 4923 -11245 4949 -11211
rect 4987 -11245 4991 -11211
rect 4991 -11245 5021 -11211
rect 5059 -11245 5093 -11211
rect 5131 -11245 5161 -11211
rect 5161 -11245 5165 -11211
rect 5203 -11245 5229 -11211
rect 5229 -11245 5237 -11211
rect 5275 -11245 5297 -11211
rect 5297 -11245 5309 -11211
rect 5347 -11245 5365 -11211
rect 5365 -11245 5381 -11211
rect 5419 -11245 5433 -11211
rect 5433 -11245 5453 -11211
rect 5491 -11245 5501 -11211
rect 5501 -11245 5525 -11211
rect 5563 -11245 5569 -11211
rect 5569 -11245 5597 -11211
rect 5635 -11245 5637 -11211
rect 5637 -11245 5669 -11211
rect 5707 -11245 5739 -11211
rect 5739 -11245 5741 -11211
rect 5779 -11245 5807 -11211
rect 5807 -11245 5813 -11211
rect 5851 -11245 5875 -11211
rect 5875 -11245 5885 -11211
rect 5923 -11245 5943 -11211
rect 5943 -11245 5957 -11211
rect 5995 -11245 6011 -11211
rect 6011 -11245 6029 -11211
rect 6067 -11245 6079 -11211
rect 6079 -11245 6101 -11211
rect 6139 -11245 6147 -11211
rect 6147 -11245 6173 -11211
rect 6211 -11245 6215 -11211
rect 6215 -11245 6245 -11211
rect 6283 -11245 6317 -11211
rect 6355 -11245 6385 -11211
rect 6385 -11245 6389 -11211
rect 6427 -11245 6453 -11211
rect 6453 -11245 6461 -11211
rect 6499 -11245 6521 -11211
rect 6521 -11245 6533 -11211
rect 6571 -11245 6589 -11211
rect 6589 -11245 6605 -11211
rect 6643 -11245 6657 -11211
rect 6657 -11245 6677 -11211
rect 6715 -11245 6725 -11211
rect 6725 -11245 6749 -11211
rect 6787 -11245 6793 -11211
rect 6793 -11245 6821 -11211
rect 6859 -11245 6861 -11211
rect 6861 -11245 6893 -11211
rect 6931 -11245 6963 -11211
rect 6963 -11245 6965 -11211
rect 7003 -11245 7031 -11211
rect 7031 -11245 7037 -11211
rect 7075 -11245 7099 -11211
rect 7099 -11245 7109 -11211
rect 7147 -11245 7167 -11211
rect 7167 -11245 7181 -11211
rect 7219 -11245 7235 -11211
rect 7235 -11245 7253 -11211
rect 7291 -11245 7303 -11211
rect 7303 -11245 7325 -11211
rect 7363 -11245 7371 -11211
rect 7371 -11245 7397 -11211
rect 7435 -11245 7439 -11211
rect 7439 -11245 7469 -11211
rect 7507 -11245 7541 -11211
rect 7579 -11245 7609 -11211
rect 7609 -11245 7613 -11211
rect 7651 -11245 7677 -11211
rect 7677 -11245 7685 -11211
rect 7723 -11245 7745 -11211
rect 7745 -11245 7757 -11211
rect 7795 -11245 7813 -11211
rect 7813 -11245 7829 -11211
rect 7867 -11245 7881 -11211
rect 7881 -11245 7901 -11211
rect 7939 -11245 7949 -11211
rect 7949 -11245 7973 -11211
rect 8011 -11245 8017 -11211
rect 8017 -11245 8045 -11211
rect 8083 -11245 8085 -11211
rect 8085 -11245 8117 -11211
rect 8155 -11245 8187 -11211
rect 8187 -11245 8189 -11211
rect 8227 -11245 8255 -11211
rect 8255 -11245 8261 -11211
rect 8299 -11245 8323 -11211
rect 8323 -11245 8333 -11211
rect 8371 -11245 8391 -11211
rect 8391 -11245 8405 -11211
rect 8443 -11245 8459 -11211
rect 8459 -11245 8477 -11211
rect 8515 -11245 8527 -11211
rect 8527 -11245 8549 -11211
rect 8587 -11245 8595 -11211
rect 8595 -11245 8621 -11211
rect 8659 -11245 8663 -11211
rect 8663 -11245 8693 -11211
rect 8731 -11245 8765 -11211
rect 8803 -11245 8833 -11211
rect 8833 -11245 8837 -11211
rect 8875 -11245 8901 -11211
rect 8901 -11245 8909 -11211
rect 8947 -11245 8969 -11211
rect 8969 -11245 8981 -11211
rect 9019 -11245 9037 -11211
rect 9037 -11245 9053 -11211
rect 9091 -11245 9105 -11211
rect 9105 -11245 9125 -11211
rect 9163 -11245 9173 -11211
rect 9173 -11245 9197 -11211
rect 9235 -11245 9241 -11211
rect 9241 -11245 9269 -11211
rect 9307 -11245 9309 -11211
rect 9309 -11245 9341 -11211
rect 9379 -11245 9411 -11211
rect 9411 -11245 9413 -11211
rect 9451 -11245 9479 -11211
rect 9479 -11245 9485 -11211
rect 9523 -11245 9547 -11211
rect 9547 -11245 9557 -11211
rect 9595 -11245 9615 -11211
rect 9615 -11245 9629 -11211
rect 9667 -11245 9683 -11211
rect 9683 -11245 9701 -11211
rect 9739 -11245 9751 -11211
rect 9751 -11245 9773 -11211
rect 9811 -11245 9819 -11211
rect 9819 -11245 9845 -11211
rect 9883 -11245 9887 -11211
rect 9887 -11245 9917 -11211
rect 9955 -11245 9989 -11211
rect 10027 -11245 10057 -11211
rect 10057 -11245 10061 -11211
rect 10099 -11245 10125 -11211
rect 10125 -11245 10133 -11211
rect 10171 -11245 10193 -11211
rect 10193 -11245 10205 -11211
rect 10243 -11245 10261 -11211
rect 10261 -11245 10277 -11211
rect 10315 -11245 10329 -11211
rect 10329 -11245 10349 -11211
rect 10387 -11245 10397 -11211
rect 10397 -11245 10421 -11211
rect 10459 -11245 10465 -11211
rect 10465 -11245 10493 -11211
rect 10531 -11245 10533 -11211
rect 10533 -11245 10565 -11211
rect 10603 -11245 10635 -11211
rect 10635 -11245 10637 -11211
rect 10675 -11245 10703 -11211
rect 10703 -11245 10709 -11211
rect 10747 -11245 10771 -11211
rect 10771 -11245 10781 -11211
rect 10819 -11245 10839 -11211
rect 10839 -11245 10853 -11211
rect 10891 -11245 10907 -11211
rect 10907 -11245 10925 -11211
rect 10963 -11245 10975 -11211
rect 10975 -11245 10997 -11211
rect 11035 -11245 11043 -11211
rect 11043 -11245 11069 -11211
rect 11107 -11245 11111 -11211
rect 11111 -11245 11141 -11211
rect 11179 -11245 11213 -11211
rect 11251 -11245 11281 -11211
rect 11281 -11245 11285 -11211
rect 11323 -11245 11349 -11211
rect 11349 -11245 11357 -11211
rect 11395 -11245 11417 -11211
rect 11417 -11245 11429 -11211
rect 11467 -11245 11485 -11211
rect 11485 -11245 11501 -11211
rect 11539 -11245 11553 -11211
rect 11553 -11245 11573 -11211
rect 11611 -11245 11621 -11211
rect 11621 -11245 11645 -11211
rect 11683 -11245 11689 -11211
rect 11689 -11245 11717 -11211
rect 11755 -11245 11757 -11211
rect 11757 -11245 11789 -11211
rect 11827 -11245 11859 -11211
rect 11859 -11245 11861 -11211
rect 11899 -11245 11927 -11211
rect 11927 -11245 11933 -11211
rect 11971 -11245 11995 -11211
rect 11995 -11245 12005 -11211
rect 12043 -11245 12063 -11211
rect 12063 -11245 12077 -11211
rect 12115 -11245 12131 -11211
rect 12131 -11245 12149 -11211
rect 12187 -11245 12199 -11211
rect 12199 -11245 12221 -11211
rect 12259 -11245 12267 -11211
rect 12267 -11245 12293 -11211
rect 12331 -11245 12335 -11211
rect 12335 -11245 12365 -11211
rect 12403 -11245 12437 -11211
rect 12475 -11245 12505 -11211
rect 12505 -11245 12509 -11211
rect 12547 -11245 12573 -11211
rect 12573 -11245 12581 -11211
rect 12619 -11245 12641 -11211
rect 12641 -11245 12653 -11211
rect 12691 -11245 12709 -11211
rect 12709 -11245 12725 -11211
rect 12763 -11245 12777 -11211
rect 12777 -11245 12797 -11211
rect 12835 -11245 12845 -11211
rect 12845 -11245 12869 -11211
rect 12907 -11245 12913 -11211
rect 12913 -11245 12941 -11211
rect 12979 -11245 12981 -11211
rect 12981 -11245 13013 -11211
rect 13051 -11245 13083 -11211
rect 13083 -11245 13085 -11211
rect 13123 -11245 13151 -11211
rect 13151 -11245 13157 -11211
rect 13195 -11245 13219 -11211
rect 13219 -11245 13229 -11211
rect 13267 -11245 13287 -11211
rect 13287 -11245 13301 -11211
rect 13339 -11245 13355 -11211
rect 13355 -11245 13373 -11211
rect 13411 -11245 13423 -11211
rect 13423 -11245 13445 -11211
rect 13483 -11245 13491 -11211
rect 13491 -11245 13517 -11211
rect 13555 -11245 13559 -11211
rect 13559 -11245 13589 -11211
rect 13627 -11245 13661 -11211
rect 13699 -11245 13729 -11211
rect 13729 -11245 13733 -11211
rect 13771 -11245 13797 -11211
rect 13797 -11245 13805 -11211
rect 13843 -11245 13865 -11211
rect 13865 -11245 13877 -11211
rect 13915 -11245 13933 -11211
rect 13933 -11245 13949 -11211
rect 13987 -11245 14001 -11211
rect 14001 -11245 14021 -11211
rect 14059 -11245 14069 -11211
rect 14069 -11245 14093 -11211
rect 14131 -11245 14137 -11211
rect 14137 -11245 14165 -11211
rect 14203 -11245 14205 -11211
rect 14205 -11245 14237 -11211
rect 14275 -11245 14307 -11211
rect 14307 -11245 14309 -11211
rect 14347 -11245 14375 -11211
rect 14375 -11245 14381 -11211
rect 14419 -11245 14443 -11211
rect 14443 -11245 14453 -11211
rect 14491 -11245 14511 -11211
rect 14511 -11245 14525 -11211
rect 14563 -11245 14579 -11211
rect 14579 -11245 14597 -11211
rect 14635 -11245 14647 -11211
rect 14647 -11245 14669 -11211
rect 14707 -11245 14715 -11211
rect 14715 -11245 14741 -11211
rect 14779 -11245 14783 -11211
rect 14783 -11245 14813 -11211
rect 14851 -11245 14885 -11211
rect 14923 -11245 14953 -11211
rect 14953 -11245 14957 -11211
rect 14995 -11245 15021 -11211
rect 15021 -11245 15029 -11211
rect 15067 -11245 15089 -11211
rect 15089 -11245 15101 -11211
rect 15139 -11245 15157 -11211
rect 15157 -11245 15173 -11211
rect 15211 -11245 15225 -11211
rect 15225 -11245 15245 -11211
rect 15283 -11245 15293 -11211
rect 15293 -11245 15317 -11211
rect 15355 -11245 15361 -11211
rect 15361 -11245 15389 -11211
rect 15427 -11245 15429 -11211
rect 15429 -11245 15461 -11211
rect 15499 -11245 15531 -11211
rect 15531 -11245 15533 -11211
rect 15571 -11245 15599 -11211
rect 15599 -11245 15605 -11211
rect 15643 -11245 15667 -11211
rect 15667 -11245 15677 -11211
rect 15715 -11245 15735 -11211
rect 15735 -11245 15749 -11211
rect 15787 -11245 15803 -11211
rect 15803 -11245 15821 -11211
rect 15859 -11245 15871 -11211
rect 15871 -11245 15893 -11211
rect 15931 -11245 15939 -11211
rect 15939 -11245 15965 -11211
rect 16003 -11245 16007 -11211
rect 16007 -11245 16037 -11211
rect 16075 -11245 16109 -11211
rect 16147 -11245 16177 -11211
rect 16177 -11245 16181 -11211
rect 16219 -11245 16245 -11211
rect 16245 -11245 16253 -11211
rect 16291 -11245 16313 -11211
rect 16313 -11245 16325 -11211
rect 16363 -11245 16381 -11211
rect 16381 -11245 16397 -11211
rect 16435 -11245 16449 -11211
rect 16449 -11245 16469 -11211
rect 16507 -11245 16517 -11211
rect 16517 -11245 16541 -11211
rect 16579 -11245 16585 -11211
rect 16585 -11245 16613 -11211
rect 16651 -11245 16653 -11211
rect 16653 -11245 16685 -11211
rect 16723 -11245 16755 -11211
rect 16755 -11245 16757 -11211
rect 16795 -11245 16823 -11211
rect 16823 -11245 16829 -11211
rect 16867 -11245 16891 -11211
rect 16891 -11245 16901 -11211
rect 16939 -11245 16959 -11211
rect 16959 -11245 16973 -11211
rect 17011 -11245 17027 -11211
rect 17027 -11245 17045 -11211
rect 17083 -11245 17095 -11211
rect 17095 -11245 17117 -11211
rect 17155 -11245 17163 -11211
rect 17163 -11245 17189 -11211
rect 17227 -11245 17231 -11211
rect 17231 -11245 17261 -11211
rect 17299 -11245 17333 -11211
rect 17371 -11245 17401 -11211
rect 17401 -11245 17405 -11211
rect 17443 -11245 17469 -11211
rect 17469 -11245 17477 -11211
rect 17515 -11245 17537 -11211
rect 17537 -11245 17549 -11211
rect 17587 -11245 17605 -11211
rect 17605 -11245 17621 -11211
rect 17659 -11245 17673 -11211
rect 17673 -11245 17693 -11211
rect 17731 -11245 17741 -11211
rect 17741 -11245 17765 -11211
rect 17803 -11245 17809 -11211
rect 17809 -11245 17837 -11211
rect 17875 -11245 17877 -11211
rect 17877 -11245 17909 -11211
rect 17947 -11245 17979 -11211
rect 17979 -11245 17981 -11211
rect 18019 -11245 18047 -11211
rect 18047 -11245 18053 -11211
rect 18091 -11245 18115 -11211
rect 18115 -11245 18125 -11211
rect 18163 -11245 18183 -11211
rect 18183 -11245 18197 -11211
rect 18235 -11245 18251 -11211
rect 18251 -11245 18269 -11211
rect 18307 -11245 18319 -11211
rect 18319 -11245 18341 -11211
rect 18379 -11245 18387 -11211
rect 18387 -11245 18413 -11211
rect 18451 -11245 18455 -11211
rect 18455 -11245 18485 -11211
rect 18523 -11245 18557 -11211
rect 18595 -11245 18625 -11211
rect 18625 -11245 18629 -11211
rect 18667 -11245 18693 -11211
rect 18693 -11245 18701 -11211
rect 18739 -11245 18761 -11211
rect 18761 -11245 18773 -11211
rect 18811 -11245 18829 -11211
rect 18829 -11245 18845 -11211
rect 18883 -11245 18897 -11211
rect 18897 -11245 18917 -11211
rect 18955 -11245 18965 -11211
rect 18965 -11245 18989 -11211
rect 19027 -11245 19033 -11211
rect 19033 -11245 19061 -11211
rect 19099 -11245 19101 -11211
rect 19101 -11245 19133 -11211
rect 19171 -11245 19203 -11211
rect 19203 -11245 19205 -11211
rect 19243 -11245 19271 -11211
rect 19271 -11245 19277 -11211
rect 19315 -11245 19339 -11211
rect 19339 -11245 19349 -11211
rect 19387 -11245 19407 -11211
rect 19407 -11245 19421 -11211
rect 19459 -11245 19475 -11211
rect 19475 -11245 19493 -11211
rect 19531 -11245 19543 -11211
rect 19543 -11245 19565 -11211
rect 19603 -11245 19611 -11211
rect 19611 -11245 19637 -11211
rect 19675 -11245 19679 -11211
rect 19679 -11245 19709 -11211
rect 19747 -11245 19781 -11211
rect 19819 -11245 19849 -11211
rect 19849 -11245 19853 -11211
rect 19891 -11245 19917 -11211
rect 19917 -11245 19925 -11211
rect 19963 -11245 19985 -11211
rect 19985 -11245 19997 -11211
rect 20035 -11245 20053 -11211
rect 20053 -11245 20069 -11211
rect 20107 -11245 20121 -11211
rect 20121 -11245 20141 -11211
rect 20179 -11245 20189 -11211
rect 20189 -11245 20213 -11211
rect 20251 -11245 20257 -11211
rect 20257 -11245 20285 -11211
rect 20323 -11245 20325 -11211
rect 20325 -11245 20357 -11211
rect 20395 -11245 20427 -11211
rect 20427 -11245 20429 -11211
rect 20467 -11245 20495 -11211
rect 20495 -11245 20501 -11211
rect 20539 -11245 20563 -11211
rect 20563 -11245 20573 -11211
rect 20611 -11245 20631 -11211
rect 20631 -11245 20645 -11211
rect 20683 -11245 20699 -11211
rect 20699 -11245 20717 -11211
rect 20755 -11245 20767 -11211
rect 20767 -11245 20789 -11211
rect 20827 -11245 20835 -11211
rect 20835 -11245 20861 -11211
rect 20899 -11245 20903 -11211
rect 20903 -11245 20933 -11211
rect 20971 -11245 21005 -11211
rect 21043 -11245 21073 -11211
rect 21073 -11245 21077 -11211
rect 21115 -11245 21141 -11211
rect 21141 -11245 21149 -11211
rect 21187 -11245 21209 -11211
rect 21209 -11245 21221 -11211
rect 21259 -11245 21277 -11211
rect 21277 -11245 21293 -11211
rect 21331 -11245 21345 -11211
rect 21345 -11245 21365 -11211
rect 21403 -11245 21413 -11211
rect 21413 -11245 21437 -11211
rect 21475 -11245 21481 -11211
rect 21481 -11245 21509 -11211
rect 21547 -11245 21549 -11211
rect 21549 -11245 21581 -11211
rect 21619 -11245 21651 -11211
rect 21651 -11245 21653 -11211
rect 21691 -11245 21719 -11211
rect 21719 -11245 21725 -11211
rect 21763 -11245 21787 -11211
rect 21787 -11245 21797 -11211
rect 21835 -11245 21855 -11211
rect 21855 -11245 21869 -11211
rect 21907 -11245 21923 -11211
rect 21923 -11245 21941 -11211
rect 21979 -11245 21991 -11211
rect 21991 -11245 22013 -11211
rect 22051 -11245 22059 -11211
rect 22059 -11245 22085 -11211
rect 22123 -11245 22127 -11211
rect 22127 -11245 22157 -11211
rect 22195 -11245 22229 -11211
rect 22267 -11245 22297 -11211
rect 22297 -11245 22301 -11211
rect 22339 -11245 22365 -11211
rect 22365 -11245 22373 -11211
rect 22411 -11245 22433 -11211
rect 22433 -11245 22445 -11211
rect 22483 -11245 22501 -11211
rect 22501 -11245 22517 -11211
rect 22555 -11245 22569 -11211
rect 22569 -11245 22589 -11211
rect 22627 -11245 22637 -11211
rect 22637 -11245 22661 -11211
rect 22699 -11245 22705 -11211
rect 22705 -11245 22733 -11211
rect 22771 -11245 22773 -11211
rect 22773 -11245 22805 -11211
rect 22843 -11245 22875 -11211
rect 22875 -11245 22877 -11211
rect 22915 -11245 22943 -11211
rect 22943 -11245 22949 -11211
rect 22987 -11245 23011 -11211
rect 23011 -11245 23021 -11211
rect 23059 -11245 23079 -11211
rect 23079 -11245 23093 -11211
rect 23131 -11245 23147 -11211
rect 23147 -11245 23165 -11211
rect 23203 -11245 23215 -11211
rect 23215 -11245 23237 -11211
rect 23275 -11245 23283 -11211
rect 23283 -11245 23309 -11211
rect 23347 -11245 23351 -11211
rect 23351 -11245 23381 -11211
rect 23419 -11245 23453 -11211
rect 23491 -11245 23521 -11211
rect 23521 -11245 23525 -11211
rect 23563 -11245 23589 -11211
rect 23589 -11245 23597 -11211
rect 23635 -11245 23657 -11211
rect 23657 -11245 23669 -11211
rect 23707 -11245 23725 -11211
rect 23725 -11245 23741 -11211
rect 23779 -11245 23793 -11211
rect 23793 -11245 23813 -11211
rect 23851 -11245 23861 -11211
rect 23861 -11245 23885 -11211
rect 23923 -11245 23929 -11211
rect 23929 -11245 23957 -11211
rect 23995 -11245 23997 -11211
rect 23997 -11245 24029 -11211
rect 24067 -11245 24099 -11211
rect 24099 -11245 24101 -11211
rect 24139 -11245 24167 -11211
rect 24167 -11245 24173 -11211
rect 24211 -11245 24235 -11211
rect 24235 -11245 24245 -11211
rect 24283 -11245 24303 -11211
rect 24303 -11245 24317 -11211
rect 24355 -11245 24371 -11211
rect 24371 -11245 24389 -11211
rect 24427 -11245 24439 -11211
rect 24439 -11245 24461 -11211
rect 24499 -11245 24507 -11211
rect 24507 -11245 24533 -11211
rect 24571 -11245 24575 -11211
rect 24575 -11245 24605 -11211
rect 24643 -11245 24677 -11211
rect 24715 -11245 24745 -11211
rect 24745 -11245 24749 -11211
rect 24787 -11245 24821 -11211
rect 2911 -11680 2921 -11646
rect 2921 -11680 2945 -11646
rect 2983 -11680 2989 -11646
rect 2989 -11680 3017 -11646
rect 3055 -11680 3057 -11646
rect 3057 -11680 3089 -11646
rect 3127 -11680 3159 -11646
rect 3159 -11680 3161 -11646
rect 3199 -11680 3227 -11646
rect 3227 -11680 3233 -11646
rect 3271 -11680 3295 -11646
rect 3295 -11680 3305 -11646
rect 3929 -11680 3939 -11646
rect 3939 -11680 3963 -11646
rect 4001 -11680 4007 -11646
rect 4007 -11680 4035 -11646
rect 4073 -11680 4075 -11646
rect 4075 -11680 4107 -11646
rect 4145 -11680 4177 -11646
rect 4177 -11680 4179 -11646
rect 4217 -11680 4245 -11646
rect 4245 -11680 4251 -11646
rect 4289 -11680 4313 -11646
rect 4313 -11680 4323 -11646
rect 4947 -11680 4957 -11646
rect 4957 -11680 4981 -11646
rect 5019 -11680 5025 -11646
rect 5025 -11680 5053 -11646
rect 5091 -11680 5093 -11646
rect 5093 -11680 5125 -11646
rect 5163 -11680 5195 -11646
rect 5195 -11680 5197 -11646
rect 5235 -11680 5263 -11646
rect 5263 -11680 5269 -11646
rect 5307 -11680 5331 -11646
rect 5331 -11680 5341 -11646
rect 5965 -11680 5975 -11646
rect 5975 -11680 5999 -11646
rect 6037 -11680 6043 -11646
rect 6043 -11680 6071 -11646
rect 6109 -11680 6111 -11646
rect 6111 -11680 6143 -11646
rect 6181 -11680 6213 -11646
rect 6213 -11680 6215 -11646
rect 6253 -11680 6281 -11646
rect 6281 -11680 6287 -11646
rect 6325 -11680 6349 -11646
rect 6349 -11680 6359 -11646
rect 6983 -11680 6993 -11646
rect 6993 -11680 7017 -11646
rect 7055 -11680 7061 -11646
rect 7061 -11680 7089 -11646
rect 7127 -11680 7129 -11646
rect 7129 -11680 7161 -11646
rect 7199 -11680 7231 -11646
rect 7231 -11680 7233 -11646
rect 7271 -11680 7299 -11646
rect 7299 -11680 7305 -11646
rect 7343 -11680 7367 -11646
rect 7367 -11680 7377 -11646
rect 8001 -11680 8011 -11646
rect 8011 -11680 8035 -11646
rect 8073 -11680 8079 -11646
rect 8079 -11680 8107 -11646
rect 8145 -11680 8147 -11646
rect 8147 -11680 8179 -11646
rect 8217 -11680 8249 -11646
rect 8249 -11680 8251 -11646
rect 8289 -11680 8317 -11646
rect 8317 -11680 8323 -11646
rect 8361 -11680 8385 -11646
rect 8385 -11680 8395 -11646
rect 9019 -11680 9029 -11646
rect 9029 -11680 9053 -11646
rect 9091 -11680 9097 -11646
rect 9097 -11680 9125 -11646
rect 9163 -11680 9165 -11646
rect 9165 -11680 9197 -11646
rect 9235 -11680 9267 -11646
rect 9267 -11680 9269 -11646
rect 9307 -11680 9335 -11646
rect 9335 -11680 9341 -11646
rect 9379 -11680 9403 -11646
rect 9403 -11680 9413 -11646
rect 10037 -11680 10047 -11646
rect 10047 -11680 10071 -11646
rect 10109 -11680 10115 -11646
rect 10115 -11680 10143 -11646
rect 10181 -11680 10183 -11646
rect 10183 -11680 10215 -11646
rect 10253 -11680 10285 -11646
rect 10285 -11680 10287 -11646
rect 10325 -11680 10353 -11646
rect 10353 -11680 10359 -11646
rect 10397 -11680 10421 -11646
rect 10421 -11680 10431 -11646
rect 11055 -11680 11065 -11646
rect 11065 -11680 11089 -11646
rect 11127 -11680 11133 -11646
rect 11133 -11680 11161 -11646
rect 11199 -11680 11201 -11646
rect 11201 -11680 11233 -11646
rect 11271 -11680 11303 -11646
rect 11303 -11680 11305 -11646
rect 11343 -11680 11371 -11646
rect 11371 -11680 11377 -11646
rect 11415 -11680 11439 -11646
rect 11439 -11680 11449 -11646
rect 12073 -11680 12083 -11646
rect 12083 -11680 12107 -11646
rect 12145 -11680 12151 -11646
rect 12151 -11680 12179 -11646
rect 12217 -11680 12219 -11646
rect 12219 -11680 12251 -11646
rect 12289 -11680 12321 -11646
rect 12321 -11680 12323 -11646
rect 12361 -11680 12389 -11646
rect 12389 -11680 12395 -11646
rect 12433 -11680 12457 -11646
rect 12457 -11680 12467 -11646
rect 13091 -11680 13101 -11646
rect 13101 -11680 13125 -11646
rect 13163 -11680 13169 -11646
rect 13169 -11680 13197 -11646
rect 13235 -11680 13237 -11646
rect 13237 -11680 13269 -11646
rect 13307 -11680 13339 -11646
rect 13339 -11680 13341 -11646
rect 13379 -11680 13407 -11646
rect 13407 -11680 13413 -11646
rect 13451 -11680 13475 -11646
rect 13475 -11680 13485 -11646
rect 14109 -11680 14119 -11646
rect 14119 -11680 14143 -11646
rect 14181 -11680 14187 -11646
rect 14187 -11680 14215 -11646
rect 14253 -11680 14255 -11646
rect 14255 -11680 14287 -11646
rect 14325 -11680 14357 -11646
rect 14357 -11680 14359 -11646
rect 14397 -11680 14425 -11646
rect 14425 -11680 14431 -11646
rect 14469 -11680 14493 -11646
rect 14493 -11680 14503 -11646
rect 15127 -11680 15137 -11646
rect 15137 -11680 15161 -11646
rect 15199 -11680 15205 -11646
rect 15205 -11680 15233 -11646
rect 15271 -11680 15273 -11646
rect 15273 -11680 15305 -11646
rect 15343 -11680 15375 -11646
rect 15375 -11680 15377 -11646
rect 15415 -11680 15443 -11646
rect 15443 -11680 15449 -11646
rect 15487 -11680 15511 -11646
rect 15511 -11680 15521 -11646
rect 16145 -11680 16155 -11646
rect 16155 -11680 16179 -11646
rect 16217 -11680 16223 -11646
rect 16223 -11680 16251 -11646
rect 16289 -11680 16291 -11646
rect 16291 -11680 16323 -11646
rect 16361 -11680 16393 -11646
rect 16393 -11680 16395 -11646
rect 16433 -11680 16461 -11646
rect 16461 -11680 16467 -11646
rect 16505 -11680 16529 -11646
rect 16529 -11680 16539 -11646
rect 17163 -11680 17173 -11646
rect 17173 -11680 17197 -11646
rect 17235 -11680 17241 -11646
rect 17241 -11680 17269 -11646
rect 17307 -11680 17309 -11646
rect 17309 -11680 17341 -11646
rect 17379 -11680 17411 -11646
rect 17411 -11680 17413 -11646
rect 17451 -11680 17479 -11646
rect 17479 -11680 17485 -11646
rect 17523 -11680 17547 -11646
rect 17547 -11680 17557 -11646
rect 18181 -11680 18191 -11646
rect 18191 -11680 18215 -11646
rect 18253 -11680 18259 -11646
rect 18259 -11680 18287 -11646
rect 18325 -11680 18327 -11646
rect 18327 -11680 18359 -11646
rect 18397 -11680 18429 -11646
rect 18429 -11680 18431 -11646
rect 18469 -11680 18497 -11646
rect 18497 -11680 18503 -11646
rect 18541 -11680 18565 -11646
rect 18565 -11680 18575 -11646
rect 19199 -11680 19209 -11646
rect 19209 -11680 19233 -11646
rect 19271 -11680 19277 -11646
rect 19277 -11680 19305 -11646
rect 19343 -11680 19345 -11646
rect 19345 -11680 19377 -11646
rect 19415 -11680 19447 -11646
rect 19447 -11680 19449 -11646
rect 19487 -11680 19515 -11646
rect 19515 -11680 19521 -11646
rect 19559 -11680 19583 -11646
rect 19583 -11680 19593 -11646
rect 20217 -11680 20227 -11646
rect 20227 -11680 20251 -11646
rect 20289 -11680 20295 -11646
rect 20295 -11680 20323 -11646
rect 20361 -11680 20363 -11646
rect 20363 -11680 20395 -11646
rect 20433 -11680 20465 -11646
rect 20465 -11680 20467 -11646
rect 20505 -11680 20533 -11646
rect 20533 -11680 20539 -11646
rect 20577 -11680 20601 -11646
rect 20601 -11680 20611 -11646
rect 21235 -11680 21245 -11646
rect 21245 -11680 21269 -11646
rect 21307 -11680 21313 -11646
rect 21313 -11680 21341 -11646
rect 21379 -11680 21381 -11646
rect 21381 -11680 21413 -11646
rect 21451 -11680 21483 -11646
rect 21483 -11680 21485 -11646
rect 21523 -11680 21551 -11646
rect 21551 -11680 21557 -11646
rect 21595 -11680 21619 -11646
rect 21619 -11680 21629 -11646
rect 22253 -11680 22263 -11646
rect 22263 -11680 22287 -11646
rect 22325 -11680 22331 -11646
rect 22331 -11680 22359 -11646
rect 22397 -11680 22399 -11646
rect 22399 -11680 22431 -11646
rect 22469 -11680 22501 -11646
rect 22501 -11680 22503 -11646
rect 22541 -11680 22569 -11646
rect 22569 -11680 22575 -11646
rect 22613 -11680 22637 -11646
rect 22637 -11680 22647 -11646
rect -12289 -12111 -12255 -12091
rect -12289 -12125 -12255 -12111
rect -12289 -12179 -12255 -12163
rect -12289 -12197 -12255 -12179
rect -12289 -12247 -12255 -12235
rect -12289 -12269 -12255 -12247
rect -12289 -12315 -12255 -12307
rect -12289 -12341 -12255 -12315
rect 2582 -11763 2616 -11749
rect 2582 -11783 2616 -11763
rect 2582 -11831 2616 -11821
rect 2582 -11855 2616 -11831
rect 2582 -11899 2616 -11893
rect 2582 -11927 2616 -11899
rect 2582 -11967 2616 -11965
rect 2582 -11999 2616 -11967
rect 2582 -12069 2616 -12037
rect 2582 -12071 2616 -12069
rect 2582 -12137 2616 -12109
rect 2582 -12143 2616 -12137
rect 2582 -12205 2616 -12181
rect 2582 -12215 2616 -12205
rect 2582 -12273 2616 -12253
rect 2582 -12287 2616 -12273
rect 3600 -11763 3634 -11749
rect 3600 -11783 3634 -11763
rect 3600 -11831 3634 -11821
rect 3600 -11855 3634 -11831
rect 3600 -11899 3634 -11893
rect 3600 -11927 3634 -11899
rect 3600 -11967 3634 -11965
rect 3600 -11999 3634 -11967
rect 3600 -12069 3634 -12037
rect 3600 -12071 3634 -12069
rect 3600 -12137 3634 -12109
rect 3600 -12143 3634 -12137
rect 3600 -12205 3634 -12181
rect 3600 -12215 3634 -12205
rect 3600 -12273 3634 -12253
rect 3600 -12287 3634 -12273
rect 4618 -11763 4652 -11749
rect 4618 -11783 4652 -11763
rect 4618 -11831 4652 -11821
rect 4618 -11855 4652 -11831
rect 4618 -11899 4652 -11893
rect 4618 -11927 4652 -11899
rect 4618 -11967 4652 -11965
rect 4618 -11999 4652 -11967
rect 4618 -12069 4652 -12037
rect 4618 -12071 4652 -12069
rect 4618 -12137 4652 -12109
rect 4618 -12143 4652 -12137
rect 4618 -12205 4652 -12181
rect 4618 -12215 4652 -12205
rect 4618 -12273 4652 -12253
rect 4618 -12287 4652 -12273
rect 5636 -11763 5670 -11749
rect 5636 -11783 5670 -11763
rect 5636 -11831 5670 -11821
rect 5636 -11855 5670 -11831
rect 5636 -11899 5670 -11893
rect 5636 -11927 5670 -11899
rect 5636 -11967 5670 -11965
rect 5636 -11999 5670 -11967
rect 5636 -12069 5670 -12037
rect 5636 -12071 5670 -12069
rect 5636 -12137 5670 -12109
rect 5636 -12143 5670 -12137
rect 5636 -12205 5670 -12181
rect 5636 -12215 5670 -12205
rect 5636 -12273 5670 -12253
rect 5636 -12287 5670 -12273
rect 6654 -11763 6688 -11749
rect 6654 -11783 6688 -11763
rect 6654 -11831 6688 -11821
rect 6654 -11855 6688 -11831
rect 6654 -11899 6688 -11893
rect 6654 -11927 6688 -11899
rect 6654 -11967 6688 -11965
rect 6654 -11999 6688 -11967
rect 6654 -12069 6688 -12037
rect 6654 -12071 6688 -12069
rect 6654 -12137 6688 -12109
rect 6654 -12143 6688 -12137
rect 6654 -12205 6688 -12181
rect 6654 -12215 6688 -12205
rect 6654 -12273 6688 -12253
rect 6654 -12287 6688 -12273
rect 7672 -11763 7706 -11749
rect 7672 -11783 7706 -11763
rect 7672 -11831 7706 -11821
rect 7672 -11855 7706 -11831
rect 7672 -11899 7706 -11893
rect 7672 -11927 7706 -11899
rect 7672 -11967 7706 -11965
rect 7672 -11999 7706 -11967
rect 7672 -12069 7706 -12037
rect 7672 -12071 7706 -12069
rect 7672 -12137 7706 -12109
rect 7672 -12143 7706 -12137
rect 7672 -12205 7706 -12181
rect 7672 -12215 7706 -12205
rect 7672 -12273 7706 -12253
rect 7672 -12287 7706 -12273
rect 8690 -11763 8724 -11749
rect 8690 -11783 8724 -11763
rect 8690 -11831 8724 -11821
rect 8690 -11855 8724 -11831
rect 8690 -11899 8724 -11893
rect 8690 -11927 8724 -11899
rect 8690 -11967 8724 -11965
rect 8690 -11999 8724 -11967
rect 8690 -12069 8724 -12037
rect 8690 -12071 8724 -12069
rect 8690 -12137 8724 -12109
rect 8690 -12143 8724 -12137
rect 8690 -12205 8724 -12181
rect 8690 -12215 8724 -12205
rect 8690 -12273 8724 -12253
rect 8690 -12287 8724 -12273
rect 9708 -11763 9742 -11749
rect 9708 -11783 9742 -11763
rect 9708 -11831 9742 -11821
rect 9708 -11855 9742 -11831
rect 9708 -11899 9742 -11893
rect 9708 -11927 9742 -11899
rect 9708 -11967 9742 -11965
rect 9708 -11999 9742 -11967
rect 9708 -12069 9742 -12037
rect 9708 -12071 9742 -12069
rect 9708 -12137 9742 -12109
rect 9708 -12143 9742 -12137
rect 9708 -12205 9742 -12181
rect 9708 -12215 9742 -12205
rect 9708 -12273 9742 -12253
rect 9708 -12287 9742 -12273
rect 10726 -11763 10760 -11749
rect 10726 -11783 10760 -11763
rect 10726 -11831 10760 -11821
rect 10726 -11855 10760 -11831
rect 10726 -11899 10760 -11893
rect 10726 -11927 10760 -11899
rect 10726 -11967 10760 -11965
rect 10726 -11999 10760 -11967
rect 10726 -12069 10760 -12037
rect 10726 -12071 10760 -12069
rect 10726 -12137 10760 -12109
rect 10726 -12143 10760 -12137
rect 10726 -12205 10760 -12181
rect 10726 -12215 10760 -12205
rect 10726 -12273 10760 -12253
rect 10726 -12287 10760 -12273
rect 11744 -11763 11778 -11749
rect 11744 -11783 11778 -11763
rect 11744 -11831 11778 -11821
rect 11744 -11855 11778 -11831
rect 11744 -11899 11778 -11893
rect 11744 -11927 11778 -11899
rect 11744 -11967 11778 -11965
rect 11744 -11999 11778 -11967
rect 11744 -12069 11778 -12037
rect 11744 -12071 11778 -12069
rect 11744 -12137 11778 -12109
rect 11744 -12143 11778 -12137
rect 11744 -12205 11778 -12181
rect 11744 -12215 11778 -12205
rect 11744 -12273 11778 -12253
rect 11744 -12287 11778 -12273
rect 12762 -11763 12796 -11749
rect 12762 -11783 12796 -11763
rect 12762 -11831 12796 -11821
rect 12762 -11855 12796 -11831
rect 12762 -11899 12796 -11893
rect 12762 -11927 12796 -11899
rect 12762 -11967 12796 -11965
rect 12762 -11999 12796 -11967
rect 12762 -12069 12796 -12037
rect 12762 -12071 12796 -12069
rect 12762 -12137 12796 -12109
rect 12762 -12143 12796 -12137
rect 12762 -12205 12796 -12181
rect 12762 -12215 12796 -12205
rect 12762 -12273 12796 -12253
rect 12762 -12287 12796 -12273
rect 13780 -11763 13814 -11749
rect 13780 -11783 13814 -11763
rect 13780 -11831 13814 -11821
rect 13780 -11855 13814 -11831
rect 13780 -11899 13814 -11893
rect 13780 -11927 13814 -11899
rect 13780 -11967 13814 -11965
rect 13780 -11999 13814 -11967
rect 13780 -12069 13814 -12037
rect 13780 -12071 13814 -12069
rect 13780 -12137 13814 -12109
rect 13780 -12143 13814 -12137
rect 13780 -12205 13814 -12181
rect 13780 -12215 13814 -12205
rect 13780 -12273 13814 -12253
rect 13780 -12287 13814 -12273
rect 14798 -11763 14832 -11749
rect 14798 -11783 14832 -11763
rect 14798 -11831 14832 -11821
rect 14798 -11855 14832 -11831
rect 14798 -11899 14832 -11893
rect 14798 -11927 14832 -11899
rect 14798 -11967 14832 -11965
rect 14798 -11999 14832 -11967
rect 14798 -12069 14832 -12037
rect 14798 -12071 14832 -12069
rect 14798 -12137 14832 -12109
rect 14798 -12143 14832 -12137
rect 14798 -12205 14832 -12181
rect 14798 -12215 14832 -12205
rect 14798 -12273 14832 -12253
rect 14798 -12287 14832 -12273
rect 15816 -11763 15850 -11749
rect 15816 -11783 15850 -11763
rect 15816 -11831 15850 -11821
rect 15816 -11855 15850 -11831
rect 15816 -11899 15850 -11893
rect 15816 -11927 15850 -11899
rect 15816 -11967 15850 -11965
rect 15816 -11999 15850 -11967
rect 15816 -12069 15850 -12037
rect 15816 -12071 15850 -12069
rect 15816 -12137 15850 -12109
rect 15816 -12143 15850 -12137
rect 15816 -12205 15850 -12181
rect 15816 -12215 15850 -12205
rect 15816 -12273 15850 -12253
rect 15816 -12287 15850 -12273
rect 16834 -11763 16868 -11749
rect 16834 -11783 16868 -11763
rect 16834 -11831 16868 -11821
rect 16834 -11855 16868 -11831
rect 16834 -11899 16868 -11893
rect 16834 -11927 16868 -11899
rect 16834 -11967 16868 -11965
rect 16834 -11999 16868 -11967
rect 16834 -12069 16868 -12037
rect 16834 -12071 16868 -12069
rect 16834 -12137 16868 -12109
rect 16834 -12143 16868 -12137
rect 16834 -12205 16868 -12181
rect 16834 -12215 16868 -12205
rect 16834 -12273 16868 -12253
rect 16834 -12287 16868 -12273
rect 17852 -11763 17886 -11749
rect 17852 -11783 17886 -11763
rect 17852 -11831 17886 -11821
rect 17852 -11855 17886 -11831
rect 17852 -11899 17886 -11893
rect 17852 -11927 17886 -11899
rect 17852 -11967 17886 -11965
rect 17852 -11999 17886 -11967
rect 17852 -12069 17886 -12037
rect 17852 -12071 17886 -12069
rect 17852 -12137 17886 -12109
rect 17852 -12143 17886 -12137
rect 17852 -12205 17886 -12181
rect 17852 -12215 17886 -12205
rect 17852 -12273 17886 -12253
rect 17852 -12287 17886 -12273
rect 18870 -11763 18904 -11749
rect 18870 -11783 18904 -11763
rect 18870 -11831 18904 -11821
rect 18870 -11855 18904 -11831
rect 18870 -11899 18904 -11893
rect 18870 -11927 18904 -11899
rect 18870 -11967 18904 -11965
rect 18870 -11999 18904 -11967
rect 18870 -12069 18904 -12037
rect 18870 -12071 18904 -12069
rect 18870 -12137 18904 -12109
rect 18870 -12143 18904 -12137
rect 18870 -12205 18904 -12181
rect 18870 -12215 18904 -12205
rect 18870 -12273 18904 -12253
rect 18870 -12287 18904 -12273
rect 19888 -11763 19922 -11749
rect 19888 -11783 19922 -11763
rect 19888 -11831 19922 -11821
rect 19888 -11855 19922 -11831
rect 19888 -11899 19922 -11893
rect 19888 -11927 19922 -11899
rect 19888 -11967 19922 -11965
rect 19888 -11999 19922 -11967
rect 19888 -12069 19922 -12037
rect 19888 -12071 19922 -12069
rect 19888 -12137 19922 -12109
rect 19888 -12143 19922 -12137
rect 19888 -12205 19922 -12181
rect 19888 -12215 19922 -12205
rect 19888 -12273 19922 -12253
rect 19888 -12287 19922 -12273
rect 20906 -11763 20940 -11749
rect 20906 -11783 20940 -11763
rect 20906 -11831 20940 -11821
rect 20906 -11855 20940 -11831
rect 20906 -11899 20940 -11893
rect 20906 -11927 20940 -11899
rect 20906 -11967 20940 -11965
rect 20906 -11999 20940 -11967
rect 20906 -12069 20940 -12037
rect 20906 -12071 20940 -12069
rect 20906 -12137 20940 -12109
rect 20906 -12143 20940 -12137
rect 20906 -12205 20940 -12181
rect 20906 -12215 20940 -12205
rect 20906 -12273 20940 -12253
rect 20906 -12287 20940 -12273
rect 21924 -11763 21958 -11749
rect 21924 -11783 21958 -11763
rect 21924 -11831 21958 -11821
rect 21924 -11855 21958 -11831
rect 21924 -11899 21958 -11893
rect 21924 -11927 21958 -11899
rect 21924 -11967 21958 -11965
rect 21924 -11999 21958 -11967
rect 21924 -12069 21958 -12037
rect 21924 -12071 21958 -12069
rect 21924 -12137 21958 -12109
rect 21924 -12143 21958 -12137
rect 21924 -12205 21958 -12181
rect 21924 -12215 21958 -12205
rect 21924 -12273 21958 -12253
rect 21924 -12287 21958 -12273
rect 22942 -11763 22976 -11749
rect 22942 -11783 22976 -11763
rect 22942 -11831 22976 -11821
rect 22942 -11855 22976 -11831
rect 22942 -11899 22976 -11893
rect 22942 -11927 22976 -11899
rect 22942 -11967 22976 -11965
rect 22942 -11999 22976 -11967
rect 22942 -12069 22976 -12037
rect 22942 -12071 22976 -12069
rect 22942 -12137 22976 -12109
rect 22942 -12143 22976 -12137
rect 22942 -12205 22976 -12181
rect 22942 -12215 22976 -12205
rect 22942 -12273 22976 -12253
rect 22942 -12287 22976 -12273
rect 24855 -12111 24889 -12091
rect 24855 -12125 24889 -12111
rect 24855 -12179 24889 -12163
rect 24855 -12197 24889 -12179
rect 24855 -12247 24889 -12235
rect 24855 -12269 24889 -12247
rect 24855 -12315 24889 -12307
rect 24855 -12341 24889 -12315
rect -12289 -12383 -12255 -12379
rect -12289 -12413 -12255 -12383
rect 2911 -12390 2921 -12356
rect 2921 -12390 2945 -12356
rect 2983 -12390 2989 -12356
rect 2989 -12390 3017 -12356
rect 3055 -12390 3057 -12356
rect 3057 -12390 3089 -12356
rect 3127 -12390 3159 -12356
rect 3159 -12390 3161 -12356
rect 3199 -12390 3227 -12356
rect 3227 -12390 3233 -12356
rect 3271 -12390 3295 -12356
rect 3295 -12390 3305 -12356
rect 3929 -12390 3939 -12356
rect 3939 -12390 3963 -12356
rect 4001 -12390 4007 -12356
rect 4007 -12390 4035 -12356
rect 4073 -12390 4075 -12356
rect 4075 -12390 4107 -12356
rect 4145 -12390 4177 -12356
rect 4177 -12390 4179 -12356
rect 4217 -12390 4245 -12356
rect 4245 -12390 4251 -12356
rect 4289 -12390 4313 -12356
rect 4313 -12390 4323 -12356
rect 4947 -12390 4957 -12356
rect 4957 -12390 4981 -12356
rect 5019 -12390 5025 -12356
rect 5025 -12390 5053 -12356
rect 5091 -12390 5093 -12356
rect 5093 -12390 5125 -12356
rect 5163 -12390 5195 -12356
rect 5195 -12390 5197 -12356
rect 5235 -12390 5263 -12356
rect 5263 -12390 5269 -12356
rect 5307 -12390 5331 -12356
rect 5331 -12390 5341 -12356
rect 5965 -12390 5975 -12356
rect 5975 -12390 5999 -12356
rect 6037 -12390 6043 -12356
rect 6043 -12390 6071 -12356
rect 6109 -12390 6111 -12356
rect 6111 -12390 6143 -12356
rect 6181 -12390 6213 -12356
rect 6213 -12390 6215 -12356
rect 6253 -12390 6281 -12356
rect 6281 -12390 6287 -12356
rect 6325 -12390 6349 -12356
rect 6349 -12390 6359 -12356
rect 6983 -12390 6993 -12356
rect 6993 -12390 7017 -12356
rect 7055 -12390 7061 -12356
rect 7061 -12390 7089 -12356
rect 7127 -12390 7129 -12356
rect 7129 -12390 7161 -12356
rect 7199 -12390 7231 -12356
rect 7231 -12390 7233 -12356
rect 7271 -12390 7299 -12356
rect 7299 -12390 7305 -12356
rect 7343 -12390 7367 -12356
rect 7367 -12390 7377 -12356
rect 8001 -12390 8011 -12356
rect 8011 -12390 8035 -12356
rect 8073 -12390 8079 -12356
rect 8079 -12390 8107 -12356
rect 8145 -12390 8147 -12356
rect 8147 -12390 8179 -12356
rect 8217 -12390 8249 -12356
rect 8249 -12390 8251 -12356
rect 8289 -12390 8317 -12356
rect 8317 -12390 8323 -12356
rect 8361 -12390 8385 -12356
rect 8385 -12390 8395 -12356
rect 9019 -12390 9029 -12356
rect 9029 -12390 9053 -12356
rect 9091 -12390 9097 -12356
rect 9097 -12390 9125 -12356
rect 9163 -12390 9165 -12356
rect 9165 -12390 9197 -12356
rect 9235 -12390 9267 -12356
rect 9267 -12390 9269 -12356
rect 9307 -12390 9335 -12356
rect 9335 -12390 9341 -12356
rect 9379 -12390 9403 -12356
rect 9403 -12390 9413 -12356
rect 10037 -12390 10047 -12356
rect 10047 -12390 10071 -12356
rect 10109 -12390 10115 -12356
rect 10115 -12390 10143 -12356
rect 10181 -12390 10183 -12356
rect 10183 -12390 10215 -12356
rect 10253 -12390 10285 -12356
rect 10285 -12390 10287 -12356
rect 10325 -12390 10353 -12356
rect 10353 -12390 10359 -12356
rect 10397 -12390 10421 -12356
rect 10421 -12390 10431 -12356
rect 11055 -12390 11065 -12356
rect 11065 -12390 11089 -12356
rect 11127 -12390 11133 -12356
rect 11133 -12390 11161 -12356
rect 11199 -12390 11201 -12356
rect 11201 -12390 11233 -12356
rect 11271 -12390 11303 -12356
rect 11303 -12390 11305 -12356
rect 11343 -12390 11371 -12356
rect 11371 -12390 11377 -12356
rect 11415 -12390 11439 -12356
rect 11439 -12390 11449 -12356
rect 12073 -12390 12083 -12356
rect 12083 -12390 12107 -12356
rect 12145 -12390 12151 -12356
rect 12151 -12390 12179 -12356
rect 12217 -12390 12219 -12356
rect 12219 -12390 12251 -12356
rect 12289 -12390 12321 -12356
rect 12321 -12390 12323 -12356
rect 12361 -12390 12389 -12356
rect 12389 -12390 12395 -12356
rect 12433 -12390 12457 -12356
rect 12457 -12390 12467 -12356
rect 13091 -12390 13101 -12356
rect 13101 -12390 13125 -12356
rect 13163 -12390 13169 -12356
rect 13169 -12390 13197 -12356
rect 13235 -12390 13237 -12356
rect 13237 -12390 13269 -12356
rect 13307 -12390 13339 -12356
rect 13339 -12390 13341 -12356
rect 13379 -12390 13407 -12356
rect 13407 -12390 13413 -12356
rect 13451 -12390 13475 -12356
rect 13475 -12390 13485 -12356
rect 14109 -12390 14119 -12356
rect 14119 -12390 14143 -12356
rect 14181 -12390 14187 -12356
rect 14187 -12390 14215 -12356
rect 14253 -12390 14255 -12356
rect 14255 -12390 14287 -12356
rect 14325 -12390 14357 -12356
rect 14357 -12390 14359 -12356
rect 14397 -12390 14425 -12356
rect 14425 -12390 14431 -12356
rect 14469 -12390 14493 -12356
rect 14493 -12390 14503 -12356
rect 15127 -12390 15137 -12356
rect 15137 -12390 15161 -12356
rect 15199 -12390 15205 -12356
rect 15205 -12390 15233 -12356
rect 15271 -12390 15273 -12356
rect 15273 -12390 15305 -12356
rect 15343 -12390 15375 -12356
rect 15375 -12390 15377 -12356
rect 15415 -12390 15443 -12356
rect 15443 -12390 15449 -12356
rect 15487 -12390 15511 -12356
rect 15511 -12390 15521 -12356
rect 16145 -12390 16155 -12356
rect 16155 -12390 16179 -12356
rect 16217 -12390 16223 -12356
rect 16223 -12390 16251 -12356
rect 16289 -12390 16291 -12356
rect 16291 -12390 16323 -12356
rect 16361 -12390 16393 -12356
rect 16393 -12390 16395 -12356
rect 16433 -12390 16461 -12356
rect 16461 -12390 16467 -12356
rect 16505 -12390 16529 -12356
rect 16529 -12390 16539 -12356
rect 17163 -12390 17173 -12356
rect 17173 -12390 17197 -12356
rect 17235 -12390 17241 -12356
rect 17241 -12390 17269 -12356
rect 17307 -12390 17309 -12356
rect 17309 -12390 17341 -12356
rect 17379 -12390 17411 -12356
rect 17411 -12390 17413 -12356
rect 17451 -12390 17479 -12356
rect 17479 -12390 17485 -12356
rect 17523 -12390 17547 -12356
rect 17547 -12390 17557 -12356
rect 18181 -12390 18191 -12356
rect 18191 -12390 18215 -12356
rect 18253 -12390 18259 -12356
rect 18259 -12390 18287 -12356
rect 18325 -12390 18327 -12356
rect 18327 -12390 18359 -12356
rect 18397 -12390 18429 -12356
rect 18429 -12390 18431 -12356
rect 18469 -12390 18497 -12356
rect 18497 -12390 18503 -12356
rect 18541 -12390 18565 -12356
rect 18565 -12390 18575 -12356
rect 19199 -12390 19209 -12356
rect 19209 -12390 19233 -12356
rect 19271 -12390 19277 -12356
rect 19277 -12390 19305 -12356
rect 19343 -12390 19345 -12356
rect 19345 -12390 19377 -12356
rect 19415 -12390 19447 -12356
rect 19447 -12390 19449 -12356
rect 19487 -12390 19515 -12356
rect 19515 -12390 19521 -12356
rect 19559 -12390 19583 -12356
rect 19583 -12390 19593 -12356
rect 20217 -12390 20227 -12356
rect 20227 -12390 20251 -12356
rect 20289 -12390 20295 -12356
rect 20295 -12390 20323 -12356
rect 20361 -12390 20363 -12356
rect 20363 -12390 20395 -12356
rect 20433 -12390 20465 -12356
rect 20465 -12390 20467 -12356
rect 20505 -12390 20533 -12356
rect 20533 -12390 20539 -12356
rect 20577 -12390 20601 -12356
rect 20601 -12390 20611 -12356
rect 21235 -12390 21245 -12356
rect 21245 -12390 21269 -12356
rect 21307 -12390 21313 -12356
rect 21313 -12390 21341 -12356
rect 21379 -12390 21381 -12356
rect 21381 -12390 21413 -12356
rect 21451 -12390 21483 -12356
rect 21483 -12390 21485 -12356
rect 21523 -12390 21551 -12356
rect 21551 -12390 21557 -12356
rect 21595 -12390 21619 -12356
rect 21619 -12390 21629 -12356
rect 22253 -12390 22263 -12356
rect 22263 -12390 22287 -12356
rect 22325 -12390 22331 -12356
rect 22331 -12390 22359 -12356
rect 22397 -12390 22399 -12356
rect 22399 -12390 22431 -12356
rect 22469 -12390 22501 -12356
rect 22501 -12390 22503 -12356
rect 22541 -12390 22569 -12356
rect 22569 -12390 22575 -12356
rect 22613 -12390 22637 -12356
rect 22637 -12390 22647 -12356
rect 24855 -12383 24889 -12379
rect 24855 -12413 24889 -12383
rect -12289 -12485 -12255 -12451
rect -8855 -12474 -8845 -12440
rect -8845 -12474 -8821 -12440
rect -8783 -12474 -8777 -12440
rect -8777 -12474 -8749 -12440
rect -8711 -12474 -8709 -12440
rect -8709 -12474 -8677 -12440
rect -8639 -12474 -8607 -12440
rect -8607 -12474 -8605 -12440
rect -8567 -12474 -8539 -12440
rect -8539 -12474 -8533 -12440
rect -8495 -12474 -8471 -12440
rect -8471 -12474 -8461 -12440
rect -7837 -12474 -7827 -12440
rect -7827 -12474 -7803 -12440
rect -7765 -12474 -7759 -12440
rect -7759 -12474 -7731 -12440
rect -7693 -12474 -7691 -12440
rect -7691 -12474 -7659 -12440
rect -7621 -12474 -7589 -12440
rect -7589 -12474 -7587 -12440
rect -7549 -12474 -7521 -12440
rect -7521 -12474 -7515 -12440
rect -7477 -12474 -7453 -12440
rect -7453 -12474 -7443 -12440
rect -6819 -12474 -6809 -12440
rect -6809 -12474 -6785 -12440
rect -6747 -12474 -6741 -12440
rect -6741 -12474 -6713 -12440
rect -6675 -12474 -6673 -12440
rect -6673 -12474 -6641 -12440
rect -6603 -12474 -6571 -12440
rect -6571 -12474 -6569 -12440
rect -6531 -12474 -6503 -12440
rect -6503 -12474 -6497 -12440
rect -6459 -12474 -6435 -12440
rect -6435 -12474 -6425 -12440
rect -5801 -12474 -5791 -12440
rect -5791 -12474 -5767 -12440
rect -5729 -12474 -5723 -12440
rect -5723 -12474 -5695 -12440
rect -5657 -12474 -5655 -12440
rect -5655 -12474 -5623 -12440
rect -5585 -12474 -5553 -12440
rect -5553 -12474 -5551 -12440
rect -5513 -12474 -5485 -12440
rect -5485 -12474 -5479 -12440
rect -5441 -12474 -5417 -12440
rect -5417 -12474 -5407 -12440
rect -4783 -12474 -4773 -12440
rect -4773 -12474 -4749 -12440
rect -4711 -12474 -4705 -12440
rect -4705 -12474 -4677 -12440
rect -4639 -12474 -4637 -12440
rect -4637 -12474 -4605 -12440
rect -4567 -12474 -4535 -12440
rect -4535 -12474 -4533 -12440
rect -4495 -12474 -4467 -12440
rect -4467 -12474 -4461 -12440
rect -4423 -12474 -4399 -12440
rect -4399 -12474 -4389 -12440
rect -3765 -12474 -3755 -12440
rect -3755 -12474 -3731 -12440
rect -3693 -12474 -3687 -12440
rect -3687 -12474 -3659 -12440
rect -3621 -12474 -3619 -12440
rect -3619 -12474 -3587 -12440
rect -3549 -12474 -3517 -12440
rect -3517 -12474 -3515 -12440
rect -3477 -12474 -3449 -12440
rect -3449 -12474 -3443 -12440
rect -3405 -12474 -3381 -12440
rect -3381 -12474 -3371 -12440
rect -2747 -12474 -2737 -12440
rect -2737 -12474 -2713 -12440
rect -2675 -12474 -2669 -12440
rect -2669 -12474 -2641 -12440
rect -2603 -12474 -2601 -12440
rect -2601 -12474 -2569 -12440
rect -2531 -12474 -2499 -12440
rect -2499 -12474 -2497 -12440
rect -2459 -12474 -2431 -12440
rect -2431 -12474 -2425 -12440
rect -2387 -12474 -2363 -12440
rect -2363 -12474 -2353 -12440
rect -1729 -12474 -1719 -12440
rect -1719 -12474 -1695 -12440
rect -1657 -12474 -1651 -12440
rect -1651 -12474 -1623 -12440
rect -1585 -12474 -1583 -12440
rect -1583 -12474 -1551 -12440
rect -1513 -12474 -1481 -12440
rect -1481 -12474 -1479 -12440
rect -1441 -12474 -1413 -12440
rect -1413 -12474 -1407 -12440
rect -1369 -12474 -1345 -12440
rect -1345 -12474 -1335 -12440
rect -711 -12474 -701 -12440
rect -701 -12474 -677 -12440
rect -639 -12474 -633 -12440
rect -633 -12474 -605 -12440
rect -567 -12474 -565 -12440
rect -565 -12474 -533 -12440
rect -495 -12474 -463 -12440
rect -463 -12474 -461 -12440
rect -423 -12474 -395 -12440
rect -395 -12474 -389 -12440
rect -351 -12474 -327 -12440
rect -327 -12474 -317 -12440
rect 24855 -12485 24889 -12451
rect -12289 -12553 -12255 -12523
rect -12289 -12557 -12255 -12553
rect -12289 -12621 -12255 -12595
rect -12289 -12629 -12255 -12621
rect -12289 -12689 -12255 -12667
rect -12289 -12701 -12255 -12689
rect -12289 -12757 -12255 -12739
rect -12289 -12773 -12255 -12757
rect -12289 -12825 -12255 -12811
rect -12289 -12845 -12255 -12825
rect -12289 -12893 -12255 -12883
rect -12289 -12917 -12255 -12893
rect -12289 -12961 -12255 -12955
rect -12289 -12989 -12255 -12961
rect -12289 -13029 -12255 -13027
rect -12289 -13061 -12255 -13029
rect -12289 -13131 -12255 -13099
rect -12289 -13133 -12255 -13131
rect -9184 -12557 -9150 -12543
rect -9184 -12577 -9150 -12557
rect -9184 -12625 -9150 -12615
rect -9184 -12649 -9150 -12625
rect -9184 -12693 -9150 -12687
rect -9184 -12721 -9150 -12693
rect -9184 -12761 -9150 -12759
rect -9184 -12793 -9150 -12761
rect -9184 -12863 -9150 -12831
rect -9184 -12865 -9150 -12863
rect -9184 -12931 -9150 -12903
rect -9184 -12937 -9150 -12931
rect -9184 -12999 -9150 -12975
rect -9184 -13009 -9150 -12999
rect -9184 -13067 -9150 -13047
rect -9184 -13081 -9150 -13067
rect -8166 -12557 -8132 -12543
rect -8166 -12577 -8132 -12557
rect -8166 -12625 -8132 -12615
rect -8166 -12649 -8132 -12625
rect -8166 -12693 -8132 -12687
rect -8166 -12721 -8132 -12693
rect -8166 -12761 -8132 -12759
rect -8166 -12793 -8132 -12761
rect -8166 -12863 -8132 -12831
rect -8166 -12865 -8132 -12863
rect -8166 -12931 -8132 -12903
rect -8166 -12937 -8132 -12931
rect -8166 -12999 -8132 -12975
rect -8166 -13009 -8132 -12999
rect -8166 -13067 -8132 -13047
rect -8166 -13081 -8132 -13067
rect -7148 -12557 -7114 -12543
rect -7148 -12577 -7114 -12557
rect -7148 -12625 -7114 -12615
rect -7148 -12649 -7114 -12625
rect -7148 -12693 -7114 -12687
rect -7148 -12721 -7114 -12693
rect -7148 -12761 -7114 -12759
rect -7148 -12793 -7114 -12761
rect -7148 -12863 -7114 -12831
rect -7148 -12865 -7114 -12863
rect -7148 -12931 -7114 -12903
rect -7148 -12937 -7114 -12931
rect -7148 -12999 -7114 -12975
rect -7148 -13009 -7114 -12999
rect -7148 -13067 -7114 -13047
rect -7148 -13081 -7114 -13067
rect -6130 -12557 -6096 -12543
rect -6130 -12577 -6096 -12557
rect -6130 -12625 -6096 -12615
rect -6130 -12649 -6096 -12625
rect -6130 -12693 -6096 -12687
rect -6130 -12721 -6096 -12693
rect -6130 -12761 -6096 -12759
rect -6130 -12793 -6096 -12761
rect -6130 -12863 -6096 -12831
rect -6130 -12865 -6096 -12863
rect -6130 -12931 -6096 -12903
rect -6130 -12937 -6096 -12931
rect -6130 -12999 -6096 -12975
rect -6130 -13009 -6096 -12999
rect -6130 -13067 -6096 -13047
rect -6130 -13081 -6096 -13067
rect -5112 -12557 -5078 -12543
rect -5112 -12577 -5078 -12557
rect -5112 -12625 -5078 -12615
rect -5112 -12649 -5078 -12625
rect -5112 -12693 -5078 -12687
rect -5112 -12721 -5078 -12693
rect -5112 -12761 -5078 -12759
rect -5112 -12793 -5078 -12761
rect -5112 -12863 -5078 -12831
rect -5112 -12865 -5078 -12863
rect -5112 -12931 -5078 -12903
rect -5112 -12937 -5078 -12931
rect -5112 -12999 -5078 -12975
rect -5112 -13009 -5078 -12999
rect -5112 -13067 -5078 -13047
rect -5112 -13081 -5078 -13067
rect -4094 -12557 -4060 -12543
rect -4094 -12577 -4060 -12557
rect -4094 -12625 -4060 -12615
rect -4094 -12649 -4060 -12625
rect -4094 -12693 -4060 -12687
rect -4094 -12721 -4060 -12693
rect -4094 -12761 -4060 -12759
rect -4094 -12793 -4060 -12761
rect -4094 -12863 -4060 -12831
rect -4094 -12865 -4060 -12863
rect -4094 -12931 -4060 -12903
rect -4094 -12937 -4060 -12931
rect -4094 -12999 -4060 -12975
rect -4094 -13009 -4060 -12999
rect -4094 -13067 -4060 -13047
rect -4094 -13081 -4060 -13067
rect -3076 -12557 -3042 -12543
rect -3076 -12577 -3042 -12557
rect -3076 -12625 -3042 -12615
rect -3076 -12649 -3042 -12625
rect -3076 -12693 -3042 -12687
rect -3076 -12721 -3042 -12693
rect -3076 -12761 -3042 -12759
rect -3076 -12793 -3042 -12761
rect -3076 -12863 -3042 -12831
rect -3076 -12865 -3042 -12863
rect -3076 -12931 -3042 -12903
rect -3076 -12937 -3042 -12931
rect -3076 -12999 -3042 -12975
rect -3076 -13009 -3042 -12999
rect -3076 -13067 -3042 -13047
rect -3076 -13081 -3042 -13067
rect -2058 -12557 -2024 -12543
rect -2058 -12577 -2024 -12557
rect -2058 -12625 -2024 -12615
rect -2058 -12649 -2024 -12625
rect -2058 -12693 -2024 -12687
rect -2058 -12721 -2024 -12693
rect -2058 -12761 -2024 -12759
rect -2058 -12793 -2024 -12761
rect -2058 -12863 -2024 -12831
rect -2058 -12865 -2024 -12863
rect -2058 -12931 -2024 -12903
rect -2058 -12937 -2024 -12931
rect -2058 -12999 -2024 -12975
rect -2058 -13009 -2024 -12999
rect -2058 -13067 -2024 -13047
rect -2058 -13081 -2024 -13067
rect -1040 -12557 -1006 -12543
rect -1040 -12577 -1006 -12557
rect -1040 -12625 -1006 -12615
rect -1040 -12649 -1006 -12625
rect -1040 -12693 -1006 -12687
rect -1040 -12721 -1006 -12693
rect -1040 -12761 -1006 -12759
rect -1040 -12793 -1006 -12761
rect -1040 -12863 -1006 -12831
rect -1040 -12865 -1006 -12863
rect -1040 -12931 -1006 -12903
rect -1040 -12937 -1006 -12931
rect -1040 -12999 -1006 -12975
rect -1040 -13009 -1006 -12999
rect -1040 -13067 -1006 -13047
rect -1040 -13081 -1006 -13067
rect -22 -12557 12 -12543
rect -22 -12577 12 -12557
rect -22 -12625 12 -12615
rect -22 -12649 12 -12625
rect -22 -12693 12 -12687
rect -22 -12721 12 -12693
rect -22 -12761 12 -12759
rect -22 -12793 12 -12761
rect -22 -12863 12 -12831
rect -22 -12865 12 -12863
rect 24855 -12553 24889 -12523
rect 24855 -12557 24889 -12553
rect 24855 -12621 24889 -12595
rect 24855 -12629 24889 -12621
rect 24855 -12689 24889 -12667
rect 24855 -12701 24889 -12689
rect 24855 -12757 24889 -12739
rect 24855 -12773 24889 -12757
rect 24855 -12825 24889 -12811
rect 24855 -12845 24889 -12825
rect -22 -12931 12 -12903
rect 2911 -12914 2921 -12880
rect 2921 -12914 2945 -12880
rect 2983 -12914 2989 -12880
rect 2989 -12914 3017 -12880
rect 3055 -12914 3057 -12880
rect 3057 -12914 3089 -12880
rect 3127 -12914 3159 -12880
rect 3159 -12914 3161 -12880
rect 3199 -12914 3227 -12880
rect 3227 -12914 3233 -12880
rect 3271 -12914 3295 -12880
rect 3295 -12914 3305 -12880
rect 3929 -12914 3939 -12880
rect 3939 -12914 3963 -12880
rect 4001 -12914 4007 -12880
rect 4007 -12914 4035 -12880
rect 4073 -12914 4075 -12880
rect 4075 -12914 4107 -12880
rect 4145 -12914 4177 -12880
rect 4177 -12914 4179 -12880
rect 4217 -12914 4245 -12880
rect 4245 -12914 4251 -12880
rect 4289 -12914 4313 -12880
rect 4313 -12914 4323 -12880
rect 4947 -12914 4957 -12880
rect 4957 -12914 4981 -12880
rect 5019 -12914 5025 -12880
rect 5025 -12914 5053 -12880
rect 5091 -12914 5093 -12880
rect 5093 -12914 5125 -12880
rect 5163 -12914 5195 -12880
rect 5195 -12914 5197 -12880
rect 5235 -12914 5263 -12880
rect 5263 -12914 5269 -12880
rect 5307 -12914 5331 -12880
rect 5331 -12914 5341 -12880
rect 5965 -12914 5975 -12880
rect 5975 -12914 5999 -12880
rect 6037 -12914 6043 -12880
rect 6043 -12914 6071 -12880
rect 6109 -12914 6111 -12880
rect 6111 -12914 6143 -12880
rect 6181 -12914 6213 -12880
rect 6213 -12914 6215 -12880
rect 6253 -12914 6281 -12880
rect 6281 -12914 6287 -12880
rect 6325 -12914 6349 -12880
rect 6349 -12914 6359 -12880
rect 6983 -12914 6993 -12880
rect 6993 -12914 7017 -12880
rect 7055 -12914 7061 -12880
rect 7061 -12914 7089 -12880
rect 7127 -12914 7129 -12880
rect 7129 -12914 7161 -12880
rect 7199 -12914 7231 -12880
rect 7231 -12914 7233 -12880
rect 7271 -12914 7299 -12880
rect 7299 -12914 7305 -12880
rect 7343 -12914 7367 -12880
rect 7367 -12914 7377 -12880
rect 8001 -12914 8011 -12880
rect 8011 -12914 8035 -12880
rect 8073 -12914 8079 -12880
rect 8079 -12914 8107 -12880
rect 8145 -12914 8147 -12880
rect 8147 -12914 8179 -12880
rect 8217 -12914 8249 -12880
rect 8249 -12914 8251 -12880
rect 8289 -12914 8317 -12880
rect 8317 -12914 8323 -12880
rect 8361 -12914 8385 -12880
rect 8385 -12914 8395 -12880
rect 9019 -12914 9029 -12880
rect 9029 -12914 9053 -12880
rect 9091 -12914 9097 -12880
rect 9097 -12914 9125 -12880
rect 9163 -12914 9165 -12880
rect 9165 -12914 9197 -12880
rect 9235 -12914 9267 -12880
rect 9267 -12914 9269 -12880
rect 9307 -12914 9335 -12880
rect 9335 -12914 9341 -12880
rect 9379 -12914 9403 -12880
rect 9403 -12914 9413 -12880
rect 10037 -12914 10047 -12880
rect 10047 -12914 10071 -12880
rect 10109 -12914 10115 -12880
rect 10115 -12914 10143 -12880
rect 10181 -12914 10183 -12880
rect 10183 -12914 10215 -12880
rect 10253 -12914 10285 -12880
rect 10285 -12914 10287 -12880
rect 10325 -12914 10353 -12880
rect 10353 -12914 10359 -12880
rect 10397 -12914 10421 -12880
rect 10421 -12914 10431 -12880
rect 11055 -12914 11065 -12880
rect 11065 -12914 11089 -12880
rect 11127 -12914 11133 -12880
rect 11133 -12914 11161 -12880
rect 11199 -12914 11201 -12880
rect 11201 -12914 11233 -12880
rect 11271 -12914 11303 -12880
rect 11303 -12914 11305 -12880
rect 11343 -12914 11371 -12880
rect 11371 -12914 11377 -12880
rect 11415 -12914 11439 -12880
rect 11439 -12914 11449 -12880
rect 12073 -12914 12083 -12880
rect 12083 -12914 12107 -12880
rect 12145 -12914 12151 -12880
rect 12151 -12914 12179 -12880
rect 12217 -12914 12219 -12880
rect 12219 -12914 12251 -12880
rect 12289 -12914 12321 -12880
rect 12321 -12914 12323 -12880
rect 12361 -12914 12389 -12880
rect 12389 -12914 12395 -12880
rect 12433 -12914 12457 -12880
rect 12457 -12914 12467 -12880
rect 13091 -12914 13101 -12880
rect 13101 -12914 13125 -12880
rect 13163 -12914 13169 -12880
rect 13169 -12914 13197 -12880
rect 13235 -12914 13237 -12880
rect 13237 -12914 13269 -12880
rect 13307 -12914 13339 -12880
rect 13339 -12914 13341 -12880
rect 13379 -12914 13407 -12880
rect 13407 -12914 13413 -12880
rect 13451 -12914 13475 -12880
rect 13475 -12914 13485 -12880
rect 14109 -12914 14119 -12880
rect 14119 -12914 14143 -12880
rect 14181 -12914 14187 -12880
rect 14187 -12914 14215 -12880
rect 14253 -12914 14255 -12880
rect 14255 -12914 14287 -12880
rect 14325 -12914 14357 -12880
rect 14357 -12914 14359 -12880
rect 14397 -12914 14425 -12880
rect 14425 -12914 14431 -12880
rect 14469 -12914 14493 -12880
rect 14493 -12914 14503 -12880
rect 15127 -12914 15137 -12880
rect 15137 -12914 15161 -12880
rect 15199 -12914 15205 -12880
rect 15205 -12914 15233 -12880
rect 15271 -12914 15273 -12880
rect 15273 -12914 15305 -12880
rect 15343 -12914 15375 -12880
rect 15375 -12914 15377 -12880
rect 15415 -12914 15443 -12880
rect 15443 -12914 15449 -12880
rect 15487 -12914 15511 -12880
rect 15511 -12914 15521 -12880
rect 16145 -12914 16155 -12880
rect 16155 -12914 16179 -12880
rect 16217 -12914 16223 -12880
rect 16223 -12914 16251 -12880
rect 16289 -12914 16291 -12880
rect 16291 -12914 16323 -12880
rect 16361 -12914 16393 -12880
rect 16393 -12914 16395 -12880
rect 16433 -12914 16461 -12880
rect 16461 -12914 16467 -12880
rect 16505 -12914 16529 -12880
rect 16529 -12914 16539 -12880
rect 17163 -12914 17173 -12880
rect 17173 -12914 17197 -12880
rect 17235 -12914 17241 -12880
rect 17241 -12914 17269 -12880
rect 17307 -12914 17309 -12880
rect 17309 -12914 17341 -12880
rect 17379 -12914 17411 -12880
rect 17411 -12914 17413 -12880
rect 17451 -12914 17479 -12880
rect 17479 -12914 17485 -12880
rect 17523 -12914 17547 -12880
rect 17547 -12914 17557 -12880
rect 18181 -12914 18191 -12880
rect 18191 -12914 18215 -12880
rect 18253 -12914 18259 -12880
rect 18259 -12914 18287 -12880
rect 18325 -12914 18327 -12880
rect 18327 -12914 18359 -12880
rect 18397 -12914 18429 -12880
rect 18429 -12914 18431 -12880
rect 18469 -12914 18497 -12880
rect 18497 -12914 18503 -12880
rect 18541 -12914 18565 -12880
rect 18565 -12914 18575 -12880
rect 19199 -12914 19209 -12880
rect 19209 -12914 19233 -12880
rect 19271 -12914 19277 -12880
rect 19277 -12914 19305 -12880
rect 19343 -12914 19345 -12880
rect 19345 -12914 19377 -12880
rect 19415 -12914 19447 -12880
rect 19447 -12914 19449 -12880
rect 19487 -12914 19515 -12880
rect 19515 -12914 19521 -12880
rect 19559 -12914 19583 -12880
rect 19583 -12914 19593 -12880
rect 20217 -12914 20227 -12880
rect 20227 -12914 20251 -12880
rect 20289 -12914 20295 -12880
rect 20295 -12914 20323 -12880
rect 20361 -12914 20363 -12880
rect 20363 -12914 20395 -12880
rect 20433 -12914 20465 -12880
rect 20465 -12914 20467 -12880
rect 20505 -12914 20533 -12880
rect 20533 -12914 20539 -12880
rect 20577 -12914 20601 -12880
rect 20601 -12914 20611 -12880
rect 21235 -12914 21245 -12880
rect 21245 -12914 21269 -12880
rect 21307 -12914 21313 -12880
rect 21313 -12914 21341 -12880
rect 21379 -12914 21381 -12880
rect 21381 -12914 21413 -12880
rect 21451 -12914 21483 -12880
rect 21483 -12914 21485 -12880
rect 21523 -12914 21551 -12880
rect 21551 -12914 21557 -12880
rect 21595 -12914 21619 -12880
rect 21619 -12914 21629 -12880
rect 22253 -12914 22263 -12880
rect 22263 -12914 22287 -12880
rect 22325 -12914 22331 -12880
rect 22331 -12914 22359 -12880
rect 22397 -12914 22399 -12880
rect 22399 -12914 22431 -12880
rect 22469 -12914 22501 -12880
rect 22501 -12914 22503 -12880
rect 22541 -12914 22569 -12880
rect 22569 -12914 22575 -12880
rect 22613 -12914 22637 -12880
rect 22637 -12914 22647 -12880
rect 24855 -12893 24889 -12883
rect 24855 -12917 24889 -12893
rect -22 -12937 12 -12931
rect -22 -12999 12 -12975
rect -22 -13009 12 -12999
rect -22 -13067 12 -13047
rect -22 -13081 12 -13067
rect 2582 -12997 2616 -12983
rect 2582 -13017 2616 -12997
rect 2582 -13065 2616 -13055
rect 2582 -13089 2616 -13065
rect 2582 -13133 2616 -13127
rect -12289 -13199 -12255 -13171
rect -12289 -13205 -12255 -13199
rect -8855 -13184 -8845 -13150
rect -8845 -13184 -8821 -13150
rect -8783 -13184 -8777 -13150
rect -8777 -13184 -8749 -13150
rect -8711 -13184 -8709 -13150
rect -8709 -13184 -8677 -13150
rect -8639 -13184 -8607 -13150
rect -8607 -13184 -8605 -13150
rect -8567 -13184 -8539 -13150
rect -8539 -13184 -8533 -13150
rect -8495 -13184 -8471 -13150
rect -8471 -13184 -8461 -13150
rect -7837 -13184 -7827 -13150
rect -7827 -13184 -7803 -13150
rect -7765 -13184 -7759 -13150
rect -7759 -13184 -7731 -13150
rect -7693 -13184 -7691 -13150
rect -7691 -13184 -7659 -13150
rect -7621 -13184 -7589 -13150
rect -7589 -13184 -7587 -13150
rect -7549 -13184 -7521 -13150
rect -7521 -13184 -7515 -13150
rect -7477 -13184 -7453 -13150
rect -7453 -13184 -7443 -13150
rect -6819 -13184 -6809 -13150
rect -6809 -13184 -6785 -13150
rect -6747 -13184 -6741 -13150
rect -6741 -13184 -6713 -13150
rect -6675 -13184 -6673 -13150
rect -6673 -13184 -6641 -13150
rect -6603 -13184 -6571 -13150
rect -6571 -13184 -6569 -13150
rect -6531 -13184 -6503 -13150
rect -6503 -13184 -6497 -13150
rect -6459 -13184 -6435 -13150
rect -6435 -13184 -6425 -13150
rect -5801 -13184 -5791 -13150
rect -5791 -13184 -5767 -13150
rect -5729 -13184 -5723 -13150
rect -5723 -13184 -5695 -13150
rect -5657 -13184 -5655 -13150
rect -5655 -13184 -5623 -13150
rect -5585 -13184 -5553 -13150
rect -5553 -13184 -5551 -13150
rect -5513 -13184 -5485 -13150
rect -5485 -13184 -5479 -13150
rect -5441 -13184 -5417 -13150
rect -5417 -13184 -5407 -13150
rect -4783 -13184 -4773 -13150
rect -4773 -13184 -4749 -13150
rect -4711 -13184 -4705 -13150
rect -4705 -13184 -4677 -13150
rect -4639 -13184 -4637 -13150
rect -4637 -13184 -4605 -13150
rect -4567 -13184 -4535 -13150
rect -4535 -13184 -4533 -13150
rect -4495 -13184 -4467 -13150
rect -4467 -13184 -4461 -13150
rect -4423 -13184 -4399 -13150
rect -4399 -13184 -4389 -13150
rect -3765 -13184 -3755 -13150
rect -3755 -13184 -3731 -13150
rect -3693 -13184 -3687 -13150
rect -3687 -13184 -3659 -13150
rect -3621 -13184 -3619 -13150
rect -3619 -13184 -3587 -13150
rect -3549 -13184 -3517 -13150
rect -3517 -13184 -3515 -13150
rect -3477 -13184 -3449 -13150
rect -3449 -13184 -3443 -13150
rect -3405 -13184 -3381 -13150
rect -3381 -13184 -3371 -13150
rect -2747 -13184 -2737 -13150
rect -2737 -13184 -2713 -13150
rect -2675 -13184 -2669 -13150
rect -2669 -13184 -2641 -13150
rect -2603 -13184 -2601 -13150
rect -2601 -13184 -2569 -13150
rect -2531 -13184 -2499 -13150
rect -2499 -13184 -2497 -13150
rect -2459 -13184 -2431 -13150
rect -2431 -13184 -2425 -13150
rect -2387 -13184 -2363 -13150
rect -2363 -13184 -2353 -13150
rect -1729 -13184 -1719 -13150
rect -1719 -13184 -1695 -13150
rect -1657 -13184 -1651 -13150
rect -1651 -13184 -1623 -13150
rect -1585 -13184 -1583 -13150
rect -1583 -13184 -1551 -13150
rect -1513 -13184 -1481 -13150
rect -1481 -13184 -1479 -13150
rect -1441 -13184 -1413 -13150
rect -1413 -13184 -1407 -13150
rect -1369 -13184 -1345 -13150
rect -1345 -13184 -1335 -13150
rect -711 -13184 -701 -13150
rect -701 -13184 -677 -13150
rect -639 -13184 -633 -13150
rect -633 -13184 -605 -13150
rect -567 -13184 -565 -13150
rect -565 -13184 -533 -13150
rect -495 -13184 -463 -13150
rect -463 -13184 -461 -13150
rect -423 -13184 -395 -13150
rect -395 -13184 -389 -13150
rect -351 -13184 -327 -13150
rect -327 -13184 -317 -13150
rect 2582 -13161 2616 -13133
rect -12289 -13267 -12255 -13243
rect -12289 -13277 -12255 -13267
rect 2582 -13201 2616 -13199
rect 2582 -13233 2616 -13201
rect -8855 -13292 -8845 -13258
rect -8845 -13292 -8821 -13258
rect -8783 -13292 -8777 -13258
rect -8777 -13292 -8749 -13258
rect -8711 -13292 -8709 -13258
rect -8709 -13292 -8677 -13258
rect -8639 -13292 -8607 -13258
rect -8607 -13292 -8605 -13258
rect -8567 -13292 -8539 -13258
rect -8539 -13292 -8533 -13258
rect -8495 -13292 -8471 -13258
rect -8471 -13292 -8461 -13258
rect -7837 -13292 -7827 -13258
rect -7827 -13292 -7803 -13258
rect -7765 -13292 -7759 -13258
rect -7759 -13292 -7731 -13258
rect -7693 -13292 -7691 -13258
rect -7691 -13292 -7659 -13258
rect -7621 -13292 -7589 -13258
rect -7589 -13292 -7587 -13258
rect -7549 -13292 -7521 -13258
rect -7521 -13292 -7515 -13258
rect -7477 -13292 -7453 -13258
rect -7453 -13292 -7443 -13258
rect -6819 -13292 -6809 -13258
rect -6809 -13292 -6785 -13258
rect -6747 -13292 -6741 -13258
rect -6741 -13292 -6713 -13258
rect -6675 -13292 -6673 -13258
rect -6673 -13292 -6641 -13258
rect -6603 -13292 -6571 -13258
rect -6571 -13292 -6569 -13258
rect -6531 -13292 -6503 -13258
rect -6503 -13292 -6497 -13258
rect -6459 -13292 -6435 -13258
rect -6435 -13292 -6425 -13258
rect -5801 -13292 -5791 -13258
rect -5791 -13292 -5767 -13258
rect -5729 -13292 -5723 -13258
rect -5723 -13292 -5695 -13258
rect -5657 -13292 -5655 -13258
rect -5655 -13292 -5623 -13258
rect -5585 -13292 -5553 -13258
rect -5553 -13292 -5551 -13258
rect -5513 -13292 -5485 -13258
rect -5485 -13292 -5479 -13258
rect -5441 -13292 -5417 -13258
rect -5417 -13292 -5407 -13258
rect -4783 -13292 -4773 -13258
rect -4773 -13292 -4749 -13258
rect -4711 -13292 -4705 -13258
rect -4705 -13292 -4677 -13258
rect -4639 -13292 -4637 -13258
rect -4637 -13292 -4605 -13258
rect -4567 -13292 -4535 -13258
rect -4535 -13292 -4533 -13258
rect -4495 -13292 -4467 -13258
rect -4467 -13292 -4461 -13258
rect -4423 -13292 -4399 -13258
rect -4399 -13292 -4389 -13258
rect -3765 -13292 -3755 -13258
rect -3755 -13292 -3731 -13258
rect -3693 -13292 -3687 -13258
rect -3687 -13292 -3659 -13258
rect -3621 -13292 -3619 -13258
rect -3619 -13292 -3587 -13258
rect -3549 -13292 -3517 -13258
rect -3517 -13292 -3515 -13258
rect -3477 -13292 -3449 -13258
rect -3449 -13292 -3443 -13258
rect -3405 -13292 -3381 -13258
rect -3381 -13292 -3371 -13258
rect -2747 -13292 -2737 -13258
rect -2737 -13292 -2713 -13258
rect -2675 -13292 -2669 -13258
rect -2669 -13292 -2641 -13258
rect -2603 -13292 -2601 -13258
rect -2601 -13292 -2569 -13258
rect -2531 -13292 -2499 -13258
rect -2499 -13292 -2497 -13258
rect -2459 -13292 -2431 -13258
rect -2431 -13292 -2425 -13258
rect -2387 -13292 -2363 -13258
rect -2363 -13292 -2353 -13258
rect -1729 -13292 -1719 -13258
rect -1719 -13292 -1695 -13258
rect -1657 -13292 -1651 -13258
rect -1651 -13292 -1623 -13258
rect -1585 -13292 -1583 -13258
rect -1583 -13292 -1551 -13258
rect -1513 -13292 -1481 -13258
rect -1481 -13292 -1479 -13258
rect -1441 -13292 -1413 -13258
rect -1413 -13292 -1407 -13258
rect -1369 -13292 -1345 -13258
rect -1345 -13292 -1335 -13258
rect -711 -13292 -701 -13258
rect -701 -13292 -677 -13258
rect -639 -13292 -633 -13258
rect -633 -13292 -605 -13258
rect -567 -13292 -565 -13258
rect -565 -13292 -533 -13258
rect -495 -13292 -463 -13258
rect -463 -13292 -461 -13258
rect -423 -13292 -395 -13258
rect -395 -13292 -389 -13258
rect -351 -13292 -327 -13258
rect -327 -13292 -317 -13258
rect -12289 -13335 -12255 -13315
rect -12289 -13349 -12255 -13335
rect 2582 -13303 2616 -13271
rect 2582 -13305 2616 -13303
rect -12289 -13403 -12255 -13387
rect -12289 -13421 -12255 -13403
rect -12289 -13471 -12255 -13459
rect -12289 -13493 -12255 -13471
rect -12289 -13539 -12255 -13531
rect -12289 -13565 -12255 -13539
rect -12289 -13607 -12255 -13603
rect -12289 -13637 -12255 -13607
rect -12289 -13709 -12255 -13675
rect -12289 -13777 -12255 -13747
rect -12289 -13781 -12255 -13777
rect -12289 -13845 -12255 -13819
rect -12289 -13853 -12255 -13845
rect -12289 -13913 -12255 -13891
rect -12289 -13925 -12255 -13913
rect -9184 -13375 -9150 -13361
rect -9184 -13395 -9150 -13375
rect -9184 -13443 -9150 -13433
rect -9184 -13467 -9150 -13443
rect -9184 -13511 -9150 -13505
rect -9184 -13539 -9150 -13511
rect -9184 -13579 -9150 -13577
rect -9184 -13611 -9150 -13579
rect -9184 -13681 -9150 -13649
rect -9184 -13683 -9150 -13681
rect -9184 -13749 -9150 -13721
rect -9184 -13755 -9150 -13749
rect -9184 -13817 -9150 -13793
rect -9184 -13827 -9150 -13817
rect -9184 -13885 -9150 -13865
rect -9184 -13899 -9150 -13885
rect -8166 -13375 -8132 -13361
rect -8166 -13395 -8132 -13375
rect -8166 -13443 -8132 -13433
rect -8166 -13467 -8132 -13443
rect -8166 -13511 -8132 -13505
rect -8166 -13539 -8132 -13511
rect -8166 -13579 -8132 -13577
rect -8166 -13611 -8132 -13579
rect -8166 -13681 -8132 -13649
rect -8166 -13683 -8132 -13681
rect -8166 -13749 -8132 -13721
rect -8166 -13755 -8132 -13749
rect -8166 -13817 -8132 -13793
rect -8166 -13827 -8132 -13817
rect -8166 -13885 -8132 -13865
rect -8166 -13899 -8132 -13885
rect -7148 -13375 -7114 -13361
rect -7148 -13395 -7114 -13375
rect -7148 -13443 -7114 -13433
rect -7148 -13467 -7114 -13443
rect -7148 -13511 -7114 -13505
rect -7148 -13539 -7114 -13511
rect -7148 -13579 -7114 -13577
rect -7148 -13611 -7114 -13579
rect -7148 -13681 -7114 -13649
rect -7148 -13683 -7114 -13681
rect -7148 -13749 -7114 -13721
rect -7148 -13755 -7114 -13749
rect -7148 -13817 -7114 -13793
rect -7148 -13827 -7114 -13817
rect -7148 -13885 -7114 -13865
rect -7148 -13899 -7114 -13885
rect -6130 -13375 -6096 -13361
rect -6130 -13395 -6096 -13375
rect -6130 -13443 -6096 -13433
rect -6130 -13467 -6096 -13443
rect -6130 -13511 -6096 -13505
rect -6130 -13539 -6096 -13511
rect -6130 -13579 -6096 -13577
rect -6130 -13611 -6096 -13579
rect -6130 -13681 -6096 -13649
rect -6130 -13683 -6096 -13681
rect -6130 -13749 -6096 -13721
rect -6130 -13755 -6096 -13749
rect -6130 -13817 -6096 -13793
rect -6130 -13827 -6096 -13817
rect -6130 -13885 -6096 -13865
rect -6130 -13899 -6096 -13885
rect -5112 -13375 -5078 -13361
rect -5112 -13395 -5078 -13375
rect -5112 -13443 -5078 -13433
rect -5112 -13467 -5078 -13443
rect -5112 -13511 -5078 -13505
rect -5112 -13539 -5078 -13511
rect -5112 -13579 -5078 -13577
rect -5112 -13611 -5078 -13579
rect -5112 -13681 -5078 -13649
rect -5112 -13683 -5078 -13681
rect -5112 -13749 -5078 -13721
rect -5112 -13755 -5078 -13749
rect -5112 -13817 -5078 -13793
rect -5112 -13827 -5078 -13817
rect -5112 -13885 -5078 -13865
rect -5112 -13899 -5078 -13885
rect -4094 -13375 -4060 -13361
rect -4094 -13395 -4060 -13375
rect -4094 -13443 -4060 -13433
rect -4094 -13467 -4060 -13443
rect -4094 -13511 -4060 -13505
rect -4094 -13539 -4060 -13511
rect -4094 -13579 -4060 -13577
rect -4094 -13611 -4060 -13579
rect -4094 -13681 -4060 -13649
rect -4094 -13683 -4060 -13681
rect -4094 -13749 -4060 -13721
rect -4094 -13755 -4060 -13749
rect -4094 -13817 -4060 -13793
rect -4094 -13827 -4060 -13817
rect -4094 -13885 -4060 -13865
rect -4094 -13899 -4060 -13885
rect -3076 -13375 -3042 -13361
rect -3076 -13395 -3042 -13375
rect -3076 -13443 -3042 -13433
rect -3076 -13467 -3042 -13443
rect -3076 -13511 -3042 -13505
rect -3076 -13539 -3042 -13511
rect -3076 -13579 -3042 -13577
rect -3076 -13611 -3042 -13579
rect -3076 -13681 -3042 -13649
rect -3076 -13683 -3042 -13681
rect -3076 -13749 -3042 -13721
rect -3076 -13755 -3042 -13749
rect -3076 -13817 -3042 -13793
rect -3076 -13827 -3042 -13817
rect -3076 -13885 -3042 -13865
rect -3076 -13899 -3042 -13885
rect -2058 -13375 -2024 -13361
rect -2058 -13395 -2024 -13375
rect -2058 -13443 -2024 -13433
rect -2058 -13467 -2024 -13443
rect -2058 -13511 -2024 -13505
rect -2058 -13539 -2024 -13511
rect -2058 -13579 -2024 -13577
rect -2058 -13611 -2024 -13579
rect -2058 -13681 -2024 -13649
rect -2058 -13683 -2024 -13681
rect -2058 -13749 -2024 -13721
rect -2058 -13755 -2024 -13749
rect -2058 -13817 -2024 -13793
rect -2058 -13827 -2024 -13817
rect -2058 -13885 -2024 -13865
rect -2058 -13899 -2024 -13885
rect -1040 -13375 -1006 -13361
rect -1040 -13395 -1006 -13375
rect -1040 -13443 -1006 -13433
rect -1040 -13467 -1006 -13443
rect -1040 -13511 -1006 -13505
rect -1040 -13539 -1006 -13511
rect -1040 -13579 -1006 -13577
rect -1040 -13611 -1006 -13579
rect -1040 -13681 -1006 -13649
rect -1040 -13683 -1006 -13681
rect -1040 -13749 -1006 -13721
rect -1040 -13755 -1006 -13749
rect -1040 -13817 -1006 -13793
rect -1040 -13827 -1006 -13817
rect -1040 -13885 -1006 -13865
rect -1040 -13899 -1006 -13885
rect -22 -13375 12 -13361
rect -22 -13395 12 -13375
rect -22 -13443 12 -13433
rect -22 -13467 12 -13443
rect -22 -13511 12 -13505
rect -22 -13539 12 -13511
rect 2582 -13371 2616 -13343
rect 2582 -13377 2616 -13371
rect 2582 -13439 2616 -13415
rect 2582 -13449 2616 -13439
rect 2582 -13507 2616 -13487
rect 2582 -13521 2616 -13507
rect 3600 -12997 3634 -12983
rect 3600 -13017 3634 -12997
rect 3600 -13065 3634 -13055
rect 3600 -13089 3634 -13065
rect 3600 -13133 3634 -13127
rect 3600 -13161 3634 -13133
rect 3600 -13201 3634 -13199
rect 3600 -13233 3634 -13201
rect 3600 -13303 3634 -13271
rect 3600 -13305 3634 -13303
rect 3600 -13371 3634 -13343
rect 3600 -13377 3634 -13371
rect 3600 -13439 3634 -13415
rect 3600 -13449 3634 -13439
rect 3600 -13507 3634 -13487
rect 3600 -13521 3634 -13507
rect 4618 -12997 4652 -12983
rect 4618 -13017 4652 -12997
rect 4618 -13065 4652 -13055
rect 4618 -13089 4652 -13065
rect 4618 -13133 4652 -13127
rect 4618 -13161 4652 -13133
rect 4618 -13201 4652 -13199
rect 4618 -13233 4652 -13201
rect 4618 -13303 4652 -13271
rect 4618 -13305 4652 -13303
rect 4618 -13371 4652 -13343
rect 4618 -13377 4652 -13371
rect 4618 -13439 4652 -13415
rect 4618 -13449 4652 -13439
rect 4618 -13507 4652 -13487
rect 4618 -13521 4652 -13507
rect 5636 -12997 5670 -12983
rect 5636 -13017 5670 -12997
rect 5636 -13065 5670 -13055
rect 5636 -13089 5670 -13065
rect 5636 -13133 5670 -13127
rect 5636 -13161 5670 -13133
rect 5636 -13201 5670 -13199
rect 5636 -13233 5670 -13201
rect 5636 -13303 5670 -13271
rect 5636 -13305 5670 -13303
rect 5636 -13371 5670 -13343
rect 5636 -13377 5670 -13371
rect 5636 -13439 5670 -13415
rect 5636 -13449 5670 -13439
rect 5636 -13507 5670 -13487
rect 5636 -13521 5670 -13507
rect 6654 -12997 6688 -12983
rect 6654 -13017 6688 -12997
rect 6654 -13065 6688 -13055
rect 6654 -13089 6688 -13065
rect 6654 -13133 6688 -13127
rect 6654 -13161 6688 -13133
rect 6654 -13201 6688 -13199
rect 6654 -13233 6688 -13201
rect 6654 -13303 6688 -13271
rect 6654 -13305 6688 -13303
rect 6654 -13371 6688 -13343
rect 6654 -13377 6688 -13371
rect 6654 -13439 6688 -13415
rect 6654 -13449 6688 -13439
rect 6654 -13507 6688 -13487
rect 6654 -13521 6688 -13507
rect 7672 -12997 7706 -12983
rect 7672 -13017 7706 -12997
rect 7672 -13065 7706 -13055
rect 7672 -13089 7706 -13065
rect 7672 -13133 7706 -13127
rect 7672 -13161 7706 -13133
rect 7672 -13201 7706 -13199
rect 7672 -13233 7706 -13201
rect 7672 -13303 7706 -13271
rect 7672 -13305 7706 -13303
rect 7672 -13371 7706 -13343
rect 7672 -13377 7706 -13371
rect 7672 -13439 7706 -13415
rect 7672 -13449 7706 -13439
rect 7672 -13507 7706 -13487
rect 7672 -13521 7706 -13507
rect 8690 -12997 8724 -12983
rect 8690 -13017 8724 -12997
rect 8690 -13065 8724 -13055
rect 8690 -13089 8724 -13065
rect 8690 -13133 8724 -13127
rect 8690 -13161 8724 -13133
rect 8690 -13201 8724 -13199
rect 8690 -13233 8724 -13201
rect 8690 -13303 8724 -13271
rect 8690 -13305 8724 -13303
rect 8690 -13371 8724 -13343
rect 8690 -13377 8724 -13371
rect 8690 -13439 8724 -13415
rect 8690 -13449 8724 -13439
rect 8690 -13507 8724 -13487
rect 8690 -13521 8724 -13507
rect 9708 -12997 9742 -12983
rect 9708 -13017 9742 -12997
rect 9708 -13065 9742 -13055
rect 9708 -13089 9742 -13065
rect 9708 -13133 9742 -13127
rect 9708 -13161 9742 -13133
rect 9708 -13201 9742 -13199
rect 9708 -13233 9742 -13201
rect 9708 -13303 9742 -13271
rect 9708 -13305 9742 -13303
rect 9708 -13371 9742 -13343
rect 9708 -13377 9742 -13371
rect 9708 -13439 9742 -13415
rect 9708 -13449 9742 -13439
rect 9708 -13507 9742 -13487
rect 9708 -13521 9742 -13507
rect 10726 -12997 10760 -12983
rect 10726 -13017 10760 -12997
rect 10726 -13065 10760 -13055
rect 10726 -13089 10760 -13065
rect 10726 -13133 10760 -13127
rect 10726 -13161 10760 -13133
rect 10726 -13201 10760 -13199
rect 10726 -13233 10760 -13201
rect 10726 -13303 10760 -13271
rect 10726 -13305 10760 -13303
rect 10726 -13371 10760 -13343
rect 10726 -13377 10760 -13371
rect 10726 -13439 10760 -13415
rect 10726 -13449 10760 -13439
rect 10726 -13507 10760 -13487
rect 10726 -13521 10760 -13507
rect 11744 -12997 11778 -12983
rect 11744 -13017 11778 -12997
rect 11744 -13065 11778 -13055
rect 11744 -13089 11778 -13065
rect 11744 -13133 11778 -13127
rect 11744 -13161 11778 -13133
rect 11744 -13201 11778 -13199
rect 11744 -13233 11778 -13201
rect 11744 -13303 11778 -13271
rect 11744 -13305 11778 -13303
rect 11744 -13371 11778 -13343
rect 11744 -13377 11778 -13371
rect 11744 -13439 11778 -13415
rect 11744 -13449 11778 -13439
rect 11744 -13507 11778 -13487
rect 11744 -13521 11778 -13507
rect 12762 -12997 12796 -12983
rect 12762 -13017 12796 -12997
rect 12762 -13065 12796 -13055
rect 12762 -13089 12796 -13065
rect 12762 -13133 12796 -13127
rect 12762 -13161 12796 -13133
rect 12762 -13201 12796 -13199
rect 12762 -13233 12796 -13201
rect 12762 -13303 12796 -13271
rect 12762 -13305 12796 -13303
rect 12762 -13371 12796 -13343
rect 12762 -13377 12796 -13371
rect 12762 -13439 12796 -13415
rect 12762 -13449 12796 -13439
rect 12762 -13507 12796 -13487
rect 12762 -13521 12796 -13507
rect 13780 -12997 13814 -12983
rect 13780 -13017 13814 -12997
rect 13780 -13065 13814 -13055
rect 13780 -13089 13814 -13065
rect 13780 -13133 13814 -13127
rect 13780 -13161 13814 -13133
rect 13780 -13201 13814 -13199
rect 13780 -13233 13814 -13201
rect 13780 -13303 13814 -13271
rect 13780 -13305 13814 -13303
rect 13780 -13371 13814 -13343
rect 13780 -13377 13814 -13371
rect 13780 -13439 13814 -13415
rect 13780 -13449 13814 -13439
rect 13780 -13507 13814 -13487
rect 13780 -13521 13814 -13507
rect 14798 -12997 14832 -12983
rect 14798 -13017 14832 -12997
rect 14798 -13065 14832 -13055
rect 14798 -13089 14832 -13065
rect 14798 -13133 14832 -13127
rect 14798 -13161 14832 -13133
rect 14798 -13201 14832 -13199
rect 14798 -13233 14832 -13201
rect 14798 -13303 14832 -13271
rect 14798 -13305 14832 -13303
rect 14798 -13371 14832 -13343
rect 14798 -13377 14832 -13371
rect 14798 -13439 14832 -13415
rect 14798 -13449 14832 -13439
rect 14798 -13507 14832 -13487
rect 14798 -13521 14832 -13507
rect 15816 -12997 15850 -12983
rect 15816 -13017 15850 -12997
rect 15816 -13065 15850 -13055
rect 15816 -13089 15850 -13065
rect 15816 -13133 15850 -13127
rect 15816 -13161 15850 -13133
rect 15816 -13201 15850 -13199
rect 15816 -13233 15850 -13201
rect 15816 -13303 15850 -13271
rect 15816 -13305 15850 -13303
rect 15816 -13371 15850 -13343
rect 15816 -13377 15850 -13371
rect 15816 -13439 15850 -13415
rect 15816 -13449 15850 -13439
rect 15816 -13507 15850 -13487
rect 15816 -13521 15850 -13507
rect 16834 -12997 16868 -12983
rect 16834 -13017 16868 -12997
rect 16834 -13065 16868 -13055
rect 16834 -13089 16868 -13065
rect 16834 -13133 16868 -13127
rect 16834 -13161 16868 -13133
rect 16834 -13201 16868 -13199
rect 16834 -13233 16868 -13201
rect 16834 -13303 16868 -13271
rect 16834 -13305 16868 -13303
rect 16834 -13371 16868 -13343
rect 16834 -13377 16868 -13371
rect 16834 -13439 16868 -13415
rect 16834 -13449 16868 -13439
rect 16834 -13507 16868 -13487
rect 16834 -13521 16868 -13507
rect 17852 -12997 17886 -12983
rect 17852 -13017 17886 -12997
rect 17852 -13065 17886 -13055
rect 17852 -13089 17886 -13065
rect 17852 -13133 17886 -13127
rect 17852 -13161 17886 -13133
rect 17852 -13201 17886 -13199
rect 17852 -13233 17886 -13201
rect 17852 -13303 17886 -13271
rect 17852 -13305 17886 -13303
rect 17852 -13371 17886 -13343
rect 17852 -13377 17886 -13371
rect 17852 -13439 17886 -13415
rect 17852 -13449 17886 -13439
rect 17852 -13507 17886 -13487
rect 17852 -13521 17886 -13507
rect 18870 -12997 18904 -12983
rect 18870 -13017 18904 -12997
rect 18870 -13065 18904 -13055
rect 18870 -13089 18904 -13065
rect 18870 -13133 18904 -13127
rect 18870 -13161 18904 -13133
rect 18870 -13201 18904 -13199
rect 18870 -13233 18904 -13201
rect 18870 -13303 18904 -13271
rect 18870 -13305 18904 -13303
rect 18870 -13371 18904 -13343
rect 18870 -13377 18904 -13371
rect 18870 -13439 18904 -13415
rect 18870 -13449 18904 -13439
rect 18870 -13507 18904 -13487
rect 18870 -13521 18904 -13507
rect 19888 -12997 19922 -12983
rect 19888 -13017 19922 -12997
rect 19888 -13065 19922 -13055
rect 19888 -13089 19922 -13065
rect 19888 -13133 19922 -13127
rect 19888 -13161 19922 -13133
rect 19888 -13201 19922 -13199
rect 19888 -13233 19922 -13201
rect 19888 -13303 19922 -13271
rect 19888 -13305 19922 -13303
rect 19888 -13371 19922 -13343
rect 19888 -13377 19922 -13371
rect 19888 -13439 19922 -13415
rect 19888 -13449 19922 -13439
rect 19888 -13507 19922 -13487
rect 19888 -13521 19922 -13507
rect 20906 -12997 20940 -12983
rect 20906 -13017 20940 -12997
rect 20906 -13065 20940 -13055
rect 20906 -13089 20940 -13065
rect 20906 -13133 20940 -13127
rect 20906 -13161 20940 -13133
rect 20906 -13201 20940 -13199
rect 20906 -13233 20940 -13201
rect 20906 -13303 20940 -13271
rect 20906 -13305 20940 -13303
rect 20906 -13371 20940 -13343
rect 20906 -13377 20940 -13371
rect 20906 -13439 20940 -13415
rect 20906 -13449 20940 -13439
rect 20906 -13507 20940 -13487
rect 20906 -13521 20940 -13507
rect 21924 -12997 21958 -12983
rect 21924 -13017 21958 -12997
rect 21924 -13065 21958 -13055
rect 21924 -13089 21958 -13065
rect 21924 -13133 21958 -13127
rect 21924 -13161 21958 -13133
rect 21924 -13201 21958 -13199
rect 21924 -13233 21958 -13201
rect 21924 -13303 21958 -13271
rect 21924 -13305 21958 -13303
rect 21924 -13371 21958 -13343
rect 21924 -13377 21958 -13371
rect 21924 -13439 21958 -13415
rect 21924 -13449 21958 -13439
rect 21924 -13507 21958 -13487
rect 21924 -13521 21958 -13507
rect 22942 -12997 22976 -12983
rect 22942 -13017 22976 -12997
rect 22942 -13065 22976 -13055
rect 22942 -13089 22976 -13065
rect 22942 -13133 22976 -13127
rect 22942 -13161 22976 -13133
rect 22942 -13201 22976 -13199
rect 22942 -13233 22976 -13201
rect 22942 -13303 22976 -13271
rect 22942 -13305 22976 -13303
rect 22942 -13371 22976 -13343
rect 22942 -13377 22976 -13371
rect 22942 -13439 22976 -13415
rect 22942 -13449 22976 -13439
rect 22942 -13507 22976 -13487
rect 22942 -13521 22976 -13507
rect 24855 -12961 24889 -12955
rect 24855 -12989 24889 -12961
rect 24855 -13029 24889 -13027
rect 24855 -13061 24889 -13029
rect 24855 -13131 24889 -13099
rect 24855 -13133 24889 -13131
rect 24855 -13199 24889 -13171
rect 24855 -13205 24889 -13199
rect 24855 -13267 24889 -13243
rect 24855 -13277 24889 -13267
rect 24855 -13335 24889 -13315
rect 24855 -13349 24889 -13335
rect 24855 -13403 24889 -13387
rect 24855 -13421 24889 -13403
rect 24855 -13471 24889 -13459
rect 24855 -13493 24889 -13471
rect -22 -13579 12 -13577
rect -22 -13611 12 -13579
rect 24855 -13539 24889 -13531
rect 24855 -13565 24889 -13539
rect 2911 -13624 2921 -13590
rect 2921 -13624 2945 -13590
rect 2983 -13624 2989 -13590
rect 2989 -13624 3017 -13590
rect 3055 -13624 3057 -13590
rect 3057 -13624 3089 -13590
rect 3127 -13624 3159 -13590
rect 3159 -13624 3161 -13590
rect 3199 -13624 3227 -13590
rect 3227 -13624 3233 -13590
rect 3271 -13624 3295 -13590
rect 3295 -13624 3305 -13590
rect 3929 -13624 3939 -13590
rect 3939 -13624 3963 -13590
rect 4001 -13624 4007 -13590
rect 4007 -13624 4035 -13590
rect 4073 -13624 4075 -13590
rect 4075 -13624 4107 -13590
rect 4145 -13624 4177 -13590
rect 4177 -13624 4179 -13590
rect 4217 -13624 4245 -13590
rect 4245 -13624 4251 -13590
rect 4289 -13624 4313 -13590
rect 4313 -13624 4323 -13590
rect 4947 -13624 4957 -13590
rect 4957 -13624 4981 -13590
rect 5019 -13624 5025 -13590
rect 5025 -13624 5053 -13590
rect 5091 -13624 5093 -13590
rect 5093 -13624 5125 -13590
rect 5163 -13624 5195 -13590
rect 5195 -13624 5197 -13590
rect 5235 -13624 5263 -13590
rect 5263 -13624 5269 -13590
rect 5307 -13624 5331 -13590
rect 5331 -13624 5341 -13590
rect 5965 -13624 5975 -13590
rect 5975 -13624 5999 -13590
rect 6037 -13624 6043 -13590
rect 6043 -13624 6071 -13590
rect 6109 -13624 6111 -13590
rect 6111 -13624 6143 -13590
rect 6181 -13624 6213 -13590
rect 6213 -13624 6215 -13590
rect 6253 -13624 6281 -13590
rect 6281 -13624 6287 -13590
rect 6325 -13624 6349 -13590
rect 6349 -13624 6359 -13590
rect 6983 -13624 6993 -13590
rect 6993 -13624 7017 -13590
rect 7055 -13624 7061 -13590
rect 7061 -13624 7089 -13590
rect 7127 -13624 7129 -13590
rect 7129 -13624 7161 -13590
rect 7199 -13624 7231 -13590
rect 7231 -13624 7233 -13590
rect 7271 -13624 7299 -13590
rect 7299 -13624 7305 -13590
rect 7343 -13624 7367 -13590
rect 7367 -13624 7377 -13590
rect 8001 -13624 8011 -13590
rect 8011 -13624 8035 -13590
rect 8073 -13624 8079 -13590
rect 8079 -13624 8107 -13590
rect 8145 -13624 8147 -13590
rect 8147 -13624 8179 -13590
rect 8217 -13624 8249 -13590
rect 8249 -13624 8251 -13590
rect 8289 -13624 8317 -13590
rect 8317 -13624 8323 -13590
rect 8361 -13624 8385 -13590
rect 8385 -13624 8395 -13590
rect 9019 -13624 9029 -13590
rect 9029 -13624 9053 -13590
rect 9091 -13624 9097 -13590
rect 9097 -13624 9125 -13590
rect 9163 -13624 9165 -13590
rect 9165 -13624 9197 -13590
rect 9235 -13624 9267 -13590
rect 9267 -13624 9269 -13590
rect 9307 -13624 9335 -13590
rect 9335 -13624 9341 -13590
rect 9379 -13624 9403 -13590
rect 9403 -13624 9413 -13590
rect 10037 -13624 10047 -13590
rect 10047 -13624 10071 -13590
rect 10109 -13624 10115 -13590
rect 10115 -13624 10143 -13590
rect 10181 -13624 10183 -13590
rect 10183 -13624 10215 -13590
rect 10253 -13624 10285 -13590
rect 10285 -13624 10287 -13590
rect 10325 -13624 10353 -13590
rect 10353 -13624 10359 -13590
rect 10397 -13624 10421 -13590
rect 10421 -13624 10431 -13590
rect 11055 -13624 11065 -13590
rect 11065 -13624 11089 -13590
rect 11127 -13624 11133 -13590
rect 11133 -13624 11161 -13590
rect 11199 -13624 11201 -13590
rect 11201 -13624 11233 -13590
rect 11271 -13624 11303 -13590
rect 11303 -13624 11305 -13590
rect 11343 -13624 11371 -13590
rect 11371 -13624 11377 -13590
rect 11415 -13624 11439 -13590
rect 11439 -13624 11449 -13590
rect 12073 -13624 12083 -13590
rect 12083 -13624 12107 -13590
rect 12145 -13624 12151 -13590
rect 12151 -13624 12179 -13590
rect 12217 -13624 12219 -13590
rect 12219 -13624 12251 -13590
rect 12289 -13624 12321 -13590
rect 12321 -13624 12323 -13590
rect 12361 -13624 12389 -13590
rect 12389 -13624 12395 -13590
rect 12433 -13624 12457 -13590
rect 12457 -13624 12467 -13590
rect 13091 -13624 13101 -13590
rect 13101 -13624 13125 -13590
rect 13163 -13624 13169 -13590
rect 13169 -13624 13197 -13590
rect 13235 -13624 13237 -13590
rect 13237 -13624 13269 -13590
rect 13307 -13624 13339 -13590
rect 13339 -13624 13341 -13590
rect 13379 -13624 13407 -13590
rect 13407 -13624 13413 -13590
rect 13451 -13624 13475 -13590
rect 13475 -13624 13485 -13590
rect 14109 -13624 14119 -13590
rect 14119 -13624 14143 -13590
rect 14181 -13624 14187 -13590
rect 14187 -13624 14215 -13590
rect 14253 -13624 14255 -13590
rect 14255 -13624 14287 -13590
rect 14325 -13624 14357 -13590
rect 14357 -13624 14359 -13590
rect 14397 -13624 14425 -13590
rect 14425 -13624 14431 -13590
rect 14469 -13624 14493 -13590
rect 14493 -13624 14503 -13590
rect 15127 -13624 15137 -13590
rect 15137 -13624 15161 -13590
rect 15199 -13624 15205 -13590
rect 15205 -13624 15233 -13590
rect 15271 -13624 15273 -13590
rect 15273 -13624 15305 -13590
rect 15343 -13624 15375 -13590
rect 15375 -13624 15377 -13590
rect 15415 -13624 15443 -13590
rect 15443 -13624 15449 -13590
rect 15487 -13624 15511 -13590
rect 15511 -13624 15521 -13590
rect 16145 -13624 16155 -13590
rect 16155 -13624 16179 -13590
rect 16217 -13624 16223 -13590
rect 16223 -13624 16251 -13590
rect 16289 -13624 16291 -13590
rect 16291 -13624 16323 -13590
rect 16361 -13624 16393 -13590
rect 16393 -13624 16395 -13590
rect 16433 -13624 16461 -13590
rect 16461 -13624 16467 -13590
rect 16505 -13624 16529 -13590
rect 16529 -13624 16539 -13590
rect 17163 -13624 17173 -13590
rect 17173 -13624 17197 -13590
rect 17235 -13624 17241 -13590
rect 17241 -13624 17269 -13590
rect 17307 -13624 17309 -13590
rect 17309 -13624 17341 -13590
rect 17379 -13624 17411 -13590
rect 17411 -13624 17413 -13590
rect 17451 -13624 17479 -13590
rect 17479 -13624 17485 -13590
rect 17523 -13624 17547 -13590
rect 17547 -13624 17557 -13590
rect 18181 -13624 18191 -13590
rect 18191 -13624 18215 -13590
rect 18253 -13624 18259 -13590
rect 18259 -13624 18287 -13590
rect 18325 -13624 18327 -13590
rect 18327 -13624 18359 -13590
rect 18397 -13624 18429 -13590
rect 18429 -13624 18431 -13590
rect 18469 -13624 18497 -13590
rect 18497 -13624 18503 -13590
rect 18541 -13624 18565 -13590
rect 18565 -13624 18575 -13590
rect 19199 -13624 19209 -13590
rect 19209 -13624 19233 -13590
rect 19271 -13624 19277 -13590
rect 19277 -13624 19305 -13590
rect 19343 -13624 19345 -13590
rect 19345 -13624 19377 -13590
rect 19415 -13624 19447 -13590
rect 19447 -13624 19449 -13590
rect 19487 -13624 19515 -13590
rect 19515 -13624 19521 -13590
rect 19559 -13624 19583 -13590
rect 19583 -13624 19593 -13590
rect 20217 -13624 20227 -13590
rect 20227 -13624 20251 -13590
rect 20289 -13624 20295 -13590
rect 20295 -13624 20323 -13590
rect 20361 -13624 20363 -13590
rect 20363 -13624 20395 -13590
rect 20433 -13624 20465 -13590
rect 20465 -13624 20467 -13590
rect 20505 -13624 20533 -13590
rect 20533 -13624 20539 -13590
rect 20577 -13624 20601 -13590
rect 20601 -13624 20611 -13590
rect 21235 -13624 21245 -13590
rect 21245 -13624 21269 -13590
rect 21307 -13624 21313 -13590
rect 21313 -13624 21341 -13590
rect 21379 -13624 21381 -13590
rect 21381 -13624 21413 -13590
rect 21451 -13624 21483 -13590
rect 21483 -13624 21485 -13590
rect 21523 -13624 21551 -13590
rect 21551 -13624 21557 -13590
rect 21595 -13624 21619 -13590
rect 21619 -13624 21629 -13590
rect 22253 -13624 22263 -13590
rect 22263 -13624 22287 -13590
rect 22325 -13624 22331 -13590
rect 22331 -13624 22359 -13590
rect 22397 -13624 22399 -13590
rect 22399 -13624 22431 -13590
rect 22469 -13624 22501 -13590
rect 22501 -13624 22503 -13590
rect 22541 -13624 22569 -13590
rect 22569 -13624 22575 -13590
rect 22613 -13624 22637 -13590
rect 22637 -13624 22647 -13590
rect -22 -13681 12 -13649
rect -22 -13683 12 -13681
rect -22 -13749 12 -13721
rect -22 -13755 12 -13749
rect -22 -13817 12 -13793
rect -22 -13827 12 -13817
rect -22 -13885 12 -13865
rect -22 -13899 12 -13885
rect 24855 -13607 24889 -13603
rect 24855 -13637 24889 -13607
rect 24855 -13709 24889 -13675
rect 24855 -13777 24889 -13747
rect 24855 -13781 24889 -13777
rect 24855 -13845 24889 -13819
rect 24855 -13853 24889 -13845
rect 24855 -13913 24889 -13891
rect 24855 -13925 24889 -13913
rect -12289 -13981 -12255 -13963
rect -12289 -13997 -12255 -13981
rect -8855 -14002 -8845 -13968
rect -8845 -14002 -8821 -13968
rect -8783 -14002 -8777 -13968
rect -8777 -14002 -8749 -13968
rect -8711 -14002 -8709 -13968
rect -8709 -14002 -8677 -13968
rect -8639 -14002 -8607 -13968
rect -8607 -14002 -8605 -13968
rect -8567 -14002 -8539 -13968
rect -8539 -14002 -8533 -13968
rect -8495 -14002 -8471 -13968
rect -8471 -14002 -8461 -13968
rect -7837 -14002 -7827 -13968
rect -7827 -14002 -7803 -13968
rect -7765 -14002 -7759 -13968
rect -7759 -14002 -7731 -13968
rect -7693 -14002 -7691 -13968
rect -7691 -14002 -7659 -13968
rect -7621 -14002 -7589 -13968
rect -7589 -14002 -7587 -13968
rect -7549 -14002 -7521 -13968
rect -7521 -14002 -7515 -13968
rect -7477 -14002 -7453 -13968
rect -7453 -14002 -7443 -13968
rect -6819 -14002 -6809 -13968
rect -6809 -14002 -6785 -13968
rect -6747 -14002 -6741 -13968
rect -6741 -14002 -6713 -13968
rect -6675 -14002 -6673 -13968
rect -6673 -14002 -6641 -13968
rect -6603 -14002 -6571 -13968
rect -6571 -14002 -6569 -13968
rect -6531 -14002 -6503 -13968
rect -6503 -14002 -6497 -13968
rect -6459 -14002 -6435 -13968
rect -6435 -14002 -6425 -13968
rect -5801 -14002 -5791 -13968
rect -5791 -14002 -5767 -13968
rect -5729 -14002 -5723 -13968
rect -5723 -14002 -5695 -13968
rect -5657 -14002 -5655 -13968
rect -5655 -14002 -5623 -13968
rect -5585 -14002 -5553 -13968
rect -5553 -14002 -5551 -13968
rect -5513 -14002 -5485 -13968
rect -5485 -14002 -5479 -13968
rect -5441 -14002 -5417 -13968
rect -5417 -14002 -5407 -13968
rect -4783 -14002 -4773 -13968
rect -4773 -14002 -4749 -13968
rect -4711 -14002 -4705 -13968
rect -4705 -14002 -4677 -13968
rect -4639 -14002 -4637 -13968
rect -4637 -14002 -4605 -13968
rect -4567 -14002 -4535 -13968
rect -4535 -14002 -4533 -13968
rect -4495 -14002 -4467 -13968
rect -4467 -14002 -4461 -13968
rect -4423 -14002 -4399 -13968
rect -4399 -14002 -4389 -13968
rect -3765 -14002 -3755 -13968
rect -3755 -14002 -3731 -13968
rect -3693 -14002 -3687 -13968
rect -3687 -14002 -3659 -13968
rect -3621 -14002 -3619 -13968
rect -3619 -14002 -3587 -13968
rect -3549 -14002 -3517 -13968
rect -3517 -14002 -3515 -13968
rect -3477 -14002 -3449 -13968
rect -3449 -14002 -3443 -13968
rect -3405 -14002 -3381 -13968
rect -3381 -14002 -3371 -13968
rect -2747 -14002 -2737 -13968
rect -2737 -14002 -2713 -13968
rect -2675 -14002 -2669 -13968
rect -2669 -14002 -2641 -13968
rect -2603 -14002 -2601 -13968
rect -2601 -14002 -2569 -13968
rect -2531 -14002 -2499 -13968
rect -2499 -14002 -2497 -13968
rect -2459 -14002 -2431 -13968
rect -2431 -14002 -2425 -13968
rect -2387 -14002 -2363 -13968
rect -2363 -14002 -2353 -13968
rect -1729 -14002 -1719 -13968
rect -1719 -14002 -1695 -13968
rect -1657 -14002 -1651 -13968
rect -1651 -14002 -1623 -13968
rect -1585 -14002 -1583 -13968
rect -1583 -14002 -1551 -13968
rect -1513 -14002 -1481 -13968
rect -1481 -14002 -1479 -13968
rect -1441 -14002 -1413 -13968
rect -1413 -14002 -1407 -13968
rect -1369 -14002 -1345 -13968
rect -1345 -14002 -1335 -13968
rect -711 -14002 -701 -13968
rect -701 -14002 -677 -13968
rect -639 -14002 -633 -13968
rect -633 -14002 -605 -13968
rect -567 -14002 -565 -13968
rect -565 -14002 -533 -13968
rect -495 -14002 -463 -13968
rect -463 -14002 -461 -13968
rect -423 -14002 -395 -13968
rect -395 -14002 -389 -13968
rect -351 -14002 -327 -13968
rect -327 -14002 -317 -13968
rect 24855 -13981 24889 -13963
rect 24855 -13997 24889 -13981
rect -12289 -14049 -12255 -14035
rect -12289 -14069 -12255 -14049
rect 24855 -14049 24889 -14035
rect 24855 -14069 24889 -14049
rect -12289 -14117 -12255 -14107
rect -12289 -14141 -12255 -14117
rect -8855 -14110 -8845 -14076
rect -8845 -14110 -8821 -14076
rect -8783 -14110 -8777 -14076
rect -8777 -14110 -8749 -14076
rect -8711 -14110 -8709 -14076
rect -8709 -14110 -8677 -14076
rect -8639 -14110 -8607 -14076
rect -8607 -14110 -8605 -14076
rect -8567 -14110 -8539 -14076
rect -8539 -14110 -8533 -14076
rect -8495 -14110 -8471 -14076
rect -8471 -14110 -8461 -14076
rect -7837 -14110 -7827 -14076
rect -7827 -14110 -7803 -14076
rect -7765 -14110 -7759 -14076
rect -7759 -14110 -7731 -14076
rect -7693 -14110 -7691 -14076
rect -7691 -14110 -7659 -14076
rect -7621 -14110 -7589 -14076
rect -7589 -14110 -7587 -14076
rect -7549 -14110 -7521 -14076
rect -7521 -14110 -7515 -14076
rect -7477 -14110 -7453 -14076
rect -7453 -14110 -7443 -14076
rect -6819 -14110 -6809 -14076
rect -6809 -14110 -6785 -14076
rect -6747 -14110 -6741 -14076
rect -6741 -14110 -6713 -14076
rect -6675 -14110 -6673 -14076
rect -6673 -14110 -6641 -14076
rect -6603 -14110 -6571 -14076
rect -6571 -14110 -6569 -14076
rect -6531 -14110 -6503 -14076
rect -6503 -14110 -6497 -14076
rect -6459 -14110 -6435 -14076
rect -6435 -14110 -6425 -14076
rect -5801 -14110 -5791 -14076
rect -5791 -14110 -5767 -14076
rect -5729 -14110 -5723 -14076
rect -5723 -14110 -5695 -14076
rect -5657 -14110 -5655 -14076
rect -5655 -14110 -5623 -14076
rect -5585 -14110 -5553 -14076
rect -5553 -14110 -5551 -14076
rect -5513 -14110 -5485 -14076
rect -5485 -14110 -5479 -14076
rect -5441 -14110 -5417 -14076
rect -5417 -14110 -5407 -14076
rect -4783 -14110 -4773 -14076
rect -4773 -14110 -4749 -14076
rect -4711 -14110 -4705 -14076
rect -4705 -14110 -4677 -14076
rect -4639 -14110 -4637 -14076
rect -4637 -14110 -4605 -14076
rect -4567 -14110 -4535 -14076
rect -4535 -14110 -4533 -14076
rect -4495 -14110 -4467 -14076
rect -4467 -14110 -4461 -14076
rect -4423 -14110 -4399 -14076
rect -4399 -14110 -4389 -14076
rect -3765 -14110 -3755 -14076
rect -3755 -14110 -3731 -14076
rect -3693 -14110 -3687 -14076
rect -3687 -14110 -3659 -14076
rect -3621 -14110 -3619 -14076
rect -3619 -14110 -3587 -14076
rect -3549 -14110 -3517 -14076
rect -3517 -14110 -3515 -14076
rect -3477 -14110 -3449 -14076
rect -3449 -14110 -3443 -14076
rect -3405 -14110 -3381 -14076
rect -3381 -14110 -3371 -14076
rect -2747 -14110 -2737 -14076
rect -2737 -14110 -2713 -14076
rect -2675 -14110 -2669 -14076
rect -2669 -14110 -2641 -14076
rect -2603 -14110 -2601 -14076
rect -2601 -14110 -2569 -14076
rect -2531 -14110 -2499 -14076
rect -2499 -14110 -2497 -14076
rect -2459 -14110 -2431 -14076
rect -2431 -14110 -2425 -14076
rect -2387 -14110 -2363 -14076
rect -2363 -14110 -2353 -14076
rect -1729 -14110 -1719 -14076
rect -1719 -14110 -1695 -14076
rect -1657 -14110 -1651 -14076
rect -1651 -14110 -1623 -14076
rect -1585 -14110 -1583 -14076
rect -1583 -14110 -1551 -14076
rect -1513 -14110 -1481 -14076
rect -1481 -14110 -1479 -14076
rect -1441 -14110 -1413 -14076
rect -1413 -14110 -1407 -14076
rect -1369 -14110 -1345 -14076
rect -1345 -14110 -1335 -14076
rect -711 -14110 -701 -14076
rect -701 -14110 -677 -14076
rect -639 -14110 -633 -14076
rect -633 -14110 -605 -14076
rect -567 -14110 -565 -14076
rect -565 -14110 -533 -14076
rect -495 -14110 -463 -14076
rect -463 -14110 -461 -14076
rect -423 -14110 -395 -14076
rect -395 -14110 -389 -14076
rect -351 -14110 -327 -14076
rect -327 -14110 -317 -14076
rect -12289 -14185 -12255 -14179
rect -12289 -14213 -12255 -14185
rect -12289 -14253 -12255 -14251
rect -12289 -14285 -12255 -14253
rect -12289 -14355 -12255 -14323
rect -12289 -14357 -12255 -14355
rect -12289 -14423 -12255 -14395
rect -12289 -14429 -12255 -14423
rect -12289 -14491 -12255 -14467
rect -12289 -14501 -12255 -14491
rect -12289 -14559 -12255 -14539
rect -12289 -14573 -12255 -14559
rect -12289 -14627 -12255 -14611
rect -12289 -14645 -12255 -14627
rect -12289 -14695 -12255 -14683
rect -12289 -14717 -12255 -14695
rect -9184 -14193 -9150 -14179
rect -9184 -14213 -9150 -14193
rect -9184 -14261 -9150 -14251
rect -9184 -14285 -9150 -14261
rect -9184 -14329 -9150 -14323
rect -9184 -14357 -9150 -14329
rect -9184 -14397 -9150 -14395
rect -9184 -14429 -9150 -14397
rect -9184 -14499 -9150 -14467
rect -9184 -14501 -9150 -14499
rect -9184 -14567 -9150 -14539
rect -9184 -14573 -9150 -14567
rect -9184 -14635 -9150 -14611
rect -9184 -14645 -9150 -14635
rect -9184 -14703 -9150 -14683
rect -9184 -14717 -9150 -14703
rect -8166 -14193 -8132 -14179
rect -8166 -14213 -8132 -14193
rect -8166 -14261 -8132 -14251
rect -8166 -14285 -8132 -14261
rect -8166 -14329 -8132 -14323
rect -8166 -14357 -8132 -14329
rect -8166 -14397 -8132 -14395
rect -8166 -14429 -8132 -14397
rect -8166 -14499 -8132 -14467
rect -8166 -14501 -8132 -14499
rect -8166 -14567 -8132 -14539
rect -8166 -14573 -8132 -14567
rect -8166 -14635 -8132 -14611
rect -8166 -14645 -8132 -14635
rect -8166 -14703 -8132 -14683
rect -8166 -14717 -8132 -14703
rect -7148 -14193 -7114 -14179
rect -7148 -14213 -7114 -14193
rect -7148 -14261 -7114 -14251
rect -7148 -14285 -7114 -14261
rect -7148 -14329 -7114 -14323
rect -7148 -14357 -7114 -14329
rect -7148 -14397 -7114 -14395
rect -7148 -14429 -7114 -14397
rect -7148 -14499 -7114 -14467
rect -7148 -14501 -7114 -14499
rect -7148 -14567 -7114 -14539
rect -7148 -14573 -7114 -14567
rect -7148 -14635 -7114 -14611
rect -7148 -14645 -7114 -14635
rect -7148 -14703 -7114 -14683
rect -7148 -14717 -7114 -14703
rect -6130 -14193 -6096 -14179
rect -6130 -14213 -6096 -14193
rect -6130 -14261 -6096 -14251
rect -6130 -14285 -6096 -14261
rect -6130 -14329 -6096 -14323
rect -6130 -14357 -6096 -14329
rect -6130 -14397 -6096 -14395
rect -6130 -14429 -6096 -14397
rect -6130 -14499 -6096 -14467
rect -6130 -14501 -6096 -14499
rect -6130 -14567 -6096 -14539
rect -6130 -14573 -6096 -14567
rect -6130 -14635 -6096 -14611
rect -6130 -14645 -6096 -14635
rect -6130 -14703 -6096 -14683
rect -6130 -14717 -6096 -14703
rect -5112 -14193 -5078 -14179
rect -5112 -14213 -5078 -14193
rect -5112 -14261 -5078 -14251
rect -5112 -14285 -5078 -14261
rect -5112 -14329 -5078 -14323
rect -5112 -14357 -5078 -14329
rect -5112 -14397 -5078 -14395
rect -5112 -14429 -5078 -14397
rect -5112 -14499 -5078 -14467
rect -5112 -14501 -5078 -14499
rect -5112 -14567 -5078 -14539
rect -5112 -14573 -5078 -14567
rect -5112 -14635 -5078 -14611
rect -5112 -14645 -5078 -14635
rect -5112 -14703 -5078 -14683
rect -5112 -14717 -5078 -14703
rect -4094 -14193 -4060 -14179
rect -4094 -14213 -4060 -14193
rect -4094 -14261 -4060 -14251
rect -4094 -14285 -4060 -14261
rect -4094 -14329 -4060 -14323
rect -4094 -14357 -4060 -14329
rect -4094 -14397 -4060 -14395
rect -4094 -14429 -4060 -14397
rect -4094 -14499 -4060 -14467
rect -4094 -14501 -4060 -14499
rect -4094 -14567 -4060 -14539
rect -4094 -14573 -4060 -14567
rect -4094 -14635 -4060 -14611
rect -4094 -14645 -4060 -14635
rect -4094 -14703 -4060 -14683
rect -4094 -14717 -4060 -14703
rect -3076 -14193 -3042 -14179
rect -3076 -14213 -3042 -14193
rect -3076 -14261 -3042 -14251
rect -3076 -14285 -3042 -14261
rect -3076 -14329 -3042 -14323
rect -3076 -14357 -3042 -14329
rect -3076 -14397 -3042 -14395
rect -3076 -14429 -3042 -14397
rect -3076 -14499 -3042 -14467
rect -3076 -14501 -3042 -14499
rect -3076 -14567 -3042 -14539
rect -3076 -14573 -3042 -14567
rect -3076 -14635 -3042 -14611
rect -3076 -14645 -3042 -14635
rect -3076 -14703 -3042 -14683
rect -3076 -14717 -3042 -14703
rect -2058 -14193 -2024 -14179
rect -2058 -14213 -2024 -14193
rect -2058 -14261 -2024 -14251
rect -2058 -14285 -2024 -14261
rect -2058 -14329 -2024 -14323
rect -2058 -14357 -2024 -14329
rect -2058 -14397 -2024 -14395
rect -2058 -14429 -2024 -14397
rect -2058 -14499 -2024 -14467
rect -2058 -14501 -2024 -14499
rect -2058 -14567 -2024 -14539
rect -2058 -14573 -2024 -14567
rect -2058 -14635 -2024 -14611
rect -2058 -14645 -2024 -14635
rect -2058 -14703 -2024 -14683
rect -2058 -14717 -2024 -14703
rect -1040 -14193 -1006 -14179
rect -1040 -14213 -1006 -14193
rect -1040 -14261 -1006 -14251
rect -1040 -14285 -1006 -14261
rect -1040 -14329 -1006 -14323
rect -1040 -14357 -1006 -14329
rect -1040 -14397 -1006 -14395
rect -1040 -14429 -1006 -14397
rect -1040 -14499 -1006 -14467
rect -1040 -14501 -1006 -14499
rect -1040 -14567 -1006 -14539
rect -1040 -14573 -1006 -14567
rect -1040 -14635 -1006 -14611
rect -1040 -14645 -1006 -14635
rect -1040 -14703 -1006 -14683
rect -1040 -14717 -1006 -14703
rect 2911 -14146 2921 -14112
rect 2921 -14146 2945 -14112
rect 2983 -14146 2989 -14112
rect 2989 -14146 3017 -14112
rect 3055 -14146 3057 -14112
rect 3057 -14146 3089 -14112
rect 3127 -14146 3159 -14112
rect 3159 -14146 3161 -14112
rect 3199 -14146 3227 -14112
rect 3227 -14146 3233 -14112
rect 3271 -14146 3295 -14112
rect 3295 -14146 3305 -14112
rect 3929 -14146 3939 -14112
rect 3939 -14146 3963 -14112
rect 4001 -14146 4007 -14112
rect 4007 -14146 4035 -14112
rect 4073 -14146 4075 -14112
rect 4075 -14146 4107 -14112
rect 4145 -14146 4177 -14112
rect 4177 -14146 4179 -14112
rect 4217 -14146 4245 -14112
rect 4245 -14146 4251 -14112
rect 4289 -14146 4313 -14112
rect 4313 -14146 4323 -14112
rect 4947 -14146 4957 -14112
rect 4957 -14146 4981 -14112
rect 5019 -14146 5025 -14112
rect 5025 -14146 5053 -14112
rect 5091 -14146 5093 -14112
rect 5093 -14146 5125 -14112
rect 5163 -14146 5195 -14112
rect 5195 -14146 5197 -14112
rect 5235 -14146 5263 -14112
rect 5263 -14146 5269 -14112
rect 5307 -14146 5331 -14112
rect 5331 -14146 5341 -14112
rect 5965 -14146 5975 -14112
rect 5975 -14146 5999 -14112
rect 6037 -14146 6043 -14112
rect 6043 -14146 6071 -14112
rect 6109 -14146 6111 -14112
rect 6111 -14146 6143 -14112
rect 6181 -14146 6213 -14112
rect 6213 -14146 6215 -14112
rect 6253 -14146 6281 -14112
rect 6281 -14146 6287 -14112
rect 6325 -14146 6349 -14112
rect 6349 -14146 6359 -14112
rect 6983 -14146 6993 -14112
rect 6993 -14146 7017 -14112
rect 7055 -14146 7061 -14112
rect 7061 -14146 7089 -14112
rect 7127 -14146 7129 -14112
rect 7129 -14146 7161 -14112
rect 7199 -14146 7231 -14112
rect 7231 -14146 7233 -14112
rect 7271 -14146 7299 -14112
rect 7299 -14146 7305 -14112
rect 7343 -14146 7367 -14112
rect 7367 -14146 7377 -14112
rect 8001 -14146 8011 -14112
rect 8011 -14146 8035 -14112
rect 8073 -14146 8079 -14112
rect 8079 -14146 8107 -14112
rect 8145 -14146 8147 -14112
rect 8147 -14146 8179 -14112
rect 8217 -14146 8249 -14112
rect 8249 -14146 8251 -14112
rect 8289 -14146 8317 -14112
rect 8317 -14146 8323 -14112
rect 8361 -14146 8385 -14112
rect 8385 -14146 8395 -14112
rect 9019 -14146 9029 -14112
rect 9029 -14146 9053 -14112
rect 9091 -14146 9097 -14112
rect 9097 -14146 9125 -14112
rect 9163 -14146 9165 -14112
rect 9165 -14146 9197 -14112
rect 9235 -14146 9267 -14112
rect 9267 -14146 9269 -14112
rect 9307 -14146 9335 -14112
rect 9335 -14146 9341 -14112
rect 9379 -14146 9403 -14112
rect 9403 -14146 9413 -14112
rect 10037 -14146 10047 -14112
rect 10047 -14146 10071 -14112
rect 10109 -14146 10115 -14112
rect 10115 -14146 10143 -14112
rect 10181 -14146 10183 -14112
rect 10183 -14146 10215 -14112
rect 10253 -14146 10285 -14112
rect 10285 -14146 10287 -14112
rect 10325 -14146 10353 -14112
rect 10353 -14146 10359 -14112
rect 10397 -14146 10421 -14112
rect 10421 -14146 10431 -14112
rect 11055 -14146 11065 -14112
rect 11065 -14146 11089 -14112
rect 11127 -14146 11133 -14112
rect 11133 -14146 11161 -14112
rect 11199 -14146 11201 -14112
rect 11201 -14146 11233 -14112
rect 11271 -14146 11303 -14112
rect 11303 -14146 11305 -14112
rect 11343 -14146 11371 -14112
rect 11371 -14146 11377 -14112
rect 11415 -14146 11439 -14112
rect 11439 -14146 11449 -14112
rect 12073 -14146 12083 -14112
rect 12083 -14146 12107 -14112
rect 12145 -14146 12151 -14112
rect 12151 -14146 12179 -14112
rect 12217 -14146 12219 -14112
rect 12219 -14146 12251 -14112
rect 12289 -14146 12321 -14112
rect 12321 -14146 12323 -14112
rect 12361 -14146 12389 -14112
rect 12389 -14146 12395 -14112
rect 12433 -14146 12457 -14112
rect 12457 -14146 12467 -14112
rect 13091 -14146 13101 -14112
rect 13101 -14146 13125 -14112
rect 13163 -14146 13169 -14112
rect 13169 -14146 13197 -14112
rect 13235 -14146 13237 -14112
rect 13237 -14146 13269 -14112
rect 13307 -14146 13339 -14112
rect 13339 -14146 13341 -14112
rect 13379 -14146 13407 -14112
rect 13407 -14146 13413 -14112
rect 13451 -14146 13475 -14112
rect 13475 -14146 13485 -14112
rect 14109 -14146 14119 -14112
rect 14119 -14146 14143 -14112
rect 14181 -14146 14187 -14112
rect 14187 -14146 14215 -14112
rect 14253 -14146 14255 -14112
rect 14255 -14146 14287 -14112
rect 14325 -14146 14357 -14112
rect 14357 -14146 14359 -14112
rect 14397 -14146 14425 -14112
rect 14425 -14146 14431 -14112
rect 14469 -14146 14493 -14112
rect 14493 -14146 14503 -14112
rect 15127 -14146 15137 -14112
rect 15137 -14146 15161 -14112
rect 15199 -14146 15205 -14112
rect 15205 -14146 15233 -14112
rect 15271 -14146 15273 -14112
rect 15273 -14146 15305 -14112
rect 15343 -14146 15375 -14112
rect 15375 -14146 15377 -14112
rect 15415 -14146 15443 -14112
rect 15443 -14146 15449 -14112
rect 15487 -14146 15511 -14112
rect 15511 -14146 15521 -14112
rect 16145 -14146 16155 -14112
rect 16155 -14146 16179 -14112
rect 16217 -14146 16223 -14112
rect 16223 -14146 16251 -14112
rect 16289 -14146 16291 -14112
rect 16291 -14146 16323 -14112
rect 16361 -14146 16393 -14112
rect 16393 -14146 16395 -14112
rect 16433 -14146 16461 -14112
rect 16461 -14146 16467 -14112
rect 16505 -14146 16529 -14112
rect 16529 -14146 16539 -14112
rect 17163 -14146 17173 -14112
rect 17173 -14146 17197 -14112
rect 17235 -14146 17241 -14112
rect 17241 -14146 17269 -14112
rect 17307 -14146 17309 -14112
rect 17309 -14146 17341 -14112
rect 17379 -14146 17411 -14112
rect 17411 -14146 17413 -14112
rect 17451 -14146 17479 -14112
rect 17479 -14146 17485 -14112
rect 17523 -14146 17547 -14112
rect 17547 -14146 17557 -14112
rect 18181 -14146 18191 -14112
rect 18191 -14146 18215 -14112
rect 18253 -14146 18259 -14112
rect 18259 -14146 18287 -14112
rect 18325 -14146 18327 -14112
rect 18327 -14146 18359 -14112
rect 18397 -14146 18429 -14112
rect 18429 -14146 18431 -14112
rect 18469 -14146 18497 -14112
rect 18497 -14146 18503 -14112
rect 18541 -14146 18565 -14112
rect 18565 -14146 18575 -14112
rect 19199 -14146 19209 -14112
rect 19209 -14146 19233 -14112
rect 19271 -14146 19277 -14112
rect 19277 -14146 19305 -14112
rect 19343 -14146 19345 -14112
rect 19345 -14146 19377 -14112
rect 19415 -14146 19447 -14112
rect 19447 -14146 19449 -14112
rect 19487 -14146 19515 -14112
rect 19515 -14146 19521 -14112
rect 19559 -14146 19583 -14112
rect 19583 -14146 19593 -14112
rect 20217 -14146 20227 -14112
rect 20227 -14146 20251 -14112
rect 20289 -14146 20295 -14112
rect 20295 -14146 20323 -14112
rect 20361 -14146 20363 -14112
rect 20363 -14146 20395 -14112
rect 20433 -14146 20465 -14112
rect 20465 -14146 20467 -14112
rect 20505 -14146 20533 -14112
rect 20533 -14146 20539 -14112
rect 20577 -14146 20601 -14112
rect 20601 -14146 20611 -14112
rect 21235 -14146 21245 -14112
rect 21245 -14146 21269 -14112
rect 21307 -14146 21313 -14112
rect 21313 -14146 21341 -14112
rect 21379 -14146 21381 -14112
rect 21381 -14146 21413 -14112
rect 21451 -14146 21483 -14112
rect 21483 -14146 21485 -14112
rect 21523 -14146 21551 -14112
rect 21551 -14146 21557 -14112
rect 21595 -14146 21619 -14112
rect 21619 -14146 21629 -14112
rect 22253 -14146 22263 -14112
rect 22263 -14146 22287 -14112
rect 22325 -14146 22331 -14112
rect 22331 -14146 22359 -14112
rect 22397 -14146 22399 -14112
rect 22399 -14146 22431 -14112
rect 22469 -14146 22501 -14112
rect 22501 -14146 22503 -14112
rect 22541 -14146 22569 -14112
rect 22569 -14146 22575 -14112
rect 22613 -14146 22637 -14112
rect 22637 -14146 22647 -14112
rect 24855 -14117 24889 -14107
rect 24855 -14141 24889 -14117
rect -22 -14193 12 -14179
rect -22 -14213 12 -14193
rect -22 -14261 12 -14251
rect -22 -14285 12 -14261
rect -22 -14329 12 -14323
rect -22 -14357 12 -14329
rect -22 -14397 12 -14395
rect -22 -14429 12 -14397
rect -22 -14499 12 -14467
rect -22 -14501 12 -14499
rect -22 -14567 12 -14539
rect -22 -14573 12 -14567
rect -22 -14635 12 -14611
rect -22 -14645 12 -14635
rect -22 -14703 12 -14683
rect -22 -14717 12 -14703
rect 2582 -14229 2616 -14215
rect 2582 -14249 2616 -14229
rect 2582 -14297 2616 -14287
rect 2582 -14321 2616 -14297
rect 2582 -14365 2616 -14359
rect 2582 -14393 2616 -14365
rect 2582 -14433 2616 -14431
rect 2582 -14465 2616 -14433
rect 2582 -14535 2616 -14503
rect 2582 -14537 2616 -14535
rect 2582 -14603 2616 -14575
rect 2582 -14609 2616 -14603
rect 2582 -14671 2616 -14647
rect 2582 -14681 2616 -14671
rect 2582 -14739 2616 -14719
rect -12289 -14763 -12255 -14755
rect -12289 -14789 -12255 -14763
rect 2582 -14753 2616 -14739
rect -8855 -14820 -8845 -14786
rect -8845 -14820 -8821 -14786
rect -8783 -14820 -8777 -14786
rect -8777 -14820 -8749 -14786
rect -8711 -14820 -8709 -14786
rect -8709 -14820 -8677 -14786
rect -8639 -14820 -8607 -14786
rect -8607 -14820 -8605 -14786
rect -8567 -14820 -8539 -14786
rect -8539 -14820 -8533 -14786
rect -8495 -14820 -8471 -14786
rect -8471 -14820 -8461 -14786
rect -7837 -14820 -7827 -14786
rect -7827 -14820 -7803 -14786
rect -7765 -14820 -7759 -14786
rect -7759 -14820 -7731 -14786
rect -7693 -14820 -7691 -14786
rect -7691 -14820 -7659 -14786
rect -7621 -14820 -7589 -14786
rect -7589 -14820 -7587 -14786
rect -7549 -14820 -7521 -14786
rect -7521 -14820 -7515 -14786
rect -7477 -14820 -7453 -14786
rect -7453 -14820 -7443 -14786
rect -6819 -14820 -6809 -14786
rect -6809 -14820 -6785 -14786
rect -6747 -14820 -6741 -14786
rect -6741 -14820 -6713 -14786
rect -6675 -14820 -6673 -14786
rect -6673 -14820 -6641 -14786
rect -6603 -14820 -6571 -14786
rect -6571 -14820 -6569 -14786
rect -6531 -14820 -6503 -14786
rect -6503 -14820 -6497 -14786
rect -6459 -14820 -6435 -14786
rect -6435 -14820 -6425 -14786
rect -5801 -14820 -5791 -14786
rect -5791 -14820 -5767 -14786
rect -5729 -14820 -5723 -14786
rect -5723 -14820 -5695 -14786
rect -5657 -14820 -5655 -14786
rect -5655 -14820 -5623 -14786
rect -5585 -14820 -5553 -14786
rect -5553 -14820 -5551 -14786
rect -5513 -14820 -5485 -14786
rect -5485 -14820 -5479 -14786
rect -5441 -14820 -5417 -14786
rect -5417 -14820 -5407 -14786
rect -4783 -14820 -4773 -14786
rect -4773 -14820 -4749 -14786
rect -4711 -14820 -4705 -14786
rect -4705 -14820 -4677 -14786
rect -4639 -14820 -4637 -14786
rect -4637 -14820 -4605 -14786
rect -4567 -14820 -4535 -14786
rect -4535 -14820 -4533 -14786
rect -4495 -14820 -4467 -14786
rect -4467 -14820 -4461 -14786
rect -4423 -14820 -4399 -14786
rect -4399 -14820 -4389 -14786
rect -3765 -14820 -3755 -14786
rect -3755 -14820 -3731 -14786
rect -3693 -14820 -3687 -14786
rect -3687 -14820 -3659 -14786
rect -3621 -14820 -3619 -14786
rect -3619 -14820 -3587 -14786
rect -3549 -14820 -3517 -14786
rect -3517 -14820 -3515 -14786
rect -3477 -14820 -3449 -14786
rect -3449 -14820 -3443 -14786
rect -3405 -14820 -3381 -14786
rect -3381 -14820 -3371 -14786
rect -2747 -14820 -2737 -14786
rect -2737 -14820 -2713 -14786
rect -2675 -14820 -2669 -14786
rect -2669 -14820 -2641 -14786
rect -2603 -14820 -2601 -14786
rect -2601 -14820 -2569 -14786
rect -2531 -14820 -2499 -14786
rect -2499 -14820 -2497 -14786
rect -2459 -14820 -2431 -14786
rect -2431 -14820 -2425 -14786
rect -2387 -14820 -2363 -14786
rect -2363 -14820 -2353 -14786
rect -1729 -14820 -1719 -14786
rect -1719 -14820 -1695 -14786
rect -1657 -14820 -1651 -14786
rect -1651 -14820 -1623 -14786
rect -1585 -14820 -1583 -14786
rect -1583 -14820 -1551 -14786
rect -1513 -14820 -1481 -14786
rect -1481 -14820 -1479 -14786
rect -1441 -14820 -1413 -14786
rect -1413 -14820 -1407 -14786
rect -1369 -14820 -1345 -14786
rect -1345 -14820 -1335 -14786
rect -711 -14820 -701 -14786
rect -701 -14820 -677 -14786
rect -639 -14820 -633 -14786
rect -633 -14820 -605 -14786
rect -567 -14820 -565 -14786
rect -565 -14820 -533 -14786
rect -495 -14820 -463 -14786
rect -463 -14820 -461 -14786
rect -423 -14820 -395 -14786
rect -395 -14820 -389 -14786
rect -351 -14820 -327 -14786
rect -327 -14820 -317 -14786
rect 3600 -14229 3634 -14215
rect 3600 -14249 3634 -14229
rect 3600 -14297 3634 -14287
rect 3600 -14321 3634 -14297
rect 3600 -14365 3634 -14359
rect 3600 -14393 3634 -14365
rect 3600 -14433 3634 -14431
rect 3600 -14465 3634 -14433
rect 3600 -14535 3634 -14503
rect 3600 -14537 3634 -14535
rect 3600 -14603 3634 -14575
rect 3600 -14609 3634 -14603
rect 3600 -14671 3634 -14647
rect 3600 -14681 3634 -14671
rect 3600 -14739 3634 -14719
rect 3600 -14753 3634 -14739
rect 4618 -14229 4652 -14215
rect 4618 -14249 4652 -14229
rect 4618 -14297 4652 -14287
rect 4618 -14321 4652 -14297
rect 4618 -14365 4652 -14359
rect 4618 -14393 4652 -14365
rect 4618 -14433 4652 -14431
rect 4618 -14465 4652 -14433
rect 4618 -14535 4652 -14503
rect 4618 -14537 4652 -14535
rect 4618 -14603 4652 -14575
rect 4618 -14609 4652 -14603
rect 4618 -14671 4652 -14647
rect 4618 -14681 4652 -14671
rect 4618 -14739 4652 -14719
rect 4618 -14753 4652 -14739
rect 5636 -14229 5670 -14215
rect 5636 -14249 5670 -14229
rect 5636 -14297 5670 -14287
rect 5636 -14321 5670 -14297
rect 5636 -14365 5670 -14359
rect 5636 -14393 5670 -14365
rect 5636 -14433 5670 -14431
rect 5636 -14465 5670 -14433
rect 5636 -14535 5670 -14503
rect 5636 -14537 5670 -14535
rect 5636 -14603 5670 -14575
rect 5636 -14609 5670 -14603
rect 5636 -14671 5670 -14647
rect 5636 -14681 5670 -14671
rect 5636 -14739 5670 -14719
rect 5636 -14753 5670 -14739
rect 6654 -14229 6688 -14215
rect 6654 -14249 6688 -14229
rect 6654 -14297 6688 -14287
rect 6654 -14321 6688 -14297
rect 6654 -14365 6688 -14359
rect 6654 -14393 6688 -14365
rect 6654 -14433 6688 -14431
rect 6654 -14465 6688 -14433
rect 6654 -14535 6688 -14503
rect 6654 -14537 6688 -14535
rect 6654 -14603 6688 -14575
rect 6654 -14609 6688 -14603
rect 6654 -14671 6688 -14647
rect 6654 -14681 6688 -14671
rect 6654 -14739 6688 -14719
rect 6654 -14753 6688 -14739
rect 7672 -14229 7706 -14215
rect 7672 -14249 7706 -14229
rect 7672 -14297 7706 -14287
rect 7672 -14321 7706 -14297
rect 7672 -14365 7706 -14359
rect 7672 -14393 7706 -14365
rect 7672 -14433 7706 -14431
rect 7672 -14465 7706 -14433
rect 7672 -14535 7706 -14503
rect 7672 -14537 7706 -14535
rect 7672 -14603 7706 -14575
rect 7672 -14609 7706 -14603
rect 7672 -14671 7706 -14647
rect 7672 -14681 7706 -14671
rect 7672 -14739 7706 -14719
rect 7672 -14753 7706 -14739
rect 8690 -14229 8724 -14215
rect 8690 -14249 8724 -14229
rect 8690 -14297 8724 -14287
rect 8690 -14321 8724 -14297
rect 8690 -14365 8724 -14359
rect 8690 -14393 8724 -14365
rect 8690 -14433 8724 -14431
rect 8690 -14465 8724 -14433
rect 8690 -14535 8724 -14503
rect 8690 -14537 8724 -14535
rect 8690 -14603 8724 -14575
rect 8690 -14609 8724 -14603
rect 8690 -14671 8724 -14647
rect 8690 -14681 8724 -14671
rect 8690 -14739 8724 -14719
rect 8690 -14753 8724 -14739
rect 9708 -14229 9742 -14215
rect 9708 -14249 9742 -14229
rect 9708 -14297 9742 -14287
rect 9708 -14321 9742 -14297
rect 9708 -14365 9742 -14359
rect 9708 -14393 9742 -14365
rect 9708 -14433 9742 -14431
rect 9708 -14465 9742 -14433
rect 9708 -14535 9742 -14503
rect 9708 -14537 9742 -14535
rect 9708 -14603 9742 -14575
rect 9708 -14609 9742 -14603
rect 9708 -14671 9742 -14647
rect 9708 -14681 9742 -14671
rect 9708 -14739 9742 -14719
rect 9708 -14753 9742 -14739
rect 10726 -14229 10760 -14215
rect 10726 -14249 10760 -14229
rect 10726 -14297 10760 -14287
rect 10726 -14321 10760 -14297
rect 10726 -14365 10760 -14359
rect 10726 -14393 10760 -14365
rect 10726 -14433 10760 -14431
rect 10726 -14465 10760 -14433
rect 10726 -14535 10760 -14503
rect 10726 -14537 10760 -14535
rect 10726 -14603 10760 -14575
rect 10726 -14609 10760 -14603
rect 10726 -14671 10760 -14647
rect 10726 -14681 10760 -14671
rect 10726 -14739 10760 -14719
rect 10726 -14753 10760 -14739
rect 11744 -14229 11778 -14215
rect 11744 -14249 11778 -14229
rect 11744 -14297 11778 -14287
rect 11744 -14321 11778 -14297
rect 11744 -14365 11778 -14359
rect 11744 -14393 11778 -14365
rect 11744 -14433 11778 -14431
rect 11744 -14465 11778 -14433
rect 11744 -14535 11778 -14503
rect 11744 -14537 11778 -14535
rect 11744 -14603 11778 -14575
rect 11744 -14609 11778 -14603
rect 11744 -14671 11778 -14647
rect 11744 -14681 11778 -14671
rect 11744 -14739 11778 -14719
rect 11744 -14753 11778 -14739
rect 12762 -14229 12796 -14215
rect 12762 -14249 12796 -14229
rect 12762 -14297 12796 -14287
rect 12762 -14321 12796 -14297
rect 12762 -14365 12796 -14359
rect 12762 -14393 12796 -14365
rect 12762 -14433 12796 -14431
rect 12762 -14465 12796 -14433
rect 12762 -14535 12796 -14503
rect 12762 -14537 12796 -14535
rect 12762 -14603 12796 -14575
rect 12762 -14609 12796 -14603
rect 12762 -14671 12796 -14647
rect 12762 -14681 12796 -14671
rect 12762 -14739 12796 -14719
rect 12762 -14753 12796 -14739
rect 13780 -14229 13814 -14215
rect 13780 -14249 13814 -14229
rect 13780 -14297 13814 -14287
rect 13780 -14321 13814 -14297
rect 13780 -14365 13814 -14359
rect 13780 -14393 13814 -14365
rect 13780 -14433 13814 -14431
rect 13780 -14465 13814 -14433
rect 13780 -14535 13814 -14503
rect 13780 -14537 13814 -14535
rect 13780 -14603 13814 -14575
rect 13780 -14609 13814 -14603
rect 13780 -14671 13814 -14647
rect 13780 -14681 13814 -14671
rect 13780 -14739 13814 -14719
rect 13780 -14753 13814 -14739
rect 14798 -14229 14832 -14215
rect 14798 -14249 14832 -14229
rect 14798 -14297 14832 -14287
rect 14798 -14321 14832 -14297
rect 14798 -14365 14832 -14359
rect 14798 -14393 14832 -14365
rect 14798 -14433 14832 -14431
rect 14798 -14465 14832 -14433
rect 14798 -14535 14832 -14503
rect 14798 -14537 14832 -14535
rect 14798 -14603 14832 -14575
rect 14798 -14609 14832 -14603
rect 14798 -14671 14832 -14647
rect 14798 -14681 14832 -14671
rect 14798 -14739 14832 -14719
rect 14798 -14753 14832 -14739
rect 15816 -14229 15850 -14215
rect 15816 -14249 15850 -14229
rect 15816 -14297 15850 -14287
rect 15816 -14321 15850 -14297
rect 15816 -14365 15850 -14359
rect 15816 -14393 15850 -14365
rect 15816 -14433 15850 -14431
rect 15816 -14465 15850 -14433
rect 15816 -14535 15850 -14503
rect 15816 -14537 15850 -14535
rect 15816 -14603 15850 -14575
rect 15816 -14609 15850 -14603
rect 15816 -14671 15850 -14647
rect 15816 -14681 15850 -14671
rect 15816 -14739 15850 -14719
rect 15816 -14753 15850 -14739
rect 16834 -14229 16868 -14215
rect 16834 -14249 16868 -14229
rect 16834 -14297 16868 -14287
rect 16834 -14321 16868 -14297
rect 16834 -14365 16868 -14359
rect 16834 -14393 16868 -14365
rect 16834 -14433 16868 -14431
rect 16834 -14465 16868 -14433
rect 16834 -14535 16868 -14503
rect 16834 -14537 16868 -14535
rect 16834 -14603 16868 -14575
rect 16834 -14609 16868 -14603
rect 16834 -14671 16868 -14647
rect 16834 -14681 16868 -14671
rect 16834 -14739 16868 -14719
rect 16834 -14753 16868 -14739
rect 17852 -14229 17886 -14215
rect 17852 -14249 17886 -14229
rect 17852 -14297 17886 -14287
rect 17852 -14321 17886 -14297
rect 17852 -14365 17886 -14359
rect 17852 -14393 17886 -14365
rect 17852 -14433 17886 -14431
rect 17852 -14465 17886 -14433
rect 17852 -14535 17886 -14503
rect 17852 -14537 17886 -14535
rect 17852 -14603 17886 -14575
rect 17852 -14609 17886 -14603
rect 17852 -14671 17886 -14647
rect 17852 -14681 17886 -14671
rect 17852 -14739 17886 -14719
rect 17852 -14753 17886 -14739
rect 18870 -14229 18904 -14215
rect 18870 -14249 18904 -14229
rect 18870 -14297 18904 -14287
rect 18870 -14321 18904 -14297
rect 18870 -14365 18904 -14359
rect 18870 -14393 18904 -14365
rect 18870 -14433 18904 -14431
rect 18870 -14465 18904 -14433
rect 18870 -14535 18904 -14503
rect 18870 -14537 18904 -14535
rect 18870 -14603 18904 -14575
rect 18870 -14609 18904 -14603
rect 18870 -14671 18904 -14647
rect 18870 -14681 18904 -14671
rect 18870 -14739 18904 -14719
rect 18870 -14753 18904 -14739
rect 19888 -14229 19922 -14215
rect 19888 -14249 19922 -14229
rect 19888 -14297 19922 -14287
rect 19888 -14321 19922 -14297
rect 19888 -14365 19922 -14359
rect 19888 -14393 19922 -14365
rect 19888 -14433 19922 -14431
rect 19888 -14465 19922 -14433
rect 19888 -14535 19922 -14503
rect 19888 -14537 19922 -14535
rect 19888 -14603 19922 -14575
rect 19888 -14609 19922 -14603
rect 19888 -14671 19922 -14647
rect 19888 -14681 19922 -14671
rect 19888 -14739 19922 -14719
rect 19888 -14753 19922 -14739
rect 20906 -14229 20940 -14215
rect 20906 -14249 20940 -14229
rect 20906 -14297 20940 -14287
rect 20906 -14321 20940 -14297
rect 20906 -14365 20940 -14359
rect 20906 -14393 20940 -14365
rect 20906 -14433 20940 -14431
rect 20906 -14465 20940 -14433
rect 20906 -14535 20940 -14503
rect 20906 -14537 20940 -14535
rect 20906 -14603 20940 -14575
rect 20906 -14609 20940 -14603
rect 20906 -14671 20940 -14647
rect 20906 -14681 20940 -14671
rect 20906 -14739 20940 -14719
rect 20906 -14753 20940 -14739
rect 21924 -14229 21958 -14215
rect 21924 -14249 21958 -14229
rect 21924 -14297 21958 -14287
rect 21924 -14321 21958 -14297
rect 21924 -14365 21958 -14359
rect 21924 -14393 21958 -14365
rect 21924 -14433 21958 -14431
rect 21924 -14465 21958 -14433
rect 21924 -14535 21958 -14503
rect 21924 -14537 21958 -14535
rect 21924 -14603 21958 -14575
rect 21924 -14609 21958 -14603
rect 21924 -14671 21958 -14647
rect 21924 -14681 21958 -14671
rect 21924 -14739 21958 -14719
rect 21924 -14753 21958 -14739
rect 22942 -14229 22976 -14215
rect 22942 -14249 22976 -14229
rect 22942 -14297 22976 -14287
rect 22942 -14321 22976 -14297
rect 22942 -14365 22976 -14359
rect 22942 -14393 22976 -14365
rect 22942 -14433 22976 -14431
rect 22942 -14465 22976 -14433
rect 22942 -14535 22976 -14503
rect 22942 -14537 22976 -14535
rect 22942 -14603 22976 -14575
rect 22942 -14609 22976 -14603
rect 22942 -14671 22976 -14647
rect 22942 -14681 22976 -14671
rect 22942 -14739 22976 -14719
rect 22942 -14753 22976 -14739
rect 24855 -14185 24889 -14179
rect 24855 -14213 24889 -14185
rect 24855 -14253 24889 -14251
rect 24855 -14285 24889 -14253
rect 24855 -14355 24889 -14323
rect 24855 -14357 24889 -14355
rect 24855 -14423 24889 -14395
rect 24855 -14429 24889 -14423
rect 24855 -14491 24889 -14467
rect 24855 -14501 24889 -14491
rect 24855 -14559 24889 -14539
rect 24855 -14573 24889 -14559
rect 24855 -14627 24889 -14611
rect 24855 -14645 24889 -14627
rect 24855 -14695 24889 -14683
rect 24855 -14717 24889 -14695
rect 24855 -14763 24889 -14755
rect 24855 -14789 24889 -14763
rect -12289 -14831 -12255 -14827
rect -12289 -14861 -12255 -14831
rect 2911 -14856 2921 -14822
rect 2921 -14856 2945 -14822
rect 2983 -14856 2989 -14822
rect 2989 -14856 3017 -14822
rect 3055 -14856 3057 -14822
rect 3057 -14856 3089 -14822
rect 3127 -14856 3159 -14822
rect 3159 -14856 3161 -14822
rect 3199 -14856 3227 -14822
rect 3227 -14856 3233 -14822
rect 3271 -14856 3295 -14822
rect 3295 -14856 3305 -14822
rect 3929 -14856 3939 -14822
rect 3939 -14856 3963 -14822
rect 4001 -14856 4007 -14822
rect 4007 -14856 4035 -14822
rect 4073 -14856 4075 -14822
rect 4075 -14856 4107 -14822
rect 4145 -14856 4177 -14822
rect 4177 -14856 4179 -14822
rect 4217 -14856 4245 -14822
rect 4245 -14856 4251 -14822
rect 4289 -14856 4313 -14822
rect 4313 -14856 4323 -14822
rect 4947 -14856 4957 -14822
rect 4957 -14856 4981 -14822
rect 5019 -14856 5025 -14822
rect 5025 -14856 5053 -14822
rect 5091 -14856 5093 -14822
rect 5093 -14856 5125 -14822
rect 5163 -14856 5195 -14822
rect 5195 -14856 5197 -14822
rect 5235 -14856 5263 -14822
rect 5263 -14856 5269 -14822
rect 5307 -14856 5331 -14822
rect 5331 -14856 5341 -14822
rect 5965 -14856 5975 -14822
rect 5975 -14856 5999 -14822
rect 6037 -14856 6043 -14822
rect 6043 -14856 6071 -14822
rect 6109 -14856 6111 -14822
rect 6111 -14856 6143 -14822
rect 6181 -14856 6213 -14822
rect 6213 -14856 6215 -14822
rect 6253 -14856 6281 -14822
rect 6281 -14856 6287 -14822
rect 6325 -14856 6349 -14822
rect 6349 -14856 6359 -14822
rect 6983 -14856 6993 -14822
rect 6993 -14856 7017 -14822
rect 7055 -14856 7061 -14822
rect 7061 -14856 7089 -14822
rect 7127 -14856 7129 -14822
rect 7129 -14856 7161 -14822
rect 7199 -14856 7231 -14822
rect 7231 -14856 7233 -14822
rect 7271 -14856 7299 -14822
rect 7299 -14856 7305 -14822
rect 7343 -14856 7367 -14822
rect 7367 -14856 7377 -14822
rect 8001 -14856 8011 -14822
rect 8011 -14856 8035 -14822
rect 8073 -14856 8079 -14822
rect 8079 -14856 8107 -14822
rect 8145 -14856 8147 -14822
rect 8147 -14856 8179 -14822
rect 8217 -14856 8249 -14822
rect 8249 -14856 8251 -14822
rect 8289 -14856 8317 -14822
rect 8317 -14856 8323 -14822
rect 8361 -14856 8385 -14822
rect 8385 -14856 8395 -14822
rect 9019 -14856 9029 -14822
rect 9029 -14856 9053 -14822
rect 9091 -14856 9097 -14822
rect 9097 -14856 9125 -14822
rect 9163 -14856 9165 -14822
rect 9165 -14856 9197 -14822
rect 9235 -14856 9267 -14822
rect 9267 -14856 9269 -14822
rect 9307 -14856 9335 -14822
rect 9335 -14856 9341 -14822
rect 9379 -14856 9403 -14822
rect 9403 -14856 9413 -14822
rect 10037 -14856 10047 -14822
rect 10047 -14856 10071 -14822
rect 10109 -14856 10115 -14822
rect 10115 -14856 10143 -14822
rect 10181 -14856 10183 -14822
rect 10183 -14856 10215 -14822
rect 10253 -14856 10285 -14822
rect 10285 -14856 10287 -14822
rect 10325 -14856 10353 -14822
rect 10353 -14856 10359 -14822
rect 10397 -14856 10421 -14822
rect 10421 -14856 10431 -14822
rect 11055 -14856 11065 -14822
rect 11065 -14856 11089 -14822
rect 11127 -14856 11133 -14822
rect 11133 -14856 11161 -14822
rect 11199 -14856 11201 -14822
rect 11201 -14856 11233 -14822
rect 11271 -14856 11303 -14822
rect 11303 -14856 11305 -14822
rect 11343 -14856 11371 -14822
rect 11371 -14856 11377 -14822
rect 11415 -14856 11439 -14822
rect 11439 -14856 11449 -14822
rect 12073 -14856 12083 -14822
rect 12083 -14856 12107 -14822
rect 12145 -14856 12151 -14822
rect 12151 -14856 12179 -14822
rect 12217 -14856 12219 -14822
rect 12219 -14856 12251 -14822
rect 12289 -14856 12321 -14822
rect 12321 -14856 12323 -14822
rect 12361 -14856 12389 -14822
rect 12389 -14856 12395 -14822
rect 12433 -14856 12457 -14822
rect 12457 -14856 12467 -14822
rect 13091 -14856 13101 -14822
rect 13101 -14856 13125 -14822
rect 13163 -14856 13169 -14822
rect 13169 -14856 13197 -14822
rect 13235 -14856 13237 -14822
rect 13237 -14856 13269 -14822
rect 13307 -14856 13339 -14822
rect 13339 -14856 13341 -14822
rect 13379 -14856 13407 -14822
rect 13407 -14856 13413 -14822
rect 13451 -14856 13475 -14822
rect 13475 -14856 13485 -14822
rect 14109 -14856 14119 -14822
rect 14119 -14856 14143 -14822
rect 14181 -14856 14187 -14822
rect 14187 -14856 14215 -14822
rect 14253 -14856 14255 -14822
rect 14255 -14856 14287 -14822
rect 14325 -14856 14357 -14822
rect 14357 -14856 14359 -14822
rect 14397 -14856 14425 -14822
rect 14425 -14856 14431 -14822
rect 14469 -14856 14493 -14822
rect 14493 -14856 14503 -14822
rect 15127 -14856 15137 -14822
rect 15137 -14856 15161 -14822
rect 15199 -14856 15205 -14822
rect 15205 -14856 15233 -14822
rect 15271 -14856 15273 -14822
rect 15273 -14856 15305 -14822
rect 15343 -14856 15375 -14822
rect 15375 -14856 15377 -14822
rect 15415 -14856 15443 -14822
rect 15443 -14856 15449 -14822
rect 15487 -14856 15511 -14822
rect 15511 -14856 15521 -14822
rect 16145 -14856 16155 -14822
rect 16155 -14856 16179 -14822
rect 16217 -14856 16223 -14822
rect 16223 -14856 16251 -14822
rect 16289 -14856 16291 -14822
rect 16291 -14856 16323 -14822
rect 16361 -14856 16393 -14822
rect 16393 -14856 16395 -14822
rect 16433 -14856 16461 -14822
rect 16461 -14856 16467 -14822
rect 16505 -14856 16529 -14822
rect 16529 -14856 16539 -14822
rect 17163 -14856 17173 -14822
rect 17173 -14856 17197 -14822
rect 17235 -14856 17241 -14822
rect 17241 -14856 17269 -14822
rect 17379 -14856 17411 -14822
rect 17411 -14856 17413 -14822
rect 17451 -14856 17479 -14822
rect 17479 -14856 17485 -14822
rect 17523 -14856 17547 -14822
rect 17547 -14856 17557 -14822
rect 18181 -14856 18191 -14822
rect 18191 -14856 18215 -14822
rect 18253 -14856 18259 -14822
rect 18259 -14856 18287 -14822
rect 18469 -14856 18497 -14822
rect 18497 -14856 18503 -14822
rect 18541 -14856 18565 -14822
rect 18565 -14856 18575 -14822
rect 19199 -14856 19209 -14822
rect 19209 -14856 19233 -14822
rect 19271 -14856 19277 -14822
rect 19277 -14856 19305 -14822
rect 19343 -14856 19345 -14822
rect 19345 -14856 19377 -14822
rect 19415 -14856 19447 -14822
rect 19447 -14856 19449 -14822
rect 19487 -14856 19515 -14822
rect 19515 -14856 19521 -14822
rect 19559 -14856 19583 -14822
rect 19583 -14856 19593 -14822
rect 20217 -14856 20227 -14822
rect 20227 -14856 20251 -14822
rect 20289 -14856 20295 -14822
rect 20295 -14856 20323 -14822
rect 20361 -14856 20363 -14822
rect 20363 -14856 20395 -14822
rect 20433 -14856 20465 -14822
rect 20465 -14856 20467 -14822
rect 20505 -14856 20533 -14822
rect 20533 -14856 20539 -14822
rect 20577 -14856 20601 -14822
rect 20601 -14856 20611 -14822
rect 21235 -14856 21245 -14822
rect 21245 -14856 21269 -14822
rect 21307 -14856 21313 -14822
rect 21313 -14856 21341 -14822
rect 21379 -14856 21381 -14822
rect 21381 -14856 21413 -14822
rect 21451 -14856 21483 -14822
rect 21483 -14856 21485 -14822
rect 21523 -14856 21551 -14822
rect 21551 -14856 21557 -14822
rect 21595 -14856 21619 -14822
rect 21619 -14856 21629 -14822
rect 22253 -14856 22263 -14822
rect 22263 -14856 22287 -14822
rect 22325 -14856 22331 -14822
rect 22331 -14856 22359 -14822
rect 22397 -14856 22399 -14822
rect 22399 -14856 22431 -14822
rect 22469 -14856 22501 -14822
rect 22501 -14856 22503 -14822
rect 22541 -14856 22569 -14822
rect 22569 -14856 22575 -14822
rect 22613 -14856 22637 -14822
rect 22637 -14856 22647 -14822
rect 24855 -14831 24889 -14827
rect 24855 -14861 24889 -14831
rect -12289 -14933 -12255 -14899
rect -8855 -14928 -8845 -14894
rect -8845 -14928 -8821 -14894
rect -8783 -14928 -8777 -14894
rect -8777 -14928 -8749 -14894
rect -8711 -14928 -8709 -14894
rect -8709 -14928 -8677 -14894
rect -8639 -14928 -8607 -14894
rect -8607 -14928 -8605 -14894
rect -8567 -14928 -8539 -14894
rect -8539 -14928 -8533 -14894
rect -8495 -14928 -8471 -14894
rect -8471 -14928 -8461 -14894
rect -7837 -14928 -7827 -14894
rect -7827 -14928 -7803 -14894
rect -7765 -14928 -7759 -14894
rect -7759 -14928 -7731 -14894
rect -7693 -14928 -7691 -14894
rect -7691 -14928 -7659 -14894
rect -7621 -14928 -7589 -14894
rect -7589 -14928 -7587 -14894
rect -7549 -14928 -7521 -14894
rect -7521 -14928 -7515 -14894
rect -7477 -14928 -7453 -14894
rect -7453 -14928 -7443 -14894
rect -6819 -14928 -6809 -14894
rect -6809 -14928 -6785 -14894
rect -6747 -14928 -6741 -14894
rect -6741 -14928 -6713 -14894
rect -6675 -14928 -6673 -14894
rect -6673 -14928 -6641 -14894
rect -6603 -14928 -6571 -14894
rect -6571 -14928 -6569 -14894
rect -6531 -14928 -6503 -14894
rect -6503 -14928 -6497 -14894
rect -6459 -14928 -6435 -14894
rect -6435 -14928 -6425 -14894
rect -5801 -14928 -5791 -14894
rect -5791 -14928 -5767 -14894
rect -5729 -14928 -5723 -14894
rect -5723 -14928 -5695 -14894
rect -5657 -14928 -5655 -14894
rect -5655 -14928 -5623 -14894
rect -5585 -14928 -5553 -14894
rect -5553 -14928 -5551 -14894
rect -5513 -14928 -5485 -14894
rect -5485 -14928 -5479 -14894
rect -5441 -14928 -5417 -14894
rect -5417 -14928 -5407 -14894
rect -4783 -14928 -4773 -14894
rect -4773 -14928 -4749 -14894
rect -4711 -14928 -4705 -14894
rect -4705 -14928 -4677 -14894
rect -4639 -14928 -4637 -14894
rect -4637 -14928 -4605 -14894
rect -4567 -14928 -4535 -14894
rect -4535 -14928 -4533 -14894
rect -4495 -14928 -4467 -14894
rect -4467 -14928 -4461 -14894
rect -4423 -14928 -4399 -14894
rect -4399 -14928 -4389 -14894
rect -3765 -14928 -3755 -14894
rect -3755 -14928 -3731 -14894
rect -3693 -14928 -3687 -14894
rect -3687 -14928 -3659 -14894
rect -3621 -14928 -3619 -14894
rect -3619 -14928 -3587 -14894
rect -3549 -14928 -3517 -14894
rect -3517 -14928 -3515 -14894
rect -3477 -14928 -3449 -14894
rect -3449 -14928 -3443 -14894
rect -3405 -14928 -3381 -14894
rect -3381 -14928 -3371 -14894
rect -2747 -14928 -2737 -14894
rect -2737 -14928 -2713 -14894
rect -2675 -14928 -2669 -14894
rect -2669 -14928 -2641 -14894
rect -2603 -14928 -2601 -14894
rect -2601 -14928 -2569 -14894
rect -2531 -14928 -2499 -14894
rect -2499 -14928 -2497 -14894
rect -2459 -14928 -2431 -14894
rect -2431 -14928 -2425 -14894
rect -2387 -14928 -2363 -14894
rect -2363 -14928 -2353 -14894
rect -1729 -14928 -1719 -14894
rect -1719 -14928 -1695 -14894
rect -1657 -14928 -1651 -14894
rect -1651 -14928 -1623 -14894
rect -1585 -14928 -1583 -14894
rect -1583 -14928 -1551 -14894
rect -1513 -14928 -1481 -14894
rect -1481 -14928 -1479 -14894
rect -1441 -14928 -1413 -14894
rect -1413 -14928 -1407 -14894
rect -1369 -14928 -1345 -14894
rect -1345 -14928 -1335 -14894
rect -711 -14928 -701 -14894
rect -701 -14928 -677 -14894
rect -639 -14928 -633 -14894
rect -633 -14928 -605 -14894
rect -567 -14928 -565 -14894
rect -565 -14928 -533 -14894
rect -495 -14928 -463 -14894
rect -463 -14928 -461 -14894
rect -423 -14928 -395 -14894
rect -395 -14928 -389 -14894
rect -351 -14928 -327 -14894
rect -327 -14928 -317 -14894
rect 24855 -14933 24889 -14899
rect -12289 -15001 -12255 -14971
rect -12289 -15005 -12255 -15001
rect -12289 -15069 -12255 -15043
rect -12289 -15077 -12255 -15069
rect -12289 -15137 -12255 -15115
rect -12289 -15149 -12255 -15137
rect -12289 -15205 -12255 -15187
rect -12289 -15221 -12255 -15205
rect -12289 -15273 -12255 -15259
rect -12289 -15293 -12255 -15273
rect -12289 -15341 -12255 -15331
rect -12289 -15365 -12255 -15341
rect -12289 -15409 -12255 -15403
rect -12289 -15437 -12255 -15409
rect -12289 -15477 -12255 -15475
rect -12289 -15509 -12255 -15477
rect -12289 -15579 -12255 -15547
rect -12289 -15581 -12255 -15579
rect -9184 -15011 -9150 -14997
rect -9184 -15031 -9150 -15011
rect -9184 -15079 -9150 -15069
rect -9184 -15103 -9150 -15079
rect -9184 -15147 -9150 -15141
rect -9184 -15175 -9150 -15147
rect -9184 -15215 -9150 -15213
rect -9184 -15247 -9150 -15215
rect -9184 -15317 -9150 -15285
rect -9184 -15319 -9150 -15317
rect -9184 -15385 -9150 -15357
rect -9184 -15391 -9150 -15385
rect -9184 -15453 -9150 -15429
rect -9184 -15463 -9150 -15453
rect -9184 -15521 -9150 -15501
rect -9184 -15535 -9150 -15521
rect -8166 -15011 -8132 -14997
rect -8166 -15031 -8132 -15011
rect -8166 -15079 -8132 -15069
rect -8166 -15103 -8132 -15079
rect -8166 -15147 -8132 -15141
rect -8166 -15175 -8132 -15147
rect -8166 -15215 -8132 -15213
rect -8166 -15247 -8132 -15215
rect -8166 -15317 -8132 -15285
rect -8166 -15319 -8132 -15317
rect -8166 -15385 -8132 -15357
rect -8166 -15391 -8132 -15385
rect -8166 -15453 -8132 -15429
rect -8166 -15463 -8132 -15453
rect -8166 -15521 -8132 -15501
rect -8166 -15535 -8132 -15521
rect -7148 -15011 -7114 -14997
rect -7148 -15031 -7114 -15011
rect -7148 -15079 -7114 -15069
rect -7148 -15103 -7114 -15079
rect -7148 -15147 -7114 -15141
rect -7148 -15175 -7114 -15147
rect -7148 -15215 -7114 -15213
rect -7148 -15247 -7114 -15215
rect -7148 -15317 -7114 -15285
rect -7148 -15319 -7114 -15317
rect -7148 -15385 -7114 -15357
rect -7148 -15391 -7114 -15385
rect -7148 -15453 -7114 -15429
rect -7148 -15463 -7114 -15453
rect -7148 -15521 -7114 -15501
rect -7148 -15535 -7114 -15521
rect -6130 -15011 -6096 -14997
rect -6130 -15031 -6096 -15011
rect -6130 -15079 -6096 -15069
rect -6130 -15103 -6096 -15079
rect -6130 -15147 -6096 -15141
rect -6130 -15175 -6096 -15147
rect -6130 -15215 -6096 -15213
rect -6130 -15247 -6096 -15215
rect -6130 -15317 -6096 -15285
rect -6130 -15319 -6096 -15317
rect -6130 -15385 -6096 -15357
rect -6130 -15391 -6096 -15385
rect -6130 -15453 -6096 -15429
rect -6130 -15463 -6096 -15453
rect -6130 -15521 -6096 -15501
rect -6130 -15535 -6096 -15521
rect -5112 -15011 -5078 -14997
rect -5112 -15031 -5078 -15011
rect -5112 -15079 -5078 -15069
rect -5112 -15103 -5078 -15079
rect -5112 -15147 -5078 -15141
rect -5112 -15175 -5078 -15147
rect -5112 -15215 -5078 -15213
rect -5112 -15247 -5078 -15215
rect -5112 -15317 -5078 -15285
rect -5112 -15319 -5078 -15317
rect -5112 -15385 -5078 -15357
rect -5112 -15391 -5078 -15385
rect -5112 -15453 -5078 -15429
rect -5112 -15463 -5078 -15453
rect -5112 -15521 -5078 -15501
rect -5112 -15535 -5078 -15521
rect -4094 -15011 -4060 -14997
rect -4094 -15031 -4060 -15011
rect -4094 -15079 -4060 -15069
rect -4094 -15103 -4060 -15079
rect -4094 -15147 -4060 -15141
rect -4094 -15175 -4060 -15147
rect -4094 -15215 -4060 -15213
rect -4094 -15247 -4060 -15215
rect -4094 -15317 -4060 -15285
rect -4094 -15319 -4060 -15317
rect -4094 -15385 -4060 -15357
rect -4094 -15391 -4060 -15385
rect -4094 -15453 -4060 -15429
rect -4094 -15463 -4060 -15453
rect -4094 -15521 -4060 -15501
rect -4094 -15535 -4060 -15521
rect -3076 -15011 -3042 -14997
rect -3076 -15031 -3042 -15011
rect -3076 -15079 -3042 -15069
rect -3076 -15103 -3042 -15079
rect -3076 -15147 -3042 -15141
rect -3076 -15175 -3042 -15147
rect -3076 -15215 -3042 -15213
rect -3076 -15247 -3042 -15215
rect -3076 -15317 -3042 -15285
rect -3076 -15319 -3042 -15317
rect -3076 -15385 -3042 -15357
rect -3076 -15391 -3042 -15385
rect -3076 -15453 -3042 -15429
rect -3076 -15463 -3042 -15453
rect -3076 -15521 -3042 -15501
rect -3076 -15535 -3042 -15521
rect -2058 -15011 -2024 -14997
rect -2058 -15031 -2024 -15011
rect -2058 -15079 -2024 -15069
rect -2058 -15103 -2024 -15079
rect -2058 -15147 -2024 -15141
rect -2058 -15175 -2024 -15147
rect -2058 -15215 -2024 -15213
rect -2058 -15247 -2024 -15215
rect -2058 -15317 -2024 -15285
rect -2058 -15319 -2024 -15317
rect -2058 -15385 -2024 -15357
rect -2058 -15391 -2024 -15385
rect -2058 -15453 -2024 -15429
rect -2058 -15463 -2024 -15453
rect -2058 -15521 -2024 -15501
rect -2058 -15535 -2024 -15521
rect -1040 -15011 -1006 -14997
rect -1040 -15031 -1006 -15011
rect -1040 -15079 -1006 -15069
rect -1040 -15103 -1006 -15079
rect -1040 -15147 -1006 -15141
rect -1040 -15175 -1006 -15147
rect -1040 -15215 -1006 -15213
rect -1040 -15247 -1006 -15215
rect -1040 -15317 -1006 -15285
rect -1040 -15319 -1006 -15317
rect -1040 -15385 -1006 -15357
rect -1040 -15391 -1006 -15385
rect -1040 -15453 -1006 -15429
rect -1040 -15463 -1006 -15453
rect -1040 -15521 -1006 -15501
rect -1040 -15535 -1006 -15521
rect -22 -15011 12 -14997
rect -22 -15031 12 -15011
rect -22 -15079 12 -15069
rect -22 -15103 12 -15079
rect -22 -15147 12 -15141
rect -22 -15175 12 -15147
rect -22 -15215 12 -15213
rect -22 -15247 12 -15215
rect -22 -15317 12 -15285
rect -22 -15319 12 -15317
rect 24855 -15001 24889 -14971
rect 24855 -15005 24889 -15001
rect 24855 -15069 24889 -15043
rect 24855 -15077 24889 -15069
rect 24855 -15137 24889 -15115
rect 24855 -15149 24889 -15137
rect 24855 -15205 24889 -15187
rect 24855 -15221 24889 -15205
rect 24855 -15273 24889 -15259
rect 24855 -15293 24889 -15273
rect -22 -15385 12 -15357
rect 2909 -15380 2919 -15346
rect 2919 -15380 2943 -15346
rect 2981 -15380 2987 -15346
rect 2987 -15380 3015 -15346
rect 3053 -15380 3055 -15346
rect 3055 -15380 3087 -15346
rect 3125 -15380 3157 -15346
rect 3157 -15380 3159 -15346
rect 3197 -15380 3225 -15346
rect 3225 -15380 3231 -15346
rect 3269 -15380 3293 -15346
rect 3293 -15380 3303 -15346
rect 3927 -15380 3937 -15346
rect 3937 -15380 3961 -15346
rect 3999 -15380 4005 -15346
rect 4005 -15380 4033 -15346
rect 4071 -15380 4073 -15346
rect 4073 -15380 4105 -15346
rect 4143 -15380 4175 -15346
rect 4175 -15380 4177 -15346
rect 4215 -15380 4243 -15346
rect 4243 -15380 4249 -15346
rect 4287 -15380 4311 -15346
rect 4311 -15380 4321 -15346
rect 4945 -15380 4955 -15346
rect 4955 -15380 4979 -15346
rect 5017 -15380 5023 -15346
rect 5023 -15380 5051 -15346
rect 5089 -15380 5091 -15346
rect 5091 -15380 5123 -15346
rect 5161 -15380 5193 -15346
rect 5193 -15380 5195 -15346
rect 5233 -15380 5261 -15346
rect 5261 -15380 5267 -15346
rect 5305 -15380 5329 -15346
rect 5329 -15380 5339 -15346
rect 5963 -15380 5973 -15346
rect 5973 -15380 5997 -15346
rect 6035 -15380 6041 -15346
rect 6041 -15380 6069 -15346
rect 6107 -15380 6109 -15346
rect 6109 -15380 6141 -15346
rect 6179 -15380 6211 -15346
rect 6211 -15380 6213 -15346
rect 6251 -15380 6279 -15346
rect 6279 -15380 6285 -15346
rect 6323 -15380 6347 -15346
rect 6347 -15380 6357 -15346
rect 6981 -15380 6991 -15346
rect 6991 -15380 7015 -15346
rect 7053 -15380 7059 -15346
rect 7059 -15380 7087 -15346
rect 7125 -15380 7127 -15346
rect 7127 -15380 7159 -15346
rect 7197 -15380 7229 -15346
rect 7229 -15380 7231 -15346
rect 7269 -15380 7297 -15346
rect 7297 -15380 7303 -15346
rect 7341 -15380 7365 -15346
rect 7365 -15380 7375 -15346
rect 7999 -15380 8009 -15346
rect 8009 -15380 8033 -15346
rect 8071 -15380 8077 -15346
rect 8077 -15380 8105 -15346
rect 8143 -15380 8145 -15346
rect 8145 -15380 8177 -15346
rect 8215 -15380 8247 -15346
rect 8247 -15380 8249 -15346
rect 8287 -15380 8315 -15346
rect 8315 -15380 8321 -15346
rect 8359 -15380 8383 -15346
rect 8383 -15380 8393 -15346
rect 9017 -15380 9027 -15346
rect 9027 -15380 9051 -15346
rect 9089 -15380 9095 -15346
rect 9095 -15380 9123 -15346
rect 9161 -15380 9163 -15346
rect 9163 -15380 9195 -15346
rect 9233 -15380 9265 -15346
rect 9265 -15380 9267 -15346
rect 9305 -15380 9333 -15346
rect 9333 -15380 9339 -15346
rect 9377 -15380 9401 -15346
rect 9401 -15380 9411 -15346
rect 10035 -15380 10045 -15346
rect 10045 -15380 10069 -15346
rect 10107 -15380 10113 -15346
rect 10113 -15380 10141 -15346
rect 10179 -15380 10181 -15346
rect 10181 -15380 10213 -15346
rect 10251 -15380 10283 -15346
rect 10283 -15380 10285 -15346
rect 10323 -15380 10351 -15346
rect 10351 -15380 10357 -15346
rect 10395 -15380 10419 -15346
rect 10419 -15380 10429 -15346
rect 11053 -15380 11063 -15346
rect 11063 -15380 11087 -15346
rect 11125 -15380 11131 -15346
rect 11131 -15380 11159 -15346
rect 11197 -15380 11199 -15346
rect 11199 -15380 11231 -15346
rect 11269 -15380 11301 -15346
rect 11301 -15380 11303 -15346
rect 11341 -15380 11369 -15346
rect 11369 -15380 11375 -15346
rect 11413 -15380 11437 -15346
rect 11437 -15380 11447 -15346
rect 12071 -15380 12081 -15346
rect 12081 -15380 12105 -15346
rect 12143 -15380 12149 -15346
rect 12149 -15380 12177 -15346
rect 12215 -15380 12217 -15346
rect 12217 -15380 12249 -15346
rect 12287 -15380 12319 -15346
rect 12319 -15380 12321 -15346
rect 12359 -15380 12387 -15346
rect 12387 -15380 12393 -15346
rect 12431 -15380 12455 -15346
rect 12455 -15380 12465 -15346
rect 13089 -15380 13099 -15346
rect 13099 -15380 13123 -15346
rect 13161 -15380 13167 -15346
rect 13167 -15380 13195 -15346
rect 13233 -15380 13235 -15346
rect 13235 -15380 13267 -15346
rect 13305 -15380 13337 -15346
rect 13337 -15380 13339 -15346
rect 13377 -15380 13405 -15346
rect 13405 -15380 13411 -15346
rect 13449 -15380 13473 -15346
rect 13473 -15380 13483 -15346
rect 14107 -15380 14117 -15346
rect 14117 -15380 14141 -15346
rect 14179 -15380 14185 -15346
rect 14185 -15380 14213 -15346
rect 14251 -15380 14253 -15346
rect 14253 -15380 14285 -15346
rect 14323 -15380 14355 -15346
rect 14355 -15380 14357 -15346
rect 14395 -15380 14423 -15346
rect 14423 -15380 14429 -15346
rect 14467 -15380 14491 -15346
rect 14491 -15380 14501 -15346
rect 15125 -15380 15135 -15346
rect 15135 -15380 15159 -15346
rect 15197 -15380 15203 -15346
rect 15203 -15380 15231 -15346
rect 15269 -15380 15271 -15346
rect 15271 -15380 15303 -15346
rect 15341 -15380 15373 -15346
rect 15373 -15380 15375 -15346
rect 15413 -15380 15441 -15346
rect 15441 -15380 15447 -15346
rect 15485 -15380 15509 -15346
rect 15509 -15380 15519 -15346
rect 16143 -15380 16153 -15346
rect 16153 -15380 16177 -15346
rect 16215 -15380 16221 -15346
rect 16221 -15380 16249 -15346
rect 16287 -15380 16289 -15346
rect 16289 -15380 16321 -15346
rect 16359 -15380 16391 -15346
rect 16391 -15380 16393 -15346
rect 16431 -15380 16459 -15346
rect 16459 -15380 16465 -15346
rect 16503 -15380 16527 -15346
rect 16527 -15380 16537 -15346
rect 17161 -15380 17171 -15346
rect 17171 -15380 17195 -15346
rect 17233 -15380 17239 -15346
rect 17239 -15380 17267 -15346
rect 17305 -15380 17307 -15346
rect 17307 -15380 17339 -15346
rect 17377 -15380 17409 -15346
rect 17409 -15380 17411 -15346
rect 17449 -15380 17477 -15346
rect 17477 -15380 17483 -15346
rect 17521 -15380 17545 -15346
rect 17545 -15380 17555 -15346
rect 18179 -15380 18189 -15346
rect 18189 -15380 18213 -15346
rect 18251 -15380 18257 -15346
rect 18257 -15380 18285 -15346
rect 18323 -15380 18325 -15346
rect 18325 -15380 18357 -15346
rect 18395 -15380 18427 -15346
rect 18427 -15380 18429 -15346
rect 18467 -15380 18495 -15346
rect 18495 -15380 18501 -15346
rect 18539 -15380 18563 -15346
rect 18563 -15380 18573 -15346
rect 19197 -15380 19207 -15346
rect 19207 -15380 19231 -15346
rect 19269 -15380 19275 -15346
rect 19275 -15380 19303 -15346
rect 19341 -15380 19343 -15346
rect 19343 -15380 19375 -15346
rect 19413 -15380 19445 -15346
rect 19445 -15380 19447 -15346
rect 19485 -15380 19513 -15346
rect 19513 -15380 19519 -15346
rect 19557 -15380 19581 -15346
rect 19581 -15380 19591 -15346
rect 20215 -15380 20225 -15346
rect 20225 -15380 20249 -15346
rect 20287 -15380 20293 -15346
rect 20293 -15380 20321 -15346
rect 20359 -15380 20361 -15346
rect 20361 -15380 20393 -15346
rect 20431 -15380 20463 -15346
rect 20463 -15380 20465 -15346
rect 20503 -15380 20531 -15346
rect 20531 -15380 20537 -15346
rect 20575 -15380 20599 -15346
rect 20599 -15380 20609 -15346
rect 21233 -15380 21243 -15346
rect 21243 -15380 21267 -15346
rect 21305 -15380 21311 -15346
rect 21311 -15380 21339 -15346
rect 21377 -15380 21379 -15346
rect 21379 -15380 21411 -15346
rect 21449 -15380 21481 -15346
rect 21481 -15380 21483 -15346
rect 21521 -15380 21549 -15346
rect 21549 -15380 21555 -15346
rect 21593 -15380 21617 -15346
rect 21617 -15380 21627 -15346
rect 22251 -15380 22261 -15346
rect 22261 -15380 22285 -15346
rect 22323 -15380 22329 -15346
rect 22329 -15380 22357 -15346
rect 22395 -15380 22397 -15346
rect 22397 -15380 22429 -15346
rect 22467 -15380 22499 -15346
rect 22499 -15380 22501 -15346
rect 22539 -15380 22567 -15346
rect 22567 -15380 22573 -15346
rect 22611 -15380 22635 -15346
rect 22635 -15380 22645 -15346
rect 24855 -15341 24889 -15331
rect 24855 -15365 24889 -15341
rect -22 -15391 12 -15385
rect -22 -15453 12 -15429
rect -22 -15463 12 -15453
rect -22 -15521 12 -15501
rect -22 -15535 12 -15521
rect 2580 -15463 2614 -15449
rect 2580 -15483 2614 -15463
rect 2580 -15531 2614 -15521
rect 2580 -15555 2614 -15531
rect 2580 -15599 2614 -15593
rect -12289 -15647 -12255 -15619
rect -12289 -15653 -12255 -15647
rect -8855 -15638 -8845 -15604
rect -8845 -15638 -8821 -15604
rect -8783 -15638 -8777 -15604
rect -8777 -15638 -8749 -15604
rect -8711 -15638 -8709 -15604
rect -8709 -15638 -8677 -15604
rect -8639 -15638 -8607 -15604
rect -8607 -15638 -8605 -15604
rect -8567 -15638 -8539 -15604
rect -8539 -15638 -8533 -15604
rect -8495 -15638 -8471 -15604
rect -8471 -15638 -8461 -15604
rect -7837 -15638 -7827 -15604
rect -7827 -15638 -7803 -15604
rect -7765 -15638 -7759 -15604
rect -7759 -15638 -7731 -15604
rect -7693 -15638 -7691 -15604
rect -7691 -15638 -7659 -15604
rect -7621 -15638 -7589 -15604
rect -7589 -15638 -7587 -15604
rect -7549 -15638 -7521 -15604
rect -7521 -15638 -7515 -15604
rect -7477 -15638 -7453 -15604
rect -7453 -15638 -7443 -15604
rect -6819 -15638 -6809 -15604
rect -6809 -15638 -6785 -15604
rect -6747 -15638 -6741 -15604
rect -6741 -15638 -6713 -15604
rect -6675 -15638 -6673 -15604
rect -6673 -15638 -6641 -15604
rect -6603 -15638 -6571 -15604
rect -6571 -15638 -6569 -15604
rect -6531 -15638 -6503 -15604
rect -6503 -15638 -6497 -15604
rect -6459 -15638 -6435 -15604
rect -6435 -15638 -6425 -15604
rect -5801 -15638 -5791 -15604
rect -5791 -15638 -5767 -15604
rect -5729 -15638 -5723 -15604
rect -5723 -15638 -5695 -15604
rect -5657 -15638 -5655 -15604
rect -5655 -15638 -5623 -15604
rect -5585 -15638 -5553 -15604
rect -5553 -15638 -5551 -15604
rect -5513 -15638 -5485 -15604
rect -5485 -15638 -5479 -15604
rect -5441 -15638 -5417 -15604
rect -5417 -15638 -5407 -15604
rect -4783 -15638 -4773 -15604
rect -4773 -15638 -4749 -15604
rect -4711 -15638 -4705 -15604
rect -4705 -15638 -4677 -15604
rect -4639 -15638 -4637 -15604
rect -4637 -15638 -4605 -15604
rect -4567 -15638 -4535 -15604
rect -4535 -15638 -4533 -15604
rect -4495 -15638 -4467 -15604
rect -4467 -15638 -4461 -15604
rect -4423 -15638 -4399 -15604
rect -4399 -15638 -4389 -15604
rect -3765 -15638 -3755 -15604
rect -3755 -15638 -3731 -15604
rect -3693 -15638 -3687 -15604
rect -3687 -15638 -3659 -15604
rect -3621 -15638 -3619 -15604
rect -3619 -15638 -3587 -15604
rect -3549 -15638 -3517 -15604
rect -3517 -15638 -3515 -15604
rect -3477 -15638 -3449 -15604
rect -3449 -15638 -3443 -15604
rect -3405 -15638 -3381 -15604
rect -3381 -15638 -3371 -15604
rect -2747 -15638 -2737 -15604
rect -2737 -15638 -2713 -15604
rect -2675 -15638 -2669 -15604
rect -2669 -15638 -2641 -15604
rect -2603 -15638 -2601 -15604
rect -2601 -15638 -2569 -15604
rect -2531 -15638 -2499 -15604
rect -2499 -15638 -2497 -15604
rect -2459 -15638 -2431 -15604
rect -2431 -15638 -2425 -15604
rect -2387 -15638 -2363 -15604
rect -2363 -15638 -2353 -15604
rect -1729 -15638 -1719 -15604
rect -1719 -15638 -1695 -15604
rect -1657 -15638 -1651 -15604
rect -1651 -15638 -1623 -15604
rect -1585 -15638 -1583 -15604
rect -1583 -15638 -1551 -15604
rect -1513 -15638 -1481 -15604
rect -1481 -15638 -1479 -15604
rect -1441 -15638 -1413 -15604
rect -1413 -15638 -1407 -15604
rect -1369 -15638 -1345 -15604
rect -1345 -15638 -1335 -15604
rect -711 -15638 -701 -15604
rect -701 -15638 -677 -15604
rect -639 -15638 -633 -15604
rect -633 -15638 -605 -15604
rect -567 -15638 -565 -15604
rect -565 -15638 -533 -15604
rect -495 -15638 -463 -15604
rect -463 -15638 -461 -15604
rect -423 -15638 -395 -15604
rect -395 -15638 -389 -15604
rect -351 -15638 -327 -15604
rect -327 -15638 -317 -15604
rect 2580 -15627 2614 -15599
rect -12289 -15715 -12255 -15691
rect -12289 -15725 -12255 -15715
rect 2580 -15667 2614 -15665
rect 2580 -15699 2614 -15667
rect -8855 -15746 -8845 -15712
rect -8845 -15746 -8821 -15712
rect -8783 -15746 -8777 -15712
rect -8777 -15746 -8749 -15712
rect -8711 -15746 -8709 -15712
rect -8709 -15746 -8677 -15712
rect -8639 -15746 -8607 -15712
rect -8607 -15746 -8605 -15712
rect -8567 -15746 -8539 -15712
rect -8539 -15746 -8533 -15712
rect -8495 -15746 -8471 -15712
rect -8471 -15746 -8461 -15712
rect -7837 -15746 -7827 -15712
rect -7827 -15746 -7803 -15712
rect -7765 -15746 -7759 -15712
rect -7759 -15746 -7731 -15712
rect -7693 -15746 -7691 -15712
rect -7691 -15746 -7659 -15712
rect -7621 -15746 -7589 -15712
rect -7589 -15746 -7587 -15712
rect -7549 -15746 -7521 -15712
rect -7521 -15746 -7515 -15712
rect -7477 -15746 -7453 -15712
rect -7453 -15746 -7443 -15712
rect -6819 -15746 -6809 -15712
rect -6809 -15746 -6785 -15712
rect -6747 -15746 -6741 -15712
rect -6741 -15746 -6713 -15712
rect -6675 -15746 -6673 -15712
rect -6673 -15746 -6641 -15712
rect -6603 -15746 -6571 -15712
rect -6571 -15746 -6569 -15712
rect -6531 -15746 -6503 -15712
rect -6503 -15746 -6497 -15712
rect -6459 -15746 -6435 -15712
rect -6435 -15746 -6425 -15712
rect -5801 -15746 -5791 -15712
rect -5791 -15746 -5767 -15712
rect -5729 -15746 -5723 -15712
rect -5723 -15746 -5695 -15712
rect -5657 -15746 -5655 -15712
rect -5655 -15746 -5623 -15712
rect -5585 -15746 -5553 -15712
rect -5553 -15746 -5551 -15712
rect -5513 -15746 -5485 -15712
rect -5485 -15746 -5479 -15712
rect -5441 -15746 -5417 -15712
rect -5417 -15746 -5407 -15712
rect -4783 -15746 -4773 -15712
rect -4773 -15746 -4749 -15712
rect -4711 -15746 -4705 -15712
rect -4705 -15746 -4677 -15712
rect -4639 -15746 -4637 -15712
rect -4637 -15746 -4605 -15712
rect -4567 -15746 -4535 -15712
rect -4535 -15746 -4533 -15712
rect -4495 -15746 -4467 -15712
rect -4467 -15746 -4461 -15712
rect -4423 -15746 -4399 -15712
rect -4399 -15746 -4389 -15712
rect -3765 -15746 -3755 -15712
rect -3755 -15746 -3731 -15712
rect -3693 -15746 -3687 -15712
rect -3687 -15746 -3659 -15712
rect -3621 -15746 -3619 -15712
rect -3619 -15746 -3587 -15712
rect -3549 -15746 -3517 -15712
rect -3517 -15746 -3515 -15712
rect -3477 -15746 -3449 -15712
rect -3449 -15746 -3443 -15712
rect -3405 -15746 -3381 -15712
rect -3381 -15746 -3371 -15712
rect -2747 -15746 -2737 -15712
rect -2737 -15746 -2713 -15712
rect -2675 -15746 -2669 -15712
rect -2669 -15746 -2641 -15712
rect -2603 -15746 -2601 -15712
rect -2601 -15746 -2569 -15712
rect -2531 -15746 -2499 -15712
rect -2499 -15746 -2497 -15712
rect -2459 -15746 -2431 -15712
rect -2431 -15746 -2425 -15712
rect -2387 -15746 -2363 -15712
rect -2363 -15746 -2353 -15712
rect -1729 -15746 -1719 -15712
rect -1719 -15746 -1695 -15712
rect -1657 -15746 -1651 -15712
rect -1651 -15746 -1623 -15712
rect -1585 -15746 -1583 -15712
rect -1583 -15746 -1551 -15712
rect -1513 -15746 -1481 -15712
rect -1481 -15746 -1479 -15712
rect -1441 -15746 -1413 -15712
rect -1413 -15746 -1407 -15712
rect -1369 -15746 -1345 -15712
rect -1345 -15746 -1335 -15712
rect -711 -15746 -701 -15712
rect -701 -15746 -677 -15712
rect -639 -15746 -633 -15712
rect -633 -15746 -605 -15712
rect -567 -15746 -565 -15712
rect -565 -15746 -533 -15712
rect -495 -15746 -463 -15712
rect -463 -15746 -461 -15712
rect -423 -15746 -395 -15712
rect -395 -15746 -389 -15712
rect -351 -15746 -327 -15712
rect -327 -15746 -317 -15712
rect -12289 -15783 -12255 -15763
rect -12289 -15797 -12255 -15783
rect 2580 -15769 2614 -15737
rect 2580 -15771 2614 -15769
rect -12289 -15851 -12255 -15835
rect -12289 -15869 -12255 -15851
rect -12289 -15919 -12255 -15907
rect -12289 -15941 -12255 -15919
rect -12289 -15987 -12255 -15979
rect -12289 -16013 -12255 -15987
rect -12289 -16055 -12255 -16051
rect -12289 -16085 -12255 -16055
rect -12289 -16157 -12255 -16123
rect -12289 -16225 -12255 -16195
rect -12289 -16229 -12255 -16225
rect -12289 -16293 -12255 -16267
rect -12289 -16301 -12255 -16293
rect -12289 -16361 -12255 -16339
rect -12289 -16373 -12255 -16361
rect -9184 -15829 -9150 -15815
rect -9184 -15849 -9150 -15829
rect -9184 -15897 -9150 -15887
rect -9184 -15921 -9150 -15897
rect -9184 -15965 -9150 -15959
rect -9184 -15993 -9150 -15965
rect -9184 -16033 -9150 -16031
rect -9184 -16065 -9150 -16033
rect -9184 -16135 -9150 -16103
rect -9184 -16137 -9150 -16135
rect -9184 -16203 -9150 -16175
rect -9184 -16209 -9150 -16203
rect -9184 -16271 -9150 -16247
rect -9184 -16281 -9150 -16271
rect -9184 -16339 -9150 -16319
rect -9184 -16353 -9150 -16339
rect -8166 -15829 -8132 -15815
rect -8166 -15849 -8132 -15829
rect -8166 -15897 -8132 -15887
rect -8166 -15921 -8132 -15897
rect -8166 -15965 -8132 -15959
rect -8166 -15993 -8132 -15965
rect -8166 -16033 -8132 -16031
rect -8166 -16065 -8132 -16033
rect -8166 -16135 -8132 -16103
rect -8166 -16137 -8132 -16135
rect -8166 -16203 -8132 -16175
rect -8166 -16209 -8132 -16203
rect -8166 -16271 -8132 -16247
rect -8166 -16281 -8132 -16271
rect -8166 -16339 -8132 -16319
rect -8166 -16353 -8132 -16339
rect -7148 -15829 -7114 -15815
rect -7148 -15849 -7114 -15829
rect -7148 -15897 -7114 -15887
rect -7148 -15921 -7114 -15897
rect -7148 -15965 -7114 -15959
rect -7148 -15993 -7114 -15965
rect -7148 -16033 -7114 -16031
rect -7148 -16065 -7114 -16033
rect -7148 -16135 -7114 -16103
rect -7148 -16137 -7114 -16135
rect -7148 -16203 -7114 -16175
rect -7148 -16209 -7114 -16203
rect -7148 -16271 -7114 -16247
rect -7148 -16281 -7114 -16271
rect -7148 -16339 -7114 -16319
rect -7148 -16353 -7114 -16339
rect -6130 -15829 -6096 -15815
rect -6130 -15849 -6096 -15829
rect -6130 -15897 -6096 -15887
rect -6130 -15921 -6096 -15897
rect -6130 -15965 -6096 -15959
rect -6130 -15993 -6096 -15965
rect -6130 -16033 -6096 -16031
rect -6130 -16065 -6096 -16033
rect -6130 -16135 -6096 -16103
rect -6130 -16137 -6096 -16135
rect -6130 -16203 -6096 -16175
rect -6130 -16209 -6096 -16203
rect -6130 -16271 -6096 -16247
rect -6130 -16281 -6096 -16271
rect -6130 -16339 -6096 -16319
rect -6130 -16353 -6096 -16339
rect -5112 -15829 -5078 -15815
rect -5112 -15849 -5078 -15829
rect -5112 -15897 -5078 -15887
rect -5112 -15921 -5078 -15897
rect -5112 -15965 -5078 -15959
rect -5112 -15993 -5078 -15965
rect -5112 -16033 -5078 -16031
rect -5112 -16065 -5078 -16033
rect -5112 -16135 -5078 -16103
rect -5112 -16137 -5078 -16135
rect -5112 -16203 -5078 -16175
rect -5112 -16209 -5078 -16203
rect -5112 -16271 -5078 -16247
rect -5112 -16281 -5078 -16271
rect -5112 -16339 -5078 -16319
rect -5112 -16353 -5078 -16339
rect -4094 -15829 -4060 -15815
rect -4094 -15849 -4060 -15829
rect -4094 -15897 -4060 -15887
rect -4094 -15921 -4060 -15897
rect -4094 -15965 -4060 -15959
rect -4094 -15993 -4060 -15965
rect -4094 -16033 -4060 -16031
rect -4094 -16065 -4060 -16033
rect -4094 -16135 -4060 -16103
rect -4094 -16137 -4060 -16135
rect -4094 -16203 -4060 -16175
rect -4094 -16209 -4060 -16203
rect -4094 -16271 -4060 -16247
rect -4094 -16281 -4060 -16271
rect -4094 -16339 -4060 -16319
rect -4094 -16353 -4060 -16339
rect -3076 -15829 -3042 -15815
rect -3076 -15849 -3042 -15829
rect -3076 -15897 -3042 -15887
rect -3076 -15921 -3042 -15897
rect -3076 -15965 -3042 -15959
rect -3076 -15993 -3042 -15965
rect -3076 -16033 -3042 -16031
rect -3076 -16065 -3042 -16033
rect -3076 -16135 -3042 -16103
rect -3076 -16137 -3042 -16135
rect -3076 -16203 -3042 -16175
rect -3076 -16209 -3042 -16203
rect -3076 -16271 -3042 -16247
rect -3076 -16281 -3042 -16271
rect -3076 -16339 -3042 -16319
rect -3076 -16353 -3042 -16339
rect -2058 -15829 -2024 -15815
rect -2058 -15849 -2024 -15829
rect -2058 -15897 -2024 -15887
rect -2058 -15921 -2024 -15897
rect -2058 -15965 -2024 -15959
rect -2058 -15993 -2024 -15965
rect -2058 -16033 -2024 -16031
rect -2058 -16065 -2024 -16033
rect -2058 -16135 -2024 -16103
rect -2058 -16137 -2024 -16135
rect -2058 -16203 -2024 -16175
rect -2058 -16209 -2024 -16203
rect -2058 -16271 -2024 -16247
rect -2058 -16281 -2024 -16271
rect -2058 -16339 -2024 -16319
rect -2058 -16353 -2024 -16339
rect -1040 -15829 -1006 -15815
rect -1040 -15849 -1006 -15829
rect -1040 -15897 -1006 -15887
rect -1040 -15921 -1006 -15897
rect -1040 -15965 -1006 -15959
rect -1040 -15993 -1006 -15965
rect -1040 -16033 -1006 -16031
rect -1040 -16065 -1006 -16033
rect -1040 -16135 -1006 -16103
rect -1040 -16137 -1006 -16135
rect -1040 -16203 -1006 -16175
rect -1040 -16209 -1006 -16203
rect -1040 -16271 -1006 -16247
rect -1040 -16281 -1006 -16271
rect -1040 -16339 -1006 -16319
rect -1040 -16353 -1006 -16339
rect -22 -15829 12 -15815
rect -22 -15849 12 -15829
rect -22 -15897 12 -15887
rect -22 -15921 12 -15897
rect -22 -15965 12 -15959
rect -22 -15993 12 -15965
rect 2580 -15837 2614 -15809
rect 2580 -15843 2614 -15837
rect 2580 -15905 2614 -15881
rect 2580 -15915 2614 -15905
rect 2580 -15973 2614 -15953
rect 2580 -15987 2614 -15973
rect 3598 -15463 3632 -15449
rect 3598 -15483 3632 -15463
rect 3598 -15531 3632 -15521
rect 3598 -15555 3632 -15531
rect 3598 -15599 3632 -15593
rect 3598 -15627 3632 -15599
rect 3598 -15667 3632 -15665
rect 3598 -15699 3632 -15667
rect 3598 -15769 3632 -15737
rect 3598 -15771 3632 -15769
rect 3598 -15837 3632 -15809
rect 3598 -15843 3632 -15837
rect 3598 -15905 3632 -15881
rect 3598 -15915 3632 -15905
rect 3598 -15973 3632 -15953
rect 3598 -15987 3632 -15973
rect 4616 -15463 4650 -15449
rect 4616 -15483 4650 -15463
rect 4616 -15531 4650 -15521
rect 4616 -15555 4650 -15531
rect 4616 -15599 4650 -15593
rect 4616 -15627 4650 -15599
rect 4616 -15667 4650 -15665
rect 4616 -15699 4650 -15667
rect 4616 -15769 4650 -15737
rect 4616 -15771 4650 -15769
rect 4616 -15837 4650 -15809
rect 4616 -15843 4650 -15837
rect 4616 -15905 4650 -15881
rect 4616 -15915 4650 -15905
rect 4616 -15973 4650 -15953
rect 4616 -15987 4650 -15973
rect 5634 -15463 5668 -15449
rect 5634 -15483 5668 -15463
rect 5634 -15531 5668 -15521
rect 5634 -15555 5668 -15531
rect 5634 -15599 5668 -15593
rect 5634 -15627 5668 -15599
rect 5634 -15667 5668 -15665
rect 5634 -15699 5668 -15667
rect 5634 -15769 5668 -15737
rect 5634 -15771 5668 -15769
rect 5634 -15837 5668 -15809
rect 5634 -15843 5668 -15837
rect 5634 -15905 5668 -15881
rect 5634 -15915 5668 -15905
rect 5634 -15973 5668 -15953
rect 5634 -15987 5668 -15973
rect 6652 -15463 6686 -15449
rect 6652 -15483 6686 -15463
rect 6652 -15531 6686 -15521
rect 6652 -15555 6686 -15531
rect 6652 -15599 6686 -15593
rect 6652 -15627 6686 -15599
rect 6652 -15667 6686 -15665
rect 6652 -15699 6686 -15667
rect 6652 -15769 6686 -15737
rect 6652 -15771 6686 -15769
rect 6652 -15837 6686 -15809
rect 6652 -15843 6686 -15837
rect 6652 -15905 6686 -15881
rect 6652 -15915 6686 -15905
rect 6652 -15973 6686 -15953
rect 6652 -15987 6686 -15973
rect 7670 -15463 7704 -15449
rect 7670 -15483 7704 -15463
rect 7670 -15531 7704 -15521
rect 7670 -15555 7704 -15531
rect 7670 -15599 7704 -15593
rect 7670 -15627 7704 -15599
rect 7670 -15667 7704 -15665
rect 7670 -15699 7704 -15667
rect 7670 -15769 7704 -15737
rect 7670 -15771 7704 -15769
rect 7670 -15837 7704 -15809
rect 7670 -15843 7704 -15837
rect 7670 -15905 7704 -15881
rect 7670 -15915 7704 -15905
rect 7670 -15973 7704 -15953
rect 7670 -15987 7704 -15973
rect 8688 -15463 8722 -15449
rect 8688 -15483 8722 -15463
rect 8688 -15531 8722 -15521
rect 8688 -15555 8722 -15531
rect 8688 -15599 8722 -15593
rect 8688 -15627 8722 -15599
rect 8688 -15667 8722 -15665
rect 8688 -15699 8722 -15667
rect 8688 -15769 8722 -15737
rect 8688 -15771 8722 -15769
rect 8688 -15837 8722 -15809
rect 8688 -15843 8722 -15837
rect 8688 -15905 8722 -15881
rect 8688 -15915 8722 -15905
rect 8688 -15973 8722 -15953
rect 8688 -15987 8722 -15973
rect 9706 -15463 9740 -15449
rect 9706 -15483 9740 -15463
rect 9706 -15531 9740 -15521
rect 9706 -15555 9740 -15531
rect 9706 -15599 9740 -15593
rect 9706 -15627 9740 -15599
rect 9706 -15667 9740 -15665
rect 9706 -15699 9740 -15667
rect 9706 -15769 9740 -15737
rect 9706 -15771 9740 -15769
rect 9706 -15837 9740 -15809
rect 9706 -15843 9740 -15837
rect 9706 -15905 9740 -15881
rect 9706 -15915 9740 -15905
rect 9706 -15973 9740 -15953
rect 9706 -15987 9740 -15973
rect 10724 -15463 10758 -15449
rect 10724 -15483 10758 -15463
rect 10724 -15531 10758 -15521
rect 10724 -15555 10758 -15531
rect 10724 -15599 10758 -15593
rect 10724 -15627 10758 -15599
rect 10724 -15667 10758 -15665
rect 10724 -15699 10758 -15667
rect 10724 -15769 10758 -15737
rect 10724 -15771 10758 -15769
rect 10724 -15837 10758 -15809
rect 10724 -15843 10758 -15837
rect 10724 -15905 10758 -15881
rect 10724 -15915 10758 -15905
rect 10724 -15973 10758 -15953
rect 10724 -15987 10758 -15973
rect 11742 -15463 11776 -15449
rect 11742 -15483 11776 -15463
rect 11742 -15531 11776 -15521
rect 11742 -15555 11776 -15531
rect 11742 -15599 11776 -15593
rect 11742 -15627 11776 -15599
rect 11742 -15667 11776 -15665
rect 11742 -15699 11776 -15667
rect 11742 -15769 11776 -15737
rect 11742 -15771 11776 -15769
rect 11742 -15837 11776 -15809
rect 11742 -15843 11776 -15837
rect 11742 -15905 11776 -15881
rect 11742 -15915 11776 -15905
rect 11742 -15973 11776 -15953
rect 11742 -15987 11776 -15973
rect 12760 -15463 12794 -15449
rect 12760 -15483 12794 -15463
rect 12760 -15531 12794 -15521
rect 12760 -15555 12794 -15531
rect 12760 -15599 12794 -15593
rect 12760 -15627 12794 -15599
rect 12760 -15667 12794 -15665
rect 12760 -15699 12794 -15667
rect 12760 -15769 12794 -15737
rect 12760 -15771 12794 -15769
rect 12760 -15837 12794 -15809
rect 12760 -15843 12794 -15837
rect 12760 -15905 12794 -15881
rect 12760 -15915 12794 -15905
rect 12760 -15973 12794 -15953
rect 12760 -15987 12794 -15973
rect 13778 -15463 13812 -15449
rect 13778 -15483 13812 -15463
rect 13778 -15531 13812 -15521
rect 13778 -15555 13812 -15531
rect 13778 -15599 13812 -15593
rect 13778 -15627 13812 -15599
rect 13778 -15667 13812 -15665
rect 13778 -15699 13812 -15667
rect 13778 -15769 13812 -15737
rect 13778 -15771 13812 -15769
rect 13778 -15837 13812 -15809
rect 13778 -15843 13812 -15837
rect 13778 -15905 13812 -15881
rect 13778 -15915 13812 -15905
rect 13778 -15973 13812 -15953
rect 13778 -15987 13812 -15973
rect 14796 -15463 14830 -15449
rect 14796 -15483 14830 -15463
rect 14796 -15531 14830 -15521
rect 14796 -15555 14830 -15531
rect 14796 -15599 14830 -15593
rect 14796 -15627 14830 -15599
rect 14796 -15667 14830 -15665
rect 14796 -15699 14830 -15667
rect 14796 -15769 14830 -15737
rect 14796 -15771 14830 -15769
rect 14796 -15837 14830 -15809
rect 14796 -15843 14830 -15837
rect 14796 -15905 14830 -15881
rect 14796 -15915 14830 -15905
rect 14796 -15973 14830 -15953
rect 14796 -15987 14830 -15973
rect 15814 -15463 15848 -15449
rect 15814 -15483 15848 -15463
rect 15814 -15531 15848 -15521
rect 15814 -15555 15848 -15531
rect 15814 -15599 15848 -15593
rect 15814 -15627 15848 -15599
rect 15814 -15667 15848 -15665
rect 15814 -15699 15848 -15667
rect 15814 -15769 15848 -15737
rect 15814 -15771 15848 -15769
rect 15814 -15837 15848 -15809
rect 15814 -15843 15848 -15837
rect 15814 -15905 15848 -15881
rect 15814 -15915 15848 -15905
rect 15814 -15973 15848 -15953
rect 15814 -15987 15848 -15973
rect 16832 -15463 16866 -15449
rect 16832 -15483 16866 -15463
rect 16832 -15531 16866 -15521
rect 16832 -15555 16866 -15531
rect 16832 -15599 16866 -15593
rect 16832 -15627 16866 -15599
rect 16832 -15667 16866 -15665
rect 16832 -15699 16866 -15667
rect 16832 -15769 16866 -15737
rect 16832 -15771 16866 -15769
rect 16832 -15837 16866 -15809
rect 16832 -15843 16866 -15837
rect 16832 -15905 16866 -15881
rect 16832 -15915 16866 -15905
rect 16832 -15973 16866 -15953
rect 16832 -15987 16866 -15973
rect 17850 -15463 17884 -15449
rect 17850 -15483 17884 -15463
rect 17850 -15531 17884 -15521
rect 17850 -15555 17884 -15531
rect 17850 -15599 17884 -15593
rect 17850 -15627 17884 -15599
rect 17850 -15667 17884 -15665
rect 17850 -15699 17884 -15667
rect 17850 -15769 17884 -15737
rect 17850 -15771 17884 -15769
rect 17850 -15837 17884 -15809
rect 17850 -15843 17884 -15837
rect 17850 -15905 17884 -15881
rect 17850 -15915 17884 -15905
rect 17850 -15973 17884 -15953
rect 17850 -15987 17884 -15973
rect 18868 -15463 18902 -15449
rect 18868 -15483 18902 -15463
rect 18868 -15531 18902 -15521
rect 18868 -15555 18902 -15531
rect 18868 -15599 18902 -15593
rect 18868 -15627 18902 -15599
rect 18868 -15667 18902 -15665
rect 18868 -15699 18902 -15667
rect 18868 -15769 18902 -15737
rect 18868 -15771 18902 -15769
rect 18868 -15837 18902 -15809
rect 18868 -15843 18902 -15837
rect 18868 -15905 18902 -15881
rect 18868 -15915 18902 -15905
rect 18868 -15973 18902 -15953
rect 18868 -15987 18902 -15973
rect 19886 -15463 19920 -15449
rect 19886 -15483 19920 -15463
rect 19886 -15531 19920 -15521
rect 19886 -15555 19920 -15531
rect 19886 -15599 19920 -15593
rect 19886 -15627 19920 -15599
rect 19886 -15667 19920 -15665
rect 19886 -15699 19920 -15667
rect 19886 -15769 19920 -15737
rect 19886 -15771 19920 -15769
rect 19886 -15837 19920 -15809
rect 19886 -15843 19920 -15837
rect 19886 -15905 19920 -15881
rect 19886 -15915 19920 -15905
rect 19886 -15973 19920 -15953
rect 19886 -15987 19920 -15973
rect 20904 -15463 20938 -15449
rect 20904 -15483 20938 -15463
rect 20904 -15531 20938 -15521
rect 20904 -15555 20938 -15531
rect 20904 -15599 20938 -15593
rect 20904 -15627 20938 -15599
rect 20904 -15667 20938 -15665
rect 20904 -15699 20938 -15667
rect 20904 -15769 20938 -15737
rect 20904 -15771 20938 -15769
rect 20904 -15837 20938 -15809
rect 20904 -15843 20938 -15837
rect 20904 -15905 20938 -15881
rect 20904 -15915 20938 -15905
rect 20904 -15973 20938 -15953
rect 20904 -15987 20938 -15973
rect 21922 -15463 21956 -15449
rect 21922 -15483 21956 -15463
rect 21922 -15531 21956 -15521
rect 21922 -15555 21956 -15531
rect 21922 -15599 21956 -15593
rect 21922 -15627 21956 -15599
rect 21922 -15667 21956 -15665
rect 21922 -15699 21956 -15667
rect 21922 -15769 21956 -15737
rect 21922 -15771 21956 -15769
rect 21922 -15837 21956 -15809
rect 21922 -15843 21956 -15837
rect 21922 -15905 21956 -15881
rect 21922 -15915 21956 -15905
rect 21922 -15973 21956 -15953
rect 21922 -15987 21956 -15973
rect 22940 -15463 22974 -15449
rect 22940 -15483 22974 -15463
rect 22940 -15531 22974 -15521
rect 22940 -15555 22974 -15531
rect 22940 -15599 22974 -15593
rect 22940 -15627 22974 -15599
rect 22940 -15667 22974 -15665
rect 22940 -15699 22974 -15667
rect 22940 -15769 22974 -15737
rect 22940 -15771 22974 -15769
rect 22940 -15837 22974 -15809
rect 22940 -15843 22974 -15837
rect 22940 -15905 22974 -15881
rect 22940 -15915 22974 -15905
rect 22940 -15973 22974 -15953
rect 22940 -15987 22974 -15973
rect 24855 -15409 24889 -15403
rect 24855 -15437 24889 -15409
rect 24855 -15477 24889 -15475
rect 24855 -15509 24889 -15477
rect 24855 -15579 24889 -15547
rect 24855 -15581 24889 -15579
rect 24855 -15647 24889 -15619
rect 24855 -15653 24889 -15647
rect 24855 -15715 24889 -15691
rect 24855 -15725 24889 -15715
rect 24855 -15783 24889 -15763
rect 24855 -15797 24889 -15783
rect 24855 -15851 24889 -15835
rect 24855 -15869 24889 -15851
rect 24855 -15919 24889 -15907
rect 24855 -15941 24889 -15919
rect 24855 -15987 24889 -15979
rect 24855 -16013 24889 -15987
rect -22 -16033 12 -16031
rect -22 -16065 12 -16033
rect 2909 -16090 2919 -16056
rect 2919 -16090 2943 -16056
rect 2981 -16090 2987 -16056
rect 2987 -16090 3015 -16056
rect 3053 -16090 3055 -16056
rect 3055 -16090 3087 -16056
rect 3125 -16090 3157 -16056
rect 3157 -16090 3159 -16056
rect 3197 -16090 3225 -16056
rect 3225 -16090 3231 -16056
rect 3269 -16090 3293 -16056
rect 3293 -16090 3303 -16056
rect 3927 -16090 3937 -16056
rect 3937 -16090 3961 -16056
rect 3999 -16090 4005 -16056
rect 4005 -16090 4033 -16056
rect 4071 -16090 4073 -16056
rect 4073 -16090 4105 -16056
rect 4143 -16090 4175 -16056
rect 4175 -16090 4177 -16056
rect 4215 -16090 4243 -16056
rect 4243 -16090 4249 -16056
rect 4287 -16090 4311 -16056
rect 4311 -16090 4321 -16056
rect 4945 -16090 4955 -16056
rect 4955 -16090 4979 -16056
rect 5017 -16090 5023 -16056
rect 5023 -16090 5051 -16056
rect 5089 -16090 5091 -16056
rect 5091 -16090 5123 -16056
rect 5161 -16090 5193 -16056
rect 5193 -16090 5195 -16056
rect 5233 -16090 5261 -16056
rect 5261 -16090 5267 -16056
rect 5305 -16090 5329 -16056
rect 5329 -16090 5339 -16056
rect 5963 -16090 5973 -16056
rect 5973 -16090 5997 -16056
rect 6035 -16090 6041 -16056
rect 6041 -16090 6069 -16056
rect 6107 -16090 6109 -16056
rect 6109 -16090 6141 -16056
rect 6179 -16090 6211 -16056
rect 6211 -16090 6213 -16056
rect 6251 -16090 6279 -16056
rect 6279 -16090 6285 -16056
rect 6323 -16090 6347 -16056
rect 6347 -16090 6357 -16056
rect 6981 -16090 6991 -16056
rect 6991 -16090 7015 -16056
rect 7053 -16090 7059 -16056
rect 7059 -16090 7087 -16056
rect 7125 -16090 7127 -16056
rect 7127 -16090 7159 -16056
rect 7197 -16090 7229 -16056
rect 7229 -16090 7231 -16056
rect 7269 -16090 7297 -16056
rect 7297 -16090 7303 -16056
rect 7341 -16090 7365 -16056
rect 7365 -16090 7375 -16056
rect 7999 -16090 8009 -16056
rect 8009 -16090 8033 -16056
rect 8071 -16090 8077 -16056
rect 8077 -16090 8105 -16056
rect 8143 -16090 8145 -16056
rect 8145 -16090 8177 -16056
rect 8215 -16090 8247 -16056
rect 8247 -16090 8249 -16056
rect 8287 -16090 8315 -16056
rect 8315 -16090 8321 -16056
rect 8359 -16090 8383 -16056
rect 8383 -16090 8393 -16056
rect 9017 -16090 9027 -16056
rect 9027 -16090 9051 -16056
rect 9089 -16090 9095 -16056
rect 9095 -16090 9123 -16056
rect 9161 -16090 9163 -16056
rect 9163 -16090 9195 -16056
rect 9233 -16090 9265 -16056
rect 9265 -16090 9267 -16056
rect 9305 -16090 9333 -16056
rect 9333 -16090 9339 -16056
rect 9377 -16090 9401 -16056
rect 9401 -16090 9411 -16056
rect 10035 -16090 10045 -16056
rect 10045 -16090 10069 -16056
rect 10107 -16090 10113 -16056
rect 10113 -16090 10141 -16056
rect 10179 -16090 10181 -16056
rect 10181 -16090 10213 -16056
rect 10251 -16090 10283 -16056
rect 10283 -16090 10285 -16056
rect 10323 -16090 10351 -16056
rect 10351 -16090 10357 -16056
rect 10395 -16090 10419 -16056
rect 10419 -16090 10429 -16056
rect 11053 -16090 11063 -16056
rect 11063 -16090 11087 -16056
rect 11125 -16090 11131 -16056
rect 11131 -16090 11159 -16056
rect 11197 -16090 11199 -16056
rect 11199 -16090 11231 -16056
rect 11269 -16090 11301 -16056
rect 11301 -16090 11303 -16056
rect 11341 -16090 11369 -16056
rect 11369 -16090 11375 -16056
rect 11413 -16090 11437 -16056
rect 11437 -16090 11447 -16056
rect 12071 -16090 12081 -16056
rect 12081 -16090 12105 -16056
rect 12143 -16090 12149 -16056
rect 12149 -16090 12177 -16056
rect 12215 -16090 12217 -16056
rect 12217 -16090 12249 -16056
rect 12287 -16090 12319 -16056
rect 12319 -16090 12321 -16056
rect 12359 -16090 12387 -16056
rect 12387 -16090 12393 -16056
rect 12431 -16090 12455 -16056
rect 12455 -16090 12465 -16056
rect 13089 -16090 13099 -16056
rect 13099 -16090 13123 -16056
rect 13161 -16090 13167 -16056
rect 13167 -16090 13195 -16056
rect 13233 -16090 13235 -16056
rect 13235 -16090 13267 -16056
rect 13305 -16090 13337 -16056
rect 13337 -16090 13339 -16056
rect 13377 -16090 13405 -16056
rect 13405 -16090 13411 -16056
rect 13449 -16090 13473 -16056
rect 13473 -16090 13483 -16056
rect 14107 -16090 14117 -16056
rect 14117 -16090 14141 -16056
rect 14179 -16090 14185 -16056
rect 14185 -16090 14213 -16056
rect 14251 -16090 14253 -16056
rect 14253 -16090 14285 -16056
rect 14323 -16090 14355 -16056
rect 14355 -16090 14357 -16056
rect 14395 -16090 14423 -16056
rect 14423 -16090 14429 -16056
rect 14467 -16090 14491 -16056
rect 14491 -16090 14501 -16056
rect 15125 -16090 15135 -16056
rect 15135 -16090 15159 -16056
rect 15197 -16090 15203 -16056
rect 15203 -16090 15231 -16056
rect 15269 -16090 15271 -16056
rect 15271 -16090 15303 -16056
rect 15341 -16090 15373 -16056
rect 15373 -16090 15375 -16056
rect 15413 -16090 15441 -16056
rect 15441 -16090 15447 -16056
rect 15485 -16090 15509 -16056
rect 15509 -16090 15519 -16056
rect 16143 -16090 16153 -16056
rect 16153 -16090 16177 -16056
rect 16215 -16090 16221 -16056
rect 16221 -16090 16249 -16056
rect 16287 -16090 16289 -16056
rect 16289 -16090 16321 -16056
rect 16359 -16090 16391 -16056
rect 16391 -16090 16393 -16056
rect 16431 -16090 16459 -16056
rect 16459 -16090 16465 -16056
rect 16503 -16090 16527 -16056
rect 16527 -16090 16537 -16056
rect 17161 -16090 17171 -16056
rect 17171 -16090 17195 -16056
rect 17233 -16090 17239 -16056
rect 17239 -16090 17267 -16056
rect 17305 -16090 17307 -16056
rect 17307 -16090 17339 -16056
rect 17377 -16090 17409 -16056
rect 17409 -16090 17411 -16056
rect 17449 -16090 17477 -16056
rect 17477 -16090 17483 -16056
rect 17521 -16090 17545 -16056
rect 17545 -16090 17555 -16056
rect 18179 -16090 18189 -16056
rect 18189 -16090 18213 -16056
rect 18251 -16090 18257 -16056
rect 18257 -16090 18285 -16056
rect 18323 -16090 18325 -16056
rect 18325 -16090 18357 -16056
rect 18395 -16090 18427 -16056
rect 18427 -16090 18429 -16056
rect 18467 -16090 18495 -16056
rect 18495 -16090 18501 -16056
rect 18539 -16090 18563 -16056
rect 18563 -16090 18573 -16056
rect 19197 -16090 19207 -16056
rect 19207 -16090 19231 -16056
rect 19269 -16090 19275 -16056
rect 19275 -16090 19303 -16056
rect 19341 -16090 19343 -16056
rect 19343 -16090 19375 -16056
rect 19413 -16090 19445 -16056
rect 19445 -16090 19447 -16056
rect 19485 -16090 19513 -16056
rect 19513 -16090 19519 -16056
rect 19557 -16090 19581 -16056
rect 19581 -16090 19591 -16056
rect 20215 -16090 20225 -16056
rect 20225 -16090 20249 -16056
rect 20287 -16090 20293 -16056
rect 20293 -16090 20321 -16056
rect 20359 -16090 20361 -16056
rect 20361 -16090 20393 -16056
rect 20431 -16090 20463 -16056
rect 20463 -16090 20465 -16056
rect 20503 -16090 20531 -16056
rect 20531 -16090 20537 -16056
rect 20575 -16090 20599 -16056
rect 20599 -16090 20609 -16056
rect 21233 -16090 21243 -16056
rect 21243 -16090 21267 -16056
rect 21305 -16090 21311 -16056
rect 21311 -16090 21339 -16056
rect 21377 -16090 21379 -16056
rect 21379 -16090 21411 -16056
rect 21449 -16090 21481 -16056
rect 21481 -16090 21483 -16056
rect 21521 -16090 21549 -16056
rect 21549 -16090 21555 -16056
rect 21593 -16090 21617 -16056
rect 21617 -16090 21627 -16056
rect 22251 -16090 22261 -16056
rect 22261 -16090 22285 -16056
rect 22323 -16090 22329 -16056
rect 22329 -16090 22357 -16056
rect 22395 -16090 22397 -16056
rect 22397 -16090 22429 -16056
rect 22467 -16090 22499 -16056
rect 22499 -16090 22501 -16056
rect 22539 -16090 22567 -16056
rect 22567 -16090 22573 -16056
rect 22611 -16090 22635 -16056
rect 22635 -16090 22645 -16056
rect 24855 -16055 24889 -16051
rect 24855 -16085 24889 -16055
rect -22 -16135 12 -16103
rect -22 -16137 12 -16135
rect -22 -16203 12 -16175
rect -22 -16209 12 -16203
rect -22 -16271 12 -16247
rect -22 -16281 12 -16271
rect -22 -16339 12 -16319
rect -22 -16353 12 -16339
rect 24855 -16157 24889 -16123
rect 24855 -16225 24889 -16195
rect 24855 -16229 24889 -16225
rect 24855 -16293 24889 -16267
rect 24855 -16301 24889 -16293
rect 24855 -16361 24889 -16339
rect 24855 -16373 24889 -16361
rect -12289 -16429 -12255 -16411
rect -12289 -16445 -12255 -16429
rect -8855 -16456 -8845 -16422
rect -8845 -16456 -8821 -16422
rect -8783 -16456 -8777 -16422
rect -8777 -16456 -8749 -16422
rect -8711 -16456 -8709 -16422
rect -8709 -16456 -8677 -16422
rect -8639 -16456 -8607 -16422
rect -8607 -16456 -8605 -16422
rect -8567 -16456 -8539 -16422
rect -8539 -16456 -8533 -16422
rect -8495 -16456 -8471 -16422
rect -8471 -16456 -8461 -16422
rect -7837 -16456 -7827 -16422
rect -7827 -16456 -7803 -16422
rect -7765 -16456 -7759 -16422
rect -7759 -16456 -7731 -16422
rect -7693 -16456 -7691 -16422
rect -7691 -16456 -7659 -16422
rect -7621 -16456 -7589 -16422
rect -7589 -16456 -7587 -16422
rect -7549 -16456 -7521 -16422
rect -7521 -16456 -7515 -16422
rect -7477 -16456 -7453 -16422
rect -7453 -16456 -7443 -16422
rect -6819 -16456 -6809 -16422
rect -6809 -16456 -6785 -16422
rect -6747 -16456 -6741 -16422
rect -6741 -16456 -6713 -16422
rect -6675 -16456 -6673 -16422
rect -6673 -16456 -6641 -16422
rect -6603 -16456 -6571 -16422
rect -6571 -16456 -6569 -16422
rect -6531 -16456 -6503 -16422
rect -6503 -16456 -6497 -16422
rect -6459 -16456 -6435 -16422
rect -6435 -16456 -6425 -16422
rect -5801 -16456 -5791 -16422
rect -5791 -16456 -5767 -16422
rect -5729 -16456 -5723 -16422
rect -5723 -16456 -5695 -16422
rect -5657 -16456 -5655 -16422
rect -5655 -16456 -5623 -16422
rect -5585 -16456 -5553 -16422
rect -5553 -16456 -5551 -16422
rect -5513 -16456 -5485 -16422
rect -5485 -16456 -5479 -16422
rect -5441 -16456 -5417 -16422
rect -5417 -16456 -5407 -16422
rect -4783 -16456 -4773 -16422
rect -4773 -16456 -4749 -16422
rect -4711 -16456 -4705 -16422
rect -4705 -16456 -4677 -16422
rect -4639 -16456 -4637 -16422
rect -4637 -16456 -4605 -16422
rect -4567 -16456 -4535 -16422
rect -4535 -16456 -4533 -16422
rect -4495 -16456 -4467 -16422
rect -4467 -16456 -4461 -16422
rect -4423 -16456 -4399 -16422
rect -4399 -16456 -4389 -16422
rect -3765 -16456 -3755 -16422
rect -3755 -16456 -3731 -16422
rect -3693 -16456 -3687 -16422
rect -3687 -16456 -3659 -16422
rect -3621 -16456 -3619 -16422
rect -3619 -16456 -3587 -16422
rect -3549 -16456 -3517 -16422
rect -3517 -16456 -3515 -16422
rect -3477 -16456 -3449 -16422
rect -3449 -16456 -3443 -16422
rect -3405 -16456 -3381 -16422
rect -3381 -16456 -3371 -16422
rect -2747 -16456 -2737 -16422
rect -2737 -16456 -2713 -16422
rect -2675 -16456 -2669 -16422
rect -2669 -16456 -2641 -16422
rect -2603 -16456 -2601 -16422
rect -2601 -16456 -2569 -16422
rect -2531 -16456 -2499 -16422
rect -2499 -16456 -2497 -16422
rect -2459 -16456 -2431 -16422
rect -2431 -16456 -2425 -16422
rect -2387 -16456 -2363 -16422
rect -2363 -16456 -2353 -16422
rect -1729 -16456 -1719 -16422
rect -1719 -16456 -1695 -16422
rect -1657 -16456 -1651 -16422
rect -1651 -16456 -1623 -16422
rect -1585 -16456 -1583 -16422
rect -1583 -16456 -1551 -16422
rect -1513 -16456 -1481 -16422
rect -1481 -16456 -1479 -16422
rect -1441 -16456 -1413 -16422
rect -1413 -16456 -1407 -16422
rect -1369 -16456 -1345 -16422
rect -1345 -16456 -1335 -16422
rect -711 -16456 -701 -16422
rect -701 -16456 -677 -16422
rect -639 -16456 -633 -16422
rect -633 -16456 -605 -16422
rect -567 -16456 -565 -16422
rect -565 -16456 -533 -16422
rect -495 -16456 -463 -16422
rect -463 -16456 -461 -16422
rect -423 -16456 -395 -16422
rect -395 -16456 -389 -16422
rect -351 -16456 -327 -16422
rect -327 -16456 -317 -16422
rect 24855 -16429 24889 -16411
rect 24855 -16445 24889 -16429
rect -12289 -16497 -12255 -16483
rect -12289 -16517 -12255 -16497
rect 24855 -16497 24889 -16483
rect 24855 -16517 24889 -16497
rect -12289 -16565 -12255 -16555
rect -12289 -16589 -12255 -16565
rect -8855 -16564 -8845 -16530
rect -8845 -16564 -8821 -16530
rect -8783 -16564 -8777 -16530
rect -8777 -16564 -8749 -16530
rect -8711 -16564 -8709 -16530
rect -8709 -16564 -8677 -16530
rect -8639 -16564 -8607 -16530
rect -8607 -16564 -8605 -16530
rect -8567 -16564 -8539 -16530
rect -8539 -16564 -8533 -16530
rect -8495 -16564 -8471 -16530
rect -8471 -16564 -8461 -16530
rect -7837 -16564 -7827 -16530
rect -7827 -16564 -7803 -16530
rect -7765 -16564 -7759 -16530
rect -7759 -16564 -7731 -16530
rect -7693 -16564 -7691 -16530
rect -7691 -16564 -7659 -16530
rect -7621 -16564 -7589 -16530
rect -7589 -16564 -7587 -16530
rect -7549 -16564 -7521 -16530
rect -7521 -16564 -7515 -16530
rect -7477 -16564 -7453 -16530
rect -7453 -16564 -7443 -16530
rect -6819 -16564 -6809 -16530
rect -6809 -16564 -6785 -16530
rect -6747 -16564 -6741 -16530
rect -6741 -16564 -6713 -16530
rect -6675 -16564 -6673 -16530
rect -6673 -16564 -6641 -16530
rect -6603 -16564 -6571 -16530
rect -6571 -16564 -6569 -16530
rect -6531 -16564 -6503 -16530
rect -6503 -16564 -6497 -16530
rect -6459 -16564 -6435 -16530
rect -6435 -16564 -6425 -16530
rect -5801 -16564 -5791 -16530
rect -5791 -16564 -5767 -16530
rect -5729 -16564 -5723 -16530
rect -5723 -16564 -5695 -16530
rect -5657 -16564 -5655 -16530
rect -5655 -16564 -5623 -16530
rect -5585 -16564 -5553 -16530
rect -5553 -16564 -5551 -16530
rect -5513 -16564 -5485 -16530
rect -5485 -16564 -5479 -16530
rect -5441 -16564 -5417 -16530
rect -5417 -16564 -5407 -16530
rect -4783 -16564 -4773 -16530
rect -4773 -16564 -4749 -16530
rect -4711 -16564 -4705 -16530
rect -4705 -16564 -4677 -16530
rect -4639 -16564 -4637 -16530
rect -4637 -16564 -4605 -16530
rect -4567 -16564 -4535 -16530
rect -4535 -16564 -4533 -16530
rect -4495 -16564 -4467 -16530
rect -4467 -16564 -4461 -16530
rect -4423 -16564 -4399 -16530
rect -4399 -16564 -4389 -16530
rect -3765 -16564 -3755 -16530
rect -3755 -16564 -3731 -16530
rect -3693 -16564 -3687 -16530
rect -3687 -16564 -3659 -16530
rect -3621 -16564 -3619 -16530
rect -3619 -16564 -3587 -16530
rect -3549 -16564 -3517 -16530
rect -3517 -16564 -3515 -16530
rect -3477 -16564 -3449 -16530
rect -3449 -16564 -3443 -16530
rect -3405 -16564 -3381 -16530
rect -3381 -16564 -3371 -16530
rect -2747 -16564 -2737 -16530
rect -2737 -16564 -2713 -16530
rect -2675 -16564 -2669 -16530
rect -2669 -16564 -2641 -16530
rect -2603 -16564 -2601 -16530
rect -2601 -16564 -2569 -16530
rect -2531 -16564 -2499 -16530
rect -2499 -16564 -2497 -16530
rect -2459 -16564 -2431 -16530
rect -2431 -16564 -2425 -16530
rect -2387 -16564 -2363 -16530
rect -2363 -16564 -2353 -16530
rect -1729 -16564 -1719 -16530
rect -1719 -16564 -1695 -16530
rect -1657 -16564 -1651 -16530
rect -1651 -16564 -1623 -16530
rect -1585 -16564 -1583 -16530
rect -1583 -16564 -1551 -16530
rect -1513 -16564 -1481 -16530
rect -1481 -16564 -1479 -16530
rect -1441 -16564 -1413 -16530
rect -1413 -16564 -1407 -16530
rect -1369 -16564 -1345 -16530
rect -1345 -16564 -1335 -16530
rect -711 -16564 -701 -16530
rect -701 -16564 -677 -16530
rect -639 -16564 -633 -16530
rect -633 -16564 -605 -16530
rect -567 -16564 -565 -16530
rect -565 -16564 -533 -16530
rect -495 -16564 -463 -16530
rect -463 -16564 -461 -16530
rect -423 -16564 -395 -16530
rect -395 -16564 -389 -16530
rect -351 -16564 -327 -16530
rect -327 -16564 -317 -16530
rect -12289 -16633 -12255 -16627
rect -12289 -16661 -12255 -16633
rect -12289 -16701 -12255 -16699
rect -12289 -16733 -12255 -16701
rect -12289 -16803 -12255 -16771
rect -12289 -16805 -12255 -16803
rect -12289 -16871 -12255 -16843
rect -12289 -16877 -12255 -16871
rect -12289 -16939 -12255 -16915
rect -12289 -16949 -12255 -16939
rect -12289 -17007 -12255 -16987
rect -12289 -17021 -12255 -17007
rect -12289 -17075 -12255 -17059
rect -12289 -17093 -12255 -17075
rect -12289 -17143 -12255 -17131
rect -12289 -17165 -12255 -17143
rect -12289 -17211 -12255 -17203
rect -12289 -17237 -12255 -17211
rect -9184 -16647 -9150 -16633
rect -9184 -16667 -9150 -16647
rect -9184 -16715 -9150 -16705
rect -9184 -16739 -9150 -16715
rect -9184 -16783 -9150 -16777
rect -9184 -16811 -9150 -16783
rect -9184 -16851 -9150 -16849
rect -9184 -16883 -9150 -16851
rect -9184 -16953 -9150 -16921
rect -9184 -16955 -9150 -16953
rect -9184 -17021 -9150 -16993
rect -9184 -17027 -9150 -17021
rect -9184 -17089 -9150 -17065
rect -9184 -17099 -9150 -17089
rect -9184 -17157 -9150 -17137
rect -9184 -17171 -9150 -17157
rect -8166 -16647 -8132 -16633
rect -8166 -16667 -8132 -16647
rect -8166 -16715 -8132 -16705
rect -8166 -16739 -8132 -16715
rect -8166 -16783 -8132 -16777
rect -8166 -16811 -8132 -16783
rect -8166 -16851 -8132 -16849
rect -8166 -16883 -8132 -16851
rect -8166 -16953 -8132 -16921
rect -8166 -16955 -8132 -16953
rect -8166 -17021 -8132 -16993
rect -8166 -17027 -8132 -17021
rect -8166 -17089 -8132 -17065
rect -8166 -17099 -8132 -17089
rect -8166 -17157 -8132 -17137
rect -8166 -17171 -8132 -17157
rect -7148 -16647 -7114 -16633
rect -7148 -16667 -7114 -16647
rect -7148 -16715 -7114 -16705
rect -7148 -16739 -7114 -16715
rect -7148 -16783 -7114 -16777
rect -7148 -16811 -7114 -16783
rect -7148 -16851 -7114 -16849
rect -7148 -16883 -7114 -16851
rect -7148 -16953 -7114 -16921
rect -7148 -16955 -7114 -16953
rect -7148 -17021 -7114 -16993
rect -7148 -17027 -7114 -17021
rect -7148 -17089 -7114 -17065
rect -7148 -17099 -7114 -17089
rect -7148 -17157 -7114 -17137
rect -7148 -17171 -7114 -17157
rect -6130 -16647 -6096 -16633
rect -6130 -16667 -6096 -16647
rect -6130 -16715 -6096 -16705
rect -6130 -16739 -6096 -16715
rect -6130 -16783 -6096 -16777
rect -6130 -16811 -6096 -16783
rect -6130 -16851 -6096 -16849
rect -6130 -16883 -6096 -16851
rect -6130 -16953 -6096 -16921
rect -6130 -16955 -6096 -16953
rect -6130 -17021 -6096 -16993
rect -6130 -17027 -6096 -17021
rect -6130 -17089 -6096 -17065
rect -6130 -17099 -6096 -17089
rect -6130 -17157 -6096 -17137
rect -6130 -17171 -6096 -17157
rect -5112 -16647 -5078 -16633
rect -5112 -16667 -5078 -16647
rect -5112 -16715 -5078 -16705
rect -5112 -16739 -5078 -16715
rect -5112 -16783 -5078 -16777
rect -5112 -16811 -5078 -16783
rect -5112 -16851 -5078 -16849
rect -5112 -16883 -5078 -16851
rect -5112 -16953 -5078 -16921
rect -5112 -16955 -5078 -16953
rect -5112 -17021 -5078 -16993
rect -5112 -17027 -5078 -17021
rect -5112 -17089 -5078 -17065
rect -5112 -17099 -5078 -17089
rect -5112 -17157 -5078 -17137
rect -5112 -17171 -5078 -17157
rect -4094 -16647 -4060 -16633
rect -4094 -16667 -4060 -16647
rect -4094 -16715 -4060 -16705
rect -4094 -16739 -4060 -16715
rect -4094 -16783 -4060 -16777
rect -4094 -16811 -4060 -16783
rect -4094 -16851 -4060 -16849
rect -4094 -16883 -4060 -16851
rect -4094 -16953 -4060 -16921
rect -4094 -16955 -4060 -16953
rect -4094 -17021 -4060 -16993
rect -4094 -17027 -4060 -17021
rect -4094 -17089 -4060 -17065
rect -4094 -17099 -4060 -17089
rect -4094 -17157 -4060 -17137
rect -4094 -17171 -4060 -17157
rect -3076 -16647 -3042 -16633
rect -3076 -16667 -3042 -16647
rect -3076 -16715 -3042 -16705
rect -3076 -16739 -3042 -16715
rect -3076 -16783 -3042 -16777
rect -3076 -16811 -3042 -16783
rect -3076 -16851 -3042 -16849
rect -3076 -16883 -3042 -16851
rect -3076 -16953 -3042 -16921
rect -3076 -16955 -3042 -16953
rect -3076 -17021 -3042 -16993
rect -3076 -17027 -3042 -17021
rect -3076 -17089 -3042 -17065
rect -3076 -17099 -3042 -17089
rect -3076 -17157 -3042 -17137
rect -3076 -17171 -3042 -17157
rect -2058 -16647 -2024 -16633
rect -2058 -16667 -2024 -16647
rect -2058 -16715 -2024 -16705
rect -2058 -16739 -2024 -16715
rect -2058 -16783 -2024 -16777
rect -2058 -16811 -2024 -16783
rect -2058 -16851 -2024 -16849
rect -2058 -16883 -2024 -16851
rect -2058 -16953 -2024 -16921
rect -2058 -16955 -2024 -16953
rect -2058 -17021 -2024 -16993
rect -2058 -17027 -2024 -17021
rect -2058 -17089 -2024 -17065
rect -2058 -17099 -2024 -17089
rect -2058 -17157 -2024 -17137
rect -2058 -17171 -2024 -17157
rect -1040 -16647 -1006 -16633
rect -1040 -16667 -1006 -16647
rect -1040 -16715 -1006 -16705
rect -1040 -16739 -1006 -16715
rect -1040 -16783 -1006 -16777
rect -1040 -16811 -1006 -16783
rect -1040 -16851 -1006 -16849
rect -1040 -16883 -1006 -16851
rect -1040 -16953 -1006 -16921
rect -1040 -16955 -1006 -16953
rect -1040 -17021 -1006 -16993
rect -1040 -17027 -1006 -17021
rect -1040 -17089 -1006 -17065
rect -1040 -17099 -1006 -17089
rect -1040 -17157 -1006 -17137
rect -1040 -17171 -1006 -17157
rect 2909 -16614 2919 -16580
rect 2919 -16614 2943 -16580
rect 2981 -16614 2987 -16580
rect 2987 -16614 3015 -16580
rect 3053 -16614 3055 -16580
rect 3055 -16614 3087 -16580
rect 3125 -16614 3157 -16580
rect 3157 -16614 3159 -16580
rect 3197 -16614 3225 -16580
rect 3225 -16614 3231 -16580
rect 3269 -16614 3293 -16580
rect 3293 -16614 3303 -16580
rect 3927 -16614 3937 -16580
rect 3937 -16614 3961 -16580
rect 3999 -16614 4005 -16580
rect 4005 -16614 4033 -16580
rect 4071 -16614 4073 -16580
rect 4073 -16614 4105 -16580
rect 4143 -16614 4175 -16580
rect 4175 -16614 4177 -16580
rect 4215 -16614 4243 -16580
rect 4243 -16614 4249 -16580
rect 4287 -16614 4311 -16580
rect 4311 -16614 4321 -16580
rect 4945 -16614 4955 -16580
rect 4955 -16614 4979 -16580
rect 5017 -16614 5023 -16580
rect 5023 -16614 5051 -16580
rect 5089 -16614 5091 -16580
rect 5091 -16614 5123 -16580
rect 5161 -16614 5193 -16580
rect 5193 -16614 5195 -16580
rect 5233 -16614 5261 -16580
rect 5261 -16614 5267 -16580
rect 5305 -16614 5329 -16580
rect 5329 -16614 5339 -16580
rect 5963 -16614 5973 -16580
rect 5973 -16614 5997 -16580
rect 6035 -16614 6041 -16580
rect 6041 -16614 6069 -16580
rect 6107 -16614 6109 -16580
rect 6109 -16614 6141 -16580
rect 6179 -16614 6211 -16580
rect 6211 -16614 6213 -16580
rect 6251 -16614 6279 -16580
rect 6279 -16614 6285 -16580
rect 6323 -16614 6347 -16580
rect 6347 -16614 6357 -16580
rect 6981 -16614 6991 -16580
rect 6991 -16614 7015 -16580
rect 7053 -16614 7059 -16580
rect 7059 -16614 7087 -16580
rect 7125 -16614 7127 -16580
rect 7127 -16614 7159 -16580
rect 7197 -16614 7229 -16580
rect 7229 -16614 7231 -16580
rect 7269 -16614 7297 -16580
rect 7297 -16614 7303 -16580
rect 7341 -16614 7365 -16580
rect 7365 -16614 7375 -16580
rect 7999 -16614 8009 -16580
rect 8009 -16614 8033 -16580
rect 8071 -16614 8077 -16580
rect 8077 -16614 8105 -16580
rect 8143 -16614 8145 -16580
rect 8145 -16614 8177 -16580
rect 8215 -16614 8247 -16580
rect 8247 -16614 8249 -16580
rect 8287 -16614 8315 -16580
rect 8315 -16614 8321 -16580
rect 8359 -16614 8383 -16580
rect 8383 -16614 8393 -16580
rect 9017 -16614 9027 -16580
rect 9027 -16614 9051 -16580
rect 9089 -16614 9095 -16580
rect 9095 -16614 9123 -16580
rect 9161 -16614 9163 -16580
rect 9163 -16614 9195 -16580
rect 9233 -16614 9265 -16580
rect 9265 -16614 9267 -16580
rect 9305 -16614 9333 -16580
rect 9333 -16614 9339 -16580
rect 9377 -16614 9401 -16580
rect 9401 -16614 9411 -16580
rect 10035 -16614 10045 -16580
rect 10045 -16614 10069 -16580
rect 10107 -16614 10113 -16580
rect 10113 -16614 10141 -16580
rect 10179 -16614 10181 -16580
rect 10181 -16614 10213 -16580
rect 10251 -16614 10283 -16580
rect 10283 -16614 10285 -16580
rect 10323 -16614 10351 -16580
rect 10351 -16614 10357 -16580
rect 10395 -16614 10419 -16580
rect 10419 -16614 10429 -16580
rect 11053 -16614 11063 -16580
rect 11063 -16614 11087 -16580
rect 11125 -16614 11131 -16580
rect 11131 -16614 11159 -16580
rect 11197 -16614 11199 -16580
rect 11199 -16614 11231 -16580
rect 11269 -16614 11301 -16580
rect 11301 -16614 11303 -16580
rect 11341 -16614 11369 -16580
rect 11369 -16614 11375 -16580
rect 11413 -16614 11437 -16580
rect 11437 -16614 11447 -16580
rect 12071 -16614 12081 -16580
rect 12081 -16614 12105 -16580
rect 12143 -16614 12149 -16580
rect 12149 -16614 12177 -16580
rect 12215 -16614 12217 -16580
rect 12217 -16614 12249 -16580
rect 12287 -16614 12319 -16580
rect 12319 -16614 12321 -16580
rect 12359 -16614 12387 -16580
rect 12387 -16614 12393 -16580
rect 12431 -16614 12455 -16580
rect 12455 -16614 12465 -16580
rect 13089 -16614 13099 -16580
rect 13099 -16614 13123 -16580
rect 13161 -16614 13167 -16580
rect 13167 -16614 13195 -16580
rect 13233 -16614 13235 -16580
rect 13235 -16614 13267 -16580
rect 13305 -16614 13337 -16580
rect 13337 -16614 13339 -16580
rect 13377 -16614 13405 -16580
rect 13405 -16614 13411 -16580
rect 13449 -16614 13473 -16580
rect 13473 -16614 13483 -16580
rect 14107 -16614 14117 -16580
rect 14117 -16614 14141 -16580
rect 14179 -16614 14185 -16580
rect 14185 -16614 14213 -16580
rect 14251 -16614 14253 -16580
rect 14253 -16614 14285 -16580
rect 14323 -16614 14355 -16580
rect 14355 -16614 14357 -16580
rect 14395 -16614 14423 -16580
rect 14423 -16614 14429 -16580
rect 14467 -16614 14491 -16580
rect 14491 -16614 14501 -16580
rect 15125 -16614 15135 -16580
rect 15135 -16614 15159 -16580
rect 15197 -16614 15203 -16580
rect 15203 -16614 15231 -16580
rect 15269 -16614 15271 -16580
rect 15271 -16614 15303 -16580
rect 15341 -16614 15373 -16580
rect 15373 -16614 15375 -16580
rect 15413 -16614 15441 -16580
rect 15441 -16614 15447 -16580
rect 15485 -16614 15509 -16580
rect 15509 -16614 15519 -16580
rect 16143 -16614 16153 -16580
rect 16153 -16614 16177 -16580
rect 16215 -16614 16221 -16580
rect 16221 -16614 16249 -16580
rect 16287 -16614 16289 -16580
rect 16289 -16614 16321 -16580
rect 16359 -16614 16391 -16580
rect 16391 -16614 16393 -16580
rect 16431 -16614 16459 -16580
rect 16459 -16614 16465 -16580
rect 16503 -16614 16527 -16580
rect 16527 -16614 16537 -16580
rect 17161 -16614 17171 -16580
rect 17171 -16614 17195 -16580
rect 17233 -16614 17239 -16580
rect 17239 -16614 17267 -16580
rect 17305 -16614 17307 -16580
rect 17307 -16614 17339 -16580
rect 17377 -16614 17409 -16580
rect 17409 -16614 17411 -16580
rect 17449 -16614 17477 -16580
rect 17477 -16614 17483 -16580
rect 17521 -16614 17545 -16580
rect 17545 -16614 17555 -16580
rect 18179 -16614 18189 -16580
rect 18189 -16614 18213 -16580
rect 18251 -16614 18257 -16580
rect 18257 -16614 18285 -16580
rect 18323 -16614 18325 -16580
rect 18325 -16614 18357 -16580
rect 18395 -16614 18427 -16580
rect 18427 -16614 18429 -16580
rect 18467 -16614 18495 -16580
rect 18495 -16614 18501 -16580
rect 18539 -16614 18563 -16580
rect 18563 -16614 18573 -16580
rect 19197 -16614 19207 -16580
rect 19207 -16614 19231 -16580
rect 19269 -16614 19275 -16580
rect 19275 -16614 19303 -16580
rect 19341 -16614 19343 -16580
rect 19343 -16614 19375 -16580
rect 19413 -16614 19445 -16580
rect 19445 -16614 19447 -16580
rect 19485 -16614 19513 -16580
rect 19513 -16614 19519 -16580
rect 19557 -16614 19581 -16580
rect 19581 -16614 19591 -16580
rect 20215 -16614 20225 -16580
rect 20225 -16614 20249 -16580
rect 20287 -16614 20293 -16580
rect 20293 -16614 20321 -16580
rect 20359 -16614 20361 -16580
rect 20361 -16614 20393 -16580
rect 20431 -16614 20463 -16580
rect 20463 -16614 20465 -16580
rect 20503 -16614 20531 -16580
rect 20531 -16614 20537 -16580
rect 20575 -16614 20599 -16580
rect 20599 -16614 20609 -16580
rect 21233 -16614 21243 -16580
rect 21243 -16614 21267 -16580
rect 21305 -16614 21311 -16580
rect 21311 -16614 21339 -16580
rect 21377 -16614 21379 -16580
rect 21379 -16614 21411 -16580
rect 21449 -16614 21481 -16580
rect 21481 -16614 21483 -16580
rect 21521 -16614 21549 -16580
rect 21549 -16614 21555 -16580
rect 21593 -16614 21617 -16580
rect 21617 -16614 21627 -16580
rect 22251 -16614 22261 -16580
rect 22261 -16614 22285 -16580
rect 22323 -16614 22329 -16580
rect 22329 -16614 22357 -16580
rect 22395 -16614 22397 -16580
rect 22397 -16614 22429 -16580
rect 22467 -16614 22499 -16580
rect 22499 -16614 22501 -16580
rect 22539 -16614 22567 -16580
rect 22567 -16614 22573 -16580
rect 22611 -16614 22635 -16580
rect 22635 -16614 22645 -16580
rect 24855 -16565 24889 -16555
rect 24855 -16589 24889 -16565
rect -22 -16647 12 -16633
rect -22 -16667 12 -16647
rect -22 -16715 12 -16705
rect -22 -16739 12 -16715
rect -22 -16783 12 -16777
rect -22 -16811 12 -16783
rect -22 -16851 12 -16849
rect -22 -16883 12 -16851
rect -22 -16953 12 -16921
rect -22 -16955 12 -16953
rect -22 -17021 12 -16993
rect -22 -17027 12 -17021
rect -22 -17089 12 -17065
rect -22 -17099 12 -17089
rect -22 -17157 12 -17137
rect -22 -17171 12 -17157
rect 2580 -16697 2614 -16683
rect 2580 -16717 2614 -16697
rect 2580 -16765 2614 -16755
rect 2580 -16789 2614 -16765
rect 2580 -16833 2614 -16827
rect 2580 -16861 2614 -16833
rect 2580 -16901 2614 -16899
rect 2580 -16933 2614 -16901
rect 2580 -17003 2614 -16971
rect 2580 -17005 2614 -17003
rect 2580 -17071 2614 -17043
rect 2580 -17077 2614 -17071
rect 2580 -17139 2614 -17115
rect 2580 -17149 2614 -17139
rect 2580 -17207 2614 -17187
rect 2580 -17221 2614 -17207
rect -8855 -17274 -8845 -17240
rect -8845 -17274 -8821 -17240
rect -8783 -17274 -8777 -17240
rect -8777 -17274 -8749 -17240
rect -8711 -17274 -8709 -17240
rect -8709 -17274 -8677 -17240
rect -8639 -17274 -8607 -17240
rect -8607 -17274 -8605 -17240
rect -8567 -17274 -8539 -17240
rect -8539 -17274 -8533 -17240
rect -8495 -17274 -8471 -17240
rect -8471 -17274 -8461 -17240
rect -7837 -17274 -7827 -17240
rect -7827 -17274 -7803 -17240
rect -7765 -17274 -7759 -17240
rect -7759 -17274 -7731 -17240
rect -7693 -17274 -7691 -17240
rect -7691 -17274 -7659 -17240
rect -7621 -17274 -7589 -17240
rect -7589 -17274 -7587 -17240
rect -7549 -17274 -7521 -17240
rect -7521 -17274 -7515 -17240
rect -7477 -17274 -7453 -17240
rect -7453 -17274 -7443 -17240
rect -6819 -17274 -6809 -17240
rect -6809 -17274 -6785 -17240
rect -6747 -17274 -6741 -17240
rect -6741 -17274 -6713 -17240
rect -6675 -17274 -6673 -17240
rect -6673 -17274 -6641 -17240
rect -6603 -17274 -6571 -17240
rect -6571 -17274 -6569 -17240
rect -6531 -17274 -6503 -17240
rect -6503 -17274 -6497 -17240
rect -6459 -17274 -6435 -17240
rect -6435 -17274 -6425 -17240
rect -5801 -17274 -5791 -17240
rect -5791 -17274 -5767 -17240
rect -5729 -17274 -5723 -17240
rect -5723 -17274 -5695 -17240
rect -5657 -17274 -5655 -17240
rect -5655 -17274 -5623 -17240
rect -5585 -17274 -5553 -17240
rect -5553 -17274 -5551 -17240
rect -5513 -17274 -5485 -17240
rect -5485 -17274 -5479 -17240
rect -5441 -17274 -5417 -17240
rect -5417 -17274 -5407 -17240
rect -4783 -17274 -4773 -17240
rect -4773 -17274 -4749 -17240
rect -4711 -17274 -4705 -17240
rect -4705 -17274 -4677 -17240
rect -4639 -17274 -4637 -17240
rect -4637 -17274 -4605 -17240
rect -4567 -17274 -4535 -17240
rect -4535 -17274 -4533 -17240
rect -4495 -17274 -4467 -17240
rect -4467 -17274 -4461 -17240
rect -4423 -17274 -4399 -17240
rect -4399 -17274 -4389 -17240
rect -3765 -17274 -3755 -17240
rect -3755 -17274 -3731 -17240
rect -3693 -17274 -3687 -17240
rect -3687 -17274 -3659 -17240
rect -3621 -17274 -3619 -17240
rect -3619 -17274 -3587 -17240
rect -3549 -17274 -3517 -17240
rect -3517 -17274 -3515 -17240
rect -3477 -17274 -3449 -17240
rect -3449 -17274 -3443 -17240
rect -3405 -17274 -3381 -17240
rect -3381 -17274 -3371 -17240
rect -2747 -17274 -2737 -17240
rect -2737 -17274 -2713 -17240
rect -2675 -17274 -2669 -17240
rect -2669 -17274 -2641 -17240
rect -2603 -17274 -2601 -17240
rect -2601 -17274 -2569 -17240
rect -2531 -17274 -2499 -17240
rect -2499 -17274 -2497 -17240
rect -2459 -17274 -2431 -17240
rect -2431 -17274 -2425 -17240
rect -2387 -17274 -2363 -17240
rect -2363 -17274 -2353 -17240
rect -1729 -17274 -1719 -17240
rect -1719 -17274 -1695 -17240
rect -1657 -17274 -1651 -17240
rect -1651 -17274 -1623 -17240
rect -1585 -17274 -1583 -17240
rect -1583 -17274 -1551 -17240
rect -1513 -17274 -1481 -17240
rect -1481 -17274 -1479 -17240
rect -1441 -17274 -1413 -17240
rect -1413 -17274 -1407 -17240
rect -1369 -17274 -1345 -17240
rect -1345 -17274 -1335 -17240
rect -711 -17274 -701 -17240
rect -701 -17274 -677 -17240
rect -639 -17274 -633 -17240
rect -633 -17274 -605 -17240
rect -567 -17274 -565 -17240
rect -565 -17274 -533 -17240
rect -495 -17274 -463 -17240
rect -463 -17274 -461 -17240
rect -423 -17274 -395 -17240
rect -395 -17274 -389 -17240
rect -351 -17274 -327 -17240
rect -327 -17274 -317 -17240
rect 3598 -16697 3632 -16683
rect 3598 -16717 3632 -16697
rect 3598 -16765 3632 -16755
rect 3598 -16789 3632 -16765
rect 3598 -16833 3632 -16827
rect 3598 -16861 3632 -16833
rect 3598 -16901 3632 -16899
rect 3598 -16933 3632 -16901
rect 3598 -17003 3632 -16971
rect 3598 -17005 3632 -17003
rect 3598 -17071 3632 -17043
rect 3598 -17077 3632 -17071
rect 3598 -17139 3632 -17115
rect 3598 -17149 3632 -17139
rect 3598 -17207 3632 -17187
rect 3598 -17221 3632 -17207
rect 4616 -16697 4650 -16683
rect 4616 -16717 4650 -16697
rect 4616 -16765 4650 -16755
rect 4616 -16789 4650 -16765
rect 4616 -16833 4650 -16827
rect 4616 -16861 4650 -16833
rect 4616 -16901 4650 -16899
rect 4616 -16933 4650 -16901
rect 4616 -17003 4650 -16971
rect 4616 -17005 4650 -17003
rect 4616 -17071 4650 -17043
rect 4616 -17077 4650 -17071
rect 4616 -17139 4650 -17115
rect 4616 -17149 4650 -17139
rect 4616 -17207 4650 -17187
rect 4616 -17221 4650 -17207
rect 5634 -16697 5668 -16683
rect 5634 -16717 5668 -16697
rect 5634 -16765 5668 -16755
rect 5634 -16789 5668 -16765
rect 5634 -16833 5668 -16827
rect 5634 -16861 5668 -16833
rect 5634 -16901 5668 -16899
rect 5634 -16933 5668 -16901
rect 5634 -17003 5668 -16971
rect 5634 -17005 5668 -17003
rect 5634 -17071 5668 -17043
rect 5634 -17077 5668 -17071
rect 5634 -17139 5668 -17115
rect 5634 -17149 5668 -17139
rect 5634 -17207 5668 -17187
rect 5634 -17221 5668 -17207
rect 6652 -16697 6686 -16683
rect 6652 -16717 6686 -16697
rect 6652 -16765 6686 -16755
rect 6652 -16789 6686 -16765
rect 6652 -16833 6686 -16827
rect 6652 -16861 6686 -16833
rect 6652 -16901 6686 -16899
rect 6652 -16933 6686 -16901
rect 6652 -17003 6686 -16971
rect 6652 -17005 6686 -17003
rect 6652 -17071 6686 -17043
rect 6652 -17077 6686 -17071
rect 6652 -17139 6686 -17115
rect 6652 -17149 6686 -17139
rect 6652 -17207 6686 -17187
rect 6652 -17221 6686 -17207
rect 7670 -16697 7704 -16683
rect 7670 -16717 7704 -16697
rect 7670 -16765 7704 -16755
rect 7670 -16789 7704 -16765
rect 7670 -16833 7704 -16827
rect 7670 -16861 7704 -16833
rect 7670 -16901 7704 -16899
rect 7670 -16933 7704 -16901
rect 7670 -17003 7704 -16971
rect 7670 -17005 7704 -17003
rect 7670 -17071 7704 -17043
rect 7670 -17077 7704 -17071
rect 7670 -17139 7704 -17115
rect 7670 -17149 7704 -17139
rect 7670 -17207 7704 -17187
rect 7670 -17221 7704 -17207
rect 8688 -16697 8722 -16683
rect 8688 -16717 8722 -16697
rect 8688 -16765 8722 -16755
rect 8688 -16789 8722 -16765
rect 8688 -16833 8722 -16827
rect 8688 -16861 8722 -16833
rect 8688 -16901 8722 -16899
rect 8688 -16933 8722 -16901
rect 8688 -17003 8722 -16971
rect 8688 -17005 8722 -17003
rect 8688 -17071 8722 -17043
rect 8688 -17077 8722 -17071
rect 8688 -17139 8722 -17115
rect 8688 -17149 8722 -17139
rect 8688 -17207 8722 -17187
rect 8688 -17221 8722 -17207
rect 9706 -16697 9740 -16683
rect 9706 -16717 9740 -16697
rect 9706 -16765 9740 -16755
rect 9706 -16789 9740 -16765
rect 9706 -16833 9740 -16827
rect 9706 -16861 9740 -16833
rect 9706 -16901 9740 -16899
rect 9706 -16933 9740 -16901
rect 9706 -17003 9740 -16971
rect 9706 -17005 9740 -17003
rect 9706 -17071 9740 -17043
rect 9706 -17077 9740 -17071
rect 9706 -17139 9740 -17115
rect 9706 -17149 9740 -17139
rect 9706 -17207 9740 -17187
rect 9706 -17221 9740 -17207
rect 10724 -16697 10758 -16683
rect 10724 -16717 10758 -16697
rect 10724 -16765 10758 -16755
rect 10724 -16789 10758 -16765
rect 10724 -16833 10758 -16827
rect 10724 -16861 10758 -16833
rect 10724 -16901 10758 -16899
rect 10724 -16933 10758 -16901
rect 10724 -17003 10758 -16971
rect 10724 -17005 10758 -17003
rect 10724 -17071 10758 -17043
rect 10724 -17077 10758 -17071
rect 10724 -17139 10758 -17115
rect 10724 -17149 10758 -17139
rect 10724 -17207 10758 -17187
rect 10724 -17221 10758 -17207
rect 11742 -16697 11776 -16683
rect 11742 -16717 11776 -16697
rect 11742 -16765 11776 -16755
rect 11742 -16789 11776 -16765
rect 11742 -16833 11776 -16827
rect 11742 -16861 11776 -16833
rect 11742 -16901 11776 -16899
rect 11742 -16933 11776 -16901
rect 11742 -17003 11776 -16971
rect 11742 -17005 11776 -17003
rect 11742 -17071 11776 -17043
rect 11742 -17077 11776 -17071
rect 11742 -17139 11776 -17115
rect 11742 -17149 11776 -17139
rect 11742 -17207 11776 -17187
rect 11742 -17221 11776 -17207
rect 12760 -16697 12794 -16683
rect 12760 -16717 12794 -16697
rect 12760 -16765 12794 -16755
rect 12760 -16789 12794 -16765
rect 12760 -16833 12794 -16827
rect 12760 -16861 12794 -16833
rect 12760 -16901 12794 -16899
rect 12760 -16933 12794 -16901
rect 12760 -17003 12794 -16971
rect 12760 -17005 12794 -17003
rect 12760 -17071 12794 -17043
rect 12760 -17077 12794 -17071
rect 12760 -17139 12794 -17115
rect 12760 -17149 12794 -17139
rect 12760 -17207 12794 -17187
rect 12760 -17221 12794 -17207
rect 13778 -16697 13812 -16683
rect 13778 -16717 13812 -16697
rect 13778 -16765 13812 -16755
rect 13778 -16789 13812 -16765
rect 13778 -16833 13812 -16827
rect 13778 -16861 13812 -16833
rect 13778 -16901 13812 -16899
rect 13778 -16933 13812 -16901
rect 13778 -17003 13812 -16971
rect 13778 -17005 13812 -17003
rect 13778 -17071 13812 -17043
rect 13778 -17077 13812 -17071
rect 13778 -17139 13812 -17115
rect 13778 -17149 13812 -17139
rect 13778 -17207 13812 -17187
rect 13778 -17221 13812 -17207
rect 14796 -16697 14830 -16683
rect 14796 -16717 14830 -16697
rect 14796 -16765 14830 -16755
rect 14796 -16789 14830 -16765
rect 14796 -16833 14830 -16827
rect 14796 -16861 14830 -16833
rect 14796 -16901 14830 -16899
rect 14796 -16933 14830 -16901
rect 14796 -17003 14830 -16971
rect 14796 -17005 14830 -17003
rect 14796 -17071 14830 -17043
rect 14796 -17077 14830 -17071
rect 14796 -17139 14830 -17115
rect 14796 -17149 14830 -17139
rect 14796 -17207 14830 -17187
rect 14796 -17221 14830 -17207
rect 15814 -16697 15848 -16683
rect 15814 -16717 15848 -16697
rect 15814 -16765 15848 -16755
rect 15814 -16789 15848 -16765
rect 15814 -16833 15848 -16827
rect 15814 -16861 15848 -16833
rect 15814 -16901 15848 -16899
rect 15814 -16933 15848 -16901
rect 15814 -17003 15848 -16971
rect 15814 -17005 15848 -17003
rect 15814 -17071 15848 -17043
rect 15814 -17077 15848 -17071
rect 15814 -17139 15848 -17115
rect 15814 -17149 15848 -17139
rect 15814 -17207 15848 -17187
rect 15814 -17221 15848 -17207
rect 16832 -16697 16866 -16683
rect 16832 -16717 16866 -16697
rect 16832 -16765 16866 -16755
rect 16832 -16789 16866 -16765
rect 16832 -16833 16866 -16827
rect 16832 -16861 16866 -16833
rect 16832 -16901 16866 -16899
rect 16832 -16933 16866 -16901
rect 16832 -17003 16866 -16971
rect 16832 -17005 16866 -17003
rect 16832 -17071 16866 -17043
rect 16832 -17077 16866 -17071
rect 16832 -17139 16866 -17115
rect 16832 -17149 16866 -17139
rect 16832 -17207 16866 -17187
rect 16832 -17221 16866 -17207
rect 17850 -16697 17884 -16683
rect 17850 -16717 17884 -16697
rect 17850 -16765 17884 -16755
rect 17850 -16789 17884 -16765
rect 17850 -16833 17884 -16827
rect 17850 -16861 17884 -16833
rect 17850 -16901 17884 -16899
rect 17850 -16933 17884 -16901
rect 17850 -17003 17884 -16971
rect 17850 -17005 17884 -17003
rect 17850 -17071 17884 -17043
rect 17850 -17077 17884 -17071
rect 17850 -17139 17884 -17115
rect 17850 -17149 17884 -17139
rect 17850 -17207 17884 -17187
rect 17850 -17221 17884 -17207
rect 18868 -16697 18902 -16683
rect 18868 -16717 18902 -16697
rect 18868 -16765 18902 -16755
rect 18868 -16789 18902 -16765
rect 18868 -16833 18902 -16827
rect 18868 -16861 18902 -16833
rect 18868 -16901 18902 -16899
rect 18868 -16933 18902 -16901
rect 18868 -17003 18902 -16971
rect 18868 -17005 18902 -17003
rect 18868 -17071 18902 -17043
rect 18868 -17077 18902 -17071
rect 18868 -17139 18902 -17115
rect 18868 -17149 18902 -17139
rect 18868 -17207 18902 -17187
rect 18868 -17221 18902 -17207
rect 19886 -16697 19920 -16683
rect 19886 -16717 19920 -16697
rect 19886 -16765 19920 -16755
rect 19886 -16789 19920 -16765
rect 19886 -16833 19920 -16827
rect 19886 -16861 19920 -16833
rect 19886 -16901 19920 -16899
rect 19886 -16933 19920 -16901
rect 19886 -17003 19920 -16971
rect 19886 -17005 19920 -17003
rect 19886 -17071 19920 -17043
rect 19886 -17077 19920 -17071
rect 19886 -17139 19920 -17115
rect 19886 -17149 19920 -17139
rect 19886 -17207 19920 -17187
rect 19886 -17221 19920 -17207
rect 20904 -16697 20938 -16683
rect 20904 -16717 20938 -16697
rect 20904 -16765 20938 -16755
rect 20904 -16789 20938 -16765
rect 20904 -16833 20938 -16827
rect 20904 -16861 20938 -16833
rect 20904 -16901 20938 -16899
rect 20904 -16933 20938 -16901
rect 20904 -17003 20938 -16971
rect 20904 -17005 20938 -17003
rect 20904 -17071 20938 -17043
rect 20904 -17077 20938 -17071
rect 20904 -17139 20938 -17115
rect 20904 -17149 20938 -17139
rect 20904 -17207 20938 -17187
rect 20904 -17221 20938 -17207
rect 21922 -16697 21956 -16683
rect 21922 -16717 21956 -16697
rect 21922 -16765 21956 -16755
rect 21922 -16789 21956 -16765
rect 21922 -16833 21956 -16827
rect 21922 -16861 21956 -16833
rect 21922 -16901 21956 -16899
rect 21922 -16933 21956 -16901
rect 21922 -17003 21956 -16971
rect 21922 -17005 21956 -17003
rect 21922 -17071 21956 -17043
rect 21922 -17077 21956 -17071
rect 21922 -17139 21956 -17115
rect 21922 -17149 21956 -17139
rect 21922 -17207 21956 -17187
rect 21922 -17221 21956 -17207
rect 22940 -16697 22974 -16683
rect 22940 -16717 22974 -16697
rect 22940 -16765 22974 -16755
rect 22940 -16789 22974 -16765
rect 22940 -16833 22974 -16827
rect 22940 -16861 22974 -16833
rect 22940 -16901 22974 -16899
rect 22940 -16933 22974 -16901
rect 22940 -17003 22974 -16971
rect 22940 -17005 22974 -17003
rect 22940 -17071 22974 -17043
rect 22940 -17077 22974 -17071
rect 22940 -17139 22974 -17115
rect 22940 -17149 22974 -17139
rect 22940 -17207 22974 -17187
rect 22940 -17221 22974 -17207
rect 24855 -16633 24889 -16627
rect 24855 -16661 24889 -16633
rect 24855 -16701 24889 -16699
rect 24855 -16733 24889 -16701
rect 24855 -16803 24889 -16771
rect 24855 -16805 24889 -16803
rect 24855 -16871 24889 -16843
rect 24855 -16877 24889 -16871
rect 24855 -16939 24889 -16915
rect 24855 -16949 24889 -16939
rect 24855 -17007 24889 -16987
rect 24855 -17021 24889 -17007
rect 24855 -17075 24889 -17059
rect 24855 -17093 24889 -17075
rect 24855 -17143 24889 -17131
rect 24855 -17165 24889 -17143
rect 24855 -17211 24889 -17203
rect 24855 -17237 24889 -17211
rect -12289 -17279 -12255 -17275
rect -12289 -17309 -12255 -17279
rect 2909 -17324 2919 -17290
rect 2919 -17324 2943 -17290
rect 2981 -17324 2987 -17290
rect 2987 -17324 3015 -17290
rect 3053 -17324 3055 -17290
rect 3055 -17324 3087 -17290
rect 3125 -17324 3157 -17290
rect 3157 -17324 3159 -17290
rect 3197 -17324 3225 -17290
rect 3225 -17324 3231 -17290
rect 3269 -17324 3293 -17290
rect 3293 -17324 3303 -17290
rect 3927 -17324 3937 -17290
rect 3937 -17324 3961 -17290
rect 3999 -17324 4005 -17290
rect 4005 -17324 4033 -17290
rect 4071 -17324 4073 -17290
rect 4073 -17324 4105 -17290
rect 4143 -17324 4175 -17290
rect 4175 -17324 4177 -17290
rect 4215 -17324 4243 -17290
rect 4243 -17324 4249 -17290
rect 4287 -17324 4311 -17290
rect 4311 -17324 4321 -17290
rect 4945 -17324 4955 -17290
rect 4955 -17324 4979 -17290
rect 5017 -17324 5023 -17290
rect 5023 -17324 5051 -17290
rect 5089 -17324 5091 -17290
rect 5091 -17324 5123 -17290
rect 5161 -17324 5193 -17290
rect 5193 -17324 5195 -17290
rect 5233 -17324 5261 -17290
rect 5261 -17324 5267 -17290
rect 5305 -17324 5329 -17290
rect 5329 -17324 5339 -17290
rect 5963 -17324 5973 -17290
rect 5973 -17324 5997 -17290
rect 6035 -17324 6041 -17290
rect 6041 -17324 6069 -17290
rect 6107 -17324 6109 -17290
rect 6109 -17324 6141 -17290
rect 6179 -17324 6211 -17290
rect 6211 -17324 6213 -17290
rect 6251 -17324 6279 -17290
rect 6279 -17324 6285 -17290
rect 6323 -17324 6347 -17290
rect 6347 -17324 6357 -17290
rect 6981 -17324 6991 -17290
rect 6991 -17324 7015 -17290
rect 7053 -17324 7059 -17290
rect 7059 -17324 7087 -17290
rect 7125 -17324 7127 -17290
rect 7127 -17324 7159 -17290
rect 7197 -17324 7229 -17290
rect 7229 -17324 7231 -17290
rect 7269 -17324 7297 -17290
rect 7297 -17324 7303 -17290
rect 7341 -17324 7365 -17290
rect 7365 -17324 7375 -17290
rect 7999 -17324 8009 -17290
rect 8009 -17324 8033 -17290
rect 8071 -17324 8077 -17290
rect 8077 -17324 8105 -17290
rect 8143 -17324 8145 -17290
rect 8145 -17324 8177 -17290
rect 8215 -17324 8247 -17290
rect 8247 -17324 8249 -17290
rect 8287 -17324 8315 -17290
rect 8315 -17324 8321 -17290
rect 8359 -17324 8383 -17290
rect 8383 -17324 8393 -17290
rect 9017 -17324 9027 -17290
rect 9027 -17324 9051 -17290
rect 9089 -17324 9095 -17290
rect 9095 -17324 9123 -17290
rect 9161 -17324 9163 -17290
rect 9163 -17324 9195 -17290
rect 9233 -17324 9265 -17290
rect 9265 -17324 9267 -17290
rect 9305 -17324 9333 -17290
rect 9333 -17324 9339 -17290
rect 9377 -17324 9401 -17290
rect 9401 -17324 9411 -17290
rect 10035 -17324 10045 -17290
rect 10045 -17324 10069 -17290
rect 10107 -17324 10113 -17290
rect 10113 -17324 10141 -17290
rect 10179 -17324 10181 -17290
rect 10181 -17324 10213 -17290
rect 10251 -17324 10283 -17290
rect 10283 -17324 10285 -17290
rect 10323 -17324 10351 -17290
rect 10351 -17324 10357 -17290
rect 10395 -17324 10419 -17290
rect 10419 -17324 10429 -17290
rect 11053 -17324 11063 -17290
rect 11063 -17324 11087 -17290
rect 11125 -17324 11131 -17290
rect 11131 -17324 11159 -17290
rect 11197 -17324 11199 -17290
rect 11199 -17324 11231 -17290
rect 11269 -17324 11301 -17290
rect 11301 -17324 11303 -17290
rect 11341 -17324 11369 -17290
rect 11369 -17324 11375 -17290
rect 11413 -17324 11437 -17290
rect 11437 -17324 11447 -17290
rect 12071 -17324 12081 -17290
rect 12081 -17324 12105 -17290
rect 12143 -17324 12149 -17290
rect 12149 -17324 12177 -17290
rect 12215 -17324 12217 -17290
rect 12217 -17324 12249 -17290
rect 12287 -17324 12319 -17290
rect 12319 -17324 12321 -17290
rect 12359 -17324 12387 -17290
rect 12387 -17324 12393 -17290
rect 12431 -17324 12455 -17290
rect 12455 -17324 12465 -17290
rect 13089 -17324 13099 -17290
rect 13099 -17324 13123 -17290
rect 13161 -17324 13167 -17290
rect 13167 -17324 13195 -17290
rect 13233 -17324 13235 -17290
rect 13235 -17324 13267 -17290
rect 13305 -17324 13337 -17290
rect 13337 -17324 13339 -17290
rect 13377 -17324 13405 -17290
rect 13405 -17324 13411 -17290
rect 13449 -17324 13473 -17290
rect 13473 -17324 13483 -17290
rect 14107 -17324 14117 -17290
rect 14117 -17324 14141 -17290
rect 14179 -17324 14185 -17290
rect 14185 -17324 14213 -17290
rect 14251 -17324 14253 -17290
rect 14253 -17324 14285 -17290
rect 14323 -17324 14355 -17290
rect 14355 -17324 14357 -17290
rect 14395 -17324 14423 -17290
rect 14423 -17324 14429 -17290
rect 14467 -17324 14491 -17290
rect 14491 -17324 14501 -17290
rect 15125 -17324 15135 -17290
rect 15135 -17324 15159 -17290
rect 15197 -17324 15203 -17290
rect 15203 -17324 15231 -17290
rect 15269 -17324 15271 -17290
rect 15271 -17324 15303 -17290
rect 15341 -17324 15373 -17290
rect 15373 -17324 15375 -17290
rect 15413 -17324 15441 -17290
rect 15441 -17324 15447 -17290
rect 15485 -17324 15509 -17290
rect 15509 -17324 15519 -17290
rect 16143 -17324 16153 -17290
rect 16153 -17324 16177 -17290
rect 16215 -17324 16221 -17290
rect 16221 -17324 16249 -17290
rect 16287 -17324 16289 -17290
rect 16289 -17324 16321 -17290
rect 16359 -17324 16391 -17290
rect 16391 -17324 16393 -17290
rect 16431 -17324 16459 -17290
rect 16459 -17324 16465 -17290
rect 16503 -17324 16527 -17290
rect 16527 -17324 16537 -17290
rect 17161 -17324 17171 -17290
rect 17171 -17324 17195 -17290
rect 17233 -17324 17239 -17290
rect 17239 -17324 17267 -17290
rect 17305 -17324 17307 -17290
rect 17307 -17324 17339 -17290
rect 17377 -17324 17409 -17290
rect 17409 -17324 17411 -17290
rect 17449 -17324 17477 -17290
rect 17477 -17324 17483 -17290
rect 17521 -17324 17545 -17290
rect 17545 -17324 17555 -17290
rect 18179 -17324 18189 -17290
rect 18189 -17324 18213 -17290
rect 18251 -17324 18257 -17290
rect 18257 -17324 18285 -17290
rect 18323 -17324 18325 -17290
rect 18325 -17324 18357 -17290
rect 18395 -17324 18427 -17290
rect 18427 -17324 18429 -17290
rect 18467 -17324 18495 -17290
rect 18495 -17324 18501 -17290
rect 18539 -17324 18563 -17290
rect 18563 -17324 18573 -17290
rect 19197 -17324 19207 -17290
rect 19207 -17324 19231 -17290
rect 19269 -17324 19275 -17290
rect 19275 -17324 19303 -17290
rect 19341 -17324 19343 -17290
rect 19343 -17324 19375 -17290
rect 19413 -17324 19445 -17290
rect 19445 -17324 19447 -17290
rect 19485 -17324 19513 -17290
rect 19513 -17324 19519 -17290
rect 19557 -17324 19581 -17290
rect 19581 -17324 19591 -17290
rect 20215 -17324 20225 -17290
rect 20225 -17324 20249 -17290
rect 20287 -17324 20293 -17290
rect 20293 -17324 20321 -17290
rect 20359 -17324 20361 -17290
rect 20361 -17324 20393 -17290
rect 20431 -17324 20463 -17290
rect 20463 -17324 20465 -17290
rect 20503 -17324 20531 -17290
rect 20531 -17324 20537 -17290
rect 20575 -17324 20599 -17290
rect 20599 -17324 20609 -17290
rect 21233 -17324 21243 -17290
rect 21243 -17324 21267 -17290
rect 21305 -17324 21311 -17290
rect 21311 -17324 21339 -17290
rect 21521 -17324 21549 -17290
rect 21549 -17324 21555 -17290
rect 21593 -17324 21617 -17290
rect 21617 -17324 21627 -17290
rect 22251 -17324 22261 -17290
rect 22261 -17324 22285 -17290
rect 22323 -17324 22329 -17290
rect 22329 -17324 22357 -17290
rect 22395 -17324 22397 -17290
rect 22397 -17324 22429 -17290
rect 22467 -17324 22499 -17290
rect 22499 -17324 22501 -17290
rect 22539 -17324 22567 -17290
rect 22567 -17324 22573 -17290
rect 22611 -17324 22635 -17290
rect 22635 -17324 22645 -17290
rect 24855 -17279 24889 -17275
rect 24855 -17309 24889 -17279
rect -12289 -17381 -12255 -17347
rect -8855 -17382 -8845 -17348
rect -8845 -17382 -8821 -17348
rect -8783 -17382 -8777 -17348
rect -8777 -17382 -8749 -17348
rect -8711 -17382 -8709 -17348
rect -8709 -17382 -8677 -17348
rect -8639 -17382 -8607 -17348
rect -8607 -17382 -8605 -17348
rect -8567 -17382 -8539 -17348
rect -8539 -17382 -8533 -17348
rect -8495 -17382 -8471 -17348
rect -8471 -17382 -8461 -17348
rect -7837 -17382 -7827 -17348
rect -7827 -17382 -7803 -17348
rect -7765 -17382 -7759 -17348
rect -7759 -17382 -7731 -17348
rect -7693 -17382 -7691 -17348
rect -7691 -17382 -7659 -17348
rect -7621 -17382 -7589 -17348
rect -7589 -17382 -7587 -17348
rect -7549 -17382 -7521 -17348
rect -7521 -17382 -7515 -17348
rect -7477 -17382 -7453 -17348
rect -7453 -17382 -7443 -17348
rect -6819 -17382 -6809 -17348
rect -6809 -17382 -6785 -17348
rect -6747 -17382 -6741 -17348
rect -6741 -17382 -6713 -17348
rect -6675 -17382 -6673 -17348
rect -6673 -17382 -6641 -17348
rect -6603 -17382 -6571 -17348
rect -6571 -17382 -6569 -17348
rect -6531 -17382 -6503 -17348
rect -6503 -17382 -6497 -17348
rect -6459 -17382 -6435 -17348
rect -6435 -17382 -6425 -17348
rect -5801 -17382 -5791 -17348
rect -5791 -17382 -5767 -17348
rect -5729 -17382 -5723 -17348
rect -5723 -17382 -5695 -17348
rect -5657 -17382 -5655 -17348
rect -5655 -17382 -5623 -17348
rect -5585 -17382 -5553 -17348
rect -5553 -17382 -5551 -17348
rect -5513 -17382 -5485 -17348
rect -5485 -17382 -5479 -17348
rect -5441 -17382 -5417 -17348
rect -5417 -17382 -5407 -17348
rect -4783 -17382 -4773 -17348
rect -4773 -17382 -4749 -17348
rect -4711 -17382 -4705 -17348
rect -4705 -17382 -4677 -17348
rect -4639 -17382 -4637 -17348
rect -4637 -17382 -4605 -17348
rect -4567 -17382 -4535 -17348
rect -4535 -17382 -4533 -17348
rect -4495 -17382 -4467 -17348
rect -4467 -17382 -4461 -17348
rect -4423 -17382 -4399 -17348
rect -4399 -17382 -4389 -17348
rect -3765 -17382 -3755 -17348
rect -3755 -17382 -3731 -17348
rect -3693 -17382 -3687 -17348
rect -3687 -17382 -3659 -17348
rect -3621 -17382 -3619 -17348
rect -3619 -17382 -3587 -17348
rect -3549 -17382 -3517 -17348
rect -3517 -17382 -3515 -17348
rect -3477 -17382 -3449 -17348
rect -3449 -17382 -3443 -17348
rect -3405 -17382 -3381 -17348
rect -3381 -17382 -3371 -17348
rect -2747 -17382 -2737 -17348
rect -2737 -17382 -2713 -17348
rect -2675 -17382 -2669 -17348
rect -2669 -17382 -2641 -17348
rect -2603 -17382 -2601 -17348
rect -2601 -17382 -2569 -17348
rect -2531 -17382 -2499 -17348
rect -2499 -17382 -2497 -17348
rect -2459 -17382 -2431 -17348
rect -2431 -17382 -2425 -17348
rect -2387 -17382 -2363 -17348
rect -2363 -17382 -2353 -17348
rect -1729 -17382 -1719 -17348
rect -1719 -17382 -1695 -17348
rect -1657 -17382 -1651 -17348
rect -1651 -17382 -1623 -17348
rect -1585 -17382 -1583 -17348
rect -1583 -17382 -1551 -17348
rect -1513 -17382 -1481 -17348
rect -1481 -17382 -1479 -17348
rect -1441 -17382 -1413 -17348
rect -1413 -17382 -1407 -17348
rect -1369 -17382 -1345 -17348
rect -1345 -17382 -1335 -17348
rect -711 -17382 -701 -17348
rect -701 -17382 -677 -17348
rect -639 -17382 -633 -17348
rect -633 -17382 -605 -17348
rect -567 -17382 -565 -17348
rect -565 -17382 -533 -17348
rect -495 -17382 -463 -17348
rect -463 -17382 -461 -17348
rect -423 -17382 -395 -17348
rect -395 -17382 -389 -17348
rect -351 -17382 -327 -17348
rect -327 -17382 -317 -17348
rect 24855 -17381 24889 -17347
rect -12289 -17449 -12255 -17419
rect -12289 -17453 -12255 -17449
rect -12289 -17517 -12255 -17491
rect -12289 -17525 -12255 -17517
rect -12289 -17585 -12255 -17563
rect -12289 -17597 -12255 -17585
rect -12289 -17653 -12255 -17635
rect -12289 -17669 -12255 -17653
rect -12289 -17721 -12255 -17707
rect -12289 -17741 -12255 -17721
rect -12289 -17789 -12255 -17779
rect -12289 -17813 -12255 -17789
rect -12289 -17857 -12255 -17851
rect -12289 -17885 -12255 -17857
rect -12289 -17925 -12255 -17923
rect -12289 -17957 -12255 -17925
rect -12289 -18027 -12255 -17995
rect -12289 -18029 -12255 -18027
rect -9184 -17465 -9150 -17451
rect -9184 -17485 -9150 -17465
rect -9184 -17533 -9150 -17523
rect -9184 -17557 -9150 -17533
rect -9184 -17601 -9150 -17595
rect -9184 -17629 -9150 -17601
rect -9184 -17669 -9150 -17667
rect -9184 -17701 -9150 -17669
rect -9184 -17771 -9150 -17739
rect -9184 -17773 -9150 -17771
rect -9184 -17839 -9150 -17811
rect -9184 -17845 -9150 -17839
rect -9184 -17907 -9150 -17883
rect -9184 -17917 -9150 -17907
rect -9184 -17975 -9150 -17955
rect -9184 -17989 -9150 -17975
rect -8166 -17465 -8132 -17451
rect -8166 -17485 -8132 -17465
rect -8166 -17533 -8132 -17523
rect -8166 -17557 -8132 -17533
rect -8166 -17601 -8132 -17595
rect -8166 -17629 -8132 -17601
rect -8166 -17669 -8132 -17667
rect -8166 -17701 -8132 -17669
rect -8166 -17771 -8132 -17739
rect -8166 -17773 -8132 -17771
rect -8166 -17839 -8132 -17811
rect -8166 -17845 -8132 -17839
rect -8166 -17907 -8132 -17883
rect -8166 -17917 -8132 -17907
rect -8166 -17975 -8132 -17955
rect -8166 -17989 -8132 -17975
rect -7148 -17465 -7114 -17451
rect -7148 -17485 -7114 -17465
rect -7148 -17533 -7114 -17523
rect -7148 -17557 -7114 -17533
rect -7148 -17601 -7114 -17595
rect -7148 -17629 -7114 -17601
rect -7148 -17669 -7114 -17667
rect -7148 -17701 -7114 -17669
rect -7148 -17771 -7114 -17739
rect -7148 -17773 -7114 -17771
rect -7148 -17839 -7114 -17811
rect -7148 -17845 -7114 -17839
rect -7148 -17907 -7114 -17883
rect -7148 -17917 -7114 -17907
rect -7148 -17975 -7114 -17955
rect -7148 -17989 -7114 -17975
rect -6130 -17465 -6096 -17451
rect -6130 -17485 -6096 -17465
rect -6130 -17533 -6096 -17523
rect -6130 -17557 -6096 -17533
rect -6130 -17601 -6096 -17595
rect -6130 -17629 -6096 -17601
rect -6130 -17669 -6096 -17667
rect -6130 -17701 -6096 -17669
rect -6130 -17771 -6096 -17739
rect -6130 -17773 -6096 -17771
rect -6130 -17839 -6096 -17811
rect -6130 -17845 -6096 -17839
rect -6130 -17907 -6096 -17883
rect -6130 -17917 -6096 -17907
rect -6130 -17975 -6096 -17955
rect -6130 -17989 -6096 -17975
rect -5112 -17465 -5078 -17451
rect -5112 -17485 -5078 -17465
rect -5112 -17533 -5078 -17523
rect -5112 -17557 -5078 -17533
rect -5112 -17601 -5078 -17595
rect -5112 -17629 -5078 -17601
rect -5112 -17669 -5078 -17667
rect -5112 -17701 -5078 -17669
rect -5112 -17771 -5078 -17739
rect -5112 -17773 -5078 -17771
rect -5112 -17839 -5078 -17811
rect -5112 -17845 -5078 -17839
rect -5112 -17907 -5078 -17883
rect -5112 -17917 -5078 -17907
rect -5112 -17975 -5078 -17955
rect -5112 -17989 -5078 -17975
rect -4094 -17465 -4060 -17451
rect -4094 -17485 -4060 -17465
rect -4094 -17533 -4060 -17523
rect -4094 -17557 -4060 -17533
rect -4094 -17601 -4060 -17595
rect -4094 -17629 -4060 -17601
rect -4094 -17669 -4060 -17667
rect -4094 -17701 -4060 -17669
rect -4094 -17771 -4060 -17739
rect -4094 -17773 -4060 -17771
rect -4094 -17839 -4060 -17811
rect -4094 -17845 -4060 -17839
rect -4094 -17907 -4060 -17883
rect -4094 -17917 -4060 -17907
rect -4094 -17975 -4060 -17955
rect -4094 -17989 -4060 -17975
rect -3076 -17465 -3042 -17451
rect -3076 -17485 -3042 -17465
rect -3076 -17533 -3042 -17523
rect -3076 -17557 -3042 -17533
rect -3076 -17601 -3042 -17595
rect -3076 -17629 -3042 -17601
rect -3076 -17669 -3042 -17667
rect -3076 -17701 -3042 -17669
rect -3076 -17771 -3042 -17739
rect -3076 -17773 -3042 -17771
rect -3076 -17839 -3042 -17811
rect -3076 -17845 -3042 -17839
rect -3076 -17907 -3042 -17883
rect -3076 -17917 -3042 -17907
rect -3076 -17975 -3042 -17955
rect -3076 -17989 -3042 -17975
rect -2058 -17465 -2024 -17451
rect -2058 -17485 -2024 -17465
rect -2058 -17533 -2024 -17523
rect -2058 -17557 -2024 -17533
rect -2058 -17601 -2024 -17595
rect -2058 -17629 -2024 -17601
rect -2058 -17669 -2024 -17667
rect -2058 -17701 -2024 -17669
rect -2058 -17771 -2024 -17739
rect -2058 -17773 -2024 -17771
rect -2058 -17839 -2024 -17811
rect -2058 -17845 -2024 -17839
rect -2058 -17907 -2024 -17883
rect -2058 -17917 -2024 -17907
rect -2058 -17975 -2024 -17955
rect -2058 -17989 -2024 -17975
rect -1040 -17465 -1006 -17451
rect -1040 -17485 -1006 -17465
rect -1040 -17533 -1006 -17523
rect -1040 -17557 -1006 -17533
rect -1040 -17601 -1006 -17595
rect -1040 -17629 -1006 -17601
rect -1040 -17669 -1006 -17667
rect -1040 -17701 -1006 -17669
rect -1040 -17771 -1006 -17739
rect -1040 -17773 -1006 -17771
rect -1040 -17839 -1006 -17811
rect -1040 -17845 -1006 -17839
rect -1040 -17907 -1006 -17883
rect -1040 -17917 -1006 -17907
rect -1040 -17975 -1006 -17955
rect -1040 -17989 -1006 -17975
rect -22 -17465 12 -17451
rect -22 -17485 12 -17465
rect -22 -17533 12 -17523
rect -22 -17557 12 -17533
rect -22 -17601 12 -17595
rect -22 -17629 12 -17601
rect -22 -17669 12 -17667
rect -22 -17701 12 -17669
rect -22 -17771 12 -17739
rect -22 -17773 12 -17771
rect -22 -17839 12 -17811
rect 24855 -17449 24889 -17419
rect 24855 -17453 24889 -17449
rect 24855 -17517 24889 -17491
rect 24855 -17525 24889 -17517
rect 24855 -17585 24889 -17563
rect 24855 -17597 24889 -17585
rect 24855 -17653 24889 -17635
rect 24855 -17669 24889 -17653
rect 24855 -17721 24889 -17707
rect 24855 -17741 24889 -17721
rect -22 -17845 12 -17839
rect 2909 -17846 2919 -17812
rect 2919 -17846 2943 -17812
rect 2981 -17846 2987 -17812
rect 2987 -17846 3015 -17812
rect 3053 -17846 3055 -17812
rect 3055 -17846 3087 -17812
rect 3125 -17846 3157 -17812
rect 3157 -17846 3159 -17812
rect 3197 -17846 3225 -17812
rect 3225 -17846 3231 -17812
rect 3269 -17846 3293 -17812
rect 3293 -17846 3303 -17812
rect 3927 -17846 3937 -17812
rect 3937 -17846 3961 -17812
rect 3999 -17846 4005 -17812
rect 4005 -17846 4033 -17812
rect 4071 -17846 4073 -17812
rect 4073 -17846 4105 -17812
rect 4143 -17846 4175 -17812
rect 4175 -17846 4177 -17812
rect 4215 -17846 4243 -17812
rect 4243 -17846 4249 -17812
rect 4287 -17846 4311 -17812
rect 4311 -17846 4321 -17812
rect 4945 -17846 4955 -17812
rect 4955 -17846 4979 -17812
rect 5017 -17846 5023 -17812
rect 5023 -17846 5051 -17812
rect 5089 -17846 5091 -17812
rect 5091 -17846 5123 -17812
rect 5161 -17846 5193 -17812
rect 5193 -17846 5195 -17812
rect 5233 -17846 5261 -17812
rect 5261 -17846 5267 -17812
rect 5305 -17846 5329 -17812
rect 5329 -17846 5339 -17812
rect 5963 -17846 5973 -17812
rect 5973 -17846 5997 -17812
rect 6035 -17846 6041 -17812
rect 6041 -17846 6069 -17812
rect 6107 -17846 6109 -17812
rect 6109 -17846 6141 -17812
rect 6179 -17846 6211 -17812
rect 6211 -17846 6213 -17812
rect 6251 -17846 6279 -17812
rect 6279 -17846 6285 -17812
rect 6323 -17846 6347 -17812
rect 6347 -17846 6357 -17812
rect 6981 -17846 6991 -17812
rect 6991 -17846 7015 -17812
rect 7053 -17846 7059 -17812
rect 7059 -17846 7087 -17812
rect 7125 -17846 7127 -17812
rect 7127 -17846 7159 -17812
rect 7197 -17846 7229 -17812
rect 7229 -17846 7231 -17812
rect 7269 -17846 7297 -17812
rect 7297 -17846 7303 -17812
rect 7341 -17846 7365 -17812
rect 7365 -17846 7375 -17812
rect 7999 -17846 8009 -17812
rect 8009 -17846 8033 -17812
rect 8071 -17846 8077 -17812
rect 8077 -17846 8105 -17812
rect 8143 -17846 8145 -17812
rect 8145 -17846 8177 -17812
rect 8215 -17846 8247 -17812
rect 8247 -17846 8249 -17812
rect 8287 -17846 8315 -17812
rect 8315 -17846 8321 -17812
rect 8359 -17846 8383 -17812
rect 8383 -17846 8393 -17812
rect 9017 -17846 9027 -17812
rect 9027 -17846 9051 -17812
rect 9089 -17846 9095 -17812
rect 9095 -17846 9123 -17812
rect 9161 -17846 9163 -17812
rect 9163 -17846 9195 -17812
rect 9233 -17846 9265 -17812
rect 9265 -17846 9267 -17812
rect 9305 -17846 9333 -17812
rect 9333 -17846 9339 -17812
rect 9377 -17846 9401 -17812
rect 9401 -17846 9411 -17812
rect 10035 -17846 10045 -17812
rect 10045 -17846 10069 -17812
rect 10107 -17846 10113 -17812
rect 10113 -17846 10141 -17812
rect 10179 -17846 10181 -17812
rect 10181 -17846 10213 -17812
rect 10251 -17846 10283 -17812
rect 10283 -17846 10285 -17812
rect 10323 -17846 10351 -17812
rect 10351 -17846 10357 -17812
rect 10395 -17846 10419 -17812
rect 10419 -17846 10429 -17812
rect 11053 -17846 11063 -17812
rect 11063 -17846 11087 -17812
rect 11125 -17846 11131 -17812
rect 11131 -17846 11159 -17812
rect 11197 -17846 11199 -17812
rect 11199 -17846 11231 -17812
rect 11269 -17846 11301 -17812
rect 11301 -17846 11303 -17812
rect 11341 -17846 11369 -17812
rect 11369 -17846 11375 -17812
rect 11413 -17846 11437 -17812
rect 11437 -17846 11447 -17812
rect 12071 -17846 12081 -17812
rect 12081 -17846 12105 -17812
rect 12143 -17846 12149 -17812
rect 12149 -17846 12177 -17812
rect 12215 -17846 12217 -17812
rect 12217 -17846 12249 -17812
rect 12287 -17846 12319 -17812
rect 12319 -17846 12321 -17812
rect 12359 -17846 12387 -17812
rect 12387 -17846 12393 -17812
rect 12431 -17846 12455 -17812
rect 12455 -17846 12465 -17812
rect 13089 -17846 13099 -17812
rect 13099 -17846 13123 -17812
rect 13161 -17846 13167 -17812
rect 13167 -17846 13195 -17812
rect 13233 -17846 13235 -17812
rect 13235 -17846 13267 -17812
rect 13305 -17846 13337 -17812
rect 13337 -17846 13339 -17812
rect 13377 -17846 13405 -17812
rect 13405 -17846 13411 -17812
rect 13449 -17846 13473 -17812
rect 13473 -17846 13483 -17812
rect 14107 -17846 14117 -17812
rect 14117 -17846 14141 -17812
rect 14179 -17846 14185 -17812
rect 14185 -17846 14213 -17812
rect 14251 -17846 14253 -17812
rect 14253 -17846 14285 -17812
rect 14323 -17846 14355 -17812
rect 14355 -17846 14357 -17812
rect 14395 -17846 14423 -17812
rect 14423 -17846 14429 -17812
rect 14467 -17846 14491 -17812
rect 14491 -17846 14501 -17812
rect 15125 -17846 15135 -17812
rect 15135 -17846 15159 -17812
rect 15197 -17846 15203 -17812
rect 15203 -17846 15231 -17812
rect 15269 -17846 15271 -17812
rect 15271 -17846 15303 -17812
rect 15341 -17846 15373 -17812
rect 15373 -17846 15375 -17812
rect 15413 -17846 15441 -17812
rect 15441 -17846 15447 -17812
rect 15485 -17846 15509 -17812
rect 15509 -17846 15519 -17812
rect 16143 -17846 16153 -17812
rect 16153 -17846 16177 -17812
rect 16215 -17846 16221 -17812
rect 16221 -17846 16249 -17812
rect 16287 -17846 16289 -17812
rect 16289 -17846 16321 -17812
rect 16359 -17846 16391 -17812
rect 16391 -17846 16393 -17812
rect 16431 -17846 16459 -17812
rect 16459 -17846 16465 -17812
rect 16503 -17846 16527 -17812
rect 16527 -17846 16537 -17812
rect 17161 -17846 17171 -17812
rect 17171 -17846 17195 -17812
rect 17233 -17846 17239 -17812
rect 17239 -17846 17267 -17812
rect 17305 -17846 17307 -17812
rect 17307 -17846 17339 -17812
rect 17377 -17846 17409 -17812
rect 17409 -17846 17411 -17812
rect 17449 -17846 17477 -17812
rect 17477 -17846 17483 -17812
rect 17521 -17846 17545 -17812
rect 17545 -17846 17555 -17812
rect 18179 -17846 18189 -17812
rect 18189 -17846 18213 -17812
rect 18251 -17846 18257 -17812
rect 18257 -17846 18285 -17812
rect 18323 -17846 18325 -17812
rect 18325 -17846 18357 -17812
rect 18395 -17846 18427 -17812
rect 18427 -17846 18429 -17812
rect 18467 -17846 18495 -17812
rect 18495 -17846 18501 -17812
rect 18539 -17846 18563 -17812
rect 18563 -17846 18573 -17812
rect 19197 -17846 19207 -17812
rect 19207 -17846 19231 -17812
rect 19269 -17846 19275 -17812
rect 19275 -17846 19303 -17812
rect 19341 -17846 19343 -17812
rect 19343 -17846 19375 -17812
rect 19413 -17846 19445 -17812
rect 19445 -17846 19447 -17812
rect 19485 -17846 19513 -17812
rect 19513 -17846 19519 -17812
rect 19557 -17846 19581 -17812
rect 19581 -17846 19591 -17812
rect 20215 -17846 20225 -17812
rect 20225 -17846 20249 -17812
rect 20287 -17846 20293 -17812
rect 20293 -17846 20321 -17812
rect 20359 -17846 20361 -17812
rect 20361 -17846 20393 -17812
rect 20431 -17846 20463 -17812
rect 20463 -17846 20465 -17812
rect 20503 -17846 20531 -17812
rect 20531 -17846 20537 -17812
rect 20575 -17846 20599 -17812
rect 20599 -17846 20609 -17812
rect 21233 -17846 21243 -17812
rect 21243 -17846 21267 -17812
rect 21305 -17846 21311 -17812
rect 21311 -17846 21339 -17812
rect 21377 -17846 21379 -17812
rect 21379 -17846 21411 -17812
rect 21449 -17846 21481 -17812
rect 21481 -17846 21483 -17812
rect 21521 -17846 21549 -17812
rect 21549 -17846 21555 -17812
rect 21593 -17846 21617 -17812
rect 21617 -17846 21627 -17812
rect 22251 -17846 22261 -17812
rect 22261 -17846 22285 -17812
rect 22323 -17846 22329 -17812
rect 22329 -17846 22357 -17812
rect 22395 -17846 22397 -17812
rect 22397 -17846 22429 -17812
rect 22467 -17846 22499 -17812
rect 22499 -17846 22501 -17812
rect 22539 -17846 22567 -17812
rect 22567 -17846 22573 -17812
rect 22611 -17846 22635 -17812
rect 22635 -17846 22645 -17812
rect 24855 -17789 24889 -17779
rect 24855 -17813 24889 -17789
rect -22 -17907 12 -17883
rect -22 -17917 12 -17907
rect -22 -17975 12 -17955
rect -22 -17989 12 -17975
rect 2580 -17929 2614 -17915
rect 2580 -17949 2614 -17929
rect 2580 -17997 2614 -17987
rect 2580 -18021 2614 -17997
rect -12289 -18095 -12255 -18067
rect -12289 -18101 -12255 -18095
rect -8855 -18092 -8845 -18058
rect -8845 -18092 -8821 -18058
rect -8783 -18092 -8777 -18058
rect -8777 -18092 -8749 -18058
rect -8711 -18092 -8709 -18058
rect -8709 -18092 -8677 -18058
rect -8639 -18092 -8607 -18058
rect -8607 -18092 -8605 -18058
rect -8567 -18092 -8539 -18058
rect -8539 -18092 -8533 -18058
rect -8495 -18092 -8471 -18058
rect -8471 -18092 -8461 -18058
rect -7837 -18092 -7827 -18058
rect -7827 -18092 -7803 -18058
rect -7765 -18092 -7759 -18058
rect -7759 -18092 -7731 -18058
rect -7693 -18092 -7691 -18058
rect -7691 -18092 -7659 -18058
rect -7621 -18092 -7589 -18058
rect -7589 -18092 -7587 -18058
rect -7549 -18092 -7521 -18058
rect -7521 -18092 -7515 -18058
rect -7477 -18092 -7453 -18058
rect -7453 -18092 -7443 -18058
rect -6819 -18092 -6809 -18058
rect -6809 -18092 -6785 -18058
rect -6747 -18092 -6741 -18058
rect -6741 -18092 -6713 -18058
rect -6675 -18092 -6673 -18058
rect -6673 -18092 -6641 -18058
rect -6603 -18092 -6571 -18058
rect -6571 -18092 -6569 -18058
rect -6531 -18092 -6503 -18058
rect -6503 -18092 -6497 -18058
rect -6459 -18092 -6435 -18058
rect -6435 -18092 -6425 -18058
rect -5801 -18092 -5791 -18058
rect -5791 -18092 -5767 -18058
rect -5729 -18092 -5723 -18058
rect -5723 -18092 -5695 -18058
rect -5657 -18092 -5655 -18058
rect -5655 -18092 -5623 -18058
rect -5585 -18092 -5553 -18058
rect -5553 -18092 -5551 -18058
rect -5513 -18092 -5485 -18058
rect -5485 -18092 -5479 -18058
rect -5441 -18092 -5417 -18058
rect -5417 -18092 -5407 -18058
rect -4783 -18092 -4773 -18058
rect -4773 -18092 -4749 -18058
rect -4711 -18092 -4705 -18058
rect -4705 -18092 -4677 -18058
rect -4639 -18092 -4637 -18058
rect -4637 -18092 -4605 -18058
rect -4567 -18092 -4535 -18058
rect -4535 -18092 -4533 -18058
rect -4495 -18092 -4467 -18058
rect -4467 -18092 -4461 -18058
rect -4423 -18092 -4399 -18058
rect -4399 -18092 -4389 -18058
rect -3765 -18092 -3755 -18058
rect -3755 -18092 -3731 -18058
rect -3693 -18092 -3687 -18058
rect -3687 -18092 -3659 -18058
rect -3621 -18092 -3619 -18058
rect -3619 -18092 -3587 -18058
rect -3549 -18092 -3517 -18058
rect -3517 -18092 -3515 -18058
rect -3477 -18092 -3449 -18058
rect -3449 -18092 -3443 -18058
rect -3405 -18092 -3381 -18058
rect -3381 -18092 -3371 -18058
rect -2747 -18092 -2737 -18058
rect -2737 -18092 -2713 -18058
rect -2675 -18092 -2669 -18058
rect -2669 -18092 -2641 -18058
rect -2603 -18092 -2601 -18058
rect -2601 -18092 -2569 -18058
rect -2531 -18092 -2499 -18058
rect -2499 -18092 -2497 -18058
rect -2459 -18092 -2431 -18058
rect -2431 -18092 -2425 -18058
rect -2387 -18092 -2363 -18058
rect -2363 -18092 -2353 -18058
rect -1729 -18092 -1719 -18058
rect -1719 -18092 -1695 -18058
rect -1657 -18092 -1651 -18058
rect -1651 -18092 -1623 -18058
rect -1585 -18092 -1583 -18058
rect -1583 -18092 -1551 -18058
rect -1513 -18092 -1481 -18058
rect -1481 -18092 -1479 -18058
rect -1441 -18092 -1413 -18058
rect -1413 -18092 -1407 -18058
rect -1369 -18092 -1345 -18058
rect -1345 -18092 -1335 -18058
rect -711 -18092 -701 -18058
rect -701 -18092 -677 -18058
rect -639 -18092 -633 -18058
rect -633 -18092 -605 -18058
rect -567 -18092 -565 -18058
rect -565 -18092 -533 -18058
rect -495 -18092 -463 -18058
rect -463 -18092 -461 -18058
rect -423 -18092 -395 -18058
rect -395 -18092 -389 -18058
rect -351 -18092 -327 -18058
rect -327 -18092 -317 -18058
rect 2580 -18065 2614 -18059
rect -12289 -18163 -12255 -18139
rect -12289 -18173 -12255 -18163
rect 2580 -18093 2614 -18065
rect 2580 -18133 2614 -18131
rect 2580 -18165 2614 -18133
rect -8855 -18200 -8845 -18166
rect -8845 -18200 -8821 -18166
rect -8783 -18200 -8777 -18166
rect -8777 -18200 -8749 -18166
rect -8711 -18200 -8709 -18166
rect -8709 -18200 -8677 -18166
rect -8639 -18200 -8607 -18166
rect -8607 -18200 -8605 -18166
rect -8567 -18200 -8539 -18166
rect -8539 -18200 -8533 -18166
rect -8495 -18200 -8471 -18166
rect -8471 -18200 -8461 -18166
rect -7837 -18200 -7827 -18166
rect -7827 -18200 -7803 -18166
rect -7765 -18200 -7759 -18166
rect -7759 -18200 -7731 -18166
rect -7693 -18200 -7691 -18166
rect -7691 -18200 -7659 -18166
rect -7621 -18200 -7589 -18166
rect -7589 -18200 -7587 -18166
rect -7549 -18200 -7521 -18166
rect -7521 -18200 -7515 -18166
rect -7477 -18200 -7453 -18166
rect -7453 -18200 -7443 -18166
rect -6819 -18200 -6809 -18166
rect -6809 -18200 -6785 -18166
rect -6747 -18200 -6741 -18166
rect -6741 -18200 -6713 -18166
rect -6675 -18200 -6673 -18166
rect -6673 -18200 -6641 -18166
rect -6603 -18200 -6571 -18166
rect -6571 -18200 -6569 -18166
rect -6531 -18200 -6503 -18166
rect -6503 -18200 -6497 -18166
rect -6459 -18200 -6435 -18166
rect -6435 -18200 -6425 -18166
rect -5801 -18200 -5791 -18166
rect -5791 -18200 -5767 -18166
rect -5729 -18200 -5723 -18166
rect -5723 -18200 -5695 -18166
rect -5657 -18200 -5655 -18166
rect -5655 -18200 -5623 -18166
rect -5585 -18200 -5553 -18166
rect -5553 -18200 -5551 -18166
rect -5513 -18200 -5485 -18166
rect -5485 -18200 -5479 -18166
rect -5441 -18200 -5417 -18166
rect -5417 -18200 -5407 -18166
rect -4783 -18200 -4773 -18166
rect -4773 -18200 -4749 -18166
rect -4711 -18200 -4705 -18166
rect -4705 -18200 -4677 -18166
rect -4639 -18200 -4637 -18166
rect -4637 -18200 -4605 -18166
rect -4567 -18200 -4535 -18166
rect -4535 -18200 -4533 -18166
rect -4495 -18200 -4467 -18166
rect -4467 -18200 -4461 -18166
rect -4423 -18200 -4399 -18166
rect -4399 -18200 -4389 -18166
rect -3765 -18200 -3755 -18166
rect -3755 -18200 -3731 -18166
rect -3693 -18200 -3687 -18166
rect -3687 -18200 -3659 -18166
rect -3621 -18200 -3619 -18166
rect -3619 -18200 -3587 -18166
rect -3549 -18200 -3517 -18166
rect -3517 -18200 -3515 -18166
rect -3477 -18200 -3449 -18166
rect -3449 -18200 -3443 -18166
rect -3405 -18200 -3381 -18166
rect -3381 -18200 -3371 -18166
rect -2747 -18200 -2737 -18166
rect -2737 -18200 -2713 -18166
rect -2675 -18200 -2669 -18166
rect -2669 -18200 -2641 -18166
rect -2603 -18200 -2601 -18166
rect -2601 -18200 -2569 -18166
rect -2531 -18200 -2499 -18166
rect -2499 -18200 -2497 -18166
rect -2459 -18200 -2431 -18166
rect -2431 -18200 -2425 -18166
rect -2387 -18200 -2363 -18166
rect -2363 -18200 -2353 -18166
rect -1729 -18200 -1719 -18166
rect -1719 -18200 -1695 -18166
rect -1657 -18200 -1651 -18166
rect -1651 -18200 -1623 -18166
rect -1585 -18200 -1583 -18166
rect -1583 -18200 -1551 -18166
rect -1513 -18200 -1481 -18166
rect -1481 -18200 -1479 -18166
rect -1441 -18200 -1413 -18166
rect -1413 -18200 -1407 -18166
rect -1369 -18200 -1345 -18166
rect -1345 -18200 -1335 -18166
rect -711 -18200 -701 -18166
rect -701 -18200 -677 -18166
rect -639 -18200 -633 -18166
rect -633 -18200 -605 -18166
rect -567 -18200 -565 -18166
rect -565 -18200 -533 -18166
rect -495 -18200 -463 -18166
rect -463 -18200 -461 -18166
rect -423 -18200 -395 -18166
rect -395 -18200 -389 -18166
rect -351 -18200 -327 -18166
rect -327 -18200 -317 -18166
rect -12289 -18231 -12255 -18211
rect -12289 -18245 -12255 -18231
rect -12289 -18299 -12255 -18283
rect -12289 -18317 -12255 -18299
rect -12289 -18367 -12255 -18355
rect -12289 -18389 -12255 -18367
rect -12289 -18435 -12255 -18427
rect -12289 -18461 -12255 -18435
rect -12289 -18503 -12255 -18499
rect -12289 -18533 -12255 -18503
rect -12289 -18605 -12255 -18571
rect -12289 -18673 -12255 -18643
rect -12289 -18677 -12255 -18673
rect -12289 -18741 -12255 -18715
rect -12289 -18749 -12255 -18741
rect -12289 -18809 -12255 -18787
rect -12289 -18821 -12255 -18809
rect -9184 -18283 -9150 -18269
rect -9184 -18303 -9150 -18283
rect -9184 -18351 -9150 -18341
rect -9184 -18375 -9150 -18351
rect -9184 -18419 -9150 -18413
rect -9184 -18447 -9150 -18419
rect -9184 -18487 -9150 -18485
rect -9184 -18519 -9150 -18487
rect -9184 -18589 -9150 -18557
rect -9184 -18591 -9150 -18589
rect -9184 -18657 -9150 -18629
rect -9184 -18663 -9150 -18657
rect -9184 -18725 -9150 -18701
rect -9184 -18735 -9150 -18725
rect -9184 -18793 -9150 -18773
rect -9184 -18807 -9150 -18793
rect -8166 -18283 -8132 -18269
rect -8166 -18303 -8132 -18283
rect -8166 -18351 -8132 -18341
rect -8166 -18375 -8132 -18351
rect -8166 -18419 -8132 -18413
rect -8166 -18447 -8132 -18419
rect -8166 -18487 -8132 -18485
rect -8166 -18519 -8132 -18487
rect -8166 -18589 -8132 -18557
rect -8166 -18591 -8132 -18589
rect -8166 -18657 -8132 -18629
rect -8166 -18663 -8132 -18657
rect -8166 -18725 -8132 -18701
rect -8166 -18735 -8132 -18725
rect -8166 -18793 -8132 -18773
rect -8166 -18807 -8132 -18793
rect -7148 -18283 -7114 -18269
rect -7148 -18303 -7114 -18283
rect -7148 -18351 -7114 -18341
rect -7148 -18375 -7114 -18351
rect -7148 -18419 -7114 -18413
rect -7148 -18447 -7114 -18419
rect -7148 -18487 -7114 -18485
rect -7148 -18519 -7114 -18487
rect -7148 -18589 -7114 -18557
rect -7148 -18591 -7114 -18589
rect -7148 -18657 -7114 -18629
rect -7148 -18663 -7114 -18657
rect -7148 -18725 -7114 -18701
rect -7148 -18735 -7114 -18725
rect -7148 -18793 -7114 -18773
rect -7148 -18807 -7114 -18793
rect -6130 -18283 -6096 -18269
rect -6130 -18303 -6096 -18283
rect -6130 -18351 -6096 -18341
rect -6130 -18375 -6096 -18351
rect -6130 -18419 -6096 -18413
rect -6130 -18447 -6096 -18419
rect -6130 -18487 -6096 -18485
rect -6130 -18519 -6096 -18487
rect -6130 -18589 -6096 -18557
rect -6130 -18591 -6096 -18589
rect -6130 -18657 -6096 -18629
rect -6130 -18663 -6096 -18657
rect -6130 -18725 -6096 -18701
rect -6130 -18735 -6096 -18725
rect -6130 -18793 -6096 -18773
rect -6130 -18807 -6096 -18793
rect -5112 -18283 -5078 -18269
rect -5112 -18303 -5078 -18283
rect -5112 -18351 -5078 -18341
rect -5112 -18375 -5078 -18351
rect -5112 -18419 -5078 -18413
rect -5112 -18447 -5078 -18419
rect -5112 -18487 -5078 -18485
rect -5112 -18519 -5078 -18487
rect -5112 -18589 -5078 -18557
rect -5112 -18591 -5078 -18589
rect -5112 -18657 -5078 -18629
rect -5112 -18663 -5078 -18657
rect -5112 -18725 -5078 -18701
rect -5112 -18735 -5078 -18725
rect -5112 -18793 -5078 -18773
rect -5112 -18807 -5078 -18793
rect -4094 -18283 -4060 -18269
rect -4094 -18303 -4060 -18283
rect -4094 -18351 -4060 -18341
rect -4094 -18375 -4060 -18351
rect -4094 -18419 -4060 -18413
rect -4094 -18447 -4060 -18419
rect -4094 -18487 -4060 -18485
rect -4094 -18519 -4060 -18487
rect -4094 -18589 -4060 -18557
rect -4094 -18591 -4060 -18589
rect -4094 -18657 -4060 -18629
rect -4094 -18663 -4060 -18657
rect -4094 -18725 -4060 -18701
rect -4094 -18735 -4060 -18725
rect -4094 -18793 -4060 -18773
rect -4094 -18807 -4060 -18793
rect -3076 -18283 -3042 -18269
rect -3076 -18303 -3042 -18283
rect -3076 -18351 -3042 -18341
rect -3076 -18375 -3042 -18351
rect -3076 -18419 -3042 -18413
rect -3076 -18447 -3042 -18419
rect -3076 -18487 -3042 -18485
rect -3076 -18519 -3042 -18487
rect -3076 -18589 -3042 -18557
rect -3076 -18591 -3042 -18589
rect -3076 -18657 -3042 -18629
rect -3076 -18663 -3042 -18657
rect -3076 -18725 -3042 -18701
rect -3076 -18735 -3042 -18725
rect -3076 -18793 -3042 -18773
rect -3076 -18807 -3042 -18793
rect -2058 -18283 -2024 -18269
rect -2058 -18303 -2024 -18283
rect -2058 -18351 -2024 -18341
rect -2058 -18375 -2024 -18351
rect -2058 -18419 -2024 -18413
rect -2058 -18447 -2024 -18419
rect -2058 -18487 -2024 -18485
rect -2058 -18519 -2024 -18487
rect -2058 -18589 -2024 -18557
rect -2058 -18591 -2024 -18589
rect -2058 -18657 -2024 -18629
rect -2058 -18663 -2024 -18657
rect -2058 -18725 -2024 -18701
rect -2058 -18735 -2024 -18725
rect -2058 -18793 -2024 -18773
rect -2058 -18807 -2024 -18793
rect -1040 -18283 -1006 -18269
rect -1040 -18303 -1006 -18283
rect -1040 -18351 -1006 -18341
rect -1040 -18375 -1006 -18351
rect -1040 -18419 -1006 -18413
rect -1040 -18447 -1006 -18419
rect -1040 -18487 -1006 -18485
rect -1040 -18519 -1006 -18487
rect -1040 -18589 -1006 -18557
rect -1040 -18591 -1006 -18589
rect -1040 -18657 -1006 -18629
rect -1040 -18663 -1006 -18657
rect -1040 -18725 -1006 -18701
rect -1040 -18735 -1006 -18725
rect -1040 -18793 -1006 -18773
rect -1040 -18807 -1006 -18793
rect -22 -18283 12 -18269
rect -22 -18303 12 -18283
rect -22 -18351 12 -18341
rect -22 -18375 12 -18351
rect -22 -18419 12 -18413
rect -22 -18447 12 -18419
rect -22 -18487 12 -18485
rect -22 -18519 12 -18487
rect 2580 -18235 2614 -18203
rect 2580 -18237 2614 -18235
rect 2580 -18303 2614 -18275
rect 2580 -18309 2614 -18303
rect 2580 -18371 2614 -18347
rect 2580 -18381 2614 -18371
rect 2580 -18439 2614 -18419
rect 2580 -18453 2614 -18439
rect 3598 -17929 3632 -17915
rect 3598 -17949 3632 -17929
rect 3598 -17997 3632 -17987
rect 3598 -18021 3632 -17997
rect 3598 -18065 3632 -18059
rect 3598 -18093 3632 -18065
rect 3598 -18133 3632 -18131
rect 3598 -18165 3632 -18133
rect 3598 -18235 3632 -18203
rect 3598 -18237 3632 -18235
rect 3598 -18303 3632 -18275
rect 3598 -18309 3632 -18303
rect 3598 -18371 3632 -18347
rect 3598 -18381 3632 -18371
rect 3598 -18439 3632 -18419
rect 3598 -18453 3632 -18439
rect 4616 -17929 4650 -17915
rect 4616 -17949 4650 -17929
rect 4616 -17997 4650 -17987
rect 4616 -18021 4650 -17997
rect 4616 -18065 4650 -18059
rect 4616 -18093 4650 -18065
rect 4616 -18133 4650 -18131
rect 4616 -18165 4650 -18133
rect 4616 -18235 4650 -18203
rect 4616 -18237 4650 -18235
rect 4616 -18303 4650 -18275
rect 4616 -18309 4650 -18303
rect 4616 -18371 4650 -18347
rect 4616 -18381 4650 -18371
rect 4616 -18439 4650 -18419
rect 4616 -18453 4650 -18439
rect 5634 -17929 5668 -17915
rect 5634 -17949 5668 -17929
rect 5634 -17997 5668 -17987
rect 5634 -18021 5668 -17997
rect 5634 -18065 5668 -18059
rect 5634 -18093 5668 -18065
rect 5634 -18133 5668 -18131
rect 5634 -18165 5668 -18133
rect 5634 -18235 5668 -18203
rect 5634 -18237 5668 -18235
rect 5634 -18303 5668 -18275
rect 5634 -18309 5668 -18303
rect 5634 -18371 5668 -18347
rect 5634 -18381 5668 -18371
rect 5634 -18439 5668 -18419
rect 5634 -18453 5668 -18439
rect 6652 -17929 6686 -17915
rect 6652 -17949 6686 -17929
rect 6652 -17997 6686 -17987
rect 6652 -18021 6686 -17997
rect 6652 -18065 6686 -18059
rect 6652 -18093 6686 -18065
rect 6652 -18133 6686 -18131
rect 6652 -18165 6686 -18133
rect 6652 -18235 6686 -18203
rect 6652 -18237 6686 -18235
rect 6652 -18303 6686 -18275
rect 6652 -18309 6686 -18303
rect 6652 -18371 6686 -18347
rect 6652 -18381 6686 -18371
rect 6652 -18439 6686 -18419
rect 6652 -18453 6686 -18439
rect 7670 -17929 7704 -17915
rect 7670 -17949 7704 -17929
rect 7670 -17997 7704 -17987
rect 7670 -18021 7704 -17997
rect 7670 -18065 7704 -18059
rect 7670 -18093 7704 -18065
rect 7670 -18133 7704 -18131
rect 7670 -18165 7704 -18133
rect 7670 -18235 7704 -18203
rect 7670 -18237 7704 -18235
rect 7670 -18303 7704 -18275
rect 7670 -18309 7704 -18303
rect 7670 -18371 7704 -18347
rect 7670 -18381 7704 -18371
rect 7670 -18439 7704 -18419
rect 7670 -18453 7704 -18439
rect 8688 -17929 8722 -17915
rect 8688 -17949 8722 -17929
rect 8688 -17997 8722 -17987
rect 8688 -18021 8722 -17997
rect 8688 -18065 8722 -18059
rect 8688 -18093 8722 -18065
rect 8688 -18133 8722 -18131
rect 8688 -18165 8722 -18133
rect 8688 -18235 8722 -18203
rect 8688 -18237 8722 -18235
rect 8688 -18303 8722 -18275
rect 8688 -18309 8722 -18303
rect 8688 -18371 8722 -18347
rect 8688 -18381 8722 -18371
rect 8688 -18439 8722 -18419
rect 8688 -18453 8722 -18439
rect 9706 -17929 9740 -17915
rect 9706 -17949 9740 -17929
rect 9706 -17997 9740 -17987
rect 9706 -18021 9740 -17997
rect 9706 -18065 9740 -18059
rect 9706 -18093 9740 -18065
rect 9706 -18133 9740 -18131
rect 9706 -18165 9740 -18133
rect 9706 -18235 9740 -18203
rect 9706 -18237 9740 -18235
rect 9706 -18303 9740 -18275
rect 9706 -18309 9740 -18303
rect 9706 -18371 9740 -18347
rect 9706 -18381 9740 -18371
rect 9706 -18439 9740 -18419
rect 9706 -18453 9740 -18439
rect 10724 -17929 10758 -17915
rect 10724 -17949 10758 -17929
rect 10724 -17997 10758 -17987
rect 10724 -18021 10758 -17997
rect 10724 -18065 10758 -18059
rect 10724 -18093 10758 -18065
rect 10724 -18133 10758 -18131
rect 10724 -18165 10758 -18133
rect 10724 -18235 10758 -18203
rect 10724 -18237 10758 -18235
rect 10724 -18303 10758 -18275
rect 10724 -18309 10758 -18303
rect 10724 -18371 10758 -18347
rect 10724 -18381 10758 -18371
rect 10724 -18439 10758 -18419
rect 10724 -18453 10758 -18439
rect 11742 -17929 11776 -17915
rect 11742 -17949 11776 -17929
rect 11742 -17997 11776 -17987
rect 11742 -18021 11776 -17997
rect 11742 -18065 11776 -18059
rect 11742 -18093 11776 -18065
rect 11742 -18133 11776 -18131
rect 11742 -18165 11776 -18133
rect 11742 -18235 11776 -18203
rect 11742 -18237 11776 -18235
rect 11742 -18303 11776 -18275
rect 11742 -18309 11776 -18303
rect 11742 -18371 11776 -18347
rect 11742 -18381 11776 -18371
rect 11742 -18439 11776 -18419
rect 11742 -18453 11776 -18439
rect 12760 -17929 12794 -17915
rect 12760 -17949 12794 -17929
rect 12760 -17997 12794 -17987
rect 12760 -18021 12794 -17997
rect 12760 -18065 12794 -18059
rect 12760 -18093 12794 -18065
rect 12760 -18133 12794 -18131
rect 12760 -18165 12794 -18133
rect 12760 -18235 12794 -18203
rect 12760 -18237 12794 -18235
rect 12760 -18303 12794 -18275
rect 12760 -18309 12794 -18303
rect 12760 -18371 12794 -18347
rect 12760 -18381 12794 -18371
rect 12760 -18439 12794 -18419
rect 12760 -18453 12794 -18439
rect 13778 -17929 13812 -17915
rect 13778 -17949 13812 -17929
rect 13778 -17997 13812 -17987
rect 13778 -18021 13812 -17997
rect 13778 -18065 13812 -18059
rect 13778 -18093 13812 -18065
rect 13778 -18133 13812 -18131
rect 13778 -18165 13812 -18133
rect 13778 -18235 13812 -18203
rect 13778 -18237 13812 -18235
rect 13778 -18303 13812 -18275
rect 13778 -18309 13812 -18303
rect 13778 -18371 13812 -18347
rect 13778 -18381 13812 -18371
rect 13778 -18439 13812 -18419
rect 13778 -18453 13812 -18439
rect 14796 -17929 14830 -17915
rect 14796 -17949 14830 -17929
rect 14796 -17997 14830 -17987
rect 14796 -18021 14830 -17997
rect 14796 -18065 14830 -18059
rect 14796 -18093 14830 -18065
rect 14796 -18133 14830 -18131
rect 14796 -18165 14830 -18133
rect 14796 -18235 14830 -18203
rect 14796 -18237 14830 -18235
rect 14796 -18303 14830 -18275
rect 14796 -18309 14830 -18303
rect 14796 -18371 14830 -18347
rect 14796 -18381 14830 -18371
rect 14796 -18439 14830 -18419
rect 14796 -18453 14830 -18439
rect 15814 -17929 15848 -17915
rect 15814 -17949 15848 -17929
rect 15814 -17997 15848 -17987
rect 15814 -18021 15848 -17997
rect 15814 -18065 15848 -18059
rect 15814 -18093 15848 -18065
rect 15814 -18133 15848 -18131
rect 15814 -18165 15848 -18133
rect 15814 -18235 15848 -18203
rect 15814 -18237 15848 -18235
rect 15814 -18303 15848 -18275
rect 15814 -18309 15848 -18303
rect 15814 -18371 15848 -18347
rect 15814 -18381 15848 -18371
rect 15814 -18439 15848 -18419
rect 15814 -18453 15848 -18439
rect 16832 -17929 16866 -17915
rect 16832 -17949 16866 -17929
rect 16832 -17997 16866 -17987
rect 16832 -18021 16866 -17997
rect 16832 -18065 16866 -18059
rect 16832 -18093 16866 -18065
rect 16832 -18133 16866 -18131
rect 16832 -18165 16866 -18133
rect 16832 -18235 16866 -18203
rect 16832 -18237 16866 -18235
rect 16832 -18303 16866 -18275
rect 16832 -18309 16866 -18303
rect 16832 -18371 16866 -18347
rect 16832 -18381 16866 -18371
rect 16832 -18439 16866 -18419
rect 16832 -18453 16866 -18439
rect 17850 -17929 17884 -17915
rect 17850 -17949 17884 -17929
rect 17850 -17997 17884 -17987
rect 17850 -18021 17884 -17997
rect 17850 -18065 17884 -18059
rect 17850 -18093 17884 -18065
rect 17850 -18133 17884 -18131
rect 17850 -18165 17884 -18133
rect 17850 -18235 17884 -18203
rect 17850 -18237 17884 -18235
rect 17850 -18303 17884 -18275
rect 17850 -18309 17884 -18303
rect 17850 -18371 17884 -18347
rect 17850 -18381 17884 -18371
rect 17850 -18439 17884 -18419
rect 17850 -18453 17884 -18439
rect 18868 -17929 18902 -17915
rect 18868 -17949 18902 -17929
rect 18868 -17997 18902 -17987
rect 18868 -18021 18902 -17997
rect 18868 -18065 18902 -18059
rect 18868 -18093 18902 -18065
rect 18868 -18133 18902 -18131
rect 18868 -18165 18902 -18133
rect 18868 -18235 18902 -18203
rect 18868 -18237 18902 -18235
rect 18868 -18303 18902 -18275
rect 18868 -18309 18902 -18303
rect 18868 -18371 18902 -18347
rect 18868 -18381 18902 -18371
rect 18868 -18439 18902 -18419
rect 18868 -18453 18902 -18439
rect 19886 -17929 19920 -17915
rect 19886 -17949 19920 -17929
rect 19886 -17997 19920 -17987
rect 19886 -18021 19920 -17997
rect 19886 -18065 19920 -18059
rect 19886 -18093 19920 -18065
rect 19886 -18133 19920 -18131
rect 19886 -18165 19920 -18133
rect 19886 -18235 19920 -18203
rect 19886 -18237 19920 -18235
rect 19886 -18303 19920 -18275
rect 19886 -18309 19920 -18303
rect 19886 -18371 19920 -18347
rect 19886 -18381 19920 -18371
rect 19886 -18439 19920 -18419
rect 19886 -18453 19920 -18439
rect 20904 -17929 20938 -17915
rect 20904 -17949 20938 -17929
rect 20904 -17997 20938 -17987
rect 20904 -18021 20938 -17997
rect 20904 -18065 20938 -18059
rect 20904 -18093 20938 -18065
rect 20904 -18133 20938 -18131
rect 20904 -18165 20938 -18133
rect 20904 -18235 20938 -18203
rect 20904 -18237 20938 -18235
rect 20904 -18303 20938 -18275
rect 20904 -18309 20938 -18303
rect 20904 -18371 20938 -18347
rect 20904 -18381 20938 -18371
rect 20904 -18439 20938 -18419
rect 20904 -18453 20938 -18439
rect 21922 -17929 21956 -17915
rect 21922 -17949 21956 -17929
rect 21922 -17997 21956 -17987
rect 21922 -18021 21956 -17997
rect 21922 -18065 21956 -18059
rect 21922 -18093 21956 -18065
rect 21922 -18133 21956 -18131
rect 21922 -18165 21956 -18133
rect 21922 -18235 21956 -18203
rect 21922 -18237 21956 -18235
rect 21922 -18303 21956 -18275
rect 21922 -18309 21956 -18303
rect 21922 -18371 21956 -18347
rect 21922 -18381 21956 -18371
rect 21922 -18439 21956 -18419
rect 21922 -18453 21956 -18439
rect 22940 -17929 22974 -17915
rect 22940 -17949 22974 -17929
rect 22940 -17997 22974 -17987
rect 22940 -18021 22974 -17997
rect 22940 -18065 22974 -18059
rect 22940 -18093 22974 -18065
rect 22940 -18133 22974 -18131
rect 22940 -18165 22974 -18133
rect 22940 -18235 22974 -18203
rect 22940 -18237 22974 -18235
rect 22940 -18303 22974 -18275
rect 22940 -18309 22974 -18303
rect 22940 -18371 22974 -18347
rect 22940 -18381 22974 -18371
rect 22940 -18439 22974 -18419
rect 22940 -18453 22974 -18439
rect 24855 -17857 24889 -17851
rect 24855 -17885 24889 -17857
rect 24855 -17925 24889 -17923
rect 24855 -17957 24889 -17925
rect 24855 -18027 24889 -17995
rect 24855 -18029 24889 -18027
rect 24855 -18095 24889 -18067
rect 24855 -18101 24889 -18095
rect 24855 -18163 24889 -18139
rect 24855 -18173 24889 -18163
rect 24855 -18231 24889 -18211
rect 24855 -18245 24889 -18231
rect 24855 -18299 24889 -18283
rect 24855 -18317 24889 -18299
rect 24855 -18367 24889 -18355
rect 24855 -18389 24889 -18367
rect 24855 -18435 24889 -18427
rect 24855 -18461 24889 -18435
rect 2909 -18556 2919 -18522
rect 2919 -18556 2943 -18522
rect 2981 -18556 2987 -18522
rect 2987 -18556 3015 -18522
rect 3053 -18556 3055 -18522
rect 3055 -18556 3087 -18522
rect 3125 -18556 3157 -18522
rect 3157 -18556 3159 -18522
rect 3197 -18556 3225 -18522
rect 3225 -18556 3231 -18522
rect 3269 -18556 3293 -18522
rect 3293 -18556 3303 -18522
rect 3927 -18556 3937 -18522
rect 3937 -18556 3961 -18522
rect 3999 -18556 4005 -18522
rect 4005 -18556 4033 -18522
rect 4071 -18556 4073 -18522
rect 4073 -18556 4105 -18522
rect 4143 -18556 4175 -18522
rect 4175 -18556 4177 -18522
rect 4215 -18556 4243 -18522
rect 4243 -18556 4249 -18522
rect 4287 -18556 4311 -18522
rect 4311 -18556 4321 -18522
rect 4945 -18556 4955 -18522
rect 4955 -18556 4979 -18522
rect 5017 -18556 5023 -18522
rect 5023 -18556 5051 -18522
rect 5089 -18556 5091 -18522
rect 5091 -18556 5123 -18522
rect 5161 -18556 5193 -18522
rect 5193 -18556 5195 -18522
rect 5233 -18556 5261 -18522
rect 5261 -18556 5267 -18522
rect 5305 -18556 5329 -18522
rect 5329 -18556 5339 -18522
rect 5963 -18556 5973 -18522
rect 5973 -18556 5997 -18522
rect 6035 -18556 6041 -18522
rect 6041 -18556 6069 -18522
rect 6107 -18556 6109 -18522
rect 6109 -18556 6141 -18522
rect 6179 -18556 6211 -18522
rect 6211 -18556 6213 -18522
rect 6251 -18556 6279 -18522
rect 6279 -18556 6285 -18522
rect 6323 -18556 6347 -18522
rect 6347 -18556 6357 -18522
rect 6981 -18556 6991 -18522
rect 6991 -18556 7015 -18522
rect 7053 -18556 7059 -18522
rect 7059 -18556 7087 -18522
rect 7125 -18556 7127 -18522
rect 7127 -18556 7159 -18522
rect 7197 -18556 7229 -18522
rect 7229 -18556 7231 -18522
rect 7269 -18556 7297 -18522
rect 7297 -18556 7303 -18522
rect 7341 -18556 7365 -18522
rect 7365 -18556 7375 -18522
rect 7999 -18556 8009 -18522
rect 8009 -18556 8033 -18522
rect 8071 -18556 8077 -18522
rect 8077 -18556 8105 -18522
rect 8143 -18556 8145 -18522
rect 8145 -18556 8177 -18522
rect 8215 -18556 8247 -18522
rect 8247 -18556 8249 -18522
rect 8287 -18556 8315 -18522
rect 8315 -18556 8321 -18522
rect 8359 -18556 8383 -18522
rect 8383 -18556 8393 -18522
rect 9017 -18556 9027 -18522
rect 9027 -18556 9051 -18522
rect 9089 -18556 9095 -18522
rect 9095 -18556 9123 -18522
rect 9161 -18556 9163 -18522
rect 9163 -18556 9195 -18522
rect 9233 -18556 9265 -18522
rect 9265 -18556 9267 -18522
rect 9305 -18556 9333 -18522
rect 9333 -18556 9339 -18522
rect 9377 -18556 9401 -18522
rect 9401 -18556 9411 -18522
rect 10035 -18556 10045 -18522
rect 10045 -18556 10069 -18522
rect 10107 -18556 10113 -18522
rect 10113 -18556 10141 -18522
rect 10179 -18556 10181 -18522
rect 10181 -18556 10213 -18522
rect 10251 -18556 10283 -18522
rect 10283 -18556 10285 -18522
rect 10323 -18556 10351 -18522
rect 10351 -18556 10357 -18522
rect 10395 -18556 10419 -18522
rect 10419 -18556 10429 -18522
rect 11053 -18556 11063 -18522
rect 11063 -18556 11087 -18522
rect 11125 -18556 11131 -18522
rect 11131 -18556 11159 -18522
rect 11197 -18556 11199 -18522
rect 11199 -18556 11231 -18522
rect 11269 -18556 11301 -18522
rect 11301 -18556 11303 -18522
rect 11341 -18556 11369 -18522
rect 11369 -18556 11375 -18522
rect 11413 -18556 11437 -18522
rect 11437 -18556 11447 -18522
rect 12071 -18556 12081 -18522
rect 12081 -18556 12105 -18522
rect 12143 -18556 12149 -18522
rect 12149 -18556 12177 -18522
rect 12215 -18556 12217 -18522
rect 12217 -18556 12249 -18522
rect 12287 -18556 12319 -18522
rect 12319 -18556 12321 -18522
rect 12359 -18556 12387 -18522
rect 12387 -18556 12393 -18522
rect 12431 -18556 12455 -18522
rect 12455 -18556 12465 -18522
rect 13089 -18556 13099 -18522
rect 13099 -18556 13123 -18522
rect 13161 -18556 13167 -18522
rect 13167 -18556 13195 -18522
rect 13233 -18556 13235 -18522
rect 13235 -18556 13267 -18522
rect 13305 -18556 13337 -18522
rect 13337 -18556 13339 -18522
rect 13377 -18556 13405 -18522
rect 13405 -18556 13411 -18522
rect 13449 -18556 13473 -18522
rect 13473 -18556 13483 -18522
rect 14107 -18556 14117 -18522
rect 14117 -18556 14141 -18522
rect 14179 -18556 14185 -18522
rect 14185 -18556 14213 -18522
rect 14251 -18556 14253 -18522
rect 14253 -18556 14285 -18522
rect 14323 -18556 14355 -18522
rect 14355 -18556 14357 -18522
rect 14395 -18556 14423 -18522
rect 14423 -18556 14429 -18522
rect 14467 -18556 14491 -18522
rect 14491 -18556 14501 -18522
rect 15125 -18556 15135 -18522
rect 15135 -18556 15159 -18522
rect 15197 -18556 15203 -18522
rect 15203 -18556 15231 -18522
rect 15269 -18556 15271 -18522
rect 15271 -18556 15303 -18522
rect 15341 -18556 15373 -18522
rect 15373 -18556 15375 -18522
rect 15413 -18556 15441 -18522
rect 15441 -18556 15447 -18522
rect 15485 -18556 15509 -18522
rect 15509 -18556 15519 -18522
rect 16143 -18556 16153 -18522
rect 16153 -18556 16177 -18522
rect 16215 -18556 16221 -18522
rect 16221 -18556 16249 -18522
rect 16287 -18556 16289 -18522
rect 16289 -18556 16321 -18522
rect 16359 -18556 16391 -18522
rect 16391 -18556 16393 -18522
rect 16431 -18556 16459 -18522
rect 16459 -18556 16465 -18522
rect 16503 -18556 16527 -18522
rect 16527 -18556 16537 -18522
rect 17161 -18556 17171 -18522
rect 17171 -18556 17195 -18522
rect 17233 -18556 17239 -18522
rect 17239 -18556 17267 -18522
rect 17305 -18556 17307 -18522
rect 17307 -18556 17339 -18522
rect 17377 -18556 17409 -18522
rect 17409 -18556 17411 -18522
rect 17449 -18556 17477 -18522
rect 17477 -18556 17483 -18522
rect 17521 -18556 17545 -18522
rect 17545 -18556 17555 -18522
rect 18179 -18556 18189 -18522
rect 18189 -18556 18213 -18522
rect 18251 -18556 18257 -18522
rect 18257 -18556 18285 -18522
rect 18323 -18556 18325 -18522
rect 18325 -18556 18357 -18522
rect 18395 -18556 18427 -18522
rect 18427 -18556 18429 -18522
rect 18467 -18556 18495 -18522
rect 18495 -18556 18501 -18522
rect 18539 -18556 18563 -18522
rect 18563 -18556 18573 -18522
rect 19197 -18556 19207 -18522
rect 19207 -18556 19231 -18522
rect 19269 -18556 19275 -18522
rect 19275 -18556 19303 -18522
rect 19341 -18556 19343 -18522
rect 19343 -18556 19375 -18522
rect 19413 -18556 19445 -18522
rect 19445 -18556 19447 -18522
rect 19485 -18556 19513 -18522
rect 19513 -18556 19519 -18522
rect 19557 -18556 19581 -18522
rect 19581 -18556 19591 -18522
rect 20215 -18556 20225 -18522
rect 20225 -18556 20249 -18522
rect 20287 -18556 20293 -18522
rect 20293 -18556 20321 -18522
rect 20359 -18556 20361 -18522
rect 20361 -18556 20393 -18522
rect 20431 -18556 20463 -18522
rect 20463 -18556 20465 -18522
rect 20503 -18556 20531 -18522
rect 20531 -18556 20537 -18522
rect 20575 -18556 20599 -18522
rect 20599 -18556 20609 -18522
rect 21233 -18556 21243 -18522
rect 21243 -18556 21267 -18522
rect 21305 -18556 21311 -18522
rect 21311 -18556 21339 -18522
rect 21377 -18556 21379 -18522
rect 21379 -18556 21411 -18522
rect 21449 -18556 21481 -18522
rect 21481 -18556 21483 -18522
rect 21521 -18556 21549 -18522
rect 21549 -18556 21555 -18522
rect 21593 -18556 21617 -18522
rect 21617 -18556 21627 -18522
rect 22251 -18556 22261 -18522
rect 22261 -18556 22285 -18522
rect 22323 -18556 22329 -18522
rect 22329 -18556 22357 -18522
rect 22395 -18556 22397 -18522
rect 22397 -18556 22429 -18522
rect 22467 -18556 22499 -18522
rect 22499 -18556 22501 -18522
rect 22539 -18556 22567 -18522
rect 22567 -18556 22573 -18522
rect 22611 -18556 22635 -18522
rect 22635 -18556 22645 -18522
rect 24855 -18503 24889 -18499
rect 24855 -18533 24889 -18503
rect -22 -18589 12 -18557
rect -22 -18591 12 -18589
rect -22 -18657 12 -18629
rect -22 -18663 12 -18657
rect -22 -18725 12 -18701
rect -22 -18735 12 -18725
rect -22 -18793 12 -18773
rect -22 -18807 12 -18793
rect 24855 -18605 24889 -18571
rect 24855 -18673 24889 -18643
rect 24855 -18677 24889 -18673
rect 24855 -18741 24889 -18715
rect 24855 -18749 24889 -18741
rect 24855 -18809 24889 -18787
rect 24855 -18821 24889 -18809
rect -12289 -18877 -12255 -18859
rect -12289 -18893 -12255 -18877
rect -8855 -18910 -8845 -18876
rect -8845 -18910 -8821 -18876
rect -8783 -18910 -8777 -18876
rect -8777 -18910 -8749 -18876
rect -8711 -18910 -8709 -18876
rect -8709 -18910 -8677 -18876
rect -8639 -18910 -8607 -18876
rect -8607 -18910 -8605 -18876
rect -8567 -18910 -8539 -18876
rect -8539 -18910 -8533 -18876
rect -8495 -18910 -8471 -18876
rect -8471 -18910 -8461 -18876
rect -7837 -18910 -7827 -18876
rect -7827 -18910 -7803 -18876
rect -7765 -18910 -7759 -18876
rect -7759 -18910 -7731 -18876
rect -7693 -18910 -7691 -18876
rect -7691 -18910 -7659 -18876
rect -7621 -18910 -7589 -18876
rect -7589 -18910 -7587 -18876
rect -7549 -18910 -7521 -18876
rect -7521 -18910 -7515 -18876
rect -7477 -18910 -7453 -18876
rect -7453 -18910 -7443 -18876
rect -6819 -18910 -6809 -18876
rect -6809 -18910 -6785 -18876
rect -6747 -18910 -6741 -18876
rect -6741 -18910 -6713 -18876
rect -6675 -18910 -6673 -18876
rect -6673 -18910 -6641 -18876
rect -6603 -18910 -6571 -18876
rect -6571 -18910 -6569 -18876
rect -6531 -18910 -6503 -18876
rect -6503 -18910 -6497 -18876
rect -6459 -18910 -6435 -18876
rect -6435 -18910 -6425 -18876
rect -5801 -18910 -5791 -18876
rect -5791 -18910 -5767 -18876
rect -5729 -18910 -5723 -18876
rect -5723 -18910 -5695 -18876
rect -5657 -18910 -5655 -18876
rect -5655 -18910 -5623 -18876
rect -5585 -18910 -5553 -18876
rect -5553 -18910 -5551 -18876
rect -5513 -18910 -5485 -18876
rect -5485 -18910 -5479 -18876
rect -5441 -18910 -5417 -18876
rect -5417 -18910 -5407 -18876
rect -4783 -18910 -4773 -18876
rect -4773 -18910 -4749 -18876
rect -4711 -18910 -4705 -18876
rect -4705 -18910 -4677 -18876
rect -4639 -18910 -4637 -18876
rect -4637 -18910 -4605 -18876
rect -4567 -18910 -4535 -18876
rect -4535 -18910 -4533 -18876
rect -4495 -18910 -4467 -18876
rect -4467 -18910 -4461 -18876
rect -4423 -18910 -4399 -18876
rect -4399 -18910 -4389 -18876
rect -3765 -18910 -3755 -18876
rect -3755 -18910 -3731 -18876
rect -3693 -18910 -3687 -18876
rect -3687 -18910 -3659 -18876
rect -3621 -18910 -3619 -18876
rect -3619 -18910 -3587 -18876
rect -3549 -18910 -3517 -18876
rect -3517 -18910 -3515 -18876
rect -3477 -18910 -3449 -18876
rect -3449 -18910 -3443 -18876
rect -3405 -18910 -3381 -18876
rect -3381 -18910 -3371 -18876
rect -2747 -18910 -2737 -18876
rect -2737 -18910 -2713 -18876
rect -2675 -18910 -2669 -18876
rect -2669 -18910 -2641 -18876
rect -2603 -18910 -2601 -18876
rect -2601 -18910 -2569 -18876
rect -2531 -18910 -2499 -18876
rect -2499 -18910 -2497 -18876
rect -2459 -18910 -2431 -18876
rect -2431 -18910 -2425 -18876
rect -2387 -18910 -2363 -18876
rect -2363 -18910 -2353 -18876
rect -1729 -18910 -1719 -18876
rect -1719 -18910 -1695 -18876
rect -1657 -18910 -1651 -18876
rect -1651 -18910 -1623 -18876
rect -1585 -18910 -1583 -18876
rect -1583 -18910 -1551 -18876
rect -1513 -18910 -1481 -18876
rect -1481 -18910 -1479 -18876
rect -1441 -18910 -1413 -18876
rect -1413 -18910 -1407 -18876
rect -1369 -18910 -1345 -18876
rect -1345 -18910 -1335 -18876
rect -711 -18910 -701 -18876
rect -701 -18910 -677 -18876
rect -639 -18910 -633 -18876
rect -633 -18910 -605 -18876
rect -567 -18910 -565 -18876
rect -565 -18910 -533 -18876
rect -495 -18910 -463 -18876
rect -463 -18910 -461 -18876
rect -423 -18910 -395 -18876
rect -395 -18910 -389 -18876
rect -351 -18910 -327 -18876
rect -327 -18910 -317 -18876
rect 24855 -18877 24889 -18859
rect 24855 -18893 24889 -18877
rect -12289 -18945 -12255 -18931
rect -12289 -18965 -12255 -18945
rect -12289 -19013 -12255 -19003
rect -12289 -19037 -12255 -19013
rect 24855 -18945 24889 -18931
rect 24855 -18965 24889 -18945
rect 24855 -19013 24889 -19003
rect 24855 -19037 24889 -19013
rect -12289 -19081 -12255 -19075
rect -12289 -19109 -12255 -19081
rect 2909 -19080 2919 -19046
rect 2919 -19080 2943 -19046
rect 2981 -19080 2987 -19046
rect 2987 -19080 3015 -19046
rect 3053 -19080 3055 -19046
rect 3055 -19080 3087 -19046
rect 3125 -19080 3157 -19046
rect 3157 -19080 3159 -19046
rect 3197 -19080 3225 -19046
rect 3225 -19080 3231 -19046
rect 3269 -19080 3293 -19046
rect 3293 -19080 3303 -19046
rect 3927 -19080 3937 -19046
rect 3937 -19080 3961 -19046
rect 3999 -19080 4005 -19046
rect 4005 -19080 4033 -19046
rect 4071 -19080 4073 -19046
rect 4073 -19080 4105 -19046
rect 4143 -19080 4175 -19046
rect 4175 -19080 4177 -19046
rect 4215 -19080 4243 -19046
rect 4243 -19080 4249 -19046
rect 4287 -19080 4311 -19046
rect 4311 -19080 4321 -19046
rect 4945 -19080 4955 -19046
rect 4955 -19080 4979 -19046
rect 5017 -19080 5023 -19046
rect 5023 -19080 5051 -19046
rect 5089 -19080 5091 -19046
rect 5091 -19080 5123 -19046
rect 5161 -19080 5193 -19046
rect 5193 -19080 5195 -19046
rect 5233 -19080 5261 -19046
rect 5261 -19080 5267 -19046
rect 5305 -19080 5329 -19046
rect 5329 -19080 5339 -19046
rect 5963 -19080 5973 -19046
rect 5973 -19080 5997 -19046
rect 6035 -19080 6041 -19046
rect 6041 -19080 6069 -19046
rect 6107 -19080 6109 -19046
rect 6109 -19080 6141 -19046
rect 6179 -19080 6211 -19046
rect 6211 -19080 6213 -19046
rect 6251 -19080 6279 -19046
rect 6279 -19080 6285 -19046
rect 6323 -19080 6347 -19046
rect 6347 -19080 6357 -19046
rect 6981 -19080 6991 -19046
rect 6991 -19080 7015 -19046
rect 7053 -19080 7059 -19046
rect 7059 -19080 7087 -19046
rect 7125 -19080 7127 -19046
rect 7127 -19080 7159 -19046
rect 7197 -19080 7229 -19046
rect 7229 -19080 7231 -19046
rect 7269 -19080 7297 -19046
rect 7297 -19080 7303 -19046
rect 7341 -19080 7365 -19046
rect 7365 -19080 7375 -19046
rect 7999 -19080 8009 -19046
rect 8009 -19080 8033 -19046
rect 8071 -19080 8077 -19046
rect 8077 -19080 8105 -19046
rect 8143 -19080 8145 -19046
rect 8145 -19080 8177 -19046
rect 8215 -19080 8247 -19046
rect 8247 -19080 8249 -19046
rect 8287 -19080 8315 -19046
rect 8315 -19080 8321 -19046
rect 8359 -19080 8383 -19046
rect 8383 -19080 8393 -19046
rect 9017 -19080 9027 -19046
rect 9027 -19080 9051 -19046
rect 9089 -19080 9095 -19046
rect 9095 -19080 9123 -19046
rect 9161 -19080 9163 -19046
rect 9163 -19080 9195 -19046
rect 9233 -19080 9265 -19046
rect 9265 -19080 9267 -19046
rect 9305 -19080 9333 -19046
rect 9333 -19080 9339 -19046
rect 9377 -19080 9401 -19046
rect 9401 -19080 9411 -19046
rect 10035 -19080 10045 -19046
rect 10045 -19080 10069 -19046
rect 10107 -19080 10113 -19046
rect 10113 -19080 10141 -19046
rect 10179 -19080 10181 -19046
rect 10181 -19080 10213 -19046
rect 10251 -19080 10283 -19046
rect 10283 -19080 10285 -19046
rect 10323 -19080 10351 -19046
rect 10351 -19080 10357 -19046
rect 10395 -19080 10419 -19046
rect 10419 -19080 10429 -19046
rect 11053 -19080 11063 -19046
rect 11063 -19080 11087 -19046
rect 11125 -19080 11131 -19046
rect 11131 -19080 11159 -19046
rect 11197 -19080 11199 -19046
rect 11199 -19080 11231 -19046
rect 11269 -19080 11301 -19046
rect 11301 -19080 11303 -19046
rect 11341 -19080 11369 -19046
rect 11369 -19080 11375 -19046
rect 11413 -19080 11437 -19046
rect 11437 -19080 11447 -19046
rect 12071 -19080 12081 -19046
rect 12081 -19080 12105 -19046
rect 12143 -19080 12149 -19046
rect 12149 -19080 12177 -19046
rect 12215 -19080 12217 -19046
rect 12217 -19080 12249 -19046
rect 12287 -19080 12319 -19046
rect 12319 -19080 12321 -19046
rect 12359 -19080 12387 -19046
rect 12387 -19080 12393 -19046
rect 12431 -19080 12455 -19046
rect 12455 -19080 12465 -19046
rect 13089 -19080 13099 -19046
rect 13099 -19080 13123 -19046
rect 13161 -19080 13167 -19046
rect 13167 -19080 13195 -19046
rect 13233 -19080 13235 -19046
rect 13235 -19080 13267 -19046
rect 13305 -19080 13337 -19046
rect 13337 -19080 13339 -19046
rect 13377 -19080 13405 -19046
rect 13405 -19080 13411 -19046
rect 13449 -19080 13473 -19046
rect 13473 -19080 13483 -19046
rect 14107 -19080 14117 -19046
rect 14117 -19080 14141 -19046
rect 14179 -19080 14185 -19046
rect 14185 -19080 14213 -19046
rect 14251 -19080 14253 -19046
rect 14253 -19080 14285 -19046
rect 14323 -19080 14355 -19046
rect 14355 -19080 14357 -19046
rect 14395 -19080 14423 -19046
rect 14423 -19080 14429 -19046
rect 14467 -19080 14491 -19046
rect 14491 -19080 14501 -19046
rect 15125 -19080 15135 -19046
rect 15135 -19080 15159 -19046
rect 15197 -19080 15203 -19046
rect 15203 -19080 15231 -19046
rect 15269 -19080 15271 -19046
rect 15271 -19080 15303 -19046
rect 15341 -19080 15373 -19046
rect 15373 -19080 15375 -19046
rect 15413 -19080 15441 -19046
rect 15441 -19080 15447 -19046
rect 15485 -19080 15509 -19046
rect 15509 -19080 15519 -19046
rect 16143 -19080 16153 -19046
rect 16153 -19080 16177 -19046
rect 16215 -19080 16221 -19046
rect 16221 -19080 16249 -19046
rect 16287 -19080 16289 -19046
rect 16289 -19080 16321 -19046
rect 16359 -19080 16391 -19046
rect 16391 -19080 16393 -19046
rect 16431 -19080 16459 -19046
rect 16459 -19080 16465 -19046
rect 16503 -19080 16527 -19046
rect 16527 -19080 16537 -19046
rect 17161 -19080 17171 -19046
rect 17171 -19080 17195 -19046
rect 17233 -19080 17239 -19046
rect 17239 -19080 17267 -19046
rect 17305 -19080 17307 -19046
rect 17307 -19080 17339 -19046
rect 17377 -19080 17409 -19046
rect 17409 -19080 17411 -19046
rect 17449 -19080 17477 -19046
rect 17477 -19080 17483 -19046
rect 17521 -19080 17545 -19046
rect 17545 -19080 17555 -19046
rect 18179 -19080 18189 -19046
rect 18189 -19080 18213 -19046
rect 18251 -19080 18257 -19046
rect 18257 -19080 18285 -19046
rect 18323 -19080 18325 -19046
rect 18325 -19080 18357 -19046
rect 18395 -19080 18427 -19046
rect 18427 -19080 18429 -19046
rect 18467 -19080 18495 -19046
rect 18495 -19080 18501 -19046
rect 18539 -19080 18563 -19046
rect 18563 -19080 18573 -19046
rect 19197 -19080 19207 -19046
rect 19207 -19080 19231 -19046
rect 19269 -19080 19275 -19046
rect 19275 -19080 19303 -19046
rect 19341 -19080 19343 -19046
rect 19343 -19080 19375 -19046
rect 19413 -19080 19445 -19046
rect 19445 -19080 19447 -19046
rect 19485 -19080 19513 -19046
rect 19513 -19080 19519 -19046
rect 19557 -19080 19581 -19046
rect 19581 -19080 19591 -19046
rect 20215 -19080 20225 -19046
rect 20225 -19080 20249 -19046
rect 20287 -19080 20293 -19046
rect 20293 -19080 20321 -19046
rect 20359 -19080 20361 -19046
rect 20361 -19080 20393 -19046
rect 20431 -19080 20463 -19046
rect 20463 -19080 20465 -19046
rect 20503 -19080 20531 -19046
rect 20531 -19080 20537 -19046
rect 20575 -19080 20599 -19046
rect 20599 -19080 20609 -19046
rect 21233 -19080 21243 -19046
rect 21243 -19080 21267 -19046
rect 21305 -19080 21311 -19046
rect 21311 -19080 21339 -19046
rect 21377 -19080 21379 -19046
rect 21379 -19080 21411 -19046
rect 21449 -19080 21481 -19046
rect 21481 -19080 21483 -19046
rect 21521 -19080 21549 -19046
rect 21549 -19080 21555 -19046
rect 21593 -19080 21617 -19046
rect 21617 -19080 21627 -19046
rect 22251 -19080 22261 -19046
rect 22261 -19080 22285 -19046
rect 22323 -19080 22329 -19046
rect 22329 -19080 22357 -19046
rect 22395 -19080 22397 -19046
rect 22397 -19080 22429 -19046
rect 22467 -19080 22499 -19046
rect 22499 -19080 22501 -19046
rect 22539 -19080 22567 -19046
rect 22567 -19080 22573 -19046
rect 22611 -19080 22635 -19046
rect 22635 -19080 22645 -19046
rect 24855 -19081 24889 -19075
rect 24855 -19109 24889 -19081
rect -12289 -19149 -12255 -19147
rect -12289 -19181 -12255 -19149
rect -12289 -19251 -12255 -19219
rect -12289 -19253 -12255 -19251
rect -12289 -19319 -12255 -19291
rect -12289 -19325 -12255 -19319
rect -12289 -19387 -12255 -19363
rect -12289 -19397 -12255 -19387
rect -12289 -19455 -12255 -19435
rect -12289 -19469 -12255 -19455
rect -12289 -19523 -12255 -19507
rect -12289 -19541 -12255 -19523
rect 2580 -19163 2614 -19149
rect 2580 -19183 2614 -19163
rect 2580 -19231 2614 -19221
rect 2580 -19255 2614 -19231
rect 2580 -19299 2614 -19293
rect 2580 -19327 2614 -19299
rect 2580 -19367 2614 -19365
rect 2580 -19399 2614 -19367
rect 2580 -19469 2614 -19437
rect 2580 -19471 2614 -19469
rect 2580 -19537 2614 -19509
rect 2580 -19543 2614 -19537
rect -12289 -19591 -12255 -19579
rect -12289 -19613 -12255 -19591
rect -2215 -19584 -2181 -19550
rect -1997 -19584 -1963 -19550
rect -1779 -19584 -1745 -19550
rect -1561 -19584 -1527 -19550
rect -1343 -19584 -1309 -19550
rect -1125 -19584 -1091 -19550
rect -907 -19584 -873 -19550
rect -689 -19584 -655 -19550
rect -471 -19584 -437 -19550
rect -253 -19584 -219 -19550
rect 2580 -19605 2614 -19581
rect 2580 -19615 2614 -19605
rect -12289 -19659 -12255 -19651
rect -12289 -19685 -12255 -19659
rect -12289 -19727 -12255 -19723
rect -12289 -19757 -12255 -19727
rect -12289 -19829 -12255 -19795
rect -2324 -19671 -2290 -19669
rect -2324 -19703 -2290 -19671
rect -2324 -19773 -2290 -19741
rect -2324 -19775 -2290 -19773
rect -2106 -19671 -2072 -19669
rect -2106 -19703 -2072 -19671
rect -2106 -19773 -2072 -19741
rect -2106 -19775 -2072 -19773
rect -1888 -19671 -1854 -19669
rect -1888 -19703 -1854 -19671
rect -1888 -19773 -1854 -19741
rect -1888 -19775 -1854 -19773
rect -1670 -19671 -1636 -19669
rect -1670 -19703 -1636 -19671
rect -1670 -19773 -1636 -19741
rect -1670 -19775 -1636 -19773
rect -1452 -19671 -1418 -19669
rect -1452 -19703 -1418 -19671
rect -1452 -19773 -1418 -19741
rect -1452 -19775 -1418 -19773
rect -1234 -19671 -1200 -19669
rect -1234 -19703 -1200 -19671
rect -1234 -19773 -1200 -19741
rect -1234 -19775 -1200 -19773
rect -1016 -19671 -982 -19669
rect -1016 -19703 -982 -19671
rect -1016 -19773 -982 -19741
rect -1016 -19775 -982 -19773
rect -798 -19671 -764 -19669
rect -798 -19703 -764 -19671
rect -798 -19773 -764 -19741
rect -798 -19775 -764 -19773
rect -580 -19671 -546 -19669
rect -580 -19703 -546 -19671
rect -580 -19773 -546 -19741
rect -580 -19775 -546 -19773
rect -362 -19671 -328 -19669
rect -362 -19703 -328 -19671
rect -362 -19773 -328 -19741
rect -362 -19775 -328 -19773
rect -144 -19671 -110 -19669
rect -144 -19703 -110 -19671
rect 2580 -19673 2614 -19653
rect 2580 -19687 2614 -19673
rect 3598 -19163 3632 -19149
rect 3598 -19183 3632 -19163
rect 3598 -19231 3632 -19221
rect 3598 -19255 3632 -19231
rect 3598 -19299 3632 -19293
rect 3598 -19327 3632 -19299
rect 3598 -19367 3632 -19365
rect 3598 -19399 3632 -19367
rect 3598 -19469 3632 -19437
rect 3598 -19471 3632 -19469
rect 3598 -19537 3632 -19509
rect 3598 -19543 3632 -19537
rect 3598 -19605 3632 -19581
rect 3598 -19615 3632 -19605
rect 3598 -19673 3632 -19653
rect 3598 -19687 3632 -19673
rect 4616 -19163 4650 -19149
rect 4616 -19183 4650 -19163
rect 4616 -19231 4650 -19221
rect 4616 -19255 4650 -19231
rect 4616 -19299 4650 -19293
rect 4616 -19327 4650 -19299
rect 4616 -19367 4650 -19365
rect 4616 -19399 4650 -19367
rect 4616 -19469 4650 -19437
rect 4616 -19471 4650 -19469
rect 4616 -19537 4650 -19509
rect 4616 -19543 4650 -19537
rect 4616 -19605 4650 -19581
rect 4616 -19615 4650 -19605
rect 4616 -19673 4650 -19653
rect 4616 -19687 4650 -19673
rect 5634 -19163 5668 -19149
rect 5634 -19183 5668 -19163
rect 5634 -19231 5668 -19221
rect 5634 -19255 5668 -19231
rect 5634 -19299 5668 -19293
rect 5634 -19327 5668 -19299
rect 5634 -19367 5668 -19365
rect 5634 -19399 5668 -19367
rect 5634 -19469 5668 -19437
rect 5634 -19471 5668 -19469
rect 5634 -19537 5668 -19509
rect 5634 -19543 5668 -19537
rect 5634 -19605 5668 -19581
rect 5634 -19615 5668 -19605
rect 5634 -19673 5668 -19653
rect 5634 -19687 5668 -19673
rect 6652 -19163 6686 -19149
rect 6652 -19183 6686 -19163
rect 6652 -19231 6686 -19221
rect 6652 -19255 6686 -19231
rect 6652 -19299 6686 -19293
rect 6652 -19327 6686 -19299
rect 6652 -19367 6686 -19365
rect 6652 -19399 6686 -19367
rect 6652 -19469 6686 -19437
rect 6652 -19471 6686 -19469
rect 6652 -19537 6686 -19509
rect 6652 -19543 6686 -19537
rect 6652 -19605 6686 -19581
rect 6652 -19615 6686 -19605
rect 6652 -19673 6686 -19653
rect 6652 -19687 6686 -19673
rect 7670 -19163 7704 -19149
rect 7670 -19183 7704 -19163
rect 7670 -19231 7704 -19221
rect 7670 -19255 7704 -19231
rect 7670 -19299 7704 -19293
rect 7670 -19327 7704 -19299
rect 7670 -19367 7704 -19365
rect 7670 -19399 7704 -19367
rect 7670 -19469 7704 -19437
rect 7670 -19471 7704 -19469
rect 7670 -19537 7704 -19509
rect 7670 -19543 7704 -19537
rect 7670 -19605 7704 -19581
rect 7670 -19615 7704 -19605
rect 7670 -19673 7704 -19653
rect 7670 -19687 7704 -19673
rect 8688 -19163 8722 -19149
rect 8688 -19183 8722 -19163
rect 8688 -19231 8722 -19221
rect 8688 -19255 8722 -19231
rect 8688 -19299 8722 -19293
rect 8688 -19327 8722 -19299
rect 8688 -19367 8722 -19365
rect 8688 -19399 8722 -19367
rect 8688 -19469 8722 -19437
rect 8688 -19471 8722 -19469
rect 8688 -19537 8722 -19509
rect 8688 -19543 8722 -19537
rect 8688 -19605 8722 -19581
rect 8688 -19615 8722 -19605
rect 8688 -19673 8722 -19653
rect 8688 -19687 8722 -19673
rect 9706 -19163 9740 -19149
rect 9706 -19183 9740 -19163
rect 9706 -19231 9740 -19221
rect 9706 -19255 9740 -19231
rect 9706 -19299 9740 -19293
rect 9706 -19327 9740 -19299
rect 9706 -19367 9740 -19365
rect 9706 -19399 9740 -19367
rect 9706 -19469 9740 -19437
rect 9706 -19471 9740 -19469
rect 9706 -19537 9740 -19509
rect 9706 -19543 9740 -19537
rect 9706 -19605 9740 -19581
rect 9706 -19615 9740 -19605
rect 9706 -19673 9740 -19653
rect 9706 -19687 9740 -19673
rect 10724 -19163 10758 -19149
rect 10724 -19183 10758 -19163
rect 10724 -19231 10758 -19221
rect 10724 -19255 10758 -19231
rect 10724 -19299 10758 -19293
rect 10724 -19327 10758 -19299
rect 10724 -19367 10758 -19365
rect 10724 -19399 10758 -19367
rect 10724 -19469 10758 -19437
rect 10724 -19471 10758 -19469
rect 10724 -19537 10758 -19509
rect 10724 -19543 10758 -19537
rect 10724 -19605 10758 -19581
rect 10724 -19615 10758 -19605
rect 10724 -19673 10758 -19653
rect 10724 -19687 10758 -19673
rect 11742 -19163 11776 -19149
rect 11742 -19183 11776 -19163
rect 11742 -19231 11776 -19221
rect 11742 -19255 11776 -19231
rect 11742 -19299 11776 -19293
rect 11742 -19327 11776 -19299
rect 11742 -19367 11776 -19365
rect 11742 -19399 11776 -19367
rect 11742 -19469 11776 -19437
rect 11742 -19471 11776 -19469
rect 11742 -19537 11776 -19509
rect 11742 -19543 11776 -19537
rect 11742 -19605 11776 -19581
rect 11742 -19615 11776 -19605
rect 11742 -19673 11776 -19653
rect 11742 -19687 11776 -19673
rect 12760 -19163 12794 -19149
rect 12760 -19183 12794 -19163
rect 12760 -19231 12794 -19221
rect 12760 -19255 12794 -19231
rect 12760 -19299 12794 -19293
rect 12760 -19327 12794 -19299
rect 12760 -19367 12794 -19365
rect 12760 -19399 12794 -19367
rect 12760 -19469 12794 -19437
rect 12760 -19471 12794 -19469
rect 12760 -19537 12794 -19509
rect 12760 -19543 12794 -19537
rect 12760 -19605 12794 -19581
rect 12760 -19615 12794 -19605
rect 12760 -19673 12794 -19653
rect 12760 -19687 12794 -19673
rect 13778 -19163 13812 -19149
rect 13778 -19183 13812 -19163
rect 13778 -19231 13812 -19221
rect 13778 -19255 13812 -19231
rect 13778 -19299 13812 -19293
rect 13778 -19327 13812 -19299
rect 13778 -19367 13812 -19365
rect 13778 -19399 13812 -19367
rect 13778 -19469 13812 -19437
rect 13778 -19471 13812 -19469
rect 13778 -19537 13812 -19509
rect 13778 -19543 13812 -19537
rect 13778 -19605 13812 -19581
rect 13778 -19615 13812 -19605
rect 13778 -19673 13812 -19653
rect 13778 -19687 13812 -19673
rect 14796 -19163 14830 -19149
rect 14796 -19183 14830 -19163
rect 14796 -19231 14830 -19221
rect 14796 -19255 14830 -19231
rect 14796 -19299 14830 -19293
rect 14796 -19327 14830 -19299
rect 14796 -19367 14830 -19365
rect 14796 -19399 14830 -19367
rect 14796 -19469 14830 -19437
rect 14796 -19471 14830 -19469
rect 14796 -19537 14830 -19509
rect 14796 -19543 14830 -19537
rect 14796 -19605 14830 -19581
rect 14796 -19615 14830 -19605
rect 14796 -19673 14830 -19653
rect 14796 -19687 14830 -19673
rect 15814 -19163 15848 -19149
rect 15814 -19183 15848 -19163
rect 15814 -19231 15848 -19221
rect 15814 -19255 15848 -19231
rect 15814 -19299 15848 -19293
rect 15814 -19327 15848 -19299
rect 15814 -19367 15848 -19365
rect 15814 -19399 15848 -19367
rect 15814 -19469 15848 -19437
rect 15814 -19471 15848 -19469
rect 15814 -19537 15848 -19509
rect 15814 -19543 15848 -19537
rect 15814 -19605 15848 -19581
rect 15814 -19615 15848 -19605
rect 15814 -19673 15848 -19653
rect 15814 -19687 15848 -19673
rect 16832 -19163 16866 -19149
rect 16832 -19183 16866 -19163
rect 16832 -19231 16866 -19221
rect 16832 -19255 16866 -19231
rect 16832 -19299 16866 -19293
rect 16832 -19327 16866 -19299
rect 16832 -19367 16866 -19365
rect 16832 -19399 16866 -19367
rect 16832 -19469 16866 -19437
rect 16832 -19471 16866 -19469
rect 16832 -19537 16866 -19509
rect 16832 -19543 16866 -19537
rect 16832 -19605 16866 -19581
rect 16832 -19615 16866 -19605
rect 16832 -19673 16866 -19653
rect 16832 -19687 16866 -19673
rect 17850 -19163 17884 -19149
rect 17850 -19183 17884 -19163
rect 17850 -19231 17884 -19221
rect 17850 -19255 17884 -19231
rect 17850 -19299 17884 -19293
rect 17850 -19327 17884 -19299
rect 17850 -19367 17884 -19365
rect 17850 -19399 17884 -19367
rect 17850 -19469 17884 -19437
rect 17850 -19471 17884 -19469
rect 17850 -19537 17884 -19509
rect 17850 -19543 17884 -19537
rect 17850 -19605 17884 -19581
rect 17850 -19615 17884 -19605
rect 17850 -19673 17884 -19653
rect 17850 -19687 17884 -19673
rect 18868 -19163 18902 -19149
rect 18868 -19183 18902 -19163
rect 18868 -19231 18902 -19221
rect 18868 -19255 18902 -19231
rect 18868 -19299 18902 -19293
rect 18868 -19327 18902 -19299
rect 18868 -19367 18902 -19365
rect 18868 -19399 18902 -19367
rect 18868 -19469 18902 -19437
rect 18868 -19471 18902 -19469
rect 18868 -19537 18902 -19509
rect 18868 -19543 18902 -19537
rect 18868 -19605 18902 -19581
rect 18868 -19615 18902 -19605
rect 18868 -19673 18902 -19653
rect 18868 -19687 18902 -19673
rect 19886 -19163 19920 -19149
rect 19886 -19183 19920 -19163
rect 19886 -19231 19920 -19221
rect 19886 -19255 19920 -19231
rect 19886 -19299 19920 -19293
rect 19886 -19327 19920 -19299
rect 19886 -19367 19920 -19365
rect 19886 -19399 19920 -19367
rect 19886 -19469 19920 -19437
rect 19886 -19471 19920 -19469
rect 19886 -19537 19920 -19509
rect 19886 -19543 19920 -19537
rect 19886 -19605 19920 -19581
rect 19886 -19615 19920 -19605
rect 19886 -19673 19920 -19653
rect 19886 -19687 19920 -19673
rect 20904 -19163 20938 -19149
rect 20904 -19183 20938 -19163
rect 20904 -19231 20938 -19221
rect 20904 -19255 20938 -19231
rect 20904 -19299 20938 -19293
rect 20904 -19327 20938 -19299
rect 20904 -19367 20938 -19365
rect 20904 -19399 20938 -19367
rect 20904 -19469 20938 -19437
rect 20904 -19471 20938 -19469
rect 20904 -19537 20938 -19509
rect 20904 -19543 20938 -19537
rect 20904 -19605 20938 -19581
rect 20904 -19615 20938 -19605
rect 20904 -19673 20938 -19653
rect 20904 -19687 20938 -19673
rect 21922 -19163 21956 -19149
rect 21922 -19183 21956 -19163
rect 21922 -19231 21956 -19221
rect 21922 -19255 21956 -19231
rect 21922 -19299 21956 -19293
rect 21922 -19327 21956 -19299
rect 21922 -19367 21956 -19365
rect 21922 -19399 21956 -19367
rect 21922 -19469 21956 -19437
rect 21922 -19471 21956 -19469
rect 21922 -19537 21956 -19509
rect 21922 -19543 21956 -19537
rect 21922 -19605 21956 -19581
rect 21922 -19615 21956 -19605
rect 21922 -19673 21956 -19653
rect 21922 -19687 21956 -19673
rect 22940 -19163 22974 -19149
rect 22940 -19183 22974 -19163
rect 22940 -19231 22974 -19221
rect 22940 -19255 22974 -19231
rect 22940 -19299 22974 -19293
rect 22940 -19327 22974 -19299
rect 22940 -19367 22974 -19365
rect 22940 -19399 22974 -19367
rect 22940 -19469 22974 -19437
rect 22940 -19471 22974 -19469
rect 22940 -19537 22974 -19509
rect 22940 -19543 22974 -19537
rect 22940 -19605 22974 -19581
rect 22940 -19615 22974 -19605
rect 22940 -19673 22974 -19653
rect 22940 -19687 22974 -19673
rect 24855 -19149 24889 -19147
rect 24855 -19181 24889 -19149
rect 24855 -19251 24889 -19219
rect 24855 -19253 24889 -19251
rect 24855 -19319 24889 -19291
rect 24855 -19325 24889 -19319
rect 24855 -19387 24889 -19363
rect 24855 -19397 24889 -19387
rect 24855 -19455 24889 -19435
rect 24855 -19469 24889 -19455
rect 24855 -19523 24889 -19507
rect 24855 -19541 24889 -19523
rect 24855 -19591 24889 -19579
rect 24855 -19613 24889 -19591
rect 24855 -19659 24889 -19651
rect 24855 -19685 24889 -19659
rect -144 -19773 -110 -19741
rect -144 -19775 -110 -19773
rect 2909 -19790 2919 -19756
rect 2919 -19790 2943 -19756
rect 2981 -19790 2987 -19756
rect 2987 -19790 3015 -19756
rect 3053 -19790 3055 -19756
rect 3055 -19790 3087 -19756
rect 3125 -19790 3157 -19756
rect 3157 -19790 3159 -19756
rect 3197 -19790 3225 -19756
rect 3225 -19790 3231 -19756
rect 3269 -19790 3293 -19756
rect 3293 -19790 3303 -19756
rect 3927 -19790 3937 -19756
rect 3937 -19790 3961 -19756
rect 3999 -19790 4005 -19756
rect 4005 -19790 4033 -19756
rect 4071 -19790 4073 -19756
rect 4073 -19790 4105 -19756
rect 4143 -19790 4175 -19756
rect 4175 -19790 4177 -19756
rect 4215 -19790 4243 -19756
rect 4243 -19790 4249 -19756
rect 4287 -19790 4311 -19756
rect 4311 -19790 4321 -19756
rect 4945 -19790 4955 -19756
rect 4955 -19790 4979 -19756
rect 5017 -19790 5023 -19756
rect 5023 -19790 5051 -19756
rect 5089 -19790 5091 -19756
rect 5091 -19790 5123 -19756
rect 5161 -19790 5193 -19756
rect 5193 -19790 5195 -19756
rect 5233 -19790 5261 -19756
rect 5261 -19790 5267 -19756
rect 5305 -19790 5329 -19756
rect 5329 -19790 5339 -19756
rect 5963 -19790 5973 -19756
rect 5973 -19790 5997 -19756
rect 6035 -19790 6041 -19756
rect 6041 -19790 6069 -19756
rect 6107 -19790 6109 -19756
rect 6109 -19790 6141 -19756
rect 6179 -19790 6211 -19756
rect 6211 -19790 6213 -19756
rect 6251 -19790 6279 -19756
rect 6279 -19790 6285 -19756
rect 6323 -19790 6347 -19756
rect 6347 -19790 6357 -19756
rect 6981 -19790 6991 -19756
rect 6991 -19790 7015 -19756
rect 7053 -19790 7059 -19756
rect 7059 -19790 7087 -19756
rect 7125 -19790 7127 -19756
rect 7127 -19790 7159 -19756
rect 7197 -19790 7229 -19756
rect 7229 -19790 7231 -19756
rect 7269 -19790 7297 -19756
rect 7297 -19790 7303 -19756
rect 7341 -19790 7365 -19756
rect 7365 -19790 7375 -19756
rect 7999 -19790 8009 -19756
rect 8009 -19790 8033 -19756
rect 8071 -19790 8077 -19756
rect 8077 -19790 8105 -19756
rect 8143 -19790 8145 -19756
rect 8145 -19790 8177 -19756
rect 8215 -19790 8247 -19756
rect 8247 -19790 8249 -19756
rect 8287 -19790 8315 -19756
rect 8315 -19790 8321 -19756
rect 8359 -19790 8383 -19756
rect 8383 -19790 8393 -19756
rect 9017 -19790 9027 -19756
rect 9027 -19790 9051 -19756
rect 9089 -19790 9095 -19756
rect 9095 -19790 9123 -19756
rect 9161 -19790 9163 -19756
rect 9163 -19790 9195 -19756
rect 9233 -19790 9265 -19756
rect 9265 -19790 9267 -19756
rect 9305 -19790 9333 -19756
rect 9333 -19790 9339 -19756
rect 9377 -19790 9401 -19756
rect 9401 -19790 9411 -19756
rect 10035 -19790 10045 -19756
rect 10045 -19790 10069 -19756
rect 10107 -19790 10113 -19756
rect 10113 -19790 10141 -19756
rect 10179 -19790 10181 -19756
rect 10181 -19790 10213 -19756
rect 10251 -19790 10283 -19756
rect 10283 -19790 10285 -19756
rect 10323 -19790 10351 -19756
rect 10351 -19790 10357 -19756
rect 10395 -19790 10419 -19756
rect 10419 -19790 10429 -19756
rect 11053 -19790 11063 -19756
rect 11063 -19790 11087 -19756
rect 11125 -19790 11131 -19756
rect 11131 -19790 11159 -19756
rect 11197 -19790 11199 -19756
rect 11199 -19790 11231 -19756
rect 11269 -19790 11301 -19756
rect 11301 -19790 11303 -19756
rect 11341 -19790 11369 -19756
rect 11369 -19790 11375 -19756
rect 11413 -19790 11437 -19756
rect 11437 -19790 11447 -19756
rect 12071 -19790 12081 -19756
rect 12081 -19790 12105 -19756
rect 12143 -19790 12149 -19756
rect 12149 -19790 12177 -19756
rect 12215 -19790 12217 -19756
rect 12217 -19790 12249 -19756
rect 12287 -19790 12319 -19756
rect 12319 -19790 12321 -19756
rect 12359 -19790 12387 -19756
rect 12387 -19790 12393 -19756
rect 12431 -19790 12455 -19756
rect 12455 -19790 12465 -19756
rect 13089 -19790 13099 -19756
rect 13099 -19790 13123 -19756
rect 13161 -19790 13167 -19756
rect 13167 -19790 13195 -19756
rect 13233 -19790 13235 -19756
rect 13235 -19790 13267 -19756
rect 13305 -19790 13337 -19756
rect 13337 -19790 13339 -19756
rect 13377 -19790 13405 -19756
rect 13405 -19790 13411 -19756
rect 13449 -19790 13473 -19756
rect 13473 -19790 13483 -19756
rect 14107 -19790 14117 -19756
rect 14117 -19790 14141 -19756
rect 14179 -19790 14185 -19756
rect 14185 -19790 14213 -19756
rect 14251 -19790 14253 -19756
rect 14253 -19790 14285 -19756
rect 14323 -19790 14355 -19756
rect 14355 -19790 14357 -19756
rect 14395 -19790 14423 -19756
rect 14423 -19790 14429 -19756
rect 14467 -19790 14491 -19756
rect 14491 -19790 14501 -19756
rect 15125 -19790 15135 -19756
rect 15135 -19790 15159 -19756
rect 15197 -19790 15203 -19756
rect 15203 -19790 15231 -19756
rect 15269 -19790 15271 -19756
rect 15271 -19790 15303 -19756
rect 15341 -19790 15373 -19756
rect 15373 -19790 15375 -19756
rect 15413 -19790 15441 -19756
rect 15441 -19790 15447 -19756
rect 15485 -19790 15509 -19756
rect 15509 -19790 15519 -19756
rect 16143 -19790 16153 -19756
rect 16153 -19790 16177 -19756
rect 16215 -19790 16221 -19756
rect 16221 -19790 16249 -19756
rect 16287 -19790 16289 -19756
rect 16289 -19790 16321 -19756
rect 16359 -19790 16391 -19756
rect 16391 -19790 16393 -19756
rect 16431 -19790 16459 -19756
rect 16459 -19790 16465 -19756
rect 16503 -19790 16527 -19756
rect 16527 -19790 16537 -19756
rect 17161 -19790 17171 -19756
rect 17171 -19790 17195 -19756
rect 17233 -19790 17239 -19756
rect 17239 -19790 17267 -19756
rect 17305 -19790 17307 -19756
rect 17307 -19790 17339 -19756
rect 17377 -19790 17409 -19756
rect 17409 -19790 17411 -19756
rect 17449 -19790 17477 -19756
rect 17477 -19790 17483 -19756
rect 17521 -19790 17545 -19756
rect 17545 -19790 17555 -19756
rect 18179 -19790 18189 -19756
rect 18189 -19790 18213 -19756
rect 18251 -19790 18257 -19756
rect 18257 -19790 18285 -19756
rect 18323 -19790 18325 -19756
rect 18325 -19790 18357 -19756
rect 18395 -19790 18427 -19756
rect 18427 -19790 18429 -19756
rect 18467 -19790 18495 -19756
rect 18495 -19790 18501 -19756
rect 18539 -19790 18563 -19756
rect 18563 -19790 18573 -19756
rect 19197 -19790 19207 -19756
rect 19207 -19790 19231 -19756
rect 19269 -19790 19275 -19756
rect 19275 -19790 19303 -19756
rect 19341 -19790 19343 -19756
rect 19343 -19790 19375 -19756
rect 19413 -19790 19445 -19756
rect 19445 -19790 19447 -19756
rect 19485 -19790 19513 -19756
rect 19513 -19790 19519 -19756
rect 19557 -19790 19581 -19756
rect 19581 -19790 19591 -19756
rect 20215 -19790 20225 -19756
rect 20225 -19790 20249 -19756
rect 20287 -19790 20293 -19756
rect 20293 -19790 20321 -19756
rect 20359 -19790 20361 -19756
rect 20361 -19790 20393 -19756
rect 20431 -19790 20463 -19756
rect 20463 -19790 20465 -19756
rect 20503 -19790 20531 -19756
rect 20531 -19790 20537 -19756
rect 20575 -19790 20599 -19756
rect 20599 -19790 20609 -19756
rect 21233 -19790 21243 -19756
rect 21243 -19790 21267 -19756
rect 21305 -19790 21311 -19756
rect 21311 -19790 21339 -19756
rect 21377 -19790 21379 -19756
rect 21379 -19790 21411 -19756
rect 21449 -19790 21481 -19756
rect 21481 -19790 21483 -19756
rect 21521 -19790 21549 -19756
rect 21549 -19790 21555 -19756
rect 21593 -19790 21617 -19756
rect 21617 -19790 21627 -19756
rect 22251 -19790 22261 -19756
rect 22261 -19790 22285 -19756
rect 22323 -19790 22329 -19756
rect 22329 -19790 22357 -19756
rect 22395 -19790 22397 -19756
rect 22397 -19790 22429 -19756
rect 22467 -19790 22499 -19756
rect 22499 -19790 22501 -19756
rect 22539 -19790 22567 -19756
rect 22567 -19790 22573 -19756
rect 22611 -19790 22635 -19756
rect 22635 -19790 22645 -19756
rect 24855 -19727 24889 -19723
rect 24855 -19757 24889 -19727
rect 24855 -19829 24889 -19795
rect -12289 -19897 -12255 -19867
rect -12289 -19901 -12255 -19897
rect -2215 -19894 -2181 -19860
rect -1997 -19894 -1963 -19860
rect -1779 -19894 -1745 -19860
rect -1561 -19894 -1527 -19860
rect -1343 -19894 -1309 -19860
rect -1125 -19894 -1091 -19860
rect -907 -19894 -873 -19860
rect -689 -19894 -655 -19860
rect -471 -19894 -437 -19860
rect -253 -19894 -219 -19860
rect -12289 -19965 -12255 -19939
rect -12289 -19973 -12255 -19965
rect -12289 -20033 -12255 -20011
rect -12289 -20045 -12255 -20033
rect -12289 -20101 -12255 -20083
rect -12289 -20117 -12255 -20101
rect -12289 -20169 -12255 -20155
rect -12289 -20189 -12255 -20169
rect -12289 -20237 -12255 -20227
rect -12289 -20261 -12255 -20237
rect -12289 -20305 -12255 -20299
rect -12289 -20333 -12255 -20305
rect 24855 -19897 24889 -19867
rect 24855 -19901 24889 -19897
rect 24855 -19965 24889 -19939
rect 24855 -19973 24889 -19965
rect 24855 -20033 24889 -20011
rect 24855 -20045 24889 -20033
rect 24855 -20101 24889 -20083
rect 24855 -20117 24889 -20101
rect 24855 -20169 24889 -20155
rect 24855 -20189 24889 -20169
rect 24855 -20237 24889 -20227
rect 24855 -20261 24889 -20237
rect 2909 -20314 2919 -20280
rect 2919 -20314 2943 -20280
rect 2981 -20314 2987 -20280
rect 2987 -20314 3015 -20280
rect 3053 -20314 3055 -20280
rect 3055 -20314 3087 -20280
rect 3125 -20314 3157 -20280
rect 3157 -20314 3159 -20280
rect 3197 -20314 3225 -20280
rect 3225 -20314 3231 -20280
rect 3269 -20314 3293 -20280
rect 3293 -20314 3303 -20280
rect 3927 -20314 3937 -20280
rect 3937 -20314 3961 -20280
rect 3999 -20314 4005 -20280
rect 4005 -20314 4033 -20280
rect 4071 -20314 4073 -20280
rect 4073 -20314 4105 -20280
rect 4143 -20314 4175 -20280
rect 4175 -20314 4177 -20280
rect 4215 -20314 4243 -20280
rect 4243 -20314 4249 -20280
rect 4287 -20314 4311 -20280
rect 4311 -20314 4321 -20280
rect 4945 -20314 4955 -20280
rect 4955 -20314 4979 -20280
rect 5017 -20314 5023 -20280
rect 5023 -20314 5051 -20280
rect 5089 -20314 5091 -20280
rect 5091 -20314 5123 -20280
rect 5161 -20314 5193 -20280
rect 5193 -20314 5195 -20280
rect 5233 -20314 5261 -20280
rect 5261 -20314 5267 -20280
rect 5305 -20314 5329 -20280
rect 5329 -20314 5339 -20280
rect 5963 -20314 5973 -20280
rect 5973 -20314 5997 -20280
rect 6035 -20314 6041 -20280
rect 6041 -20314 6069 -20280
rect 6107 -20314 6109 -20280
rect 6109 -20314 6141 -20280
rect 6179 -20314 6211 -20280
rect 6211 -20314 6213 -20280
rect 6251 -20314 6279 -20280
rect 6279 -20314 6285 -20280
rect 6323 -20314 6347 -20280
rect 6347 -20314 6357 -20280
rect 6981 -20314 6991 -20280
rect 6991 -20314 7015 -20280
rect 7053 -20314 7059 -20280
rect 7059 -20314 7087 -20280
rect 7125 -20314 7127 -20280
rect 7127 -20314 7159 -20280
rect 7197 -20314 7229 -20280
rect 7229 -20314 7231 -20280
rect 7269 -20314 7297 -20280
rect 7297 -20314 7303 -20280
rect 7341 -20314 7365 -20280
rect 7365 -20314 7375 -20280
rect 7999 -20314 8009 -20280
rect 8009 -20314 8033 -20280
rect 8071 -20314 8077 -20280
rect 8077 -20314 8105 -20280
rect 8143 -20314 8145 -20280
rect 8145 -20314 8177 -20280
rect 8215 -20314 8247 -20280
rect 8247 -20314 8249 -20280
rect 8287 -20314 8315 -20280
rect 8315 -20314 8321 -20280
rect 8359 -20314 8383 -20280
rect 8383 -20314 8393 -20280
rect 9017 -20314 9027 -20280
rect 9027 -20314 9051 -20280
rect 9089 -20314 9095 -20280
rect 9095 -20314 9123 -20280
rect 9161 -20314 9163 -20280
rect 9163 -20314 9195 -20280
rect 9233 -20314 9265 -20280
rect 9265 -20314 9267 -20280
rect 9305 -20314 9333 -20280
rect 9333 -20314 9339 -20280
rect 9377 -20314 9401 -20280
rect 9401 -20314 9411 -20280
rect 10035 -20314 10045 -20280
rect 10045 -20314 10069 -20280
rect 10107 -20314 10113 -20280
rect 10113 -20314 10141 -20280
rect 10179 -20314 10181 -20280
rect 10181 -20314 10213 -20280
rect 10251 -20314 10283 -20280
rect 10283 -20314 10285 -20280
rect 10323 -20314 10351 -20280
rect 10351 -20314 10357 -20280
rect 10395 -20314 10419 -20280
rect 10419 -20314 10429 -20280
rect 11053 -20314 11063 -20280
rect 11063 -20314 11087 -20280
rect 11125 -20314 11131 -20280
rect 11131 -20314 11159 -20280
rect 11197 -20314 11199 -20280
rect 11199 -20314 11231 -20280
rect 11269 -20314 11301 -20280
rect 11301 -20314 11303 -20280
rect 11341 -20314 11369 -20280
rect 11369 -20314 11375 -20280
rect 11413 -20314 11437 -20280
rect 11437 -20314 11447 -20280
rect 12071 -20314 12081 -20280
rect 12081 -20314 12105 -20280
rect 12143 -20314 12149 -20280
rect 12149 -20314 12177 -20280
rect 12215 -20314 12217 -20280
rect 12217 -20314 12249 -20280
rect 12287 -20314 12319 -20280
rect 12319 -20314 12321 -20280
rect 12359 -20314 12387 -20280
rect 12387 -20314 12393 -20280
rect 12431 -20314 12455 -20280
rect 12455 -20314 12465 -20280
rect 13089 -20314 13099 -20280
rect 13099 -20314 13123 -20280
rect 13161 -20314 13167 -20280
rect 13167 -20314 13195 -20280
rect 13233 -20314 13235 -20280
rect 13235 -20314 13267 -20280
rect 13305 -20314 13337 -20280
rect 13337 -20314 13339 -20280
rect 13377 -20314 13405 -20280
rect 13405 -20314 13411 -20280
rect 13449 -20314 13473 -20280
rect 13473 -20314 13483 -20280
rect 14107 -20314 14117 -20280
rect 14117 -20314 14141 -20280
rect 14179 -20314 14185 -20280
rect 14185 -20314 14213 -20280
rect 14251 -20314 14253 -20280
rect 14253 -20314 14285 -20280
rect 14323 -20314 14355 -20280
rect 14355 -20314 14357 -20280
rect 14395 -20314 14423 -20280
rect 14423 -20314 14429 -20280
rect 14467 -20314 14491 -20280
rect 14491 -20314 14501 -20280
rect 15125 -20314 15135 -20280
rect 15135 -20314 15159 -20280
rect 15197 -20314 15203 -20280
rect 15203 -20314 15231 -20280
rect 15269 -20314 15271 -20280
rect 15271 -20314 15303 -20280
rect 15341 -20314 15373 -20280
rect 15373 -20314 15375 -20280
rect 15413 -20314 15441 -20280
rect 15441 -20314 15447 -20280
rect 15485 -20314 15509 -20280
rect 15509 -20314 15519 -20280
rect 16143 -20314 16153 -20280
rect 16153 -20314 16177 -20280
rect 16215 -20314 16221 -20280
rect 16221 -20314 16249 -20280
rect 16287 -20314 16289 -20280
rect 16289 -20314 16321 -20280
rect 16359 -20314 16391 -20280
rect 16391 -20314 16393 -20280
rect 16431 -20314 16459 -20280
rect 16459 -20314 16465 -20280
rect 16503 -20314 16527 -20280
rect 16527 -20314 16537 -20280
rect 17161 -20314 17171 -20280
rect 17171 -20314 17195 -20280
rect 17233 -20314 17239 -20280
rect 17239 -20314 17267 -20280
rect 17305 -20314 17307 -20280
rect 17307 -20314 17339 -20280
rect 17377 -20314 17409 -20280
rect 17409 -20314 17411 -20280
rect 17449 -20314 17477 -20280
rect 17477 -20314 17483 -20280
rect 17521 -20314 17545 -20280
rect 17545 -20314 17555 -20280
rect 18179 -20314 18189 -20280
rect 18189 -20314 18213 -20280
rect 18251 -20314 18257 -20280
rect 18257 -20314 18285 -20280
rect 18323 -20314 18325 -20280
rect 18325 -20314 18357 -20280
rect 18395 -20314 18427 -20280
rect 18427 -20314 18429 -20280
rect 18467 -20314 18495 -20280
rect 18495 -20314 18501 -20280
rect 18539 -20314 18563 -20280
rect 18563 -20314 18573 -20280
rect 19197 -20314 19207 -20280
rect 19207 -20314 19231 -20280
rect 19269 -20314 19275 -20280
rect 19275 -20314 19303 -20280
rect 19341 -20314 19343 -20280
rect 19343 -20314 19375 -20280
rect 19413 -20314 19445 -20280
rect 19445 -20314 19447 -20280
rect 19485 -20314 19513 -20280
rect 19513 -20314 19519 -20280
rect 19557 -20314 19581 -20280
rect 19581 -20314 19591 -20280
rect 20215 -20314 20225 -20280
rect 20225 -20314 20249 -20280
rect 20287 -20314 20293 -20280
rect 20293 -20314 20321 -20280
rect 20359 -20314 20361 -20280
rect 20361 -20314 20393 -20280
rect 20431 -20314 20463 -20280
rect 20463 -20314 20465 -20280
rect 20503 -20314 20531 -20280
rect 20531 -20314 20537 -20280
rect 20575 -20314 20599 -20280
rect 20599 -20314 20609 -20280
rect 21233 -20314 21243 -20280
rect 21243 -20314 21267 -20280
rect 21305 -20314 21311 -20280
rect 21311 -20314 21339 -20280
rect 21377 -20314 21379 -20280
rect 21379 -20314 21411 -20280
rect 21449 -20314 21481 -20280
rect 21481 -20314 21483 -20280
rect 21521 -20314 21549 -20280
rect 21549 -20314 21555 -20280
rect 21593 -20314 21617 -20280
rect 21617 -20314 21627 -20280
rect 22251 -20314 22261 -20280
rect 22261 -20314 22285 -20280
rect 22323 -20314 22329 -20280
rect 22329 -20314 22357 -20280
rect 22395 -20314 22397 -20280
rect 22397 -20314 22429 -20280
rect 22467 -20314 22499 -20280
rect 22499 -20314 22501 -20280
rect 22539 -20314 22567 -20280
rect 22567 -20314 22573 -20280
rect 22611 -20314 22635 -20280
rect 22635 -20314 22645 -20280
rect -12289 -20373 -12255 -20371
rect -12289 -20405 -12255 -20373
rect 24855 -20305 24889 -20299
rect 24855 -20333 24889 -20305
rect -2215 -20416 -2181 -20382
rect -1997 -20416 -1963 -20382
rect -1779 -20416 -1745 -20382
rect -1561 -20416 -1527 -20382
rect -1343 -20416 -1309 -20382
rect -1125 -20416 -1091 -20382
rect -907 -20416 -873 -20382
rect -689 -20416 -655 -20382
rect -471 -20416 -437 -20382
rect -253 -20416 -219 -20382
rect 2580 -20397 2614 -20383
rect -12289 -20475 -12255 -20443
rect -12289 -20477 -12255 -20475
rect 2580 -20417 2614 -20397
rect -12289 -20543 -12255 -20515
rect -12289 -20549 -12255 -20543
rect -12289 -20611 -12255 -20587
rect -12289 -20621 -12255 -20611
rect -2324 -20503 -2290 -20501
rect -2324 -20535 -2290 -20503
rect -2324 -20605 -2290 -20573
rect -2324 -20607 -2290 -20605
rect -2106 -20503 -2072 -20501
rect -2106 -20535 -2072 -20503
rect -2106 -20605 -2072 -20573
rect -2106 -20607 -2072 -20605
rect -1888 -20503 -1854 -20501
rect -1888 -20535 -1854 -20503
rect -1888 -20605 -1854 -20573
rect -1888 -20607 -1854 -20605
rect -1670 -20503 -1636 -20501
rect -1670 -20535 -1636 -20503
rect -1670 -20605 -1636 -20573
rect -1670 -20607 -1636 -20605
rect -1452 -20503 -1418 -20501
rect -1452 -20535 -1418 -20503
rect -1452 -20605 -1418 -20573
rect -1452 -20607 -1418 -20605
rect -1234 -20503 -1200 -20501
rect -1234 -20535 -1200 -20503
rect -1234 -20605 -1200 -20573
rect -1234 -20607 -1200 -20605
rect -1016 -20503 -982 -20501
rect -1016 -20535 -982 -20503
rect -1016 -20605 -982 -20573
rect -1016 -20607 -982 -20605
rect -798 -20503 -764 -20501
rect -798 -20535 -764 -20503
rect -798 -20605 -764 -20573
rect -798 -20607 -764 -20605
rect -580 -20503 -546 -20501
rect -580 -20535 -546 -20503
rect -580 -20605 -546 -20573
rect -580 -20607 -546 -20605
rect -362 -20503 -328 -20501
rect -362 -20535 -328 -20503
rect -362 -20605 -328 -20573
rect -362 -20607 -328 -20605
rect -144 -20503 -110 -20501
rect -144 -20535 -110 -20503
rect -144 -20605 -110 -20573
rect -144 -20607 -110 -20605
rect 2580 -20465 2614 -20455
rect 2580 -20489 2614 -20465
rect 2580 -20533 2614 -20527
rect 2580 -20561 2614 -20533
rect 2580 -20601 2614 -20599
rect 2580 -20633 2614 -20601
rect -12289 -20679 -12255 -20659
rect -12289 -20693 -12255 -20679
rect -2215 -20726 -2181 -20692
rect -1997 -20726 -1963 -20692
rect -1779 -20726 -1745 -20692
rect -1561 -20726 -1527 -20692
rect -1343 -20726 -1309 -20692
rect -1125 -20726 -1091 -20692
rect -907 -20726 -873 -20692
rect -689 -20726 -655 -20692
rect -471 -20726 -437 -20692
rect -253 -20726 -219 -20692
rect 2580 -20703 2614 -20671
rect 2580 -20705 2614 -20703
rect -12289 -20747 -12255 -20731
rect -12289 -20765 -12255 -20747
rect -12289 -20815 -12255 -20803
rect -12289 -20837 -12255 -20815
rect -12289 -20883 -12255 -20875
rect -12289 -20909 -12255 -20883
rect -12289 -20951 -12255 -20947
rect -12289 -20981 -12255 -20951
rect 2580 -20771 2614 -20743
rect 2580 -20777 2614 -20771
rect 2580 -20839 2614 -20815
rect 2580 -20849 2614 -20839
rect 2580 -20907 2614 -20887
rect 2580 -20921 2614 -20907
rect 3598 -20397 3632 -20383
rect 3598 -20417 3632 -20397
rect 3598 -20465 3632 -20455
rect 3598 -20489 3632 -20465
rect 3598 -20533 3632 -20527
rect 3598 -20561 3632 -20533
rect 3598 -20601 3632 -20599
rect 3598 -20633 3632 -20601
rect 3598 -20703 3632 -20671
rect 3598 -20705 3632 -20703
rect 3598 -20771 3632 -20743
rect 3598 -20777 3632 -20771
rect 3598 -20839 3632 -20815
rect 3598 -20849 3632 -20839
rect 3598 -20907 3632 -20887
rect 3598 -20921 3632 -20907
rect 4616 -20397 4650 -20383
rect 4616 -20417 4650 -20397
rect 4616 -20465 4650 -20455
rect 4616 -20489 4650 -20465
rect 4616 -20533 4650 -20527
rect 4616 -20561 4650 -20533
rect 4616 -20601 4650 -20599
rect 4616 -20633 4650 -20601
rect 4616 -20703 4650 -20671
rect 4616 -20705 4650 -20703
rect 4616 -20771 4650 -20743
rect 4616 -20777 4650 -20771
rect 4616 -20839 4650 -20815
rect 4616 -20849 4650 -20839
rect 4616 -20907 4650 -20887
rect 4616 -20921 4650 -20907
rect 5634 -20397 5668 -20383
rect 5634 -20417 5668 -20397
rect 5634 -20465 5668 -20455
rect 5634 -20489 5668 -20465
rect 5634 -20533 5668 -20527
rect 5634 -20561 5668 -20533
rect 5634 -20601 5668 -20599
rect 5634 -20633 5668 -20601
rect 5634 -20703 5668 -20671
rect 5634 -20705 5668 -20703
rect 5634 -20771 5668 -20743
rect 5634 -20777 5668 -20771
rect 5634 -20839 5668 -20815
rect 5634 -20849 5668 -20839
rect 5634 -20907 5668 -20887
rect 5634 -20921 5668 -20907
rect 6652 -20397 6686 -20383
rect 6652 -20417 6686 -20397
rect 6652 -20465 6686 -20455
rect 6652 -20489 6686 -20465
rect 6652 -20533 6686 -20527
rect 6652 -20561 6686 -20533
rect 6652 -20601 6686 -20599
rect 6652 -20633 6686 -20601
rect 6652 -20703 6686 -20671
rect 6652 -20705 6686 -20703
rect 6652 -20771 6686 -20743
rect 6652 -20777 6686 -20771
rect 6652 -20839 6686 -20815
rect 6652 -20849 6686 -20839
rect 6652 -20907 6686 -20887
rect 6652 -20921 6686 -20907
rect 7670 -20397 7704 -20383
rect 7670 -20417 7704 -20397
rect 7670 -20465 7704 -20455
rect 7670 -20489 7704 -20465
rect 7670 -20533 7704 -20527
rect 7670 -20561 7704 -20533
rect 7670 -20601 7704 -20599
rect 7670 -20633 7704 -20601
rect 7670 -20703 7704 -20671
rect 7670 -20705 7704 -20703
rect 7670 -20771 7704 -20743
rect 7670 -20777 7704 -20771
rect 7670 -20839 7704 -20815
rect 7670 -20849 7704 -20839
rect 7670 -20907 7704 -20887
rect 7670 -20921 7704 -20907
rect 8688 -20397 8722 -20383
rect 8688 -20417 8722 -20397
rect 8688 -20465 8722 -20455
rect 8688 -20489 8722 -20465
rect 8688 -20533 8722 -20527
rect 8688 -20561 8722 -20533
rect 8688 -20601 8722 -20599
rect 8688 -20633 8722 -20601
rect 8688 -20703 8722 -20671
rect 8688 -20705 8722 -20703
rect 8688 -20771 8722 -20743
rect 8688 -20777 8722 -20771
rect 8688 -20839 8722 -20815
rect 8688 -20849 8722 -20839
rect 8688 -20907 8722 -20887
rect 8688 -20921 8722 -20907
rect 9706 -20397 9740 -20383
rect 9706 -20417 9740 -20397
rect 9706 -20465 9740 -20455
rect 9706 -20489 9740 -20465
rect 9706 -20533 9740 -20527
rect 9706 -20561 9740 -20533
rect 9706 -20601 9740 -20599
rect 9706 -20633 9740 -20601
rect 9706 -20703 9740 -20671
rect 9706 -20705 9740 -20703
rect 9706 -20771 9740 -20743
rect 9706 -20777 9740 -20771
rect 9706 -20839 9740 -20815
rect 9706 -20849 9740 -20839
rect 9706 -20907 9740 -20887
rect 9706 -20921 9740 -20907
rect 10724 -20397 10758 -20383
rect 10724 -20417 10758 -20397
rect 10724 -20465 10758 -20455
rect 10724 -20489 10758 -20465
rect 10724 -20533 10758 -20527
rect 10724 -20561 10758 -20533
rect 10724 -20601 10758 -20599
rect 10724 -20633 10758 -20601
rect 10724 -20703 10758 -20671
rect 10724 -20705 10758 -20703
rect 10724 -20771 10758 -20743
rect 10724 -20777 10758 -20771
rect 10724 -20839 10758 -20815
rect 10724 -20849 10758 -20839
rect 10724 -20907 10758 -20887
rect 10724 -20921 10758 -20907
rect 11742 -20397 11776 -20383
rect 11742 -20417 11776 -20397
rect 11742 -20465 11776 -20455
rect 11742 -20489 11776 -20465
rect 11742 -20533 11776 -20527
rect 11742 -20561 11776 -20533
rect 11742 -20601 11776 -20599
rect 11742 -20633 11776 -20601
rect 11742 -20703 11776 -20671
rect 11742 -20705 11776 -20703
rect 11742 -20771 11776 -20743
rect 11742 -20777 11776 -20771
rect 11742 -20839 11776 -20815
rect 11742 -20849 11776 -20839
rect 11742 -20907 11776 -20887
rect 11742 -20921 11776 -20907
rect 12760 -20397 12794 -20383
rect 12760 -20417 12794 -20397
rect 12760 -20465 12794 -20455
rect 12760 -20489 12794 -20465
rect 12760 -20533 12794 -20527
rect 12760 -20561 12794 -20533
rect 12760 -20601 12794 -20599
rect 12760 -20633 12794 -20601
rect 12760 -20703 12794 -20671
rect 12760 -20705 12794 -20703
rect 12760 -20771 12794 -20743
rect 12760 -20777 12794 -20771
rect 12760 -20839 12794 -20815
rect 12760 -20849 12794 -20839
rect 12760 -20907 12794 -20887
rect 12760 -20921 12794 -20907
rect 13778 -20397 13812 -20383
rect 13778 -20417 13812 -20397
rect 13778 -20465 13812 -20455
rect 13778 -20489 13812 -20465
rect 13778 -20533 13812 -20527
rect 13778 -20561 13812 -20533
rect 13778 -20601 13812 -20599
rect 13778 -20633 13812 -20601
rect 13778 -20703 13812 -20671
rect 13778 -20705 13812 -20703
rect 13778 -20771 13812 -20743
rect 13778 -20777 13812 -20771
rect 13778 -20839 13812 -20815
rect 13778 -20849 13812 -20839
rect 13778 -20907 13812 -20887
rect 13778 -20921 13812 -20907
rect 14796 -20397 14830 -20383
rect 14796 -20417 14830 -20397
rect 14796 -20465 14830 -20455
rect 14796 -20489 14830 -20465
rect 14796 -20533 14830 -20527
rect 14796 -20561 14830 -20533
rect 14796 -20601 14830 -20599
rect 14796 -20633 14830 -20601
rect 14796 -20703 14830 -20671
rect 14796 -20705 14830 -20703
rect 14796 -20771 14830 -20743
rect 14796 -20777 14830 -20771
rect 14796 -20839 14830 -20815
rect 14796 -20849 14830 -20839
rect 14796 -20907 14830 -20887
rect 14796 -20921 14830 -20907
rect 15814 -20397 15848 -20383
rect 15814 -20417 15848 -20397
rect 15814 -20465 15848 -20455
rect 15814 -20489 15848 -20465
rect 15814 -20533 15848 -20527
rect 15814 -20561 15848 -20533
rect 15814 -20601 15848 -20599
rect 15814 -20633 15848 -20601
rect 15814 -20703 15848 -20671
rect 15814 -20705 15848 -20703
rect 15814 -20771 15848 -20743
rect 15814 -20777 15848 -20771
rect 15814 -20839 15848 -20815
rect 15814 -20849 15848 -20839
rect 15814 -20907 15848 -20887
rect 15814 -20921 15848 -20907
rect 16832 -20397 16866 -20383
rect 16832 -20417 16866 -20397
rect 16832 -20465 16866 -20455
rect 16832 -20489 16866 -20465
rect 16832 -20533 16866 -20527
rect 16832 -20561 16866 -20533
rect 16832 -20601 16866 -20599
rect 16832 -20633 16866 -20601
rect 16832 -20703 16866 -20671
rect 16832 -20705 16866 -20703
rect 16832 -20771 16866 -20743
rect 16832 -20777 16866 -20771
rect 16832 -20839 16866 -20815
rect 16832 -20849 16866 -20839
rect 16832 -20907 16866 -20887
rect 16832 -20921 16866 -20907
rect 17850 -20397 17884 -20383
rect 17850 -20417 17884 -20397
rect 17850 -20465 17884 -20455
rect 17850 -20489 17884 -20465
rect 17850 -20533 17884 -20527
rect 17850 -20561 17884 -20533
rect 17850 -20601 17884 -20599
rect 17850 -20633 17884 -20601
rect 17850 -20703 17884 -20671
rect 17850 -20705 17884 -20703
rect 17850 -20771 17884 -20743
rect 17850 -20777 17884 -20771
rect 17850 -20839 17884 -20815
rect 17850 -20849 17884 -20839
rect 17850 -20907 17884 -20887
rect 17850 -20921 17884 -20907
rect 18868 -20397 18902 -20383
rect 18868 -20417 18902 -20397
rect 18868 -20465 18902 -20455
rect 18868 -20489 18902 -20465
rect 18868 -20533 18902 -20527
rect 18868 -20561 18902 -20533
rect 18868 -20601 18902 -20599
rect 18868 -20633 18902 -20601
rect 18868 -20703 18902 -20671
rect 18868 -20705 18902 -20703
rect 18868 -20771 18902 -20743
rect 18868 -20777 18902 -20771
rect 18868 -20839 18902 -20815
rect 18868 -20849 18902 -20839
rect 18868 -20907 18902 -20887
rect 18868 -20921 18902 -20907
rect 19886 -20397 19920 -20383
rect 19886 -20417 19920 -20397
rect 19886 -20465 19920 -20455
rect 19886 -20489 19920 -20465
rect 19886 -20533 19920 -20527
rect 19886 -20561 19920 -20533
rect 19886 -20601 19920 -20599
rect 19886 -20633 19920 -20601
rect 19886 -20703 19920 -20671
rect 19886 -20705 19920 -20703
rect 19886 -20771 19920 -20743
rect 19886 -20777 19920 -20771
rect 19886 -20839 19920 -20815
rect 19886 -20849 19920 -20839
rect 19886 -20907 19920 -20887
rect 19886 -20921 19920 -20907
rect 20904 -20397 20938 -20383
rect 20904 -20417 20938 -20397
rect 20904 -20465 20938 -20455
rect 20904 -20489 20938 -20465
rect 20904 -20533 20938 -20527
rect 20904 -20561 20938 -20533
rect 20904 -20601 20938 -20599
rect 20904 -20633 20938 -20601
rect 20904 -20703 20938 -20671
rect 20904 -20705 20938 -20703
rect 20904 -20771 20938 -20743
rect 20904 -20777 20938 -20771
rect 20904 -20839 20938 -20815
rect 20904 -20849 20938 -20839
rect 20904 -20907 20938 -20887
rect 20904 -20921 20938 -20907
rect 21922 -20397 21956 -20383
rect 21922 -20417 21956 -20397
rect 21922 -20465 21956 -20455
rect 21922 -20489 21956 -20465
rect 21922 -20533 21956 -20527
rect 21922 -20561 21956 -20533
rect 21922 -20601 21956 -20599
rect 21922 -20633 21956 -20601
rect 21922 -20703 21956 -20671
rect 21922 -20705 21956 -20703
rect 21922 -20771 21956 -20743
rect 21922 -20777 21956 -20771
rect 21922 -20839 21956 -20815
rect 21922 -20849 21956 -20839
rect 21922 -20907 21956 -20887
rect 21922 -20921 21956 -20907
rect 22940 -20397 22974 -20383
rect 22940 -20417 22974 -20397
rect 22940 -20465 22974 -20455
rect 22940 -20489 22974 -20465
rect 22940 -20533 22974 -20527
rect 22940 -20561 22974 -20533
rect 22940 -20601 22974 -20599
rect 22940 -20633 22974 -20601
rect 22940 -20703 22974 -20671
rect 22940 -20705 22974 -20703
rect 22940 -20771 22974 -20743
rect 22940 -20777 22974 -20771
rect 22940 -20839 22974 -20815
rect 22940 -20849 22974 -20839
rect 22940 -20907 22974 -20887
rect 22940 -20921 22974 -20907
rect 24855 -20373 24889 -20371
rect 24855 -20405 24889 -20373
rect 24855 -20475 24889 -20443
rect 24855 -20477 24889 -20475
rect 24855 -20543 24889 -20515
rect 24855 -20549 24889 -20543
rect 24855 -20611 24889 -20587
rect 24855 -20621 24889 -20611
rect 24855 -20679 24889 -20659
rect 24855 -20693 24889 -20679
rect 24855 -20747 24889 -20731
rect 24855 -20765 24889 -20747
rect 24855 -20815 24889 -20803
rect 24855 -20837 24889 -20815
rect 24855 -20883 24889 -20875
rect 24855 -20909 24889 -20883
rect 24855 -20951 24889 -20947
rect 24855 -20981 24889 -20951
rect -12289 -21053 -12255 -21019
rect 2909 -21024 2919 -20990
rect 2919 -21024 2943 -20990
rect 2981 -21024 2987 -20990
rect 2987 -21024 3015 -20990
rect 3053 -21024 3055 -20990
rect 3055 -21024 3087 -20990
rect 3125 -21024 3157 -20990
rect 3157 -21024 3159 -20990
rect 3197 -21024 3225 -20990
rect 3225 -21024 3231 -20990
rect 3269 -21024 3293 -20990
rect 3293 -21024 3303 -20990
rect 3927 -21024 3937 -20990
rect 3937 -21024 3961 -20990
rect 3999 -21024 4005 -20990
rect 4005 -21024 4033 -20990
rect 4071 -21024 4073 -20990
rect 4073 -21024 4105 -20990
rect 4143 -21024 4175 -20990
rect 4175 -21024 4177 -20990
rect 4215 -21024 4243 -20990
rect 4243 -21024 4249 -20990
rect 4287 -21024 4311 -20990
rect 4311 -21024 4321 -20990
rect 4945 -21024 4955 -20990
rect 4955 -21024 4979 -20990
rect 5017 -21024 5023 -20990
rect 5023 -21024 5051 -20990
rect 5089 -21024 5091 -20990
rect 5091 -21024 5123 -20990
rect 5161 -21024 5193 -20990
rect 5193 -21024 5195 -20990
rect 5233 -21024 5261 -20990
rect 5261 -21024 5267 -20990
rect 5305 -21024 5329 -20990
rect 5329 -21024 5339 -20990
rect 5963 -21024 5973 -20990
rect 5973 -21024 5997 -20990
rect 6035 -21024 6041 -20990
rect 6041 -21024 6069 -20990
rect 6107 -21024 6109 -20990
rect 6109 -21024 6141 -20990
rect 6179 -21024 6211 -20990
rect 6211 -21024 6213 -20990
rect 6251 -21024 6279 -20990
rect 6279 -21024 6285 -20990
rect 6323 -21024 6347 -20990
rect 6347 -21024 6357 -20990
rect 6981 -21024 6991 -20990
rect 6991 -21024 7015 -20990
rect 7053 -21024 7059 -20990
rect 7059 -21024 7087 -20990
rect 7125 -21024 7127 -20990
rect 7127 -21024 7159 -20990
rect 7197 -21024 7229 -20990
rect 7229 -21024 7231 -20990
rect 7269 -21024 7297 -20990
rect 7297 -21024 7303 -20990
rect 7341 -21024 7365 -20990
rect 7365 -21024 7375 -20990
rect 7999 -21024 8009 -20990
rect 8009 -21024 8033 -20990
rect 8071 -21024 8077 -20990
rect 8077 -21024 8105 -20990
rect 8143 -21024 8145 -20990
rect 8145 -21024 8177 -20990
rect 8215 -21024 8247 -20990
rect 8247 -21024 8249 -20990
rect 8287 -21024 8315 -20990
rect 8315 -21024 8321 -20990
rect 8359 -21024 8383 -20990
rect 8383 -21024 8393 -20990
rect 9017 -21024 9027 -20990
rect 9027 -21024 9051 -20990
rect 9089 -21024 9095 -20990
rect 9095 -21024 9123 -20990
rect 9161 -21024 9163 -20990
rect 9163 -21024 9195 -20990
rect 9233 -21024 9265 -20990
rect 9265 -21024 9267 -20990
rect 9305 -21024 9333 -20990
rect 9333 -21024 9339 -20990
rect 9377 -21024 9401 -20990
rect 9401 -21024 9411 -20990
rect 10035 -21024 10045 -20990
rect 10045 -21024 10069 -20990
rect 10107 -21024 10113 -20990
rect 10113 -21024 10141 -20990
rect 10179 -21024 10181 -20990
rect 10181 -21024 10213 -20990
rect 10251 -21024 10283 -20990
rect 10283 -21024 10285 -20990
rect 10323 -21024 10351 -20990
rect 10351 -21024 10357 -20990
rect 10395 -21024 10419 -20990
rect 10419 -21024 10429 -20990
rect 11053 -21024 11063 -20990
rect 11063 -21024 11087 -20990
rect 11125 -21024 11131 -20990
rect 11131 -21024 11159 -20990
rect 11197 -21024 11199 -20990
rect 11199 -21024 11231 -20990
rect 11269 -21024 11301 -20990
rect 11301 -21024 11303 -20990
rect 11341 -21024 11369 -20990
rect 11369 -21024 11375 -20990
rect 11413 -21024 11437 -20990
rect 11437 -21024 11447 -20990
rect 12071 -21024 12081 -20990
rect 12081 -21024 12105 -20990
rect 12143 -21024 12149 -20990
rect 12149 -21024 12177 -20990
rect 12215 -21024 12217 -20990
rect 12217 -21024 12249 -20990
rect 12287 -21024 12319 -20990
rect 12319 -21024 12321 -20990
rect 12359 -21024 12387 -20990
rect 12387 -21024 12393 -20990
rect 12431 -21024 12455 -20990
rect 12455 -21024 12465 -20990
rect 13089 -21024 13099 -20990
rect 13099 -21024 13123 -20990
rect 13161 -21024 13167 -20990
rect 13167 -21024 13195 -20990
rect 13233 -21024 13235 -20990
rect 13235 -21024 13267 -20990
rect 13305 -21024 13337 -20990
rect 13337 -21024 13339 -20990
rect 13377 -21024 13405 -20990
rect 13405 -21024 13411 -20990
rect 13449 -21024 13473 -20990
rect 13473 -21024 13483 -20990
rect 14107 -21024 14117 -20990
rect 14117 -21024 14141 -20990
rect 14179 -21024 14185 -20990
rect 14185 -21024 14213 -20990
rect 14251 -21024 14253 -20990
rect 14253 -21024 14285 -20990
rect 14323 -21024 14355 -20990
rect 14355 -21024 14357 -20990
rect 14395 -21024 14423 -20990
rect 14423 -21024 14429 -20990
rect 14467 -21024 14491 -20990
rect 14491 -21024 14501 -20990
rect 15125 -21024 15135 -20990
rect 15135 -21024 15159 -20990
rect 15197 -21024 15203 -20990
rect 15203 -21024 15231 -20990
rect 15269 -21024 15271 -20990
rect 15271 -21024 15303 -20990
rect 15341 -21024 15373 -20990
rect 15373 -21024 15375 -20990
rect 15413 -21024 15441 -20990
rect 15441 -21024 15447 -20990
rect 15485 -21024 15509 -20990
rect 15509 -21024 15519 -20990
rect 16143 -21024 16153 -20990
rect 16153 -21024 16177 -20990
rect 16215 -21024 16221 -20990
rect 16221 -21024 16249 -20990
rect 16287 -21024 16289 -20990
rect 16289 -21024 16321 -20990
rect 16359 -21024 16391 -20990
rect 16391 -21024 16393 -20990
rect 16431 -21024 16459 -20990
rect 16459 -21024 16465 -20990
rect 16503 -21024 16527 -20990
rect 16527 -21024 16537 -20990
rect 17161 -21024 17171 -20990
rect 17171 -21024 17195 -20990
rect 17233 -21024 17239 -20990
rect 17239 -21024 17267 -20990
rect 17305 -21024 17307 -20990
rect 17307 -21024 17339 -20990
rect 17377 -21024 17409 -20990
rect 17409 -21024 17411 -20990
rect 17449 -21024 17477 -20990
rect 17477 -21024 17483 -20990
rect 17521 -21024 17545 -20990
rect 17545 -21024 17555 -20990
rect 18179 -21024 18189 -20990
rect 18189 -21024 18213 -20990
rect 18251 -21024 18257 -20990
rect 18257 -21024 18285 -20990
rect 18323 -21024 18325 -20990
rect 18325 -21024 18357 -20990
rect 18395 -21024 18427 -20990
rect 18427 -21024 18429 -20990
rect 18467 -21024 18495 -20990
rect 18495 -21024 18501 -20990
rect 18539 -21024 18563 -20990
rect 18563 -21024 18573 -20990
rect 19197 -21024 19207 -20990
rect 19207 -21024 19231 -20990
rect 19269 -21024 19275 -20990
rect 19275 -21024 19303 -20990
rect 19341 -21024 19343 -20990
rect 19343 -21024 19375 -20990
rect 19413 -21024 19445 -20990
rect 19445 -21024 19447 -20990
rect 19485 -21024 19513 -20990
rect 19513 -21024 19519 -20990
rect 19557 -21024 19581 -20990
rect 19581 -21024 19591 -20990
rect 20215 -21024 20225 -20990
rect 20225 -21024 20249 -20990
rect 20287 -21024 20293 -20990
rect 20293 -21024 20321 -20990
rect 20359 -21024 20361 -20990
rect 20361 -21024 20393 -20990
rect 20431 -21024 20463 -20990
rect 20463 -21024 20465 -20990
rect 20503 -21024 20531 -20990
rect 20531 -21024 20537 -20990
rect 20575 -21024 20599 -20990
rect 20599 -21024 20609 -20990
rect 21233 -21024 21243 -20990
rect 21243 -21024 21267 -20990
rect 21305 -21024 21311 -20990
rect 21311 -21024 21339 -20990
rect 21377 -21024 21379 -20990
rect 21379 -21024 21411 -20990
rect 21449 -21024 21481 -20990
rect 21481 -21024 21483 -20990
rect 21521 -21024 21549 -20990
rect 21549 -21024 21555 -20990
rect 21593 -21024 21617 -20990
rect 21617 -21024 21627 -20990
rect 22251 -21024 22261 -20990
rect 22261 -21024 22285 -20990
rect 22323 -21024 22329 -20990
rect 22329 -21024 22357 -20990
rect 22395 -21024 22397 -20990
rect 22397 -21024 22429 -20990
rect 22467 -21024 22499 -20990
rect 22499 -21024 22501 -20990
rect 22539 -21024 22567 -20990
rect 22567 -21024 22573 -20990
rect 22611 -21024 22635 -20990
rect 22635 -21024 22645 -20990
rect -12289 -21121 -12255 -21091
rect -12289 -21125 -12255 -21121
rect -12289 -21189 -12255 -21163
rect -12289 -21197 -12255 -21189
rect -12289 -21257 -12255 -21235
rect -12289 -21269 -12255 -21257
rect -12289 -21325 -12255 -21307
rect -12289 -21341 -12255 -21325
rect -12289 -21393 -12255 -21379
rect -12289 -21413 -12255 -21393
rect -12289 -21461 -12255 -21451
rect -12289 -21485 -12255 -21461
rect -12289 -21529 -12255 -21523
rect -12289 -21557 -12255 -21529
rect 24855 -21053 24889 -21019
rect 24855 -21121 24889 -21091
rect 24855 -21125 24889 -21121
rect 24855 -21189 24889 -21163
rect 24855 -21197 24889 -21189
rect 24855 -21257 24889 -21235
rect 24855 -21269 24889 -21257
rect 24855 -21325 24889 -21307
rect 24855 -21341 24889 -21325
rect 24855 -21393 24889 -21379
rect 24855 -21413 24889 -21393
rect 24855 -21461 24889 -21451
rect 24855 -21485 24889 -21461
rect 2909 -21546 2919 -21512
rect 2919 -21546 2943 -21512
rect 2981 -21546 2987 -21512
rect 2987 -21546 3015 -21512
rect 3053 -21546 3055 -21512
rect 3055 -21546 3087 -21512
rect 3125 -21546 3157 -21512
rect 3157 -21546 3159 -21512
rect 3197 -21546 3225 -21512
rect 3225 -21546 3231 -21512
rect 3269 -21546 3293 -21512
rect 3293 -21546 3303 -21512
rect 3927 -21546 3937 -21512
rect 3937 -21546 3961 -21512
rect 3999 -21546 4005 -21512
rect 4005 -21546 4033 -21512
rect 4071 -21546 4073 -21512
rect 4073 -21546 4105 -21512
rect 4143 -21546 4175 -21512
rect 4175 -21546 4177 -21512
rect 4215 -21546 4243 -21512
rect 4243 -21546 4249 -21512
rect 4287 -21546 4311 -21512
rect 4311 -21546 4321 -21512
rect 4945 -21546 4955 -21512
rect 4955 -21546 4979 -21512
rect 5017 -21546 5023 -21512
rect 5023 -21546 5051 -21512
rect 5089 -21546 5091 -21512
rect 5091 -21546 5123 -21512
rect 5161 -21546 5193 -21512
rect 5193 -21546 5195 -21512
rect 5233 -21546 5261 -21512
rect 5261 -21546 5267 -21512
rect 5305 -21546 5329 -21512
rect 5329 -21546 5339 -21512
rect 5963 -21546 5973 -21512
rect 5973 -21546 5997 -21512
rect 6035 -21546 6041 -21512
rect 6041 -21546 6069 -21512
rect 6107 -21546 6109 -21512
rect 6109 -21546 6141 -21512
rect 6179 -21546 6211 -21512
rect 6211 -21546 6213 -21512
rect 6251 -21546 6279 -21512
rect 6279 -21546 6285 -21512
rect 6323 -21546 6347 -21512
rect 6347 -21546 6357 -21512
rect 6981 -21546 6991 -21512
rect 6991 -21546 7015 -21512
rect 7053 -21546 7059 -21512
rect 7059 -21546 7087 -21512
rect 7125 -21546 7127 -21512
rect 7127 -21546 7159 -21512
rect 7197 -21546 7229 -21512
rect 7229 -21546 7231 -21512
rect 7269 -21546 7297 -21512
rect 7297 -21546 7303 -21512
rect 7341 -21546 7365 -21512
rect 7365 -21546 7375 -21512
rect 7999 -21546 8009 -21512
rect 8009 -21546 8033 -21512
rect 8071 -21546 8077 -21512
rect 8077 -21546 8105 -21512
rect 8143 -21546 8145 -21512
rect 8145 -21546 8177 -21512
rect 8215 -21546 8247 -21512
rect 8247 -21546 8249 -21512
rect 8287 -21546 8315 -21512
rect 8315 -21546 8321 -21512
rect 8359 -21546 8383 -21512
rect 8383 -21546 8393 -21512
rect 9017 -21546 9027 -21512
rect 9027 -21546 9051 -21512
rect 9089 -21546 9095 -21512
rect 9095 -21546 9123 -21512
rect 9161 -21546 9163 -21512
rect 9163 -21546 9195 -21512
rect 9233 -21546 9265 -21512
rect 9265 -21546 9267 -21512
rect 9305 -21546 9333 -21512
rect 9333 -21546 9339 -21512
rect 9377 -21546 9401 -21512
rect 9401 -21546 9411 -21512
rect 10035 -21546 10045 -21512
rect 10045 -21546 10069 -21512
rect 10107 -21546 10113 -21512
rect 10113 -21546 10141 -21512
rect 10179 -21546 10181 -21512
rect 10181 -21546 10213 -21512
rect 10251 -21546 10283 -21512
rect 10283 -21546 10285 -21512
rect 10323 -21546 10351 -21512
rect 10351 -21546 10357 -21512
rect 10395 -21546 10419 -21512
rect 10419 -21546 10429 -21512
rect 11053 -21546 11063 -21512
rect 11063 -21546 11087 -21512
rect 11125 -21546 11131 -21512
rect 11131 -21546 11159 -21512
rect 11197 -21546 11199 -21512
rect 11199 -21546 11231 -21512
rect 11269 -21546 11301 -21512
rect 11301 -21546 11303 -21512
rect 11341 -21546 11369 -21512
rect 11369 -21546 11375 -21512
rect 11413 -21546 11437 -21512
rect 11437 -21546 11447 -21512
rect 12071 -21546 12081 -21512
rect 12081 -21546 12105 -21512
rect 12143 -21546 12149 -21512
rect 12149 -21546 12177 -21512
rect 12215 -21546 12217 -21512
rect 12217 -21546 12249 -21512
rect 12287 -21546 12319 -21512
rect 12319 -21546 12321 -21512
rect 12359 -21546 12387 -21512
rect 12387 -21546 12393 -21512
rect 12431 -21546 12455 -21512
rect 12455 -21546 12465 -21512
rect 13089 -21546 13099 -21512
rect 13099 -21546 13123 -21512
rect 13161 -21546 13167 -21512
rect 13167 -21546 13195 -21512
rect 13233 -21546 13235 -21512
rect 13235 -21546 13267 -21512
rect 13305 -21546 13337 -21512
rect 13337 -21546 13339 -21512
rect 13377 -21546 13405 -21512
rect 13405 -21546 13411 -21512
rect 13449 -21546 13473 -21512
rect 13473 -21546 13483 -21512
rect 14107 -21546 14117 -21512
rect 14117 -21546 14141 -21512
rect 14179 -21546 14185 -21512
rect 14185 -21546 14213 -21512
rect 14251 -21546 14253 -21512
rect 14253 -21546 14285 -21512
rect 14323 -21546 14355 -21512
rect 14355 -21546 14357 -21512
rect 14395 -21546 14423 -21512
rect 14423 -21546 14429 -21512
rect 14467 -21546 14491 -21512
rect 14491 -21546 14501 -21512
rect 15125 -21546 15135 -21512
rect 15135 -21546 15159 -21512
rect 15197 -21546 15203 -21512
rect 15203 -21546 15231 -21512
rect 15269 -21546 15271 -21512
rect 15271 -21546 15303 -21512
rect 15341 -21546 15373 -21512
rect 15373 -21546 15375 -21512
rect 15413 -21546 15441 -21512
rect 15441 -21546 15447 -21512
rect 15485 -21546 15509 -21512
rect 15509 -21546 15519 -21512
rect 16143 -21546 16153 -21512
rect 16153 -21546 16177 -21512
rect 16215 -21546 16221 -21512
rect 16221 -21546 16249 -21512
rect 16287 -21546 16289 -21512
rect 16289 -21546 16321 -21512
rect 16359 -21546 16391 -21512
rect 16391 -21546 16393 -21512
rect 16431 -21546 16459 -21512
rect 16459 -21546 16465 -21512
rect 16503 -21546 16527 -21512
rect 16527 -21546 16537 -21512
rect 17161 -21546 17171 -21512
rect 17171 -21546 17195 -21512
rect 17233 -21546 17239 -21512
rect 17239 -21546 17267 -21512
rect 17305 -21546 17307 -21512
rect 17307 -21546 17339 -21512
rect 17377 -21546 17409 -21512
rect 17409 -21546 17411 -21512
rect 17449 -21546 17477 -21512
rect 17477 -21546 17483 -21512
rect 17521 -21546 17545 -21512
rect 17545 -21546 17555 -21512
rect 18179 -21546 18189 -21512
rect 18189 -21546 18213 -21512
rect 18251 -21546 18257 -21512
rect 18257 -21546 18285 -21512
rect 18323 -21546 18325 -21512
rect 18325 -21546 18357 -21512
rect 18395 -21546 18427 -21512
rect 18427 -21546 18429 -21512
rect 18467 -21546 18495 -21512
rect 18495 -21546 18501 -21512
rect 18539 -21546 18563 -21512
rect 18563 -21546 18573 -21512
rect 19197 -21546 19207 -21512
rect 19207 -21546 19231 -21512
rect 19269 -21546 19275 -21512
rect 19275 -21546 19303 -21512
rect 19341 -21546 19343 -21512
rect 19343 -21546 19375 -21512
rect 19413 -21546 19445 -21512
rect 19445 -21546 19447 -21512
rect 19485 -21546 19513 -21512
rect 19513 -21546 19519 -21512
rect 19557 -21546 19581 -21512
rect 19581 -21546 19591 -21512
rect 20215 -21546 20225 -21512
rect 20225 -21546 20249 -21512
rect 20287 -21546 20293 -21512
rect 20293 -21546 20321 -21512
rect 20359 -21546 20361 -21512
rect 20361 -21546 20393 -21512
rect 20431 -21546 20463 -21512
rect 20463 -21546 20465 -21512
rect 20503 -21546 20531 -21512
rect 20531 -21546 20537 -21512
rect 20575 -21546 20599 -21512
rect 20599 -21546 20609 -21512
rect 21233 -21546 21243 -21512
rect 21243 -21546 21267 -21512
rect 21305 -21546 21311 -21512
rect 21311 -21546 21339 -21512
rect 21377 -21546 21379 -21512
rect 21379 -21546 21411 -21512
rect 21449 -21546 21481 -21512
rect 21481 -21546 21483 -21512
rect 21521 -21546 21549 -21512
rect 21549 -21546 21555 -21512
rect 21593 -21546 21617 -21512
rect 21617 -21546 21627 -21512
rect 22251 -21546 22261 -21512
rect 22261 -21546 22285 -21512
rect 22323 -21546 22329 -21512
rect 22329 -21546 22357 -21512
rect 22395 -21546 22397 -21512
rect 22397 -21546 22429 -21512
rect 22467 -21546 22499 -21512
rect 22499 -21546 22501 -21512
rect 22539 -21546 22567 -21512
rect 22567 -21546 22573 -21512
rect 22611 -21546 22635 -21512
rect 22635 -21546 22645 -21512
rect -12289 -21597 -12255 -21595
rect -12289 -21629 -12255 -21597
rect 24855 -21529 24889 -21523
rect 24855 -21557 24889 -21529
rect -12289 -21699 -12255 -21667
rect -12289 -21701 -12255 -21699
rect 2580 -21629 2614 -21615
rect 2580 -21649 2614 -21629
rect 2580 -21697 2614 -21687
rect -12289 -21767 -12255 -21739
rect -12289 -21773 -12255 -21767
rect -9076 -21743 -9066 -21709
rect -9066 -21743 -9042 -21709
rect -9004 -21743 -8998 -21709
rect -8998 -21743 -8970 -21709
rect -8932 -21743 -8930 -21709
rect -8930 -21743 -8898 -21709
rect -8860 -21743 -8828 -21709
rect -8828 -21743 -8826 -21709
rect -8788 -21743 -8760 -21709
rect -8760 -21743 -8754 -21709
rect -8716 -21743 -8692 -21709
rect -8692 -21743 -8682 -21709
rect -8058 -21743 -8048 -21709
rect -8048 -21743 -8024 -21709
rect -7986 -21743 -7980 -21709
rect -7980 -21743 -7952 -21709
rect -7914 -21743 -7912 -21709
rect -7912 -21743 -7880 -21709
rect -7842 -21743 -7810 -21709
rect -7810 -21743 -7808 -21709
rect -7770 -21743 -7742 -21709
rect -7742 -21743 -7736 -21709
rect -7698 -21743 -7674 -21709
rect -7674 -21743 -7664 -21709
rect -7040 -21743 -7030 -21709
rect -7030 -21743 -7006 -21709
rect -6968 -21743 -6962 -21709
rect -6962 -21743 -6934 -21709
rect -6896 -21743 -6894 -21709
rect -6894 -21743 -6862 -21709
rect -6824 -21743 -6792 -21709
rect -6792 -21743 -6790 -21709
rect -6752 -21743 -6724 -21709
rect -6724 -21743 -6718 -21709
rect -6680 -21743 -6656 -21709
rect -6656 -21743 -6646 -21709
rect -6022 -21743 -6012 -21709
rect -6012 -21743 -5988 -21709
rect -5950 -21743 -5944 -21709
rect -5944 -21743 -5916 -21709
rect -5878 -21743 -5876 -21709
rect -5876 -21743 -5844 -21709
rect -5806 -21743 -5774 -21709
rect -5774 -21743 -5772 -21709
rect -5734 -21743 -5706 -21709
rect -5706 -21743 -5700 -21709
rect -5662 -21743 -5638 -21709
rect -5638 -21743 -5628 -21709
rect -5004 -21743 -4994 -21709
rect -4994 -21743 -4970 -21709
rect -4932 -21743 -4926 -21709
rect -4926 -21743 -4898 -21709
rect -4860 -21743 -4858 -21709
rect -4858 -21743 -4826 -21709
rect -4788 -21743 -4756 -21709
rect -4756 -21743 -4754 -21709
rect -4716 -21743 -4688 -21709
rect -4688 -21743 -4682 -21709
rect -4644 -21743 -4620 -21709
rect -4620 -21743 -4610 -21709
rect -3986 -21743 -3976 -21709
rect -3976 -21743 -3952 -21709
rect -3914 -21743 -3908 -21709
rect -3908 -21743 -3880 -21709
rect -3842 -21743 -3840 -21709
rect -3840 -21743 -3808 -21709
rect -3770 -21743 -3738 -21709
rect -3738 -21743 -3736 -21709
rect -3698 -21743 -3670 -21709
rect -3670 -21743 -3664 -21709
rect -3626 -21743 -3602 -21709
rect -3602 -21743 -3592 -21709
rect -2261 -21742 -2227 -21708
rect -1963 -21742 -1929 -21708
rect -1665 -21742 -1631 -21708
rect -1367 -21742 -1333 -21708
rect -1069 -21742 -1035 -21708
rect -771 -21742 -737 -21708
rect -473 -21742 -439 -21708
rect -175 -21742 -141 -21708
rect 123 -21742 157 -21708
rect 421 -21742 455 -21708
rect 719 -21742 753 -21708
rect 2580 -21721 2614 -21697
rect 2580 -21765 2614 -21759
rect -12289 -21835 -12255 -21811
rect -12289 -21845 -12255 -21835
rect -12289 -21903 -12255 -21883
rect -12289 -21917 -12255 -21903
rect -12289 -21971 -12255 -21955
rect -12289 -21989 -12255 -21971
rect -12289 -22039 -12255 -22027
rect -12289 -22061 -12255 -22039
rect -12289 -22107 -12255 -22099
rect -12289 -22133 -12255 -22107
rect -12289 -22175 -12255 -22171
rect -12289 -22205 -12255 -22175
rect -12289 -22277 -12255 -22243
rect -12289 -22345 -12255 -22315
rect -12289 -22349 -12255 -22345
rect -12289 -22413 -12255 -22387
rect -12289 -22421 -12255 -22413
rect -9405 -21826 -9371 -21812
rect -9405 -21846 -9371 -21826
rect -9405 -21894 -9371 -21884
rect -9405 -21918 -9371 -21894
rect -9405 -21962 -9371 -21956
rect -9405 -21990 -9371 -21962
rect -9405 -22030 -9371 -22028
rect -9405 -22062 -9371 -22030
rect -9405 -22132 -9371 -22100
rect -9405 -22134 -9371 -22132
rect -9405 -22200 -9371 -22172
rect -9405 -22206 -9371 -22200
rect -9405 -22268 -9371 -22244
rect -9405 -22278 -9371 -22268
rect -9405 -22336 -9371 -22316
rect -9405 -22350 -9371 -22336
rect -8387 -21826 -8353 -21812
rect -8387 -21846 -8353 -21826
rect -8387 -21894 -8353 -21884
rect -8387 -21918 -8353 -21894
rect -8387 -21962 -8353 -21956
rect -8387 -21990 -8353 -21962
rect -8387 -22030 -8353 -22028
rect -8387 -22062 -8353 -22030
rect -8387 -22132 -8353 -22100
rect -8387 -22134 -8353 -22132
rect -8387 -22200 -8353 -22172
rect -8387 -22206 -8353 -22200
rect -8387 -22268 -8353 -22244
rect -8387 -22278 -8353 -22268
rect -8387 -22336 -8353 -22316
rect -8387 -22350 -8353 -22336
rect -7369 -21826 -7335 -21812
rect -7369 -21846 -7335 -21826
rect -7369 -21894 -7335 -21884
rect -7369 -21918 -7335 -21894
rect -7369 -21962 -7335 -21956
rect -7369 -21990 -7335 -21962
rect -7369 -22030 -7335 -22028
rect -7369 -22062 -7335 -22030
rect -7369 -22132 -7335 -22100
rect -7369 -22134 -7335 -22132
rect -7369 -22200 -7335 -22172
rect -7369 -22206 -7335 -22200
rect -7369 -22268 -7335 -22244
rect -7369 -22278 -7335 -22268
rect -7369 -22336 -7335 -22316
rect -7369 -22350 -7335 -22336
rect -6351 -21826 -6317 -21812
rect -6351 -21846 -6317 -21826
rect -6351 -21894 -6317 -21884
rect -6351 -21918 -6317 -21894
rect -6351 -21962 -6317 -21956
rect -6351 -21990 -6317 -21962
rect -6351 -22030 -6317 -22028
rect -6351 -22062 -6317 -22030
rect -6351 -22132 -6317 -22100
rect -6351 -22134 -6317 -22132
rect -6351 -22200 -6317 -22172
rect -6351 -22206 -6317 -22200
rect -6351 -22268 -6317 -22244
rect -6351 -22278 -6317 -22268
rect -6351 -22336 -6317 -22316
rect -6351 -22350 -6317 -22336
rect -5333 -21826 -5299 -21812
rect -5333 -21846 -5299 -21826
rect -5333 -21894 -5299 -21884
rect -5333 -21918 -5299 -21894
rect -5333 -21962 -5299 -21956
rect -5333 -21990 -5299 -21962
rect -5333 -22030 -5299 -22028
rect -5333 -22062 -5299 -22030
rect -5333 -22132 -5299 -22100
rect -5333 -22134 -5299 -22132
rect -5333 -22200 -5299 -22172
rect -5333 -22206 -5299 -22200
rect -5333 -22268 -5299 -22244
rect -5333 -22278 -5299 -22268
rect -5333 -22336 -5299 -22316
rect -5333 -22350 -5299 -22336
rect -4315 -21826 -4281 -21812
rect -4315 -21846 -4281 -21826
rect -4315 -21894 -4281 -21884
rect -4315 -21918 -4281 -21894
rect -4315 -21962 -4281 -21956
rect -4315 -21990 -4281 -21962
rect -4315 -22030 -4281 -22028
rect -4315 -22062 -4281 -22030
rect -4315 -22132 -4281 -22100
rect -4315 -22134 -4281 -22132
rect -4315 -22200 -4281 -22172
rect -4315 -22206 -4281 -22200
rect -4315 -22268 -4281 -22244
rect -4315 -22278 -4281 -22268
rect -4315 -22336 -4281 -22316
rect -4315 -22350 -4281 -22336
rect -3297 -21826 -3263 -21812
rect -3297 -21846 -3263 -21826
rect -3297 -21894 -3263 -21884
rect -3297 -21918 -3263 -21894
rect -3297 -21962 -3263 -21956
rect -3297 -21990 -3263 -21962
rect -3297 -22030 -3263 -22028
rect -3297 -22062 -3263 -22030
rect -3297 -22132 -3263 -22100
rect -3297 -22134 -3263 -22132
rect -3297 -22200 -3263 -22172
rect -3297 -22206 -3263 -22200
rect -3297 -22268 -3263 -22244
rect -3297 -22278 -3263 -22268
rect -3297 -22336 -3263 -22316
rect -3297 -22350 -3263 -22336
rect -2410 -21825 -2376 -21811
rect -2410 -21845 -2376 -21825
rect -2410 -21893 -2376 -21883
rect -2410 -21917 -2376 -21893
rect -2410 -21961 -2376 -21955
rect -2410 -21989 -2376 -21961
rect -2410 -22029 -2376 -22027
rect -2410 -22061 -2376 -22029
rect -2410 -22131 -2376 -22099
rect -2410 -22133 -2376 -22131
rect -2410 -22199 -2376 -22171
rect -2410 -22205 -2376 -22199
rect -2410 -22267 -2376 -22243
rect -2410 -22277 -2376 -22267
rect -2410 -22335 -2376 -22315
rect -2410 -22349 -2376 -22335
rect -2112 -21825 -2078 -21811
rect -2112 -21845 -2078 -21825
rect -2112 -21893 -2078 -21883
rect -2112 -21917 -2078 -21893
rect -2112 -21961 -2078 -21955
rect -2112 -21989 -2078 -21961
rect -2112 -22029 -2078 -22027
rect -2112 -22061 -2078 -22029
rect -2112 -22131 -2078 -22099
rect -2112 -22133 -2078 -22131
rect -2112 -22199 -2078 -22171
rect -2112 -22205 -2078 -22199
rect -2112 -22267 -2078 -22243
rect -2112 -22277 -2078 -22267
rect -2112 -22335 -2078 -22315
rect -2112 -22349 -2078 -22335
rect -1814 -21825 -1780 -21811
rect -1814 -21845 -1780 -21825
rect -1814 -21893 -1780 -21883
rect -1814 -21917 -1780 -21893
rect -1814 -21961 -1780 -21955
rect -1814 -21989 -1780 -21961
rect -1814 -22029 -1780 -22027
rect -1814 -22061 -1780 -22029
rect -1814 -22131 -1780 -22099
rect -1814 -22133 -1780 -22131
rect -1814 -22199 -1780 -22171
rect -1814 -22205 -1780 -22199
rect -1814 -22267 -1780 -22243
rect -1814 -22277 -1780 -22267
rect -1814 -22335 -1780 -22315
rect -1814 -22349 -1780 -22335
rect -1516 -21825 -1482 -21811
rect -1516 -21845 -1482 -21825
rect -1516 -21893 -1482 -21883
rect -1516 -21917 -1482 -21893
rect -1516 -21961 -1482 -21955
rect -1516 -21989 -1482 -21961
rect -1516 -22029 -1482 -22027
rect -1516 -22061 -1482 -22029
rect -1516 -22131 -1482 -22099
rect -1516 -22133 -1482 -22131
rect -1516 -22199 -1482 -22171
rect -1516 -22205 -1482 -22199
rect -1516 -22267 -1482 -22243
rect -1516 -22277 -1482 -22267
rect -1516 -22335 -1482 -22315
rect -1516 -22349 -1482 -22335
rect -1218 -21825 -1184 -21811
rect -1218 -21845 -1184 -21825
rect -1218 -21893 -1184 -21883
rect -1218 -21917 -1184 -21893
rect -1218 -21961 -1184 -21955
rect -1218 -21989 -1184 -21961
rect -1218 -22029 -1184 -22027
rect -1218 -22061 -1184 -22029
rect -1218 -22131 -1184 -22099
rect -1218 -22133 -1184 -22131
rect -1218 -22199 -1184 -22171
rect -1218 -22205 -1184 -22199
rect -1218 -22267 -1184 -22243
rect -1218 -22277 -1184 -22267
rect -1218 -22335 -1184 -22315
rect -1218 -22349 -1184 -22335
rect -920 -21825 -886 -21811
rect -920 -21845 -886 -21825
rect -920 -21893 -886 -21883
rect -920 -21917 -886 -21893
rect -920 -21961 -886 -21955
rect -920 -21989 -886 -21961
rect -920 -22029 -886 -22027
rect -920 -22061 -886 -22029
rect -920 -22131 -886 -22099
rect -920 -22133 -886 -22131
rect -920 -22199 -886 -22171
rect -920 -22205 -886 -22199
rect -920 -22267 -886 -22243
rect -920 -22277 -886 -22267
rect -920 -22335 -886 -22315
rect -920 -22349 -886 -22335
rect -622 -21825 -588 -21811
rect -622 -21845 -588 -21825
rect -622 -21893 -588 -21883
rect -622 -21917 -588 -21893
rect -622 -21961 -588 -21955
rect -622 -21989 -588 -21961
rect -622 -22029 -588 -22027
rect -622 -22061 -588 -22029
rect -622 -22131 -588 -22099
rect -622 -22133 -588 -22131
rect -622 -22199 -588 -22171
rect -622 -22205 -588 -22199
rect -622 -22267 -588 -22243
rect -622 -22277 -588 -22267
rect -622 -22335 -588 -22315
rect -622 -22349 -588 -22335
rect -324 -21825 -290 -21811
rect -324 -21845 -290 -21825
rect -324 -21893 -290 -21883
rect -324 -21917 -290 -21893
rect -324 -21961 -290 -21955
rect -324 -21989 -290 -21961
rect -324 -22029 -290 -22027
rect -324 -22061 -290 -22029
rect -324 -22131 -290 -22099
rect -324 -22133 -290 -22131
rect -324 -22199 -290 -22171
rect -324 -22205 -290 -22199
rect -324 -22267 -290 -22243
rect -324 -22277 -290 -22267
rect -324 -22335 -290 -22315
rect -324 -22349 -290 -22335
rect -26 -21825 8 -21811
rect -26 -21845 8 -21825
rect -26 -21893 8 -21883
rect -26 -21917 8 -21893
rect -26 -21961 8 -21955
rect -26 -21989 8 -21961
rect -26 -22029 8 -22027
rect -26 -22061 8 -22029
rect -26 -22131 8 -22099
rect -26 -22133 8 -22131
rect -26 -22199 8 -22171
rect -26 -22205 8 -22199
rect -26 -22267 8 -22243
rect -26 -22277 8 -22267
rect -26 -22335 8 -22315
rect -26 -22349 8 -22335
rect 272 -21825 306 -21811
rect 272 -21845 306 -21825
rect 272 -21893 306 -21883
rect 272 -21917 306 -21893
rect 272 -21961 306 -21955
rect 272 -21989 306 -21961
rect 272 -22029 306 -22027
rect 272 -22061 306 -22029
rect 272 -22131 306 -22099
rect 272 -22133 306 -22131
rect 272 -22199 306 -22171
rect 272 -22205 306 -22199
rect 272 -22267 306 -22243
rect 272 -22277 306 -22267
rect 272 -22335 306 -22315
rect 272 -22349 306 -22335
rect 570 -21825 604 -21811
rect 570 -21845 604 -21825
rect 570 -21893 604 -21883
rect 570 -21917 604 -21893
rect 570 -21961 604 -21955
rect 570 -21989 604 -21961
rect 570 -22029 604 -22027
rect 570 -22061 604 -22029
rect 570 -22131 604 -22099
rect 570 -22133 604 -22131
rect 570 -22199 604 -22171
rect 570 -22205 604 -22199
rect 570 -22267 604 -22243
rect 570 -22277 604 -22267
rect 570 -22335 604 -22315
rect 570 -22349 604 -22335
rect 868 -21825 902 -21811
rect 868 -21845 902 -21825
rect 868 -21893 902 -21883
rect 868 -21917 902 -21893
rect 868 -21961 902 -21955
rect 868 -21989 902 -21961
rect 868 -22029 902 -22027
rect 868 -22061 902 -22029
rect 868 -22131 902 -22099
rect 868 -22133 902 -22131
rect 868 -22199 902 -22171
rect 2580 -21793 2614 -21765
rect 2580 -21833 2614 -21831
rect 2580 -21865 2614 -21833
rect 2580 -21935 2614 -21903
rect 2580 -21937 2614 -21935
rect 2580 -22003 2614 -21975
rect 2580 -22009 2614 -22003
rect 2580 -22071 2614 -22047
rect 2580 -22081 2614 -22071
rect 2580 -22139 2614 -22119
rect 2580 -22153 2614 -22139
rect 3598 -21629 3632 -21615
rect 3598 -21649 3632 -21629
rect 3598 -21697 3632 -21687
rect 3598 -21721 3632 -21697
rect 3598 -21765 3632 -21759
rect 3598 -21793 3632 -21765
rect 3598 -21833 3632 -21831
rect 3598 -21865 3632 -21833
rect 3598 -21935 3632 -21903
rect 3598 -21937 3632 -21935
rect 3598 -22003 3632 -21975
rect 3598 -22009 3632 -22003
rect 3598 -22071 3632 -22047
rect 3598 -22081 3632 -22071
rect 3598 -22139 3632 -22119
rect 3598 -22153 3632 -22139
rect 4616 -21629 4650 -21615
rect 4616 -21649 4650 -21629
rect 4616 -21697 4650 -21687
rect 4616 -21721 4650 -21697
rect 4616 -21765 4650 -21759
rect 4616 -21793 4650 -21765
rect 4616 -21833 4650 -21831
rect 4616 -21865 4650 -21833
rect 4616 -21935 4650 -21903
rect 4616 -21937 4650 -21935
rect 4616 -22003 4650 -21975
rect 4616 -22009 4650 -22003
rect 4616 -22071 4650 -22047
rect 4616 -22081 4650 -22071
rect 4616 -22139 4650 -22119
rect 4616 -22153 4650 -22139
rect 5634 -21629 5668 -21615
rect 5634 -21649 5668 -21629
rect 5634 -21697 5668 -21687
rect 5634 -21721 5668 -21697
rect 5634 -21765 5668 -21759
rect 5634 -21793 5668 -21765
rect 5634 -21833 5668 -21831
rect 5634 -21865 5668 -21833
rect 5634 -21935 5668 -21903
rect 5634 -21937 5668 -21935
rect 5634 -22003 5668 -21975
rect 5634 -22009 5668 -22003
rect 5634 -22071 5668 -22047
rect 5634 -22081 5668 -22071
rect 5634 -22139 5668 -22119
rect 5634 -22153 5668 -22139
rect 6652 -21629 6686 -21615
rect 6652 -21649 6686 -21629
rect 6652 -21697 6686 -21687
rect 6652 -21721 6686 -21697
rect 6652 -21765 6686 -21759
rect 6652 -21793 6686 -21765
rect 6652 -21833 6686 -21831
rect 6652 -21865 6686 -21833
rect 6652 -21935 6686 -21903
rect 6652 -21937 6686 -21935
rect 6652 -22003 6686 -21975
rect 6652 -22009 6686 -22003
rect 6652 -22071 6686 -22047
rect 6652 -22081 6686 -22071
rect 6652 -22139 6686 -22119
rect 6652 -22153 6686 -22139
rect 7670 -21629 7704 -21615
rect 7670 -21649 7704 -21629
rect 7670 -21697 7704 -21687
rect 7670 -21721 7704 -21697
rect 7670 -21765 7704 -21759
rect 7670 -21793 7704 -21765
rect 7670 -21833 7704 -21831
rect 7670 -21865 7704 -21833
rect 7670 -21935 7704 -21903
rect 7670 -21937 7704 -21935
rect 7670 -22003 7704 -21975
rect 7670 -22009 7704 -22003
rect 7670 -22071 7704 -22047
rect 7670 -22081 7704 -22071
rect 7670 -22139 7704 -22119
rect 7670 -22153 7704 -22139
rect 8688 -21629 8722 -21615
rect 8688 -21649 8722 -21629
rect 8688 -21697 8722 -21687
rect 8688 -21721 8722 -21697
rect 8688 -21765 8722 -21759
rect 8688 -21793 8722 -21765
rect 8688 -21833 8722 -21831
rect 8688 -21865 8722 -21833
rect 8688 -21935 8722 -21903
rect 8688 -21937 8722 -21935
rect 8688 -22003 8722 -21975
rect 8688 -22009 8722 -22003
rect 8688 -22071 8722 -22047
rect 8688 -22081 8722 -22071
rect 8688 -22139 8722 -22119
rect 8688 -22153 8722 -22139
rect 9706 -21629 9740 -21615
rect 9706 -21649 9740 -21629
rect 9706 -21697 9740 -21687
rect 9706 -21721 9740 -21697
rect 9706 -21765 9740 -21759
rect 9706 -21793 9740 -21765
rect 9706 -21833 9740 -21831
rect 9706 -21865 9740 -21833
rect 9706 -21935 9740 -21903
rect 9706 -21937 9740 -21935
rect 9706 -22003 9740 -21975
rect 9706 -22009 9740 -22003
rect 9706 -22071 9740 -22047
rect 9706 -22081 9740 -22071
rect 9706 -22139 9740 -22119
rect 9706 -22153 9740 -22139
rect 10724 -21629 10758 -21615
rect 10724 -21649 10758 -21629
rect 10724 -21697 10758 -21687
rect 10724 -21721 10758 -21697
rect 10724 -21765 10758 -21759
rect 10724 -21793 10758 -21765
rect 10724 -21833 10758 -21831
rect 10724 -21865 10758 -21833
rect 10724 -21935 10758 -21903
rect 10724 -21937 10758 -21935
rect 10724 -22003 10758 -21975
rect 10724 -22009 10758 -22003
rect 10724 -22071 10758 -22047
rect 10724 -22081 10758 -22071
rect 10724 -22139 10758 -22119
rect 10724 -22153 10758 -22139
rect 11742 -21629 11776 -21615
rect 11742 -21649 11776 -21629
rect 11742 -21697 11776 -21687
rect 11742 -21721 11776 -21697
rect 11742 -21765 11776 -21759
rect 11742 -21793 11776 -21765
rect 11742 -21833 11776 -21831
rect 11742 -21865 11776 -21833
rect 11742 -21935 11776 -21903
rect 11742 -21937 11776 -21935
rect 11742 -22003 11776 -21975
rect 11742 -22009 11776 -22003
rect 11742 -22071 11776 -22047
rect 11742 -22081 11776 -22071
rect 11742 -22139 11776 -22119
rect 11742 -22153 11776 -22139
rect 12760 -21629 12794 -21615
rect 12760 -21649 12794 -21629
rect 12760 -21697 12794 -21687
rect 12760 -21721 12794 -21697
rect 12760 -21765 12794 -21759
rect 12760 -21793 12794 -21765
rect 12760 -21833 12794 -21831
rect 12760 -21865 12794 -21833
rect 12760 -21935 12794 -21903
rect 12760 -21937 12794 -21935
rect 12760 -22003 12794 -21975
rect 12760 -22009 12794 -22003
rect 12760 -22071 12794 -22047
rect 12760 -22081 12794 -22071
rect 12760 -22139 12794 -22119
rect 12760 -22153 12794 -22139
rect 13778 -21629 13812 -21615
rect 13778 -21649 13812 -21629
rect 13778 -21697 13812 -21687
rect 13778 -21721 13812 -21697
rect 13778 -21765 13812 -21759
rect 13778 -21793 13812 -21765
rect 13778 -21833 13812 -21831
rect 13778 -21865 13812 -21833
rect 13778 -21935 13812 -21903
rect 13778 -21937 13812 -21935
rect 13778 -22003 13812 -21975
rect 13778 -22009 13812 -22003
rect 13778 -22071 13812 -22047
rect 13778 -22081 13812 -22071
rect 13778 -22139 13812 -22119
rect 13778 -22153 13812 -22139
rect 14796 -21629 14830 -21615
rect 14796 -21649 14830 -21629
rect 14796 -21697 14830 -21687
rect 14796 -21721 14830 -21697
rect 14796 -21765 14830 -21759
rect 14796 -21793 14830 -21765
rect 14796 -21833 14830 -21831
rect 14796 -21865 14830 -21833
rect 14796 -21935 14830 -21903
rect 14796 -21937 14830 -21935
rect 14796 -22003 14830 -21975
rect 14796 -22009 14830 -22003
rect 14796 -22071 14830 -22047
rect 14796 -22081 14830 -22071
rect 14796 -22139 14830 -22119
rect 14796 -22153 14830 -22139
rect 15814 -21629 15848 -21615
rect 15814 -21649 15848 -21629
rect 15814 -21697 15848 -21687
rect 15814 -21721 15848 -21697
rect 15814 -21765 15848 -21759
rect 15814 -21793 15848 -21765
rect 15814 -21833 15848 -21831
rect 15814 -21865 15848 -21833
rect 15814 -21935 15848 -21903
rect 15814 -21937 15848 -21935
rect 15814 -22003 15848 -21975
rect 15814 -22009 15848 -22003
rect 15814 -22071 15848 -22047
rect 15814 -22081 15848 -22071
rect 15814 -22139 15848 -22119
rect 15814 -22153 15848 -22139
rect 16832 -21629 16866 -21615
rect 16832 -21649 16866 -21629
rect 16832 -21697 16866 -21687
rect 16832 -21721 16866 -21697
rect 16832 -21765 16866 -21759
rect 16832 -21793 16866 -21765
rect 16832 -21833 16866 -21831
rect 16832 -21865 16866 -21833
rect 16832 -21935 16866 -21903
rect 16832 -21937 16866 -21935
rect 16832 -22003 16866 -21975
rect 16832 -22009 16866 -22003
rect 16832 -22071 16866 -22047
rect 16832 -22081 16866 -22071
rect 16832 -22139 16866 -22119
rect 16832 -22153 16866 -22139
rect 17850 -21629 17884 -21615
rect 17850 -21649 17884 -21629
rect 17850 -21697 17884 -21687
rect 17850 -21721 17884 -21697
rect 17850 -21765 17884 -21759
rect 17850 -21793 17884 -21765
rect 17850 -21833 17884 -21831
rect 17850 -21865 17884 -21833
rect 17850 -21935 17884 -21903
rect 17850 -21937 17884 -21935
rect 17850 -22003 17884 -21975
rect 17850 -22009 17884 -22003
rect 17850 -22071 17884 -22047
rect 17850 -22081 17884 -22071
rect 17850 -22139 17884 -22119
rect 17850 -22153 17884 -22139
rect 18868 -21629 18902 -21615
rect 18868 -21649 18902 -21629
rect 18868 -21697 18902 -21687
rect 18868 -21721 18902 -21697
rect 18868 -21765 18902 -21759
rect 18868 -21793 18902 -21765
rect 18868 -21833 18902 -21831
rect 18868 -21865 18902 -21833
rect 18868 -21935 18902 -21903
rect 18868 -21937 18902 -21935
rect 18868 -22003 18902 -21975
rect 18868 -22009 18902 -22003
rect 18868 -22071 18902 -22047
rect 18868 -22081 18902 -22071
rect 18868 -22139 18902 -22119
rect 18868 -22153 18902 -22139
rect 19886 -21629 19920 -21615
rect 19886 -21649 19920 -21629
rect 19886 -21697 19920 -21687
rect 19886 -21721 19920 -21697
rect 19886 -21765 19920 -21759
rect 19886 -21793 19920 -21765
rect 19886 -21833 19920 -21831
rect 19886 -21865 19920 -21833
rect 19886 -21935 19920 -21903
rect 19886 -21937 19920 -21935
rect 19886 -22003 19920 -21975
rect 19886 -22009 19920 -22003
rect 19886 -22071 19920 -22047
rect 19886 -22081 19920 -22071
rect 19886 -22139 19920 -22119
rect 19886 -22153 19920 -22139
rect 20904 -21629 20938 -21615
rect 20904 -21649 20938 -21629
rect 20904 -21697 20938 -21687
rect 20904 -21721 20938 -21697
rect 20904 -21765 20938 -21759
rect 20904 -21793 20938 -21765
rect 20904 -21833 20938 -21831
rect 20904 -21865 20938 -21833
rect 20904 -21935 20938 -21903
rect 20904 -21937 20938 -21935
rect 20904 -22003 20938 -21975
rect 20904 -22009 20938 -22003
rect 20904 -22071 20938 -22047
rect 20904 -22081 20938 -22071
rect 20904 -22139 20938 -22119
rect 20904 -22153 20938 -22139
rect 21922 -21629 21956 -21615
rect 21922 -21649 21956 -21629
rect 21922 -21697 21956 -21687
rect 21922 -21721 21956 -21697
rect 21922 -21765 21956 -21759
rect 21922 -21793 21956 -21765
rect 21922 -21833 21956 -21831
rect 21922 -21865 21956 -21833
rect 21922 -21935 21956 -21903
rect 21922 -21937 21956 -21935
rect 21922 -22003 21956 -21975
rect 21922 -22009 21956 -22003
rect 21922 -22071 21956 -22047
rect 21922 -22081 21956 -22071
rect 21922 -22139 21956 -22119
rect 21922 -22153 21956 -22139
rect 22940 -21629 22974 -21615
rect 22940 -21649 22974 -21629
rect 22940 -21697 22974 -21687
rect 22940 -21721 22974 -21697
rect 22940 -21765 22974 -21759
rect 22940 -21793 22974 -21765
rect 22940 -21833 22974 -21831
rect 22940 -21865 22974 -21833
rect 22940 -21935 22974 -21903
rect 22940 -21937 22974 -21935
rect 22940 -22003 22974 -21975
rect 22940 -22009 22974 -22003
rect 22940 -22071 22974 -22047
rect 22940 -22081 22974 -22071
rect 22940 -22139 22974 -22119
rect 22940 -22153 22974 -22139
rect 24855 -21597 24889 -21595
rect 24855 -21629 24889 -21597
rect 24855 -21699 24889 -21667
rect 24855 -21701 24889 -21699
rect 24855 -21767 24889 -21739
rect 24855 -21773 24889 -21767
rect 24855 -21835 24889 -21811
rect 24855 -21845 24889 -21835
rect 24855 -21903 24889 -21883
rect 24855 -21917 24889 -21903
rect 24855 -21971 24889 -21955
rect 24855 -21989 24889 -21971
rect 24855 -22039 24889 -22027
rect 24855 -22061 24889 -22039
rect 24855 -22107 24889 -22099
rect 24855 -22133 24889 -22107
rect 868 -22205 902 -22199
rect 24855 -22175 24889 -22171
rect 24855 -22205 24889 -22175
rect 868 -22267 902 -22243
rect 2909 -22256 2919 -22222
rect 2919 -22256 2943 -22222
rect 2981 -22256 2987 -22222
rect 2987 -22256 3015 -22222
rect 3053 -22256 3055 -22222
rect 3055 -22256 3087 -22222
rect 3125 -22256 3157 -22222
rect 3157 -22256 3159 -22222
rect 3197 -22256 3225 -22222
rect 3225 -22256 3231 -22222
rect 3269 -22256 3293 -22222
rect 3293 -22256 3303 -22222
rect 3927 -22256 3937 -22222
rect 3937 -22256 3961 -22222
rect 3999 -22256 4005 -22222
rect 4005 -22256 4033 -22222
rect 4071 -22256 4073 -22222
rect 4073 -22256 4105 -22222
rect 4143 -22256 4175 -22222
rect 4175 -22256 4177 -22222
rect 4215 -22256 4243 -22222
rect 4243 -22256 4249 -22222
rect 4287 -22256 4311 -22222
rect 4311 -22256 4321 -22222
rect 4945 -22256 4955 -22222
rect 4955 -22256 4979 -22222
rect 5017 -22256 5023 -22222
rect 5023 -22256 5051 -22222
rect 5089 -22256 5091 -22222
rect 5091 -22256 5123 -22222
rect 5161 -22256 5193 -22222
rect 5193 -22256 5195 -22222
rect 5233 -22256 5261 -22222
rect 5261 -22256 5267 -22222
rect 5305 -22256 5329 -22222
rect 5329 -22256 5339 -22222
rect 5963 -22256 5973 -22222
rect 5973 -22256 5997 -22222
rect 6035 -22256 6041 -22222
rect 6041 -22256 6069 -22222
rect 6107 -22256 6109 -22222
rect 6109 -22256 6141 -22222
rect 6179 -22256 6211 -22222
rect 6211 -22256 6213 -22222
rect 6251 -22256 6279 -22222
rect 6279 -22256 6285 -22222
rect 6323 -22256 6347 -22222
rect 6347 -22256 6357 -22222
rect 6981 -22256 6991 -22222
rect 6991 -22256 7015 -22222
rect 7053 -22256 7059 -22222
rect 7059 -22256 7087 -22222
rect 7125 -22256 7127 -22222
rect 7127 -22256 7159 -22222
rect 7197 -22256 7229 -22222
rect 7229 -22256 7231 -22222
rect 7269 -22256 7297 -22222
rect 7297 -22256 7303 -22222
rect 7341 -22256 7365 -22222
rect 7365 -22256 7375 -22222
rect 7999 -22256 8009 -22222
rect 8009 -22256 8033 -22222
rect 8071 -22256 8077 -22222
rect 8077 -22256 8105 -22222
rect 8143 -22256 8145 -22222
rect 8145 -22256 8177 -22222
rect 8215 -22256 8247 -22222
rect 8247 -22256 8249 -22222
rect 8287 -22256 8315 -22222
rect 8315 -22256 8321 -22222
rect 8359 -22256 8383 -22222
rect 8383 -22256 8393 -22222
rect 9017 -22256 9027 -22222
rect 9027 -22256 9051 -22222
rect 9089 -22256 9095 -22222
rect 9095 -22256 9123 -22222
rect 9161 -22256 9163 -22222
rect 9163 -22256 9195 -22222
rect 9233 -22256 9265 -22222
rect 9265 -22256 9267 -22222
rect 9305 -22256 9333 -22222
rect 9333 -22256 9339 -22222
rect 9377 -22256 9401 -22222
rect 9401 -22256 9411 -22222
rect 10035 -22256 10045 -22222
rect 10045 -22256 10069 -22222
rect 10107 -22256 10113 -22222
rect 10113 -22256 10141 -22222
rect 10179 -22256 10181 -22222
rect 10181 -22256 10213 -22222
rect 10251 -22256 10283 -22222
rect 10283 -22256 10285 -22222
rect 10323 -22256 10351 -22222
rect 10351 -22256 10357 -22222
rect 10395 -22256 10419 -22222
rect 10419 -22256 10429 -22222
rect 11053 -22256 11063 -22222
rect 11063 -22256 11087 -22222
rect 11125 -22256 11131 -22222
rect 11131 -22256 11159 -22222
rect 11197 -22256 11199 -22222
rect 11199 -22256 11231 -22222
rect 11269 -22256 11301 -22222
rect 11301 -22256 11303 -22222
rect 11341 -22256 11369 -22222
rect 11369 -22256 11375 -22222
rect 11413 -22256 11437 -22222
rect 11437 -22256 11447 -22222
rect 12071 -22256 12081 -22222
rect 12081 -22256 12105 -22222
rect 12143 -22256 12149 -22222
rect 12149 -22256 12177 -22222
rect 12215 -22256 12217 -22222
rect 12217 -22256 12249 -22222
rect 12287 -22256 12319 -22222
rect 12319 -22256 12321 -22222
rect 12359 -22256 12387 -22222
rect 12387 -22256 12393 -22222
rect 12431 -22256 12455 -22222
rect 12455 -22256 12465 -22222
rect 13089 -22256 13099 -22222
rect 13099 -22256 13123 -22222
rect 13161 -22256 13167 -22222
rect 13167 -22256 13195 -22222
rect 13233 -22256 13235 -22222
rect 13235 -22256 13267 -22222
rect 13305 -22256 13337 -22222
rect 13337 -22256 13339 -22222
rect 13377 -22256 13405 -22222
rect 13405 -22256 13411 -22222
rect 13449 -22256 13473 -22222
rect 13473 -22256 13483 -22222
rect 14107 -22256 14117 -22222
rect 14117 -22256 14141 -22222
rect 14179 -22256 14185 -22222
rect 14185 -22256 14213 -22222
rect 14251 -22256 14253 -22222
rect 14253 -22256 14285 -22222
rect 14323 -22256 14355 -22222
rect 14355 -22256 14357 -22222
rect 14395 -22256 14423 -22222
rect 14423 -22256 14429 -22222
rect 14467 -22256 14491 -22222
rect 14491 -22256 14501 -22222
rect 15125 -22256 15135 -22222
rect 15135 -22256 15159 -22222
rect 15197 -22256 15203 -22222
rect 15203 -22256 15231 -22222
rect 15269 -22256 15271 -22222
rect 15271 -22256 15303 -22222
rect 15341 -22256 15373 -22222
rect 15373 -22256 15375 -22222
rect 15413 -22256 15441 -22222
rect 15441 -22256 15447 -22222
rect 15485 -22256 15509 -22222
rect 15509 -22256 15519 -22222
rect 16143 -22256 16153 -22222
rect 16153 -22256 16177 -22222
rect 16215 -22256 16221 -22222
rect 16221 -22256 16249 -22222
rect 16287 -22256 16289 -22222
rect 16289 -22256 16321 -22222
rect 16359 -22256 16391 -22222
rect 16391 -22256 16393 -22222
rect 16431 -22256 16459 -22222
rect 16459 -22256 16465 -22222
rect 16503 -22256 16527 -22222
rect 16527 -22256 16537 -22222
rect 17161 -22256 17171 -22222
rect 17171 -22256 17195 -22222
rect 17233 -22256 17239 -22222
rect 17239 -22256 17267 -22222
rect 17305 -22256 17307 -22222
rect 17307 -22256 17339 -22222
rect 17377 -22256 17409 -22222
rect 17409 -22256 17411 -22222
rect 17449 -22256 17477 -22222
rect 17477 -22256 17483 -22222
rect 17521 -22256 17545 -22222
rect 17545 -22256 17555 -22222
rect 18179 -22256 18189 -22222
rect 18189 -22256 18213 -22222
rect 18251 -22256 18257 -22222
rect 18257 -22256 18285 -22222
rect 18323 -22256 18325 -22222
rect 18325 -22256 18357 -22222
rect 18395 -22256 18427 -22222
rect 18427 -22256 18429 -22222
rect 18467 -22256 18495 -22222
rect 18495 -22256 18501 -22222
rect 18539 -22256 18563 -22222
rect 18563 -22256 18573 -22222
rect 19197 -22256 19207 -22222
rect 19207 -22256 19231 -22222
rect 19269 -22256 19275 -22222
rect 19275 -22256 19303 -22222
rect 19341 -22256 19343 -22222
rect 19343 -22256 19375 -22222
rect 19413 -22256 19445 -22222
rect 19445 -22256 19447 -22222
rect 19485 -22256 19513 -22222
rect 19513 -22256 19519 -22222
rect 19557 -22256 19581 -22222
rect 19581 -22256 19591 -22222
rect 20215 -22256 20225 -22222
rect 20225 -22256 20249 -22222
rect 20287 -22256 20293 -22222
rect 20293 -22256 20321 -22222
rect 20359 -22256 20361 -22222
rect 20361 -22256 20393 -22222
rect 20431 -22256 20463 -22222
rect 20463 -22256 20465 -22222
rect 20503 -22256 20531 -22222
rect 20531 -22256 20537 -22222
rect 20575 -22256 20599 -22222
rect 20599 -22256 20609 -22222
rect 21233 -22256 21243 -22222
rect 21243 -22256 21267 -22222
rect 21305 -22256 21311 -22222
rect 21311 -22256 21339 -22222
rect 21521 -22256 21549 -22222
rect 21549 -22256 21555 -22222
rect 21593 -22256 21617 -22222
rect 21617 -22256 21627 -22222
rect 22251 -22256 22261 -22222
rect 22261 -22256 22285 -22222
rect 22323 -22256 22329 -22222
rect 22329 -22256 22357 -22222
rect 22395 -22256 22397 -22222
rect 22397 -22256 22429 -22222
rect 22467 -22256 22499 -22222
rect 22499 -22256 22501 -22222
rect 22539 -22256 22567 -22222
rect 22567 -22256 22573 -22222
rect 22611 -22256 22635 -22222
rect 22635 -22256 22645 -22222
rect 868 -22277 902 -22267
rect 868 -22335 902 -22315
rect 868 -22349 902 -22335
rect 24855 -22277 24889 -22243
rect 24855 -22345 24889 -22315
rect 24855 -22349 24889 -22345
rect -12289 -22481 -12255 -22459
rect -12289 -22493 -12255 -22481
rect -9076 -22453 -9066 -22419
rect -9066 -22453 -9042 -22419
rect -9004 -22453 -8998 -22419
rect -8998 -22453 -8970 -22419
rect -8932 -22453 -8930 -22419
rect -8930 -22453 -8898 -22419
rect -8860 -22453 -8828 -22419
rect -8828 -22453 -8826 -22419
rect -8788 -22453 -8760 -22419
rect -8760 -22453 -8754 -22419
rect -8716 -22453 -8692 -22419
rect -8692 -22453 -8682 -22419
rect -8058 -22453 -8048 -22419
rect -8048 -22453 -8024 -22419
rect -7986 -22453 -7980 -22419
rect -7980 -22453 -7952 -22419
rect -7914 -22453 -7912 -22419
rect -7912 -22453 -7880 -22419
rect -7842 -22453 -7810 -22419
rect -7810 -22453 -7808 -22419
rect -7770 -22453 -7742 -22419
rect -7742 -22453 -7736 -22419
rect -7698 -22453 -7674 -22419
rect -7674 -22453 -7664 -22419
rect -7040 -22453 -7030 -22419
rect -7030 -22453 -7006 -22419
rect -6968 -22453 -6962 -22419
rect -6962 -22453 -6934 -22419
rect -6896 -22453 -6894 -22419
rect -6894 -22453 -6862 -22419
rect -6824 -22453 -6792 -22419
rect -6792 -22453 -6790 -22419
rect -6752 -22453 -6724 -22419
rect -6724 -22453 -6718 -22419
rect -6680 -22453 -6656 -22419
rect -6656 -22453 -6646 -22419
rect -6022 -22453 -6012 -22419
rect -6012 -22453 -5988 -22419
rect -5950 -22453 -5944 -22419
rect -5944 -22453 -5916 -22419
rect -5878 -22453 -5876 -22419
rect -5876 -22453 -5844 -22419
rect -5806 -22453 -5774 -22419
rect -5774 -22453 -5772 -22419
rect -5734 -22453 -5706 -22419
rect -5706 -22453 -5700 -22419
rect -5662 -22453 -5638 -22419
rect -5638 -22453 -5628 -22419
rect -5004 -22453 -4994 -22419
rect -4994 -22453 -4970 -22419
rect -4932 -22453 -4926 -22419
rect -4926 -22453 -4898 -22419
rect -4860 -22453 -4858 -22419
rect -4858 -22453 -4826 -22419
rect -4788 -22453 -4756 -22419
rect -4756 -22453 -4754 -22419
rect -4716 -22453 -4688 -22419
rect -4688 -22453 -4682 -22419
rect -4644 -22453 -4620 -22419
rect -4620 -22453 -4610 -22419
rect -3986 -22453 -3976 -22419
rect -3976 -22453 -3952 -22419
rect -3914 -22453 -3908 -22419
rect -3908 -22453 -3880 -22419
rect -3842 -22453 -3840 -22419
rect -3840 -22453 -3808 -22419
rect -3770 -22453 -3738 -22419
rect -3738 -22453 -3736 -22419
rect -3698 -22453 -3670 -22419
rect -3670 -22453 -3664 -22419
rect -3626 -22453 -3602 -22419
rect -3602 -22453 -3592 -22419
rect -2261 -22452 -2227 -22418
rect -1963 -22452 -1929 -22418
rect -1665 -22452 -1631 -22418
rect -1367 -22452 -1333 -22418
rect -1069 -22452 -1035 -22418
rect -771 -22452 -737 -22418
rect -473 -22452 -439 -22418
rect -175 -22452 -141 -22418
rect 123 -22452 157 -22418
rect 421 -22452 455 -22418
rect 719 -22452 753 -22418
rect 24855 -22413 24889 -22387
rect 24855 -22421 24889 -22413
rect -12289 -22549 -12255 -22531
rect -12289 -22565 -12255 -22549
rect -12289 -22617 -12255 -22603
rect -12289 -22637 -12255 -22617
rect -12289 -22685 -12255 -22675
rect -12289 -22709 -12255 -22685
rect -12289 -22753 -12255 -22747
rect -12289 -22781 -12255 -22753
rect 24855 -22481 24889 -22459
rect 24855 -22493 24889 -22481
rect 24855 -22549 24889 -22531
rect 24855 -22565 24889 -22549
rect 24855 -22617 24889 -22603
rect 24855 -22637 24889 -22617
rect 24855 -22685 24889 -22675
rect 24855 -22709 24889 -22685
rect 2909 -22780 2919 -22746
rect 2919 -22780 2943 -22746
rect 2981 -22780 2987 -22746
rect 2987 -22780 3015 -22746
rect 3053 -22780 3055 -22746
rect 3055 -22780 3087 -22746
rect 3125 -22780 3157 -22746
rect 3157 -22780 3159 -22746
rect 3197 -22780 3225 -22746
rect 3225 -22780 3231 -22746
rect 3269 -22780 3293 -22746
rect 3293 -22780 3303 -22746
rect 3927 -22780 3937 -22746
rect 3937 -22780 3961 -22746
rect 3999 -22780 4005 -22746
rect 4005 -22780 4033 -22746
rect 4071 -22780 4073 -22746
rect 4073 -22780 4105 -22746
rect 4143 -22780 4175 -22746
rect 4175 -22780 4177 -22746
rect 4215 -22780 4243 -22746
rect 4243 -22780 4249 -22746
rect 4287 -22780 4311 -22746
rect 4311 -22780 4321 -22746
rect 4945 -22780 4955 -22746
rect 4955 -22780 4979 -22746
rect 5017 -22780 5023 -22746
rect 5023 -22780 5051 -22746
rect 5089 -22780 5091 -22746
rect 5091 -22780 5123 -22746
rect 5161 -22780 5193 -22746
rect 5193 -22780 5195 -22746
rect 5233 -22780 5261 -22746
rect 5261 -22780 5267 -22746
rect 5305 -22780 5329 -22746
rect 5329 -22780 5339 -22746
rect 5963 -22780 5973 -22746
rect 5973 -22780 5997 -22746
rect 6035 -22780 6041 -22746
rect 6041 -22780 6069 -22746
rect 6107 -22780 6109 -22746
rect 6109 -22780 6141 -22746
rect 6179 -22780 6211 -22746
rect 6211 -22780 6213 -22746
rect 6251 -22780 6279 -22746
rect 6279 -22780 6285 -22746
rect 6323 -22780 6347 -22746
rect 6347 -22780 6357 -22746
rect 6981 -22780 6991 -22746
rect 6991 -22780 7015 -22746
rect 7053 -22780 7059 -22746
rect 7059 -22780 7087 -22746
rect 7125 -22780 7127 -22746
rect 7127 -22780 7159 -22746
rect 7197 -22780 7229 -22746
rect 7229 -22780 7231 -22746
rect 7269 -22780 7297 -22746
rect 7297 -22780 7303 -22746
rect 7341 -22780 7365 -22746
rect 7365 -22780 7375 -22746
rect 7999 -22780 8009 -22746
rect 8009 -22780 8033 -22746
rect 8071 -22780 8077 -22746
rect 8077 -22780 8105 -22746
rect 8143 -22780 8145 -22746
rect 8145 -22780 8177 -22746
rect 8215 -22780 8247 -22746
rect 8247 -22780 8249 -22746
rect 8287 -22780 8315 -22746
rect 8315 -22780 8321 -22746
rect 8359 -22780 8383 -22746
rect 8383 -22780 8393 -22746
rect 9017 -22780 9027 -22746
rect 9027 -22780 9051 -22746
rect 9089 -22780 9095 -22746
rect 9095 -22780 9123 -22746
rect 9161 -22780 9163 -22746
rect 9163 -22780 9195 -22746
rect 9233 -22780 9265 -22746
rect 9265 -22780 9267 -22746
rect 9305 -22780 9333 -22746
rect 9333 -22780 9339 -22746
rect 9377 -22780 9401 -22746
rect 9401 -22780 9411 -22746
rect 10035 -22780 10045 -22746
rect 10045 -22780 10069 -22746
rect 10107 -22780 10113 -22746
rect 10113 -22780 10141 -22746
rect 10179 -22780 10181 -22746
rect 10181 -22780 10213 -22746
rect 10251 -22780 10283 -22746
rect 10283 -22780 10285 -22746
rect 10323 -22780 10351 -22746
rect 10351 -22780 10357 -22746
rect 10395 -22780 10419 -22746
rect 10419 -22780 10429 -22746
rect 11053 -22780 11063 -22746
rect 11063 -22780 11087 -22746
rect 11125 -22780 11131 -22746
rect 11131 -22780 11159 -22746
rect 11197 -22780 11199 -22746
rect 11199 -22780 11231 -22746
rect 11269 -22780 11301 -22746
rect 11301 -22780 11303 -22746
rect 11341 -22780 11369 -22746
rect 11369 -22780 11375 -22746
rect 11413 -22780 11437 -22746
rect 11437 -22780 11447 -22746
rect 12071 -22780 12081 -22746
rect 12081 -22780 12105 -22746
rect 12143 -22780 12149 -22746
rect 12149 -22780 12177 -22746
rect 12215 -22780 12217 -22746
rect 12217 -22780 12249 -22746
rect 12287 -22780 12319 -22746
rect 12319 -22780 12321 -22746
rect 12359 -22780 12387 -22746
rect 12387 -22780 12393 -22746
rect 12431 -22780 12455 -22746
rect 12455 -22780 12465 -22746
rect 13089 -22780 13099 -22746
rect 13099 -22780 13123 -22746
rect 13161 -22780 13167 -22746
rect 13167 -22780 13195 -22746
rect 13233 -22780 13235 -22746
rect 13235 -22780 13267 -22746
rect 13305 -22780 13337 -22746
rect 13337 -22780 13339 -22746
rect 13377 -22780 13405 -22746
rect 13405 -22780 13411 -22746
rect 13449 -22780 13473 -22746
rect 13473 -22780 13483 -22746
rect 14107 -22780 14117 -22746
rect 14117 -22780 14141 -22746
rect 14179 -22780 14185 -22746
rect 14185 -22780 14213 -22746
rect 14251 -22780 14253 -22746
rect 14253 -22780 14285 -22746
rect 14323 -22780 14355 -22746
rect 14355 -22780 14357 -22746
rect 14395 -22780 14423 -22746
rect 14423 -22780 14429 -22746
rect 14467 -22780 14491 -22746
rect 14491 -22780 14501 -22746
rect 15125 -22780 15135 -22746
rect 15135 -22780 15159 -22746
rect 15197 -22780 15203 -22746
rect 15203 -22780 15231 -22746
rect 15269 -22780 15271 -22746
rect 15271 -22780 15303 -22746
rect 15341 -22780 15373 -22746
rect 15373 -22780 15375 -22746
rect 15413 -22780 15441 -22746
rect 15441 -22780 15447 -22746
rect 15485 -22780 15509 -22746
rect 15509 -22780 15519 -22746
rect 16143 -22780 16153 -22746
rect 16153 -22780 16177 -22746
rect 16215 -22780 16221 -22746
rect 16221 -22780 16249 -22746
rect 16287 -22780 16289 -22746
rect 16289 -22780 16321 -22746
rect 16359 -22780 16391 -22746
rect 16391 -22780 16393 -22746
rect 16431 -22780 16459 -22746
rect 16459 -22780 16465 -22746
rect 16503 -22780 16527 -22746
rect 16527 -22780 16537 -22746
rect 17161 -22780 17171 -22746
rect 17171 -22780 17195 -22746
rect 17233 -22780 17239 -22746
rect 17239 -22780 17267 -22746
rect 17305 -22780 17307 -22746
rect 17307 -22780 17339 -22746
rect 17377 -22780 17409 -22746
rect 17409 -22780 17411 -22746
rect 17449 -22780 17477 -22746
rect 17477 -22780 17483 -22746
rect 17521 -22780 17545 -22746
rect 17545 -22780 17555 -22746
rect 18179 -22780 18189 -22746
rect 18189 -22780 18213 -22746
rect 18251 -22780 18257 -22746
rect 18257 -22780 18285 -22746
rect 18323 -22780 18325 -22746
rect 18325 -22780 18357 -22746
rect 18395 -22780 18427 -22746
rect 18427 -22780 18429 -22746
rect 18467 -22780 18495 -22746
rect 18495 -22780 18501 -22746
rect 18539 -22780 18563 -22746
rect 18563 -22780 18573 -22746
rect 19197 -22780 19207 -22746
rect 19207 -22780 19231 -22746
rect 19269 -22780 19275 -22746
rect 19275 -22780 19303 -22746
rect 19341 -22780 19343 -22746
rect 19343 -22780 19375 -22746
rect 19413 -22780 19445 -22746
rect 19445 -22780 19447 -22746
rect 19485 -22780 19513 -22746
rect 19513 -22780 19519 -22746
rect 19557 -22780 19581 -22746
rect 19581 -22780 19591 -22746
rect 20215 -22780 20225 -22746
rect 20225 -22780 20249 -22746
rect 20287 -22780 20293 -22746
rect 20293 -22780 20321 -22746
rect 20359 -22780 20361 -22746
rect 20361 -22780 20393 -22746
rect 20431 -22780 20463 -22746
rect 20463 -22780 20465 -22746
rect 20503 -22780 20531 -22746
rect 20531 -22780 20537 -22746
rect 20575 -22780 20599 -22746
rect 20599 -22780 20609 -22746
rect 21233 -22780 21243 -22746
rect 21243 -22780 21267 -22746
rect 21305 -22780 21311 -22746
rect 21311 -22780 21339 -22746
rect 21377 -22780 21379 -22746
rect 21379 -22780 21411 -22746
rect 21449 -22780 21481 -22746
rect 21481 -22780 21483 -22746
rect 21521 -22780 21549 -22746
rect 21549 -22780 21555 -22746
rect 21593 -22780 21617 -22746
rect 21617 -22780 21627 -22746
rect 22251 -22780 22261 -22746
rect 22261 -22780 22285 -22746
rect 22323 -22780 22329 -22746
rect 22329 -22780 22357 -22746
rect 22395 -22780 22397 -22746
rect 22397 -22780 22429 -22746
rect 22467 -22780 22499 -22746
rect 22499 -22780 22501 -22746
rect 22539 -22780 22567 -22746
rect 22567 -22780 22573 -22746
rect 22611 -22780 22635 -22746
rect 22635 -22780 22645 -22746
rect 24855 -22753 24889 -22747
rect 24855 -22781 24889 -22753
rect -12289 -22821 -12255 -22819
rect -12289 -22853 -12255 -22821
rect -9077 -22856 -9067 -22822
rect -9067 -22856 -9043 -22822
rect -9005 -22856 -8999 -22822
rect -8999 -22856 -8971 -22822
rect -8933 -22856 -8931 -22822
rect -8931 -22856 -8899 -22822
rect -8861 -22856 -8829 -22822
rect -8829 -22856 -8827 -22822
rect -8789 -22856 -8761 -22822
rect -8761 -22856 -8755 -22822
rect -8717 -22856 -8693 -22822
rect -8693 -22856 -8683 -22822
rect -8059 -22856 -8049 -22822
rect -8049 -22856 -8025 -22822
rect -7987 -22856 -7981 -22822
rect -7981 -22856 -7953 -22822
rect -7915 -22856 -7913 -22822
rect -7913 -22856 -7881 -22822
rect -7843 -22856 -7811 -22822
rect -7811 -22856 -7809 -22822
rect -7771 -22856 -7743 -22822
rect -7743 -22856 -7737 -22822
rect -7699 -22856 -7675 -22822
rect -7675 -22856 -7665 -22822
rect -7041 -22856 -7031 -22822
rect -7031 -22856 -7007 -22822
rect -6969 -22856 -6963 -22822
rect -6963 -22856 -6935 -22822
rect -6897 -22856 -6895 -22822
rect -6895 -22856 -6863 -22822
rect -6825 -22856 -6793 -22822
rect -6793 -22856 -6791 -22822
rect -6753 -22856 -6725 -22822
rect -6725 -22856 -6719 -22822
rect -6681 -22856 -6657 -22822
rect -6657 -22856 -6647 -22822
rect -6023 -22856 -6013 -22822
rect -6013 -22856 -5989 -22822
rect -5951 -22856 -5945 -22822
rect -5945 -22856 -5917 -22822
rect -5879 -22856 -5877 -22822
rect -5877 -22856 -5845 -22822
rect -5807 -22856 -5775 -22822
rect -5775 -22856 -5773 -22822
rect -5735 -22856 -5707 -22822
rect -5707 -22856 -5701 -22822
rect -5663 -22856 -5639 -22822
rect -5639 -22856 -5629 -22822
rect -5005 -22856 -4995 -22822
rect -4995 -22856 -4971 -22822
rect -4933 -22856 -4927 -22822
rect -4927 -22856 -4899 -22822
rect -4861 -22856 -4859 -22822
rect -4859 -22856 -4827 -22822
rect -4789 -22856 -4757 -22822
rect -4757 -22856 -4755 -22822
rect -4717 -22856 -4689 -22822
rect -4689 -22856 -4683 -22822
rect -4645 -22856 -4621 -22822
rect -4621 -22856 -4611 -22822
rect -3987 -22856 -3977 -22822
rect -3977 -22856 -3953 -22822
rect -3915 -22856 -3909 -22822
rect -3909 -22856 -3881 -22822
rect -3843 -22856 -3841 -22822
rect -3841 -22856 -3809 -22822
rect -3771 -22856 -3739 -22822
rect -3739 -22856 -3737 -22822
rect -3699 -22856 -3671 -22822
rect -3671 -22856 -3665 -22822
rect -3627 -22856 -3603 -22822
rect -3603 -22856 -3593 -22822
rect -2261 -22854 -2227 -22820
rect -1963 -22854 -1929 -22820
rect -1665 -22854 -1631 -22820
rect -1367 -22854 -1333 -22820
rect -1069 -22854 -1035 -22820
rect -771 -22854 -737 -22820
rect -473 -22854 -439 -22820
rect -175 -22854 -141 -22820
rect 123 -22854 157 -22820
rect 421 -22854 455 -22820
rect 719 -22854 753 -22820
rect 2580 -22863 2614 -22849
rect 2580 -22883 2614 -22863
rect -12289 -22923 -12255 -22891
rect -12289 -22925 -12255 -22923
rect -12289 -22991 -12255 -22963
rect -12289 -22997 -12255 -22991
rect -12289 -23059 -12255 -23035
rect -12289 -23069 -12255 -23059
rect -12289 -23127 -12255 -23107
rect -12289 -23141 -12255 -23127
rect -12289 -23195 -12255 -23179
rect -12289 -23213 -12255 -23195
rect -12289 -23263 -12255 -23251
rect -12289 -23285 -12255 -23263
rect -12289 -23331 -12255 -23323
rect -12289 -23357 -12255 -23331
rect -12289 -23399 -12255 -23395
rect -12289 -23429 -12255 -23399
rect -12289 -23501 -12255 -23467
rect -9406 -22939 -9372 -22925
rect -9406 -22959 -9372 -22939
rect -9406 -23007 -9372 -22997
rect -9406 -23031 -9372 -23007
rect -9406 -23075 -9372 -23069
rect -9406 -23103 -9372 -23075
rect -9406 -23143 -9372 -23141
rect -9406 -23175 -9372 -23143
rect -9406 -23245 -9372 -23213
rect -9406 -23247 -9372 -23245
rect -9406 -23313 -9372 -23285
rect -9406 -23319 -9372 -23313
rect -9406 -23381 -9372 -23357
rect -9406 -23391 -9372 -23381
rect -9406 -23449 -9372 -23429
rect -9406 -23463 -9372 -23449
rect -8388 -22939 -8354 -22925
rect -8388 -22959 -8354 -22939
rect -8388 -23007 -8354 -22997
rect -8388 -23031 -8354 -23007
rect -8388 -23075 -8354 -23069
rect -8388 -23103 -8354 -23075
rect -8388 -23143 -8354 -23141
rect -8388 -23175 -8354 -23143
rect -8388 -23245 -8354 -23213
rect -8388 -23247 -8354 -23245
rect -8388 -23313 -8354 -23285
rect -8388 -23319 -8354 -23313
rect -8388 -23381 -8354 -23357
rect -8388 -23391 -8354 -23381
rect -8388 -23449 -8354 -23429
rect -8388 -23463 -8354 -23449
rect -7370 -22939 -7336 -22925
rect -7370 -22959 -7336 -22939
rect -7370 -23007 -7336 -22997
rect -7370 -23031 -7336 -23007
rect -7370 -23075 -7336 -23069
rect -7370 -23103 -7336 -23075
rect -7370 -23143 -7336 -23141
rect -7370 -23175 -7336 -23143
rect -7370 -23245 -7336 -23213
rect -7370 -23247 -7336 -23245
rect -7370 -23313 -7336 -23285
rect -7370 -23319 -7336 -23313
rect -7370 -23381 -7336 -23357
rect -7370 -23391 -7336 -23381
rect -7370 -23449 -7336 -23429
rect -7370 -23463 -7336 -23449
rect -6352 -22939 -6318 -22925
rect -6352 -22959 -6318 -22939
rect -6352 -23007 -6318 -22997
rect -6352 -23031 -6318 -23007
rect -6352 -23075 -6318 -23069
rect -6352 -23103 -6318 -23075
rect -6352 -23143 -6318 -23141
rect -6352 -23175 -6318 -23143
rect -6352 -23245 -6318 -23213
rect -6352 -23247 -6318 -23245
rect -6352 -23313 -6318 -23285
rect -6352 -23319 -6318 -23313
rect -6352 -23381 -6318 -23357
rect -6352 -23391 -6318 -23381
rect -6352 -23449 -6318 -23429
rect -6352 -23463 -6318 -23449
rect -5334 -22939 -5300 -22925
rect -5334 -22959 -5300 -22939
rect -5334 -23007 -5300 -22997
rect -5334 -23031 -5300 -23007
rect -5334 -23075 -5300 -23069
rect -5334 -23103 -5300 -23075
rect -5334 -23143 -5300 -23141
rect -5334 -23175 -5300 -23143
rect -5334 -23245 -5300 -23213
rect -5334 -23247 -5300 -23245
rect -5334 -23313 -5300 -23285
rect -5334 -23319 -5300 -23313
rect -5334 -23381 -5300 -23357
rect -5334 -23391 -5300 -23381
rect -5334 -23449 -5300 -23429
rect -5334 -23463 -5300 -23449
rect -4316 -22939 -4282 -22925
rect -4316 -22959 -4282 -22939
rect -4316 -23007 -4282 -22997
rect -4316 -23031 -4282 -23007
rect -4316 -23075 -4282 -23069
rect -4316 -23103 -4282 -23075
rect -4316 -23143 -4282 -23141
rect -4316 -23175 -4282 -23143
rect -4316 -23245 -4282 -23213
rect -4316 -23247 -4282 -23245
rect -4316 -23313 -4282 -23285
rect -4316 -23319 -4282 -23313
rect -4316 -23381 -4282 -23357
rect -4316 -23391 -4282 -23381
rect -4316 -23449 -4282 -23429
rect -4316 -23463 -4282 -23449
rect -3298 -22939 -3264 -22925
rect -3298 -22959 -3264 -22939
rect -3298 -23007 -3264 -22997
rect -3298 -23031 -3264 -23007
rect -3298 -23075 -3264 -23069
rect -3298 -23103 -3264 -23075
rect -3298 -23143 -3264 -23141
rect -3298 -23175 -3264 -23143
rect -3298 -23245 -3264 -23213
rect -3298 -23247 -3264 -23245
rect -3298 -23313 -3264 -23285
rect -3298 -23319 -3264 -23313
rect -3298 -23381 -3264 -23357
rect -3298 -23391 -3264 -23381
rect -3298 -23449 -3264 -23429
rect -3298 -23463 -3264 -23449
rect -2410 -22937 -2376 -22923
rect -2410 -22957 -2376 -22937
rect -2410 -23005 -2376 -22995
rect -2410 -23029 -2376 -23005
rect -2410 -23073 -2376 -23067
rect -2410 -23101 -2376 -23073
rect -2410 -23141 -2376 -23139
rect -2410 -23173 -2376 -23141
rect -2410 -23243 -2376 -23211
rect -2410 -23245 -2376 -23243
rect -2410 -23311 -2376 -23283
rect -2410 -23317 -2376 -23311
rect -2410 -23379 -2376 -23355
rect -2410 -23389 -2376 -23379
rect -2410 -23447 -2376 -23427
rect -2410 -23461 -2376 -23447
rect -2112 -22937 -2078 -22923
rect -2112 -22957 -2078 -22937
rect -2112 -23005 -2078 -22995
rect -2112 -23029 -2078 -23005
rect -2112 -23073 -2078 -23067
rect -2112 -23101 -2078 -23073
rect -2112 -23141 -2078 -23139
rect -2112 -23173 -2078 -23141
rect -2112 -23243 -2078 -23211
rect -2112 -23245 -2078 -23243
rect -2112 -23311 -2078 -23283
rect -2112 -23317 -2078 -23311
rect -2112 -23379 -2078 -23355
rect -2112 -23389 -2078 -23379
rect -2112 -23447 -2078 -23427
rect -2112 -23461 -2078 -23447
rect -1814 -22937 -1780 -22923
rect -1814 -22957 -1780 -22937
rect -1814 -23005 -1780 -22995
rect -1814 -23029 -1780 -23005
rect -1814 -23073 -1780 -23067
rect -1814 -23101 -1780 -23073
rect -1814 -23141 -1780 -23139
rect -1814 -23173 -1780 -23141
rect -1814 -23243 -1780 -23211
rect -1814 -23245 -1780 -23243
rect -1814 -23311 -1780 -23283
rect -1814 -23317 -1780 -23311
rect -1814 -23379 -1780 -23355
rect -1814 -23389 -1780 -23379
rect -1814 -23447 -1780 -23427
rect -1814 -23461 -1780 -23447
rect -1516 -22937 -1482 -22923
rect -1516 -22957 -1482 -22937
rect -1516 -23005 -1482 -22995
rect -1516 -23029 -1482 -23005
rect -1516 -23073 -1482 -23067
rect -1516 -23101 -1482 -23073
rect -1516 -23141 -1482 -23139
rect -1516 -23173 -1482 -23141
rect -1516 -23243 -1482 -23211
rect -1516 -23245 -1482 -23243
rect -1516 -23311 -1482 -23283
rect -1516 -23317 -1482 -23311
rect -1516 -23379 -1482 -23355
rect -1516 -23389 -1482 -23379
rect -1516 -23447 -1482 -23427
rect -1516 -23461 -1482 -23447
rect -1218 -22937 -1184 -22923
rect -1218 -22957 -1184 -22937
rect -1218 -23005 -1184 -22995
rect -1218 -23029 -1184 -23005
rect -1218 -23073 -1184 -23067
rect -1218 -23101 -1184 -23073
rect -1218 -23141 -1184 -23139
rect -1218 -23173 -1184 -23141
rect -1218 -23243 -1184 -23211
rect -1218 -23245 -1184 -23243
rect -1218 -23311 -1184 -23283
rect -1218 -23317 -1184 -23311
rect -1218 -23379 -1184 -23355
rect -1218 -23389 -1184 -23379
rect -1218 -23447 -1184 -23427
rect -1218 -23461 -1184 -23447
rect -920 -22937 -886 -22923
rect -920 -22957 -886 -22937
rect -920 -23005 -886 -22995
rect -920 -23029 -886 -23005
rect -920 -23073 -886 -23067
rect -920 -23101 -886 -23073
rect -920 -23141 -886 -23139
rect -920 -23173 -886 -23141
rect -920 -23243 -886 -23211
rect -920 -23245 -886 -23243
rect -920 -23311 -886 -23283
rect -920 -23317 -886 -23311
rect -920 -23379 -886 -23355
rect -920 -23389 -886 -23379
rect -920 -23447 -886 -23427
rect -920 -23461 -886 -23447
rect -622 -22937 -588 -22923
rect -622 -22957 -588 -22937
rect -622 -23005 -588 -22995
rect -622 -23029 -588 -23005
rect -622 -23073 -588 -23067
rect -622 -23101 -588 -23073
rect -622 -23141 -588 -23139
rect -622 -23173 -588 -23141
rect -622 -23243 -588 -23211
rect -622 -23245 -588 -23243
rect -622 -23311 -588 -23283
rect -622 -23317 -588 -23311
rect -622 -23379 -588 -23355
rect -622 -23389 -588 -23379
rect -622 -23447 -588 -23427
rect -622 -23461 -588 -23447
rect -324 -22937 -290 -22923
rect -324 -22957 -290 -22937
rect -324 -23005 -290 -22995
rect -324 -23029 -290 -23005
rect -324 -23073 -290 -23067
rect -324 -23101 -290 -23073
rect -324 -23141 -290 -23139
rect -324 -23173 -290 -23141
rect -324 -23243 -290 -23211
rect -324 -23245 -290 -23243
rect -324 -23311 -290 -23283
rect -324 -23317 -290 -23311
rect -324 -23379 -290 -23355
rect -324 -23389 -290 -23379
rect -324 -23447 -290 -23427
rect -324 -23461 -290 -23447
rect -26 -22937 8 -22923
rect -26 -22957 8 -22937
rect -26 -23005 8 -22995
rect -26 -23029 8 -23005
rect -26 -23073 8 -23067
rect -26 -23101 8 -23073
rect -26 -23141 8 -23139
rect -26 -23173 8 -23141
rect -26 -23243 8 -23211
rect -26 -23245 8 -23243
rect -26 -23311 8 -23283
rect -26 -23317 8 -23311
rect -26 -23379 8 -23355
rect -26 -23389 8 -23379
rect -26 -23447 8 -23427
rect -26 -23461 8 -23447
rect 272 -22937 306 -22923
rect 272 -22957 306 -22937
rect 272 -23005 306 -22995
rect 272 -23029 306 -23005
rect 272 -23073 306 -23067
rect 272 -23101 306 -23073
rect 272 -23141 306 -23139
rect 272 -23173 306 -23141
rect 272 -23243 306 -23211
rect 272 -23245 306 -23243
rect 272 -23311 306 -23283
rect 272 -23317 306 -23311
rect 272 -23379 306 -23355
rect 272 -23389 306 -23379
rect 272 -23447 306 -23427
rect 272 -23461 306 -23447
rect 570 -22937 604 -22923
rect 570 -22957 604 -22937
rect 570 -23005 604 -22995
rect 570 -23029 604 -23005
rect 570 -23073 604 -23067
rect 570 -23101 604 -23073
rect 570 -23141 604 -23139
rect 570 -23173 604 -23141
rect 570 -23243 604 -23211
rect 570 -23245 604 -23243
rect 570 -23311 604 -23283
rect 570 -23317 604 -23311
rect 570 -23379 604 -23355
rect 570 -23389 604 -23379
rect 570 -23447 604 -23427
rect 570 -23461 604 -23447
rect 868 -22937 902 -22923
rect 868 -22957 902 -22937
rect 868 -23005 902 -22995
rect 868 -23029 902 -23005
rect 868 -23073 902 -23067
rect 868 -23101 902 -23073
rect 868 -23141 902 -23139
rect 868 -23173 902 -23141
rect 868 -23243 902 -23211
rect 868 -23245 902 -23243
rect 868 -23311 902 -23283
rect 868 -23317 902 -23311
rect 868 -23379 902 -23355
rect 868 -23389 902 -23379
rect 2580 -22931 2614 -22921
rect 2580 -22955 2614 -22931
rect 2580 -22999 2614 -22993
rect 2580 -23027 2614 -22999
rect 2580 -23067 2614 -23065
rect 2580 -23099 2614 -23067
rect 2580 -23169 2614 -23137
rect 2580 -23171 2614 -23169
rect 2580 -23237 2614 -23209
rect 2580 -23243 2614 -23237
rect 2580 -23305 2614 -23281
rect 2580 -23315 2614 -23305
rect 2580 -23373 2614 -23353
rect 2580 -23387 2614 -23373
rect 3598 -22863 3632 -22849
rect 3598 -22883 3632 -22863
rect 3598 -22931 3632 -22921
rect 3598 -22955 3632 -22931
rect 3598 -22999 3632 -22993
rect 3598 -23027 3632 -22999
rect 3598 -23067 3632 -23065
rect 3598 -23099 3632 -23067
rect 3598 -23169 3632 -23137
rect 3598 -23171 3632 -23169
rect 3598 -23237 3632 -23209
rect 3598 -23243 3632 -23237
rect 3598 -23305 3632 -23281
rect 3598 -23315 3632 -23305
rect 3598 -23373 3632 -23353
rect 3598 -23387 3632 -23373
rect 4616 -22863 4650 -22849
rect 4616 -22883 4650 -22863
rect 4616 -22931 4650 -22921
rect 4616 -22955 4650 -22931
rect 4616 -22999 4650 -22993
rect 4616 -23027 4650 -22999
rect 4616 -23067 4650 -23065
rect 4616 -23099 4650 -23067
rect 4616 -23169 4650 -23137
rect 4616 -23171 4650 -23169
rect 4616 -23237 4650 -23209
rect 4616 -23243 4650 -23237
rect 4616 -23305 4650 -23281
rect 4616 -23315 4650 -23305
rect 4616 -23373 4650 -23353
rect 4616 -23387 4650 -23373
rect 5634 -22863 5668 -22849
rect 5634 -22883 5668 -22863
rect 5634 -22931 5668 -22921
rect 5634 -22955 5668 -22931
rect 5634 -22999 5668 -22993
rect 5634 -23027 5668 -22999
rect 5634 -23067 5668 -23065
rect 5634 -23099 5668 -23067
rect 5634 -23169 5668 -23137
rect 5634 -23171 5668 -23169
rect 5634 -23237 5668 -23209
rect 5634 -23243 5668 -23237
rect 5634 -23305 5668 -23281
rect 5634 -23315 5668 -23305
rect 5634 -23373 5668 -23353
rect 5634 -23387 5668 -23373
rect 6652 -22863 6686 -22849
rect 6652 -22883 6686 -22863
rect 6652 -22931 6686 -22921
rect 6652 -22955 6686 -22931
rect 6652 -22999 6686 -22993
rect 6652 -23027 6686 -22999
rect 6652 -23067 6686 -23065
rect 6652 -23099 6686 -23067
rect 6652 -23169 6686 -23137
rect 6652 -23171 6686 -23169
rect 6652 -23237 6686 -23209
rect 6652 -23243 6686 -23237
rect 6652 -23305 6686 -23281
rect 6652 -23315 6686 -23305
rect 6652 -23373 6686 -23353
rect 6652 -23387 6686 -23373
rect 7670 -22863 7704 -22849
rect 7670 -22883 7704 -22863
rect 7670 -22931 7704 -22921
rect 7670 -22955 7704 -22931
rect 7670 -22999 7704 -22993
rect 7670 -23027 7704 -22999
rect 7670 -23067 7704 -23065
rect 7670 -23099 7704 -23067
rect 7670 -23169 7704 -23137
rect 7670 -23171 7704 -23169
rect 7670 -23237 7704 -23209
rect 7670 -23243 7704 -23237
rect 7670 -23305 7704 -23281
rect 7670 -23315 7704 -23305
rect 7670 -23373 7704 -23353
rect 7670 -23387 7704 -23373
rect 8688 -22863 8722 -22849
rect 8688 -22883 8722 -22863
rect 8688 -22931 8722 -22921
rect 8688 -22955 8722 -22931
rect 8688 -22999 8722 -22993
rect 8688 -23027 8722 -22999
rect 8688 -23067 8722 -23065
rect 8688 -23099 8722 -23067
rect 8688 -23169 8722 -23137
rect 8688 -23171 8722 -23169
rect 8688 -23237 8722 -23209
rect 8688 -23243 8722 -23237
rect 8688 -23305 8722 -23281
rect 8688 -23315 8722 -23305
rect 8688 -23373 8722 -23353
rect 8688 -23387 8722 -23373
rect 9706 -22863 9740 -22849
rect 9706 -22883 9740 -22863
rect 9706 -22931 9740 -22921
rect 9706 -22955 9740 -22931
rect 9706 -22999 9740 -22993
rect 9706 -23027 9740 -22999
rect 9706 -23067 9740 -23065
rect 9706 -23099 9740 -23067
rect 9706 -23169 9740 -23137
rect 9706 -23171 9740 -23169
rect 9706 -23237 9740 -23209
rect 9706 -23243 9740 -23237
rect 9706 -23305 9740 -23281
rect 9706 -23315 9740 -23305
rect 9706 -23373 9740 -23353
rect 9706 -23387 9740 -23373
rect 10724 -22863 10758 -22849
rect 10724 -22883 10758 -22863
rect 10724 -22931 10758 -22921
rect 10724 -22955 10758 -22931
rect 10724 -22999 10758 -22993
rect 10724 -23027 10758 -22999
rect 10724 -23067 10758 -23065
rect 10724 -23099 10758 -23067
rect 10724 -23169 10758 -23137
rect 10724 -23171 10758 -23169
rect 10724 -23237 10758 -23209
rect 10724 -23243 10758 -23237
rect 10724 -23305 10758 -23281
rect 10724 -23315 10758 -23305
rect 10724 -23373 10758 -23353
rect 10724 -23387 10758 -23373
rect 11742 -22863 11776 -22849
rect 11742 -22883 11776 -22863
rect 11742 -22931 11776 -22921
rect 11742 -22955 11776 -22931
rect 11742 -22999 11776 -22993
rect 11742 -23027 11776 -22999
rect 11742 -23067 11776 -23065
rect 11742 -23099 11776 -23067
rect 11742 -23169 11776 -23137
rect 11742 -23171 11776 -23169
rect 11742 -23237 11776 -23209
rect 11742 -23243 11776 -23237
rect 11742 -23305 11776 -23281
rect 11742 -23315 11776 -23305
rect 11742 -23373 11776 -23353
rect 11742 -23387 11776 -23373
rect 12760 -22863 12794 -22849
rect 12760 -22883 12794 -22863
rect 12760 -22931 12794 -22921
rect 12760 -22955 12794 -22931
rect 12760 -22999 12794 -22993
rect 12760 -23027 12794 -22999
rect 12760 -23067 12794 -23065
rect 12760 -23099 12794 -23067
rect 12760 -23169 12794 -23137
rect 12760 -23171 12794 -23169
rect 12760 -23237 12794 -23209
rect 12760 -23243 12794 -23237
rect 12760 -23305 12794 -23281
rect 12760 -23315 12794 -23305
rect 12760 -23373 12794 -23353
rect 12760 -23387 12794 -23373
rect 13778 -22863 13812 -22849
rect 13778 -22883 13812 -22863
rect 13778 -22931 13812 -22921
rect 13778 -22955 13812 -22931
rect 13778 -22999 13812 -22993
rect 13778 -23027 13812 -22999
rect 13778 -23067 13812 -23065
rect 13778 -23099 13812 -23067
rect 13778 -23169 13812 -23137
rect 13778 -23171 13812 -23169
rect 13778 -23237 13812 -23209
rect 13778 -23243 13812 -23237
rect 13778 -23305 13812 -23281
rect 13778 -23315 13812 -23305
rect 13778 -23373 13812 -23353
rect 13778 -23387 13812 -23373
rect 14796 -22863 14830 -22849
rect 14796 -22883 14830 -22863
rect 14796 -22931 14830 -22921
rect 14796 -22955 14830 -22931
rect 14796 -22999 14830 -22993
rect 14796 -23027 14830 -22999
rect 14796 -23067 14830 -23065
rect 14796 -23099 14830 -23067
rect 14796 -23169 14830 -23137
rect 14796 -23171 14830 -23169
rect 14796 -23237 14830 -23209
rect 14796 -23243 14830 -23237
rect 14796 -23305 14830 -23281
rect 14796 -23315 14830 -23305
rect 14796 -23373 14830 -23353
rect 14796 -23387 14830 -23373
rect 15814 -22863 15848 -22849
rect 15814 -22883 15848 -22863
rect 15814 -22931 15848 -22921
rect 15814 -22955 15848 -22931
rect 15814 -22999 15848 -22993
rect 15814 -23027 15848 -22999
rect 15814 -23067 15848 -23065
rect 15814 -23099 15848 -23067
rect 15814 -23169 15848 -23137
rect 15814 -23171 15848 -23169
rect 15814 -23237 15848 -23209
rect 15814 -23243 15848 -23237
rect 15814 -23305 15848 -23281
rect 15814 -23315 15848 -23305
rect 15814 -23373 15848 -23353
rect 15814 -23387 15848 -23373
rect 16832 -22863 16866 -22849
rect 16832 -22883 16866 -22863
rect 16832 -22931 16866 -22921
rect 16832 -22955 16866 -22931
rect 16832 -22999 16866 -22993
rect 16832 -23027 16866 -22999
rect 16832 -23067 16866 -23065
rect 16832 -23099 16866 -23067
rect 16832 -23169 16866 -23137
rect 16832 -23171 16866 -23169
rect 16832 -23237 16866 -23209
rect 16832 -23243 16866 -23237
rect 16832 -23305 16866 -23281
rect 16832 -23315 16866 -23305
rect 16832 -23373 16866 -23353
rect 16832 -23387 16866 -23373
rect 17850 -22863 17884 -22849
rect 17850 -22883 17884 -22863
rect 17850 -22931 17884 -22921
rect 17850 -22955 17884 -22931
rect 17850 -22999 17884 -22993
rect 17850 -23027 17884 -22999
rect 17850 -23067 17884 -23065
rect 17850 -23099 17884 -23067
rect 17850 -23169 17884 -23137
rect 17850 -23171 17884 -23169
rect 17850 -23237 17884 -23209
rect 17850 -23243 17884 -23237
rect 17850 -23305 17884 -23281
rect 17850 -23315 17884 -23305
rect 17850 -23373 17884 -23353
rect 17850 -23387 17884 -23373
rect 18868 -22863 18902 -22849
rect 18868 -22883 18902 -22863
rect 18868 -22931 18902 -22921
rect 18868 -22955 18902 -22931
rect 18868 -22999 18902 -22993
rect 18868 -23027 18902 -22999
rect 18868 -23067 18902 -23065
rect 18868 -23099 18902 -23067
rect 18868 -23169 18902 -23137
rect 18868 -23171 18902 -23169
rect 18868 -23237 18902 -23209
rect 18868 -23243 18902 -23237
rect 18868 -23305 18902 -23281
rect 18868 -23315 18902 -23305
rect 18868 -23373 18902 -23353
rect 18868 -23387 18902 -23373
rect 19886 -22863 19920 -22849
rect 19886 -22883 19920 -22863
rect 19886 -22931 19920 -22921
rect 19886 -22955 19920 -22931
rect 19886 -22999 19920 -22993
rect 19886 -23027 19920 -22999
rect 19886 -23067 19920 -23065
rect 19886 -23099 19920 -23067
rect 19886 -23169 19920 -23137
rect 19886 -23171 19920 -23169
rect 19886 -23237 19920 -23209
rect 19886 -23243 19920 -23237
rect 19886 -23305 19920 -23281
rect 19886 -23315 19920 -23305
rect 19886 -23373 19920 -23353
rect 19886 -23387 19920 -23373
rect 20904 -22863 20938 -22849
rect 20904 -22883 20938 -22863
rect 20904 -22931 20938 -22921
rect 20904 -22955 20938 -22931
rect 20904 -22999 20938 -22993
rect 20904 -23027 20938 -22999
rect 20904 -23067 20938 -23065
rect 20904 -23099 20938 -23067
rect 20904 -23169 20938 -23137
rect 20904 -23171 20938 -23169
rect 20904 -23237 20938 -23209
rect 20904 -23243 20938 -23237
rect 20904 -23305 20938 -23281
rect 20904 -23315 20938 -23305
rect 20904 -23373 20938 -23353
rect 20904 -23387 20938 -23373
rect 21922 -22863 21956 -22849
rect 21922 -22883 21956 -22863
rect 21922 -22931 21956 -22921
rect 21922 -22955 21956 -22931
rect 21922 -22999 21956 -22993
rect 21922 -23027 21956 -22999
rect 21922 -23067 21956 -23065
rect 21922 -23099 21956 -23067
rect 21922 -23169 21956 -23137
rect 21922 -23171 21956 -23169
rect 21922 -23237 21956 -23209
rect 21922 -23243 21956 -23237
rect 21922 -23305 21956 -23281
rect 21922 -23315 21956 -23305
rect 21922 -23373 21956 -23353
rect 21922 -23387 21956 -23373
rect 22940 -22863 22974 -22849
rect 22940 -22883 22974 -22863
rect 22940 -22931 22974 -22921
rect 22940 -22955 22974 -22931
rect 22940 -22999 22974 -22993
rect 22940 -23027 22974 -22999
rect 22940 -23067 22974 -23065
rect 22940 -23099 22974 -23067
rect 22940 -23169 22974 -23137
rect 22940 -23171 22974 -23169
rect 22940 -23237 22974 -23209
rect 22940 -23243 22974 -23237
rect 22940 -23305 22974 -23281
rect 22940 -23315 22974 -23305
rect 22940 -23373 22974 -23353
rect 22940 -23387 22974 -23373
rect 24855 -22821 24889 -22819
rect 24855 -22853 24889 -22821
rect 24855 -22923 24889 -22891
rect 24855 -22925 24889 -22923
rect 24855 -22991 24889 -22963
rect 24855 -22997 24889 -22991
rect 24855 -23059 24889 -23035
rect 24855 -23069 24889 -23059
rect 24855 -23127 24889 -23107
rect 24855 -23141 24889 -23127
rect 24855 -23195 24889 -23179
rect 24855 -23213 24889 -23195
rect 24855 -23263 24889 -23251
rect 24855 -23285 24889 -23263
rect 24855 -23331 24889 -23323
rect 24855 -23357 24889 -23331
rect 868 -23447 902 -23427
rect 868 -23461 902 -23447
rect 24855 -23399 24889 -23395
rect 24855 -23429 24889 -23399
rect 2909 -23490 2919 -23456
rect 2919 -23490 2943 -23456
rect 2981 -23490 2987 -23456
rect 2987 -23490 3015 -23456
rect 3053 -23490 3055 -23456
rect 3055 -23490 3087 -23456
rect 3125 -23490 3157 -23456
rect 3157 -23490 3159 -23456
rect 3197 -23490 3225 -23456
rect 3225 -23490 3231 -23456
rect 3269 -23490 3293 -23456
rect 3293 -23490 3303 -23456
rect 3927 -23490 3937 -23456
rect 3937 -23490 3961 -23456
rect 3999 -23490 4005 -23456
rect 4005 -23490 4033 -23456
rect 4071 -23490 4073 -23456
rect 4073 -23490 4105 -23456
rect 4143 -23490 4175 -23456
rect 4175 -23490 4177 -23456
rect 4215 -23490 4243 -23456
rect 4243 -23490 4249 -23456
rect 4287 -23490 4311 -23456
rect 4311 -23490 4321 -23456
rect 4945 -23490 4955 -23456
rect 4955 -23490 4979 -23456
rect 5017 -23490 5023 -23456
rect 5023 -23490 5051 -23456
rect 5089 -23490 5091 -23456
rect 5091 -23490 5123 -23456
rect 5161 -23490 5193 -23456
rect 5193 -23490 5195 -23456
rect 5233 -23490 5261 -23456
rect 5261 -23490 5267 -23456
rect 5305 -23490 5329 -23456
rect 5329 -23490 5339 -23456
rect 5963 -23490 5973 -23456
rect 5973 -23490 5997 -23456
rect 6035 -23490 6041 -23456
rect 6041 -23490 6069 -23456
rect 6107 -23490 6109 -23456
rect 6109 -23490 6141 -23456
rect 6179 -23490 6211 -23456
rect 6211 -23490 6213 -23456
rect 6251 -23490 6279 -23456
rect 6279 -23490 6285 -23456
rect 6323 -23490 6347 -23456
rect 6347 -23490 6357 -23456
rect 6981 -23490 6991 -23456
rect 6991 -23490 7015 -23456
rect 7053 -23490 7059 -23456
rect 7059 -23490 7087 -23456
rect 7125 -23490 7127 -23456
rect 7127 -23490 7159 -23456
rect 7197 -23490 7229 -23456
rect 7229 -23490 7231 -23456
rect 7269 -23490 7297 -23456
rect 7297 -23490 7303 -23456
rect 7341 -23490 7365 -23456
rect 7365 -23490 7375 -23456
rect 7999 -23490 8009 -23456
rect 8009 -23490 8033 -23456
rect 8071 -23490 8077 -23456
rect 8077 -23490 8105 -23456
rect 8143 -23490 8145 -23456
rect 8145 -23490 8177 -23456
rect 8215 -23490 8247 -23456
rect 8247 -23490 8249 -23456
rect 8287 -23490 8315 -23456
rect 8315 -23490 8321 -23456
rect 8359 -23490 8383 -23456
rect 8383 -23490 8393 -23456
rect 9017 -23490 9027 -23456
rect 9027 -23490 9051 -23456
rect 9089 -23490 9095 -23456
rect 9095 -23490 9123 -23456
rect 9161 -23490 9163 -23456
rect 9163 -23490 9195 -23456
rect 9233 -23490 9265 -23456
rect 9265 -23490 9267 -23456
rect 9305 -23490 9333 -23456
rect 9333 -23490 9339 -23456
rect 9377 -23490 9401 -23456
rect 9401 -23490 9411 -23456
rect 10035 -23490 10045 -23456
rect 10045 -23490 10069 -23456
rect 10107 -23490 10113 -23456
rect 10113 -23490 10141 -23456
rect 10179 -23490 10181 -23456
rect 10181 -23490 10213 -23456
rect 10251 -23490 10283 -23456
rect 10283 -23490 10285 -23456
rect 10323 -23490 10351 -23456
rect 10351 -23490 10357 -23456
rect 10395 -23490 10419 -23456
rect 10419 -23490 10429 -23456
rect 11053 -23490 11063 -23456
rect 11063 -23490 11087 -23456
rect 11125 -23490 11131 -23456
rect 11131 -23490 11159 -23456
rect 11197 -23490 11199 -23456
rect 11199 -23490 11231 -23456
rect 11269 -23490 11301 -23456
rect 11301 -23490 11303 -23456
rect 11341 -23490 11369 -23456
rect 11369 -23490 11375 -23456
rect 11413 -23490 11437 -23456
rect 11437 -23490 11447 -23456
rect 12071 -23490 12081 -23456
rect 12081 -23490 12105 -23456
rect 12143 -23490 12149 -23456
rect 12149 -23490 12177 -23456
rect 12215 -23490 12217 -23456
rect 12217 -23490 12249 -23456
rect 12287 -23490 12319 -23456
rect 12319 -23490 12321 -23456
rect 12359 -23490 12387 -23456
rect 12387 -23490 12393 -23456
rect 12431 -23490 12455 -23456
rect 12455 -23490 12465 -23456
rect 13089 -23490 13099 -23456
rect 13099 -23490 13123 -23456
rect 13161 -23490 13167 -23456
rect 13167 -23490 13195 -23456
rect 13233 -23490 13235 -23456
rect 13235 -23490 13267 -23456
rect 13305 -23490 13337 -23456
rect 13337 -23490 13339 -23456
rect 13377 -23490 13405 -23456
rect 13405 -23490 13411 -23456
rect 13449 -23490 13473 -23456
rect 13473 -23490 13483 -23456
rect 14107 -23490 14117 -23456
rect 14117 -23490 14141 -23456
rect 14179 -23490 14185 -23456
rect 14185 -23490 14213 -23456
rect 14251 -23490 14253 -23456
rect 14253 -23490 14285 -23456
rect 14323 -23490 14355 -23456
rect 14355 -23490 14357 -23456
rect 14395 -23490 14423 -23456
rect 14423 -23490 14429 -23456
rect 14467 -23490 14491 -23456
rect 14491 -23490 14501 -23456
rect 15125 -23490 15135 -23456
rect 15135 -23490 15159 -23456
rect 15197 -23490 15203 -23456
rect 15203 -23490 15231 -23456
rect 15269 -23490 15271 -23456
rect 15271 -23490 15303 -23456
rect 15341 -23490 15373 -23456
rect 15373 -23490 15375 -23456
rect 15413 -23490 15441 -23456
rect 15441 -23490 15447 -23456
rect 15485 -23490 15509 -23456
rect 15509 -23490 15519 -23456
rect 16143 -23490 16153 -23456
rect 16153 -23490 16177 -23456
rect 16215 -23490 16221 -23456
rect 16221 -23490 16249 -23456
rect 16287 -23490 16289 -23456
rect 16289 -23490 16321 -23456
rect 16359 -23490 16391 -23456
rect 16391 -23490 16393 -23456
rect 16431 -23490 16459 -23456
rect 16459 -23490 16465 -23456
rect 16503 -23490 16527 -23456
rect 16527 -23490 16537 -23456
rect 17161 -23490 17171 -23456
rect 17171 -23490 17195 -23456
rect 17233 -23490 17239 -23456
rect 17239 -23490 17267 -23456
rect 17305 -23490 17307 -23456
rect 17307 -23490 17339 -23456
rect 17377 -23490 17409 -23456
rect 17409 -23490 17411 -23456
rect 17449 -23490 17477 -23456
rect 17477 -23490 17483 -23456
rect 17521 -23490 17545 -23456
rect 17545 -23490 17555 -23456
rect 18179 -23490 18189 -23456
rect 18189 -23490 18213 -23456
rect 18251 -23490 18257 -23456
rect 18257 -23490 18285 -23456
rect 18323 -23490 18325 -23456
rect 18325 -23490 18357 -23456
rect 18395 -23490 18427 -23456
rect 18427 -23490 18429 -23456
rect 18467 -23490 18495 -23456
rect 18495 -23490 18501 -23456
rect 18539 -23490 18563 -23456
rect 18563 -23490 18573 -23456
rect 19197 -23490 19207 -23456
rect 19207 -23490 19231 -23456
rect 19269 -23490 19275 -23456
rect 19275 -23490 19303 -23456
rect 19341 -23490 19343 -23456
rect 19343 -23490 19375 -23456
rect 19413 -23490 19445 -23456
rect 19445 -23490 19447 -23456
rect 19485 -23490 19513 -23456
rect 19513 -23490 19519 -23456
rect 19557 -23490 19581 -23456
rect 19581 -23490 19591 -23456
rect 20215 -23490 20225 -23456
rect 20225 -23490 20249 -23456
rect 20287 -23490 20293 -23456
rect 20293 -23490 20321 -23456
rect 20359 -23490 20361 -23456
rect 20361 -23490 20393 -23456
rect 20431 -23490 20463 -23456
rect 20463 -23490 20465 -23456
rect 20503 -23490 20531 -23456
rect 20531 -23490 20537 -23456
rect 20575 -23490 20599 -23456
rect 20599 -23490 20609 -23456
rect 21233 -23490 21243 -23456
rect 21243 -23490 21267 -23456
rect 21305 -23490 21311 -23456
rect 21311 -23490 21339 -23456
rect 21377 -23490 21379 -23456
rect 21379 -23490 21411 -23456
rect 21449 -23490 21481 -23456
rect 21481 -23490 21483 -23456
rect 21521 -23490 21549 -23456
rect 21549 -23490 21555 -23456
rect 21593 -23490 21617 -23456
rect 21617 -23490 21627 -23456
rect 22251 -23490 22261 -23456
rect 22261 -23490 22285 -23456
rect 22323 -23490 22329 -23456
rect 22329 -23490 22357 -23456
rect 22395 -23490 22397 -23456
rect 22397 -23490 22429 -23456
rect 22467 -23490 22499 -23456
rect 22499 -23490 22501 -23456
rect 22539 -23490 22567 -23456
rect 22567 -23490 22573 -23456
rect 22611 -23490 22635 -23456
rect 22635 -23490 22645 -23456
rect 24855 -23501 24889 -23467
rect -12289 -23569 -12255 -23539
rect -12289 -23573 -12255 -23569
rect -9077 -23566 -9067 -23532
rect -9067 -23566 -9043 -23532
rect -9005 -23566 -8999 -23532
rect -8999 -23566 -8971 -23532
rect -8933 -23566 -8931 -23532
rect -8931 -23566 -8899 -23532
rect -8861 -23566 -8829 -23532
rect -8829 -23566 -8827 -23532
rect -8789 -23566 -8761 -23532
rect -8761 -23566 -8755 -23532
rect -8717 -23566 -8693 -23532
rect -8693 -23566 -8683 -23532
rect -8059 -23566 -8049 -23532
rect -8049 -23566 -8025 -23532
rect -7987 -23566 -7981 -23532
rect -7981 -23566 -7953 -23532
rect -7915 -23566 -7913 -23532
rect -7913 -23566 -7881 -23532
rect -7843 -23566 -7811 -23532
rect -7811 -23566 -7809 -23532
rect -7771 -23566 -7743 -23532
rect -7743 -23566 -7737 -23532
rect -7699 -23566 -7675 -23532
rect -7675 -23566 -7665 -23532
rect -7041 -23566 -7031 -23532
rect -7031 -23566 -7007 -23532
rect -6969 -23566 -6963 -23532
rect -6963 -23566 -6935 -23532
rect -6897 -23566 -6895 -23532
rect -6895 -23566 -6863 -23532
rect -6825 -23566 -6793 -23532
rect -6793 -23566 -6791 -23532
rect -6753 -23566 -6725 -23532
rect -6725 -23566 -6719 -23532
rect -6681 -23566 -6657 -23532
rect -6657 -23566 -6647 -23532
rect -6023 -23566 -6013 -23532
rect -6013 -23566 -5989 -23532
rect -5951 -23566 -5945 -23532
rect -5945 -23566 -5917 -23532
rect -5879 -23566 -5877 -23532
rect -5877 -23566 -5845 -23532
rect -5807 -23566 -5775 -23532
rect -5775 -23566 -5773 -23532
rect -5735 -23566 -5707 -23532
rect -5707 -23566 -5701 -23532
rect -5663 -23566 -5639 -23532
rect -5639 -23566 -5629 -23532
rect -5005 -23566 -4995 -23532
rect -4995 -23566 -4971 -23532
rect -4933 -23566 -4927 -23532
rect -4927 -23566 -4899 -23532
rect -4861 -23566 -4859 -23532
rect -4859 -23566 -4827 -23532
rect -4789 -23566 -4757 -23532
rect -4757 -23566 -4755 -23532
rect -4717 -23566 -4689 -23532
rect -4689 -23566 -4683 -23532
rect -4645 -23566 -4621 -23532
rect -4621 -23566 -4611 -23532
rect -3987 -23566 -3977 -23532
rect -3977 -23566 -3953 -23532
rect -3915 -23566 -3909 -23532
rect -3909 -23566 -3881 -23532
rect -3843 -23566 -3841 -23532
rect -3841 -23566 -3809 -23532
rect -3771 -23566 -3739 -23532
rect -3739 -23566 -3737 -23532
rect -3699 -23566 -3671 -23532
rect -3671 -23566 -3665 -23532
rect -3627 -23566 -3603 -23532
rect -3603 -23566 -3593 -23532
rect -2261 -23564 -2227 -23530
rect -1963 -23564 -1929 -23530
rect -1665 -23564 -1631 -23530
rect -1367 -23564 -1333 -23530
rect -1069 -23564 -1035 -23530
rect -771 -23564 -737 -23530
rect -473 -23564 -439 -23530
rect -175 -23564 -141 -23530
rect 123 -23564 157 -23530
rect 421 -23564 455 -23530
rect 719 -23564 753 -23530
rect -12289 -23637 -12255 -23611
rect -12289 -23645 -12255 -23637
rect -12289 -23705 -12255 -23683
rect -12289 -23717 -12255 -23705
rect -12289 -23773 -12255 -23755
rect -12289 -23789 -12255 -23773
rect -12289 -23841 -12255 -23827
rect -12289 -23861 -12255 -23841
rect -12289 -23909 -12255 -23899
rect -12289 -23933 -12255 -23909
rect 24855 -23569 24889 -23539
rect 24855 -23573 24889 -23569
rect 24855 -23637 24889 -23611
rect 24855 -23645 24889 -23637
rect 24855 -23705 24889 -23683
rect 24855 -23717 24889 -23705
rect 24855 -23773 24889 -23755
rect 24855 -23789 24889 -23773
rect 24855 -23841 24889 -23827
rect 24855 -23861 24889 -23841
rect -12289 -23977 -12255 -23971
rect -12289 -24005 -12255 -23977
rect -9076 -23967 -9066 -23933
rect -9066 -23967 -9042 -23933
rect -9004 -23967 -8998 -23933
rect -8998 -23967 -8970 -23933
rect -8932 -23967 -8930 -23933
rect -8930 -23967 -8898 -23933
rect -8860 -23967 -8828 -23933
rect -8828 -23967 -8826 -23933
rect -8788 -23967 -8760 -23933
rect -8760 -23967 -8754 -23933
rect -8716 -23967 -8692 -23933
rect -8692 -23967 -8682 -23933
rect -8058 -23967 -8048 -23933
rect -8048 -23967 -8024 -23933
rect -7986 -23967 -7980 -23933
rect -7980 -23967 -7952 -23933
rect -7914 -23967 -7912 -23933
rect -7912 -23967 -7880 -23933
rect -7842 -23967 -7810 -23933
rect -7810 -23967 -7808 -23933
rect -7770 -23967 -7742 -23933
rect -7742 -23967 -7736 -23933
rect -7698 -23967 -7674 -23933
rect -7674 -23967 -7664 -23933
rect -7040 -23967 -7030 -23933
rect -7030 -23967 -7006 -23933
rect -6968 -23967 -6962 -23933
rect -6962 -23967 -6934 -23933
rect -6896 -23967 -6894 -23933
rect -6894 -23967 -6862 -23933
rect -6824 -23967 -6792 -23933
rect -6792 -23967 -6790 -23933
rect -6752 -23967 -6724 -23933
rect -6724 -23967 -6718 -23933
rect -6680 -23967 -6656 -23933
rect -6656 -23967 -6646 -23933
rect -6022 -23967 -6012 -23933
rect -6012 -23967 -5988 -23933
rect -5950 -23967 -5944 -23933
rect -5944 -23967 -5916 -23933
rect -5878 -23967 -5876 -23933
rect -5876 -23967 -5844 -23933
rect -5806 -23967 -5774 -23933
rect -5774 -23967 -5772 -23933
rect -5734 -23967 -5706 -23933
rect -5706 -23967 -5700 -23933
rect -5662 -23967 -5638 -23933
rect -5638 -23967 -5628 -23933
rect -5004 -23967 -4994 -23933
rect -4994 -23967 -4970 -23933
rect -4932 -23967 -4926 -23933
rect -4926 -23967 -4898 -23933
rect -4860 -23967 -4858 -23933
rect -4858 -23967 -4826 -23933
rect -4788 -23967 -4756 -23933
rect -4756 -23967 -4754 -23933
rect -4716 -23967 -4688 -23933
rect -4688 -23967 -4682 -23933
rect -4644 -23967 -4620 -23933
rect -4620 -23967 -4610 -23933
rect -3986 -23967 -3976 -23933
rect -3976 -23967 -3952 -23933
rect -3914 -23967 -3908 -23933
rect -3908 -23967 -3880 -23933
rect -3842 -23967 -3840 -23933
rect -3840 -23967 -3808 -23933
rect -3770 -23967 -3738 -23933
rect -3738 -23967 -3736 -23933
rect -3698 -23967 -3670 -23933
rect -3670 -23967 -3664 -23933
rect -3626 -23967 -3602 -23933
rect -3602 -23967 -3592 -23933
rect -2263 -23966 -2229 -23932
rect -1965 -23966 -1931 -23932
rect -1667 -23966 -1633 -23932
rect -1369 -23966 -1335 -23932
rect -1071 -23966 -1037 -23932
rect -773 -23966 -739 -23932
rect -475 -23966 -441 -23932
rect -177 -23966 -143 -23932
rect 121 -23966 155 -23932
rect 419 -23966 453 -23932
rect 717 -23966 751 -23932
rect 24855 -23909 24889 -23899
rect 24855 -23933 24889 -23909
rect -12289 -24045 -12255 -24043
rect -12289 -24077 -12255 -24045
rect -12289 -24147 -12255 -24115
rect -12289 -24149 -12255 -24147
rect -12289 -24215 -12255 -24187
rect -12289 -24221 -12255 -24215
rect -12289 -24283 -12255 -24259
rect -12289 -24293 -12255 -24283
rect -12289 -24351 -12255 -24331
rect -12289 -24365 -12255 -24351
rect -12289 -24419 -12255 -24403
rect -12289 -24437 -12255 -24419
rect -12289 -24487 -12255 -24475
rect -12289 -24509 -12255 -24487
rect -12289 -24555 -12255 -24547
rect -12289 -24581 -12255 -24555
rect -9405 -24050 -9371 -24036
rect -9405 -24070 -9371 -24050
rect -9405 -24118 -9371 -24108
rect -9405 -24142 -9371 -24118
rect -9405 -24186 -9371 -24180
rect -9405 -24214 -9371 -24186
rect -9405 -24254 -9371 -24252
rect -9405 -24286 -9371 -24254
rect -9405 -24356 -9371 -24324
rect -9405 -24358 -9371 -24356
rect -9405 -24424 -9371 -24396
rect -9405 -24430 -9371 -24424
rect -9405 -24492 -9371 -24468
rect -9405 -24502 -9371 -24492
rect -9405 -24560 -9371 -24540
rect -9405 -24574 -9371 -24560
rect -8387 -24050 -8353 -24036
rect -8387 -24070 -8353 -24050
rect -8387 -24118 -8353 -24108
rect -8387 -24142 -8353 -24118
rect -8387 -24186 -8353 -24180
rect -8387 -24214 -8353 -24186
rect -8387 -24254 -8353 -24252
rect -8387 -24286 -8353 -24254
rect -8387 -24356 -8353 -24324
rect -8387 -24358 -8353 -24356
rect -8387 -24424 -8353 -24396
rect -8387 -24430 -8353 -24424
rect -8387 -24492 -8353 -24468
rect -8387 -24502 -8353 -24492
rect -8387 -24560 -8353 -24540
rect -8387 -24574 -8353 -24560
rect -7369 -24050 -7335 -24036
rect -7369 -24070 -7335 -24050
rect -7369 -24118 -7335 -24108
rect -7369 -24142 -7335 -24118
rect -7369 -24186 -7335 -24180
rect -7369 -24214 -7335 -24186
rect -7369 -24254 -7335 -24252
rect -7369 -24286 -7335 -24254
rect -7369 -24356 -7335 -24324
rect -7369 -24358 -7335 -24356
rect -7369 -24424 -7335 -24396
rect -7369 -24430 -7335 -24424
rect -7369 -24492 -7335 -24468
rect -7369 -24502 -7335 -24492
rect -7369 -24560 -7335 -24540
rect -7369 -24574 -7335 -24560
rect -6351 -24050 -6317 -24036
rect -6351 -24070 -6317 -24050
rect -6351 -24118 -6317 -24108
rect -6351 -24142 -6317 -24118
rect -6351 -24186 -6317 -24180
rect -6351 -24214 -6317 -24186
rect -6351 -24254 -6317 -24252
rect -6351 -24286 -6317 -24254
rect -6351 -24356 -6317 -24324
rect -6351 -24358 -6317 -24356
rect -6351 -24424 -6317 -24396
rect -6351 -24430 -6317 -24424
rect -6351 -24492 -6317 -24468
rect -6351 -24502 -6317 -24492
rect -6351 -24560 -6317 -24540
rect -6351 -24574 -6317 -24560
rect -5333 -24050 -5299 -24036
rect -5333 -24070 -5299 -24050
rect -5333 -24118 -5299 -24108
rect -5333 -24142 -5299 -24118
rect -5333 -24186 -5299 -24180
rect -5333 -24214 -5299 -24186
rect -5333 -24254 -5299 -24252
rect -5333 -24286 -5299 -24254
rect -5333 -24356 -5299 -24324
rect -5333 -24358 -5299 -24356
rect -5333 -24424 -5299 -24396
rect -5333 -24430 -5299 -24424
rect -5333 -24492 -5299 -24468
rect -5333 -24502 -5299 -24492
rect -5333 -24560 -5299 -24540
rect -5333 -24574 -5299 -24560
rect -4315 -24050 -4281 -24036
rect -4315 -24070 -4281 -24050
rect -4315 -24118 -4281 -24108
rect -4315 -24142 -4281 -24118
rect -4315 -24186 -4281 -24180
rect -4315 -24214 -4281 -24186
rect -4315 -24254 -4281 -24252
rect -4315 -24286 -4281 -24254
rect -4315 -24356 -4281 -24324
rect -4315 -24358 -4281 -24356
rect -4315 -24424 -4281 -24396
rect -4315 -24430 -4281 -24424
rect -4315 -24492 -4281 -24468
rect -4315 -24502 -4281 -24492
rect -4315 -24560 -4281 -24540
rect -4315 -24574 -4281 -24560
rect -3297 -24050 -3263 -24036
rect -3297 -24070 -3263 -24050
rect -3297 -24118 -3263 -24108
rect -3297 -24142 -3263 -24118
rect -3297 -24186 -3263 -24180
rect -3297 -24214 -3263 -24186
rect -3297 -24254 -3263 -24252
rect -3297 -24286 -3263 -24254
rect -3297 -24356 -3263 -24324
rect -3297 -24358 -3263 -24356
rect -3297 -24424 -3263 -24396
rect -3297 -24430 -3263 -24424
rect -3297 -24492 -3263 -24468
rect -3297 -24502 -3263 -24492
rect -3297 -24560 -3263 -24540
rect -3297 -24574 -3263 -24560
rect -2412 -24049 -2378 -24035
rect -2412 -24069 -2378 -24049
rect -2412 -24117 -2378 -24107
rect -2412 -24141 -2378 -24117
rect -2412 -24185 -2378 -24179
rect -2412 -24213 -2378 -24185
rect -2412 -24253 -2378 -24251
rect -2412 -24285 -2378 -24253
rect -2412 -24355 -2378 -24323
rect -2412 -24357 -2378 -24355
rect -2412 -24423 -2378 -24395
rect -2412 -24429 -2378 -24423
rect -2412 -24491 -2378 -24467
rect -2412 -24501 -2378 -24491
rect -2412 -24559 -2378 -24539
rect -2412 -24573 -2378 -24559
rect -2114 -24049 -2080 -24035
rect -2114 -24069 -2080 -24049
rect -2114 -24117 -2080 -24107
rect -2114 -24141 -2080 -24117
rect -2114 -24185 -2080 -24179
rect -2114 -24213 -2080 -24185
rect -2114 -24253 -2080 -24251
rect -2114 -24285 -2080 -24253
rect -2114 -24355 -2080 -24323
rect -2114 -24357 -2080 -24355
rect -2114 -24423 -2080 -24395
rect -2114 -24429 -2080 -24423
rect -2114 -24491 -2080 -24467
rect -2114 -24501 -2080 -24491
rect -2114 -24559 -2080 -24539
rect -2114 -24573 -2080 -24559
rect -1816 -24049 -1782 -24035
rect -1816 -24069 -1782 -24049
rect -1816 -24117 -1782 -24107
rect -1816 -24141 -1782 -24117
rect -1816 -24185 -1782 -24179
rect -1816 -24213 -1782 -24185
rect -1816 -24253 -1782 -24251
rect -1816 -24285 -1782 -24253
rect -1816 -24355 -1782 -24323
rect -1816 -24357 -1782 -24355
rect -1816 -24423 -1782 -24395
rect -1816 -24429 -1782 -24423
rect -1816 -24491 -1782 -24467
rect -1816 -24501 -1782 -24491
rect -1816 -24559 -1782 -24539
rect -1816 -24573 -1782 -24559
rect -1518 -24049 -1484 -24035
rect -1518 -24069 -1484 -24049
rect -1518 -24117 -1484 -24107
rect -1518 -24141 -1484 -24117
rect -1518 -24185 -1484 -24179
rect -1518 -24213 -1484 -24185
rect -1518 -24253 -1484 -24251
rect -1518 -24285 -1484 -24253
rect -1518 -24355 -1484 -24323
rect -1518 -24357 -1484 -24355
rect -1518 -24423 -1484 -24395
rect -1518 -24429 -1484 -24423
rect -1518 -24491 -1484 -24467
rect -1518 -24501 -1484 -24491
rect -1518 -24559 -1484 -24539
rect -1518 -24573 -1484 -24559
rect -1220 -24049 -1186 -24035
rect -1220 -24069 -1186 -24049
rect -1220 -24117 -1186 -24107
rect -1220 -24141 -1186 -24117
rect -1220 -24185 -1186 -24179
rect -1220 -24213 -1186 -24185
rect -1220 -24253 -1186 -24251
rect -1220 -24285 -1186 -24253
rect -1220 -24355 -1186 -24323
rect -1220 -24357 -1186 -24355
rect -1220 -24423 -1186 -24395
rect -1220 -24429 -1186 -24423
rect -1220 -24491 -1186 -24467
rect -1220 -24501 -1186 -24491
rect -1220 -24559 -1186 -24539
rect -1220 -24573 -1186 -24559
rect -922 -24049 -888 -24035
rect -922 -24069 -888 -24049
rect -922 -24117 -888 -24107
rect -922 -24141 -888 -24117
rect -922 -24185 -888 -24179
rect -922 -24213 -888 -24185
rect -922 -24253 -888 -24251
rect -922 -24285 -888 -24253
rect -922 -24355 -888 -24323
rect -922 -24357 -888 -24355
rect -922 -24423 -888 -24395
rect -922 -24429 -888 -24423
rect -922 -24491 -888 -24467
rect -922 -24501 -888 -24491
rect -922 -24559 -888 -24539
rect -922 -24573 -888 -24559
rect -624 -24049 -590 -24035
rect -624 -24069 -590 -24049
rect -624 -24117 -590 -24107
rect -624 -24141 -590 -24117
rect -624 -24185 -590 -24179
rect -624 -24213 -590 -24185
rect -624 -24253 -590 -24251
rect -624 -24285 -590 -24253
rect -624 -24355 -590 -24323
rect -624 -24357 -590 -24355
rect -624 -24423 -590 -24395
rect -624 -24429 -590 -24423
rect -624 -24491 -590 -24467
rect -624 -24501 -590 -24491
rect -624 -24559 -590 -24539
rect -624 -24573 -590 -24559
rect -326 -24049 -292 -24035
rect -326 -24069 -292 -24049
rect -326 -24117 -292 -24107
rect -326 -24141 -292 -24117
rect -326 -24185 -292 -24179
rect -326 -24213 -292 -24185
rect -326 -24253 -292 -24251
rect -326 -24285 -292 -24253
rect -326 -24355 -292 -24323
rect -326 -24357 -292 -24355
rect -326 -24423 -292 -24395
rect -326 -24429 -292 -24423
rect -326 -24491 -292 -24467
rect -326 -24501 -292 -24491
rect -326 -24559 -292 -24539
rect -326 -24573 -292 -24559
rect -28 -24049 6 -24035
rect -28 -24069 6 -24049
rect -28 -24117 6 -24107
rect -28 -24141 6 -24117
rect -28 -24185 6 -24179
rect -28 -24213 6 -24185
rect -28 -24253 6 -24251
rect -28 -24285 6 -24253
rect -28 -24355 6 -24323
rect -28 -24357 6 -24355
rect -28 -24423 6 -24395
rect -28 -24429 6 -24423
rect -28 -24491 6 -24467
rect -28 -24501 6 -24491
rect -28 -24559 6 -24539
rect -28 -24573 6 -24559
rect 270 -24049 304 -24035
rect 270 -24069 304 -24049
rect 270 -24117 304 -24107
rect 270 -24141 304 -24117
rect 270 -24185 304 -24179
rect 270 -24213 304 -24185
rect 270 -24253 304 -24251
rect 270 -24285 304 -24253
rect 270 -24355 304 -24323
rect 270 -24357 304 -24355
rect 270 -24423 304 -24395
rect 270 -24429 304 -24423
rect 270 -24491 304 -24467
rect 270 -24501 304 -24491
rect 270 -24559 304 -24539
rect 270 -24573 304 -24559
rect 568 -24049 602 -24035
rect 568 -24069 602 -24049
rect 568 -24117 602 -24107
rect 568 -24141 602 -24117
rect 568 -24185 602 -24179
rect 568 -24213 602 -24185
rect 568 -24253 602 -24251
rect 568 -24285 602 -24253
rect 568 -24355 602 -24323
rect 568 -24357 602 -24355
rect 568 -24423 602 -24395
rect 568 -24429 602 -24423
rect 568 -24491 602 -24467
rect 568 -24501 602 -24491
rect 568 -24559 602 -24539
rect 568 -24573 602 -24559
rect 2909 -24014 2919 -23980
rect 2919 -24014 2943 -23980
rect 2981 -24014 2987 -23980
rect 2987 -24014 3015 -23980
rect 3053 -24014 3055 -23980
rect 3055 -24014 3087 -23980
rect 3125 -24014 3157 -23980
rect 3157 -24014 3159 -23980
rect 3197 -24014 3225 -23980
rect 3225 -24014 3231 -23980
rect 3269 -24014 3293 -23980
rect 3293 -24014 3303 -23980
rect 3927 -24014 3937 -23980
rect 3937 -24014 3961 -23980
rect 3999 -24014 4005 -23980
rect 4005 -24014 4033 -23980
rect 4071 -24014 4073 -23980
rect 4073 -24014 4105 -23980
rect 4143 -24014 4175 -23980
rect 4175 -24014 4177 -23980
rect 4215 -24014 4243 -23980
rect 4243 -24014 4249 -23980
rect 4287 -24014 4311 -23980
rect 4311 -24014 4321 -23980
rect 4945 -24014 4955 -23980
rect 4955 -24014 4979 -23980
rect 5017 -24014 5023 -23980
rect 5023 -24014 5051 -23980
rect 5089 -24014 5091 -23980
rect 5091 -24014 5123 -23980
rect 5161 -24014 5193 -23980
rect 5193 -24014 5195 -23980
rect 5233 -24014 5261 -23980
rect 5261 -24014 5267 -23980
rect 5305 -24014 5329 -23980
rect 5329 -24014 5339 -23980
rect 5963 -24014 5973 -23980
rect 5973 -24014 5997 -23980
rect 6035 -24014 6041 -23980
rect 6041 -24014 6069 -23980
rect 6107 -24014 6109 -23980
rect 6109 -24014 6141 -23980
rect 6179 -24014 6211 -23980
rect 6211 -24014 6213 -23980
rect 6251 -24014 6279 -23980
rect 6279 -24014 6285 -23980
rect 6323 -24014 6347 -23980
rect 6347 -24014 6357 -23980
rect 6981 -24014 6991 -23980
rect 6991 -24014 7015 -23980
rect 7053 -24014 7059 -23980
rect 7059 -24014 7087 -23980
rect 7125 -24014 7127 -23980
rect 7127 -24014 7159 -23980
rect 7197 -24014 7229 -23980
rect 7229 -24014 7231 -23980
rect 7269 -24014 7297 -23980
rect 7297 -24014 7303 -23980
rect 7341 -24014 7365 -23980
rect 7365 -24014 7375 -23980
rect 7999 -24014 8009 -23980
rect 8009 -24014 8033 -23980
rect 8071 -24014 8077 -23980
rect 8077 -24014 8105 -23980
rect 8143 -24014 8145 -23980
rect 8145 -24014 8177 -23980
rect 8215 -24014 8247 -23980
rect 8247 -24014 8249 -23980
rect 8287 -24014 8315 -23980
rect 8315 -24014 8321 -23980
rect 8359 -24014 8383 -23980
rect 8383 -24014 8393 -23980
rect 9017 -24014 9027 -23980
rect 9027 -24014 9051 -23980
rect 9089 -24014 9095 -23980
rect 9095 -24014 9123 -23980
rect 9161 -24014 9163 -23980
rect 9163 -24014 9195 -23980
rect 9233 -24014 9265 -23980
rect 9265 -24014 9267 -23980
rect 9305 -24014 9333 -23980
rect 9333 -24014 9339 -23980
rect 9377 -24014 9401 -23980
rect 9401 -24014 9411 -23980
rect 10035 -24014 10045 -23980
rect 10045 -24014 10069 -23980
rect 10107 -24014 10113 -23980
rect 10113 -24014 10141 -23980
rect 10179 -24014 10181 -23980
rect 10181 -24014 10213 -23980
rect 10251 -24014 10283 -23980
rect 10283 -24014 10285 -23980
rect 10323 -24014 10351 -23980
rect 10351 -24014 10357 -23980
rect 10395 -24014 10419 -23980
rect 10419 -24014 10429 -23980
rect 11053 -24014 11063 -23980
rect 11063 -24014 11087 -23980
rect 11125 -24014 11131 -23980
rect 11131 -24014 11159 -23980
rect 11197 -24014 11199 -23980
rect 11199 -24014 11231 -23980
rect 11269 -24014 11301 -23980
rect 11301 -24014 11303 -23980
rect 11341 -24014 11369 -23980
rect 11369 -24014 11375 -23980
rect 11413 -24014 11437 -23980
rect 11437 -24014 11447 -23980
rect 12071 -24014 12081 -23980
rect 12081 -24014 12105 -23980
rect 12143 -24014 12149 -23980
rect 12149 -24014 12177 -23980
rect 12215 -24014 12217 -23980
rect 12217 -24014 12249 -23980
rect 12287 -24014 12319 -23980
rect 12319 -24014 12321 -23980
rect 12359 -24014 12387 -23980
rect 12387 -24014 12393 -23980
rect 12431 -24014 12455 -23980
rect 12455 -24014 12465 -23980
rect 13089 -24014 13099 -23980
rect 13099 -24014 13123 -23980
rect 13161 -24014 13167 -23980
rect 13167 -24014 13195 -23980
rect 13233 -24014 13235 -23980
rect 13235 -24014 13267 -23980
rect 13305 -24014 13337 -23980
rect 13337 -24014 13339 -23980
rect 13377 -24014 13405 -23980
rect 13405 -24014 13411 -23980
rect 13449 -24014 13473 -23980
rect 13473 -24014 13483 -23980
rect 14107 -24014 14117 -23980
rect 14117 -24014 14141 -23980
rect 14179 -24014 14185 -23980
rect 14185 -24014 14213 -23980
rect 14251 -24014 14253 -23980
rect 14253 -24014 14285 -23980
rect 14323 -24014 14355 -23980
rect 14355 -24014 14357 -23980
rect 14395 -24014 14423 -23980
rect 14423 -24014 14429 -23980
rect 14467 -24014 14491 -23980
rect 14491 -24014 14501 -23980
rect 15125 -24014 15135 -23980
rect 15135 -24014 15159 -23980
rect 15197 -24014 15203 -23980
rect 15203 -24014 15231 -23980
rect 15269 -24014 15271 -23980
rect 15271 -24014 15303 -23980
rect 15341 -24014 15373 -23980
rect 15373 -24014 15375 -23980
rect 15413 -24014 15441 -23980
rect 15441 -24014 15447 -23980
rect 15485 -24014 15509 -23980
rect 15509 -24014 15519 -23980
rect 16143 -24014 16153 -23980
rect 16153 -24014 16177 -23980
rect 16215 -24014 16221 -23980
rect 16221 -24014 16249 -23980
rect 16287 -24014 16289 -23980
rect 16289 -24014 16321 -23980
rect 16359 -24014 16391 -23980
rect 16391 -24014 16393 -23980
rect 16431 -24014 16459 -23980
rect 16459 -24014 16465 -23980
rect 16503 -24014 16527 -23980
rect 16527 -24014 16537 -23980
rect 17161 -24014 17171 -23980
rect 17171 -24014 17195 -23980
rect 17233 -24014 17239 -23980
rect 17239 -24014 17267 -23980
rect 17305 -24014 17307 -23980
rect 17307 -24014 17339 -23980
rect 17377 -24014 17409 -23980
rect 17409 -24014 17411 -23980
rect 17449 -24014 17477 -23980
rect 17477 -24014 17483 -23980
rect 17521 -24014 17545 -23980
rect 17545 -24014 17555 -23980
rect 18179 -24014 18189 -23980
rect 18189 -24014 18213 -23980
rect 18251 -24014 18257 -23980
rect 18257 -24014 18285 -23980
rect 18323 -24014 18325 -23980
rect 18325 -24014 18357 -23980
rect 18395 -24014 18427 -23980
rect 18427 -24014 18429 -23980
rect 18467 -24014 18495 -23980
rect 18495 -24014 18501 -23980
rect 18539 -24014 18563 -23980
rect 18563 -24014 18573 -23980
rect 19197 -24014 19207 -23980
rect 19207 -24014 19231 -23980
rect 19269 -24014 19275 -23980
rect 19275 -24014 19303 -23980
rect 19341 -24014 19343 -23980
rect 19343 -24014 19375 -23980
rect 19413 -24014 19445 -23980
rect 19445 -24014 19447 -23980
rect 19485 -24014 19513 -23980
rect 19513 -24014 19519 -23980
rect 19557 -24014 19581 -23980
rect 19581 -24014 19591 -23980
rect 20215 -24014 20225 -23980
rect 20225 -24014 20249 -23980
rect 20287 -24014 20293 -23980
rect 20293 -24014 20321 -23980
rect 20359 -24014 20361 -23980
rect 20361 -24014 20393 -23980
rect 20431 -24014 20463 -23980
rect 20463 -24014 20465 -23980
rect 20503 -24014 20531 -23980
rect 20531 -24014 20537 -23980
rect 20575 -24014 20599 -23980
rect 20599 -24014 20609 -23980
rect 21233 -24014 21243 -23980
rect 21243 -24014 21267 -23980
rect 21305 -24014 21311 -23980
rect 21311 -24014 21339 -23980
rect 21377 -24014 21379 -23980
rect 21379 -24014 21411 -23980
rect 21449 -24014 21481 -23980
rect 21481 -24014 21483 -23980
rect 21521 -24014 21549 -23980
rect 21549 -24014 21555 -23980
rect 21593 -24014 21617 -23980
rect 21617 -24014 21627 -23980
rect 22251 -24014 22261 -23980
rect 22261 -24014 22285 -23980
rect 22323 -24014 22329 -23980
rect 22329 -24014 22357 -23980
rect 22395 -24014 22397 -23980
rect 22397 -24014 22429 -23980
rect 22467 -24014 22499 -23980
rect 22499 -24014 22501 -23980
rect 22539 -24014 22567 -23980
rect 22567 -24014 22573 -23980
rect 22611 -24014 22635 -23980
rect 22635 -24014 22645 -23980
rect 24855 -23977 24889 -23971
rect 24855 -24005 24889 -23977
rect 866 -24049 900 -24035
rect 866 -24069 900 -24049
rect 866 -24117 900 -24107
rect 866 -24141 900 -24117
rect 866 -24185 900 -24179
rect 866 -24213 900 -24185
rect 866 -24253 900 -24251
rect 866 -24285 900 -24253
rect 866 -24355 900 -24323
rect 866 -24357 900 -24355
rect 866 -24423 900 -24395
rect 866 -24429 900 -24423
rect 866 -24491 900 -24467
rect 866 -24501 900 -24491
rect 866 -24559 900 -24539
rect 866 -24573 900 -24559
rect 2580 -24097 2614 -24083
rect 2580 -24117 2614 -24097
rect 2580 -24165 2614 -24155
rect 2580 -24189 2614 -24165
rect 2580 -24233 2614 -24227
rect 2580 -24261 2614 -24233
rect 2580 -24301 2614 -24299
rect 2580 -24333 2614 -24301
rect 2580 -24403 2614 -24371
rect 2580 -24405 2614 -24403
rect 2580 -24471 2614 -24443
rect 2580 -24477 2614 -24471
rect 2580 -24539 2614 -24515
rect 2580 -24549 2614 -24539
rect 2580 -24607 2614 -24587
rect -12289 -24623 -12255 -24619
rect -12289 -24653 -12255 -24623
rect 2580 -24621 2614 -24607
rect -9076 -24677 -9066 -24643
rect -9066 -24677 -9042 -24643
rect -9004 -24677 -8998 -24643
rect -8998 -24677 -8970 -24643
rect -8932 -24677 -8930 -24643
rect -8930 -24677 -8898 -24643
rect -8860 -24677 -8828 -24643
rect -8828 -24677 -8826 -24643
rect -8788 -24677 -8760 -24643
rect -8760 -24677 -8754 -24643
rect -8716 -24677 -8692 -24643
rect -8692 -24677 -8682 -24643
rect -8058 -24677 -8048 -24643
rect -8048 -24677 -8024 -24643
rect -7986 -24677 -7980 -24643
rect -7980 -24677 -7952 -24643
rect -7914 -24677 -7912 -24643
rect -7912 -24677 -7880 -24643
rect -7842 -24677 -7810 -24643
rect -7810 -24677 -7808 -24643
rect -7770 -24677 -7742 -24643
rect -7742 -24677 -7736 -24643
rect -7698 -24677 -7674 -24643
rect -7674 -24677 -7664 -24643
rect -7040 -24677 -7030 -24643
rect -7030 -24677 -7006 -24643
rect -6968 -24677 -6962 -24643
rect -6962 -24677 -6934 -24643
rect -6896 -24677 -6894 -24643
rect -6894 -24677 -6862 -24643
rect -6824 -24677 -6792 -24643
rect -6792 -24677 -6790 -24643
rect -6752 -24677 -6724 -24643
rect -6724 -24677 -6718 -24643
rect -6680 -24677 -6656 -24643
rect -6656 -24677 -6646 -24643
rect -6022 -24677 -6012 -24643
rect -6012 -24677 -5988 -24643
rect -5950 -24677 -5944 -24643
rect -5944 -24677 -5916 -24643
rect -5878 -24677 -5876 -24643
rect -5876 -24677 -5844 -24643
rect -5806 -24677 -5774 -24643
rect -5774 -24677 -5772 -24643
rect -5734 -24677 -5706 -24643
rect -5706 -24677 -5700 -24643
rect -5662 -24677 -5638 -24643
rect -5638 -24677 -5628 -24643
rect -5004 -24677 -4994 -24643
rect -4994 -24677 -4970 -24643
rect -4932 -24677 -4926 -24643
rect -4926 -24677 -4898 -24643
rect -4860 -24677 -4858 -24643
rect -4858 -24677 -4826 -24643
rect -4788 -24677 -4756 -24643
rect -4756 -24677 -4754 -24643
rect -4716 -24677 -4688 -24643
rect -4688 -24677 -4682 -24643
rect -4644 -24677 -4620 -24643
rect -4620 -24677 -4610 -24643
rect -3986 -24677 -3976 -24643
rect -3976 -24677 -3952 -24643
rect -3914 -24677 -3908 -24643
rect -3908 -24677 -3880 -24643
rect -3842 -24677 -3840 -24643
rect -3840 -24677 -3808 -24643
rect -3770 -24677 -3738 -24643
rect -3738 -24677 -3736 -24643
rect -3698 -24677 -3670 -24643
rect -3670 -24677 -3664 -24643
rect -3626 -24677 -3602 -24643
rect -3602 -24677 -3592 -24643
rect -2263 -24676 -2229 -24642
rect -1965 -24676 -1931 -24642
rect -1667 -24676 -1633 -24642
rect -1369 -24676 -1335 -24642
rect -1071 -24676 -1037 -24642
rect -773 -24676 -739 -24642
rect -475 -24676 -441 -24642
rect -177 -24676 -143 -24642
rect 121 -24676 155 -24642
rect 419 -24676 453 -24642
rect 717 -24676 751 -24642
rect 3598 -24097 3632 -24083
rect 3598 -24117 3632 -24097
rect 3598 -24165 3632 -24155
rect 3598 -24189 3632 -24165
rect 3598 -24233 3632 -24227
rect 3598 -24261 3632 -24233
rect 3598 -24301 3632 -24299
rect 3598 -24333 3632 -24301
rect 3598 -24403 3632 -24371
rect 3598 -24405 3632 -24403
rect 3598 -24471 3632 -24443
rect 3598 -24477 3632 -24471
rect 3598 -24539 3632 -24515
rect 3598 -24549 3632 -24539
rect 3598 -24607 3632 -24587
rect 3598 -24621 3632 -24607
rect 4616 -24097 4650 -24083
rect 4616 -24117 4650 -24097
rect 4616 -24165 4650 -24155
rect 4616 -24189 4650 -24165
rect 4616 -24233 4650 -24227
rect 4616 -24261 4650 -24233
rect 4616 -24301 4650 -24299
rect 4616 -24333 4650 -24301
rect 4616 -24403 4650 -24371
rect 4616 -24405 4650 -24403
rect 4616 -24471 4650 -24443
rect 4616 -24477 4650 -24471
rect 4616 -24539 4650 -24515
rect 4616 -24549 4650 -24539
rect 4616 -24607 4650 -24587
rect 4616 -24621 4650 -24607
rect 5634 -24097 5668 -24083
rect 5634 -24117 5668 -24097
rect 5634 -24165 5668 -24155
rect 5634 -24189 5668 -24165
rect 5634 -24233 5668 -24227
rect 5634 -24261 5668 -24233
rect 5634 -24301 5668 -24299
rect 5634 -24333 5668 -24301
rect 5634 -24403 5668 -24371
rect 5634 -24405 5668 -24403
rect 5634 -24471 5668 -24443
rect 5634 -24477 5668 -24471
rect 5634 -24539 5668 -24515
rect 5634 -24549 5668 -24539
rect 5634 -24607 5668 -24587
rect 5634 -24621 5668 -24607
rect 6652 -24097 6686 -24083
rect 6652 -24117 6686 -24097
rect 6652 -24165 6686 -24155
rect 6652 -24189 6686 -24165
rect 6652 -24233 6686 -24227
rect 6652 -24261 6686 -24233
rect 6652 -24301 6686 -24299
rect 6652 -24333 6686 -24301
rect 6652 -24403 6686 -24371
rect 6652 -24405 6686 -24403
rect 6652 -24471 6686 -24443
rect 6652 -24477 6686 -24471
rect 6652 -24539 6686 -24515
rect 6652 -24549 6686 -24539
rect 6652 -24607 6686 -24587
rect 6652 -24621 6686 -24607
rect 7670 -24097 7704 -24083
rect 7670 -24117 7704 -24097
rect 7670 -24165 7704 -24155
rect 7670 -24189 7704 -24165
rect 7670 -24233 7704 -24227
rect 7670 -24261 7704 -24233
rect 7670 -24301 7704 -24299
rect 7670 -24333 7704 -24301
rect 7670 -24403 7704 -24371
rect 7670 -24405 7704 -24403
rect 7670 -24471 7704 -24443
rect 7670 -24477 7704 -24471
rect 7670 -24539 7704 -24515
rect 7670 -24549 7704 -24539
rect 7670 -24607 7704 -24587
rect 7670 -24621 7704 -24607
rect 8688 -24097 8722 -24083
rect 8688 -24117 8722 -24097
rect 8688 -24165 8722 -24155
rect 8688 -24189 8722 -24165
rect 8688 -24233 8722 -24227
rect 8688 -24261 8722 -24233
rect 8688 -24301 8722 -24299
rect 8688 -24333 8722 -24301
rect 8688 -24403 8722 -24371
rect 8688 -24405 8722 -24403
rect 8688 -24471 8722 -24443
rect 8688 -24477 8722 -24471
rect 8688 -24539 8722 -24515
rect 8688 -24549 8722 -24539
rect 8688 -24607 8722 -24587
rect 8688 -24621 8722 -24607
rect 9706 -24097 9740 -24083
rect 9706 -24117 9740 -24097
rect 9706 -24165 9740 -24155
rect 9706 -24189 9740 -24165
rect 9706 -24233 9740 -24227
rect 9706 -24261 9740 -24233
rect 9706 -24301 9740 -24299
rect 9706 -24333 9740 -24301
rect 9706 -24403 9740 -24371
rect 9706 -24405 9740 -24403
rect 9706 -24471 9740 -24443
rect 9706 -24477 9740 -24471
rect 9706 -24539 9740 -24515
rect 9706 -24549 9740 -24539
rect 9706 -24607 9740 -24587
rect 9706 -24621 9740 -24607
rect 10724 -24097 10758 -24083
rect 10724 -24117 10758 -24097
rect 10724 -24165 10758 -24155
rect 10724 -24189 10758 -24165
rect 10724 -24233 10758 -24227
rect 10724 -24261 10758 -24233
rect 10724 -24301 10758 -24299
rect 10724 -24333 10758 -24301
rect 10724 -24403 10758 -24371
rect 10724 -24405 10758 -24403
rect 10724 -24471 10758 -24443
rect 10724 -24477 10758 -24471
rect 10724 -24539 10758 -24515
rect 10724 -24549 10758 -24539
rect 10724 -24607 10758 -24587
rect 10724 -24621 10758 -24607
rect 11742 -24097 11776 -24083
rect 11742 -24117 11776 -24097
rect 11742 -24165 11776 -24155
rect 11742 -24189 11776 -24165
rect 11742 -24233 11776 -24227
rect 11742 -24261 11776 -24233
rect 11742 -24301 11776 -24299
rect 11742 -24333 11776 -24301
rect 11742 -24403 11776 -24371
rect 11742 -24405 11776 -24403
rect 11742 -24471 11776 -24443
rect 11742 -24477 11776 -24471
rect 11742 -24539 11776 -24515
rect 11742 -24549 11776 -24539
rect 11742 -24607 11776 -24587
rect 11742 -24621 11776 -24607
rect 12760 -24097 12794 -24083
rect 12760 -24117 12794 -24097
rect 12760 -24165 12794 -24155
rect 12760 -24189 12794 -24165
rect 12760 -24233 12794 -24227
rect 12760 -24261 12794 -24233
rect 12760 -24301 12794 -24299
rect 12760 -24333 12794 -24301
rect 12760 -24403 12794 -24371
rect 12760 -24405 12794 -24403
rect 12760 -24471 12794 -24443
rect 12760 -24477 12794 -24471
rect 12760 -24539 12794 -24515
rect 12760 -24549 12794 -24539
rect 12760 -24607 12794 -24587
rect 12760 -24621 12794 -24607
rect 13778 -24097 13812 -24083
rect 13778 -24117 13812 -24097
rect 13778 -24165 13812 -24155
rect 13778 -24189 13812 -24165
rect 13778 -24233 13812 -24227
rect 13778 -24261 13812 -24233
rect 13778 -24301 13812 -24299
rect 13778 -24333 13812 -24301
rect 13778 -24403 13812 -24371
rect 13778 -24405 13812 -24403
rect 13778 -24471 13812 -24443
rect 13778 -24477 13812 -24471
rect 13778 -24539 13812 -24515
rect 13778 -24549 13812 -24539
rect 13778 -24607 13812 -24587
rect 13778 -24621 13812 -24607
rect 14796 -24097 14830 -24083
rect 14796 -24117 14830 -24097
rect 14796 -24165 14830 -24155
rect 14796 -24189 14830 -24165
rect 14796 -24233 14830 -24227
rect 14796 -24261 14830 -24233
rect 14796 -24301 14830 -24299
rect 14796 -24333 14830 -24301
rect 14796 -24403 14830 -24371
rect 14796 -24405 14830 -24403
rect 14796 -24471 14830 -24443
rect 14796 -24477 14830 -24471
rect 14796 -24539 14830 -24515
rect 14796 -24549 14830 -24539
rect 14796 -24607 14830 -24587
rect 14796 -24621 14830 -24607
rect 15814 -24097 15848 -24083
rect 15814 -24117 15848 -24097
rect 15814 -24165 15848 -24155
rect 15814 -24189 15848 -24165
rect 15814 -24233 15848 -24227
rect 15814 -24261 15848 -24233
rect 15814 -24301 15848 -24299
rect 15814 -24333 15848 -24301
rect 15814 -24403 15848 -24371
rect 15814 -24405 15848 -24403
rect 15814 -24471 15848 -24443
rect 15814 -24477 15848 -24471
rect 15814 -24539 15848 -24515
rect 15814 -24549 15848 -24539
rect 15814 -24607 15848 -24587
rect 15814 -24621 15848 -24607
rect 16832 -24097 16866 -24083
rect 16832 -24117 16866 -24097
rect 16832 -24165 16866 -24155
rect 16832 -24189 16866 -24165
rect 16832 -24233 16866 -24227
rect 16832 -24261 16866 -24233
rect 16832 -24301 16866 -24299
rect 16832 -24333 16866 -24301
rect 16832 -24403 16866 -24371
rect 16832 -24405 16866 -24403
rect 16832 -24471 16866 -24443
rect 16832 -24477 16866 -24471
rect 16832 -24539 16866 -24515
rect 16832 -24549 16866 -24539
rect 16832 -24607 16866 -24587
rect 16832 -24621 16866 -24607
rect 17850 -24097 17884 -24083
rect 17850 -24117 17884 -24097
rect 17850 -24165 17884 -24155
rect 17850 -24189 17884 -24165
rect 17850 -24233 17884 -24227
rect 17850 -24261 17884 -24233
rect 17850 -24301 17884 -24299
rect 17850 -24333 17884 -24301
rect 17850 -24403 17884 -24371
rect 17850 -24405 17884 -24403
rect 17850 -24471 17884 -24443
rect 17850 -24477 17884 -24471
rect 17850 -24539 17884 -24515
rect 17850 -24549 17884 -24539
rect 17850 -24607 17884 -24587
rect 17850 -24621 17884 -24607
rect 18868 -24097 18902 -24083
rect 18868 -24117 18902 -24097
rect 18868 -24165 18902 -24155
rect 18868 -24189 18902 -24165
rect 18868 -24233 18902 -24227
rect 18868 -24261 18902 -24233
rect 18868 -24301 18902 -24299
rect 18868 -24333 18902 -24301
rect 18868 -24403 18902 -24371
rect 18868 -24405 18902 -24403
rect 18868 -24471 18902 -24443
rect 18868 -24477 18902 -24471
rect 18868 -24539 18902 -24515
rect 18868 -24549 18902 -24539
rect 18868 -24607 18902 -24587
rect 18868 -24621 18902 -24607
rect 19886 -24097 19920 -24083
rect 19886 -24117 19920 -24097
rect 19886 -24165 19920 -24155
rect 19886 -24189 19920 -24165
rect 19886 -24233 19920 -24227
rect 19886 -24261 19920 -24233
rect 19886 -24301 19920 -24299
rect 19886 -24333 19920 -24301
rect 19886 -24403 19920 -24371
rect 19886 -24405 19920 -24403
rect 19886 -24471 19920 -24443
rect 19886 -24477 19920 -24471
rect 19886 -24539 19920 -24515
rect 19886 -24549 19920 -24539
rect 19886 -24607 19920 -24587
rect 19886 -24621 19920 -24607
rect 20904 -24097 20938 -24083
rect 20904 -24117 20938 -24097
rect 20904 -24165 20938 -24155
rect 20904 -24189 20938 -24165
rect 20904 -24233 20938 -24227
rect 20904 -24261 20938 -24233
rect 20904 -24301 20938 -24299
rect 20904 -24333 20938 -24301
rect 20904 -24403 20938 -24371
rect 20904 -24405 20938 -24403
rect 20904 -24471 20938 -24443
rect 20904 -24477 20938 -24471
rect 20904 -24539 20938 -24515
rect 20904 -24549 20938 -24539
rect 20904 -24607 20938 -24587
rect 20904 -24621 20938 -24607
rect 21922 -24097 21956 -24083
rect 21922 -24117 21956 -24097
rect 21922 -24165 21956 -24155
rect 21922 -24189 21956 -24165
rect 21922 -24233 21956 -24227
rect 21922 -24261 21956 -24233
rect 21922 -24301 21956 -24299
rect 21922 -24333 21956 -24301
rect 21922 -24403 21956 -24371
rect 21922 -24405 21956 -24403
rect 21922 -24471 21956 -24443
rect 21922 -24477 21956 -24471
rect 21922 -24539 21956 -24515
rect 21922 -24549 21956 -24539
rect 21922 -24607 21956 -24587
rect 21922 -24621 21956 -24607
rect 22940 -24097 22974 -24083
rect 22940 -24117 22974 -24097
rect 22940 -24165 22974 -24155
rect 22940 -24189 22974 -24165
rect 22940 -24233 22974 -24227
rect 22940 -24261 22974 -24233
rect 22940 -24301 22974 -24299
rect 22940 -24333 22974 -24301
rect 22940 -24403 22974 -24371
rect 22940 -24405 22974 -24403
rect 22940 -24471 22974 -24443
rect 22940 -24477 22974 -24471
rect 22940 -24539 22974 -24515
rect 22940 -24549 22974 -24539
rect 22940 -24607 22974 -24587
rect 22940 -24621 22974 -24607
rect 24855 -24045 24889 -24043
rect 24855 -24077 24889 -24045
rect 24855 -24147 24889 -24115
rect 24855 -24149 24889 -24147
rect 24855 -24215 24889 -24187
rect 24855 -24221 24889 -24215
rect 24855 -24283 24889 -24259
rect 24855 -24293 24889 -24283
rect 24855 -24351 24889 -24331
rect 24855 -24365 24889 -24351
rect 24855 -24419 24889 -24403
rect 24855 -24437 24889 -24419
rect 24855 -24487 24889 -24475
rect 24855 -24509 24889 -24487
rect 24855 -24555 24889 -24547
rect 24855 -24581 24889 -24555
rect 24855 -24623 24889 -24619
rect 24855 -24653 24889 -24623
rect -12289 -24725 -12255 -24691
rect 2909 -24724 2919 -24690
rect 2919 -24724 2943 -24690
rect 2981 -24724 2987 -24690
rect 2987 -24724 3015 -24690
rect 3053 -24724 3055 -24690
rect 3055 -24724 3087 -24690
rect 3125 -24724 3157 -24690
rect 3157 -24724 3159 -24690
rect 3197 -24724 3225 -24690
rect 3225 -24724 3231 -24690
rect 3269 -24724 3293 -24690
rect 3293 -24724 3303 -24690
rect 3927 -24724 3937 -24690
rect 3937 -24724 3961 -24690
rect 3999 -24724 4005 -24690
rect 4005 -24724 4033 -24690
rect 4071 -24724 4073 -24690
rect 4073 -24724 4105 -24690
rect 4143 -24724 4175 -24690
rect 4175 -24724 4177 -24690
rect 4215 -24724 4243 -24690
rect 4243 -24724 4249 -24690
rect 4287 -24724 4311 -24690
rect 4311 -24724 4321 -24690
rect 4945 -24724 4955 -24690
rect 4955 -24724 4979 -24690
rect 5017 -24724 5023 -24690
rect 5023 -24724 5051 -24690
rect 5089 -24724 5091 -24690
rect 5091 -24724 5123 -24690
rect 5161 -24724 5193 -24690
rect 5193 -24724 5195 -24690
rect 5233 -24724 5261 -24690
rect 5261 -24724 5267 -24690
rect 5305 -24724 5329 -24690
rect 5329 -24724 5339 -24690
rect 5963 -24724 5973 -24690
rect 5973 -24724 5997 -24690
rect 6035 -24724 6041 -24690
rect 6041 -24724 6069 -24690
rect 6107 -24724 6109 -24690
rect 6109 -24724 6141 -24690
rect 6179 -24724 6211 -24690
rect 6211 -24724 6213 -24690
rect 6251 -24724 6279 -24690
rect 6279 -24724 6285 -24690
rect 6323 -24724 6347 -24690
rect 6347 -24724 6357 -24690
rect 6981 -24724 6991 -24690
rect 6991 -24724 7015 -24690
rect 7053 -24724 7059 -24690
rect 7059 -24724 7087 -24690
rect 7125 -24724 7127 -24690
rect 7127 -24724 7159 -24690
rect 7197 -24724 7229 -24690
rect 7229 -24724 7231 -24690
rect 7269 -24724 7297 -24690
rect 7297 -24724 7303 -24690
rect 7341 -24724 7365 -24690
rect 7365 -24724 7375 -24690
rect 7999 -24724 8009 -24690
rect 8009 -24724 8033 -24690
rect 8071 -24724 8077 -24690
rect 8077 -24724 8105 -24690
rect 8143 -24724 8145 -24690
rect 8145 -24724 8177 -24690
rect 8215 -24724 8247 -24690
rect 8247 -24724 8249 -24690
rect 8287 -24724 8315 -24690
rect 8315 -24724 8321 -24690
rect 8359 -24724 8383 -24690
rect 8383 -24724 8393 -24690
rect 9017 -24724 9027 -24690
rect 9027 -24724 9051 -24690
rect 9089 -24724 9095 -24690
rect 9095 -24724 9123 -24690
rect 9161 -24724 9163 -24690
rect 9163 -24724 9195 -24690
rect 9233 -24724 9265 -24690
rect 9265 -24724 9267 -24690
rect 9305 -24724 9333 -24690
rect 9333 -24724 9339 -24690
rect 9377 -24724 9401 -24690
rect 9401 -24724 9411 -24690
rect 10035 -24724 10045 -24690
rect 10045 -24724 10069 -24690
rect 10107 -24724 10113 -24690
rect 10113 -24724 10141 -24690
rect 10179 -24724 10181 -24690
rect 10181 -24724 10213 -24690
rect 10251 -24724 10283 -24690
rect 10283 -24724 10285 -24690
rect 10323 -24724 10351 -24690
rect 10351 -24724 10357 -24690
rect 10395 -24724 10419 -24690
rect 10419 -24724 10429 -24690
rect 11053 -24724 11063 -24690
rect 11063 -24724 11087 -24690
rect 11125 -24724 11131 -24690
rect 11131 -24724 11159 -24690
rect 11197 -24724 11199 -24690
rect 11199 -24724 11231 -24690
rect 11269 -24724 11301 -24690
rect 11301 -24724 11303 -24690
rect 11341 -24724 11369 -24690
rect 11369 -24724 11375 -24690
rect 11413 -24724 11437 -24690
rect 11437 -24724 11447 -24690
rect 12071 -24724 12081 -24690
rect 12081 -24724 12105 -24690
rect 12143 -24724 12149 -24690
rect 12149 -24724 12177 -24690
rect 12215 -24724 12217 -24690
rect 12217 -24724 12249 -24690
rect 12287 -24724 12319 -24690
rect 12319 -24724 12321 -24690
rect 12359 -24724 12387 -24690
rect 12387 -24724 12393 -24690
rect 12431 -24724 12455 -24690
rect 12455 -24724 12465 -24690
rect 13089 -24724 13099 -24690
rect 13099 -24724 13123 -24690
rect 13161 -24724 13167 -24690
rect 13167 -24724 13195 -24690
rect 13233 -24724 13235 -24690
rect 13235 -24724 13267 -24690
rect 13305 -24724 13337 -24690
rect 13337 -24724 13339 -24690
rect 13377 -24724 13405 -24690
rect 13405 -24724 13411 -24690
rect 13449 -24724 13473 -24690
rect 13473 -24724 13483 -24690
rect 14107 -24724 14117 -24690
rect 14117 -24724 14141 -24690
rect 14179 -24724 14185 -24690
rect 14185 -24724 14213 -24690
rect 14251 -24724 14253 -24690
rect 14253 -24724 14285 -24690
rect 14323 -24724 14355 -24690
rect 14355 -24724 14357 -24690
rect 14395 -24724 14423 -24690
rect 14423 -24724 14429 -24690
rect 14467 -24724 14491 -24690
rect 14491 -24724 14501 -24690
rect 15125 -24724 15135 -24690
rect 15135 -24724 15159 -24690
rect 15197 -24724 15203 -24690
rect 15203 -24724 15231 -24690
rect 15269 -24724 15271 -24690
rect 15271 -24724 15303 -24690
rect 15341 -24724 15373 -24690
rect 15373 -24724 15375 -24690
rect 15413 -24724 15441 -24690
rect 15441 -24724 15447 -24690
rect 15485 -24724 15509 -24690
rect 15509 -24724 15519 -24690
rect 16143 -24724 16153 -24690
rect 16153 -24724 16177 -24690
rect 16215 -24724 16221 -24690
rect 16221 -24724 16249 -24690
rect 16287 -24724 16289 -24690
rect 16289 -24724 16321 -24690
rect 16359 -24724 16391 -24690
rect 16391 -24724 16393 -24690
rect 16431 -24724 16459 -24690
rect 16459 -24724 16465 -24690
rect 16503 -24724 16527 -24690
rect 16527 -24724 16537 -24690
rect 17161 -24724 17171 -24690
rect 17171 -24724 17195 -24690
rect 17233 -24724 17239 -24690
rect 17239 -24724 17267 -24690
rect 17305 -24724 17307 -24690
rect 17307 -24724 17339 -24690
rect 17377 -24724 17409 -24690
rect 17409 -24724 17411 -24690
rect 17449 -24724 17477 -24690
rect 17477 -24724 17483 -24690
rect 17521 -24724 17545 -24690
rect 17545 -24724 17555 -24690
rect 18179 -24724 18189 -24690
rect 18189 -24724 18213 -24690
rect 18251 -24724 18257 -24690
rect 18257 -24724 18285 -24690
rect 18323 -24724 18325 -24690
rect 18325 -24724 18357 -24690
rect 18395 -24724 18427 -24690
rect 18427 -24724 18429 -24690
rect 18467 -24724 18495 -24690
rect 18495 -24724 18501 -24690
rect 18539 -24724 18563 -24690
rect 18563 -24724 18573 -24690
rect 19197 -24724 19207 -24690
rect 19207 -24724 19231 -24690
rect 19269 -24724 19275 -24690
rect 19275 -24724 19303 -24690
rect 19341 -24724 19343 -24690
rect 19343 -24724 19375 -24690
rect 19413 -24724 19445 -24690
rect 19445 -24724 19447 -24690
rect 19485 -24724 19513 -24690
rect 19513 -24724 19519 -24690
rect 19557 -24724 19581 -24690
rect 19581 -24724 19591 -24690
rect 20215 -24724 20225 -24690
rect 20225 -24724 20249 -24690
rect 20287 -24724 20293 -24690
rect 20293 -24724 20321 -24690
rect 20359 -24724 20361 -24690
rect 20361 -24724 20393 -24690
rect 20431 -24724 20463 -24690
rect 20463 -24724 20465 -24690
rect 20503 -24724 20531 -24690
rect 20531 -24724 20537 -24690
rect 20575 -24724 20599 -24690
rect 20599 -24724 20609 -24690
rect 21233 -24724 21243 -24690
rect 21243 -24724 21267 -24690
rect 21305 -24724 21311 -24690
rect 21311 -24724 21339 -24690
rect 21377 -24724 21379 -24690
rect 21379 -24724 21411 -24690
rect 21449 -24724 21481 -24690
rect 21481 -24724 21483 -24690
rect 21521 -24724 21549 -24690
rect 21549 -24724 21555 -24690
rect 21593 -24724 21617 -24690
rect 21617 -24724 21627 -24690
rect 22251 -24724 22261 -24690
rect 22261 -24724 22285 -24690
rect 22323 -24724 22329 -24690
rect 22329 -24724 22357 -24690
rect 22395 -24724 22397 -24690
rect 22397 -24724 22429 -24690
rect 22467 -24724 22499 -24690
rect 22499 -24724 22501 -24690
rect 22539 -24724 22567 -24690
rect 22567 -24724 22573 -24690
rect 22611 -24724 22635 -24690
rect 22635 -24724 22645 -24690
rect -12289 -24793 -12255 -24763
rect -12289 -24797 -12255 -24793
rect -12289 -24861 -12255 -24835
rect -12289 -24869 -12255 -24861
rect -12289 -24929 -12255 -24907
rect -12289 -24941 -12255 -24929
rect -12289 -24997 -12255 -24979
rect -12289 -25013 -12255 -24997
rect -12289 -25065 -12255 -25051
rect -12289 -25085 -12255 -25065
rect 24855 -24725 24889 -24691
rect 24855 -24793 24889 -24763
rect 24855 -24797 24889 -24793
rect 24855 -24861 24889 -24835
rect 24855 -24869 24889 -24861
rect 24855 -24929 24889 -24907
rect 24855 -24941 24889 -24929
rect 24855 -24997 24889 -24979
rect 24855 -25013 24889 -24997
rect -9077 -25080 -9067 -25046
rect -9067 -25080 -9043 -25046
rect -9005 -25080 -8999 -25046
rect -8999 -25080 -8971 -25046
rect -8933 -25080 -8931 -25046
rect -8931 -25080 -8899 -25046
rect -8861 -25080 -8829 -25046
rect -8829 -25080 -8827 -25046
rect -8789 -25080 -8761 -25046
rect -8761 -25080 -8755 -25046
rect -8717 -25080 -8693 -25046
rect -8693 -25080 -8683 -25046
rect -8059 -25080 -8049 -25046
rect -8049 -25080 -8025 -25046
rect -7987 -25080 -7981 -25046
rect -7981 -25080 -7953 -25046
rect -7915 -25080 -7913 -25046
rect -7913 -25080 -7881 -25046
rect -7843 -25080 -7811 -25046
rect -7811 -25080 -7809 -25046
rect -7771 -25080 -7743 -25046
rect -7743 -25080 -7737 -25046
rect -7699 -25080 -7675 -25046
rect -7675 -25080 -7665 -25046
rect -7041 -25080 -7031 -25046
rect -7031 -25080 -7007 -25046
rect -6969 -25080 -6963 -25046
rect -6963 -25080 -6935 -25046
rect -6897 -25080 -6895 -25046
rect -6895 -25080 -6863 -25046
rect -6825 -25080 -6793 -25046
rect -6793 -25080 -6791 -25046
rect -6753 -25080 -6725 -25046
rect -6725 -25080 -6719 -25046
rect -6681 -25080 -6657 -25046
rect -6657 -25080 -6647 -25046
rect -6023 -25080 -6013 -25046
rect -6013 -25080 -5989 -25046
rect -5951 -25080 -5945 -25046
rect -5945 -25080 -5917 -25046
rect -5879 -25080 -5877 -25046
rect -5877 -25080 -5845 -25046
rect -5807 -25080 -5775 -25046
rect -5775 -25080 -5773 -25046
rect -5735 -25080 -5707 -25046
rect -5707 -25080 -5701 -25046
rect -5663 -25080 -5639 -25046
rect -5639 -25080 -5629 -25046
rect -5005 -25080 -4995 -25046
rect -4995 -25080 -4971 -25046
rect -4933 -25080 -4927 -25046
rect -4927 -25080 -4899 -25046
rect -4861 -25080 -4859 -25046
rect -4859 -25080 -4827 -25046
rect -4789 -25080 -4757 -25046
rect -4757 -25080 -4755 -25046
rect -4717 -25080 -4689 -25046
rect -4689 -25080 -4683 -25046
rect -4645 -25080 -4621 -25046
rect -4621 -25080 -4611 -25046
rect -3987 -25080 -3977 -25046
rect -3977 -25080 -3953 -25046
rect -3915 -25080 -3909 -25046
rect -3909 -25080 -3881 -25046
rect -3843 -25080 -3841 -25046
rect -3841 -25080 -3809 -25046
rect -3771 -25080 -3739 -25046
rect -3739 -25080 -3737 -25046
rect -3699 -25080 -3671 -25046
rect -3671 -25080 -3665 -25046
rect -3627 -25080 -3603 -25046
rect -3603 -25080 -3593 -25046
rect -2263 -25076 -2229 -25042
rect -1965 -25076 -1931 -25042
rect -1667 -25076 -1633 -25042
rect -1369 -25076 -1335 -25042
rect -1071 -25076 -1037 -25042
rect -773 -25076 -739 -25042
rect -475 -25076 -441 -25042
rect -177 -25076 -143 -25042
rect 121 -25076 155 -25042
rect 419 -25076 453 -25042
rect 717 -25076 751 -25042
rect -12289 -25133 -12255 -25123
rect -12289 -25157 -12255 -25133
rect 24855 -25065 24889 -25051
rect 24855 -25085 24889 -25065
rect -12289 -25201 -12255 -25195
rect -12289 -25229 -12255 -25201
rect -12289 -25269 -12255 -25267
rect -12289 -25301 -12255 -25269
rect -12289 -25371 -12255 -25339
rect -12289 -25373 -12255 -25371
rect -12289 -25439 -12255 -25411
rect -12289 -25445 -12255 -25439
rect -12289 -25507 -12255 -25483
rect -12289 -25517 -12255 -25507
rect -12289 -25575 -12255 -25555
rect -12289 -25589 -12255 -25575
rect -12289 -25643 -12255 -25627
rect -12289 -25661 -12255 -25643
rect -12289 -25711 -12255 -25699
rect -12289 -25733 -12255 -25711
rect -9406 -25163 -9372 -25149
rect -9406 -25183 -9372 -25163
rect -9406 -25231 -9372 -25221
rect -9406 -25255 -9372 -25231
rect -9406 -25299 -9372 -25293
rect -9406 -25327 -9372 -25299
rect -9406 -25367 -9372 -25365
rect -9406 -25399 -9372 -25367
rect -9406 -25469 -9372 -25437
rect -9406 -25471 -9372 -25469
rect -9406 -25537 -9372 -25509
rect -9406 -25543 -9372 -25537
rect -9406 -25605 -9372 -25581
rect -9406 -25615 -9372 -25605
rect -9406 -25673 -9372 -25653
rect -9406 -25687 -9372 -25673
rect -8388 -25163 -8354 -25149
rect -8388 -25183 -8354 -25163
rect -8388 -25231 -8354 -25221
rect -8388 -25255 -8354 -25231
rect -8388 -25299 -8354 -25293
rect -8388 -25327 -8354 -25299
rect -8388 -25367 -8354 -25365
rect -8388 -25399 -8354 -25367
rect -8388 -25469 -8354 -25437
rect -8388 -25471 -8354 -25469
rect -8388 -25537 -8354 -25509
rect -8388 -25543 -8354 -25537
rect -8388 -25605 -8354 -25581
rect -8388 -25615 -8354 -25605
rect -8388 -25673 -8354 -25653
rect -8388 -25687 -8354 -25673
rect -7370 -25163 -7336 -25149
rect -7370 -25183 -7336 -25163
rect -7370 -25231 -7336 -25221
rect -7370 -25255 -7336 -25231
rect -7370 -25299 -7336 -25293
rect -7370 -25327 -7336 -25299
rect -7370 -25367 -7336 -25365
rect -7370 -25399 -7336 -25367
rect -7370 -25469 -7336 -25437
rect -7370 -25471 -7336 -25469
rect -7370 -25537 -7336 -25509
rect -7370 -25543 -7336 -25537
rect -7370 -25605 -7336 -25581
rect -7370 -25615 -7336 -25605
rect -7370 -25673 -7336 -25653
rect -7370 -25687 -7336 -25673
rect -6352 -25163 -6318 -25149
rect -6352 -25183 -6318 -25163
rect -6352 -25231 -6318 -25221
rect -6352 -25255 -6318 -25231
rect -6352 -25299 -6318 -25293
rect -6352 -25327 -6318 -25299
rect -6352 -25367 -6318 -25365
rect -6352 -25399 -6318 -25367
rect -6352 -25469 -6318 -25437
rect -6352 -25471 -6318 -25469
rect -6352 -25537 -6318 -25509
rect -6352 -25543 -6318 -25537
rect -6352 -25605 -6318 -25581
rect -6352 -25615 -6318 -25605
rect -6352 -25673 -6318 -25653
rect -6352 -25687 -6318 -25673
rect -5334 -25163 -5300 -25149
rect -5334 -25183 -5300 -25163
rect -5334 -25231 -5300 -25221
rect -5334 -25255 -5300 -25231
rect -5334 -25299 -5300 -25293
rect -5334 -25327 -5300 -25299
rect -5334 -25367 -5300 -25365
rect -5334 -25399 -5300 -25367
rect -5334 -25469 -5300 -25437
rect -5334 -25471 -5300 -25469
rect -5334 -25537 -5300 -25509
rect -5334 -25543 -5300 -25537
rect -5334 -25605 -5300 -25581
rect -5334 -25615 -5300 -25605
rect -5334 -25673 -5300 -25653
rect -5334 -25687 -5300 -25673
rect -4316 -25163 -4282 -25149
rect -4316 -25183 -4282 -25163
rect -4316 -25231 -4282 -25221
rect -4316 -25255 -4282 -25231
rect -4316 -25299 -4282 -25293
rect -4316 -25327 -4282 -25299
rect -4316 -25367 -4282 -25365
rect -4316 -25399 -4282 -25367
rect -4316 -25469 -4282 -25437
rect -4316 -25471 -4282 -25469
rect -4316 -25537 -4282 -25509
rect -4316 -25543 -4282 -25537
rect -4316 -25605 -4282 -25581
rect -4316 -25615 -4282 -25605
rect -4316 -25673 -4282 -25653
rect -4316 -25687 -4282 -25673
rect -3298 -25163 -3264 -25149
rect -3298 -25183 -3264 -25163
rect -3298 -25231 -3264 -25221
rect -3298 -25255 -3264 -25231
rect -3298 -25299 -3264 -25293
rect -3298 -25327 -3264 -25299
rect -3298 -25367 -3264 -25365
rect -3298 -25399 -3264 -25367
rect -3298 -25469 -3264 -25437
rect -3298 -25471 -3264 -25469
rect -3298 -25537 -3264 -25509
rect -3298 -25543 -3264 -25537
rect -3298 -25605 -3264 -25581
rect -3298 -25615 -3264 -25605
rect -3298 -25673 -3264 -25653
rect -3298 -25687 -3264 -25673
rect -2412 -25159 -2378 -25145
rect -2412 -25179 -2378 -25159
rect -2412 -25227 -2378 -25217
rect -2412 -25251 -2378 -25227
rect -2412 -25295 -2378 -25289
rect -2412 -25323 -2378 -25295
rect -2412 -25363 -2378 -25361
rect -2412 -25395 -2378 -25363
rect -2412 -25465 -2378 -25433
rect -2412 -25467 -2378 -25465
rect -2412 -25533 -2378 -25505
rect -2412 -25539 -2378 -25533
rect -2412 -25601 -2378 -25577
rect -2412 -25611 -2378 -25601
rect -2412 -25669 -2378 -25649
rect -2412 -25683 -2378 -25669
rect -2114 -25159 -2080 -25145
rect -2114 -25179 -2080 -25159
rect -2114 -25227 -2080 -25217
rect -2114 -25251 -2080 -25227
rect -2114 -25295 -2080 -25289
rect -2114 -25323 -2080 -25295
rect -2114 -25363 -2080 -25361
rect -2114 -25395 -2080 -25363
rect -2114 -25465 -2080 -25433
rect -2114 -25467 -2080 -25465
rect -2114 -25533 -2080 -25505
rect -2114 -25539 -2080 -25533
rect -2114 -25601 -2080 -25577
rect -2114 -25611 -2080 -25601
rect -2114 -25669 -2080 -25649
rect -2114 -25683 -2080 -25669
rect -1816 -25159 -1782 -25145
rect -1816 -25179 -1782 -25159
rect -1816 -25227 -1782 -25217
rect -1816 -25251 -1782 -25227
rect -1816 -25295 -1782 -25289
rect -1816 -25323 -1782 -25295
rect -1816 -25363 -1782 -25361
rect -1816 -25395 -1782 -25363
rect -1816 -25465 -1782 -25433
rect -1816 -25467 -1782 -25465
rect -1816 -25533 -1782 -25505
rect -1816 -25539 -1782 -25533
rect -1816 -25601 -1782 -25577
rect -1816 -25611 -1782 -25601
rect -1816 -25669 -1782 -25649
rect -1816 -25683 -1782 -25669
rect -1518 -25159 -1484 -25145
rect -1518 -25179 -1484 -25159
rect -1518 -25227 -1484 -25217
rect -1518 -25251 -1484 -25227
rect -1518 -25295 -1484 -25289
rect -1518 -25323 -1484 -25295
rect -1518 -25363 -1484 -25361
rect -1518 -25395 -1484 -25363
rect -1518 -25465 -1484 -25433
rect -1518 -25467 -1484 -25465
rect -1518 -25533 -1484 -25505
rect -1518 -25539 -1484 -25533
rect -1518 -25601 -1484 -25577
rect -1518 -25611 -1484 -25601
rect -1518 -25669 -1484 -25649
rect -1518 -25683 -1484 -25669
rect -1220 -25159 -1186 -25145
rect -1220 -25179 -1186 -25159
rect -1220 -25227 -1186 -25217
rect -1220 -25251 -1186 -25227
rect -1220 -25295 -1186 -25289
rect -1220 -25323 -1186 -25295
rect -1220 -25363 -1186 -25361
rect -1220 -25395 -1186 -25363
rect -1220 -25465 -1186 -25433
rect -1220 -25467 -1186 -25465
rect -1220 -25533 -1186 -25505
rect -1220 -25539 -1186 -25533
rect -1220 -25601 -1186 -25577
rect -1220 -25611 -1186 -25601
rect -1220 -25669 -1186 -25649
rect -1220 -25683 -1186 -25669
rect -922 -25159 -888 -25145
rect -922 -25179 -888 -25159
rect -922 -25227 -888 -25217
rect -922 -25251 -888 -25227
rect -922 -25295 -888 -25289
rect -922 -25323 -888 -25295
rect -922 -25363 -888 -25361
rect -922 -25395 -888 -25363
rect -922 -25465 -888 -25433
rect -922 -25467 -888 -25465
rect -922 -25533 -888 -25505
rect -922 -25539 -888 -25533
rect -922 -25601 -888 -25577
rect -922 -25611 -888 -25601
rect -922 -25669 -888 -25649
rect -922 -25683 -888 -25669
rect -624 -25159 -590 -25145
rect -624 -25179 -590 -25159
rect -624 -25227 -590 -25217
rect -624 -25251 -590 -25227
rect -624 -25295 -590 -25289
rect -624 -25323 -590 -25295
rect -624 -25363 -590 -25361
rect -624 -25395 -590 -25363
rect -624 -25465 -590 -25433
rect -624 -25467 -590 -25465
rect -624 -25533 -590 -25505
rect -624 -25539 -590 -25533
rect -624 -25601 -590 -25577
rect -624 -25611 -590 -25601
rect -624 -25669 -590 -25649
rect -624 -25683 -590 -25669
rect -326 -25159 -292 -25145
rect -326 -25179 -292 -25159
rect -326 -25227 -292 -25217
rect -326 -25251 -292 -25227
rect -326 -25295 -292 -25289
rect -326 -25323 -292 -25295
rect -326 -25363 -292 -25361
rect -326 -25395 -292 -25363
rect -326 -25465 -292 -25433
rect -326 -25467 -292 -25465
rect -326 -25533 -292 -25505
rect -326 -25539 -292 -25533
rect -326 -25601 -292 -25577
rect -326 -25611 -292 -25601
rect -326 -25669 -292 -25649
rect -326 -25683 -292 -25669
rect -28 -25159 6 -25145
rect -28 -25179 6 -25159
rect -28 -25227 6 -25217
rect -28 -25251 6 -25227
rect -28 -25295 6 -25289
rect -28 -25323 6 -25295
rect -28 -25363 6 -25361
rect -28 -25395 6 -25363
rect -28 -25465 6 -25433
rect -28 -25467 6 -25465
rect -28 -25533 6 -25505
rect -28 -25539 6 -25533
rect -28 -25601 6 -25577
rect -28 -25611 6 -25601
rect -28 -25669 6 -25649
rect -28 -25683 6 -25669
rect 270 -25159 304 -25145
rect 270 -25179 304 -25159
rect 270 -25227 304 -25217
rect 270 -25251 304 -25227
rect 270 -25295 304 -25289
rect 270 -25323 304 -25295
rect 270 -25363 304 -25361
rect 270 -25395 304 -25363
rect 270 -25465 304 -25433
rect 270 -25467 304 -25465
rect 270 -25533 304 -25505
rect 270 -25539 304 -25533
rect 270 -25601 304 -25577
rect 270 -25611 304 -25601
rect 270 -25669 304 -25649
rect 270 -25683 304 -25669
rect 568 -25159 602 -25145
rect 568 -25179 602 -25159
rect 568 -25227 602 -25217
rect 568 -25251 602 -25227
rect 568 -25295 602 -25289
rect 568 -25323 602 -25295
rect 568 -25363 602 -25361
rect 568 -25395 602 -25363
rect 568 -25465 602 -25433
rect 568 -25467 602 -25465
rect 568 -25533 602 -25505
rect 568 -25539 602 -25533
rect 568 -25601 602 -25577
rect 568 -25611 602 -25601
rect 568 -25669 602 -25649
rect 568 -25683 602 -25669
rect 866 -25159 900 -25145
rect 866 -25179 900 -25159
rect 24855 -25133 24889 -25123
rect 24855 -25157 24889 -25133
rect 866 -25227 900 -25217
rect 866 -25251 900 -25227
rect 2909 -25246 2919 -25212
rect 2919 -25246 2943 -25212
rect 2981 -25246 2987 -25212
rect 2987 -25246 3015 -25212
rect 3053 -25246 3055 -25212
rect 3055 -25246 3087 -25212
rect 3125 -25246 3157 -25212
rect 3157 -25246 3159 -25212
rect 3197 -25246 3225 -25212
rect 3225 -25246 3231 -25212
rect 3269 -25246 3293 -25212
rect 3293 -25246 3303 -25212
rect 3927 -25246 3937 -25212
rect 3937 -25246 3961 -25212
rect 3999 -25246 4005 -25212
rect 4005 -25246 4033 -25212
rect 4071 -25246 4073 -25212
rect 4073 -25246 4105 -25212
rect 4143 -25246 4175 -25212
rect 4175 -25246 4177 -25212
rect 4215 -25246 4243 -25212
rect 4243 -25246 4249 -25212
rect 4287 -25246 4311 -25212
rect 4311 -25246 4321 -25212
rect 4945 -25246 4955 -25212
rect 4955 -25246 4979 -25212
rect 5017 -25246 5023 -25212
rect 5023 -25246 5051 -25212
rect 5089 -25246 5091 -25212
rect 5091 -25246 5123 -25212
rect 5161 -25246 5193 -25212
rect 5193 -25246 5195 -25212
rect 5233 -25246 5261 -25212
rect 5261 -25246 5267 -25212
rect 5305 -25246 5329 -25212
rect 5329 -25246 5339 -25212
rect 5963 -25246 5973 -25212
rect 5973 -25246 5997 -25212
rect 6035 -25246 6041 -25212
rect 6041 -25246 6069 -25212
rect 6107 -25246 6109 -25212
rect 6109 -25246 6141 -25212
rect 6179 -25246 6211 -25212
rect 6211 -25246 6213 -25212
rect 6251 -25246 6279 -25212
rect 6279 -25246 6285 -25212
rect 6323 -25246 6347 -25212
rect 6347 -25246 6357 -25212
rect 6981 -25246 6991 -25212
rect 6991 -25246 7015 -25212
rect 7053 -25246 7059 -25212
rect 7059 -25246 7087 -25212
rect 7125 -25246 7127 -25212
rect 7127 -25246 7159 -25212
rect 7197 -25246 7229 -25212
rect 7229 -25246 7231 -25212
rect 7269 -25246 7297 -25212
rect 7297 -25246 7303 -25212
rect 7341 -25246 7365 -25212
rect 7365 -25246 7375 -25212
rect 7999 -25246 8009 -25212
rect 8009 -25246 8033 -25212
rect 8071 -25246 8077 -25212
rect 8077 -25246 8105 -25212
rect 8143 -25246 8145 -25212
rect 8145 -25246 8177 -25212
rect 8215 -25246 8247 -25212
rect 8247 -25246 8249 -25212
rect 8287 -25246 8315 -25212
rect 8315 -25246 8321 -25212
rect 8359 -25246 8383 -25212
rect 8383 -25246 8393 -25212
rect 9017 -25246 9027 -25212
rect 9027 -25246 9051 -25212
rect 9089 -25246 9095 -25212
rect 9095 -25246 9123 -25212
rect 9161 -25246 9163 -25212
rect 9163 -25246 9195 -25212
rect 9233 -25246 9265 -25212
rect 9265 -25246 9267 -25212
rect 9305 -25246 9333 -25212
rect 9333 -25246 9339 -25212
rect 9377 -25246 9401 -25212
rect 9401 -25246 9411 -25212
rect 10035 -25246 10045 -25212
rect 10045 -25246 10069 -25212
rect 10107 -25246 10113 -25212
rect 10113 -25246 10141 -25212
rect 10179 -25246 10181 -25212
rect 10181 -25246 10213 -25212
rect 10251 -25246 10283 -25212
rect 10283 -25246 10285 -25212
rect 10323 -25246 10351 -25212
rect 10351 -25246 10357 -25212
rect 10395 -25246 10419 -25212
rect 10419 -25246 10429 -25212
rect 11053 -25246 11063 -25212
rect 11063 -25246 11087 -25212
rect 11125 -25246 11131 -25212
rect 11131 -25246 11159 -25212
rect 11197 -25246 11199 -25212
rect 11199 -25246 11231 -25212
rect 11269 -25246 11301 -25212
rect 11301 -25246 11303 -25212
rect 11341 -25246 11369 -25212
rect 11369 -25246 11375 -25212
rect 11413 -25246 11437 -25212
rect 11437 -25246 11447 -25212
rect 12071 -25246 12081 -25212
rect 12081 -25246 12105 -25212
rect 12143 -25246 12149 -25212
rect 12149 -25246 12177 -25212
rect 12215 -25246 12217 -25212
rect 12217 -25246 12249 -25212
rect 12287 -25246 12319 -25212
rect 12319 -25246 12321 -25212
rect 12359 -25246 12387 -25212
rect 12387 -25246 12393 -25212
rect 12431 -25246 12455 -25212
rect 12455 -25246 12465 -25212
rect 13089 -25246 13099 -25212
rect 13099 -25246 13123 -25212
rect 13161 -25246 13167 -25212
rect 13167 -25246 13195 -25212
rect 13233 -25246 13235 -25212
rect 13235 -25246 13267 -25212
rect 13305 -25246 13337 -25212
rect 13337 -25246 13339 -25212
rect 13377 -25246 13405 -25212
rect 13405 -25246 13411 -25212
rect 13449 -25246 13473 -25212
rect 13473 -25246 13483 -25212
rect 14107 -25246 14117 -25212
rect 14117 -25246 14141 -25212
rect 14179 -25246 14185 -25212
rect 14185 -25246 14213 -25212
rect 14251 -25246 14253 -25212
rect 14253 -25246 14285 -25212
rect 14323 -25246 14355 -25212
rect 14355 -25246 14357 -25212
rect 14395 -25246 14423 -25212
rect 14423 -25246 14429 -25212
rect 14467 -25246 14491 -25212
rect 14491 -25246 14501 -25212
rect 15125 -25246 15135 -25212
rect 15135 -25246 15159 -25212
rect 15197 -25246 15203 -25212
rect 15203 -25246 15231 -25212
rect 15269 -25246 15271 -25212
rect 15271 -25246 15303 -25212
rect 15341 -25246 15373 -25212
rect 15373 -25246 15375 -25212
rect 15413 -25246 15441 -25212
rect 15441 -25246 15447 -25212
rect 15485 -25246 15509 -25212
rect 15509 -25246 15519 -25212
rect 16143 -25246 16153 -25212
rect 16153 -25246 16177 -25212
rect 16215 -25246 16221 -25212
rect 16221 -25246 16249 -25212
rect 16287 -25246 16289 -25212
rect 16289 -25246 16321 -25212
rect 16359 -25246 16391 -25212
rect 16391 -25246 16393 -25212
rect 16431 -25246 16459 -25212
rect 16459 -25246 16465 -25212
rect 16503 -25246 16527 -25212
rect 16527 -25246 16537 -25212
rect 17161 -25246 17171 -25212
rect 17171 -25246 17195 -25212
rect 17233 -25246 17239 -25212
rect 17239 -25246 17267 -25212
rect 17305 -25246 17307 -25212
rect 17307 -25246 17339 -25212
rect 17377 -25246 17409 -25212
rect 17409 -25246 17411 -25212
rect 17449 -25246 17477 -25212
rect 17477 -25246 17483 -25212
rect 17521 -25246 17545 -25212
rect 17545 -25246 17555 -25212
rect 18179 -25246 18189 -25212
rect 18189 -25246 18213 -25212
rect 18251 -25246 18257 -25212
rect 18257 -25246 18285 -25212
rect 18323 -25246 18325 -25212
rect 18325 -25246 18357 -25212
rect 18395 -25246 18427 -25212
rect 18427 -25246 18429 -25212
rect 18467 -25246 18495 -25212
rect 18495 -25246 18501 -25212
rect 18539 -25246 18563 -25212
rect 18563 -25246 18573 -25212
rect 19197 -25246 19207 -25212
rect 19207 -25246 19231 -25212
rect 19269 -25246 19275 -25212
rect 19275 -25246 19303 -25212
rect 19341 -25246 19343 -25212
rect 19343 -25246 19375 -25212
rect 19413 -25246 19445 -25212
rect 19445 -25246 19447 -25212
rect 19485 -25246 19513 -25212
rect 19513 -25246 19519 -25212
rect 19557 -25246 19581 -25212
rect 19581 -25246 19591 -25212
rect 20215 -25246 20225 -25212
rect 20225 -25246 20249 -25212
rect 20287 -25246 20293 -25212
rect 20293 -25246 20321 -25212
rect 20359 -25246 20361 -25212
rect 20361 -25246 20393 -25212
rect 20431 -25246 20463 -25212
rect 20463 -25246 20465 -25212
rect 20503 -25246 20531 -25212
rect 20531 -25246 20537 -25212
rect 20575 -25246 20599 -25212
rect 20599 -25246 20609 -25212
rect 21233 -25246 21243 -25212
rect 21243 -25246 21267 -25212
rect 21305 -25246 21311 -25212
rect 21311 -25246 21339 -25212
rect 21377 -25246 21379 -25212
rect 21379 -25246 21411 -25212
rect 21449 -25246 21481 -25212
rect 21481 -25246 21483 -25212
rect 21521 -25246 21549 -25212
rect 21549 -25246 21555 -25212
rect 21593 -25246 21617 -25212
rect 21617 -25246 21627 -25212
rect 22251 -25246 22261 -25212
rect 22261 -25246 22285 -25212
rect 22323 -25246 22329 -25212
rect 22329 -25246 22357 -25212
rect 22395 -25246 22397 -25212
rect 22397 -25246 22429 -25212
rect 22467 -25246 22499 -25212
rect 22499 -25246 22501 -25212
rect 22539 -25246 22567 -25212
rect 22567 -25246 22573 -25212
rect 22611 -25246 22635 -25212
rect 22635 -25246 22645 -25212
rect 24855 -25201 24889 -25195
rect 24855 -25229 24889 -25201
rect 866 -25295 900 -25289
rect 866 -25323 900 -25295
rect 866 -25363 900 -25361
rect 866 -25395 900 -25363
rect 866 -25465 900 -25433
rect 866 -25467 900 -25465
rect 866 -25533 900 -25505
rect 866 -25539 900 -25533
rect 866 -25601 900 -25577
rect 866 -25611 900 -25601
rect 866 -25669 900 -25649
rect 866 -25683 900 -25669
rect 2580 -25329 2614 -25315
rect 2580 -25349 2614 -25329
rect 2580 -25397 2614 -25387
rect 2580 -25421 2614 -25397
rect 2580 -25465 2614 -25459
rect 2580 -25493 2614 -25465
rect 2580 -25533 2614 -25531
rect 2580 -25565 2614 -25533
rect 2580 -25635 2614 -25603
rect 2580 -25637 2614 -25635
rect 2580 -25703 2614 -25675
rect 2580 -25709 2614 -25703
rect -12289 -25779 -12255 -25771
rect -12289 -25805 -12255 -25779
rect -9077 -25790 -9067 -25756
rect -9067 -25790 -9043 -25756
rect -9005 -25790 -8999 -25756
rect -8999 -25790 -8971 -25756
rect -8933 -25790 -8931 -25756
rect -8931 -25790 -8899 -25756
rect -8861 -25790 -8829 -25756
rect -8829 -25790 -8827 -25756
rect -8789 -25790 -8761 -25756
rect -8761 -25790 -8755 -25756
rect -8717 -25790 -8693 -25756
rect -8693 -25790 -8683 -25756
rect -8059 -25790 -8049 -25756
rect -8049 -25790 -8025 -25756
rect -7987 -25790 -7981 -25756
rect -7981 -25790 -7953 -25756
rect -7915 -25790 -7913 -25756
rect -7913 -25790 -7881 -25756
rect -7843 -25790 -7811 -25756
rect -7811 -25790 -7809 -25756
rect -7771 -25790 -7743 -25756
rect -7743 -25790 -7737 -25756
rect -7699 -25790 -7675 -25756
rect -7675 -25790 -7665 -25756
rect -7041 -25790 -7031 -25756
rect -7031 -25790 -7007 -25756
rect -6969 -25790 -6963 -25756
rect -6963 -25790 -6935 -25756
rect -6897 -25790 -6895 -25756
rect -6895 -25790 -6863 -25756
rect -6825 -25790 -6793 -25756
rect -6793 -25790 -6791 -25756
rect -6753 -25790 -6725 -25756
rect -6725 -25790 -6719 -25756
rect -6681 -25790 -6657 -25756
rect -6657 -25790 -6647 -25756
rect -6023 -25790 -6013 -25756
rect -6013 -25790 -5989 -25756
rect -5951 -25790 -5945 -25756
rect -5945 -25790 -5917 -25756
rect -5879 -25790 -5877 -25756
rect -5877 -25790 -5845 -25756
rect -5807 -25790 -5775 -25756
rect -5775 -25790 -5773 -25756
rect -5735 -25790 -5707 -25756
rect -5707 -25790 -5701 -25756
rect -5663 -25790 -5639 -25756
rect -5639 -25790 -5629 -25756
rect -5005 -25790 -4995 -25756
rect -4995 -25790 -4971 -25756
rect -4933 -25790 -4927 -25756
rect -4927 -25790 -4899 -25756
rect -4861 -25790 -4859 -25756
rect -4859 -25790 -4827 -25756
rect -4789 -25790 -4757 -25756
rect -4757 -25790 -4755 -25756
rect -4717 -25790 -4689 -25756
rect -4689 -25790 -4683 -25756
rect -4645 -25790 -4621 -25756
rect -4621 -25790 -4611 -25756
rect -3987 -25790 -3977 -25756
rect -3977 -25790 -3953 -25756
rect -3915 -25790 -3909 -25756
rect -3909 -25790 -3881 -25756
rect -3843 -25790 -3841 -25756
rect -3841 -25790 -3809 -25756
rect -3771 -25790 -3739 -25756
rect -3739 -25790 -3737 -25756
rect -3699 -25790 -3671 -25756
rect -3671 -25790 -3665 -25756
rect -3627 -25790 -3603 -25756
rect -3603 -25790 -3593 -25756
rect -2263 -25786 -2229 -25752
rect -1965 -25786 -1931 -25752
rect -1667 -25786 -1633 -25752
rect -1369 -25786 -1335 -25752
rect -1071 -25786 -1037 -25752
rect -773 -25786 -739 -25752
rect -475 -25786 -441 -25752
rect -177 -25786 -143 -25752
rect 121 -25786 155 -25752
rect 419 -25786 453 -25752
rect 717 -25786 751 -25752
rect 2580 -25771 2614 -25747
rect 2580 -25781 2614 -25771
rect -12289 -25847 -12255 -25843
rect -12289 -25877 -12255 -25847
rect 2580 -25839 2614 -25819
rect 3598 -25329 3632 -25315
rect 3598 -25349 3632 -25329
rect 3598 -25397 3632 -25387
rect 3598 -25421 3632 -25397
rect 3598 -25465 3632 -25459
rect 3598 -25493 3632 -25465
rect 3598 -25533 3632 -25531
rect 3598 -25565 3632 -25533
rect 3598 -25635 3632 -25603
rect 3598 -25637 3632 -25635
rect 3598 -25703 3632 -25675
rect 3598 -25709 3632 -25703
rect 3598 -25771 3632 -25747
rect 3598 -25781 3632 -25771
rect 2580 -25853 2614 -25839
rect 3598 -25839 3632 -25819
rect 4616 -25329 4650 -25315
rect 4616 -25349 4650 -25329
rect 4616 -25397 4650 -25387
rect 4616 -25421 4650 -25397
rect 4616 -25465 4650 -25459
rect 4616 -25493 4650 -25465
rect 4616 -25533 4650 -25531
rect 4616 -25565 4650 -25533
rect 4616 -25635 4650 -25603
rect 4616 -25637 4650 -25635
rect 4616 -25703 4650 -25675
rect 4616 -25709 4650 -25703
rect 4616 -25771 4650 -25747
rect 4616 -25781 4650 -25771
rect 3598 -25853 3632 -25839
rect 4616 -25839 4650 -25819
rect 4616 -25853 4650 -25839
rect 5634 -25329 5668 -25315
rect 5634 -25349 5668 -25329
rect 5634 -25397 5668 -25387
rect 5634 -25421 5668 -25397
rect 5634 -25465 5668 -25459
rect 5634 -25493 5668 -25465
rect 5634 -25533 5668 -25531
rect 5634 -25565 5668 -25533
rect 5634 -25635 5668 -25603
rect 5634 -25637 5668 -25635
rect 5634 -25703 5668 -25675
rect 5634 -25709 5668 -25703
rect 5634 -25771 5668 -25747
rect 5634 -25781 5668 -25771
rect 5634 -25839 5668 -25819
rect 5634 -25853 5668 -25839
rect 6652 -25329 6686 -25315
rect 6652 -25349 6686 -25329
rect 6652 -25397 6686 -25387
rect 6652 -25421 6686 -25397
rect 6652 -25465 6686 -25459
rect 6652 -25493 6686 -25465
rect 6652 -25533 6686 -25531
rect 6652 -25565 6686 -25533
rect 6652 -25635 6686 -25603
rect 6652 -25637 6686 -25635
rect 6652 -25703 6686 -25675
rect 6652 -25709 6686 -25703
rect 6652 -25771 6686 -25747
rect 6652 -25781 6686 -25771
rect 6652 -25839 6686 -25819
rect 7670 -25329 7704 -25315
rect 7670 -25349 7704 -25329
rect 7670 -25397 7704 -25387
rect 7670 -25421 7704 -25397
rect 7670 -25465 7704 -25459
rect 7670 -25493 7704 -25465
rect 7670 -25533 7704 -25531
rect 7670 -25565 7704 -25533
rect 7670 -25635 7704 -25603
rect 7670 -25637 7704 -25635
rect 7670 -25703 7704 -25675
rect 7670 -25709 7704 -25703
rect 7670 -25771 7704 -25747
rect 7670 -25781 7704 -25771
rect 6652 -25853 6686 -25839
rect 7670 -25839 7704 -25819
rect 8688 -25329 8722 -25315
rect 8688 -25349 8722 -25329
rect 8688 -25397 8722 -25387
rect 8688 -25421 8722 -25397
rect 8688 -25465 8722 -25459
rect 8688 -25493 8722 -25465
rect 8688 -25533 8722 -25531
rect 8688 -25565 8722 -25533
rect 8688 -25635 8722 -25603
rect 8688 -25637 8722 -25635
rect 8688 -25703 8722 -25675
rect 8688 -25709 8722 -25703
rect 8688 -25771 8722 -25747
rect 8688 -25781 8722 -25771
rect 7670 -25853 7704 -25839
rect 8688 -25839 8722 -25819
rect 8688 -25853 8722 -25839
rect 9706 -25329 9740 -25315
rect 9706 -25349 9740 -25329
rect 9706 -25397 9740 -25387
rect 9706 -25421 9740 -25397
rect 9706 -25465 9740 -25459
rect 9706 -25493 9740 -25465
rect 9706 -25533 9740 -25531
rect 9706 -25565 9740 -25533
rect 9706 -25635 9740 -25603
rect 9706 -25637 9740 -25635
rect 9706 -25703 9740 -25675
rect 9706 -25709 9740 -25703
rect 9706 -25771 9740 -25747
rect 9706 -25781 9740 -25771
rect 9706 -25839 9740 -25819
rect 9706 -25853 9740 -25839
rect 10724 -25329 10758 -25315
rect 10724 -25349 10758 -25329
rect 10724 -25397 10758 -25387
rect 10724 -25421 10758 -25397
rect 10724 -25465 10758 -25459
rect 10724 -25493 10758 -25465
rect 10724 -25533 10758 -25531
rect 10724 -25565 10758 -25533
rect 10724 -25635 10758 -25603
rect 10724 -25637 10758 -25635
rect 10724 -25703 10758 -25675
rect 10724 -25709 10758 -25703
rect 10724 -25771 10758 -25747
rect 10724 -25781 10758 -25771
rect 10724 -25839 10758 -25819
rect 10724 -25853 10758 -25839
rect 11742 -25329 11776 -25315
rect 11742 -25349 11776 -25329
rect 11742 -25397 11776 -25387
rect 11742 -25421 11776 -25397
rect 11742 -25465 11776 -25459
rect 11742 -25493 11776 -25465
rect 11742 -25533 11776 -25531
rect 11742 -25565 11776 -25533
rect 11742 -25635 11776 -25603
rect 11742 -25637 11776 -25635
rect 11742 -25703 11776 -25675
rect 11742 -25709 11776 -25703
rect 11742 -25771 11776 -25747
rect 11742 -25781 11776 -25771
rect 11742 -25839 11776 -25819
rect 11742 -25853 11776 -25839
rect 12760 -25329 12794 -25315
rect 12760 -25349 12794 -25329
rect 12760 -25397 12794 -25387
rect 12760 -25421 12794 -25397
rect 12760 -25465 12794 -25459
rect 12760 -25493 12794 -25465
rect 12760 -25533 12794 -25531
rect 12760 -25565 12794 -25533
rect 12760 -25635 12794 -25603
rect 12760 -25637 12794 -25635
rect 12760 -25703 12794 -25675
rect 12760 -25709 12794 -25703
rect 12760 -25771 12794 -25747
rect 12760 -25781 12794 -25771
rect 12760 -25839 12794 -25819
rect 13778 -25329 13812 -25315
rect 13778 -25349 13812 -25329
rect 13778 -25397 13812 -25387
rect 13778 -25421 13812 -25397
rect 13778 -25465 13812 -25459
rect 13778 -25493 13812 -25465
rect 13778 -25533 13812 -25531
rect 13778 -25565 13812 -25533
rect 13778 -25635 13812 -25603
rect 13778 -25637 13812 -25635
rect 13778 -25703 13812 -25675
rect 13778 -25709 13812 -25703
rect 13778 -25771 13812 -25747
rect 13778 -25781 13812 -25771
rect 12760 -25853 12794 -25839
rect 13778 -25839 13812 -25819
rect 14796 -25329 14830 -25315
rect 14796 -25349 14830 -25329
rect 14796 -25397 14830 -25387
rect 14796 -25421 14830 -25397
rect 14796 -25465 14830 -25459
rect 14796 -25493 14830 -25465
rect 14796 -25533 14830 -25531
rect 14796 -25565 14830 -25533
rect 14796 -25635 14830 -25603
rect 14796 -25637 14830 -25635
rect 14796 -25703 14830 -25675
rect 14796 -25709 14830 -25703
rect 14796 -25771 14830 -25747
rect 14796 -25781 14830 -25771
rect 13778 -25853 13812 -25839
rect 14796 -25839 14830 -25819
rect 14796 -25853 14830 -25839
rect 15814 -25329 15848 -25315
rect 15814 -25349 15848 -25329
rect 15814 -25397 15848 -25387
rect 15814 -25421 15848 -25397
rect 15814 -25465 15848 -25459
rect 15814 -25493 15848 -25465
rect 15814 -25533 15848 -25531
rect 15814 -25565 15848 -25533
rect 15814 -25635 15848 -25603
rect 15814 -25637 15848 -25635
rect 15814 -25703 15848 -25675
rect 15814 -25709 15848 -25703
rect 15814 -25771 15848 -25747
rect 15814 -25781 15848 -25771
rect 15814 -25839 15848 -25819
rect 15814 -25853 15848 -25839
rect 16832 -25329 16866 -25315
rect 16832 -25349 16866 -25329
rect 16832 -25397 16866 -25387
rect 16832 -25421 16866 -25397
rect 16832 -25465 16866 -25459
rect 16832 -25493 16866 -25465
rect 16832 -25533 16866 -25531
rect 16832 -25565 16866 -25533
rect 16832 -25635 16866 -25603
rect 16832 -25637 16866 -25635
rect 16832 -25703 16866 -25675
rect 16832 -25709 16866 -25703
rect 16832 -25771 16866 -25747
rect 16832 -25781 16866 -25771
rect 16832 -25839 16866 -25819
rect 17850 -25329 17884 -25315
rect 17850 -25349 17884 -25329
rect 17850 -25397 17884 -25387
rect 17850 -25421 17884 -25397
rect 17850 -25465 17884 -25459
rect 17850 -25493 17884 -25465
rect 17850 -25533 17884 -25531
rect 17850 -25565 17884 -25533
rect 17850 -25635 17884 -25603
rect 17850 -25637 17884 -25635
rect 17850 -25703 17884 -25675
rect 17850 -25709 17884 -25703
rect 17850 -25771 17884 -25747
rect 17850 -25781 17884 -25771
rect 16832 -25853 16866 -25839
rect 17850 -25839 17884 -25819
rect 18868 -25329 18902 -25315
rect 18868 -25349 18902 -25329
rect 18868 -25397 18902 -25387
rect 18868 -25421 18902 -25397
rect 18868 -25465 18902 -25459
rect 18868 -25493 18902 -25465
rect 18868 -25533 18902 -25531
rect 18868 -25565 18902 -25533
rect 18868 -25635 18902 -25603
rect 18868 -25637 18902 -25635
rect 18868 -25703 18902 -25675
rect 18868 -25709 18902 -25703
rect 18868 -25771 18902 -25747
rect 18868 -25781 18902 -25771
rect 17850 -25853 17884 -25839
rect 18868 -25839 18902 -25819
rect 18868 -25853 18902 -25839
rect 19886 -25329 19920 -25315
rect 19886 -25349 19920 -25329
rect 19886 -25397 19920 -25387
rect 19886 -25421 19920 -25397
rect 19886 -25465 19920 -25459
rect 19886 -25493 19920 -25465
rect 19886 -25533 19920 -25531
rect 19886 -25565 19920 -25533
rect 19886 -25635 19920 -25603
rect 19886 -25637 19920 -25635
rect 19886 -25703 19920 -25675
rect 19886 -25709 19920 -25703
rect 19886 -25771 19920 -25747
rect 19886 -25781 19920 -25771
rect 19886 -25839 19920 -25819
rect 19886 -25853 19920 -25839
rect 20904 -25329 20938 -25315
rect 20904 -25349 20938 -25329
rect 20904 -25397 20938 -25387
rect 20904 -25421 20938 -25397
rect 20904 -25465 20938 -25459
rect 20904 -25493 20938 -25465
rect 20904 -25533 20938 -25531
rect 20904 -25565 20938 -25533
rect 20904 -25635 20938 -25603
rect 20904 -25637 20938 -25635
rect 20904 -25703 20938 -25675
rect 20904 -25709 20938 -25703
rect 20904 -25771 20938 -25747
rect 20904 -25781 20938 -25771
rect 20904 -25839 20938 -25819
rect 21922 -25329 21956 -25315
rect 21922 -25349 21956 -25329
rect 21922 -25397 21956 -25387
rect 21922 -25421 21956 -25397
rect 21922 -25465 21956 -25459
rect 21922 -25493 21956 -25465
rect 21922 -25533 21956 -25531
rect 21922 -25565 21956 -25533
rect 21922 -25635 21956 -25603
rect 21922 -25637 21956 -25635
rect 21922 -25703 21956 -25675
rect 21922 -25709 21956 -25703
rect 21922 -25771 21956 -25747
rect 21922 -25781 21956 -25771
rect 20904 -25853 20938 -25839
rect 21922 -25839 21956 -25819
rect 22940 -25329 22974 -25315
rect 22940 -25349 22974 -25329
rect 22940 -25397 22974 -25387
rect 22940 -25421 22974 -25397
rect 22940 -25465 22974 -25459
rect 22940 -25493 22974 -25465
rect 22940 -25533 22974 -25531
rect 22940 -25565 22974 -25533
rect 22940 -25635 22974 -25603
rect 22940 -25637 22974 -25635
rect 22940 -25703 22974 -25675
rect 22940 -25709 22974 -25703
rect 22940 -25771 22974 -25747
rect 22940 -25781 22974 -25771
rect 21922 -25853 21956 -25839
rect 22940 -25839 22974 -25819
rect 22940 -25853 22974 -25839
rect 24855 -25269 24889 -25267
rect 24855 -25301 24889 -25269
rect 24855 -25371 24889 -25339
rect 24855 -25373 24889 -25371
rect 24855 -25439 24889 -25411
rect 24855 -25445 24889 -25439
rect 24855 -25507 24889 -25483
rect 24855 -25517 24889 -25507
rect 24855 -25575 24889 -25555
rect 24855 -25589 24889 -25575
rect 24855 -25643 24889 -25627
rect 24855 -25661 24889 -25643
rect 24855 -25711 24889 -25699
rect 24855 -25733 24889 -25711
rect 24855 -25779 24889 -25771
rect 24855 -25805 24889 -25779
rect 24855 -25847 24889 -25843
rect 24855 -25877 24889 -25847
rect -12289 -25949 -12255 -25915
rect 2909 -25956 2919 -25922
rect 2919 -25956 2943 -25922
rect 2981 -25956 2987 -25922
rect 2987 -25956 3015 -25922
rect 3053 -25956 3055 -25922
rect 3055 -25956 3087 -25922
rect 3125 -25956 3157 -25922
rect 3157 -25956 3159 -25922
rect 3197 -25956 3225 -25922
rect 3225 -25956 3231 -25922
rect 3269 -25956 3293 -25922
rect 3293 -25956 3303 -25922
rect 3927 -25956 3937 -25922
rect 3937 -25956 3961 -25922
rect 3999 -25956 4005 -25922
rect 4005 -25956 4033 -25922
rect 4071 -25956 4073 -25922
rect 4073 -25956 4105 -25922
rect 4143 -25956 4175 -25922
rect 4175 -25956 4177 -25922
rect 4215 -25956 4243 -25922
rect 4243 -25956 4249 -25922
rect 4287 -25956 4311 -25922
rect 4311 -25956 4321 -25922
rect 4945 -25956 4955 -25922
rect 4955 -25956 4979 -25922
rect 5017 -25956 5023 -25922
rect 5023 -25956 5051 -25922
rect 5089 -25956 5091 -25922
rect 5091 -25956 5123 -25922
rect 5161 -25956 5193 -25922
rect 5193 -25956 5195 -25922
rect 5233 -25956 5261 -25922
rect 5261 -25956 5267 -25922
rect 5305 -25956 5329 -25922
rect 5329 -25956 5339 -25922
rect 5963 -25956 5973 -25922
rect 5973 -25956 5997 -25922
rect 6035 -25956 6041 -25922
rect 6041 -25956 6069 -25922
rect 6107 -25956 6109 -25922
rect 6109 -25956 6141 -25922
rect 6179 -25956 6211 -25922
rect 6211 -25956 6213 -25922
rect 6251 -25956 6279 -25922
rect 6279 -25956 6285 -25922
rect 6323 -25956 6347 -25922
rect 6347 -25956 6357 -25922
rect 6981 -25956 6991 -25922
rect 6991 -25956 7015 -25922
rect 7053 -25956 7059 -25922
rect 7059 -25956 7087 -25922
rect 7125 -25956 7127 -25922
rect 7127 -25956 7159 -25922
rect 7197 -25956 7229 -25922
rect 7229 -25956 7231 -25922
rect 7269 -25956 7297 -25922
rect 7297 -25956 7303 -25922
rect 7341 -25956 7365 -25922
rect 7365 -25956 7375 -25922
rect 7999 -25956 8009 -25922
rect 8009 -25956 8033 -25922
rect 8071 -25956 8077 -25922
rect 8077 -25956 8105 -25922
rect 8143 -25956 8145 -25922
rect 8145 -25956 8177 -25922
rect 8215 -25956 8247 -25922
rect 8247 -25956 8249 -25922
rect 8287 -25956 8315 -25922
rect 8315 -25956 8321 -25922
rect 8359 -25956 8383 -25922
rect 8383 -25956 8393 -25922
rect 9017 -25956 9027 -25922
rect 9027 -25956 9051 -25922
rect 9089 -25956 9095 -25922
rect 9095 -25956 9123 -25922
rect 9161 -25956 9163 -25922
rect 9163 -25956 9195 -25922
rect 9233 -25956 9265 -25922
rect 9265 -25956 9267 -25922
rect 9305 -25956 9333 -25922
rect 9333 -25956 9339 -25922
rect 9377 -25956 9401 -25922
rect 9401 -25956 9411 -25922
rect 10035 -25956 10045 -25922
rect 10045 -25956 10069 -25922
rect 10107 -25956 10113 -25922
rect 10113 -25956 10141 -25922
rect 10179 -25956 10181 -25922
rect 10181 -25956 10213 -25922
rect 10251 -25956 10283 -25922
rect 10283 -25956 10285 -25922
rect 10323 -25956 10351 -25922
rect 10351 -25956 10357 -25922
rect 10395 -25956 10419 -25922
rect 10419 -25956 10429 -25922
rect 11053 -25956 11063 -25922
rect 11063 -25956 11087 -25922
rect 11125 -25956 11131 -25922
rect 11131 -25956 11159 -25922
rect 11197 -25956 11199 -25922
rect 11199 -25956 11231 -25922
rect 11269 -25956 11301 -25922
rect 11301 -25956 11303 -25922
rect 11341 -25956 11369 -25922
rect 11369 -25956 11375 -25922
rect 11413 -25956 11437 -25922
rect 11437 -25956 11447 -25922
rect 12071 -25956 12081 -25922
rect 12081 -25956 12105 -25922
rect 12143 -25956 12149 -25922
rect 12149 -25956 12177 -25922
rect 12215 -25956 12217 -25922
rect 12217 -25956 12249 -25922
rect 12287 -25956 12319 -25922
rect 12319 -25956 12321 -25922
rect 12359 -25956 12387 -25922
rect 12387 -25956 12393 -25922
rect 12431 -25956 12455 -25922
rect 12455 -25956 12465 -25922
rect 13089 -25956 13099 -25922
rect 13099 -25956 13123 -25922
rect 13161 -25956 13167 -25922
rect 13167 -25956 13195 -25922
rect 13233 -25956 13235 -25922
rect 13235 -25956 13267 -25922
rect 13305 -25956 13337 -25922
rect 13337 -25956 13339 -25922
rect 13377 -25956 13405 -25922
rect 13405 -25956 13411 -25922
rect 13449 -25956 13473 -25922
rect 13473 -25956 13483 -25922
rect 14107 -25956 14117 -25922
rect 14117 -25956 14141 -25922
rect 14179 -25956 14185 -25922
rect 14185 -25956 14213 -25922
rect 14251 -25956 14253 -25922
rect 14253 -25956 14285 -25922
rect 14323 -25956 14355 -25922
rect 14355 -25956 14357 -25922
rect 14395 -25956 14423 -25922
rect 14423 -25956 14429 -25922
rect 14467 -25956 14491 -25922
rect 14491 -25956 14501 -25922
rect 15125 -25956 15135 -25922
rect 15135 -25956 15159 -25922
rect 15197 -25956 15203 -25922
rect 15203 -25956 15231 -25922
rect 15269 -25956 15271 -25922
rect 15271 -25956 15303 -25922
rect 15341 -25956 15373 -25922
rect 15373 -25956 15375 -25922
rect 15413 -25956 15441 -25922
rect 15441 -25956 15447 -25922
rect 15485 -25956 15509 -25922
rect 15509 -25956 15519 -25922
rect 16143 -25956 16153 -25922
rect 16153 -25956 16177 -25922
rect 16215 -25956 16221 -25922
rect 16221 -25956 16249 -25922
rect 16287 -25956 16289 -25922
rect 16289 -25956 16321 -25922
rect 16359 -25956 16391 -25922
rect 16391 -25956 16393 -25922
rect 16431 -25956 16459 -25922
rect 16459 -25956 16465 -25922
rect 16503 -25956 16527 -25922
rect 16527 -25956 16537 -25922
rect 17161 -25956 17171 -25922
rect 17171 -25956 17195 -25922
rect 17233 -25956 17239 -25922
rect 17239 -25956 17267 -25922
rect 17305 -25956 17307 -25922
rect 17307 -25956 17339 -25922
rect 17377 -25956 17409 -25922
rect 17409 -25956 17411 -25922
rect 17449 -25956 17477 -25922
rect 17477 -25956 17483 -25922
rect 17521 -25956 17545 -25922
rect 17545 -25956 17555 -25922
rect 18179 -25956 18189 -25922
rect 18189 -25956 18213 -25922
rect 18251 -25956 18257 -25922
rect 18257 -25956 18285 -25922
rect 18323 -25956 18325 -25922
rect 18325 -25956 18357 -25922
rect 18395 -25956 18427 -25922
rect 18427 -25956 18429 -25922
rect 18467 -25956 18495 -25922
rect 18495 -25956 18501 -25922
rect 18539 -25956 18563 -25922
rect 18563 -25956 18573 -25922
rect 19197 -25956 19207 -25922
rect 19207 -25956 19231 -25922
rect 19269 -25956 19275 -25922
rect 19275 -25956 19303 -25922
rect 19341 -25956 19343 -25922
rect 19343 -25956 19375 -25922
rect 19413 -25956 19445 -25922
rect 19445 -25956 19447 -25922
rect 19485 -25956 19513 -25922
rect 19513 -25956 19519 -25922
rect 19557 -25956 19581 -25922
rect 19581 -25956 19591 -25922
rect 20215 -25956 20225 -25922
rect 20225 -25956 20249 -25922
rect 20287 -25956 20293 -25922
rect 20293 -25956 20321 -25922
rect 20359 -25956 20361 -25922
rect 20361 -25956 20393 -25922
rect 20431 -25956 20463 -25922
rect 20463 -25956 20465 -25922
rect 20503 -25956 20531 -25922
rect 20531 -25956 20537 -25922
rect 20575 -25956 20599 -25922
rect 20599 -25956 20609 -25922
rect 21233 -25956 21243 -25922
rect 21243 -25956 21267 -25922
rect 21305 -25956 21311 -25922
rect 21311 -25956 21339 -25922
rect 21377 -25956 21379 -25922
rect 21379 -25956 21411 -25922
rect 21449 -25956 21481 -25922
rect 21481 -25956 21483 -25922
rect 21521 -25956 21549 -25922
rect 21549 -25956 21555 -25922
rect 21593 -25956 21617 -25922
rect 21617 -25956 21627 -25922
rect 22251 -25956 22261 -25922
rect 22261 -25956 22285 -25922
rect 22323 -25956 22329 -25922
rect 22329 -25956 22357 -25922
rect 22395 -25956 22397 -25922
rect 22397 -25956 22429 -25922
rect 22467 -25956 22499 -25922
rect 22499 -25956 22501 -25922
rect 22539 -25956 22567 -25922
rect 22567 -25956 22573 -25922
rect 22611 -25956 22635 -25922
rect 22635 -25956 22645 -25922
rect 24855 -25949 24889 -25915
rect -12289 -26017 -12255 -25987
rect -12289 -26021 -12255 -26017
rect -12289 -26085 -12255 -26059
rect -12289 -26093 -12255 -26085
rect -12289 -26153 -12255 -26131
rect -12289 -26165 -12255 -26153
rect -12289 -26221 -12255 -26203
rect -12289 -26237 -12255 -26221
rect -12289 -26289 -12255 -26275
rect -12289 -26309 -12255 -26289
rect 24855 -26017 24889 -25987
rect 24855 -26021 24889 -26017
rect 24855 -26085 24889 -26059
rect 24855 -26093 24889 -26085
rect 24855 -26153 24889 -26131
rect 24855 -26165 24889 -26153
rect 24855 -26221 24889 -26203
rect 24855 -26237 24889 -26221
rect 24855 -26289 24889 -26275
rect 24855 -26309 24889 -26289
rect -12221 -27189 -12187 -27155
rect -12149 -27189 -12145 -27155
rect -12145 -27189 -12115 -27155
rect -12077 -27189 -12043 -27155
rect -12005 -27189 -11975 -27155
rect -11975 -27189 -11971 -27155
rect -11933 -27189 -11907 -27155
rect -11907 -27189 -11899 -27155
rect -11861 -27189 -11839 -27155
rect -11839 -27189 -11827 -27155
rect -11789 -27189 -11771 -27155
rect -11771 -27189 -11755 -27155
rect -11717 -27189 -11703 -27155
rect -11703 -27189 -11683 -27155
rect -11645 -27189 -11635 -27155
rect -11635 -27189 -11611 -27155
rect -11573 -27189 -11567 -27155
rect -11567 -27189 -11539 -27155
rect -11501 -27189 -11499 -27155
rect -11499 -27189 -11467 -27155
rect -11429 -27189 -11397 -27155
rect -11397 -27189 -11395 -27155
rect -11357 -27189 -11329 -27155
rect -11329 -27189 -11323 -27155
rect -11285 -27189 -11261 -27155
rect -11261 -27189 -11251 -27155
rect -11213 -27189 -11193 -27155
rect -11193 -27189 -11179 -27155
rect -11141 -27189 -11125 -27155
rect -11125 -27189 -11107 -27155
rect -11069 -27189 -11057 -27155
rect -11057 -27189 -11035 -27155
rect -10997 -27189 -10989 -27155
rect -10989 -27189 -10963 -27155
rect -10925 -27189 -10921 -27155
rect -10921 -27189 -10891 -27155
rect -10853 -27189 -10819 -27155
rect -10781 -27189 -10751 -27155
rect -10751 -27189 -10747 -27155
rect -10709 -27189 -10683 -27155
rect -10683 -27189 -10675 -27155
rect -10637 -27189 -10615 -27155
rect -10615 -27189 -10603 -27155
rect -10565 -27189 -10547 -27155
rect -10547 -27189 -10531 -27155
rect -10493 -27189 -10479 -27155
rect -10479 -27189 -10459 -27155
rect -10421 -27189 -10411 -27155
rect -10411 -27189 -10387 -27155
rect -10349 -27189 -10343 -27155
rect -10343 -27189 -10315 -27155
rect -10277 -27189 -10275 -27155
rect -10275 -27189 -10243 -27155
rect -10205 -27189 -10173 -27155
rect -10173 -27189 -10171 -27155
rect -10133 -27189 -10105 -27155
rect -10105 -27189 -10099 -27155
rect -10061 -27189 -10037 -27155
rect -10037 -27189 -10027 -27155
rect -9989 -27189 -9969 -27155
rect -9969 -27189 -9955 -27155
rect -9917 -27189 -9901 -27155
rect -9901 -27189 -9883 -27155
rect -9845 -27189 -9833 -27155
rect -9833 -27189 -9811 -27155
rect -9773 -27189 -9765 -27155
rect -9765 -27189 -9739 -27155
rect -9701 -27189 -9697 -27155
rect -9697 -27189 -9667 -27155
rect -9629 -27189 -9595 -27155
rect -9557 -27189 -9527 -27155
rect -9527 -27189 -9523 -27155
rect -9485 -27189 -9459 -27155
rect -9459 -27189 -9451 -27155
rect -9413 -27189 -9391 -27155
rect -9391 -27189 -9379 -27155
rect -9341 -27189 -9323 -27155
rect -9323 -27189 -9307 -27155
rect -9269 -27189 -9255 -27155
rect -9255 -27189 -9235 -27155
rect -9197 -27189 -9187 -27155
rect -9187 -27189 -9163 -27155
rect -9125 -27189 -9119 -27155
rect -9119 -27189 -9091 -27155
rect -9053 -27189 -9051 -27155
rect -9051 -27189 -9019 -27155
rect -8981 -27189 -8949 -27155
rect -8949 -27189 -8947 -27155
rect -8909 -27189 -8881 -27155
rect -8881 -27189 -8875 -27155
rect -8837 -27189 -8813 -27155
rect -8813 -27189 -8803 -27155
rect -8765 -27189 -8745 -27155
rect -8745 -27189 -8731 -27155
rect -8693 -27189 -8677 -27155
rect -8677 -27189 -8659 -27155
rect -8621 -27189 -8609 -27155
rect -8609 -27189 -8587 -27155
rect -8549 -27189 -8541 -27155
rect -8541 -27189 -8515 -27155
rect -8477 -27189 -8473 -27155
rect -8473 -27189 -8443 -27155
rect -8405 -27189 -8371 -27155
rect -8333 -27189 -8303 -27155
rect -8303 -27189 -8299 -27155
rect -8261 -27189 -8235 -27155
rect -8235 -27189 -8227 -27155
rect -8189 -27189 -8167 -27155
rect -8167 -27189 -8155 -27155
rect -8117 -27189 -8099 -27155
rect -8099 -27189 -8083 -27155
rect -8045 -27189 -8031 -27155
rect -8031 -27189 -8011 -27155
rect -7973 -27189 -7963 -27155
rect -7963 -27189 -7939 -27155
rect -7901 -27189 -7895 -27155
rect -7895 -27189 -7867 -27155
rect -7829 -27189 -7827 -27155
rect -7827 -27189 -7795 -27155
rect -7757 -27189 -7725 -27155
rect -7725 -27189 -7723 -27155
rect -7685 -27189 -7657 -27155
rect -7657 -27189 -7651 -27155
rect -7613 -27189 -7589 -27155
rect -7589 -27189 -7579 -27155
rect -7541 -27189 -7521 -27155
rect -7521 -27189 -7507 -27155
rect -7469 -27189 -7453 -27155
rect -7453 -27189 -7435 -27155
rect -7397 -27189 -7385 -27155
rect -7385 -27189 -7363 -27155
rect -7325 -27189 -7317 -27155
rect -7317 -27189 -7291 -27155
rect -7253 -27189 -7249 -27155
rect -7249 -27189 -7219 -27155
rect -7181 -27189 -7147 -27155
rect -7109 -27189 -7079 -27155
rect -7079 -27189 -7075 -27155
rect -7037 -27189 -7011 -27155
rect -7011 -27189 -7003 -27155
rect -6965 -27189 -6943 -27155
rect -6943 -27189 -6931 -27155
rect -6893 -27189 -6875 -27155
rect -6875 -27189 -6859 -27155
rect -6821 -27189 -6807 -27155
rect -6807 -27189 -6787 -27155
rect -6749 -27189 -6739 -27155
rect -6739 -27189 -6715 -27155
rect -6677 -27189 -6671 -27155
rect -6671 -27189 -6643 -27155
rect -6605 -27189 -6603 -27155
rect -6603 -27189 -6571 -27155
rect -6533 -27189 -6501 -27155
rect -6501 -27189 -6499 -27155
rect -6461 -27189 -6433 -27155
rect -6433 -27189 -6427 -27155
rect -6389 -27189 -6365 -27155
rect -6365 -27189 -6355 -27155
rect -6317 -27189 -6297 -27155
rect -6297 -27189 -6283 -27155
rect -6245 -27189 -6229 -27155
rect -6229 -27189 -6211 -27155
rect -6173 -27189 -6161 -27155
rect -6161 -27189 -6139 -27155
rect -6101 -27189 -6093 -27155
rect -6093 -27189 -6067 -27155
rect -6029 -27189 -6025 -27155
rect -6025 -27189 -5995 -27155
rect -5957 -27189 -5923 -27155
rect -5885 -27189 -5855 -27155
rect -5855 -27189 -5851 -27155
rect -5813 -27189 -5787 -27155
rect -5787 -27189 -5779 -27155
rect -5741 -27189 -5719 -27155
rect -5719 -27189 -5707 -27155
rect -5669 -27189 -5651 -27155
rect -5651 -27189 -5635 -27155
rect -5597 -27189 -5583 -27155
rect -5583 -27189 -5563 -27155
rect -5525 -27189 -5515 -27155
rect -5515 -27189 -5491 -27155
rect -5453 -27189 -5447 -27155
rect -5447 -27189 -5419 -27155
rect -5381 -27189 -5379 -27155
rect -5379 -27189 -5347 -27155
rect -5309 -27189 -5277 -27155
rect -5277 -27189 -5275 -27155
rect -5237 -27189 -5209 -27155
rect -5209 -27189 -5203 -27155
rect -5165 -27189 -5141 -27155
rect -5141 -27189 -5131 -27155
rect -5093 -27189 -5073 -27155
rect -5073 -27189 -5059 -27155
rect -5021 -27189 -5005 -27155
rect -5005 -27189 -4987 -27155
rect -4949 -27189 -4937 -27155
rect -4937 -27189 -4915 -27155
rect -4877 -27189 -4869 -27155
rect -4869 -27189 -4843 -27155
rect -4805 -27189 -4801 -27155
rect -4801 -27189 -4771 -27155
rect -4733 -27189 -4699 -27155
rect -4661 -27189 -4631 -27155
rect -4631 -27189 -4627 -27155
rect -4589 -27189 -4563 -27155
rect -4563 -27189 -4555 -27155
rect -4517 -27189 -4495 -27155
rect -4495 -27189 -4483 -27155
rect -4445 -27189 -4427 -27155
rect -4427 -27189 -4411 -27155
rect -4373 -27189 -4359 -27155
rect -4359 -27189 -4339 -27155
rect -4301 -27189 -4291 -27155
rect -4291 -27189 -4267 -27155
rect -4229 -27189 -4223 -27155
rect -4223 -27189 -4195 -27155
rect -4157 -27189 -4155 -27155
rect -4155 -27189 -4123 -27155
rect -4085 -27189 -4053 -27155
rect -4053 -27189 -4051 -27155
rect -4013 -27189 -3985 -27155
rect -3985 -27189 -3979 -27155
rect -3941 -27189 -3917 -27155
rect -3917 -27189 -3907 -27155
rect -3869 -27189 -3849 -27155
rect -3849 -27189 -3835 -27155
rect -3797 -27189 -3781 -27155
rect -3781 -27189 -3763 -27155
rect -3725 -27189 -3713 -27155
rect -3713 -27189 -3691 -27155
rect -3653 -27189 -3645 -27155
rect -3645 -27189 -3619 -27155
rect -3581 -27189 -3577 -27155
rect -3577 -27189 -3547 -27155
rect -3509 -27189 -3475 -27155
rect -3437 -27189 -3407 -27155
rect -3407 -27189 -3403 -27155
rect -3365 -27189 -3339 -27155
rect -3339 -27189 -3331 -27155
rect -3293 -27189 -3271 -27155
rect -3271 -27189 -3259 -27155
rect -3221 -27189 -3203 -27155
rect -3203 -27189 -3187 -27155
rect -3149 -27189 -3135 -27155
rect -3135 -27189 -3115 -27155
rect -3077 -27189 -3067 -27155
rect -3067 -27189 -3043 -27155
rect -3005 -27189 -2999 -27155
rect -2999 -27189 -2971 -27155
rect -2933 -27189 -2931 -27155
rect -2931 -27189 -2899 -27155
rect -2861 -27189 -2829 -27155
rect -2829 -27189 -2827 -27155
rect -2789 -27189 -2761 -27155
rect -2761 -27189 -2755 -27155
rect -2717 -27189 -2693 -27155
rect -2693 -27189 -2683 -27155
rect -2645 -27189 -2625 -27155
rect -2625 -27189 -2611 -27155
rect -2573 -27189 -2557 -27155
rect -2557 -27189 -2539 -27155
rect -2501 -27189 -2489 -27155
rect -2489 -27189 -2467 -27155
rect -2429 -27189 -2421 -27155
rect -2421 -27189 -2395 -27155
rect -2357 -27189 -2353 -27155
rect -2353 -27189 -2323 -27155
rect -2285 -27189 -2251 -27155
rect -2213 -27189 -2183 -27155
rect -2183 -27189 -2179 -27155
rect -2141 -27189 -2115 -27155
rect -2115 -27189 -2107 -27155
rect -2069 -27189 -2047 -27155
rect -2047 -27189 -2035 -27155
rect -1997 -27189 -1979 -27155
rect -1979 -27189 -1963 -27155
rect -1925 -27189 -1911 -27155
rect -1911 -27189 -1891 -27155
rect -1853 -27189 -1843 -27155
rect -1843 -27189 -1819 -27155
rect -1781 -27189 -1775 -27155
rect -1775 -27189 -1747 -27155
rect -1709 -27189 -1707 -27155
rect -1707 -27189 -1675 -27155
rect -1637 -27189 -1605 -27155
rect -1605 -27189 -1603 -27155
rect -1565 -27189 -1537 -27155
rect -1537 -27189 -1531 -27155
rect -1493 -27189 -1469 -27155
rect -1469 -27189 -1459 -27155
rect -1421 -27189 -1401 -27155
rect -1401 -27189 -1387 -27155
rect -1349 -27189 -1333 -27155
rect -1333 -27189 -1315 -27155
rect -1277 -27189 -1265 -27155
rect -1265 -27189 -1243 -27155
rect -1205 -27189 -1197 -27155
rect -1197 -27189 -1171 -27155
rect -1133 -27189 -1129 -27155
rect -1129 -27189 -1099 -27155
rect -1061 -27189 -1027 -27155
rect -989 -27189 -959 -27155
rect -959 -27189 -955 -27155
rect -917 -27189 -891 -27155
rect -891 -27189 -883 -27155
rect -845 -27189 -823 -27155
rect -823 -27189 -811 -27155
rect -773 -27189 -755 -27155
rect -755 -27189 -739 -27155
rect -701 -27189 -687 -27155
rect -687 -27189 -667 -27155
rect -629 -27189 -619 -27155
rect -619 -27189 -595 -27155
rect -557 -27189 -551 -27155
rect -551 -27189 -523 -27155
rect -485 -27189 -483 -27155
rect -483 -27189 -451 -27155
rect -413 -27189 -381 -27155
rect -381 -27189 -379 -27155
rect -341 -27189 -313 -27155
rect -313 -27189 -307 -27155
rect -269 -27189 -245 -27155
rect -245 -27189 -235 -27155
rect -197 -27189 -177 -27155
rect -177 -27189 -163 -27155
rect -125 -27189 -109 -27155
rect -109 -27189 -91 -27155
rect -53 -27189 -41 -27155
rect -41 -27189 -19 -27155
rect 19 -27189 27 -27155
rect 27 -27189 53 -27155
rect 91 -27189 95 -27155
rect 95 -27189 125 -27155
rect 163 -27189 197 -27155
rect 235 -27189 265 -27155
rect 265 -27189 269 -27155
rect 307 -27189 333 -27155
rect 333 -27189 341 -27155
rect 379 -27189 401 -27155
rect 401 -27189 413 -27155
rect 451 -27189 469 -27155
rect 469 -27189 485 -27155
rect 523 -27189 537 -27155
rect 537 -27189 557 -27155
rect 595 -27189 605 -27155
rect 605 -27189 629 -27155
rect 667 -27189 673 -27155
rect 673 -27189 701 -27155
rect 739 -27189 741 -27155
rect 741 -27189 773 -27155
rect 811 -27189 843 -27155
rect 843 -27189 845 -27155
rect 883 -27189 911 -27155
rect 911 -27189 917 -27155
rect 955 -27189 979 -27155
rect 979 -27189 989 -27155
rect 1027 -27189 1047 -27155
rect 1047 -27189 1061 -27155
rect 1099 -27189 1115 -27155
rect 1115 -27189 1133 -27155
rect 1171 -27189 1183 -27155
rect 1183 -27189 1205 -27155
rect 1243 -27189 1251 -27155
rect 1251 -27189 1277 -27155
rect 1315 -27189 1319 -27155
rect 1319 -27189 1349 -27155
rect 1387 -27189 1421 -27155
rect 1459 -27189 1489 -27155
rect 1489 -27189 1493 -27155
rect 1531 -27189 1557 -27155
rect 1557 -27189 1565 -27155
rect 1603 -27189 1625 -27155
rect 1625 -27189 1637 -27155
rect 1675 -27189 1693 -27155
rect 1693 -27189 1709 -27155
rect 1747 -27189 1761 -27155
rect 1761 -27189 1781 -27155
rect 1819 -27189 1829 -27155
rect 1829 -27189 1853 -27155
rect 1891 -27189 1897 -27155
rect 1897 -27189 1925 -27155
rect 1963 -27189 1965 -27155
rect 1965 -27189 1997 -27155
rect 2035 -27189 2067 -27155
rect 2067 -27189 2069 -27155
rect 2107 -27189 2135 -27155
rect 2135 -27189 2141 -27155
rect 2179 -27189 2203 -27155
rect 2203 -27189 2213 -27155
rect 2251 -27189 2271 -27155
rect 2271 -27189 2285 -27155
rect 2323 -27189 2339 -27155
rect 2339 -27189 2357 -27155
rect 2395 -27189 2407 -27155
rect 2407 -27189 2429 -27155
rect 2467 -27189 2475 -27155
rect 2475 -27189 2501 -27155
rect 2539 -27189 2543 -27155
rect 2543 -27189 2573 -27155
rect 2611 -27189 2645 -27155
rect 2683 -27189 2713 -27155
rect 2713 -27189 2717 -27155
rect 2755 -27189 2781 -27155
rect 2781 -27189 2789 -27155
rect 2827 -27189 2849 -27155
rect 2849 -27189 2861 -27155
rect 2899 -27189 2917 -27155
rect 2917 -27189 2933 -27155
rect 2971 -27189 2985 -27155
rect 2985 -27189 3005 -27155
rect 3043 -27189 3053 -27155
rect 3053 -27189 3077 -27155
rect 3115 -27189 3121 -27155
rect 3121 -27189 3149 -27155
rect 3187 -27189 3189 -27155
rect 3189 -27189 3221 -27155
rect 3259 -27189 3291 -27155
rect 3291 -27189 3293 -27155
rect 3331 -27189 3359 -27155
rect 3359 -27189 3365 -27155
rect 3403 -27189 3427 -27155
rect 3427 -27189 3437 -27155
rect 3475 -27189 3495 -27155
rect 3495 -27189 3509 -27155
rect 3547 -27189 3563 -27155
rect 3563 -27189 3581 -27155
rect 3619 -27189 3631 -27155
rect 3631 -27189 3653 -27155
rect 3691 -27189 3699 -27155
rect 3699 -27189 3725 -27155
rect 3763 -27189 3767 -27155
rect 3767 -27189 3797 -27155
rect 3835 -27189 3869 -27155
rect 3907 -27189 3937 -27155
rect 3937 -27189 3941 -27155
rect 3979 -27189 4005 -27155
rect 4005 -27189 4013 -27155
rect 4051 -27189 4073 -27155
rect 4073 -27189 4085 -27155
rect 4123 -27189 4141 -27155
rect 4141 -27189 4157 -27155
rect 4195 -27189 4209 -27155
rect 4209 -27189 4229 -27155
rect 4267 -27189 4277 -27155
rect 4277 -27189 4301 -27155
rect 4339 -27189 4345 -27155
rect 4345 -27189 4373 -27155
rect 4411 -27189 4413 -27155
rect 4413 -27189 4445 -27155
rect 4483 -27189 4515 -27155
rect 4515 -27189 4517 -27155
rect 4555 -27189 4583 -27155
rect 4583 -27189 4589 -27155
rect 4627 -27189 4651 -27155
rect 4651 -27189 4661 -27155
rect 4699 -27189 4719 -27155
rect 4719 -27189 4733 -27155
rect 4771 -27189 4787 -27155
rect 4787 -27189 4805 -27155
rect 4843 -27189 4855 -27155
rect 4855 -27189 4877 -27155
rect 4915 -27189 4923 -27155
rect 4923 -27189 4949 -27155
rect 4987 -27189 4991 -27155
rect 4991 -27189 5021 -27155
rect 5059 -27189 5093 -27155
rect 5131 -27189 5161 -27155
rect 5161 -27189 5165 -27155
rect 5203 -27189 5229 -27155
rect 5229 -27189 5237 -27155
rect 5275 -27189 5297 -27155
rect 5297 -27189 5309 -27155
rect 5347 -27189 5365 -27155
rect 5365 -27189 5381 -27155
rect 5419 -27189 5433 -27155
rect 5433 -27189 5453 -27155
rect 5491 -27189 5501 -27155
rect 5501 -27189 5525 -27155
rect 5563 -27189 5569 -27155
rect 5569 -27189 5597 -27155
rect 5635 -27189 5637 -27155
rect 5637 -27189 5669 -27155
rect 5707 -27189 5739 -27155
rect 5739 -27189 5741 -27155
rect 5779 -27189 5807 -27155
rect 5807 -27189 5813 -27155
rect 5851 -27189 5875 -27155
rect 5875 -27189 5885 -27155
rect 5923 -27189 5943 -27155
rect 5943 -27189 5957 -27155
rect 5995 -27189 6011 -27155
rect 6011 -27189 6029 -27155
rect 6067 -27189 6079 -27155
rect 6079 -27189 6101 -27155
rect 6139 -27189 6147 -27155
rect 6147 -27189 6173 -27155
rect 6211 -27189 6215 -27155
rect 6215 -27189 6245 -27155
rect 6283 -27189 6317 -27155
rect 6355 -27189 6385 -27155
rect 6385 -27189 6389 -27155
rect 6427 -27189 6453 -27155
rect 6453 -27189 6461 -27155
rect 6499 -27189 6521 -27155
rect 6521 -27189 6533 -27155
rect 6571 -27189 6589 -27155
rect 6589 -27189 6605 -27155
rect 6643 -27189 6657 -27155
rect 6657 -27189 6677 -27155
rect 6715 -27189 6725 -27155
rect 6725 -27189 6749 -27155
rect 6787 -27189 6793 -27155
rect 6793 -27189 6821 -27155
rect 6859 -27189 6861 -27155
rect 6861 -27189 6893 -27155
rect 6931 -27189 6963 -27155
rect 6963 -27189 6965 -27155
rect 7003 -27189 7031 -27155
rect 7031 -27189 7037 -27155
rect 7075 -27189 7099 -27155
rect 7099 -27189 7109 -27155
rect 7147 -27189 7167 -27155
rect 7167 -27189 7181 -27155
rect 7219 -27189 7235 -27155
rect 7235 -27189 7253 -27155
rect 7291 -27189 7303 -27155
rect 7303 -27189 7325 -27155
rect 7363 -27189 7371 -27155
rect 7371 -27189 7397 -27155
rect 7435 -27189 7439 -27155
rect 7439 -27189 7469 -27155
rect 7507 -27189 7541 -27155
rect 7579 -27189 7609 -27155
rect 7609 -27189 7613 -27155
rect 7651 -27189 7677 -27155
rect 7677 -27189 7685 -27155
rect 7723 -27189 7745 -27155
rect 7745 -27189 7757 -27155
rect 7795 -27189 7813 -27155
rect 7813 -27189 7829 -27155
rect 7867 -27189 7881 -27155
rect 7881 -27189 7901 -27155
rect 7939 -27189 7949 -27155
rect 7949 -27189 7973 -27155
rect 8011 -27189 8017 -27155
rect 8017 -27189 8045 -27155
rect 8083 -27189 8085 -27155
rect 8085 -27189 8117 -27155
rect 8155 -27189 8187 -27155
rect 8187 -27189 8189 -27155
rect 8227 -27189 8255 -27155
rect 8255 -27189 8261 -27155
rect 8299 -27189 8323 -27155
rect 8323 -27189 8333 -27155
rect 8371 -27189 8391 -27155
rect 8391 -27189 8405 -27155
rect 8443 -27189 8459 -27155
rect 8459 -27189 8477 -27155
rect 8515 -27189 8527 -27155
rect 8527 -27189 8549 -27155
rect 8587 -27189 8595 -27155
rect 8595 -27189 8621 -27155
rect 8659 -27189 8663 -27155
rect 8663 -27189 8693 -27155
rect 8731 -27189 8765 -27155
rect 8803 -27189 8833 -27155
rect 8833 -27189 8837 -27155
rect 8875 -27189 8901 -27155
rect 8901 -27189 8909 -27155
rect 8947 -27189 8969 -27155
rect 8969 -27189 8981 -27155
rect 9019 -27189 9037 -27155
rect 9037 -27189 9053 -27155
rect 9091 -27189 9105 -27155
rect 9105 -27189 9125 -27155
rect 9163 -27189 9173 -27155
rect 9173 -27189 9197 -27155
rect 9235 -27189 9241 -27155
rect 9241 -27189 9269 -27155
rect 9307 -27189 9309 -27155
rect 9309 -27189 9341 -27155
rect 9379 -27189 9411 -27155
rect 9411 -27189 9413 -27155
rect 9451 -27189 9479 -27155
rect 9479 -27189 9485 -27155
rect 9523 -27189 9547 -27155
rect 9547 -27189 9557 -27155
rect 9595 -27189 9615 -27155
rect 9615 -27189 9629 -27155
rect 9667 -27189 9683 -27155
rect 9683 -27189 9701 -27155
rect 9739 -27189 9751 -27155
rect 9751 -27189 9773 -27155
rect 9811 -27189 9819 -27155
rect 9819 -27189 9845 -27155
rect 9883 -27189 9887 -27155
rect 9887 -27189 9917 -27155
rect 9955 -27189 9989 -27155
rect 10027 -27189 10057 -27155
rect 10057 -27189 10061 -27155
rect 10099 -27189 10125 -27155
rect 10125 -27189 10133 -27155
rect 10171 -27189 10193 -27155
rect 10193 -27189 10205 -27155
rect 10243 -27189 10261 -27155
rect 10261 -27189 10277 -27155
rect 10315 -27189 10329 -27155
rect 10329 -27189 10349 -27155
rect 10387 -27189 10397 -27155
rect 10397 -27189 10421 -27155
rect 10459 -27189 10465 -27155
rect 10465 -27189 10493 -27155
rect 10531 -27189 10533 -27155
rect 10533 -27189 10565 -27155
rect 10603 -27189 10635 -27155
rect 10635 -27189 10637 -27155
rect 10675 -27189 10703 -27155
rect 10703 -27189 10709 -27155
rect 10747 -27189 10771 -27155
rect 10771 -27189 10781 -27155
rect 10819 -27189 10839 -27155
rect 10839 -27189 10853 -27155
rect 10891 -27189 10907 -27155
rect 10907 -27189 10925 -27155
rect 10963 -27189 10975 -27155
rect 10975 -27189 10997 -27155
rect 11035 -27189 11043 -27155
rect 11043 -27189 11069 -27155
rect 11107 -27189 11111 -27155
rect 11111 -27189 11141 -27155
rect 11179 -27189 11213 -27155
rect 11251 -27189 11281 -27155
rect 11281 -27189 11285 -27155
rect 11323 -27189 11349 -27155
rect 11349 -27189 11357 -27155
rect 11395 -27189 11417 -27155
rect 11417 -27189 11429 -27155
rect 11467 -27189 11485 -27155
rect 11485 -27189 11501 -27155
rect 11539 -27189 11553 -27155
rect 11553 -27189 11573 -27155
rect 11611 -27189 11621 -27155
rect 11621 -27189 11645 -27155
rect 11683 -27189 11689 -27155
rect 11689 -27189 11717 -27155
rect 11755 -27189 11757 -27155
rect 11757 -27189 11789 -27155
rect 11827 -27189 11859 -27155
rect 11859 -27189 11861 -27155
rect 11899 -27189 11927 -27155
rect 11927 -27189 11933 -27155
rect 11971 -27189 11995 -27155
rect 11995 -27189 12005 -27155
rect 12043 -27189 12063 -27155
rect 12063 -27189 12077 -27155
rect 12115 -27189 12131 -27155
rect 12131 -27189 12149 -27155
rect 12187 -27189 12199 -27155
rect 12199 -27189 12221 -27155
rect 12259 -27189 12267 -27155
rect 12267 -27189 12293 -27155
rect 12331 -27189 12335 -27155
rect 12335 -27189 12365 -27155
rect 12403 -27189 12437 -27155
rect 12475 -27189 12505 -27155
rect 12505 -27189 12509 -27155
rect 12547 -27189 12573 -27155
rect 12573 -27189 12581 -27155
rect 12619 -27189 12641 -27155
rect 12641 -27189 12653 -27155
rect 12691 -27189 12709 -27155
rect 12709 -27189 12725 -27155
rect 12763 -27189 12777 -27155
rect 12777 -27189 12797 -27155
rect 12835 -27189 12845 -27155
rect 12845 -27189 12869 -27155
rect 12907 -27189 12913 -27155
rect 12913 -27189 12941 -27155
rect 12979 -27189 12981 -27155
rect 12981 -27189 13013 -27155
rect 13051 -27189 13083 -27155
rect 13083 -27189 13085 -27155
rect 13123 -27189 13151 -27155
rect 13151 -27189 13157 -27155
rect 13195 -27189 13219 -27155
rect 13219 -27189 13229 -27155
rect 13267 -27189 13287 -27155
rect 13287 -27189 13301 -27155
rect 13339 -27189 13355 -27155
rect 13355 -27189 13373 -27155
rect 13411 -27189 13423 -27155
rect 13423 -27189 13445 -27155
rect 13483 -27189 13491 -27155
rect 13491 -27189 13517 -27155
rect 13555 -27189 13559 -27155
rect 13559 -27189 13589 -27155
rect 13627 -27189 13661 -27155
rect 13699 -27189 13729 -27155
rect 13729 -27189 13733 -27155
rect 13771 -27189 13797 -27155
rect 13797 -27189 13805 -27155
rect 13843 -27189 13865 -27155
rect 13865 -27189 13877 -27155
rect 13915 -27189 13933 -27155
rect 13933 -27189 13949 -27155
rect 13987 -27189 14001 -27155
rect 14001 -27189 14021 -27155
rect 14059 -27189 14069 -27155
rect 14069 -27189 14093 -27155
rect 14131 -27189 14137 -27155
rect 14137 -27189 14165 -27155
rect 14203 -27189 14205 -27155
rect 14205 -27189 14237 -27155
rect 14275 -27189 14307 -27155
rect 14307 -27189 14309 -27155
rect 14347 -27189 14375 -27155
rect 14375 -27189 14381 -27155
rect 14419 -27189 14443 -27155
rect 14443 -27189 14453 -27155
rect 14491 -27189 14511 -27155
rect 14511 -27189 14525 -27155
rect 14563 -27189 14579 -27155
rect 14579 -27189 14597 -27155
rect 14635 -27189 14647 -27155
rect 14647 -27189 14669 -27155
rect 14707 -27189 14715 -27155
rect 14715 -27189 14741 -27155
rect 14779 -27189 14783 -27155
rect 14783 -27189 14813 -27155
rect 14851 -27189 14885 -27155
rect 14923 -27189 14953 -27155
rect 14953 -27189 14957 -27155
rect 14995 -27189 15021 -27155
rect 15021 -27189 15029 -27155
rect 15067 -27189 15089 -27155
rect 15089 -27189 15101 -27155
rect 15139 -27189 15157 -27155
rect 15157 -27189 15173 -27155
rect 15211 -27189 15225 -27155
rect 15225 -27189 15245 -27155
rect 15283 -27189 15293 -27155
rect 15293 -27189 15317 -27155
rect 15355 -27189 15361 -27155
rect 15361 -27189 15389 -27155
rect 15427 -27189 15429 -27155
rect 15429 -27189 15461 -27155
rect 15499 -27189 15531 -27155
rect 15531 -27189 15533 -27155
rect 15571 -27189 15599 -27155
rect 15599 -27189 15605 -27155
rect 15643 -27189 15667 -27155
rect 15667 -27189 15677 -27155
rect 15715 -27189 15735 -27155
rect 15735 -27189 15749 -27155
rect 15787 -27189 15803 -27155
rect 15803 -27189 15821 -27155
rect 15859 -27189 15871 -27155
rect 15871 -27189 15893 -27155
rect 15931 -27189 15939 -27155
rect 15939 -27189 15965 -27155
rect 16003 -27189 16007 -27155
rect 16007 -27189 16037 -27155
rect 16075 -27189 16109 -27155
rect 16147 -27189 16177 -27155
rect 16177 -27189 16181 -27155
rect 16219 -27189 16245 -27155
rect 16245 -27189 16253 -27155
rect 16291 -27189 16313 -27155
rect 16313 -27189 16325 -27155
rect 16363 -27189 16381 -27155
rect 16381 -27189 16397 -27155
rect 16435 -27189 16449 -27155
rect 16449 -27189 16469 -27155
rect 16507 -27189 16517 -27155
rect 16517 -27189 16541 -27155
rect 16579 -27189 16585 -27155
rect 16585 -27189 16613 -27155
rect 16651 -27189 16653 -27155
rect 16653 -27189 16685 -27155
rect 16723 -27189 16755 -27155
rect 16755 -27189 16757 -27155
rect 16795 -27189 16823 -27155
rect 16823 -27189 16829 -27155
rect 16867 -27189 16891 -27155
rect 16891 -27189 16901 -27155
rect 16939 -27189 16959 -27155
rect 16959 -27189 16973 -27155
rect 17011 -27189 17027 -27155
rect 17027 -27189 17045 -27155
rect 17083 -27189 17095 -27155
rect 17095 -27189 17117 -27155
rect 17155 -27189 17163 -27155
rect 17163 -27189 17189 -27155
rect 17227 -27189 17231 -27155
rect 17231 -27189 17261 -27155
rect 17299 -27189 17333 -27155
rect 17371 -27189 17401 -27155
rect 17401 -27189 17405 -27155
rect 17443 -27189 17469 -27155
rect 17469 -27189 17477 -27155
rect 17515 -27189 17537 -27155
rect 17537 -27189 17549 -27155
rect 17587 -27189 17605 -27155
rect 17605 -27189 17621 -27155
rect 17659 -27189 17673 -27155
rect 17673 -27189 17693 -27155
rect 17731 -27189 17741 -27155
rect 17741 -27189 17765 -27155
rect 17803 -27189 17809 -27155
rect 17809 -27189 17837 -27155
rect 17875 -27189 17877 -27155
rect 17877 -27189 17909 -27155
rect 17947 -27189 17979 -27155
rect 17979 -27189 17981 -27155
rect 18019 -27189 18047 -27155
rect 18047 -27189 18053 -27155
rect 18091 -27189 18115 -27155
rect 18115 -27189 18125 -27155
rect 18163 -27189 18183 -27155
rect 18183 -27189 18197 -27155
rect 18235 -27189 18251 -27155
rect 18251 -27189 18269 -27155
rect 18307 -27189 18319 -27155
rect 18319 -27189 18341 -27155
rect 18379 -27189 18387 -27155
rect 18387 -27189 18413 -27155
rect 18451 -27189 18455 -27155
rect 18455 -27189 18485 -27155
rect 18523 -27189 18557 -27155
rect 18595 -27189 18625 -27155
rect 18625 -27189 18629 -27155
rect 18667 -27189 18693 -27155
rect 18693 -27189 18701 -27155
rect 18739 -27189 18761 -27155
rect 18761 -27189 18773 -27155
rect 18811 -27189 18829 -27155
rect 18829 -27189 18845 -27155
rect 18883 -27189 18897 -27155
rect 18897 -27189 18917 -27155
rect 18955 -27189 18965 -27155
rect 18965 -27189 18989 -27155
rect 19027 -27189 19033 -27155
rect 19033 -27189 19061 -27155
rect 19099 -27189 19101 -27155
rect 19101 -27189 19133 -27155
rect 19171 -27189 19203 -27155
rect 19203 -27189 19205 -27155
rect 19243 -27189 19271 -27155
rect 19271 -27189 19277 -27155
rect 19315 -27189 19339 -27155
rect 19339 -27189 19349 -27155
rect 19387 -27189 19407 -27155
rect 19407 -27189 19421 -27155
rect 19459 -27189 19475 -27155
rect 19475 -27189 19493 -27155
rect 19531 -27189 19543 -27155
rect 19543 -27189 19565 -27155
rect 19603 -27189 19611 -27155
rect 19611 -27189 19637 -27155
rect 19675 -27189 19679 -27155
rect 19679 -27189 19709 -27155
rect 19747 -27189 19781 -27155
rect 19819 -27189 19849 -27155
rect 19849 -27189 19853 -27155
rect 19891 -27189 19917 -27155
rect 19917 -27189 19925 -27155
rect 19963 -27189 19985 -27155
rect 19985 -27189 19997 -27155
rect 20035 -27189 20053 -27155
rect 20053 -27189 20069 -27155
rect 20107 -27189 20121 -27155
rect 20121 -27189 20141 -27155
rect 20179 -27189 20189 -27155
rect 20189 -27189 20213 -27155
rect 20251 -27189 20257 -27155
rect 20257 -27189 20285 -27155
rect 20323 -27189 20325 -27155
rect 20325 -27189 20357 -27155
rect 20395 -27189 20427 -27155
rect 20427 -27189 20429 -27155
rect 20467 -27189 20495 -27155
rect 20495 -27189 20501 -27155
rect 20539 -27189 20563 -27155
rect 20563 -27189 20573 -27155
rect 20611 -27189 20631 -27155
rect 20631 -27189 20645 -27155
rect 20683 -27189 20699 -27155
rect 20699 -27189 20717 -27155
rect 20755 -27189 20767 -27155
rect 20767 -27189 20789 -27155
rect 20827 -27189 20835 -27155
rect 20835 -27189 20861 -27155
rect 20899 -27189 20903 -27155
rect 20903 -27189 20933 -27155
rect 20971 -27189 21005 -27155
rect 21043 -27189 21073 -27155
rect 21073 -27189 21077 -27155
rect 21115 -27189 21141 -27155
rect 21141 -27189 21149 -27155
rect 21187 -27189 21209 -27155
rect 21209 -27189 21221 -27155
rect 21259 -27189 21277 -27155
rect 21277 -27189 21293 -27155
rect 21331 -27189 21345 -27155
rect 21345 -27189 21365 -27155
rect 21403 -27189 21413 -27155
rect 21413 -27189 21437 -27155
rect 21475 -27189 21481 -27155
rect 21481 -27189 21509 -27155
rect 21547 -27189 21549 -27155
rect 21549 -27189 21581 -27155
rect 21619 -27189 21651 -27155
rect 21651 -27189 21653 -27155
rect 21691 -27189 21719 -27155
rect 21719 -27189 21725 -27155
rect 21763 -27189 21787 -27155
rect 21787 -27189 21797 -27155
rect 21835 -27189 21855 -27155
rect 21855 -27189 21869 -27155
rect 21907 -27189 21923 -27155
rect 21923 -27189 21941 -27155
rect 21979 -27189 21991 -27155
rect 21991 -27189 22013 -27155
rect 22051 -27189 22059 -27155
rect 22059 -27189 22085 -27155
rect 22123 -27189 22127 -27155
rect 22127 -27189 22157 -27155
rect 22195 -27189 22229 -27155
rect 22267 -27189 22297 -27155
rect 22297 -27189 22301 -27155
rect 22339 -27189 22365 -27155
rect 22365 -27189 22373 -27155
rect 22411 -27189 22433 -27155
rect 22433 -27189 22445 -27155
rect 22483 -27189 22501 -27155
rect 22501 -27189 22517 -27155
rect 22555 -27189 22569 -27155
rect 22569 -27189 22589 -27155
rect 22627 -27189 22637 -27155
rect 22637 -27189 22661 -27155
rect 22699 -27189 22705 -27155
rect 22705 -27189 22733 -27155
rect 22771 -27189 22773 -27155
rect 22773 -27189 22805 -27155
rect 22843 -27189 22875 -27155
rect 22875 -27189 22877 -27155
rect 22915 -27189 22943 -27155
rect 22943 -27189 22949 -27155
rect 22987 -27189 23011 -27155
rect 23011 -27189 23021 -27155
rect 23059 -27189 23079 -27155
rect 23079 -27189 23093 -27155
rect 23131 -27189 23147 -27155
rect 23147 -27189 23165 -27155
rect 23203 -27189 23215 -27155
rect 23215 -27189 23237 -27155
rect 23275 -27189 23283 -27155
rect 23283 -27189 23309 -27155
rect 23347 -27189 23351 -27155
rect 23351 -27189 23381 -27155
rect 23419 -27189 23453 -27155
rect 23491 -27189 23521 -27155
rect 23521 -27189 23525 -27155
rect 23563 -27189 23589 -27155
rect 23589 -27189 23597 -27155
rect 23635 -27189 23657 -27155
rect 23657 -27189 23669 -27155
rect 23707 -27189 23725 -27155
rect 23725 -27189 23741 -27155
rect 23779 -27189 23793 -27155
rect 23793 -27189 23813 -27155
rect 23851 -27189 23861 -27155
rect 23861 -27189 23885 -27155
rect 23923 -27189 23929 -27155
rect 23929 -27189 23957 -27155
rect 23995 -27189 23997 -27155
rect 23997 -27189 24029 -27155
rect 24067 -27189 24099 -27155
rect 24099 -27189 24101 -27155
rect 24139 -27189 24167 -27155
rect 24167 -27189 24173 -27155
rect 24211 -27189 24235 -27155
rect 24235 -27189 24245 -27155
rect 24283 -27189 24303 -27155
rect 24303 -27189 24317 -27155
rect 24355 -27189 24371 -27155
rect 24371 -27189 24389 -27155
rect 24427 -27189 24439 -27155
rect 24439 -27189 24461 -27155
rect 24499 -27189 24507 -27155
rect 24507 -27189 24533 -27155
rect 24571 -27189 24575 -27155
rect 24575 -27189 24605 -27155
rect 24643 -27189 24677 -27155
rect 24715 -27189 24745 -27155
rect 24745 -27189 24749 -27155
rect 24787 -27189 24821 -27155
<< metal1 >>
rect 372 1689 24828 1728
rect 372 1655 487 1689
rect 521 1655 559 1689
rect 593 1655 631 1689
rect 665 1655 703 1689
rect 737 1655 775 1689
rect 809 1655 847 1689
rect 881 1655 919 1689
rect 953 1655 991 1689
rect 1025 1655 1063 1689
rect 1097 1655 1135 1689
rect 1169 1655 1207 1689
rect 1241 1655 1279 1689
rect 1313 1655 1351 1689
rect 1385 1655 1423 1689
rect 1457 1655 1495 1689
rect 1529 1655 1567 1689
rect 1601 1655 1639 1689
rect 1673 1655 1711 1689
rect 1745 1655 1783 1689
rect 1817 1655 1855 1689
rect 1889 1655 1927 1689
rect 1961 1655 1999 1689
rect 2033 1655 2071 1689
rect 2105 1655 2143 1689
rect 2177 1655 2215 1689
rect 2249 1655 2287 1689
rect 2321 1655 2359 1689
rect 2393 1655 2431 1689
rect 2465 1655 2503 1689
rect 2537 1655 2575 1689
rect 2609 1655 2647 1689
rect 2681 1655 2719 1689
rect 2753 1655 2791 1689
rect 2825 1655 2863 1689
rect 2897 1655 2935 1689
rect 2969 1655 3007 1689
rect 3041 1655 3079 1689
rect 3113 1655 3151 1689
rect 3185 1655 3223 1689
rect 3257 1655 3295 1689
rect 3329 1655 3367 1689
rect 3401 1655 3439 1689
rect 3473 1655 3511 1689
rect 3545 1655 3583 1689
rect 3617 1655 3655 1689
rect 3689 1655 3727 1689
rect 3761 1655 3799 1689
rect 3833 1655 3871 1689
rect 3905 1655 3943 1689
rect 3977 1655 4015 1689
rect 4049 1655 4087 1689
rect 4121 1655 4159 1689
rect 4193 1655 4231 1689
rect 4265 1655 4303 1689
rect 4337 1655 4375 1689
rect 4409 1655 4447 1689
rect 4481 1655 4519 1689
rect 4553 1655 4591 1689
rect 4625 1655 4663 1689
rect 4697 1655 4735 1689
rect 4769 1655 4807 1689
rect 4841 1655 4879 1689
rect 4913 1655 4951 1689
rect 4985 1655 5023 1689
rect 5057 1655 5095 1689
rect 5129 1655 5167 1689
rect 5201 1655 5239 1689
rect 5273 1655 5311 1689
rect 5345 1655 5383 1689
rect 5417 1655 5455 1689
rect 5489 1655 5527 1689
rect 5561 1655 5599 1689
rect 5633 1655 5671 1689
rect 5705 1655 5743 1689
rect 5777 1655 5815 1689
rect 5849 1655 5887 1689
rect 5921 1655 5959 1689
rect 5993 1655 6031 1689
rect 6065 1655 6103 1689
rect 6137 1655 6175 1689
rect 6209 1655 6247 1689
rect 6281 1655 6319 1689
rect 6353 1655 6391 1689
rect 6425 1655 6463 1689
rect 6497 1655 6535 1689
rect 6569 1655 6607 1689
rect 6641 1655 6679 1689
rect 6713 1655 6751 1689
rect 6785 1655 6823 1689
rect 6857 1655 6895 1689
rect 6929 1655 6967 1689
rect 7001 1655 7039 1689
rect 7073 1655 7111 1689
rect 7145 1655 7183 1689
rect 7217 1655 7255 1689
rect 7289 1655 7327 1689
rect 7361 1655 7399 1689
rect 7433 1655 7471 1689
rect 7505 1655 7543 1689
rect 7577 1655 7615 1689
rect 7649 1655 7687 1689
rect 7721 1655 7759 1689
rect 7793 1655 7831 1689
rect 7865 1655 7903 1689
rect 7937 1655 7975 1689
rect 8009 1655 8047 1689
rect 8081 1655 8119 1689
rect 8153 1655 8191 1689
rect 8225 1655 8263 1689
rect 8297 1655 8335 1689
rect 8369 1655 8407 1689
rect 8441 1655 8479 1689
rect 8513 1655 8551 1689
rect 8585 1655 8623 1689
rect 8657 1655 8695 1689
rect 8729 1655 8767 1689
rect 8801 1655 8839 1689
rect 8873 1655 8911 1689
rect 8945 1655 8983 1689
rect 9017 1655 9055 1689
rect 9089 1655 9127 1689
rect 9161 1655 9199 1689
rect 9233 1655 9271 1689
rect 9305 1655 9343 1689
rect 9377 1655 9415 1689
rect 9449 1655 9487 1689
rect 9521 1655 9559 1689
rect 9593 1655 9631 1689
rect 9665 1655 9703 1689
rect 9737 1655 9775 1689
rect 9809 1655 9847 1689
rect 9881 1655 9919 1689
rect 9953 1655 9991 1689
rect 10025 1655 10063 1689
rect 10097 1655 10135 1689
rect 10169 1655 10207 1689
rect 10241 1655 10279 1689
rect 10313 1655 10351 1689
rect 10385 1655 10423 1689
rect 10457 1655 10495 1689
rect 10529 1655 10567 1689
rect 10601 1655 10639 1689
rect 10673 1655 10711 1689
rect 10745 1655 10783 1689
rect 10817 1655 10855 1689
rect 10889 1655 10927 1689
rect 10961 1655 10999 1689
rect 11033 1655 11071 1689
rect 11105 1655 11143 1689
rect 11177 1655 11215 1689
rect 11249 1655 11287 1689
rect 11321 1655 11359 1689
rect 11393 1655 11431 1689
rect 11465 1655 11503 1689
rect 11537 1655 11575 1689
rect 11609 1655 11647 1689
rect 11681 1655 11719 1689
rect 11753 1655 11791 1689
rect 11825 1655 11863 1689
rect 11897 1655 11935 1689
rect 11969 1655 12007 1689
rect 12041 1655 12079 1689
rect 12113 1655 12151 1689
rect 12185 1655 12223 1689
rect 12257 1655 12295 1689
rect 12329 1655 12367 1689
rect 12401 1655 12439 1689
rect 12473 1655 12511 1689
rect 12545 1655 12583 1689
rect 12617 1655 12655 1689
rect 12689 1655 12727 1689
rect 12761 1655 12799 1689
rect 12833 1655 12871 1689
rect 12905 1655 12943 1689
rect 12977 1655 13015 1689
rect 13049 1655 13087 1689
rect 13121 1655 13159 1689
rect 13193 1655 13231 1689
rect 13265 1655 13303 1689
rect 13337 1655 13375 1689
rect 13409 1655 13447 1689
rect 13481 1655 13519 1689
rect 13553 1655 13591 1689
rect 13625 1655 13663 1689
rect 13697 1655 13735 1689
rect 13769 1655 13807 1689
rect 13841 1655 13879 1689
rect 13913 1655 13951 1689
rect 13985 1655 14023 1689
rect 14057 1655 14095 1689
rect 14129 1655 14167 1689
rect 14201 1655 14239 1689
rect 14273 1655 14311 1689
rect 14345 1655 14383 1689
rect 14417 1655 14455 1689
rect 14489 1655 14527 1689
rect 14561 1655 14599 1689
rect 14633 1655 14671 1689
rect 14705 1655 14743 1689
rect 14777 1655 14815 1689
rect 14849 1655 14887 1689
rect 14921 1655 14959 1689
rect 14993 1655 15031 1689
rect 15065 1655 15103 1689
rect 15137 1655 15175 1689
rect 15209 1655 15247 1689
rect 15281 1655 15319 1689
rect 15353 1655 15391 1689
rect 15425 1655 15463 1689
rect 15497 1655 15535 1689
rect 15569 1655 15607 1689
rect 15641 1655 15679 1689
rect 15713 1655 15751 1689
rect 15785 1655 15823 1689
rect 15857 1655 15895 1689
rect 15929 1655 15967 1689
rect 16001 1655 16039 1689
rect 16073 1655 16111 1689
rect 16145 1655 16183 1689
rect 16217 1655 16255 1689
rect 16289 1655 16327 1689
rect 16361 1655 16399 1689
rect 16433 1655 16471 1689
rect 16505 1655 16543 1689
rect 16577 1655 16615 1689
rect 16649 1655 16687 1689
rect 16721 1655 16759 1689
rect 16793 1655 16831 1689
rect 16865 1655 16903 1689
rect 16937 1655 16975 1689
rect 17009 1655 17047 1689
rect 17081 1655 17119 1689
rect 17153 1655 17191 1689
rect 17225 1655 17263 1689
rect 17297 1655 17335 1689
rect 17369 1655 17407 1689
rect 17441 1655 17479 1689
rect 17513 1655 17551 1689
rect 17585 1655 17623 1689
rect 17657 1655 17695 1689
rect 17729 1655 17767 1689
rect 17801 1655 17839 1689
rect 17873 1655 17911 1689
rect 17945 1655 17983 1689
rect 18017 1655 18055 1689
rect 18089 1655 18127 1689
rect 18161 1655 18199 1689
rect 18233 1655 18271 1689
rect 18305 1655 18343 1689
rect 18377 1655 18415 1689
rect 18449 1655 18487 1689
rect 18521 1655 18559 1689
rect 18593 1655 18631 1689
rect 18665 1655 18703 1689
rect 18737 1655 18775 1689
rect 18809 1655 18847 1689
rect 18881 1655 18919 1689
rect 18953 1655 18991 1689
rect 19025 1655 19063 1689
rect 19097 1655 19135 1689
rect 19169 1655 19207 1689
rect 19241 1655 19279 1689
rect 19313 1655 19351 1689
rect 19385 1655 19423 1689
rect 19457 1655 19495 1689
rect 19529 1655 19567 1689
rect 19601 1655 19639 1689
rect 19673 1655 19711 1689
rect 19745 1655 19783 1689
rect 19817 1655 19855 1689
rect 19889 1655 19927 1689
rect 19961 1655 19999 1689
rect 20033 1655 20071 1689
rect 20105 1655 20143 1689
rect 20177 1655 20215 1689
rect 20249 1655 20287 1689
rect 20321 1655 20359 1689
rect 20393 1655 20431 1689
rect 20465 1655 20503 1689
rect 20537 1655 20575 1689
rect 20609 1655 20647 1689
rect 20681 1655 20719 1689
rect 20753 1655 20791 1689
rect 20825 1655 20863 1689
rect 20897 1655 20935 1689
rect 20969 1655 21007 1689
rect 21041 1655 21079 1689
rect 21113 1655 21151 1689
rect 21185 1655 21223 1689
rect 21257 1655 21295 1689
rect 21329 1655 21367 1689
rect 21401 1655 21439 1689
rect 21473 1655 21511 1689
rect 21545 1655 21583 1689
rect 21617 1655 21655 1689
rect 21689 1655 21727 1689
rect 21761 1655 21799 1689
rect 21833 1655 21871 1689
rect 21905 1655 21943 1689
rect 21977 1655 22015 1689
rect 22049 1655 22087 1689
rect 22121 1655 22159 1689
rect 22193 1655 22231 1689
rect 22265 1655 22303 1689
rect 22337 1655 22375 1689
rect 22409 1655 22447 1689
rect 22481 1655 22519 1689
rect 22553 1655 22591 1689
rect 22625 1655 22663 1689
rect 22697 1655 22735 1689
rect 22769 1655 22807 1689
rect 22841 1655 22879 1689
rect 22913 1655 22951 1689
rect 22985 1655 23023 1689
rect 23057 1655 23095 1689
rect 23129 1655 23167 1689
rect 23201 1655 23239 1689
rect 23273 1655 23311 1689
rect 23345 1655 23383 1689
rect 23417 1655 23455 1689
rect 23489 1655 23527 1689
rect 23561 1655 23599 1689
rect 23633 1655 23671 1689
rect 23705 1655 23743 1689
rect 23777 1655 23815 1689
rect 23849 1655 23887 1689
rect 23921 1655 23959 1689
rect 23993 1655 24031 1689
rect 24065 1655 24103 1689
rect 24137 1655 24175 1689
rect 24209 1655 24247 1689
rect 24281 1655 24319 1689
rect 24353 1655 24391 1689
rect 24425 1655 24463 1689
rect 24497 1655 24535 1689
rect 24569 1655 24607 1689
rect 24641 1655 24679 1689
rect 24713 1655 24828 1689
rect 372 1616 24828 1655
rect 372 1588 1094 1616
rect 372 1344 502 1588
rect 1066 1344 1094 1588
rect 372 1316 1094 1344
rect 24106 1588 24828 1616
rect 24106 1344 24134 1588
rect 24698 1344 24828 1588
rect 24106 1316 24828 1344
rect 372 1081 484 1316
rect 372 1047 411 1081
rect 445 1047 484 1081
rect 372 1009 484 1047
rect 372 975 411 1009
rect 445 975 484 1009
rect 3998 1217 20878 1266
rect 3998 1037 4075 1217
rect 20831 1037 20878 1217
rect 3998 1000 20878 1037
rect 24716 1081 24828 1316
rect 24716 1047 24755 1081
rect 24789 1047 24828 1081
rect 24716 1009 24828 1047
rect 3998 998 8352 1000
rect 372 937 484 975
rect 372 903 411 937
rect 445 903 484 937
rect 372 865 484 903
rect 372 831 411 865
rect 445 831 484 865
rect 372 793 484 831
rect 372 759 411 793
rect 445 759 484 793
rect 372 721 484 759
rect 372 687 411 721
rect 445 687 484 721
rect 372 649 484 687
rect 372 615 411 649
rect 445 615 484 649
rect 372 577 484 615
rect 372 543 411 577
rect 445 543 484 577
rect 372 505 484 543
rect 372 471 411 505
rect 445 471 484 505
rect 372 433 484 471
rect 372 399 411 433
rect 445 399 484 433
rect 372 361 484 399
rect 372 327 411 361
rect 445 327 484 361
rect 372 289 484 327
rect 372 255 411 289
rect 445 255 484 289
rect 372 217 484 255
rect 372 183 411 217
rect 445 183 484 217
rect 372 145 484 183
rect 372 111 411 145
rect 445 111 484 145
rect 372 73 484 111
rect 372 39 411 73
rect 445 39 484 73
rect 372 1 484 39
rect 372 -33 411 1
rect 445 -33 484 1
rect 372 -71 484 -33
rect 372 -105 411 -71
rect 445 -105 484 -71
rect 372 -143 484 -105
rect 372 -177 411 -143
rect 445 -177 484 -143
rect 372 -215 484 -177
rect 372 -249 411 -215
rect 445 -249 484 -215
rect 372 -287 484 -249
rect 372 -321 411 -287
rect 445 -321 484 -287
rect 372 -359 484 -321
rect 372 -393 411 -359
rect 445 -393 484 -359
rect 372 -431 484 -393
rect 372 -465 411 -431
rect 445 -465 484 -431
rect 372 -503 484 -465
rect 372 -537 411 -503
rect 445 -537 484 -503
rect 372 -575 484 -537
rect 372 -609 411 -575
rect 445 -609 484 -575
rect 372 -647 484 -609
rect 372 -681 411 -647
rect 445 -681 484 -647
rect 372 -719 484 -681
rect 372 -753 411 -719
rect 445 -753 484 -719
rect 372 -791 484 -753
rect 372 -825 411 -791
rect 445 -825 484 -791
rect 372 -863 484 -825
rect 372 -897 411 -863
rect 445 -897 484 -863
rect 372 -935 484 -897
rect 372 -969 411 -935
rect 445 -969 484 -935
rect 372 -1007 484 -969
rect 372 -1041 411 -1007
rect 445 -1041 484 -1007
rect 372 -1079 484 -1041
rect 372 -1113 411 -1079
rect 445 -1113 484 -1079
rect 372 -1151 484 -1113
rect 372 -1185 411 -1151
rect 445 -1185 484 -1151
rect 372 -1223 484 -1185
rect 372 -1257 411 -1223
rect 445 -1257 484 -1223
rect 372 -1295 484 -1257
rect 372 -1329 411 -1295
rect 445 -1329 484 -1295
rect 372 -1367 484 -1329
rect 372 -1401 411 -1367
rect 445 -1401 484 -1367
rect 372 -1439 484 -1401
rect 372 -1473 411 -1439
rect 445 -1473 484 -1439
rect 372 -1511 484 -1473
rect 372 -1545 411 -1511
rect 445 -1545 484 -1511
rect 372 -1583 484 -1545
rect 372 -1617 411 -1583
rect 445 -1617 484 -1583
rect 372 -1655 484 -1617
rect 372 -1689 411 -1655
rect 445 -1689 484 -1655
rect 372 -1727 484 -1689
rect 372 -1761 411 -1727
rect 445 -1761 484 -1727
rect 372 -1799 484 -1761
rect 372 -1833 411 -1799
rect 445 -1833 484 -1799
rect 372 -1871 484 -1833
rect 372 -1905 411 -1871
rect 445 -1905 484 -1871
rect 372 -1943 484 -1905
rect 372 -1977 411 -1943
rect 445 -1977 484 -1943
rect 372 -2015 484 -1977
rect 372 -2049 411 -2015
rect 445 -2049 484 -2015
rect 372 -2087 484 -2049
rect 372 -2121 411 -2087
rect 445 -2121 484 -2087
rect 372 -2159 484 -2121
rect 372 -2193 411 -2159
rect 445 -2193 484 -2159
rect 372 -2231 484 -2193
rect 372 -2265 411 -2231
rect 445 -2265 484 -2231
rect 372 -2303 484 -2265
rect 372 -2337 411 -2303
rect 445 -2337 484 -2303
rect 372 -2375 484 -2337
rect 372 -2409 411 -2375
rect 445 -2409 484 -2375
rect 372 -2447 484 -2409
rect 372 -2481 411 -2447
rect 445 -2481 484 -2447
rect 372 -2519 484 -2481
rect 372 -2553 411 -2519
rect 445 -2553 484 -2519
rect 372 -2591 484 -2553
rect 372 -2625 411 -2591
rect 445 -2625 484 -2591
rect 372 -2663 484 -2625
rect 372 -2697 411 -2663
rect 445 -2697 484 -2663
rect 372 -2735 484 -2697
rect 372 -2769 411 -2735
rect 445 -2769 484 -2735
rect 372 -2807 484 -2769
rect 372 -2841 411 -2807
rect 445 -2841 484 -2807
rect 372 -2879 484 -2841
rect 372 -2913 411 -2879
rect 445 -2913 484 -2879
rect 372 -2951 484 -2913
rect 372 -2985 411 -2951
rect 445 -2985 484 -2951
rect 372 -3023 484 -2985
rect 372 -3057 411 -3023
rect 445 -3057 484 -3023
rect 372 -3095 484 -3057
rect 372 -3129 411 -3095
rect 445 -3129 484 -3095
rect 372 -3167 484 -3129
rect 372 -3201 411 -3167
rect 445 -3201 484 -3167
rect 372 -3239 484 -3201
rect 372 -3273 411 -3239
rect 445 -3273 484 -3239
rect 372 -3311 484 -3273
rect 372 -3345 411 -3311
rect 445 -3345 484 -3311
rect 372 -3383 484 -3345
rect 372 -3417 411 -3383
rect 445 -3417 484 -3383
rect 372 -3455 484 -3417
rect 372 -3489 411 -3455
rect 445 -3489 484 -3455
rect 372 -3527 484 -3489
rect 372 -3561 411 -3527
rect 445 -3561 484 -3527
rect 372 -3599 484 -3561
rect 372 -3633 411 -3599
rect 445 -3633 484 -3599
rect 372 -3671 484 -3633
rect 372 -3705 411 -3671
rect 445 -3705 484 -3671
rect 372 -3743 484 -3705
rect 372 -3777 411 -3743
rect 445 -3777 484 -3743
rect 372 -3815 484 -3777
rect 372 -3849 411 -3815
rect 445 -3849 484 -3815
rect 372 -3887 484 -3849
rect 372 -3921 411 -3887
rect 445 -3921 484 -3887
rect 372 -3959 484 -3921
rect 372 -3993 411 -3959
rect 445 -3993 484 -3959
rect 372 -4031 484 -3993
rect 372 -4065 411 -4031
rect 445 -4065 484 -4031
rect 372 -4103 484 -4065
rect 372 -4137 411 -4103
rect 445 -4137 484 -4103
rect 372 -4175 484 -4137
rect 372 -4209 411 -4175
rect 445 -4209 484 -4175
rect 372 -4247 484 -4209
rect 372 -4281 411 -4247
rect 445 -4281 484 -4247
rect 372 -4319 484 -4281
rect 372 -4353 411 -4319
rect 445 -4353 484 -4319
rect 372 -4391 484 -4353
rect 372 -4425 411 -4391
rect 445 -4425 484 -4391
rect 372 -4463 484 -4425
rect 372 -4497 411 -4463
rect 445 -4497 484 -4463
rect 372 -4535 484 -4497
rect 372 -4569 411 -4535
rect 445 -4569 484 -4535
rect 372 -4607 484 -4569
rect 372 -4641 411 -4607
rect 445 -4641 484 -4607
rect 372 -4679 484 -4641
rect 372 -4713 411 -4679
rect 445 -4713 484 -4679
rect 372 -4751 484 -4713
rect 3614 -4562 4002 -4502
rect 3614 -4729 3674 -4562
rect 3716 -4603 3776 -4562
rect 3708 -4609 3796 -4603
rect 3708 -4643 3735 -4609
rect 3769 -4643 3796 -4609
rect 3708 -4649 3796 -4643
rect 3614 -4730 3626 -4729
rect 372 -4785 411 -4751
rect 445 -4785 484 -4751
rect 372 -4823 484 -4785
rect 372 -4857 411 -4823
rect 445 -4857 484 -4823
rect 372 -4895 484 -4857
rect 372 -4929 411 -4895
rect 445 -4929 484 -4895
rect 372 -4967 484 -4929
rect 372 -5001 411 -4967
rect 445 -5001 484 -4967
rect 372 -5039 484 -5001
rect 372 -5073 411 -5039
rect 445 -5073 484 -5039
rect 372 -5111 484 -5073
rect 3620 -4763 3626 -4730
rect 3660 -4730 3674 -4729
rect 3832 -4729 3892 -4562
rect 3942 -4603 4002 -4562
rect 3926 -4609 4014 -4603
rect 3926 -4643 3953 -4609
rect 3987 -4643 4014 -4609
rect 3926 -4649 4014 -4643
rect 3660 -4763 3666 -4730
rect 3832 -4734 3844 -4729
rect 3620 -4801 3666 -4763
rect 3620 -4835 3626 -4801
rect 3660 -4835 3666 -4801
rect 3620 -4873 3666 -4835
rect 3620 -4907 3626 -4873
rect 3660 -4907 3666 -4873
rect 3620 -4945 3666 -4907
rect 3620 -4979 3626 -4945
rect 3660 -4979 3666 -4945
rect 3620 -5017 3666 -4979
rect 3620 -5051 3626 -5017
rect 3660 -5051 3666 -5017
rect 3838 -4763 3844 -4734
rect 3878 -4734 3892 -4729
rect 4048 -4729 4108 998
rect 4150 -4506 4222 -4502
rect 4150 -4558 4160 -4506
rect 4212 -4558 4222 -4506
rect 4150 -4562 4222 -4558
rect 4262 -4506 4334 -4502
rect 4262 -4558 4272 -4506
rect 4324 -4558 4334 -4506
rect 4262 -4562 4334 -4558
rect 4372 -4506 4444 -4502
rect 4372 -4558 4382 -4506
rect 4434 -4558 4444 -4506
rect 4372 -4562 4444 -4558
rect 4156 -4603 4216 -4562
rect 4144 -4609 4232 -4603
rect 4144 -4643 4171 -4609
rect 4205 -4643 4232 -4609
rect 4144 -4649 4232 -4643
rect 4268 -4728 4328 -4562
rect 4378 -4603 4438 -4562
rect 4362 -4609 4376 -4603
rect 4378 -4609 4450 -4603
rect 4362 -4643 4389 -4609
rect 4423 -4643 4450 -4609
rect 4362 -4649 4450 -4643
rect 3878 -4763 3884 -4734
rect 3838 -4801 3884 -4763
rect 3838 -4835 3844 -4801
rect 3878 -4835 3884 -4801
rect 3838 -4873 3884 -4835
rect 3838 -4907 3844 -4873
rect 3878 -4907 3884 -4873
rect 3838 -4945 3884 -4907
rect 3838 -4979 3844 -4945
rect 3878 -4979 3884 -4945
rect 3838 -5017 3884 -4979
rect 3838 -5048 3844 -5017
rect 3620 -5090 3666 -5051
rect 3832 -5051 3844 -5048
rect 3878 -5048 3884 -5017
rect 4048 -4763 4062 -4729
rect 4096 -4763 4108 -4729
rect 4048 -4801 4108 -4763
rect 4048 -4835 4062 -4801
rect 4096 -4835 4108 -4801
rect 4048 -4873 4108 -4835
rect 4048 -4907 4062 -4873
rect 4096 -4907 4108 -4873
rect 4048 -4945 4108 -4907
rect 4048 -4979 4062 -4945
rect 4096 -4979 4108 -4945
rect 4048 -5017 4108 -4979
rect 3878 -5051 3892 -5048
rect 372 -5145 411 -5111
rect 445 -5145 484 -5111
rect 372 -5183 484 -5145
rect 3708 -5137 3796 -5131
rect 3708 -5171 3735 -5137
rect 3769 -5171 3796 -5137
rect 3708 -5177 3796 -5171
rect 372 -5217 411 -5183
rect 445 -5217 484 -5183
rect 3832 -5214 3892 -5051
rect 4048 -5051 4062 -5017
rect 4096 -5051 4108 -5017
rect 3926 -5137 4014 -5131
rect 3926 -5171 3953 -5137
rect 3987 -5171 4014 -5137
rect 3926 -5177 4014 -5171
rect 3942 -5214 4002 -5177
rect 372 -5255 484 -5217
rect 372 -5289 411 -5255
rect 445 -5289 484 -5255
rect 3486 -5218 3558 -5214
rect 3486 -5270 3496 -5218
rect 3548 -5270 3558 -5218
rect 3486 -5274 3558 -5270
rect 3826 -5218 3898 -5214
rect 3826 -5270 3836 -5218
rect 3888 -5270 3898 -5218
rect 3826 -5274 3898 -5270
rect 3936 -5218 4008 -5214
rect 3936 -5270 3946 -5218
rect 3998 -5270 4008 -5218
rect 3936 -5274 4008 -5270
rect 372 -5327 484 -5289
rect 372 -5361 411 -5327
rect 445 -5361 484 -5327
rect 372 -5399 484 -5361
rect 372 -5433 411 -5399
rect 445 -5433 484 -5399
rect 372 -5471 484 -5433
rect 372 -5505 411 -5471
rect 445 -5505 484 -5471
rect 372 -5543 484 -5505
rect 372 -5577 411 -5543
rect 445 -5577 484 -5543
rect 372 -5615 484 -5577
rect 372 -5649 411 -5615
rect 445 -5649 484 -5615
rect 372 -5687 484 -5649
rect 372 -5721 411 -5687
rect 445 -5721 484 -5687
rect 372 -5759 484 -5721
rect 372 -5793 411 -5759
rect 445 -5793 484 -5759
rect 372 -5831 484 -5793
rect 372 -5865 411 -5831
rect 445 -5865 484 -5831
rect 372 -5903 484 -5865
rect 372 -5937 411 -5903
rect 445 -5937 484 -5903
rect 372 -5975 484 -5937
rect 372 -6009 411 -5975
rect 445 -6009 484 -5975
rect 372 -6047 484 -6009
rect 372 -6081 411 -6047
rect 445 -6081 484 -6047
rect 372 -6119 484 -6081
rect 372 -6153 411 -6119
rect 445 -6153 484 -6119
rect 372 -6191 484 -6153
rect 372 -6225 411 -6191
rect 445 -6225 484 -6191
rect 2104 -6164 2176 -6160
rect 2104 -6216 2114 -6164
rect 2166 -6216 2176 -6164
rect 2104 -6220 2176 -6216
rect 372 -6263 484 -6225
rect 372 -6297 411 -6263
rect 445 -6297 484 -6263
rect 372 -6335 484 -6297
rect 372 -6369 411 -6335
rect 445 -6369 484 -6335
rect 372 -6407 484 -6369
rect 372 -6441 411 -6407
rect 445 -6441 484 -6407
rect 372 -6479 484 -6441
rect 372 -6513 411 -6479
rect 445 -6513 484 -6479
rect 372 -6551 484 -6513
rect 372 -6585 411 -6551
rect 445 -6585 484 -6551
rect 372 -6623 484 -6585
rect 372 -6657 411 -6623
rect 445 -6657 484 -6623
rect 372 -6695 484 -6657
rect 372 -6729 411 -6695
rect 445 -6729 484 -6695
rect 372 -6767 484 -6729
rect 372 -6801 411 -6767
rect 445 -6801 484 -6767
rect 372 -6839 484 -6801
rect 372 -6873 411 -6839
rect 445 -6873 484 -6839
rect 372 -6911 484 -6873
rect 372 -6945 411 -6911
rect 445 -6945 484 -6911
rect 372 -6983 484 -6945
rect 372 -7017 411 -6983
rect 445 -7017 484 -6983
rect 372 -7055 484 -7017
rect 372 -7089 411 -7055
rect 445 -7089 484 -7055
rect 372 -7127 484 -7089
rect 372 -7161 411 -7127
rect 445 -7161 484 -7127
rect 372 -7199 484 -7161
rect 372 -7233 411 -7199
rect 445 -7233 484 -7199
rect 372 -7271 484 -7233
rect 372 -7305 411 -7271
rect 445 -7305 484 -7271
rect 372 -7343 484 -7305
rect 372 -7377 411 -7343
rect 445 -7377 484 -7343
rect 372 -7415 484 -7377
rect 372 -7449 411 -7415
rect 445 -7449 484 -7415
rect 372 -7487 484 -7449
rect 372 -7521 411 -7487
rect 445 -7521 484 -7487
rect 372 -7559 484 -7521
rect 372 -7593 411 -7559
rect 445 -7593 484 -7559
rect 372 -7631 484 -7593
rect 372 -7665 411 -7631
rect 445 -7665 484 -7631
rect 372 -7703 484 -7665
rect 372 -7737 411 -7703
rect 445 -7737 484 -7703
rect 372 -7775 484 -7737
rect 372 -7809 411 -7775
rect 445 -7809 484 -7775
rect 372 -7847 484 -7809
rect 372 -7881 411 -7847
rect 445 -7881 484 -7847
rect 372 -7919 484 -7881
rect 372 -7953 411 -7919
rect 445 -7953 484 -7919
rect 372 -7991 484 -7953
rect 372 -8025 411 -7991
rect 445 -8025 484 -7991
rect 372 -8063 484 -8025
rect 372 -8097 411 -8063
rect 445 -8097 484 -8063
rect 372 -8135 484 -8097
rect 372 -8169 411 -8135
rect 445 -8169 484 -8135
rect 372 -8207 484 -8169
rect 372 -8241 411 -8207
rect 445 -8241 484 -8207
rect 372 -8776 484 -8241
rect 2110 -8392 2170 -6220
rect 3492 -7002 3552 -5274
rect 4048 -5320 4108 -5051
rect 4274 -4729 4320 -4728
rect 4274 -4763 4280 -4729
rect 4314 -4763 4320 -4729
rect 4274 -4801 4320 -4763
rect 4274 -4835 4280 -4801
rect 4314 -4835 4320 -4801
rect 4274 -4873 4320 -4835
rect 4274 -4907 4280 -4873
rect 4314 -4907 4320 -4873
rect 4274 -4945 4320 -4907
rect 4274 -4979 4280 -4945
rect 4314 -4979 4320 -4945
rect 4274 -5017 4320 -4979
rect 4274 -5051 4280 -5017
rect 4314 -5051 4320 -5017
rect 4274 -5090 4320 -5051
rect 4484 -4729 4544 998
rect 4580 -4609 4668 -4603
rect 4580 -4643 4607 -4609
rect 4641 -4643 4668 -4609
rect 4580 -4649 4668 -4643
rect 4798 -4609 4886 -4603
rect 4798 -4643 4825 -4609
rect 4859 -4643 4886 -4609
rect 4798 -4649 4886 -4643
rect 4484 -4763 4498 -4729
rect 4532 -4763 4544 -4729
rect 4484 -4801 4544 -4763
rect 4484 -4835 4498 -4801
rect 4532 -4835 4544 -4801
rect 4484 -4873 4544 -4835
rect 4484 -4907 4498 -4873
rect 4532 -4907 4544 -4873
rect 4484 -4945 4544 -4907
rect 4484 -4979 4498 -4945
rect 4532 -4979 4544 -4945
rect 4484 -5017 4544 -4979
rect 4484 -5051 4498 -5017
rect 4532 -5051 4544 -5017
rect 4710 -4729 4756 -4690
rect 4710 -4763 4716 -4729
rect 4750 -4763 4756 -4729
rect 4710 -4801 4756 -4763
rect 4710 -4835 4716 -4801
rect 4750 -4835 4756 -4801
rect 4710 -4873 4756 -4835
rect 4710 -4907 4716 -4873
rect 4750 -4907 4756 -4873
rect 4710 -4945 4756 -4907
rect 4710 -4979 4716 -4945
rect 4750 -4979 4756 -4945
rect 4710 -5017 4756 -4979
rect 4710 -5046 4716 -5017
rect 4144 -5137 4232 -5131
rect 4144 -5171 4171 -5137
rect 4205 -5171 4232 -5137
rect 4144 -5177 4232 -5171
rect 4362 -5137 4450 -5131
rect 4362 -5171 4389 -5137
rect 4423 -5171 4450 -5137
rect 4362 -5177 4450 -5171
rect 4484 -5320 4544 -5051
rect 4704 -5051 4716 -5046
rect 4750 -5046 4756 -5017
rect 4922 -4729 4982 998
rect 5022 -4506 5094 -4502
rect 5022 -4558 5032 -4506
rect 5084 -4558 5094 -4506
rect 5022 -4562 5094 -4558
rect 5132 -4506 5204 -4502
rect 5132 -4558 5142 -4506
rect 5194 -4558 5204 -4506
rect 5132 -4562 5204 -4558
rect 5240 -4506 5312 -4502
rect 5240 -4558 5250 -4506
rect 5302 -4558 5312 -4506
rect 5240 -4562 5312 -4558
rect 5028 -4603 5088 -4562
rect 5016 -4609 5088 -4603
rect 5090 -4609 5104 -4603
rect 5016 -4643 5043 -4609
rect 5077 -4643 5104 -4609
rect 5016 -4649 5104 -4643
rect 4922 -4763 4934 -4729
rect 4968 -4763 4982 -4729
rect 5138 -4729 5198 -4562
rect 5246 -4603 5306 -4562
rect 5234 -4609 5306 -4603
rect 5308 -4609 5322 -4603
rect 5234 -4643 5261 -4609
rect 5295 -4643 5322 -4609
rect 5234 -4649 5322 -4643
rect 5138 -4730 5152 -4729
rect 4922 -4801 4982 -4763
rect 4922 -4835 4934 -4801
rect 4968 -4835 4982 -4801
rect 4922 -4873 4982 -4835
rect 4922 -4907 4934 -4873
rect 4968 -4907 4982 -4873
rect 4922 -4945 4982 -4907
rect 4922 -4979 4934 -4945
rect 4968 -4979 4982 -4945
rect 4922 -5017 4982 -4979
rect 4750 -5051 4764 -5046
rect 4580 -5137 4668 -5131
rect 4580 -5171 4607 -5137
rect 4641 -5171 4668 -5137
rect 4580 -5177 4668 -5171
rect 4592 -5214 4652 -5177
rect 4704 -5214 4764 -5051
rect 4922 -5051 4934 -5017
rect 4968 -5051 4982 -5017
rect 4798 -5137 4886 -5131
rect 4798 -5171 4825 -5137
rect 4859 -5171 4886 -5137
rect 4798 -5177 4886 -5171
rect 4812 -5214 4872 -5177
rect 4586 -5218 4658 -5214
rect 4586 -5270 4596 -5218
rect 4648 -5270 4658 -5218
rect 4586 -5274 4658 -5270
rect 4698 -5218 4770 -5214
rect 4698 -5270 4708 -5218
rect 4760 -5270 4770 -5218
rect 4698 -5274 4770 -5270
rect 4806 -5218 4878 -5214
rect 4806 -5270 4816 -5218
rect 4868 -5270 4878 -5218
rect 4806 -5274 4878 -5270
rect 4922 -5320 4982 -5051
rect 5146 -4763 5152 -4730
rect 5186 -4730 5198 -4729
rect 5356 -4729 5416 998
rect 7980 880 8052 884
rect 7980 828 7990 880
rect 8042 828 8052 880
rect 7980 824 8052 828
rect 6474 608 7552 668
rect 6474 388 6534 608
rect 6978 492 7038 608
rect 7492 402 7552 608
rect 7986 484 8046 824
rect 8512 638 8572 1000
rect 9062 880 9134 884
rect 9062 828 9072 880
rect 9124 828 9134 880
rect 9062 824 9134 828
rect 10020 880 10092 884
rect 10020 828 10030 880
rect 10082 828 10092 880
rect 10020 824 10092 828
rect 8506 634 8578 638
rect 8506 582 8516 634
rect 8568 582 8578 634
rect 8506 578 8578 582
rect 8512 404 8572 578
rect 9068 482 9128 824
rect 10026 478 10086 824
rect 10548 638 10608 1000
rect 11056 880 11128 884
rect 11056 828 11066 880
rect 11118 828 11128 880
rect 11056 824 11128 828
rect 12062 880 12134 884
rect 12062 828 12072 880
rect 12124 828 12134 880
rect 12062 824 12134 828
rect 10542 634 10614 638
rect 10542 582 10552 634
rect 10604 582 10614 634
rect 10542 578 10614 582
rect 10548 404 10608 578
rect 11062 478 11122 824
rect 11560 746 11632 750
rect 11560 694 11570 746
rect 11622 694 11632 746
rect 11560 690 11632 694
rect 11566 400 11626 690
rect 12068 488 12128 824
rect 12586 640 12646 1000
rect 13084 880 13156 884
rect 13084 828 13094 880
rect 13146 828 13156 880
rect 13084 824 13156 828
rect 14102 880 14174 884
rect 14102 828 14112 880
rect 14164 828 14174 880
rect 14102 824 14174 828
rect 12580 636 12652 640
rect 12580 584 12590 636
rect 12642 584 12652 636
rect 12580 580 12652 584
rect 12586 388 12646 580
rect 13090 488 13150 824
rect 14108 482 14168 824
rect 14618 640 14678 1000
rect 15126 880 15198 884
rect 15126 828 15136 880
rect 15188 828 15198 880
rect 15126 824 15198 828
rect 16138 880 16210 884
rect 16138 828 16148 880
rect 16200 828 16210 880
rect 16138 824 16210 828
rect 14610 636 14682 640
rect 14610 584 14620 636
rect 14672 584 14682 636
rect 14610 580 14682 584
rect 14618 388 14678 580
rect 15132 488 15192 824
rect 16144 488 16204 824
rect 16658 642 16718 1000
rect 17156 880 17228 884
rect 17156 828 17166 880
rect 17218 828 17228 880
rect 17156 824 17228 828
rect 18168 880 18240 884
rect 18168 828 18178 880
rect 18230 828 18240 880
rect 18168 824 18240 828
rect 16652 638 16724 642
rect 16652 586 16662 638
rect 16714 586 16724 638
rect 16652 582 16724 586
rect 16658 390 16718 582
rect 17162 488 17222 824
rect 17664 746 17736 750
rect 17664 694 17674 746
rect 17726 694 17736 746
rect 17664 690 17736 694
rect 17670 386 17730 690
rect 18174 482 18234 824
rect 18690 642 18750 1000
rect 19196 880 19268 884
rect 19196 828 19206 880
rect 19258 828 19268 880
rect 19196 824 19268 828
rect 20208 880 20280 884
rect 20208 828 20218 880
rect 20270 828 20280 880
rect 20208 824 20280 828
rect 18684 638 18756 642
rect 18684 586 18694 638
rect 18746 586 18756 638
rect 18684 582 18756 586
rect 18690 400 18750 582
rect 19202 488 19262 824
rect 20214 488 20274 824
rect 20726 642 20786 1000
rect 24716 975 24755 1009
rect 24789 975 24828 1009
rect 24716 937 24828 975
rect 24716 903 24755 937
rect 24789 903 24828 937
rect 21226 880 21298 884
rect 21226 828 21236 880
rect 21288 828 21298 880
rect 21226 824 21298 828
rect 24716 865 24828 903
rect 24716 831 24755 865
rect 24789 831 24828 865
rect 20720 638 20792 642
rect 20720 586 20730 638
rect 20782 586 20792 638
rect 20720 582 20792 586
rect 20726 396 20786 582
rect 21232 482 21292 824
rect 24716 793 24828 831
rect 24716 759 24755 793
rect 24789 759 24828 793
rect 24716 721 24828 759
rect 24716 687 24755 721
rect 24789 687 24828 721
rect 21746 590 22826 650
rect 21746 398 21806 590
rect 22248 488 22308 590
rect 22766 382 22826 590
rect 24716 649 24828 687
rect 24716 615 24755 649
rect 24789 615 24828 649
rect 24716 577 24828 615
rect 24716 543 24755 577
rect 24789 543 24828 577
rect 24716 505 24828 543
rect 24716 471 24755 505
rect 24789 471 24828 505
rect 24716 433 24828 471
rect 24716 399 24755 433
rect 24789 399 24828 433
rect 24716 361 24828 399
rect 24716 327 24755 361
rect 24789 327 24828 361
rect 24716 289 24828 327
rect 24716 255 24755 289
rect 24789 255 24828 289
rect 24716 217 24828 255
rect 24716 183 24755 217
rect 24789 183 24828 217
rect 24716 145 24828 183
rect 24716 111 24755 145
rect 24789 111 24828 145
rect 24716 73 24828 111
rect 24716 39 24755 73
rect 24789 39 24828 73
rect 24716 1 24828 39
rect 24716 -33 24755 1
rect 24789 -33 24828 1
rect 24716 -71 24828 -33
rect 7494 -294 7554 -112
rect 6324 -298 6396 -294
rect 6324 -350 6334 -298
rect 6386 -350 6396 -298
rect 6324 -354 6396 -350
rect 7488 -298 7560 -294
rect 7488 -350 7498 -298
rect 7550 -350 7560 -298
rect 7488 -354 7560 -350
rect 6194 -502 6266 -498
rect 6194 -554 6204 -502
rect 6256 -554 6266 -502
rect 6194 -558 6266 -554
rect 6200 -3426 6260 -558
rect 6330 -2968 6390 -354
rect 7488 -502 7560 -498
rect 7488 -554 7498 -502
rect 7550 -554 7560 -502
rect 7488 -558 7560 -554
rect 7494 -746 7554 -558
rect 7998 -658 8058 -200
rect 8514 -748 8574 -108
rect 9020 -652 9080 -194
rect 9530 -398 9590 -120
rect 9524 -402 9596 -398
rect 9524 -454 9534 -402
rect 9586 -454 9596 -402
rect 9524 -458 9596 -454
rect 10050 -652 10110 -194
rect 10538 -738 10602 -90
rect 11050 -646 11110 -188
rect 11560 -402 11632 -398
rect 11560 -454 11570 -402
rect 11622 -454 11632 -402
rect 11560 -458 11632 -454
rect 11566 -746 11626 -458
rect 12068 -652 12128 -194
rect 12574 -742 12638 -94
rect 13092 -656 13152 -198
rect 13604 -294 13664 -108
rect 13598 -298 13670 -294
rect 13598 -350 13608 -298
rect 13660 -350 13670 -298
rect 13598 -354 13670 -350
rect 13594 -502 13666 -498
rect 13594 -554 13604 -502
rect 13656 -554 13666 -502
rect 13594 -558 13666 -554
rect 13600 -734 13660 -558
rect 14110 -650 14170 -192
rect 14616 -740 14680 -92
rect 15126 -658 15186 -195
rect 15638 -294 15698 -110
rect 15632 -298 15704 -294
rect 15632 -350 15642 -298
rect 15694 -350 15704 -298
rect 15632 -354 15704 -350
rect 15630 -502 15702 -498
rect 15630 -554 15640 -502
rect 15692 -554 15702 -502
rect 15630 -558 15702 -554
rect 15636 -740 15696 -558
rect 16138 -658 16198 -195
rect 16654 -756 16718 -108
rect 17144 -658 17204 -195
rect 17672 -300 17732 -116
rect 17672 -360 17874 -300
rect 17666 -402 17738 -398
rect 17666 -454 17676 -402
rect 17728 -454 17738 -402
rect 17666 -458 17738 -454
rect 17672 -732 17732 -458
rect 17814 -502 17874 -360
rect 17808 -506 17880 -502
rect 17808 -558 17818 -506
rect 17870 -558 17880 -506
rect 17808 -562 17880 -558
rect 18162 -658 18222 -195
rect 18690 -752 18750 -100
rect 24716 -105 24755 -71
rect 24789 -105 24828 -71
rect 19180 -658 19240 -195
rect 19706 -398 19766 -116
rect 19700 -402 19772 -398
rect 19700 -454 19710 -402
rect 19762 -454 19772 -402
rect 19700 -458 19772 -454
rect 19702 -506 19774 -502
rect 19702 -558 19712 -506
rect 19764 -558 19774 -506
rect 19702 -562 19774 -558
rect 19708 -736 19768 -562
rect 20180 -658 20240 -195
rect 20730 -744 20790 -110
rect 21210 -652 21270 -189
rect 21746 -294 21806 -108
rect 24716 -143 24828 -105
rect 24716 -177 24755 -143
rect 24789 -177 24828 -143
rect 24716 -215 24828 -177
rect 24716 -249 24755 -215
rect 24789 -249 24828 -215
rect 24716 -287 24828 -249
rect 21740 -298 21812 -294
rect 21740 -350 21750 -298
rect 21802 -350 21812 -298
rect 21740 -354 21812 -350
rect 22878 -298 22950 -294
rect 22878 -350 22888 -298
rect 22940 -350 22950 -298
rect 22878 -354 22950 -350
rect 24716 -321 24755 -287
rect 24789 -321 24828 -287
rect 21750 -570 22820 -510
rect 21750 -736 21810 -570
rect 22256 -644 22316 -570
rect 22760 -742 22820 -570
rect 14618 -1238 14678 -1236
rect 6476 -1434 6536 -1248
rect 6988 -1434 7048 -1346
rect 7494 -1434 7554 -1254
rect 10546 -1258 10606 -1256
rect 6476 -1494 7554 -1434
rect 7488 -1642 7548 -1636
rect 6478 -1702 7548 -1642
rect 6478 -1876 6538 -1702
rect 6988 -1778 7048 -1702
rect 7488 -1876 7548 -1702
rect 7980 -1788 8040 -1330
rect 8510 -1432 8570 -1258
rect 8504 -1436 8576 -1432
rect 8504 -1488 8514 -1436
rect 8566 -1488 8576 -1436
rect 8504 -1492 8576 -1488
rect 8510 -1896 8570 -1492
rect 9026 -1788 9086 -1330
rect 9528 -1528 9588 -1264
rect 10546 -1432 10610 -1258
rect 10540 -1436 10612 -1432
rect 10540 -1488 10550 -1436
rect 10602 -1488 10612 -1436
rect 10540 -1492 10612 -1488
rect 9522 -1532 9594 -1528
rect 9522 -1584 9532 -1532
rect 9584 -1584 9594 -1532
rect 9522 -1588 9594 -1584
rect 10226 -1536 10302 -1530
rect 10226 -1588 10238 -1536
rect 10290 -1588 10302 -1536
rect 10226 -1594 10302 -1588
rect 10232 -1624 10296 -1594
rect 9530 -1688 10296 -1624
rect 9530 -1890 9594 -1688
rect 10546 -1892 10610 -1492
rect 11074 -1782 11134 -1324
rect 11564 -1530 11628 -1248
rect 12580 -1250 12640 -1248
rect 11398 -1536 11628 -1530
rect 11398 -1588 11410 -1536
rect 11462 -1588 11628 -1536
rect 11398 -1594 11628 -1588
rect 11560 -1642 11632 -1638
rect 11560 -1694 11570 -1642
rect 11622 -1694 11632 -1642
rect 11560 -1698 11632 -1694
rect 11566 -1880 11626 -1698
rect 12092 -1792 12152 -1334
rect 12580 -1432 12644 -1250
rect 12574 -1436 12646 -1432
rect 12574 -1488 12584 -1436
rect 12636 -1488 12646 -1436
rect 12574 -1492 12646 -1488
rect 12580 -1904 12644 -1492
rect 13092 -1788 13152 -1330
rect 14120 -1798 14180 -1340
rect 14618 -1434 14682 -1238
rect 16654 -1242 16714 -1240
rect 14612 -1438 14684 -1434
rect 14612 -1490 14622 -1438
rect 14674 -1490 14684 -1438
rect 14612 -1494 14684 -1490
rect 14618 -1884 14682 -1494
rect 15138 -1788 15198 -1325
rect 15638 -1532 15698 -1254
rect 15632 -1536 15704 -1532
rect 15632 -1588 15642 -1536
rect 15694 -1588 15704 -1536
rect 15632 -1592 15704 -1588
rect 16138 -1792 16198 -1329
rect 16654 -1434 16718 -1242
rect 16648 -1438 16720 -1434
rect 16648 -1490 16658 -1438
rect 16710 -1490 16720 -1438
rect 16648 -1494 16720 -1490
rect 16654 -1896 16718 -1494
rect 17144 -1792 17204 -1329
rect 17666 -1642 17738 -1638
rect 17666 -1694 17676 -1642
rect 17728 -1694 17738 -1642
rect 17666 -1698 17738 -1694
rect 17672 -1880 17732 -1698
rect 18186 -1792 18246 -1329
rect 18690 -1434 18750 -1248
rect 18684 -1438 18756 -1434
rect 18684 -1490 18694 -1438
rect 18746 -1490 18756 -1438
rect 18684 -1494 18756 -1490
rect 18690 -1898 18750 -1494
rect 19186 -1788 19246 -1325
rect 19708 -1638 19768 -1248
rect 20724 -1254 20784 -1252
rect 19702 -1642 19774 -1638
rect 19702 -1694 19712 -1642
rect 19764 -1694 19774 -1642
rect 19702 -1698 19774 -1694
rect 20212 -1792 20272 -1329
rect 20724 -1436 20788 -1254
rect 20718 -1440 20790 -1436
rect 20718 -1492 20728 -1440
rect 20780 -1492 20790 -1440
rect 20718 -1496 20790 -1492
rect 20724 -1890 20788 -1496
rect 21210 -1794 21270 -1331
rect 21746 -1532 21806 -1254
rect 21740 -1536 21812 -1532
rect 21740 -1588 21750 -1536
rect 21802 -1588 21812 -1536
rect 21740 -1592 21812 -1588
rect 21748 -1646 21808 -1644
rect 21748 -1706 22820 -1646
rect 21748 -1870 21808 -1706
rect 22252 -1782 22312 -1706
rect 22760 -1894 22820 -1706
rect 7488 -2818 7552 -2378
rect 8510 -2570 8570 -2384
rect 10546 -2396 10606 -2394
rect 8504 -2574 8576 -2570
rect 8504 -2626 8514 -2574
rect 8566 -2626 8576 -2574
rect 8504 -2630 8576 -2626
rect 9526 -2680 9590 -2396
rect 9520 -2686 9596 -2680
rect 9520 -2738 9532 -2686
rect 9584 -2738 9596 -2686
rect 9520 -2744 9596 -2738
rect 7482 -2824 7558 -2818
rect 7482 -2876 7494 -2824
rect 7546 -2876 7558 -2824
rect 7482 -2882 7558 -2876
rect 6324 -2972 6396 -2968
rect 6324 -3024 6334 -2972
rect 6386 -3024 6396 -2972
rect 6324 -3028 6396 -3024
rect 7312 -2972 7372 -2962
rect 7312 -3024 7316 -2972
rect 7368 -3024 7372 -2972
rect 6916 -3308 6976 -3298
rect 6916 -3360 6920 -3308
rect 6972 -3360 6976 -3308
rect 6200 -3486 6862 -3426
rect 6042 -4506 6114 -4502
rect 5576 -4570 5856 -4510
rect 6042 -4558 6052 -4506
rect 6104 -4558 6114 -4506
rect 6042 -4562 6114 -4558
rect 5452 -4609 5540 -4603
rect 5452 -4643 5479 -4609
rect 5513 -4643 5540 -4609
rect 5452 -4649 5540 -4643
rect 5576 -4726 5636 -4570
rect 5684 -4603 5744 -4570
rect 5670 -4609 5758 -4603
rect 5670 -4643 5697 -4609
rect 5731 -4643 5758 -4609
rect 5670 -4649 5758 -4643
rect 5186 -4763 5192 -4730
rect 5146 -4801 5192 -4763
rect 5146 -4835 5152 -4801
rect 5186 -4835 5192 -4801
rect 5146 -4873 5192 -4835
rect 5146 -4907 5152 -4873
rect 5186 -4907 5192 -4873
rect 5146 -4945 5192 -4907
rect 5146 -4979 5152 -4945
rect 5186 -4979 5192 -4945
rect 5146 -5017 5192 -4979
rect 5146 -5051 5152 -5017
rect 5186 -5051 5192 -5017
rect 5146 -5090 5192 -5051
rect 5356 -4763 5370 -4729
rect 5404 -4763 5416 -4729
rect 5356 -4801 5416 -4763
rect 5356 -4835 5370 -4801
rect 5404 -4835 5416 -4801
rect 5356 -4873 5416 -4835
rect 5356 -4907 5370 -4873
rect 5404 -4907 5416 -4873
rect 5356 -4945 5416 -4907
rect 5356 -4979 5370 -4945
rect 5404 -4979 5416 -4945
rect 5356 -5017 5416 -4979
rect 5356 -5051 5370 -5017
rect 5404 -5051 5416 -5017
rect 5582 -4729 5628 -4726
rect 5582 -4763 5588 -4729
rect 5622 -4763 5628 -4729
rect 5796 -4729 5856 -4570
rect 5796 -4734 5806 -4729
rect 5582 -4801 5628 -4763
rect 5582 -4835 5588 -4801
rect 5622 -4835 5628 -4801
rect 5582 -4873 5628 -4835
rect 5582 -4907 5588 -4873
rect 5622 -4907 5628 -4873
rect 5582 -4945 5628 -4907
rect 5582 -4979 5588 -4945
rect 5622 -4979 5628 -4945
rect 5582 -5017 5628 -4979
rect 5582 -5032 5588 -5017
rect 5016 -5137 5104 -5131
rect 5016 -5171 5043 -5137
rect 5077 -5171 5104 -5137
rect 5016 -5177 5104 -5171
rect 5234 -5137 5322 -5131
rect 5234 -5171 5261 -5137
rect 5295 -5171 5322 -5137
rect 5234 -5177 5322 -5171
rect 5356 -5320 5416 -5051
rect 5574 -5051 5588 -5032
rect 5622 -5032 5628 -5017
rect 5800 -4763 5806 -4734
rect 5840 -4734 5856 -4729
rect 5840 -4763 5846 -4734
rect 5800 -4801 5846 -4763
rect 5800 -4835 5806 -4801
rect 5840 -4835 5846 -4801
rect 5800 -4873 5846 -4835
rect 5800 -4907 5806 -4873
rect 5840 -4907 5846 -4873
rect 5800 -4945 5846 -4907
rect 5800 -4979 5806 -4945
rect 5840 -4979 5846 -4945
rect 5800 -5017 5846 -4979
rect 5622 -5051 5634 -5032
rect 5452 -5137 5540 -5131
rect 5452 -5171 5479 -5137
rect 5513 -5171 5540 -5137
rect 5452 -5177 5540 -5171
rect 5464 -5214 5524 -5177
rect 5574 -5214 5634 -5051
rect 5800 -5051 5806 -5017
rect 5840 -5051 5846 -5017
rect 5800 -5090 5846 -5051
rect 5670 -5137 5758 -5131
rect 5670 -5171 5697 -5137
rect 5731 -5171 5758 -5137
rect 5670 -5177 5758 -5171
rect 5458 -5218 5530 -5214
rect 5458 -5270 5468 -5218
rect 5520 -5270 5530 -5218
rect 5458 -5274 5530 -5270
rect 5568 -5218 5640 -5214
rect 5568 -5270 5578 -5218
rect 5630 -5270 5640 -5218
rect 5568 -5274 5640 -5270
rect 4042 -5324 4114 -5320
rect 4042 -5376 4052 -5324
rect 4104 -5376 4114 -5324
rect 4042 -5380 4114 -5376
rect 4478 -5324 4550 -5320
rect 4478 -5376 4488 -5324
rect 4540 -5376 4550 -5324
rect 4478 -5380 4550 -5376
rect 4916 -5324 4988 -5320
rect 4916 -5376 4926 -5324
rect 4978 -5376 4988 -5324
rect 4916 -5380 4988 -5376
rect 5350 -5324 5422 -5320
rect 5350 -5376 5360 -5324
rect 5412 -5376 5422 -5324
rect 5350 -5380 5422 -5376
rect 3616 -5498 3892 -5438
rect 3616 -5667 3676 -5498
rect 3720 -5541 3780 -5498
rect 3708 -5547 3796 -5541
rect 3708 -5581 3735 -5547
rect 3769 -5581 3796 -5547
rect 3708 -5587 3796 -5581
rect 3616 -5674 3626 -5667
rect 3620 -5701 3626 -5674
rect 3660 -5674 3676 -5667
rect 3832 -5667 3892 -5498
rect 3926 -5547 4014 -5541
rect 3926 -5581 3953 -5547
rect 3987 -5581 4014 -5547
rect 3926 -5587 4014 -5581
rect 3832 -5670 3844 -5667
rect 3660 -5701 3666 -5674
rect 3620 -5739 3666 -5701
rect 3620 -5773 3626 -5739
rect 3660 -5773 3666 -5739
rect 3620 -5811 3666 -5773
rect 3620 -5845 3626 -5811
rect 3660 -5845 3666 -5811
rect 3620 -5883 3666 -5845
rect 3620 -5917 3626 -5883
rect 3660 -5917 3666 -5883
rect 3620 -5955 3666 -5917
rect 3620 -5989 3626 -5955
rect 3660 -5989 3666 -5955
rect 3838 -5701 3844 -5670
rect 3878 -5670 3892 -5667
rect 4048 -5667 4108 -5380
rect 4262 -5440 4334 -5436
rect 4262 -5492 4272 -5440
rect 4324 -5492 4334 -5440
rect 4262 -5496 4334 -5492
rect 4144 -5547 4232 -5541
rect 4144 -5581 4171 -5547
rect 4205 -5581 4232 -5547
rect 4144 -5587 4232 -5581
rect 4268 -5666 4328 -5496
rect 4362 -5547 4450 -5541
rect 4362 -5581 4389 -5547
rect 4423 -5581 4450 -5547
rect 4362 -5587 4450 -5581
rect 4048 -5668 4062 -5667
rect 3878 -5701 3884 -5670
rect 3838 -5739 3884 -5701
rect 3838 -5773 3844 -5739
rect 3878 -5773 3884 -5739
rect 3838 -5811 3884 -5773
rect 3838 -5845 3844 -5811
rect 3878 -5845 3884 -5811
rect 3838 -5883 3884 -5845
rect 3838 -5917 3844 -5883
rect 3878 -5917 3884 -5883
rect 3838 -5955 3884 -5917
rect 3838 -5982 3844 -5955
rect 3620 -6028 3666 -5989
rect 3832 -5989 3844 -5982
rect 3878 -5982 3884 -5955
rect 4056 -5701 4062 -5668
rect 4096 -5668 4108 -5667
rect 4274 -5667 4320 -5666
rect 4096 -5701 4102 -5668
rect 4056 -5739 4102 -5701
rect 4056 -5773 4062 -5739
rect 4096 -5773 4102 -5739
rect 4056 -5811 4102 -5773
rect 4056 -5845 4062 -5811
rect 4096 -5845 4102 -5811
rect 4056 -5883 4102 -5845
rect 4056 -5917 4062 -5883
rect 4096 -5917 4102 -5883
rect 4056 -5955 4102 -5917
rect 4056 -5974 4062 -5955
rect 3878 -5989 3892 -5982
rect 3708 -6075 3796 -6069
rect 3708 -6109 3735 -6075
rect 3769 -6109 3796 -6075
rect 3708 -6115 3796 -6109
rect 3832 -6160 3892 -5989
rect 4048 -5989 4062 -5974
rect 4096 -5974 4102 -5955
rect 4274 -5701 4280 -5667
rect 4314 -5701 4320 -5667
rect 4484 -5667 4544 -5380
rect 4580 -5547 4668 -5541
rect 4580 -5581 4607 -5547
rect 4641 -5581 4668 -5547
rect 4580 -5587 4668 -5581
rect 4798 -5547 4886 -5541
rect 4798 -5581 4825 -5547
rect 4859 -5581 4886 -5547
rect 4798 -5587 4886 -5581
rect 4484 -5670 4498 -5667
rect 4274 -5739 4320 -5701
rect 4274 -5773 4280 -5739
rect 4314 -5773 4320 -5739
rect 4274 -5811 4320 -5773
rect 4274 -5845 4280 -5811
rect 4314 -5845 4320 -5811
rect 4274 -5883 4320 -5845
rect 4274 -5917 4280 -5883
rect 4314 -5917 4320 -5883
rect 4274 -5955 4320 -5917
rect 4096 -5989 4108 -5974
rect 3926 -6075 4014 -6069
rect 3926 -6109 3953 -6075
rect 3987 -6109 4014 -6075
rect 3926 -6115 4014 -6109
rect 3826 -6164 3898 -6160
rect 3826 -6216 3836 -6164
rect 3888 -6216 3898 -6164
rect 3826 -6220 3898 -6216
rect 3942 -6358 4002 -6115
rect 4048 -6264 4108 -5989
rect 4274 -5989 4280 -5955
rect 4314 -5989 4320 -5955
rect 4492 -5701 4498 -5670
rect 4532 -5670 4544 -5667
rect 4710 -5667 4756 -5628
rect 4532 -5701 4538 -5670
rect 4492 -5739 4538 -5701
rect 4492 -5773 4498 -5739
rect 4532 -5773 4538 -5739
rect 4492 -5811 4538 -5773
rect 4492 -5845 4498 -5811
rect 4532 -5845 4538 -5811
rect 4492 -5883 4538 -5845
rect 4492 -5917 4498 -5883
rect 4532 -5917 4538 -5883
rect 4492 -5955 4538 -5917
rect 4492 -5984 4498 -5955
rect 4274 -6028 4320 -5989
rect 4484 -5989 4498 -5984
rect 4532 -5984 4538 -5955
rect 4710 -5701 4716 -5667
rect 4750 -5701 4756 -5667
rect 4922 -5667 4982 -5380
rect 5132 -5440 5204 -5436
rect 5132 -5492 5142 -5440
rect 5194 -5492 5204 -5440
rect 5132 -5496 5204 -5492
rect 5016 -5547 5104 -5541
rect 5016 -5581 5043 -5547
rect 5077 -5581 5104 -5547
rect 5016 -5587 5104 -5581
rect 4922 -5674 4934 -5667
rect 4710 -5739 4756 -5701
rect 4710 -5773 4716 -5739
rect 4750 -5773 4756 -5739
rect 4710 -5811 4756 -5773
rect 4710 -5845 4716 -5811
rect 4750 -5845 4756 -5811
rect 4710 -5883 4756 -5845
rect 4710 -5917 4716 -5883
rect 4750 -5917 4756 -5883
rect 4710 -5955 4756 -5917
rect 4710 -5980 4716 -5955
rect 4532 -5989 4544 -5984
rect 4144 -6075 4232 -6069
rect 4144 -6109 4171 -6075
rect 4205 -6109 4232 -6075
rect 4144 -6115 4232 -6109
rect 4362 -6075 4450 -6069
rect 4362 -6109 4389 -6075
rect 4423 -6109 4450 -6075
rect 4362 -6115 4450 -6109
rect 4042 -6268 4114 -6264
rect 4042 -6320 4052 -6268
rect 4104 -6320 4114 -6268
rect 4042 -6324 4114 -6320
rect 3614 -6362 4002 -6358
rect 3614 -6366 4008 -6362
rect 3614 -6418 3946 -6366
rect 3998 -6418 4008 -6366
rect 3614 -6604 3674 -6418
rect 3720 -6479 3780 -6418
rect 3708 -6485 3796 -6479
rect 3708 -6519 3735 -6485
rect 3769 -6519 3796 -6485
rect 3708 -6525 3796 -6519
rect 3620 -6605 3666 -6604
rect 3620 -6639 3626 -6605
rect 3660 -6639 3666 -6605
rect 3834 -6605 3894 -6418
rect 3936 -6422 4008 -6418
rect 3942 -6479 4002 -6422
rect 3926 -6485 4014 -6479
rect 3926 -6519 3953 -6485
rect 3987 -6519 4014 -6485
rect 3926 -6525 4014 -6519
rect 3834 -6616 3844 -6605
rect 3620 -6677 3666 -6639
rect 3620 -6711 3626 -6677
rect 3660 -6711 3666 -6677
rect 3620 -6749 3666 -6711
rect 3620 -6783 3626 -6749
rect 3660 -6783 3666 -6749
rect 3620 -6821 3666 -6783
rect 3620 -6855 3626 -6821
rect 3660 -6855 3666 -6821
rect 3620 -6893 3666 -6855
rect 3620 -6927 3626 -6893
rect 3660 -6927 3666 -6893
rect 3620 -6966 3666 -6927
rect 3838 -6639 3844 -6616
rect 3878 -6616 3894 -6605
rect 4048 -6605 4108 -6324
rect 4156 -6362 4216 -6115
rect 4260 -6164 4332 -6160
rect 4260 -6216 4270 -6164
rect 4322 -6216 4332 -6164
rect 4260 -6220 4332 -6216
rect 4150 -6366 4222 -6362
rect 4150 -6418 4160 -6366
rect 4212 -6418 4222 -6366
rect 4150 -6422 4222 -6418
rect 4156 -6479 4216 -6422
rect 4144 -6485 4232 -6479
rect 4144 -6519 4171 -6485
rect 4205 -6519 4232 -6485
rect 4144 -6525 4232 -6519
rect 4048 -6612 4062 -6605
rect 3878 -6639 3884 -6616
rect 3838 -6677 3884 -6639
rect 3838 -6711 3844 -6677
rect 3878 -6711 3884 -6677
rect 3838 -6749 3884 -6711
rect 3838 -6783 3844 -6749
rect 3878 -6783 3884 -6749
rect 3838 -6821 3884 -6783
rect 3838 -6855 3844 -6821
rect 3878 -6855 3884 -6821
rect 3838 -6893 3884 -6855
rect 3838 -6927 3844 -6893
rect 3878 -6927 3884 -6893
rect 3838 -6928 3884 -6927
rect 4056 -6639 4062 -6612
rect 4096 -6612 4108 -6605
rect 4266 -6605 4326 -6220
rect 4376 -6362 4436 -6115
rect 4484 -6264 4544 -5989
rect 4702 -5989 4716 -5980
rect 4750 -5980 4756 -5955
rect 4928 -5701 4934 -5674
rect 4968 -5674 4982 -5667
rect 5138 -5667 5198 -5496
rect 5234 -5547 5322 -5541
rect 5234 -5581 5261 -5547
rect 5295 -5581 5322 -5547
rect 5234 -5587 5322 -5581
rect 5356 -5662 5416 -5380
rect 5576 -5480 5856 -5420
rect 5452 -5547 5540 -5541
rect 5452 -5581 5479 -5547
rect 5513 -5581 5540 -5547
rect 5452 -5587 5540 -5581
rect 5138 -5672 5152 -5667
rect 4968 -5701 4974 -5674
rect 4928 -5739 4974 -5701
rect 4928 -5773 4934 -5739
rect 4968 -5773 4974 -5739
rect 4928 -5811 4974 -5773
rect 4928 -5845 4934 -5811
rect 4968 -5845 4974 -5811
rect 4928 -5883 4974 -5845
rect 4928 -5917 4934 -5883
rect 4968 -5917 4974 -5883
rect 4928 -5955 4974 -5917
rect 4750 -5989 4762 -5980
rect 4928 -5988 4934 -5955
rect 4580 -6075 4668 -6069
rect 4580 -6109 4607 -6075
rect 4641 -6109 4668 -6075
rect 4580 -6115 4668 -6109
rect 4478 -6268 4550 -6264
rect 4478 -6320 4488 -6268
rect 4540 -6320 4550 -6268
rect 4478 -6324 4550 -6320
rect 4370 -6366 4442 -6362
rect 4370 -6418 4380 -6366
rect 4432 -6418 4442 -6366
rect 4370 -6422 4442 -6418
rect 4376 -6479 4436 -6422
rect 4362 -6485 4450 -6479
rect 4362 -6519 4389 -6485
rect 4423 -6519 4450 -6485
rect 4362 -6525 4450 -6519
rect 4266 -6612 4280 -6605
rect 4096 -6639 4102 -6612
rect 4056 -6677 4102 -6639
rect 4056 -6711 4062 -6677
rect 4096 -6711 4102 -6677
rect 4056 -6749 4102 -6711
rect 4056 -6783 4062 -6749
rect 4096 -6783 4102 -6749
rect 4056 -6821 4102 -6783
rect 4056 -6855 4062 -6821
rect 4096 -6855 4102 -6821
rect 4056 -6893 4102 -6855
rect 4056 -6927 4062 -6893
rect 4096 -6927 4102 -6893
rect 3492 -7054 3496 -7002
rect 3548 -7054 3552 -7002
rect 3708 -7013 3796 -7007
rect 3708 -7047 3735 -7013
rect 3769 -7047 3796 -7013
rect 3708 -7053 3796 -7047
rect 3492 -7314 3552 -7054
rect 3832 -7098 3892 -6928
rect 4056 -6930 4102 -6927
rect 4274 -6639 4280 -6612
rect 4314 -6612 4326 -6605
rect 4484 -6605 4544 -6324
rect 4594 -6362 4654 -6115
rect 4702 -6160 4762 -5989
rect 4922 -5989 4934 -5988
rect 4968 -5988 4974 -5955
rect 5146 -5701 5152 -5672
rect 5186 -5672 5198 -5667
rect 5364 -5667 5410 -5662
rect 5576 -5664 5636 -5480
rect 5686 -5541 5746 -5480
rect 5670 -5547 5758 -5541
rect 5670 -5581 5697 -5547
rect 5731 -5581 5758 -5547
rect 5670 -5587 5758 -5581
rect 5186 -5701 5192 -5672
rect 5146 -5739 5192 -5701
rect 5146 -5773 5152 -5739
rect 5186 -5773 5192 -5739
rect 5146 -5811 5192 -5773
rect 5146 -5845 5152 -5811
rect 5186 -5845 5192 -5811
rect 5146 -5883 5192 -5845
rect 5146 -5917 5152 -5883
rect 5186 -5917 5192 -5883
rect 5146 -5955 5192 -5917
rect 4968 -5989 4982 -5988
rect 4798 -6075 4886 -6069
rect 4798 -6109 4825 -6075
rect 4859 -6109 4886 -6075
rect 4798 -6115 4886 -6109
rect 4696 -6164 4768 -6160
rect 4696 -6216 4706 -6164
rect 4758 -6216 4768 -6164
rect 4696 -6220 4768 -6216
rect 4810 -6362 4870 -6115
rect 4922 -6264 4982 -5989
rect 5146 -5989 5152 -5955
rect 5186 -5989 5192 -5955
rect 5364 -5701 5370 -5667
rect 5404 -5701 5410 -5667
rect 5364 -5739 5410 -5701
rect 5364 -5773 5370 -5739
rect 5404 -5773 5410 -5739
rect 5364 -5811 5410 -5773
rect 5364 -5845 5370 -5811
rect 5404 -5845 5410 -5811
rect 5364 -5883 5410 -5845
rect 5364 -5917 5370 -5883
rect 5404 -5917 5410 -5883
rect 5364 -5955 5410 -5917
rect 5364 -5986 5370 -5955
rect 5146 -6028 5192 -5989
rect 5356 -5989 5370 -5986
rect 5404 -5986 5410 -5955
rect 5582 -5667 5628 -5664
rect 5582 -5701 5588 -5667
rect 5622 -5701 5628 -5667
rect 5796 -5667 5856 -5480
rect 5926 -5440 5998 -5436
rect 5926 -5492 5936 -5440
rect 5988 -5492 5998 -5440
rect 5926 -5496 5998 -5492
rect 5796 -5676 5806 -5667
rect 5582 -5739 5628 -5701
rect 5582 -5773 5588 -5739
rect 5622 -5773 5628 -5739
rect 5582 -5811 5628 -5773
rect 5582 -5845 5588 -5811
rect 5622 -5845 5628 -5811
rect 5582 -5883 5628 -5845
rect 5582 -5917 5588 -5883
rect 5622 -5917 5628 -5883
rect 5582 -5955 5628 -5917
rect 5582 -5980 5588 -5955
rect 5404 -5989 5416 -5986
rect 5016 -6075 5104 -6069
rect 5016 -6109 5043 -6075
rect 5077 -6109 5104 -6075
rect 5016 -6115 5104 -6109
rect 5234 -6075 5322 -6069
rect 5234 -6109 5261 -6075
rect 5295 -6109 5322 -6075
rect 5234 -6115 5322 -6109
rect 4916 -6268 4988 -6264
rect 4916 -6320 4926 -6268
rect 4978 -6320 4988 -6268
rect 4916 -6324 4988 -6320
rect 4588 -6366 4660 -6362
rect 4588 -6418 4598 -6366
rect 4650 -6418 4660 -6366
rect 4588 -6422 4660 -6418
rect 4698 -6366 4770 -6362
rect 4698 -6418 4708 -6366
rect 4760 -6418 4770 -6366
rect 4698 -6422 4770 -6418
rect 4804 -6366 4876 -6362
rect 4804 -6418 4814 -6366
rect 4866 -6418 4876 -6366
rect 4804 -6422 4876 -6418
rect 4594 -6479 4654 -6422
rect 4580 -6485 4668 -6479
rect 4580 -6519 4607 -6485
rect 4641 -6519 4668 -6485
rect 4580 -6525 4668 -6519
rect 4314 -6639 4320 -6612
rect 4484 -6614 4498 -6605
rect 4274 -6677 4320 -6639
rect 4274 -6711 4280 -6677
rect 4314 -6711 4320 -6677
rect 4274 -6749 4320 -6711
rect 4274 -6783 4280 -6749
rect 4314 -6783 4320 -6749
rect 4274 -6821 4320 -6783
rect 4274 -6855 4280 -6821
rect 4314 -6855 4320 -6821
rect 4274 -6893 4320 -6855
rect 4274 -6927 4280 -6893
rect 4314 -6927 4320 -6893
rect 4492 -6639 4498 -6614
rect 4532 -6614 4544 -6605
rect 4704 -6605 4764 -6422
rect 4810 -6479 4870 -6422
rect 4798 -6485 4886 -6479
rect 4798 -6519 4825 -6485
rect 4859 -6519 4886 -6485
rect 4798 -6525 4886 -6519
rect 4704 -6606 4716 -6605
rect 4532 -6639 4538 -6614
rect 4492 -6677 4538 -6639
rect 4492 -6711 4498 -6677
rect 4532 -6711 4538 -6677
rect 4492 -6749 4538 -6711
rect 4492 -6783 4498 -6749
rect 4532 -6783 4538 -6749
rect 4492 -6821 4538 -6783
rect 4492 -6855 4498 -6821
rect 4532 -6855 4538 -6821
rect 4492 -6893 4538 -6855
rect 4492 -6916 4498 -6893
rect 3926 -7013 4014 -7007
rect 3926 -7047 3953 -7013
rect 3987 -7047 4014 -7013
rect 3926 -7053 4014 -7047
rect 3826 -7102 3898 -7098
rect 3826 -7154 3836 -7102
rect 3888 -7154 3898 -7102
rect 3826 -7158 3898 -7154
rect 4048 -7196 4108 -6930
rect 4274 -6966 4320 -6927
rect 4484 -6927 4498 -6916
rect 4532 -6916 4538 -6893
rect 4710 -6639 4716 -6606
rect 4750 -6606 4764 -6605
rect 4922 -6605 4982 -6324
rect 5028 -6362 5088 -6115
rect 5132 -6164 5204 -6160
rect 5132 -6216 5142 -6164
rect 5194 -6216 5204 -6164
rect 5132 -6220 5204 -6216
rect 5022 -6366 5094 -6362
rect 5022 -6418 5032 -6366
rect 5084 -6418 5094 -6366
rect 5022 -6422 5094 -6418
rect 5028 -6479 5088 -6422
rect 5016 -6485 5104 -6479
rect 5016 -6519 5043 -6485
rect 5077 -6519 5104 -6485
rect 5016 -6525 5104 -6519
rect 5138 -6604 5198 -6220
rect 5246 -6362 5306 -6115
rect 5356 -6264 5416 -5989
rect 5576 -5989 5588 -5980
rect 5622 -5980 5628 -5955
rect 5800 -5701 5806 -5676
rect 5840 -5676 5856 -5667
rect 5840 -5701 5846 -5676
rect 5800 -5739 5846 -5701
rect 5800 -5773 5806 -5739
rect 5840 -5773 5846 -5739
rect 5800 -5811 5846 -5773
rect 5800 -5845 5806 -5811
rect 5840 -5845 5846 -5811
rect 5800 -5883 5846 -5845
rect 5800 -5917 5806 -5883
rect 5840 -5917 5846 -5883
rect 5800 -5955 5846 -5917
rect 5622 -5989 5636 -5980
rect 5452 -6075 5540 -6069
rect 5452 -6109 5479 -6075
rect 5513 -6109 5540 -6075
rect 5452 -6115 5540 -6109
rect 5350 -6268 5422 -6264
rect 5350 -6320 5360 -6268
rect 5412 -6320 5422 -6268
rect 5350 -6324 5422 -6320
rect 5240 -6366 5312 -6362
rect 5240 -6418 5250 -6366
rect 5302 -6418 5312 -6366
rect 5240 -6422 5312 -6418
rect 5246 -6479 5306 -6422
rect 5234 -6485 5322 -6479
rect 5234 -6519 5261 -6485
rect 5295 -6519 5322 -6485
rect 5234 -6525 5322 -6519
rect 4750 -6639 4756 -6606
rect 4922 -6618 4934 -6605
rect 4710 -6677 4756 -6639
rect 4710 -6711 4716 -6677
rect 4750 -6711 4756 -6677
rect 4710 -6749 4756 -6711
rect 4710 -6783 4716 -6749
rect 4750 -6783 4756 -6749
rect 4710 -6821 4756 -6783
rect 4710 -6855 4716 -6821
rect 4750 -6855 4756 -6821
rect 4710 -6893 4756 -6855
rect 4532 -6927 4544 -6916
rect 4710 -6924 4716 -6893
rect 4144 -7013 4232 -7007
rect 4144 -7047 4171 -7013
rect 4205 -7047 4232 -7013
rect 4144 -7053 4232 -7047
rect 4362 -7013 4450 -7007
rect 4362 -7047 4389 -7013
rect 4423 -7047 4450 -7013
rect 4362 -7053 4450 -7047
rect 4484 -7196 4544 -6927
rect 4702 -6927 4716 -6924
rect 4750 -6924 4756 -6893
rect 4928 -6639 4934 -6618
rect 4968 -6618 4982 -6605
rect 5146 -6605 5192 -6604
rect 4968 -6639 4974 -6618
rect 4928 -6677 4974 -6639
rect 4928 -6711 4934 -6677
rect 4968 -6711 4974 -6677
rect 4928 -6749 4974 -6711
rect 4928 -6783 4934 -6749
rect 4968 -6783 4974 -6749
rect 4928 -6821 4974 -6783
rect 4928 -6855 4934 -6821
rect 4968 -6855 4974 -6821
rect 4928 -6893 4974 -6855
rect 4928 -6920 4934 -6893
rect 4750 -6927 4762 -6924
rect 4580 -7013 4668 -7007
rect 4580 -7047 4607 -7013
rect 4641 -7047 4668 -7013
rect 4580 -7053 4668 -7047
rect 4702 -7098 4762 -6927
rect 4922 -6927 4934 -6920
rect 4968 -6920 4974 -6893
rect 5146 -6639 5152 -6605
rect 5186 -6639 5192 -6605
rect 5356 -6605 5416 -6324
rect 5462 -6362 5522 -6115
rect 5576 -6160 5636 -5989
rect 5800 -5989 5806 -5955
rect 5840 -5989 5846 -5955
rect 5800 -6028 5846 -5989
rect 5670 -6075 5758 -6069
rect 5670 -6109 5697 -6075
rect 5731 -6109 5758 -6075
rect 5670 -6115 5758 -6109
rect 5570 -6164 5642 -6160
rect 5570 -6216 5580 -6164
rect 5632 -6216 5642 -6164
rect 5570 -6220 5642 -6216
rect 5456 -6366 5856 -6362
rect 5456 -6418 5466 -6366
rect 5518 -6418 5856 -6366
rect 5456 -6422 5856 -6418
rect 5462 -6479 5522 -6422
rect 5452 -6485 5540 -6479
rect 5452 -6519 5479 -6485
rect 5513 -6519 5540 -6485
rect 5452 -6525 5540 -6519
rect 5574 -6596 5634 -6422
rect 5682 -6479 5742 -6422
rect 5670 -6485 5758 -6479
rect 5670 -6519 5697 -6485
rect 5731 -6519 5758 -6485
rect 5670 -6525 5758 -6519
rect 5356 -6606 5370 -6605
rect 5146 -6677 5192 -6639
rect 5146 -6711 5152 -6677
rect 5186 -6711 5192 -6677
rect 5146 -6749 5192 -6711
rect 5146 -6783 5152 -6749
rect 5186 -6783 5192 -6749
rect 5146 -6821 5192 -6783
rect 5146 -6855 5152 -6821
rect 5186 -6855 5192 -6821
rect 5146 -6893 5192 -6855
rect 4968 -6927 4982 -6920
rect 4798 -7013 4886 -7007
rect 4798 -7047 4825 -7013
rect 4859 -7047 4886 -7013
rect 4798 -7053 4886 -7047
rect 4696 -7102 4768 -7098
rect 4696 -7154 4706 -7102
rect 4758 -7154 4768 -7102
rect 4696 -7158 4768 -7154
rect 4922 -7196 4982 -6927
rect 5146 -6927 5152 -6893
rect 5186 -6927 5192 -6893
rect 5364 -6639 5370 -6606
rect 5404 -6606 5416 -6605
rect 5582 -6605 5628 -6596
rect 5796 -6600 5856 -6422
rect 5404 -6639 5410 -6606
rect 5364 -6677 5410 -6639
rect 5364 -6711 5370 -6677
rect 5404 -6711 5410 -6677
rect 5364 -6749 5410 -6711
rect 5364 -6783 5370 -6749
rect 5404 -6783 5410 -6749
rect 5364 -6821 5410 -6783
rect 5364 -6855 5370 -6821
rect 5404 -6855 5410 -6821
rect 5364 -6893 5410 -6855
rect 5364 -6920 5370 -6893
rect 5146 -6966 5192 -6927
rect 5356 -6927 5370 -6920
rect 5404 -6920 5410 -6893
rect 5582 -6639 5588 -6605
rect 5622 -6639 5628 -6605
rect 5582 -6677 5628 -6639
rect 5582 -6711 5588 -6677
rect 5622 -6711 5628 -6677
rect 5582 -6749 5628 -6711
rect 5582 -6783 5588 -6749
rect 5622 -6783 5628 -6749
rect 5582 -6821 5628 -6783
rect 5582 -6855 5588 -6821
rect 5622 -6855 5628 -6821
rect 5582 -6893 5628 -6855
rect 5582 -6920 5588 -6893
rect 5404 -6927 5416 -6920
rect 5016 -7013 5104 -7007
rect 5016 -7047 5043 -7013
rect 5077 -7047 5104 -7013
rect 5016 -7053 5104 -7047
rect 5234 -7013 5322 -7007
rect 5234 -7047 5261 -7013
rect 5295 -7047 5322 -7013
rect 5234 -7053 5322 -7047
rect 5356 -7196 5416 -6927
rect 5576 -6927 5588 -6920
rect 5622 -6920 5628 -6893
rect 5800 -6605 5846 -6600
rect 5800 -6639 5806 -6605
rect 5840 -6639 5846 -6605
rect 5800 -6677 5846 -6639
rect 5800 -6711 5806 -6677
rect 5840 -6711 5846 -6677
rect 5800 -6749 5846 -6711
rect 5800 -6783 5806 -6749
rect 5840 -6783 5846 -6749
rect 5800 -6821 5846 -6783
rect 5800 -6855 5806 -6821
rect 5840 -6855 5846 -6821
rect 5800 -6893 5846 -6855
rect 5622 -6927 5636 -6920
rect 5452 -7013 5540 -7007
rect 5452 -7047 5479 -7013
rect 5513 -7047 5540 -7013
rect 5452 -7053 5540 -7047
rect 5576 -7098 5636 -6927
rect 5800 -6927 5806 -6893
rect 5840 -6927 5846 -6893
rect 5800 -6966 5846 -6927
rect 5670 -7013 5758 -7007
rect 5670 -7047 5697 -7013
rect 5731 -7047 5758 -7013
rect 5670 -7053 5758 -7047
rect 5932 -7098 5992 -5496
rect 5570 -7102 5642 -7098
rect 5570 -7154 5580 -7102
rect 5632 -7154 5642 -7102
rect 5570 -7158 5642 -7154
rect 5926 -7102 5998 -7098
rect 5926 -7154 5936 -7102
rect 5988 -7154 5998 -7102
rect 5926 -7158 5998 -7154
rect 4042 -7200 4114 -7196
rect 4042 -7252 4052 -7200
rect 4104 -7252 4114 -7200
rect 4042 -7256 4114 -7252
rect 4478 -7200 4550 -7196
rect 4478 -7252 4488 -7200
rect 4540 -7252 4550 -7200
rect 4478 -7256 4550 -7252
rect 4916 -7200 4988 -7196
rect 4916 -7252 4926 -7200
rect 4978 -7252 4988 -7200
rect 4916 -7256 4988 -7252
rect 5350 -7200 5422 -7196
rect 5350 -7252 5360 -7200
rect 5412 -7252 5422 -7200
rect 5350 -7256 5422 -7252
rect 3486 -7318 3558 -7314
rect 3486 -7370 3496 -7318
rect 3548 -7370 3558 -7318
rect 3486 -7374 3558 -7370
rect 3616 -7376 4002 -7316
rect 3616 -7543 3676 -7376
rect 3722 -7417 3782 -7376
rect 3708 -7423 3796 -7417
rect 3708 -7457 3735 -7423
rect 3769 -7457 3796 -7423
rect 3708 -7463 3796 -7457
rect 3832 -7540 3892 -7376
rect 3942 -7417 4002 -7376
rect 3926 -7423 4014 -7417
rect 3926 -7457 3953 -7423
rect 3987 -7457 4014 -7423
rect 3926 -7463 4014 -7457
rect 3616 -7546 3626 -7543
rect 3620 -7577 3626 -7546
rect 3660 -7546 3676 -7543
rect 3838 -7543 3884 -7540
rect 3660 -7577 3666 -7546
rect 3620 -7615 3666 -7577
rect 3620 -7649 3626 -7615
rect 3660 -7649 3666 -7615
rect 3620 -7687 3666 -7649
rect 3620 -7721 3626 -7687
rect 3660 -7721 3666 -7687
rect 3620 -7759 3666 -7721
rect 3620 -7793 3626 -7759
rect 3660 -7793 3666 -7759
rect 3620 -7831 3666 -7793
rect 3620 -7865 3626 -7831
rect 3660 -7865 3666 -7831
rect 3838 -7577 3844 -7543
rect 3878 -7577 3884 -7543
rect 4048 -7543 4108 -7256
rect 4152 -7318 4224 -7314
rect 4152 -7370 4162 -7318
rect 4214 -7370 4224 -7318
rect 4152 -7374 4224 -7370
rect 4260 -7318 4332 -7314
rect 4260 -7370 4270 -7318
rect 4322 -7370 4332 -7318
rect 4260 -7374 4332 -7370
rect 4368 -7318 4440 -7314
rect 4368 -7370 4378 -7318
rect 4430 -7370 4440 -7318
rect 4368 -7374 4440 -7370
rect 4158 -7417 4218 -7374
rect 4144 -7423 4232 -7417
rect 4144 -7457 4171 -7423
rect 4205 -7457 4232 -7423
rect 4144 -7463 4232 -7457
rect 4266 -7540 4326 -7374
rect 4374 -7417 4434 -7374
rect 4362 -7423 4450 -7417
rect 4362 -7457 4389 -7423
rect 4423 -7457 4450 -7423
rect 4362 -7463 4450 -7457
rect 4048 -7544 4062 -7543
rect 3838 -7615 3884 -7577
rect 3838 -7649 3844 -7615
rect 3878 -7649 3884 -7615
rect 3838 -7687 3884 -7649
rect 3838 -7721 3844 -7687
rect 3878 -7721 3884 -7687
rect 3838 -7759 3884 -7721
rect 3838 -7793 3844 -7759
rect 3878 -7793 3884 -7759
rect 3838 -7831 3884 -7793
rect 3838 -7864 3844 -7831
rect 3620 -7904 3666 -7865
rect 3832 -7865 3844 -7864
rect 3878 -7864 3884 -7831
rect 4056 -7577 4062 -7544
rect 4096 -7544 4108 -7543
rect 4274 -7543 4320 -7540
rect 4096 -7577 4102 -7544
rect 4056 -7615 4102 -7577
rect 4056 -7649 4062 -7615
rect 4096 -7649 4102 -7615
rect 4056 -7687 4102 -7649
rect 4056 -7721 4062 -7687
rect 4096 -7721 4102 -7687
rect 4056 -7759 4102 -7721
rect 4056 -7793 4062 -7759
rect 4096 -7793 4102 -7759
rect 4056 -7831 4102 -7793
rect 3878 -7865 3892 -7864
rect 3708 -7951 3796 -7945
rect 3708 -7985 3735 -7951
rect 3769 -7985 3796 -7951
rect 3708 -7991 3796 -7985
rect 3832 -8034 3892 -7865
rect 4056 -7865 4062 -7831
rect 4096 -7865 4102 -7831
rect 4056 -7904 4102 -7865
rect 4274 -7577 4280 -7543
rect 4314 -7577 4320 -7543
rect 4484 -7543 4544 -7256
rect 4580 -7423 4668 -7417
rect 4580 -7457 4607 -7423
rect 4641 -7457 4668 -7423
rect 4580 -7463 4668 -7457
rect 4798 -7423 4886 -7417
rect 4798 -7457 4825 -7423
rect 4859 -7457 4886 -7423
rect 4798 -7463 4886 -7457
rect 4484 -7546 4498 -7543
rect 4274 -7615 4320 -7577
rect 4274 -7649 4280 -7615
rect 4314 -7649 4320 -7615
rect 4274 -7687 4320 -7649
rect 4274 -7721 4280 -7687
rect 4314 -7721 4320 -7687
rect 4274 -7759 4320 -7721
rect 4274 -7793 4280 -7759
rect 4314 -7793 4320 -7759
rect 4274 -7831 4320 -7793
rect 4274 -7865 4280 -7831
rect 4314 -7865 4320 -7831
rect 4274 -7904 4320 -7865
rect 4492 -7577 4498 -7546
rect 4532 -7546 4544 -7543
rect 4710 -7543 4756 -7504
rect 4532 -7577 4538 -7546
rect 4492 -7615 4538 -7577
rect 4492 -7649 4498 -7615
rect 4532 -7649 4538 -7615
rect 4492 -7687 4538 -7649
rect 4492 -7721 4498 -7687
rect 4532 -7721 4538 -7687
rect 4492 -7759 4538 -7721
rect 4492 -7793 4498 -7759
rect 4532 -7793 4538 -7759
rect 4492 -7831 4538 -7793
rect 4492 -7865 4498 -7831
rect 4532 -7865 4538 -7831
rect 4710 -7577 4716 -7543
rect 4750 -7577 4756 -7543
rect 4922 -7543 4982 -7256
rect 5014 -7318 5086 -7314
rect 5014 -7370 5024 -7318
rect 5076 -7370 5086 -7318
rect 5014 -7374 5086 -7370
rect 5132 -7318 5204 -7314
rect 5132 -7370 5142 -7318
rect 5194 -7370 5204 -7318
rect 5132 -7374 5204 -7370
rect 5241 -7319 5311 -7316
rect 5241 -7371 5250 -7319
rect 5302 -7371 5311 -7319
rect 5241 -7374 5311 -7371
rect 5020 -7417 5080 -7374
rect 5016 -7423 5104 -7417
rect 5016 -7457 5043 -7423
rect 5077 -7457 5104 -7423
rect 5016 -7463 5104 -7457
rect 4922 -7550 4934 -7543
rect 4710 -7615 4756 -7577
rect 4710 -7649 4716 -7615
rect 4750 -7649 4756 -7615
rect 4710 -7687 4756 -7649
rect 4710 -7721 4716 -7687
rect 4750 -7721 4756 -7687
rect 4710 -7759 4756 -7721
rect 4710 -7793 4716 -7759
rect 4750 -7793 4756 -7759
rect 4710 -7831 4756 -7793
rect 4710 -7862 4716 -7831
rect 4492 -7904 4538 -7865
rect 4702 -7865 4716 -7862
rect 4750 -7862 4756 -7831
rect 4928 -7577 4934 -7550
rect 4968 -7550 4982 -7543
rect 5138 -7543 5198 -7374
rect 5247 -7417 5305 -7374
rect 5234 -7423 5322 -7417
rect 5234 -7457 5261 -7423
rect 5295 -7457 5322 -7423
rect 5234 -7463 5322 -7457
rect 5356 -7538 5416 -7256
rect 5576 -7366 5856 -7306
rect 5452 -7423 5540 -7417
rect 5452 -7457 5479 -7423
rect 5513 -7457 5540 -7423
rect 5452 -7463 5540 -7457
rect 4968 -7577 4974 -7550
rect 5138 -7556 5152 -7543
rect 4928 -7615 4974 -7577
rect 4928 -7649 4934 -7615
rect 4968 -7649 4974 -7615
rect 4928 -7687 4974 -7649
rect 4928 -7721 4934 -7687
rect 4968 -7721 4974 -7687
rect 4928 -7759 4974 -7721
rect 4928 -7793 4934 -7759
rect 4968 -7793 4974 -7759
rect 4928 -7831 4974 -7793
rect 4750 -7865 4762 -7862
rect 3926 -7951 4014 -7945
rect 3926 -7985 3953 -7951
rect 3987 -7985 4014 -7951
rect 3926 -7991 3940 -7985
rect 3942 -7991 4014 -7985
rect 4144 -7951 4232 -7945
rect 4144 -7985 4171 -7951
rect 4205 -7985 4232 -7951
rect 4144 -7991 4232 -7985
rect 4362 -7951 4450 -7945
rect 4362 -7985 4389 -7951
rect 4423 -7985 4450 -7951
rect 4362 -7991 4450 -7985
rect 4580 -7951 4668 -7945
rect 4580 -7985 4607 -7951
rect 4641 -7985 4668 -7951
rect 4580 -7991 4592 -7985
rect 4596 -7991 4668 -7985
rect 3942 -8034 4002 -7991
rect 4596 -8034 4656 -7991
rect 4702 -8034 4762 -7865
rect 4928 -7865 4934 -7831
rect 4968 -7865 4974 -7831
rect 4928 -7904 4974 -7865
rect 5146 -7577 5152 -7556
rect 5186 -7556 5198 -7543
rect 5364 -7543 5410 -7538
rect 5576 -7540 5636 -7366
rect 5682 -7417 5742 -7366
rect 5670 -7423 5758 -7417
rect 5670 -7457 5697 -7423
rect 5731 -7457 5758 -7423
rect 5670 -7463 5758 -7457
rect 5186 -7577 5192 -7556
rect 5146 -7615 5192 -7577
rect 5146 -7649 5152 -7615
rect 5186 -7649 5192 -7615
rect 5146 -7687 5192 -7649
rect 5146 -7721 5152 -7687
rect 5186 -7721 5192 -7687
rect 5146 -7759 5192 -7721
rect 5146 -7793 5152 -7759
rect 5186 -7793 5192 -7759
rect 5146 -7831 5192 -7793
rect 5146 -7865 5152 -7831
rect 5186 -7865 5192 -7831
rect 5146 -7904 5192 -7865
rect 5364 -7577 5370 -7543
rect 5404 -7577 5410 -7543
rect 5364 -7615 5410 -7577
rect 5364 -7649 5370 -7615
rect 5404 -7649 5410 -7615
rect 5364 -7687 5410 -7649
rect 5364 -7721 5370 -7687
rect 5404 -7721 5410 -7687
rect 5364 -7759 5410 -7721
rect 5364 -7793 5370 -7759
rect 5404 -7793 5410 -7759
rect 5364 -7831 5410 -7793
rect 5364 -7865 5370 -7831
rect 5404 -7865 5410 -7831
rect 5582 -7543 5628 -7540
rect 5582 -7577 5588 -7543
rect 5622 -7577 5628 -7543
rect 5796 -7543 5856 -7366
rect 5796 -7544 5806 -7543
rect 5582 -7615 5628 -7577
rect 5582 -7649 5588 -7615
rect 5622 -7649 5628 -7615
rect 5582 -7687 5628 -7649
rect 5582 -7721 5588 -7687
rect 5622 -7721 5628 -7687
rect 5582 -7759 5628 -7721
rect 5582 -7793 5588 -7759
rect 5622 -7793 5628 -7759
rect 5582 -7831 5628 -7793
rect 5582 -7858 5588 -7831
rect 5364 -7904 5410 -7865
rect 5576 -7865 5588 -7858
rect 5622 -7858 5628 -7831
rect 5800 -7577 5806 -7544
rect 5840 -7544 5856 -7543
rect 5840 -7577 5846 -7544
rect 5800 -7615 5846 -7577
rect 5800 -7649 5806 -7615
rect 5840 -7649 5846 -7615
rect 5800 -7687 5846 -7649
rect 5800 -7721 5806 -7687
rect 5840 -7721 5846 -7687
rect 5800 -7759 5846 -7721
rect 5800 -7793 5806 -7759
rect 5840 -7793 5846 -7759
rect 5800 -7831 5846 -7793
rect 5622 -7865 5636 -7858
rect 4798 -7951 4886 -7945
rect 4798 -7985 4825 -7951
rect 4859 -7985 4886 -7951
rect 4798 -7991 4872 -7985
rect 4874 -7991 4886 -7985
rect 5016 -7951 5104 -7945
rect 5016 -7985 5043 -7951
rect 5077 -7985 5104 -7951
rect 5016 -7991 5104 -7985
rect 5234 -7951 5322 -7945
rect 5234 -7985 5261 -7951
rect 5295 -7985 5322 -7951
rect 5234 -7991 5322 -7985
rect 5452 -7951 5540 -7945
rect 5452 -7985 5479 -7951
rect 5513 -7985 5540 -7951
rect 5452 -7991 5540 -7985
rect 4812 -8034 4872 -7991
rect 5464 -8034 5524 -7991
rect 5576 -8034 5636 -7865
rect 5800 -7865 5806 -7831
rect 5840 -7865 5846 -7831
rect 5800 -7904 5846 -7865
rect 5670 -7951 5758 -7945
rect 5670 -7985 5697 -7951
rect 5731 -7985 5758 -7951
rect 5670 -7991 5758 -7985
rect 6048 -8034 6108 -4562
rect 6802 -5608 6862 -3486
rect 6796 -5612 6868 -5608
rect 6796 -5664 6806 -5612
rect 6858 -5664 6868 -5612
rect 6796 -5668 6868 -5664
rect 6916 -5712 6976 -3360
rect 7312 -3404 7372 -3024
rect 9526 -3114 9590 -2744
rect 10032 -2752 10092 -2480
rect 10546 -2570 10610 -2396
rect 10540 -2574 10612 -2570
rect 10540 -2626 10550 -2574
rect 10602 -2626 10612 -2574
rect 10540 -2630 10612 -2626
rect 11074 -2752 11134 -2480
rect 10032 -2812 11134 -2752
rect 9520 -3120 9596 -3114
rect 9520 -3172 9532 -3120
rect 9584 -3172 9596 -3120
rect 9520 -3178 9596 -3172
rect 10032 -3216 10092 -2812
rect 9494 -3276 10092 -3216
rect 7306 -3408 7378 -3404
rect 7306 -3460 7316 -3408
rect 7368 -3460 7378 -3408
rect 7306 -3464 7378 -3460
rect 8472 -3408 8544 -3404
rect 8472 -3460 8482 -3408
rect 8534 -3460 8544 -3408
rect 8472 -3464 8544 -3460
rect 7038 -4454 7110 -4450
rect 7038 -4506 7048 -4454
rect 7100 -4506 7110 -4454
rect 7038 -4510 7110 -4506
rect 6910 -5716 6982 -5712
rect 6910 -5768 6920 -5716
rect 6972 -5768 6982 -5716
rect 6910 -5772 6982 -5768
rect 3826 -8038 3898 -8034
rect 3826 -8090 3836 -8038
rect 3888 -8090 3898 -8038
rect 3826 -8094 3898 -8090
rect 3936 -8038 4008 -8034
rect 3936 -8090 3946 -8038
rect 3998 -8090 4008 -8038
rect 3936 -8094 4008 -8090
rect 4590 -8038 4662 -8034
rect 4590 -8090 4600 -8038
rect 4652 -8090 4662 -8038
rect 4590 -8094 4662 -8090
rect 4696 -8038 4768 -8034
rect 4696 -8090 4706 -8038
rect 4758 -8090 4768 -8038
rect 4696 -8094 4768 -8090
rect 4806 -8038 4878 -8034
rect 4806 -8090 4816 -8038
rect 4868 -8090 4878 -8038
rect 4806 -8094 4878 -8090
rect 5458 -8038 5530 -8034
rect 5458 -8090 5468 -8038
rect 5520 -8090 5530 -8038
rect 5458 -8094 5530 -8090
rect 5570 -8038 5642 -8034
rect 5570 -8090 5580 -8038
rect 5632 -8090 5642 -8038
rect 5570 -8094 5642 -8090
rect 6042 -8038 6114 -8034
rect 6042 -8090 6052 -8038
rect 6104 -8090 6114 -8038
rect 6042 -8094 6114 -8090
rect 7044 -8122 7104 -4510
rect 7174 -4552 7246 -4548
rect 7174 -4604 7184 -4552
rect 7236 -4604 7246 -4552
rect 7174 -4608 7246 -4604
rect 7038 -8126 7110 -8122
rect 7038 -8178 7048 -8126
rect 7100 -8178 7110 -8126
rect 7038 -8182 7110 -8178
rect 7180 -8252 7240 -4608
rect 7312 -7072 7372 -3464
rect 8478 -3644 8538 -3464
rect 9494 -3664 9554 -3276
rect 11564 -3304 11624 -2372
rect 14618 -2376 14678 -2374
rect 12580 -2388 12640 -2386
rect 12580 -2566 12644 -2388
rect 12040 -2578 12100 -2568
rect 12040 -2630 12044 -2578
rect 12096 -2630 12100 -2578
rect 11558 -3308 11630 -3304
rect 11558 -3360 11568 -3308
rect 11620 -3360 11630 -3308
rect 11558 -3364 11630 -3360
rect 10508 -3408 10580 -3404
rect 10508 -3460 10518 -3408
rect 10570 -3460 10580 -3408
rect 10508 -3464 10580 -3460
rect 10514 -3642 10574 -3464
rect 12040 -3562 12100 -2630
rect 12548 -2570 12644 -2566
rect 12548 -2575 12646 -2570
rect 12548 -2627 12568 -2575
rect 12620 -2627 12646 -2575
rect 12548 -2630 12646 -2627
rect 13034 -2574 13106 -2570
rect 13034 -2626 13044 -2574
rect 13096 -2626 13106 -2574
rect 13034 -2630 13106 -2626
rect 7460 -4352 7520 -4158
rect 7974 -4352 8034 -4256
rect 8476 -4352 8536 -4170
rect 7460 -4412 8536 -4352
rect 8476 -4662 8548 -4658
rect 8476 -4714 8486 -4662
rect 8538 -4714 8548 -4662
rect 8476 -4718 8548 -4714
rect 8482 -4900 8542 -4718
rect 8966 -4816 9026 -4248
rect 9496 -4352 9556 -4170
rect 9490 -4356 9562 -4352
rect 9490 -4408 9500 -4356
rect 9552 -4408 9562 -4356
rect 9490 -4412 9562 -4408
rect 9496 -4548 9556 -4412
rect 9490 -4552 9562 -4548
rect 9490 -4604 9500 -4552
rect 9552 -4604 9562 -4552
rect 9490 -4608 9562 -4604
rect 10004 -4821 10064 -4247
rect 10510 -4550 10582 -4546
rect 10510 -4602 10520 -4550
rect 10572 -4602 10582 -4550
rect 10510 -4606 10582 -4602
rect 10516 -4658 10576 -4606
rect 10510 -4662 10582 -4658
rect 10510 -4714 10520 -4662
rect 10572 -4714 10582 -4662
rect 10510 -4718 10582 -4714
rect 10516 -4896 10576 -4718
rect 11010 -4821 11070 -4247
rect 11532 -4352 11592 -4166
rect 12042 -4348 12102 -4252
rect 12548 -4348 12608 -2630
rect 13040 -3558 13100 -2630
rect 13598 -2818 13662 -2388
rect 14618 -2562 14682 -2376
rect 16654 -2380 16714 -2378
rect 14084 -2572 14144 -2562
rect 14084 -2624 14088 -2572
rect 14140 -2624 14144 -2572
rect 13592 -2824 13668 -2818
rect 13592 -2876 13604 -2824
rect 13656 -2876 13668 -2824
rect 13592 -2882 13668 -2876
rect 13598 -3108 13662 -2882
rect 13598 -3160 13604 -3108
rect 13656 -3160 13662 -3108
rect 13598 -3172 13662 -3160
rect 14084 -3572 14144 -2624
rect 14586 -2572 14682 -2562
rect 15100 -2572 15160 -2562
rect 14586 -2574 14684 -2572
rect 14586 -2626 14606 -2574
rect 14658 -2626 14684 -2574
rect 14586 -2632 14684 -2626
rect 15100 -2624 15104 -2572
rect 15156 -2624 15160 -2572
rect 13062 -4348 13122 -4256
rect 13568 -4348 13628 -4170
rect 14072 -4348 14132 -4254
rect 14586 -4348 14646 -2632
rect 15100 -3562 15160 -2624
rect 15634 -2818 15698 -2384
rect 16128 -2572 16188 -2562
rect 16654 -2568 16718 -2380
rect 18690 -2392 18750 -2390
rect 16128 -2624 16132 -2572
rect 16184 -2624 16188 -2572
rect 15628 -2824 15704 -2818
rect 15628 -2876 15640 -2824
rect 15692 -2876 15704 -2824
rect 15628 -2882 15704 -2876
rect 16128 -3562 16188 -2624
rect 16622 -2572 16718 -2568
rect 16622 -2577 16720 -2572
rect 16622 -2629 16642 -2577
rect 16694 -2629 16720 -2577
rect 16622 -2632 16720 -2629
rect 17150 -2582 17210 -2572
rect 15094 -4348 15154 -4256
rect 15602 -4348 15662 -4168
rect 16116 -4348 16176 -4256
rect 16622 -4348 16682 -2632
rect 17150 -2634 17154 -2582
rect 17206 -2634 17210 -2582
rect 17150 -3566 17210 -2634
rect 17638 -2578 17698 -2568
rect 17638 -2630 17642 -2578
rect 17694 -2630 17698 -2578
rect 17142 -4348 17202 -4255
rect 17638 -4348 17698 -2630
rect 18150 -2582 18210 -2572
rect 18690 -2574 18754 -2392
rect 18150 -2634 18154 -2582
rect 18206 -2634 18210 -2582
rect 18684 -2578 18756 -2574
rect 18684 -2630 18694 -2578
rect 18746 -2630 18756 -2578
rect 18684 -2634 18756 -2630
rect 18150 -3572 18210 -2634
rect 19706 -2680 19770 -2386
rect 20724 -2392 20784 -2390
rect 20724 -2574 20788 -2392
rect 20718 -2578 20790 -2574
rect 20718 -2630 20728 -2578
rect 20780 -2630 20790 -2578
rect 20718 -2634 20790 -2630
rect 19700 -2686 19776 -2680
rect 19700 -2738 19712 -2686
rect 19764 -2738 19776 -2686
rect 19700 -2744 19776 -2738
rect 21742 -2818 21806 -2390
rect 21736 -2824 21812 -2818
rect 21736 -2876 21748 -2824
rect 21800 -2876 21812 -2824
rect 21736 -2882 21812 -2876
rect 21714 -3102 21774 -3092
rect 21714 -3154 21718 -3102
rect 21770 -3154 21774 -3102
rect 21714 -3400 21774 -3154
rect 22884 -3108 22944 -354
rect 22884 -3160 22888 -3108
rect 22940 -3160 22944 -3108
rect 22884 -3170 22944 -3160
rect 24716 -359 24828 -321
rect 24716 -393 24755 -359
rect 24789 -393 24828 -359
rect 24716 -431 24828 -393
rect 24716 -465 24755 -431
rect 24789 -465 24828 -431
rect 24716 -503 24828 -465
rect 24716 -537 24755 -503
rect 24789 -537 24828 -503
rect 24716 -575 24828 -537
rect 24716 -609 24755 -575
rect 24789 -609 24828 -575
rect 24716 -647 24828 -609
rect 24716 -681 24755 -647
rect 24789 -681 24828 -647
rect 24716 -719 24828 -681
rect 24716 -753 24755 -719
rect 24789 -753 24828 -719
rect 24716 -791 24828 -753
rect 24716 -825 24755 -791
rect 24789 -825 24828 -791
rect 24716 -863 24828 -825
rect 24716 -897 24755 -863
rect 24789 -897 24828 -863
rect 24716 -935 24828 -897
rect 24716 -969 24755 -935
rect 24789 -969 24828 -935
rect 24716 -1007 24828 -969
rect 24716 -1041 24755 -1007
rect 24789 -1041 24828 -1007
rect 24716 -1079 24828 -1041
rect 24716 -1113 24755 -1079
rect 24789 -1113 24828 -1079
rect 24716 -1151 24828 -1113
rect 24716 -1185 24755 -1151
rect 24789 -1185 24828 -1151
rect 24716 -1223 24828 -1185
rect 24716 -1257 24755 -1223
rect 24789 -1257 24828 -1223
rect 24716 -1295 24828 -1257
rect 24716 -1329 24755 -1295
rect 24789 -1329 24828 -1295
rect 24716 -1367 24828 -1329
rect 24716 -1401 24755 -1367
rect 24789 -1401 24828 -1367
rect 24716 -1439 24828 -1401
rect 24716 -1473 24755 -1439
rect 24789 -1473 24828 -1439
rect 24716 -1511 24828 -1473
rect 24716 -1545 24755 -1511
rect 24789 -1545 24828 -1511
rect 24716 -1583 24828 -1545
rect 24716 -1617 24755 -1583
rect 24789 -1617 24828 -1583
rect 24716 -1655 24828 -1617
rect 24716 -1689 24755 -1655
rect 24789 -1689 24828 -1655
rect 24716 -1727 24828 -1689
rect 24716 -1761 24755 -1727
rect 24789 -1761 24828 -1727
rect 24716 -1799 24828 -1761
rect 24716 -1833 24755 -1799
rect 24789 -1833 24828 -1799
rect 24716 -1871 24828 -1833
rect 24716 -1905 24755 -1871
rect 24789 -1905 24828 -1871
rect 24716 -1943 24828 -1905
rect 24716 -1977 24755 -1943
rect 24789 -1977 24828 -1943
rect 24716 -2015 24828 -1977
rect 24716 -2049 24755 -2015
rect 24789 -2049 24828 -2015
rect 24716 -2087 24828 -2049
rect 24716 -2121 24755 -2087
rect 24789 -2121 24828 -2087
rect 24716 -2159 24828 -2121
rect 24716 -2193 24755 -2159
rect 24789 -2193 24828 -2159
rect 24716 -2231 24828 -2193
rect 24716 -2265 24755 -2231
rect 24789 -2265 24828 -2231
rect 24716 -2303 24828 -2265
rect 24716 -2337 24755 -2303
rect 24789 -2337 24828 -2303
rect 24716 -2375 24828 -2337
rect 24716 -2409 24755 -2375
rect 24789 -2409 24828 -2375
rect 24716 -2447 24828 -2409
rect 24716 -2481 24755 -2447
rect 24789 -2481 24828 -2447
rect 24716 -2519 24828 -2481
rect 24716 -2553 24755 -2519
rect 24789 -2553 24828 -2519
rect 24716 -2591 24828 -2553
rect 24716 -2625 24755 -2591
rect 24789 -2625 24828 -2591
rect 24716 -2663 24828 -2625
rect 24716 -2697 24755 -2663
rect 24789 -2697 24828 -2663
rect 24716 -2735 24828 -2697
rect 24716 -2769 24755 -2735
rect 24789 -2769 24828 -2735
rect 24716 -2807 24828 -2769
rect 24716 -2841 24755 -2807
rect 24789 -2841 24828 -2807
rect 24716 -2879 24828 -2841
rect 24716 -2913 24755 -2879
rect 24789 -2913 24828 -2879
rect 24716 -2951 24828 -2913
rect 24716 -2985 24755 -2951
rect 24789 -2985 24828 -2951
rect 24716 -3023 24828 -2985
rect 24716 -3057 24755 -3023
rect 24789 -3057 24828 -3023
rect 24716 -3095 24828 -3057
rect 24716 -3129 24755 -3095
rect 24789 -3129 24828 -3095
rect 24716 -3167 24828 -3129
rect 24716 -3201 24755 -3167
rect 24789 -3201 24828 -3167
rect 24716 -3239 24828 -3201
rect 24716 -3273 24755 -3239
rect 24789 -3273 24828 -3239
rect 24716 -3311 24828 -3273
rect 24716 -3345 24755 -3311
rect 24789 -3345 24828 -3311
rect 24716 -3383 24828 -3345
rect 18654 -3408 18726 -3404
rect 18654 -3460 18664 -3408
rect 18716 -3460 18726 -3408
rect 18654 -3464 18726 -3460
rect 20688 -3408 20760 -3404
rect 20688 -3460 20698 -3408
rect 20750 -3460 20760 -3408
rect 20688 -3464 20760 -3460
rect 21714 -3460 22790 -3400
rect 18660 -3646 18720 -3464
rect 20694 -3642 20754 -3464
rect 21714 -3654 21774 -3460
rect 22228 -3556 22288 -3460
rect 22730 -3642 22790 -3460
rect 23132 -3408 23204 -3404
rect 23132 -3460 23142 -3408
rect 23194 -3460 23204 -3408
rect 23132 -3464 23204 -3460
rect 24716 -3417 24755 -3383
rect 24789 -3417 24828 -3383
rect 24716 -3455 24828 -3417
rect 18154 -4348 18214 -4258
rect 11526 -4356 11598 -4352
rect 11526 -4408 11536 -4356
rect 11588 -4408 11598 -4356
rect 12042 -4408 18214 -4348
rect 11526 -4412 11598 -4408
rect 12548 -4508 12608 -4408
rect 17638 -4508 17698 -4408
rect 12548 -4568 17698 -4508
rect 12548 -4918 12608 -4568
rect 13566 -4664 13638 -4660
rect 13566 -4716 13576 -4664
rect 13628 -4716 13638 -4664
rect 13566 -4720 13638 -4716
rect 14076 -4706 15134 -4646
rect 13572 -4902 13632 -4720
rect 14076 -4818 14136 -4706
rect 15076 -4744 15134 -4706
rect 15600 -4664 15672 -4660
rect 15600 -4716 15610 -4664
rect 15662 -4716 15672 -4664
rect 15600 -4720 15672 -4716
rect 15076 -4818 15136 -4744
rect 15606 -4904 15666 -4720
rect 17638 -4894 17698 -4568
rect 18656 -4664 18728 -4660
rect 18656 -4716 18666 -4664
rect 18718 -4716 18728 -4664
rect 18656 -4720 18728 -4716
rect 18662 -4902 18722 -4720
rect 19162 -4821 19222 -4247
rect 19676 -4352 19736 -4170
rect 19670 -4356 19742 -4352
rect 19670 -4408 19680 -4356
rect 19732 -4408 19742 -4356
rect 19670 -4412 19742 -4408
rect 20186 -4821 20246 -4247
rect 20690 -4664 20762 -4660
rect 20690 -4716 20700 -4664
rect 20752 -4716 20762 -4664
rect 20690 -4720 20762 -4716
rect 20696 -4898 20756 -4720
rect 21192 -4815 21252 -4241
rect 21712 -4352 21772 -4166
rect 21706 -4356 21778 -4352
rect 21706 -4408 21716 -4356
rect 21768 -4408 21778 -4356
rect 21706 -4412 21778 -4408
rect 22972 -4550 23044 -4546
rect 22972 -4602 22982 -4550
rect 23034 -4602 23044 -4550
rect 22972 -4606 23044 -4602
rect 21714 -4714 22790 -4654
rect 21714 -4908 21774 -4714
rect 22228 -4810 22288 -4714
rect 22730 -4896 22790 -4714
rect 7464 -5608 7524 -5414
rect 7978 -5608 8038 -5512
rect 8480 -5608 8540 -5426
rect 7464 -5668 8540 -5608
rect 7462 -5970 8538 -5910
rect 7462 -6164 7522 -5970
rect 7976 -6066 8036 -5970
rect 8478 -6152 8538 -5970
rect 8960 -6076 9020 -5502
rect 9498 -5716 9558 -5424
rect 9498 -5768 9502 -5716
rect 9554 -5768 9558 -5716
rect 9498 -5778 9558 -5768
rect 9492 -5920 9564 -5916
rect 9492 -5972 9502 -5920
rect 9554 -5972 9564 -5920
rect 9492 -5976 9564 -5972
rect 9498 -6154 9558 -5976
rect 9998 -6077 10058 -5502
rect 11004 -6077 11064 -5502
rect 11534 -5712 11594 -5420
rect 12054 -5604 12114 -5511
rect 12550 -5604 12610 -5420
rect 13066 -5604 13126 -5514
rect 12054 -5664 13126 -5604
rect 13562 -5612 13634 -5608
rect 13562 -5664 13572 -5612
rect 13624 -5664 13634 -5612
rect 11528 -5716 11600 -5712
rect 11528 -5768 11538 -5716
rect 11590 -5768 11600 -5716
rect 11528 -5772 11600 -5768
rect 11526 -5818 11598 -5814
rect 11526 -5870 11536 -5818
rect 11588 -5870 11598 -5818
rect 11526 -5874 11598 -5870
rect 11532 -5916 11592 -5874
rect 11526 -5920 11598 -5916
rect 11526 -5972 11536 -5920
rect 11588 -5972 11598 -5920
rect 11526 -5976 11598 -5972
rect 11532 -6158 11592 -5976
rect 12550 -6168 12610 -5664
rect 13562 -5668 13634 -5664
rect 13568 -6154 13628 -5668
rect 14070 -6082 14130 -5508
rect 14588 -5608 14648 -5426
rect 14582 -5612 14654 -5608
rect 14582 -5664 14592 -5612
rect 14644 -5664 14654 -5612
rect 14582 -5668 14654 -5664
rect 14582 -5918 14654 -5914
rect 14582 -5970 14592 -5918
rect 14644 -5970 14654 -5918
rect 14582 -5974 14654 -5970
rect 14588 -6152 14648 -5974
rect 15100 -6070 15160 -5496
rect 15606 -5914 15666 -5422
rect 15600 -5918 15672 -5914
rect 15600 -5970 15610 -5918
rect 15662 -5970 15672 -5918
rect 15600 -5974 15672 -5970
rect 16112 -6070 16172 -5496
rect 16624 -5608 16684 -5422
rect 17142 -5606 17202 -5513
rect 17638 -5606 17698 -5422
rect 18154 -5606 18214 -5516
rect 16618 -5612 16690 -5608
rect 16618 -5664 16628 -5612
rect 16680 -5664 16690 -5612
rect 16618 -5668 16690 -5664
rect 17142 -5666 18214 -5606
rect 16616 -5918 16688 -5914
rect 16616 -5970 16626 -5918
rect 16678 -5970 16688 -5918
rect 16616 -5974 16688 -5970
rect 16622 -6156 16682 -5974
rect 17638 -6160 17698 -5666
rect 18652 -5716 18724 -5712
rect 18652 -5768 18662 -5716
rect 18714 -5768 18724 -5716
rect 18652 -5772 18724 -5768
rect 18658 -6162 18718 -5772
rect 19156 -6077 19216 -5502
rect 19520 -5598 19592 -5594
rect 19520 -5650 19530 -5598
rect 19582 -5650 19592 -5598
rect 19520 -5654 19592 -5650
rect 19526 -5914 19586 -5654
rect 19674 -5704 19734 -5414
rect 19668 -5708 19740 -5704
rect 19668 -5760 19678 -5708
rect 19730 -5760 19740 -5708
rect 19668 -5764 19740 -5760
rect 19520 -5918 19592 -5914
rect 19520 -5970 19530 -5918
rect 19582 -5970 19592 -5918
rect 19520 -5974 19592 -5970
rect 19672 -5916 19744 -5912
rect 19672 -5968 19682 -5916
rect 19734 -5968 19744 -5916
rect 19672 -5972 19744 -5968
rect 19678 -6150 19738 -5972
rect 20180 -6077 20240 -5502
rect 20694 -5814 20754 -5422
rect 20688 -5818 20760 -5814
rect 20688 -5870 20698 -5818
rect 20750 -5870 20760 -5818
rect 20688 -5874 20760 -5870
rect 21186 -6071 21246 -5496
rect 21714 -5704 21774 -5410
rect 21708 -5708 21780 -5704
rect 21708 -5760 21718 -5708
rect 21770 -5760 21780 -5708
rect 21708 -5764 21780 -5760
rect 22840 -5708 22912 -5704
rect 22840 -5760 22850 -5708
rect 22902 -5760 22912 -5708
rect 22840 -5764 22912 -5760
rect 21706 -5916 21778 -5912
rect 21706 -5968 21716 -5916
rect 21768 -5968 21778 -5916
rect 21706 -5972 21778 -5968
rect 21712 -6154 21772 -5972
rect 8480 -6864 8540 -6678
rect 8474 -6868 8546 -6864
rect 8474 -6920 8484 -6868
rect 8536 -6920 8546 -6868
rect 8474 -6924 8546 -6920
rect 7306 -7076 7378 -7072
rect 7306 -7128 7316 -7076
rect 7368 -7128 7378 -7076
rect 7306 -7132 7378 -7128
rect 7462 -7230 8538 -7170
rect 7462 -7424 7522 -7230
rect 7976 -7326 8036 -7230
rect 8478 -7412 8538 -7230
rect 8972 -7326 9032 -6752
rect 9488 -7178 9560 -7174
rect 9488 -7230 9498 -7178
rect 9550 -7230 9560 -7178
rect 9488 -7234 9560 -7230
rect 9494 -7412 9554 -7234
rect 10010 -7326 10070 -6752
rect 10516 -6864 10576 -6682
rect 10510 -6868 10582 -6864
rect 10510 -6920 10520 -6868
rect 10572 -6920 10582 -6868
rect 10510 -6924 10582 -6920
rect 10516 -6972 10576 -6924
rect 10510 -6976 10582 -6972
rect 10510 -7028 10520 -6976
rect 10572 -7028 10582 -6976
rect 10510 -7032 10582 -7028
rect 11016 -7022 11076 -6752
rect 12052 -6856 12112 -6763
rect 12548 -6856 12608 -6672
rect 13064 -6856 13124 -6766
rect 12052 -6916 13124 -6856
rect 13570 -6862 13630 -6676
rect 13564 -6866 13636 -6862
rect 11016 -7082 11792 -7022
rect 11016 -7326 11076 -7082
rect 11732 -7168 11792 -7082
rect 11726 -7172 11798 -7168
rect 11522 -7178 11594 -7174
rect 11522 -7230 11532 -7178
rect 11584 -7230 11594 -7178
rect 11726 -7224 11736 -7172
rect 11788 -7224 11798 -7172
rect 11726 -7228 11798 -7224
rect 11522 -7234 11594 -7230
rect 11528 -7416 11588 -7234
rect 12548 -7444 12608 -6916
rect 13564 -6918 13574 -6866
rect 13626 -6918 13636 -6866
rect 13564 -6922 13636 -6918
rect 14080 -6994 14140 -6764
rect 15096 -6994 15156 -6756
rect 15606 -6862 15666 -6680
rect 15600 -6866 15672 -6862
rect 15600 -6918 15610 -6866
rect 15662 -6918 15672 -6866
rect 15600 -6922 15672 -6918
rect 16110 -6994 16170 -6760
rect 17140 -6858 17200 -6765
rect 17636 -6858 17696 -6674
rect 18152 -6858 18212 -6768
rect 17140 -6918 18212 -6858
rect 18660 -6860 18720 -6674
rect 18654 -6864 18726 -6860
rect 18654 -6916 18664 -6864
rect 18716 -6916 18726 -6864
rect 14080 -7054 16894 -6994
rect 13566 -7168 13626 -7162
rect 14080 -7168 14140 -7054
rect 13566 -7172 14140 -7168
rect 13566 -7224 13570 -7172
rect 13622 -7224 14140 -7172
rect 13566 -7228 14140 -7224
rect 14580 -7176 14652 -7172
rect 14580 -7228 14590 -7176
rect 14642 -7228 14652 -7176
rect 13566 -7234 13626 -7228
rect 14580 -7232 14652 -7228
rect 16614 -7176 16686 -7172
rect 16834 -7176 16894 -7054
rect 16614 -7228 16624 -7176
rect 16676 -7228 16686 -7176
rect 16614 -7232 16686 -7228
rect 16828 -7180 16900 -7176
rect 16828 -7232 16838 -7180
rect 16890 -7232 16900 -7180
rect 14586 -7410 14646 -7232
rect 16620 -7414 16680 -7232
rect 16828 -7236 16900 -7232
rect 17636 -7424 17696 -6918
rect 18654 -6920 18726 -6916
rect 19168 -7170 19228 -6752
rect 19168 -7180 19230 -7170
rect 19168 -7232 19174 -7180
rect 19226 -7232 19230 -7180
rect 19168 -7242 19230 -7232
rect 19676 -7178 19748 -7174
rect 19676 -7230 19686 -7178
rect 19738 -7230 19748 -7178
rect 19676 -7234 19748 -7230
rect 19168 -7326 19228 -7242
rect 19682 -7412 19742 -7234
rect 20192 -7326 20252 -6752
rect 20696 -6860 20756 -6678
rect 20690 -6864 20762 -6860
rect 20690 -6916 20700 -6864
rect 20752 -6916 20762 -6864
rect 20690 -6920 20762 -6916
rect 21198 -7320 21258 -6746
rect 21712 -6864 21772 -6670
rect 22226 -6864 22286 -6768
rect 22728 -6864 22788 -6682
rect 21712 -6924 22788 -6864
rect 22846 -6972 22906 -5764
rect 22978 -5912 23038 -4606
rect 22972 -5916 23044 -5912
rect 22972 -5968 22982 -5916
rect 23034 -5968 23044 -5916
rect 22972 -5972 23044 -5968
rect 22840 -6976 22912 -6972
rect 22840 -7028 22850 -6976
rect 22902 -7028 22912 -6976
rect 22840 -7032 22912 -7028
rect 21710 -7178 21782 -7174
rect 21710 -7230 21720 -7178
rect 21772 -7230 21782 -7178
rect 21710 -7234 21782 -7230
rect 21716 -7416 21776 -7234
rect 8476 -8122 8536 -7936
rect 8470 -8126 8542 -8122
rect 8470 -8178 8480 -8126
rect 8532 -8178 8542 -8126
rect 8470 -8182 8542 -8178
rect 8984 -8236 9044 -8024
rect 10008 -8236 10068 -8016
rect 10512 -8122 10572 -7940
rect 10506 -8126 10578 -8122
rect 10506 -8178 10516 -8126
rect 10568 -8178 10578 -8126
rect 10506 -8182 10578 -8178
rect 11014 -8236 11074 -8016
rect 7174 -8256 7246 -8252
rect 7174 -8308 7184 -8256
rect 7236 -8308 7246 -8256
rect 7174 -8312 7246 -8308
rect 8984 -8296 11074 -8236
rect 2104 -8396 2176 -8392
rect 2104 -8448 2114 -8396
rect 2166 -8448 2176 -8396
rect 2104 -8452 2176 -8448
rect 1954 -8498 2014 -8492
rect 7180 -8498 7240 -8312
rect 1954 -8502 7240 -8498
rect 1954 -8554 1958 -8502
rect 2010 -8554 7240 -8502
rect 1954 -8558 7240 -8554
rect 1954 -8564 2014 -8558
rect 1184 -8616 1244 -8610
rect 8984 -8616 9044 -8296
rect 11014 -8546 11074 -8296
rect 11534 -8392 11594 -7926
rect 12052 -8116 12112 -8021
rect 12548 -8116 12608 -7930
rect 13064 -8116 13124 -8024
rect 13570 -8116 13630 -7918
rect 14080 -8116 14140 -8024
rect 14586 -8116 14646 -7938
rect 15096 -8116 15156 -8024
rect 15604 -8116 15664 -7924
rect 16106 -8116 16166 -8024
rect 16622 -8116 16682 -7934
rect 17140 -8116 17200 -8023
rect 17636 -8116 17696 -7932
rect 18152 -8116 18212 -8026
rect 12052 -8176 18212 -8116
rect 18664 -8122 18724 -7936
rect 18658 -8126 18730 -8122
rect 18658 -8178 18668 -8126
rect 18720 -8178 18730 -8126
rect 18658 -8182 18730 -8178
rect 19172 -8234 19232 -8008
rect 20192 -8234 20252 -8016
rect 20700 -8122 20760 -7940
rect 20694 -8126 20766 -8122
rect 20694 -8178 20704 -8126
rect 20756 -8178 20766 -8126
rect 20694 -8182 20766 -8178
rect 21194 -8234 21254 -8016
rect 21714 -8118 21774 -7924
rect 22228 -8118 22288 -8022
rect 22730 -8118 22790 -7936
rect 21714 -8178 22790 -8118
rect 19172 -8294 21254 -8234
rect 11528 -8396 11600 -8392
rect 11528 -8448 11538 -8396
rect 11590 -8448 11600 -8396
rect 11528 -8452 11600 -8448
rect 19172 -8546 19232 -8294
rect 23138 -8392 23198 -3464
rect 24716 -3489 24755 -3455
rect 24789 -3489 24828 -3455
rect 24716 -3527 24828 -3489
rect 24716 -3561 24755 -3527
rect 24789 -3561 24828 -3527
rect 24716 -3599 24828 -3561
rect 24716 -3633 24755 -3599
rect 24789 -3633 24828 -3599
rect 24716 -3671 24828 -3633
rect 24716 -3705 24755 -3671
rect 24789 -3705 24828 -3671
rect 24716 -3743 24828 -3705
rect 24716 -3777 24755 -3743
rect 24789 -3777 24828 -3743
rect 24716 -3815 24828 -3777
rect 24716 -3849 24755 -3815
rect 24789 -3849 24828 -3815
rect 24716 -3887 24828 -3849
rect 24716 -3921 24755 -3887
rect 24789 -3921 24828 -3887
rect 24716 -3959 24828 -3921
rect 24716 -3993 24755 -3959
rect 24789 -3993 24828 -3959
rect 24716 -4031 24828 -3993
rect 24716 -4065 24755 -4031
rect 24789 -4065 24828 -4031
rect 24716 -4103 24828 -4065
rect 24716 -4137 24755 -4103
rect 24789 -4137 24828 -4103
rect 24716 -4175 24828 -4137
rect 24716 -4209 24755 -4175
rect 24789 -4209 24828 -4175
rect 24716 -4247 24828 -4209
rect 24716 -4281 24755 -4247
rect 24789 -4281 24828 -4247
rect 24716 -4319 24828 -4281
rect 24716 -4353 24755 -4319
rect 24789 -4353 24828 -4319
rect 24716 -4391 24828 -4353
rect 24716 -4425 24755 -4391
rect 24789 -4425 24828 -4391
rect 24716 -4463 24828 -4425
rect 24716 -4497 24755 -4463
rect 24789 -4497 24828 -4463
rect 24716 -4535 24828 -4497
rect 24716 -4569 24755 -4535
rect 24789 -4569 24828 -4535
rect 24716 -4607 24828 -4569
rect 24716 -4641 24755 -4607
rect 24789 -4641 24828 -4607
rect 24716 -4679 24828 -4641
rect 24716 -4713 24755 -4679
rect 24789 -4713 24828 -4679
rect 24716 -4751 24828 -4713
rect 24716 -4785 24755 -4751
rect 24789 -4785 24828 -4751
rect 24716 -4823 24828 -4785
rect 24716 -4857 24755 -4823
rect 24789 -4857 24828 -4823
rect 24716 -4895 24828 -4857
rect 24716 -4929 24755 -4895
rect 24789 -4929 24828 -4895
rect 24716 -4967 24828 -4929
rect 24716 -5001 24755 -4967
rect 24789 -5001 24828 -4967
rect 24716 -5039 24828 -5001
rect 24716 -5073 24755 -5039
rect 24789 -5073 24828 -5039
rect 24716 -5111 24828 -5073
rect 24716 -5145 24755 -5111
rect 24789 -5145 24828 -5111
rect 24716 -5183 24828 -5145
rect 24716 -5217 24755 -5183
rect 24789 -5217 24828 -5183
rect 24716 -5255 24828 -5217
rect 24716 -5289 24755 -5255
rect 24789 -5289 24828 -5255
rect 24716 -5327 24828 -5289
rect 24716 -5361 24755 -5327
rect 24789 -5361 24828 -5327
rect 24716 -5399 24828 -5361
rect 24716 -5433 24755 -5399
rect 24789 -5433 24828 -5399
rect 24716 -5471 24828 -5433
rect 24716 -5505 24755 -5471
rect 24789 -5505 24828 -5471
rect 24716 -5543 24828 -5505
rect 24716 -5577 24755 -5543
rect 24789 -5577 24828 -5543
rect 24716 -5615 24828 -5577
rect 24716 -5649 24755 -5615
rect 24789 -5649 24828 -5615
rect 24716 -5687 24828 -5649
rect 24716 -5721 24755 -5687
rect 24789 -5721 24828 -5687
rect 24716 -5759 24828 -5721
rect 24716 -5793 24755 -5759
rect 24789 -5793 24828 -5759
rect 24716 -5831 24828 -5793
rect 24716 -5865 24755 -5831
rect 24789 -5865 24828 -5831
rect 24716 -5903 24828 -5865
rect 24716 -5937 24755 -5903
rect 24789 -5937 24828 -5903
rect 24716 -5975 24828 -5937
rect 24716 -6009 24755 -5975
rect 24789 -6009 24828 -5975
rect 24716 -6047 24828 -6009
rect 24716 -6081 24755 -6047
rect 24789 -6081 24828 -6047
rect 24716 -6119 24828 -6081
rect 24716 -6153 24755 -6119
rect 24789 -6153 24828 -6119
rect 24716 -6191 24828 -6153
rect 24716 -6225 24755 -6191
rect 24789 -6225 24828 -6191
rect 24716 -6263 24828 -6225
rect 24716 -6297 24755 -6263
rect 24789 -6297 24828 -6263
rect 24716 -6335 24828 -6297
rect 24716 -6369 24755 -6335
rect 24789 -6369 24828 -6335
rect 24716 -6407 24828 -6369
rect 24716 -6441 24755 -6407
rect 24789 -6441 24828 -6407
rect 24716 -6479 24828 -6441
rect 24716 -6513 24755 -6479
rect 24789 -6513 24828 -6479
rect 24716 -6551 24828 -6513
rect 24716 -6585 24755 -6551
rect 24789 -6585 24828 -6551
rect 24716 -6623 24828 -6585
rect 24716 -6657 24755 -6623
rect 24789 -6657 24828 -6623
rect 24716 -6695 24828 -6657
rect 24716 -6729 24755 -6695
rect 24789 -6729 24828 -6695
rect 24716 -6767 24828 -6729
rect 24716 -6801 24755 -6767
rect 24789 -6801 24828 -6767
rect 24716 -6839 24828 -6801
rect 24716 -6873 24755 -6839
rect 24789 -6873 24828 -6839
rect 24716 -6911 24828 -6873
rect 24716 -6945 24755 -6911
rect 24789 -6945 24828 -6911
rect 24716 -6983 24828 -6945
rect 24716 -7017 24755 -6983
rect 24789 -7017 24828 -6983
rect 24716 -7055 24828 -7017
rect 24716 -7089 24755 -7055
rect 24789 -7089 24828 -7055
rect 24716 -7127 24828 -7089
rect 24716 -7161 24755 -7127
rect 24789 -7161 24828 -7127
rect 24716 -7199 24828 -7161
rect 24716 -7233 24755 -7199
rect 24789 -7233 24828 -7199
rect 24716 -7271 24828 -7233
rect 24716 -7305 24755 -7271
rect 24789 -7305 24828 -7271
rect 24716 -7343 24828 -7305
rect 24716 -7377 24755 -7343
rect 24789 -7377 24828 -7343
rect 24716 -7415 24828 -7377
rect 24716 -7449 24755 -7415
rect 24789 -7449 24828 -7415
rect 24716 -7487 24828 -7449
rect 24716 -7521 24755 -7487
rect 24789 -7521 24828 -7487
rect 24716 -7559 24828 -7521
rect 24716 -7593 24755 -7559
rect 24789 -7593 24828 -7559
rect 24716 -7631 24828 -7593
rect 24716 -7665 24755 -7631
rect 24789 -7665 24828 -7631
rect 24716 -7703 24828 -7665
rect 24716 -7737 24755 -7703
rect 24789 -7737 24828 -7703
rect 24716 -7775 24828 -7737
rect 24716 -7809 24755 -7775
rect 24789 -7809 24828 -7775
rect 24716 -7847 24828 -7809
rect 24716 -7881 24755 -7847
rect 24789 -7881 24828 -7847
rect 24716 -7919 24828 -7881
rect 24716 -7953 24755 -7919
rect 24789 -7953 24828 -7919
rect 24716 -7991 24828 -7953
rect 24716 -8025 24755 -7991
rect 24789 -8025 24828 -7991
rect 24716 -8063 24828 -8025
rect 24716 -8097 24755 -8063
rect 24789 -8097 24828 -8063
rect 24716 -8135 24828 -8097
rect 24716 -8169 24755 -8135
rect 24789 -8169 24828 -8135
rect 24716 -8207 24828 -8169
rect 24716 -8241 24755 -8207
rect 24789 -8241 24828 -8207
rect 23132 -8396 23204 -8392
rect 23132 -8448 23142 -8396
rect 23194 -8448 23204 -8396
rect 23132 -8452 23204 -8448
rect 11014 -8606 19232 -8546
rect 1184 -8620 9044 -8616
rect 1184 -8672 1188 -8620
rect 1240 -8672 9044 -8620
rect 1184 -8676 9044 -8672
rect 1184 -8682 1244 -8676
rect 24716 -8776 24828 -8241
rect 372 -8815 24828 -8776
rect 372 -8849 487 -8815
rect 521 -8849 559 -8815
rect 593 -8849 631 -8815
rect 665 -8849 703 -8815
rect 737 -8849 775 -8815
rect 809 -8849 847 -8815
rect 881 -8849 919 -8815
rect 953 -8849 991 -8815
rect 1025 -8849 1063 -8815
rect 1097 -8849 1135 -8815
rect 1169 -8849 1207 -8815
rect 1241 -8849 1279 -8815
rect 1313 -8849 1351 -8815
rect 1385 -8849 1423 -8815
rect 1457 -8849 1495 -8815
rect 1529 -8849 1567 -8815
rect 1601 -8849 1639 -8815
rect 1673 -8849 1711 -8815
rect 1745 -8849 1783 -8815
rect 1817 -8849 1855 -8815
rect 1889 -8849 1927 -8815
rect 1961 -8849 1999 -8815
rect 2033 -8849 2071 -8815
rect 2105 -8849 2143 -8815
rect 2177 -8849 2215 -8815
rect 2249 -8849 2287 -8815
rect 2321 -8849 2359 -8815
rect 2393 -8849 2431 -8815
rect 2465 -8849 2503 -8815
rect 2537 -8849 2575 -8815
rect 2609 -8849 2647 -8815
rect 2681 -8849 2719 -8815
rect 2753 -8849 2791 -8815
rect 2825 -8849 2863 -8815
rect 2897 -8849 2935 -8815
rect 2969 -8849 3007 -8815
rect 3041 -8849 3079 -8815
rect 3113 -8849 3151 -8815
rect 3185 -8849 3223 -8815
rect 3257 -8849 3295 -8815
rect 3329 -8849 3367 -8815
rect 3401 -8849 3439 -8815
rect 3473 -8849 3511 -8815
rect 3545 -8849 3583 -8815
rect 3617 -8849 3655 -8815
rect 3689 -8849 3727 -8815
rect 3761 -8849 3799 -8815
rect 3833 -8849 3871 -8815
rect 3905 -8849 3943 -8815
rect 3977 -8849 4015 -8815
rect 4049 -8849 4087 -8815
rect 4121 -8849 4159 -8815
rect 4193 -8849 4231 -8815
rect 4265 -8849 4303 -8815
rect 4337 -8849 4375 -8815
rect 4409 -8849 4447 -8815
rect 4481 -8849 4519 -8815
rect 4553 -8849 4591 -8815
rect 4625 -8849 4663 -8815
rect 4697 -8849 4735 -8815
rect 4769 -8849 4807 -8815
rect 4841 -8849 4879 -8815
rect 4913 -8849 4951 -8815
rect 4985 -8849 5023 -8815
rect 5057 -8849 5095 -8815
rect 5129 -8849 5167 -8815
rect 5201 -8849 5239 -8815
rect 5273 -8849 5311 -8815
rect 5345 -8849 5383 -8815
rect 5417 -8849 5455 -8815
rect 5489 -8849 5527 -8815
rect 5561 -8849 5599 -8815
rect 5633 -8849 5671 -8815
rect 5705 -8849 5743 -8815
rect 5777 -8849 5815 -8815
rect 5849 -8849 5887 -8815
rect 5921 -8849 5959 -8815
rect 5993 -8849 6031 -8815
rect 6065 -8849 6103 -8815
rect 6137 -8849 6175 -8815
rect 6209 -8849 6247 -8815
rect 6281 -8849 6319 -8815
rect 6353 -8849 6391 -8815
rect 6425 -8849 6463 -8815
rect 6497 -8849 6535 -8815
rect 6569 -8849 6607 -8815
rect 6641 -8849 6679 -8815
rect 6713 -8849 6751 -8815
rect 6785 -8849 6823 -8815
rect 6857 -8849 6895 -8815
rect 6929 -8849 6967 -8815
rect 7001 -8849 7039 -8815
rect 7073 -8849 7111 -8815
rect 7145 -8849 7183 -8815
rect 7217 -8849 7255 -8815
rect 7289 -8849 7327 -8815
rect 7361 -8849 7399 -8815
rect 7433 -8849 7471 -8815
rect 7505 -8849 7543 -8815
rect 7577 -8849 7615 -8815
rect 7649 -8849 7687 -8815
rect 7721 -8849 7759 -8815
rect 7793 -8849 7831 -8815
rect 7865 -8849 7903 -8815
rect 7937 -8849 7975 -8815
rect 8009 -8849 8047 -8815
rect 8081 -8849 8119 -8815
rect 8153 -8849 8191 -8815
rect 8225 -8849 8263 -8815
rect 8297 -8849 8335 -8815
rect 8369 -8849 8407 -8815
rect 8441 -8849 8479 -8815
rect 8513 -8849 8551 -8815
rect 8585 -8849 8623 -8815
rect 8657 -8849 8695 -8815
rect 8729 -8849 8767 -8815
rect 8801 -8849 8839 -8815
rect 8873 -8849 8911 -8815
rect 8945 -8849 8983 -8815
rect 9017 -8849 9055 -8815
rect 9089 -8849 9127 -8815
rect 9161 -8849 9199 -8815
rect 9233 -8849 9271 -8815
rect 9305 -8849 9343 -8815
rect 9377 -8849 9415 -8815
rect 9449 -8849 9487 -8815
rect 9521 -8849 9559 -8815
rect 9593 -8849 9631 -8815
rect 9665 -8849 9703 -8815
rect 9737 -8849 9775 -8815
rect 9809 -8849 9847 -8815
rect 9881 -8849 9919 -8815
rect 9953 -8849 9991 -8815
rect 10025 -8849 10063 -8815
rect 10097 -8849 10135 -8815
rect 10169 -8849 10207 -8815
rect 10241 -8849 10279 -8815
rect 10313 -8849 10351 -8815
rect 10385 -8849 10423 -8815
rect 10457 -8849 10495 -8815
rect 10529 -8849 10567 -8815
rect 10601 -8849 10639 -8815
rect 10673 -8849 10711 -8815
rect 10745 -8849 10783 -8815
rect 10817 -8849 10855 -8815
rect 10889 -8849 10927 -8815
rect 10961 -8849 10999 -8815
rect 11033 -8849 11071 -8815
rect 11105 -8849 11143 -8815
rect 11177 -8849 11215 -8815
rect 11249 -8849 11287 -8815
rect 11321 -8849 11359 -8815
rect 11393 -8849 11431 -8815
rect 11465 -8849 11503 -8815
rect 11537 -8849 11575 -8815
rect 11609 -8849 11647 -8815
rect 11681 -8849 11719 -8815
rect 11753 -8849 11791 -8815
rect 11825 -8849 11863 -8815
rect 11897 -8849 11935 -8815
rect 11969 -8849 12007 -8815
rect 12041 -8849 12079 -8815
rect 12113 -8849 12151 -8815
rect 12185 -8849 12223 -8815
rect 12257 -8849 12295 -8815
rect 12329 -8849 12367 -8815
rect 12401 -8849 12439 -8815
rect 12473 -8849 12511 -8815
rect 12545 -8849 12583 -8815
rect 12617 -8849 12655 -8815
rect 12689 -8849 12727 -8815
rect 12761 -8849 12799 -8815
rect 12833 -8849 12871 -8815
rect 12905 -8849 12943 -8815
rect 12977 -8849 13015 -8815
rect 13049 -8849 13087 -8815
rect 13121 -8849 13159 -8815
rect 13193 -8849 13231 -8815
rect 13265 -8849 13303 -8815
rect 13337 -8849 13375 -8815
rect 13409 -8849 13447 -8815
rect 13481 -8849 13519 -8815
rect 13553 -8849 13591 -8815
rect 13625 -8849 13663 -8815
rect 13697 -8849 13735 -8815
rect 13769 -8849 13807 -8815
rect 13841 -8849 13879 -8815
rect 13913 -8849 13951 -8815
rect 13985 -8849 14023 -8815
rect 14057 -8849 14095 -8815
rect 14129 -8849 14167 -8815
rect 14201 -8849 14239 -8815
rect 14273 -8849 14311 -8815
rect 14345 -8849 14383 -8815
rect 14417 -8849 14455 -8815
rect 14489 -8849 14527 -8815
rect 14561 -8849 14599 -8815
rect 14633 -8849 14671 -8815
rect 14705 -8849 14743 -8815
rect 14777 -8849 14815 -8815
rect 14849 -8849 14887 -8815
rect 14921 -8849 14959 -8815
rect 14993 -8849 15031 -8815
rect 15065 -8849 15103 -8815
rect 15137 -8849 15175 -8815
rect 15209 -8849 15247 -8815
rect 15281 -8849 15319 -8815
rect 15353 -8849 15391 -8815
rect 15425 -8849 15463 -8815
rect 15497 -8849 15535 -8815
rect 15569 -8849 15607 -8815
rect 15641 -8849 15679 -8815
rect 15713 -8849 15751 -8815
rect 15785 -8849 15823 -8815
rect 15857 -8849 15895 -8815
rect 15929 -8849 15967 -8815
rect 16001 -8849 16039 -8815
rect 16073 -8849 16111 -8815
rect 16145 -8849 16183 -8815
rect 16217 -8849 16255 -8815
rect 16289 -8849 16327 -8815
rect 16361 -8849 16399 -8815
rect 16433 -8849 16471 -8815
rect 16505 -8849 16543 -8815
rect 16577 -8849 16615 -8815
rect 16649 -8849 16687 -8815
rect 16721 -8849 16759 -8815
rect 16793 -8849 16831 -8815
rect 16865 -8849 16903 -8815
rect 16937 -8849 16975 -8815
rect 17009 -8849 17047 -8815
rect 17081 -8849 17119 -8815
rect 17153 -8849 17191 -8815
rect 17225 -8849 17263 -8815
rect 17297 -8849 17335 -8815
rect 17369 -8849 17407 -8815
rect 17441 -8849 17479 -8815
rect 17513 -8849 17551 -8815
rect 17585 -8849 17623 -8815
rect 17657 -8849 17695 -8815
rect 17729 -8849 17767 -8815
rect 17801 -8849 17839 -8815
rect 17873 -8849 17911 -8815
rect 17945 -8849 17983 -8815
rect 18017 -8849 18055 -8815
rect 18089 -8849 18127 -8815
rect 18161 -8849 18199 -8815
rect 18233 -8849 18271 -8815
rect 18305 -8849 18343 -8815
rect 18377 -8849 18415 -8815
rect 18449 -8849 18487 -8815
rect 18521 -8849 18559 -8815
rect 18593 -8849 18631 -8815
rect 18665 -8849 18703 -8815
rect 18737 -8849 18775 -8815
rect 18809 -8849 18847 -8815
rect 18881 -8849 18919 -8815
rect 18953 -8849 18991 -8815
rect 19025 -8849 19063 -8815
rect 19097 -8849 19135 -8815
rect 19169 -8849 19207 -8815
rect 19241 -8849 19279 -8815
rect 19313 -8849 19351 -8815
rect 19385 -8849 19423 -8815
rect 19457 -8849 19495 -8815
rect 19529 -8849 19567 -8815
rect 19601 -8849 19639 -8815
rect 19673 -8849 19711 -8815
rect 19745 -8849 19783 -8815
rect 19817 -8849 19855 -8815
rect 19889 -8849 19927 -8815
rect 19961 -8849 19999 -8815
rect 20033 -8849 20071 -8815
rect 20105 -8849 20143 -8815
rect 20177 -8849 20215 -8815
rect 20249 -8849 20287 -8815
rect 20321 -8849 20359 -8815
rect 20393 -8849 20431 -8815
rect 20465 -8849 20503 -8815
rect 20537 -8849 20575 -8815
rect 20609 -8849 20647 -8815
rect 20681 -8849 20719 -8815
rect 20753 -8849 20791 -8815
rect 20825 -8849 20863 -8815
rect 20897 -8849 20935 -8815
rect 20969 -8849 21007 -8815
rect 21041 -8849 21079 -8815
rect 21113 -8849 21151 -8815
rect 21185 -8849 21223 -8815
rect 21257 -8849 21295 -8815
rect 21329 -8849 21367 -8815
rect 21401 -8849 21439 -8815
rect 21473 -8849 21511 -8815
rect 21545 -8849 21583 -8815
rect 21617 -8849 21655 -8815
rect 21689 -8849 21727 -8815
rect 21761 -8849 21799 -8815
rect 21833 -8849 21871 -8815
rect 21905 -8849 21943 -8815
rect 21977 -8849 22015 -8815
rect 22049 -8849 22087 -8815
rect 22121 -8849 22159 -8815
rect 22193 -8849 22231 -8815
rect 22265 -8849 22303 -8815
rect 22337 -8849 22375 -8815
rect 22409 -8849 22447 -8815
rect 22481 -8849 22519 -8815
rect 22553 -8849 22591 -8815
rect 22625 -8849 22663 -8815
rect 22697 -8849 22735 -8815
rect 22769 -8849 22807 -8815
rect 22841 -8849 22879 -8815
rect 22913 -8849 22951 -8815
rect 22985 -8849 23023 -8815
rect 23057 -8849 23095 -8815
rect 23129 -8849 23167 -8815
rect 23201 -8849 23239 -8815
rect 23273 -8849 23311 -8815
rect 23345 -8849 23383 -8815
rect 23417 -8849 23455 -8815
rect 23489 -8849 23527 -8815
rect 23561 -8849 23599 -8815
rect 23633 -8849 23671 -8815
rect 23705 -8849 23743 -8815
rect 23777 -8849 23815 -8815
rect 23849 -8849 23887 -8815
rect 23921 -8849 23959 -8815
rect 23993 -8849 24031 -8815
rect 24065 -8849 24103 -8815
rect 24137 -8849 24175 -8815
rect 24209 -8849 24247 -8815
rect 24281 -8849 24319 -8815
rect 24353 -8849 24391 -8815
rect 24425 -8849 24463 -8815
rect 24497 -8849 24535 -8815
rect 24569 -8849 24607 -8815
rect 24641 -8849 24679 -8815
rect 24713 -8849 24828 -8815
rect 372 -8888 24828 -8849
rect -645 -11172 -523 -11167
rect -12328 -11200 24928 -11172
rect -12328 -11202 -5014 -11200
rect -12328 -11211 -12008 -11202
rect -11956 -11211 -10214 -11202
rect -10162 -11211 -7614 -11202
rect -7562 -11211 -5014 -11202
rect -4962 -11211 -2414 -11200
rect -2362 -11211 -610 -11200
rect -558 -11211 24928 -11200
rect -12328 -11245 -12221 -11211
rect -12187 -11245 -12149 -11211
rect -12115 -11245 -12077 -11211
rect -12043 -11245 -12008 -11211
rect -11956 -11245 -11933 -11211
rect -11899 -11245 -11861 -11211
rect -11827 -11245 -11789 -11211
rect -11755 -11245 -11717 -11211
rect -11683 -11245 -11645 -11211
rect -11611 -11245 -11573 -11211
rect -11539 -11245 -11501 -11211
rect -11467 -11245 -11429 -11211
rect -11395 -11245 -11357 -11211
rect -11323 -11245 -11285 -11211
rect -11251 -11245 -11213 -11211
rect -11179 -11245 -11141 -11211
rect -11107 -11245 -11069 -11211
rect -11035 -11245 -10997 -11211
rect -10963 -11245 -10925 -11211
rect -10891 -11245 -10853 -11211
rect -10819 -11245 -10781 -11211
rect -10747 -11245 -10709 -11211
rect -10675 -11245 -10637 -11211
rect -10603 -11245 -10565 -11211
rect -10531 -11245 -10493 -11211
rect -10459 -11245 -10421 -11211
rect -10387 -11245 -10349 -11211
rect -10315 -11245 -10277 -11211
rect -10243 -11245 -10214 -11211
rect -10162 -11245 -10133 -11211
rect -10099 -11245 -10061 -11211
rect -10027 -11245 -9989 -11211
rect -9955 -11245 -9917 -11211
rect -9883 -11245 -9845 -11211
rect -9811 -11245 -9773 -11211
rect -9739 -11245 -9701 -11211
rect -9667 -11245 -9629 -11211
rect -9595 -11245 -9557 -11211
rect -9523 -11245 -9485 -11211
rect -9451 -11245 -9413 -11211
rect -9379 -11245 -9341 -11211
rect -9307 -11245 -9269 -11211
rect -9235 -11245 -9197 -11211
rect -9163 -11245 -9125 -11211
rect -9091 -11245 -9053 -11211
rect -9019 -11245 -8981 -11211
rect -8947 -11245 -8909 -11211
rect -8875 -11245 -8837 -11211
rect -8803 -11245 -8765 -11211
rect -8731 -11245 -8693 -11211
rect -8659 -11245 -8621 -11211
rect -8587 -11245 -8549 -11211
rect -8515 -11245 -8477 -11211
rect -8443 -11245 -8405 -11211
rect -8371 -11245 -8333 -11211
rect -8299 -11245 -8261 -11211
rect -8227 -11245 -8189 -11211
rect -8155 -11245 -8117 -11211
rect -8083 -11245 -8045 -11211
rect -8011 -11245 -7973 -11211
rect -7939 -11245 -7901 -11211
rect -7867 -11245 -7829 -11211
rect -7795 -11245 -7757 -11211
rect -7723 -11245 -7685 -11211
rect -7651 -11245 -7614 -11211
rect -7562 -11245 -7541 -11211
rect -7507 -11245 -7469 -11211
rect -7435 -11245 -7397 -11211
rect -7363 -11245 -7325 -11211
rect -7291 -11245 -7253 -11211
rect -7219 -11245 -7181 -11211
rect -7147 -11245 -7109 -11211
rect -7075 -11245 -7037 -11211
rect -7003 -11245 -6965 -11211
rect -6931 -11245 -6893 -11211
rect -6859 -11245 -6821 -11211
rect -6787 -11245 -6749 -11211
rect -6715 -11245 -6677 -11211
rect -6643 -11245 -6605 -11211
rect -6571 -11245 -6533 -11211
rect -6499 -11245 -6461 -11211
rect -6427 -11245 -6389 -11211
rect -6355 -11245 -6317 -11211
rect -6283 -11245 -6245 -11211
rect -6211 -11245 -6173 -11211
rect -6139 -11245 -6101 -11211
rect -6067 -11245 -6029 -11211
rect -5995 -11245 -5957 -11211
rect -5923 -11245 -5885 -11211
rect -5851 -11245 -5813 -11211
rect -5779 -11245 -5741 -11211
rect -5707 -11245 -5669 -11211
rect -5635 -11245 -5597 -11211
rect -5563 -11245 -5525 -11211
rect -5491 -11245 -5453 -11211
rect -5419 -11245 -5381 -11211
rect -5347 -11245 -5309 -11211
rect -5275 -11245 -5237 -11211
rect -5203 -11245 -5165 -11211
rect -5131 -11245 -5093 -11211
rect -5059 -11245 -5021 -11211
rect -4962 -11245 -4949 -11211
rect -4915 -11245 -4877 -11211
rect -4843 -11245 -4805 -11211
rect -4771 -11245 -4733 -11211
rect -4699 -11245 -4661 -11211
rect -4627 -11245 -4589 -11211
rect -4555 -11245 -4517 -11211
rect -4483 -11245 -4445 -11211
rect -4411 -11245 -4373 -11211
rect -4339 -11245 -4301 -11211
rect -4267 -11245 -4229 -11211
rect -4195 -11245 -4157 -11211
rect -4123 -11245 -4085 -11211
rect -4051 -11245 -4013 -11211
rect -3979 -11245 -3941 -11211
rect -3907 -11245 -3869 -11211
rect -3835 -11245 -3797 -11211
rect -3763 -11245 -3725 -11211
rect -3691 -11245 -3653 -11211
rect -3619 -11245 -3581 -11211
rect -3547 -11245 -3509 -11211
rect -3475 -11245 -3437 -11211
rect -3403 -11245 -3365 -11211
rect -3331 -11245 -3293 -11211
rect -3259 -11245 -3221 -11211
rect -3187 -11245 -3149 -11211
rect -3115 -11245 -3077 -11211
rect -3043 -11245 -3005 -11211
rect -2971 -11245 -2933 -11211
rect -2899 -11245 -2861 -11211
rect -2827 -11245 -2789 -11211
rect -2755 -11245 -2717 -11211
rect -2683 -11245 -2645 -11211
rect -2611 -11245 -2573 -11211
rect -2539 -11245 -2501 -11211
rect -2467 -11245 -2429 -11211
rect -2362 -11245 -2357 -11211
rect -2323 -11245 -2285 -11211
rect -2251 -11245 -2213 -11211
rect -2179 -11245 -2141 -11211
rect -2107 -11245 -2069 -11211
rect -2035 -11245 -1997 -11211
rect -1963 -11245 -1925 -11211
rect -1891 -11245 -1853 -11211
rect -1819 -11245 -1781 -11211
rect -1747 -11245 -1709 -11211
rect -1675 -11245 -1637 -11211
rect -1603 -11245 -1565 -11211
rect -1531 -11245 -1493 -11211
rect -1459 -11245 -1421 -11211
rect -1387 -11245 -1349 -11211
rect -1315 -11245 -1277 -11211
rect -1243 -11245 -1205 -11211
rect -1171 -11245 -1133 -11211
rect -1099 -11245 -1061 -11211
rect -1027 -11245 -989 -11211
rect -955 -11245 -917 -11211
rect -883 -11245 -845 -11211
rect -811 -11245 -773 -11211
rect -739 -11245 -701 -11211
rect -667 -11245 -629 -11211
rect -558 -11245 -557 -11211
rect -523 -11245 -485 -11211
rect -451 -11245 -413 -11211
rect -379 -11245 -341 -11211
rect -307 -11245 -269 -11211
rect -235 -11245 -197 -11211
rect -163 -11245 -125 -11211
rect -91 -11245 -53 -11211
rect -19 -11245 19 -11211
rect 53 -11245 91 -11211
rect 125 -11245 163 -11211
rect 197 -11245 235 -11211
rect 269 -11245 307 -11211
rect 341 -11245 379 -11211
rect 413 -11245 451 -11211
rect 485 -11245 523 -11211
rect 557 -11245 595 -11211
rect 629 -11245 667 -11211
rect 701 -11245 739 -11211
rect 773 -11245 811 -11211
rect 845 -11245 883 -11211
rect 917 -11245 955 -11211
rect 989 -11245 1027 -11211
rect 1061 -11245 1099 -11211
rect 1133 -11245 1171 -11211
rect 1205 -11245 1243 -11211
rect 1277 -11245 1315 -11211
rect 1349 -11245 1387 -11211
rect 1421 -11245 1459 -11211
rect 1493 -11245 1531 -11211
rect 1565 -11245 1603 -11211
rect 1637 -11245 1675 -11211
rect 1709 -11245 1747 -11211
rect 1781 -11245 1819 -11211
rect 1853 -11245 1891 -11211
rect 1925 -11245 1963 -11211
rect 1997 -11245 2035 -11211
rect 2069 -11245 2107 -11211
rect 2141 -11245 2179 -11211
rect 2213 -11245 2251 -11211
rect 2285 -11245 2323 -11211
rect 2357 -11245 2395 -11211
rect 2429 -11245 2467 -11211
rect 2501 -11245 2539 -11211
rect 2573 -11245 2611 -11211
rect 2645 -11245 2683 -11211
rect 2717 -11245 2755 -11211
rect 2789 -11245 2827 -11211
rect 2861 -11245 2899 -11211
rect 2933 -11245 2971 -11211
rect 3005 -11245 3043 -11211
rect 3077 -11245 3115 -11211
rect 3149 -11245 3187 -11211
rect 3221 -11245 3259 -11211
rect 3293 -11245 3331 -11211
rect 3365 -11245 3403 -11211
rect 3437 -11245 3475 -11211
rect 3509 -11245 3547 -11211
rect 3581 -11245 3619 -11211
rect 3653 -11245 3691 -11211
rect 3725 -11245 3763 -11211
rect 3797 -11245 3835 -11211
rect 3869 -11245 3907 -11211
rect 3941 -11245 3979 -11211
rect 4013 -11245 4051 -11211
rect 4085 -11245 4123 -11211
rect 4157 -11245 4195 -11211
rect 4229 -11245 4267 -11211
rect 4301 -11245 4339 -11211
rect 4373 -11245 4411 -11211
rect 4445 -11245 4483 -11211
rect 4517 -11245 4555 -11211
rect 4589 -11245 4627 -11211
rect 4661 -11245 4699 -11211
rect 4733 -11245 4771 -11211
rect 4805 -11245 4843 -11211
rect 4877 -11245 4915 -11211
rect 4949 -11245 4987 -11211
rect 5021 -11245 5059 -11211
rect 5093 -11245 5131 -11211
rect 5165 -11245 5203 -11211
rect 5237 -11245 5275 -11211
rect 5309 -11245 5347 -11211
rect 5381 -11245 5419 -11211
rect 5453 -11245 5491 -11211
rect 5525 -11245 5563 -11211
rect 5597 -11245 5635 -11211
rect 5669 -11245 5707 -11211
rect 5741 -11245 5779 -11211
rect 5813 -11245 5851 -11211
rect 5885 -11245 5923 -11211
rect 5957 -11245 5995 -11211
rect 6029 -11245 6067 -11211
rect 6101 -11245 6139 -11211
rect 6173 -11245 6211 -11211
rect 6245 -11245 6283 -11211
rect 6317 -11245 6355 -11211
rect 6389 -11245 6427 -11211
rect 6461 -11245 6499 -11211
rect 6533 -11245 6571 -11211
rect 6605 -11245 6643 -11211
rect 6677 -11245 6715 -11211
rect 6749 -11245 6787 -11211
rect 6821 -11245 6859 -11211
rect 6893 -11245 6931 -11211
rect 6965 -11245 7003 -11211
rect 7037 -11245 7075 -11211
rect 7109 -11245 7147 -11211
rect 7181 -11245 7219 -11211
rect 7253 -11245 7291 -11211
rect 7325 -11245 7363 -11211
rect 7397 -11245 7435 -11211
rect 7469 -11245 7507 -11211
rect 7541 -11245 7579 -11211
rect 7613 -11245 7651 -11211
rect 7685 -11245 7723 -11211
rect 7757 -11245 7795 -11211
rect 7829 -11245 7867 -11211
rect 7901 -11245 7939 -11211
rect 7973 -11245 8011 -11211
rect 8045 -11245 8083 -11211
rect 8117 -11245 8155 -11211
rect 8189 -11245 8227 -11211
rect 8261 -11245 8299 -11211
rect 8333 -11245 8371 -11211
rect 8405 -11245 8443 -11211
rect 8477 -11245 8515 -11211
rect 8549 -11245 8587 -11211
rect 8621 -11245 8659 -11211
rect 8693 -11245 8731 -11211
rect 8765 -11245 8803 -11211
rect 8837 -11245 8875 -11211
rect 8909 -11245 8947 -11211
rect 8981 -11245 9019 -11211
rect 9053 -11245 9091 -11211
rect 9125 -11245 9163 -11211
rect 9197 -11245 9235 -11211
rect 9269 -11245 9307 -11211
rect 9341 -11245 9379 -11211
rect 9413 -11245 9451 -11211
rect 9485 -11245 9523 -11211
rect 9557 -11245 9595 -11211
rect 9629 -11245 9667 -11211
rect 9701 -11245 9739 -11211
rect 9773 -11245 9811 -11211
rect 9845 -11245 9883 -11211
rect 9917 -11245 9955 -11211
rect 9989 -11245 10027 -11211
rect 10061 -11245 10099 -11211
rect 10133 -11245 10171 -11211
rect 10205 -11245 10243 -11211
rect 10277 -11245 10315 -11211
rect 10349 -11245 10387 -11211
rect 10421 -11245 10459 -11211
rect 10493 -11245 10531 -11211
rect 10565 -11245 10603 -11211
rect 10637 -11245 10675 -11211
rect 10709 -11245 10747 -11211
rect 10781 -11245 10819 -11211
rect 10853 -11245 10891 -11211
rect 10925 -11245 10963 -11211
rect 10997 -11245 11035 -11211
rect 11069 -11245 11107 -11211
rect 11141 -11245 11179 -11211
rect 11213 -11245 11251 -11211
rect 11285 -11245 11323 -11211
rect 11357 -11245 11395 -11211
rect 11429 -11245 11467 -11211
rect 11501 -11245 11539 -11211
rect 11573 -11245 11611 -11211
rect 11645 -11245 11683 -11211
rect 11717 -11245 11755 -11211
rect 11789 -11245 11827 -11211
rect 11861 -11245 11899 -11211
rect 11933 -11245 11971 -11211
rect 12005 -11245 12043 -11211
rect 12077 -11245 12115 -11211
rect 12149 -11245 12187 -11211
rect 12221 -11245 12259 -11211
rect 12293 -11245 12331 -11211
rect 12365 -11245 12403 -11211
rect 12437 -11245 12475 -11211
rect 12509 -11245 12547 -11211
rect 12581 -11245 12619 -11211
rect 12653 -11245 12691 -11211
rect 12725 -11245 12763 -11211
rect 12797 -11245 12835 -11211
rect 12869 -11245 12907 -11211
rect 12941 -11245 12979 -11211
rect 13013 -11245 13051 -11211
rect 13085 -11245 13123 -11211
rect 13157 -11245 13195 -11211
rect 13229 -11245 13267 -11211
rect 13301 -11245 13339 -11211
rect 13373 -11245 13411 -11211
rect 13445 -11245 13483 -11211
rect 13517 -11245 13555 -11211
rect 13589 -11245 13627 -11211
rect 13661 -11245 13699 -11211
rect 13733 -11245 13771 -11211
rect 13805 -11245 13843 -11211
rect 13877 -11245 13915 -11211
rect 13949 -11245 13987 -11211
rect 14021 -11245 14059 -11211
rect 14093 -11245 14131 -11211
rect 14165 -11245 14203 -11211
rect 14237 -11245 14275 -11211
rect 14309 -11245 14347 -11211
rect 14381 -11245 14419 -11211
rect 14453 -11245 14491 -11211
rect 14525 -11245 14563 -11211
rect 14597 -11245 14635 -11211
rect 14669 -11245 14707 -11211
rect 14741 -11245 14779 -11211
rect 14813 -11245 14851 -11211
rect 14885 -11245 14923 -11211
rect 14957 -11245 14995 -11211
rect 15029 -11245 15067 -11211
rect 15101 -11245 15139 -11211
rect 15173 -11245 15211 -11211
rect 15245 -11245 15283 -11211
rect 15317 -11245 15355 -11211
rect 15389 -11245 15427 -11211
rect 15461 -11245 15499 -11211
rect 15533 -11245 15571 -11211
rect 15605 -11245 15643 -11211
rect 15677 -11245 15715 -11211
rect 15749 -11245 15787 -11211
rect 15821 -11245 15859 -11211
rect 15893 -11245 15931 -11211
rect 15965 -11245 16003 -11211
rect 16037 -11245 16075 -11211
rect 16109 -11245 16147 -11211
rect 16181 -11245 16219 -11211
rect 16253 -11245 16291 -11211
rect 16325 -11245 16363 -11211
rect 16397 -11245 16435 -11211
rect 16469 -11245 16507 -11211
rect 16541 -11245 16579 -11211
rect 16613 -11245 16651 -11211
rect 16685 -11245 16723 -11211
rect 16757 -11245 16795 -11211
rect 16829 -11245 16867 -11211
rect 16901 -11245 16939 -11211
rect 16973 -11245 17011 -11211
rect 17045 -11245 17083 -11211
rect 17117 -11245 17155 -11211
rect 17189 -11245 17227 -11211
rect 17261 -11245 17299 -11211
rect 17333 -11245 17371 -11211
rect 17405 -11245 17443 -11211
rect 17477 -11245 17515 -11211
rect 17549 -11245 17587 -11211
rect 17621 -11245 17659 -11211
rect 17693 -11245 17731 -11211
rect 17765 -11245 17803 -11211
rect 17837 -11245 17875 -11211
rect 17909 -11245 17947 -11211
rect 17981 -11245 18019 -11211
rect 18053 -11245 18091 -11211
rect 18125 -11245 18163 -11211
rect 18197 -11245 18235 -11211
rect 18269 -11245 18307 -11211
rect 18341 -11245 18379 -11211
rect 18413 -11245 18451 -11211
rect 18485 -11245 18523 -11211
rect 18557 -11245 18595 -11211
rect 18629 -11245 18667 -11211
rect 18701 -11245 18739 -11211
rect 18773 -11245 18811 -11211
rect 18845 -11245 18883 -11211
rect 18917 -11245 18955 -11211
rect 18989 -11245 19027 -11211
rect 19061 -11245 19099 -11211
rect 19133 -11245 19171 -11211
rect 19205 -11245 19243 -11211
rect 19277 -11245 19315 -11211
rect 19349 -11245 19387 -11211
rect 19421 -11245 19459 -11211
rect 19493 -11245 19531 -11211
rect 19565 -11245 19603 -11211
rect 19637 -11245 19675 -11211
rect 19709 -11245 19747 -11211
rect 19781 -11245 19819 -11211
rect 19853 -11245 19891 -11211
rect 19925 -11245 19963 -11211
rect 19997 -11245 20035 -11211
rect 20069 -11245 20107 -11211
rect 20141 -11245 20179 -11211
rect 20213 -11245 20251 -11211
rect 20285 -11245 20323 -11211
rect 20357 -11245 20395 -11211
rect 20429 -11245 20467 -11211
rect 20501 -11245 20539 -11211
rect 20573 -11245 20611 -11211
rect 20645 -11245 20683 -11211
rect 20717 -11245 20755 -11211
rect 20789 -11245 20827 -11211
rect 20861 -11245 20899 -11211
rect 20933 -11245 20971 -11211
rect 21005 -11245 21043 -11211
rect 21077 -11245 21115 -11211
rect 21149 -11245 21187 -11211
rect 21221 -11245 21259 -11211
rect 21293 -11245 21331 -11211
rect 21365 -11245 21403 -11211
rect 21437 -11245 21475 -11211
rect 21509 -11245 21547 -11211
rect 21581 -11245 21619 -11211
rect 21653 -11245 21691 -11211
rect 21725 -11245 21763 -11211
rect 21797 -11245 21835 -11211
rect 21869 -11245 21907 -11211
rect 21941 -11245 21979 -11211
rect 22013 -11245 22051 -11211
rect 22085 -11245 22123 -11211
rect 22157 -11245 22195 -11211
rect 22229 -11245 22267 -11211
rect 22301 -11245 22339 -11211
rect 22373 -11245 22411 -11211
rect 22445 -11245 22483 -11211
rect 22517 -11245 22555 -11211
rect 22589 -11245 22627 -11211
rect 22661 -11245 22699 -11211
rect 22733 -11245 22771 -11211
rect 22805 -11245 22843 -11211
rect 22877 -11245 22915 -11211
rect 22949 -11245 22987 -11211
rect 23021 -11245 23059 -11211
rect 23093 -11245 23131 -11211
rect 23165 -11245 23203 -11211
rect 23237 -11245 23275 -11211
rect 23309 -11245 23347 -11211
rect 23381 -11245 23419 -11211
rect 23453 -11245 23491 -11211
rect 23525 -11245 23563 -11211
rect 23597 -11245 23635 -11211
rect 23669 -11245 23707 -11211
rect 23741 -11245 23779 -11211
rect 23813 -11245 23851 -11211
rect 23885 -11245 23923 -11211
rect 23957 -11245 23995 -11211
rect 24029 -11245 24067 -11211
rect 24101 -11245 24139 -11211
rect 24173 -11245 24211 -11211
rect 24245 -11245 24283 -11211
rect 24317 -11245 24355 -11211
rect 24389 -11245 24427 -11211
rect 24461 -11245 24499 -11211
rect 24533 -11245 24571 -11211
rect 24605 -11245 24643 -11211
rect 24677 -11245 24715 -11211
rect 24749 -11245 24787 -11211
rect 24821 -11245 24928 -11211
rect -12328 -11254 -12008 -11245
rect -11956 -11254 -10214 -11245
rect -10162 -11254 -7614 -11245
rect -7562 -11252 -5014 -11245
rect -4962 -11252 -2414 -11245
rect -2362 -11252 -610 -11245
rect -558 -11252 24928 -11245
rect -7562 -11254 24928 -11252
rect -12328 -11284 24928 -11254
rect -12328 -12091 -12216 -11284
rect 1948 -11352 2020 -11348
rect 1948 -11404 1958 -11352
rect 2010 -11404 2020 -11352
rect 1948 -11408 2020 -11404
rect 2104 -11352 2176 -11348
rect 2104 -11404 2114 -11352
rect 2166 -11404 2176 -11352
rect 2104 -11408 2176 -11404
rect 2336 -11360 2396 -11350
rect -12328 -12125 -12289 -12091
rect -12255 -12125 -12216 -12091
rect -12328 -12163 -12216 -12125
rect -12328 -12197 -12289 -12163
rect -12255 -12197 -12216 -12163
rect 1954 -12186 2014 -11408
rect -12328 -12235 -12216 -12197
rect -12328 -12269 -12289 -12235
rect -12255 -12269 -12216 -12235
rect -12328 -12307 -12216 -12269
rect -12328 -12341 -12289 -12307
rect -12255 -12341 -12216 -12307
rect -2072 -12246 2014 -12186
rect -2072 -12324 -2012 -12246
rect -12328 -12379 -12216 -12341
rect -12328 -12413 -12289 -12379
rect -12255 -12413 -12216 -12379
rect -12328 -12451 -12216 -12413
rect -12328 -12485 -12289 -12451
rect -12255 -12485 -12216 -12451
rect -12328 -12523 -12216 -12485
rect -12328 -12557 -12289 -12523
rect -12255 -12557 -12216 -12523
rect -9196 -12384 -2012 -12324
rect -9196 -12543 -9136 -12384
rect -8686 -12434 -8626 -12384
rect -8902 -12440 -8414 -12434
rect -8902 -12474 -8855 -12440
rect -8821 -12474 -8783 -12440
rect -8749 -12474 -8711 -12440
rect -8677 -12474 -8639 -12440
rect -8605 -12474 -8567 -12440
rect -8533 -12474 -8495 -12440
rect -8461 -12474 -8414 -12440
rect -8902 -12480 -8414 -12474
rect -9196 -12554 -9184 -12543
rect -12328 -12595 -12216 -12557
rect -12328 -12629 -12289 -12595
rect -12255 -12629 -12216 -12595
rect -12328 -12667 -12216 -12629
rect -12328 -12701 -12289 -12667
rect -12255 -12701 -12216 -12667
rect -12328 -12739 -12216 -12701
rect -12328 -12773 -12289 -12739
rect -12255 -12773 -12216 -12739
rect -12328 -12811 -12216 -12773
rect -12328 -12845 -12289 -12811
rect -12255 -12845 -12216 -12811
rect -12328 -12883 -12216 -12845
rect -12328 -12917 -12289 -12883
rect -12255 -12917 -12216 -12883
rect -12328 -12955 -12216 -12917
rect -12328 -12989 -12289 -12955
rect -12255 -12989 -12216 -12955
rect -12328 -13027 -12216 -12989
rect -12328 -13061 -12289 -13027
rect -12255 -13061 -12216 -13027
rect -12328 -13099 -12216 -13061
rect -9190 -12577 -9184 -12554
rect -9150 -12554 -9136 -12543
rect -8180 -12543 -8120 -12384
rect -7678 -12434 -7618 -12384
rect -6650 -12434 -6590 -12384
rect -7884 -12440 -7396 -12434
rect -7884 -12474 -7837 -12440
rect -7803 -12474 -7765 -12440
rect -7731 -12474 -7693 -12440
rect -7659 -12474 -7621 -12440
rect -7587 -12474 -7549 -12440
rect -7515 -12474 -7477 -12440
rect -7443 -12474 -7396 -12440
rect -7884 -12480 -7396 -12474
rect -6866 -12440 -6378 -12434
rect -6866 -12474 -6819 -12440
rect -6785 -12474 -6747 -12440
rect -6713 -12474 -6675 -12440
rect -6641 -12474 -6603 -12440
rect -6569 -12474 -6531 -12440
rect -6497 -12474 -6459 -12440
rect -6425 -12474 -6378 -12440
rect -6866 -12480 -6378 -12474
rect -8180 -12548 -8166 -12543
rect -9150 -12577 -9144 -12554
rect -9190 -12615 -9144 -12577
rect -9190 -12649 -9184 -12615
rect -9150 -12649 -9144 -12615
rect -9190 -12687 -9144 -12649
rect -9190 -12721 -9184 -12687
rect -9150 -12721 -9144 -12687
rect -9190 -12759 -9144 -12721
rect -9190 -12793 -9184 -12759
rect -9150 -12793 -9144 -12759
rect -9190 -12831 -9144 -12793
rect -9190 -12865 -9184 -12831
rect -9150 -12865 -9144 -12831
rect -9190 -12903 -9144 -12865
rect -9190 -12937 -9184 -12903
rect -9150 -12937 -9144 -12903
rect -9190 -12975 -9144 -12937
rect -9190 -13009 -9184 -12975
rect -9150 -13009 -9144 -12975
rect -9190 -13047 -9144 -13009
rect -9190 -13081 -9184 -13047
rect -9150 -13081 -9144 -13047
rect -8172 -12577 -8166 -12548
rect -8132 -12548 -8120 -12543
rect -7154 -12543 -7108 -12512
rect -8132 -12577 -8126 -12548
rect -8172 -12615 -8126 -12577
rect -8172 -12649 -8166 -12615
rect -8132 -12649 -8126 -12615
rect -8172 -12687 -8126 -12649
rect -8172 -12721 -8166 -12687
rect -8132 -12721 -8126 -12687
rect -8172 -12759 -8126 -12721
rect -8172 -12793 -8166 -12759
rect -8132 -12793 -8126 -12759
rect -8172 -12831 -8126 -12793
rect -8172 -12865 -8166 -12831
rect -8132 -12865 -8126 -12831
rect -8172 -12903 -8126 -12865
rect -8172 -12937 -8166 -12903
rect -8132 -12937 -8126 -12903
rect -8172 -12975 -8126 -12937
rect -8172 -13009 -8166 -12975
rect -8132 -13009 -8126 -12975
rect -8172 -13047 -8126 -13009
rect -8172 -13078 -8166 -13047
rect -9190 -13082 -9144 -13081
rect -8180 -13081 -8166 -13078
rect -8132 -13078 -8126 -13047
rect -7154 -12577 -7148 -12543
rect -7114 -12577 -7108 -12543
rect -6142 -12543 -6082 -12384
rect -5636 -12434 -5576 -12384
rect -4622 -12434 -4562 -12384
rect -5848 -12440 -5360 -12434
rect -5848 -12474 -5801 -12440
rect -5767 -12474 -5729 -12440
rect -5695 -12474 -5657 -12440
rect -5623 -12474 -5585 -12440
rect -5551 -12474 -5513 -12440
rect -5479 -12474 -5441 -12440
rect -5407 -12474 -5360 -12440
rect -5848 -12480 -5360 -12474
rect -4830 -12440 -4342 -12434
rect -4830 -12474 -4783 -12440
rect -4749 -12474 -4711 -12440
rect -4677 -12474 -4639 -12440
rect -4605 -12474 -4567 -12440
rect -4533 -12474 -4495 -12440
rect -4461 -12474 -4423 -12440
rect -4389 -12474 -4342 -12440
rect -4830 -12480 -4342 -12474
rect -6142 -12562 -6130 -12543
rect -7154 -12615 -7108 -12577
rect -7154 -12649 -7148 -12615
rect -7114 -12649 -7108 -12615
rect -7154 -12687 -7108 -12649
rect -7154 -12721 -7148 -12687
rect -7114 -12721 -7108 -12687
rect -7154 -12759 -7108 -12721
rect -7154 -12793 -7148 -12759
rect -7114 -12793 -7108 -12759
rect -7154 -12831 -7108 -12793
rect -7154 -12865 -7148 -12831
rect -7114 -12865 -7108 -12831
rect -7154 -12903 -7108 -12865
rect -7154 -12937 -7148 -12903
rect -7114 -12937 -7108 -12903
rect -7154 -12975 -7108 -12937
rect -7154 -13009 -7148 -12975
rect -7114 -13009 -7108 -12975
rect -7154 -13047 -7108 -13009
rect -7154 -13076 -7148 -13047
rect -8132 -13081 -8120 -13078
rect -12328 -13133 -12289 -13099
rect -12255 -13133 -12216 -13099
rect -12328 -13171 -12216 -13133
rect -12328 -13205 -12289 -13171
rect -12255 -13205 -12216 -13171
rect -12328 -13243 -12216 -13205
rect -12328 -13277 -12289 -13243
rect -12255 -13277 -12216 -13243
rect -12328 -13315 -12216 -13277
rect -12328 -13349 -12289 -13315
rect -12255 -13349 -12216 -13315
rect -12328 -13387 -12216 -13349
rect -9200 -13361 -9140 -13082
rect -8902 -13150 -8414 -13144
rect -8902 -13184 -8855 -13150
rect -8821 -13184 -8783 -13150
rect -8749 -13184 -8711 -13150
rect -8677 -13184 -8639 -13150
rect -8605 -13184 -8567 -13150
rect -8533 -13184 -8495 -13150
rect -8461 -13184 -8414 -13150
rect -8902 -13190 -8414 -13184
rect -8686 -13252 -8626 -13190
rect -8902 -13258 -8414 -13252
rect -8902 -13292 -8855 -13258
rect -8821 -13292 -8783 -13258
rect -8749 -13292 -8711 -13258
rect -8677 -13292 -8639 -13258
rect -8605 -13292 -8567 -13258
rect -8533 -13292 -8495 -13258
rect -8461 -13292 -8414 -13258
rect -8902 -13298 -8414 -13292
rect -9200 -13372 -9184 -13361
rect -12328 -13421 -12289 -13387
rect -12255 -13421 -12216 -13387
rect -12328 -13459 -12216 -13421
rect -12328 -13493 -12289 -13459
rect -12255 -13493 -12216 -13459
rect -12328 -13531 -12216 -13493
rect -12328 -13565 -12289 -13531
rect -12255 -13565 -12216 -13531
rect -12328 -13603 -12216 -13565
rect -12328 -13637 -12289 -13603
rect -12255 -13637 -12216 -13603
rect -12328 -13675 -12216 -13637
rect -12328 -13709 -12289 -13675
rect -12255 -13709 -12216 -13675
rect -12328 -13747 -12216 -13709
rect -12328 -13781 -12289 -13747
rect -12255 -13781 -12216 -13747
rect -12328 -13819 -12216 -13781
rect -12328 -13853 -12289 -13819
rect -12255 -13853 -12216 -13819
rect -12328 -13891 -12216 -13853
rect -12328 -13925 -12289 -13891
rect -12255 -13925 -12216 -13891
rect -9190 -13395 -9184 -13372
rect -9150 -13372 -9140 -13361
rect -8180 -13361 -8120 -13081
rect -7160 -13081 -7148 -13076
rect -7114 -13076 -7108 -13047
rect -6136 -12577 -6130 -12562
rect -6096 -12562 -6082 -12543
rect -5118 -12543 -5072 -12512
rect -4106 -12524 -4046 -12384
rect -3590 -12434 -3530 -12384
rect -2584 -12434 -2524 -12384
rect -3812 -12440 -3324 -12434
rect -3812 -12474 -3765 -12440
rect -3731 -12474 -3693 -12440
rect -3659 -12474 -3621 -12440
rect -3587 -12474 -3549 -12440
rect -3515 -12474 -3477 -12440
rect -3443 -12474 -3405 -12440
rect -3371 -12474 -3324 -12440
rect -3812 -12480 -3324 -12474
rect -2794 -12440 -2306 -12434
rect -2794 -12474 -2747 -12440
rect -2713 -12474 -2675 -12440
rect -2641 -12474 -2603 -12440
rect -2569 -12474 -2531 -12440
rect -2497 -12474 -2459 -12440
rect -2425 -12474 -2387 -12440
rect -2353 -12474 -2306 -12440
rect -2794 -12480 -2306 -12474
rect -6096 -12577 -6090 -12562
rect -6136 -12615 -6090 -12577
rect -6136 -12649 -6130 -12615
rect -6096 -12649 -6090 -12615
rect -6136 -12687 -6090 -12649
rect -6136 -12721 -6130 -12687
rect -6096 -12721 -6090 -12687
rect -6136 -12759 -6090 -12721
rect -6136 -12793 -6130 -12759
rect -6096 -12793 -6090 -12759
rect -6136 -12831 -6090 -12793
rect -6136 -12865 -6130 -12831
rect -6096 -12865 -6090 -12831
rect -6136 -12903 -6090 -12865
rect -6136 -12937 -6130 -12903
rect -6096 -12937 -6090 -12903
rect -6136 -12975 -6090 -12937
rect -6136 -13009 -6130 -12975
rect -6096 -13009 -6090 -12975
rect -6136 -13047 -6090 -13009
rect -7114 -13081 -7100 -13076
rect -6136 -13080 -6130 -13047
rect -7884 -13150 -7396 -13144
rect -7884 -13184 -7837 -13150
rect -7803 -13184 -7765 -13150
rect -7731 -13184 -7693 -13150
rect -7659 -13184 -7621 -13150
rect -7587 -13184 -7549 -13150
rect -7515 -13184 -7477 -13150
rect -7443 -13184 -7396 -13150
rect -7884 -13190 -7396 -13184
rect -7682 -13252 -7622 -13190
rect -7884 -13258 -7396 -13252
rect -7884 -13292 -7837 -13258
rect -7803 -13292 -7765 -13258
rect -7731 -13292 -7693 -13258
rect -7659 -13292 -7621 -13258
rect -7587 -13292 -7549 -13258
rect -7515 -13292 -7477 -13258
rect -7443 -13292 -7396 -13258
rect -7884 -13298 -7396 -13292
rect -8180 -13368 -8166 -13361
rect -9150 -13395 -9144 -13372
rect -9190 -13433 -9144 -13395
rect -9190 -13467 -9184 -13433
rect -9150 -13467 -9144 -13433
rect -9190 -13505 -9144 -13467
rect -9190 -13539 -9184 -13505
rect -9150 -13539 -9144 -13505
rect -9190 -13577 -9144 -13539
rect -9190 -13611 -9184 -13577
rect -9150 -13611 -9144 -13577
rect -9190 -13649 -9144 -13611
rect -9190 -13683 -9184 -13649
rect -9150 -13683 -9144 -13649
rect -9190 -13721 -9144 -13683
rect -9190 -13755 -9184 -13721
rect -9150 -13755 -9144 -13721
rect -9190 -13793 -9144 -13755
rect -9190 -13827 -9184 -13793
rect -9150 -13827 -9144 -13793
rect -9190 -13865 -9144 -13827
rect -9190 -13896 -9184 -13865
rect -12328 -13963 -12216 -13925
rect -12328 -13997 -12289 -13963
rect -12255 -13997 -12216 -13963
rect -12328 -14035 -12216 -13997
rect -12328 -14069 -12289 -14035
rect -12255 -14069 -12216 -14035
rect -12328 -14107 -12216 -14069
rect -12328 -14141 -12289 -14107
rect -12255 -14141 -12216 -14107
rect -12328 -14179 -12216 -14141
rect -12328 -14213 -12289 -14179
rect -12255 -14213 -12216 -14179
rect -9198 -13899 -9184 -13896
rect -9150 -13896 -9144 -13865
rect -8172 -13395 -8166 -13368
rect -8132 -13368 -8120 -13361
rect -7160 -13361 -7100 -13081
rect -6142 -13081 -6130 -13080
rect -6096 -13080 -6090 -13047
rect -5118 -12577 -5112 -12543
rect -5078 -12577 -5072 -12543
rect -4108 -12543 -4046 -12524
rect -4108 -12558 -4094 -12543
rect -4106 -12570 -4094 -12558
rect -5118 -12615 -5072 -12577
rect -5118 -12649 -5112 -12615
rect -5078 -12649 -5072 -12615
rect -5118 -12687 -5072 -12649
rect -5118 -12721 -5112 -12687
rect -5078 -12721 -5072 -12687
rect -5118 -12759 -5072 -12721
rect -5118 -12793 -5112 -12759
rect -5078 -12793 -5072 -12759
rect -5118 -12831 -5072 -12793
rect -5118 -12865 -5112 -12831
rect -5078 -12865 -5072 -12831
rect -5118 -12903 -5072 -12865
rect -5118 -12937 -5112 -12903
rect -5078 -12937 -5072 -12903
rect -5118 -12975 -5072 -12937
rect -5118 -13009 -5112 -12975
rect -5078 -13009 -5072 -12975
rect -5118 -13047 -5072 -13009
rect -5118 -13072 -5112 -13047
rect -6096 -13081 -6082 -13080
rect -6866 -13150 -6378 -13144
rect -6866 -13184 -6819 -13150
rect -6785 -13184 -6747 -13150
rect -6713 -13184 -6675 -13150
rect -6641 -13184 -6603 -13150
rect -6569 -13184 -6531 -13150
rect -6497 -13184 -6459 -13150
rect -6425 -13184 -6378 -13150
rect -6866 -13190 -6378 -13184
rect -6652 -13252 -6592 -13190
rect -6866 -13258 -6378 -13252
rect -6866 -13292 -6819 -13258
rect -6785 -13292 -6747 -13258
rect -6713 -13292 -6675 -13258
rect -6641 -13292 -6603 -13258
rect -6569 -13292 -6531 -13258
rect -6497 -13292 -6459 -13258
rect -6425 -13292 -6378 -13258
rect -6866 -13298 -6378 -13292
rect -7160 -13366 -7148 -13361
rect -8132 -13395 -8126 -13368
rect -8172 -13433 -8126 -13395
rect -8172 -13467 -8166 -13433
rect -8132 -13467 -8126 -13433
rect -8172 -13505 -8126 -13467
rect -8172 -13539 -8166 -13505
rect -8132 -13539 -8126 -13505
rect -8172 -13577 -8126 -13539
rect -8172 -13611 -8166 -13577
rect -8132 -13611 -8126 -13577
rect -8172 -13649 -8126 -13611
rect -8172 -13683 -8166 -13649
rect -8132 -13683 -8126 -13649
rect -8172 -13721 -8126 -13683
rect -8172 -13755 -8166 -13721
rect -8132 -13755 -8126 -13721
rect -8172 -13793 -8126 -13755
rect -8172 -13827 -8166 -13793
rect -8132 -13827 -8126 -13793
rect -8172 -13865 -8126 -13827
rect -8172 -13892 -8166 -13865
rect -9150 -13899 -9138 -13896
rect -9198 -14179 -9138 -13899
rect -8178 -13899 -8166 -13892
rect -8132 -13892 -8126 -13865
rect -7154 -13395 -7148 -13366
rect -7114 -13366 -7100 -13361
rect -6142 -13361 -6082 -13081
rect -5122 -13081 -5112 -13072
rect -5078 -13072 -5072 -13047
rect -4100 -12577 -4094 -12570
rect -4060 -12570 -4046 -12543
rect -3082 -12543 -3036 -12512
rect -4060 -12577 -4054 -12570
rect -4100 -12615 -4054 -12577
rect -4100 -12649 -4094 -12615
rect -4060 -12649 -4054 -12615
rect -4100 -12687 -4054 -12649
rect -4100 -12721 -4094 -12687
rect -4060 -12721 -4054 -12687
rect -4100 -12759 -4054 -12721
rect -4100 -12793 -4094 -12759
rect -4060 -12793 -4054 -12759
rect -4100 -12831 -4054 -12793
rect -4100 -12865 -4094 -12831
rect -4060 -12865 -4054 -12831
rect -4100 -12903 -4054 -12865
rect -4100 -12937 -4094 -12903
rect -4060 -12937 -4054 -12903
rect -4100 -12975 -4054 -12937
rect -4100 -13009 -4094 -12975
rect -4060 -13009 -4054 -12975
rect -4100 -13047 -4054 -13009
rect -5078 -13081 -5062 -13072
rect -4100 -13080 -4094 -13047
rect -5848 -13150 -5360 -13144
rect -5848 -13184 -5801 -13150
rect -5767 -13184 -5729 -13150
rect -5695 -13184 -5657 -13150
rect -5623 -13184 -5585 -13150
rect -5551 -13184 -5513 -13150
rect -5479 -13184 -5441 -13150
rect -5407 -13184 -5360 -13150
rect -5848 -13190 -5360 -13184
rect -5650 -13252 -5590 -13190
rect -5848 -13258 -5360 -13252
rect -5848 -13292 -5801 -13258
rect -5767 -13292 -5729 -13258
rect -5695 -13292 -5657 -13258
rect -5623 -13292 -5585 -13258
rect -5551 -13292 -5513 -13258
rect -5479 -13292 -5441 -13258
rect -5407 -13292 -5360 -13258
rect -5848 -13298 -5360 -13292
rect -7114 -13395 -7108 -13366
rect -6142 -13370 -6130 -13361
rect -7154 -13433 -7108 -13395
rect -7154 -13467 -7148 -13433
rect -7114 -13467 -7108 -13433
rect -7154 -13505 -7108 -13467
rect -7154 -13539 -7148 -13505
rect -7114 -13539 -7108 -13505
rect -7154 -13577 -7108 -13539
rect -7154 -13611 -7148 -13577
rect -7114 -13611 -7108 -13577
rect -7154 -13649 -7108 -13611
rect -7154 -13683 -7148 -13649
rect -7114 -13683 -7108 -13649
rect -7154 -13721 -7108 -13683
rect -7154 -13755 -7148 -13721
rect -7114 -13755 -7108 -13721
rect -7154 -13793 -7108 -13755
rect -7154 -13827 -7148 -13793
rect -7114 -13827 -7108 -13793
rect -7154 -13865 -7108 -13827
rect -7154 -13890 -7148 -13865
rect -8132 -13899 -8118 -13892
rect -8902 -13968 -8414 -13962
rect -8902 -14002 -8855 -13968
rect -8821 -14002 -8783 -13968
rect -8749 -14002 -8711 -13968
rect -8677 -14002 -8639 -13968
rect -8605 -14002 -8567 -13968
rect -8533 -14002 -8495 -13968
rect -8461 -14002 -8414 -13968
rect -8902 -14008 -8414 -14002
rect -8686 -14070 -8626 -14008
rect -8902 -14076 -8414 -14070
rect -8902 -14110 -8855 -14076
rect -8821 -14110 -8783 -14076
rect -8749 -14110 -8711 -14076
rect -8677 -14110 -8639 -14076
rect -8605 -14110 -8567 -14076
rect -8533 -14110 -8495 -14076
rect -8461 -14110 -8414 -14076
rect -8902 -14116 -8414 -14110
rect -9198 -14186 -9184 -14179
rect -12328 -14251 -12216 -14213
rect -12328 -14285 -12289 -14251
rect -12255 -14285 -12216 -14251
rect -12328 -14323 -12216 -14285
rect -12328 -14357 -12289 -14323
rect -12255 -14357 -12216 -14323
rect -12328 -14395 -12216 -14357
rect -12328 -14429 -12289 -14395
rect -12255 -14429 -12216 -14395
rect -12328 -14467 -12216 -14429
rect -12328 -14501 -12289 -14467
rect -12255 -14501 -12216 -14467
rect -12328 -14539 -12216 -14501
rect -12328 -14573 -12289 -14539
rect -12255 -14573 -12216 -14539
rect -12328 -14611 -12216 -14573
rect -12328 -14645 -12289 -14611
rect -12255 -14645 -12216 -14611
rect -12328 -14683 -12216 -14645
rect -12328 -14717 -12289 -14683
rect -12255 -14717 -12216 -14683
rect -12328 -14755 -12216 -14717
rect -9190 -14213 -9184 -14186
rect -9150 -14186 -9138 -14179
rect -8178 -14179 -8118 -13899
rect -7158 -13899 -7148 -13890
rect -7114 -13890 -7108 -13865
rect -6136 -13395 -6130 -13370
rect -6096 -13370 -6082 -13361
rect -5122 -13361 -5062 -13081
rect -4110 -13081 -4094 -13080
rect -4060 -13080 -4054 -13047
rect -3082 -12577 -3076 -12543
rect -3042 -12577 -3036 -12543
rect -2072 -12543 -2012 -12384
rect -1562 -12434 -1502 -12246
rect 1184 -12334 1244 -12328
rect -32 -12338 1244 -12334
rect -32 -12390 1188 -12338
rect 1240 -12390 1244 -12338
rect -32 -12394 1244 -12390
rect -1776 -12440 -1288 -12434
rect -1776 -12474 -1729 -12440
rect -1695 -12474 -1657 -12440
rect -1623 -12474 -1585 -12440
rect -1551 -12474 -1513 -12440
rect -1479 -12474 -1441 -12440
rect -1407 -12474 -1369 -12440
rect -1335 -12474 -1288 -12440
rect -1776 -12480 -1288 -12474
rect -758 -12440 -270 -12434
rect -758 -12474 -711 -12440
rect -677 -12474 -639 -12440
rect -605 -12474 -567 -12440
rect -533 -12474 -495 -12440
rect -461 -12474 -423 -12440
rect -389 -12474 -351 -12440
rect -317 -12474 -270 -12440
rect -758 -12480 -270 -12474
rect -2072 -12560 -2058 -12543
rect -3082 -12615 -3036 -12577
rect -3082 -12649 -3076 -12615
rect -3042 -12649 -3036 -12615
rect -3082 -12687 -3036 -12649
rect -3082 -12721 -3076 -12687
rect -3042 -12721 -3036 -12687
rect -3082 -12759 -3036 -12721
rect -3082 -12793 -3076 -12759
rect -3042 -12793 -3036 -12759
rect -3082 -12831 -3036 -12793
rect -3082 -12865 -3076 -12831
rect -3042 -12865 -3036 -12831
rect -3082 -12903 -3036 -12865
rect -3082 -12937 -3076 -12903
rect -3042 -12937 -3036 -12903
rect -3082 -12975 -3036 -12937
rect -3082 -13009 -3076 -12975
rect -3042 -13009 -3036 -12975
rect -3082 -13047 -3036 -13009
rect -3082 -13080 -3076 -13047
rect -4060 -13081 -4050 -13080
rect -4830 -13150 -4342 -13144
rect -4830 -13184 -4783 -13150
rect -4749 -13184 -4711 -13150
rect -4677 -13184 -4639 -13150
rect -4605 -13184 -4567 -13150
rect -4533 -13184 -4495 -13150
rect -4461 -13184 -4423 -13150
rect -4389 -13184 -4342 -13150
rect -4830 -13190 -4342 -13184
rect -4620 -13252 -4560 -13190
rect -4830 -13258 -4342 -13252
rect -4830 -13292 -4783 -13258
rect -4749 -13292 -4711 -13258
rect -4677 -13292 -4639 -13258
rect -4605 -13292 -4567 -13258
rect -4533 -13292 -4495 -13258
rect -4461 -13292 -4423 -13258
rect -4389 -13292 -4342 -13258
rect -4830 -13298 -4342 -13292
rect -5122 -13362 -5112 -13361
rect -6096 -13395 -6090 -13370
rect -6136 -13433 -6090 -13395
rect -6136 -13467 -6130 -13433
rect -6096 -13467 -6090 -13433
rect -6136 -13505 -6090 -13467
rect -6136 -13539 -6130 -13505
rect -6096 -13539 -6090 -13505
rect -6136 -13577 -6090 -13539
rect -6136 -13611 -6130 -13577
rect -6096 -13611 -6090 -13577
rect -6136 -13649 -6090 -13611
rect -6136 -13683 -6130 -13649
rect -6096 -13683 -6090 -13649
rect -6136 -13721 -6090 -13683
rect -6136 -13755 -6130 -13721
rect -6096 -13755 -6090 -13721
rect -6136 -13793 -6090 -13755
rect -6136 -13827 -6130 -13793
rect -6096 -13827 -6090 -13793
rect -6136 -13865 -6090 -13827
rect -7114 -13899 -7098 -13890
rect -6136 -13894 -6130 -13865
rect -7884 -13968 -7396 -13962
rect -7884 -14002 -7837 -13968
rect -7803 -14002 -7765 -13968
rect -7731 -14002 -7693 -13968
rect -7659 -14002 -7621 -13968
rect -7587 -14002 -7549 -13968
rect -7515 -14002 -7477 -13968
rect -7443 -14002 -7396 -13968
rect -7884 -14008 -7396 -14002
rect -7670 -14070 -7610 -14008
rect -7884 -14076 -7396 -14070
rect -7884 -14110 -7837 -14076
rect -7803 -14110 -7765 -14076
rect -7731 -14110 -7693 -14076
rect -7659 -14110 -7621 -14076
rect -7587 -14110 -7549 -14076
rect -7515 -14110 -7477 -14076
rect -7443 -14110 -7396 -14076
rect -7884 -14116 -7396 -14110
rect -8178 -14182 -8166 -14179
rect -9150 -14213 -9144 -14186
rect -9190 -14251 -9144 -14213
rect -9190 -14285 -9184 -14251
rect -9150 -14285 -9144 -14251
rect -9190 -14323 -9144 -14285
rect -9190 -14357 -9184 -14323
rect -9150 -14357 -9144 -14323
rect -9190 -14395 -9144 -14357
rect -9190 -14429 -9184 -14395
rect -9150 -14429 -9144 -14395
rect -9190 -14467 -9144 -14429
rect -9190 -14501 -9184 -14467
rect -9150 -14501 -9144 -14467
rect -9190 -14539 -9144 -14501
rect -9190 -14573 -9184 -14539
rect -9150 -14573 -9144 -14539
rect -9190 -14611 -9144 -14573
rect -9190 -14645 -9184 -14611
rect -9150 -14645 -9144 -14611
rect -9190 -14683 -9144 -14645
rect -9190 -14717 -9184 -14683
rect -9150 -14717 -9144 -14683
rect -9190 -14724 -9144 -14717
rect -8172 -14213 -8166 -14182
rect -8132 -14182 -8118 -14179
rect -7158 -14179 -7098 -13899
rect -6140 -13899 -6130 -13894
rect -6096 -13894 -6090 -13865
rect -5118 -13395 -5112 -13362
rect -5078 -13362 -5062 -13361
rect -4110 -13361 -4050 -13081
rect -3088 -13081 -3076 -13080
rect -3042 -13080 -3036 -13047
rect -2064 -12577 -2058 -12560
rect -2024 -12560 -2012 -12543
rect -1046 -12543 -1000 -12512
rect -2024 -12577 -2018 -12560
rect -2064 -12615 -2018 -12577
rect -2064 -12649 -2058 -12615
rect -2024 -12649 -2018 -12615
rect -2064 -12687 -2018 -12649
rect -2064 -12721 -2058 -12687
rect -2024 -12721 -2018 -12687
rect -2064 -12759 -2018 -12721
rect -2064 -12793 -2058 -12759
rect -2024 -12793 -2018 -12759
rect -2064 -12831 -2018 -12793
rect -2064 -12865 -2058 -12831
rect -2024 -12865 -2018 -12831
rect -2064 -12903 -2018 -12865
rect -2064 -12937 -2058 -12903
rect -2024 -12937 -2018 -12903
rect -2064 -12975 -2018 -12937
rect -2064 -13009 -2058 -12975
rect -2024 -13009 -2018 -12975
rect -2064 -13047 -2018 -13009
rect -2064 -13080 -2058 -13047
rect -3042 -13081 -3028 -13080
rect -3812 -13150 -3324 -13144
rect -3812 -13184 -3765 -13150
rect -3731 -13184 -3693 -13150
rect -3659 -13184 -3621 -13150
rect -3587 -13184 -3549 -13150
rect -3515 -13184 -3477 -13150
rect -3443 -13184 -3405 -13150
rect -3371 -13184 -3324 -13150
rect -3812 -13190 -3324 -13184
rect -3604 -13252 -3544 -13190
rect -3812 -13258 -3324 -13252
rect -3812 -13292 -3765 -13258
rect -3731 -13292 -3693 -13258
rect -3659 -13292 -3621 -13258
rect -3587 -13292 -3549 -13258
rect -3515 -13292 -3477 -13258
rect -3443 -13292 -3405 -13258
rect -3371 -13292 -3324 -13258
rect -3812 -13298 -3324 -13292
rect -5078 -13395 -5072 -13362
rect -4110 -13370 -4094 -13361
rect -5118 -13433 -5072 -13395
rect -5118 -13467 -5112 -13433
rect -5078 -13467 -5072 -13433
rect -5118 -13505 -5072 -13467
rect -5118 -13539 -5112 -13505
rect -5078 -13539 -5072 -13505
rect -5118 -13577 -5072 -13539
rect -5118 -13611 -5112 -13577
rect -5078 -13611 -5072 -13577
rect -5118 -13649 -5072 -13611
rect -5118 -13683 -5112 -13649
rect -5078 -13683 -5072 -13649
rect -5118 -13721 -5072 -13683
rect -5118 -13755 -5112 -13721
rect -5078 -13755 -5072 -13721
rect -5118 -13793 -5072 -13755
rect -5118 -13827 -5112 -13793
rect -5078 -13827 -5072 -13793
rect -5118 -13865 -5072 -13827
rect -5118 -13886 -5112 -13865
rect -6096 -13899 -6080 -13894
rect -6866 -13968 -6378 -13962
rect -6866 -14002 -6819 -13968
rect -6785 -14002 -6747 -13968
rect -6713 -14002 -6675 -13968
rect -6641 -14002 -6603 -13968
rect -6569 -14002 -6531 -13968
rect -6497 -14002 -6459 -13968
rect -6425 -14002 -6378 -13968
rect -6866 -14008 -6378 -14002
rect -6652 -14070 -6592 -14008
rect -6866 -14076 -6378 -14070
rect -6866 -14110 -6819 -14076
rect -6785 -14110 -6747 -14076
rect -6713 -14110 -6675 -14076
rect -6641 -14110 -6603 -14076
rect -6569 -14110 -6531 -14076
rect -6497 -14110 -6459 -14076
rect -6425 -14110 -6378 -14076
rect -6866 -14116 -6378 -14110
rect -7158 -14180 -7148 -14179
rect -8132 -14213 -8126 -14182
rect -8172 -14251 -8126 -14213
rect -8172 -14285 -8166 -14251
rect -8132 -14285 -8126 -14251
rect -8172 -14323 -8126 -14285
rect -8172 -14357 -8166 -14323
rect -8132 -14357 -8126 -14323
rect -8172 -14395 -8126 -14357
rect -8172 -14429 -8166 -14395
rect -8132 -14429 -8126 -14395
rect -8172 -14467 -8126 -14429
rect -8172 -14501 -8166 -14467
rect -8132 -14501 -8126 -14467
rect -8172 -14539 -8126 -14501
rect -8172 -14573 -8166 -14539
rect -8132 -14573 -8126 -14539
rect -8172 -14611 -8126 -14573
rect -8172 -14645 -8166 -14611
rect -8132 -14645 -8126 -14611
rect -8172 -14683 -8126 -14645
rect -8172 -14717 -8166 -14683
rect -8132 -14717 -8126 -14683
rect -8172 -14720 -8126 -14717
rect -7154 -14213 -7148 -14180
rect -7114 -14180 -7098 -14179
rect -6140 -14179 -6080 -13899
rect -5120 -13899 -5112 -13886
rect -5078 -13886 -5072 -13865
rect -4100 -13395 -4094 -13370
rect -4060 -13370 -4050 -13361
rect -3088 -13361 -3028 -13081
rect -2068 -13081 -2058 -13080
rect -2024 -13080 -2018 -13047
rect -1046 -12577 -1040 -12543
rect -1006 -12577 -1000 -12543
rect -32 -12543 28 -12394
rect 1184 -12400 1244 -12394
rect 1844 -12452 1916 -12448
rect 1844 -12504 1854 -12452
rect 1906 -12504 1916 -12452
rect 1844 -12508 1916 -12504
rect -32 -12576 -22 -12543
rect -1046 -12615 -1000 -12577
rect -1046 -12649 -1040 -12615
rect -1006 -12649 -1000 -12615
rect -1046 -12687 -1000 -12649
rect -1046 -12721 -1040 -12687
rect -1006 -12721 -1000 -12687
rect -1046 -12759 -1000 -12721
rect -1046 -12793 -1040 -12759
rect -1006 -12793 -1000 -12759
rect -1046 -12831 -1000 -12793
rect -1046 -12865 -1040 -12831
rect -1006 -12865 -1000 -12831
rect -1046 -12903 -1000 -12865
rect -1046 -12937 -1040 -12903
rect -1006 -12937 -1000 -12903
rect -1046 -12975 -1000 -12937
rect -1046 -13009 -1040 -12975
rect -1006 -13009 -1000 -12975
rect -1046 -13047 -1000 -13009
rect -1046 -13076 -1040 -13047
rect -2024 -13081 -2008 -13080
rect -2794 -13150 -2306 -13144
rect -2794 -13184 -2747 -13150
rect -2713 -13184 -2675 -13150
rect -2641 -13184 -2603 -13150
rect -2569 -13184 -2531 -13150
rect -2497 -13184 -2459 -13150
rect -2425 -13184 -2387 -13150
rect -2353 -13184 -2306 -13150
rect -2794 -13190 -2306 -13184
rect -2582 -13252 -2522 -13190
rect -2794 -13258 -2306 -13252
rect -2794 -13292 -2747 -13258
rect -2713 -13292 -2675 -13258
rect -2641 -13292 -2603 -13258
rect -2569 -13292 -2531 -13258
rect -2497 -13292 -2459 -13258
rect -2425 -13292 -2387 -13258
rect -2353 -13292 -2306 -13258
rect -2794 -13298 -2306 -13292
rect -3088 -13370 -3076 -13361
rect -4060 -13395 -4054 -13370
rect -4100 -13433 -4054 -13395
rect -4100 -13467 -4094 -13433
rect -4060 -13467 -4054 -13433
rect -4100 -13505 -4054 -13467
rect -4100 -13539 -4094 -13505
rect -4060 -13539 -4054 -13505
rect -4100 -13577 -4054 -13539
rect -4100 -13611 -4094 -13577
rect -4060 -13611 -4054 -13577
rect -4100 -13649 -4054 -13611
rect -4100 -13683 -4094 -13649
rect -4060 -13683 -4054 -13649
rect -4100 -13721 -4054 -13683
rect -4100 -13755 -4094 -13721
rect -4060 -13755 -4054 -13721
rect -4100 -13793 -4054 -13755
rect -4100 -13827 -4094 -13793
rect -4060 -13827 -4054 -13793
rect -4100 -13865 -4054 -13827
rect -5078 -13899 -5060 -13886
rect -4100 -13894 -4094 -13865
rect -5848 -13968 -5360 -13962
rect -5848 -14002 -5801 -13968
rect -5767 -14002 -5729 -13968
rect -5695 -14002 -5657 -13968
rect -5623 -14002 -5585 -13968
rect -5551 -14002 -5513 -13968
rect -5479 -14002 -5441 -13968
rect -5407 -14002 -5360 -13968
rect -5848 -14008 -5360 -14002
rect -5650 -14070 -5590 -14008
rect -5848 -14076 -5360 -14070
rect -5848 -14110 -5801 -14076
rect -5767 -14110 -5729 -14076
rect -5695 -14110 -5657 -14076
rect -5623 -14110 -5585 -14076
rect -5551 -14110 -5513 -14076
rect -5479 -14110 -5441 -14076
rect -5407 -14110 -5360 -14076
rect -5848 -14116 -5360 -14110
rect -5120 -14176 -5060 -13899
rect -4108 -13899 -4094 -13894
rect -4060 -13894 -4054 -13865
rect -3082 -13395 -3076 -13370
rect -3042 -13370 -3028 -13361
rect -2068 -13361 -2008 -13081
rect -1052 -13081 -1040 -13076
rect -1006 -13076 -1000 -13047
rect -28 -12577 -22 -12576
rect 12 -12576 28 -12543
rect 12 -12577 18 -12576
rect -28 -12615 18 -12577
rect -28 -12649 -22 -12615
rect 12 -12649 18 -12615
rect -28 -12687 18 -12649
rect -28 -12721 -22 -12687
rect 12 -12721 18 -12687
rect -28 -12759 18 -12721
rect -28 -12793 -22 -12759
rect 12 -12793 18 -12759
rect -28 -12831 18 -12793
rect -28 -12865 -22 -12831
rect 12 -12865 18 -12831
rect -28 -12903 18 -12865
rect -28 -12937 -22 -12903
rect 12 -12937 18 -12903
rect -28 -12975 18 -12937
rect -28 -13009 -22 -12975
rect 12 -13009 18 -12975
rect -28 -13047 18 -13009
rect -1006 -13081 -992 -13076
rect -28 -13080 -22 -13047
rect -1776 -13150 -1288 -13144
rect -1776 -13184 -1729 -13150
rect -1695 -13184 -1657 -13150
rect -1623 -13184 -1585 -13150
rect -1551 -13184 -1513 -13150
rect -1479 -13184 -1441 -13150
rect -1407 -13184 -1369 -13150
rect -1335 -13184 -1288 -13150
rect -1776 -13190 -1288 -13184
rect -1570 -13252 -1510 -13190
rect -1776 -13258 -1288 -13252
rect -1776 -13292 -1729 -13258
rect -1695 -13292 -1657 -13258
rect -1623 -13292 -1585 -13258
rect -1551 -13292 -1513 -13258
rect -1479 -13292 -1441 -13258
rect -1407 -13292 -1369 -13258
rect -1335 -13292 -1288 -13258
rect -1776 -13298 -1288 -13292
rect -2068 -13370 -2058 -13361
rect -3042 -13395 -3036 -13370
rect -3082 -13433 -3036 -13395
rect -3082 -13467 -3076 -13433
rect -3042 -13467 -3036 -13433
rect -3082 -13505 -3036 -13467
rect -3082 -13539 -3076 -13505
rect -3042 -13539 -3036 -13505
rect -3082 -13577 -3036 -13539
rect -3082 -13611 -3076 -13577
rect -3042 -13611 -3036 -13577
rect -3082 -13649 -3036 -13611
rect -3082 -13683 -3076 -13649
rect -3042 -13683 -3036 -13649
rect -3082 -13721 -3036 -13683
rect -3082 -13755 -3076 -13721
rect -3042 -13755 -3036 -13721
rect -3082 -13793 -3036 -13755
rect -3082 -13827 -3076 -13793
rect -3042 -13827 -3036 -13793
rect -3082 -13865 -3036 -13827
rect -3082 -13894 -3076 -13865
rect -4060 -13899 -4048 -13894
rect -4830 -13968 -4342 -13962
rect -4830 -14002 -4783 -13968
rect -4749 -14002 -4711 -13968
rect -4677 -14002 -4639 -13968
rect -4605 -14002 -4567 -13968
rect -4533 -14002 -4495 -13968
rect -4461 -14002 -4423 -13968
rect -4389 -14002 -4342 -13968
rect -4830 -14008 -4342 -14002
rect -4620 -14070 -4560 -14008
rect -4830 -14076 -4342 -14070
rect -4830 -14110 -4783 -14076
rect -4749 -14110 -4711 -14076
rect -4677 -14110 -4639 -14076
rect -4605 -14110 -4567 -14076
rect -4533 -14110 -4495 -14076
rect -4461 -14110 -4423 -14076
rect -4389 -14110 -4342 -14076
rect -4830 -14116 -4342 -14110
rect -7114 -14213 -7108 -14180
rect -6140 -14184 -6130 -14179
rect -7154 -14251 -7108 -14213
rect -7154 -14285 -7148 -14251
rect -7114 -14285 -7108 -14251
rect -7154 -14323 -7108 -14285
rect -7154 -14357 -7148 -14323
rect -7114 -14357 -7108 -14323
rect -7154 -14395 -7108 -14357
rect -7154 -14429 -7148 -14395
rect -7114 -14429 -7108 -14395
rect -7154 -14467 -7108 -14429
rect -7154 -14501 -7148 -14467
rect -7114 -14501 -7108 -14467
rect -7154 -14539 -7108 -14501
rect -7154 -14573 -7148 -14539
rect -7114 -14573 -7108 -14539
rect -7154 -14611 -7108 -14573
rect -7154 -14645 -7148 -14611
rect -7114 -14645 -7108 -14611
rect -7154 -14683 -7108 -14645
rect -7154 -14717 -7148 -14683
rect -7114 -14717 -7108 -14683
rect -7154 -14718 -7108 -14717
rect -6136 -14213 -6130 -14184
rect -6096 -14184 -6080 -14179
rect -5118 -14179 -5072 -14176
rect -6096 -14213 -6090 -14184
rect -6136 -14251 -6090 -14213
rect -6136 -14285 -6130 -14251
rect -6096 -14285 -6090 -14251
rect -6136 -14323 -6090 -14285
rect -6136 -14357 -6130 -14323
rect -6096 -14357 -6090 -14323
rect -6136 -14395 -6090 -14357
rect -6136 -14429 -6130 -14395
rect -6096 -14429 -6090 -14395
rect -6136 -14467 -6090 -14429
rect -6136 -14501 -6130 -14467
rect -6096 -14501 -6090 -14467
rect -6136 -14539 -6090 -14501
rect -6136 -14573 -6130 -14539
rect -6096 -14573 -6090 -14539
rect -6136 -14611 -6090 -14573
rect -6136 -14645 -6130 -14611
rect -6096 -14645 -6090 -14611
rect -6136 -14683 -6090 -14645
rect -6136 -14717 -6130 -14683
rect -6096 -14717 -6090 -14683
rect -5118 -14213 -5112 -14179
rect -5078 -14213 -5072 -14179
rect -4108 -14179 -4048 -13899
rect -3086 -13899 -3076 -13894
rect -3042 -13894 -3036 -13865
rect -2064 -13395 -2058 -13370
rect -2024 -13370 -2008 -13361
rect -1052 -13361 -992 -13081
rect -30 -13081 -22 -13080
rect 12 -13080 18 -13047
rect 12 -13081 30 -13080
rect -758 -13150 -270 -13144
rect -758 -13184 -711 -13150
rect -677 -13184 -639 -13150
rect -605 -13184 -567 -13150
rect -533 -13184 -495 -13150
rect -461 -13184 -423 -13150
rect -389 -13184 -351 -13150
rect -317 -13184 -270 -13150
rect -758 -13190 -270 -13184
rect -550 -13252 -490 -13190
rect -758 -13258 -270 -13252
rect -758 -13292 -711 -13258
rect -677 -13292 -639 -13258
rect -605 -13292 -567 -13258
rect -533 -13292 -495 -13258
rect -461 -13292 -423 -13258
rect -389 -13292 -351 -13258
rect -317 -13292 -270 -13258
rect -758 -13298 -270 -13292
rect -1052 -13366 -1040 -13361
rect -2024 -13395 -2018 -13370
rect -2064 -13433 -2018 -13395
rect -2064 -13467 -2058 -13433
rect -2024 -13467 -2018 -13433
rect -2064 -13505 -2018 -13467
rect -2064 -13539 -2058 -13505
rect -2024 -13539 -2018 -13505
rect -2064 -13577 -2018 -13539
rect -2064 -13611 -2058 -13577
rect -2024 -13611 -2018 -13577
rect -2064 -13649 -2018 -13611
rect -2064 -13683 -2058 -13649
rect -2024 -13683 -2018 -13649
rect -2064 -13721 -2018 -13683
rect -2064 -13755 -2058 -13721
rect -2024 -13755 -2018 -13721
rect -2064 -13793 -2018 -13755
rect -2064 -13827 -2058 -13793
rect -2024 -13827 -2018 -13793
rect -2064 -13865 -2018 -13827
rect -2064 -13894 -2058 -13865
rect -3042 -13899 -3026 -13894
rect -3812 -13968 -3324 -13962
rect -3812 -14002 -3765 -13968
rect -3731 -14002 -3693 -13968
rect -3659 -14002 -3621 -13968
rect -3587 -14002 -3549 -13968
rect -3515 -14002 -3477 -13968
rect -3443 -14002 -3405 -13968
rect -3371 -14002 -3324 -13968
rect -3812 -14008 -3324 -14002
rect -3604 -14070 -3544 -14008
rect -3812 -14076 -3324 -14070
rect -3812 -14110 -3765 -14076
rect -3731 -14110 -3693 -14076
rect -3659 -14110 -3621 -14076
rect -3587 -14110 -3549 -14076
rect -3515 -14110 -3477 -14076
rect -3443 -14110 -3405 -14076
rect -3371 -14110 -3324 -14076
rect -3812 -14116 -3324 -14110
rect -4108 -14184 -4094 -14179
rect -5118 -14251 -5072 -14213
rect -5118 -14285 -5112 -14251
rect -5078 -14285 -5072 -14251
rect -5118 -14323 -5072 -14285
rect -5118 -14357 -5112 -14323
rect -5078 -14357 -5072 -14323
rect -5118 -14395 -5072 -14357
rect -5118 -14429 -5112 -14395
rect -5078 -14429 -5072 -14395
rect -5118 -14467 -5072 -14429
rect -5118 -14501 -5112 -14467
rect -5078 -14501 -5072 -14467
rect -5118 -14539 -5072 -14501
rect -5118 -14573 -5112 -14539
rect -5078 -14573 -5072 -14539
rect -5118 -14611 -5072 -14573
rect -5118 -14645 -5112 -14611
rect -5078 -14645 -5072 -14611
rect -5118 -14683 -5072 -14645
rect -5118 -14714 -5112 -14683
rect -12328 -14789 -12289 -14755
rect -12255 -14789 -12216 -14755
rect -12328 -14827 -12216 -14789
rect -12328 -14861 -12289 -14827
rect -12255 -14861 -12216 -14827
rect -12328 -14899 -12216 -14861
rect -12328 -14933 -12289 -14899
rect -12255 -14933 -12216 -14899
rect -12328 -14971 -12216 -14933
rect -12328 -15005 -12289 -14971
rect -12255 -15005 -12216 -14971
rect -12328 -15043 -12216 -15005
rect -9198 -14997 -9138 -14724
rect -8902 -14786 -8414 -14780
rect -8902 -14820 -8855 -14786
rect -8821 -14820 -8783 -14786
rect -8749 -14820 -8711 -14786
rect -8677 -14820 -8639 -14786
rect -8605 -14820 -8567 -14786
rect -8533 -14820 -8495 -14786
rect -8461 -14820 -8414 -14786
rect -8902 -14826 -8414 -14820
rect -8692 -14888 -8632 -14826
rect -8902 -14894 -8414 -14888
rect -8902 -14928 -8855 -14894
rect -8821 -14928 -8783 -14894
rect -8749 -14928 -8711 -14894
rect -8677 -14928 -8639 -14894
rect -8605 -14928 -8567 -14894
rect -8533 -14928 -8495 -14894
rect -8461 -14928 -8414 -14894
rect -8902 -14934 -8414 -14928
rect -9198 -15014 -9184 -14997
rect -12328 -15077 -12289 -15043
rect -12255 -15077 -12216 -15043
rect -12328 -15115 -12216 -15077
rect -12328 -15149 -12289 -15115
rect -12255 -15149 -12216 -15115
rect -12328 -15187 -12216 -15149
rect -12328 -15221 -12289 -15187
rect -12255 -15221 -12216 -15187
rect -12328 -15259 -12216 -15221
rect -12328 -15293 -12289 -15259
rect -12255 -15293 -12216 -15259
rect -12328 -15331 -12216 -15293
rect -12328 -15365 -12289 -15331
rect -12255 -15365 -12216 -15331
rect -12328 -15403 -12216 -15365
rect -12328 -15437 -12289 -15403
rect -12255 -15437 -12216 -15403
rect -12328 -15475 -12216 -15437
rect -12328 -15509 -12289 -15475
rect -12255 -15509 -12216 -15475
rect -12328 -15547 -12216 -15509
rect -9190 -15031 -9184 -15014
rect -9150 -15014 -9138 -14997
rect -8178 -14997 -8118 -14720
rect -7884 -14786 -7396 -14780
rect -7884 -14820 -7837 -14786
rect -7803 -14820 -7765 -14786
rect -7731 -14820 -7693 -14786
rect -7659 -14820 -7621 -14786
rect -7587 -14820 -7549 -14786
rect -7515 -14820 -7477 -14786
rect -7443 -14820 -7396 -14786
rect -7884 -14826 -7396 -14820
rect -7670 -14888 -7610 -14826
rect -7884 -14894 -7396 -14888
rect -7884 -14928 -7837 -14894
rect -7803 -14928 -7765 -14894
rect -7731 -14928 -7693 -14894
rect -7659 -14928 -7621 -14894
rect -7587 -14928 -7549 -14894
rect -7515 -14928 -7477 -14894
rect -7443 -14928 -7396 -14894
rect -7884 -14934 -7396 -14928
rect -8178 -15010 -8166 -14997
rect -9150 -15031 -9144 -15014
rect -9190 -15069 -9144 -15031
rect -9190 -15103 -9184 -15069
rect -9150 -15103 -9144 -15069
rect -9190 -15141 -9144 -15103
rect -9190 -15175 -9184 -15141
rect -9150 -15175 -9144 -15141
rect -9190 -15213 -9144 -15175
rect -9190 -15247 -9184 -15213
rect -9150 -15247 -9144 -15213
rect -9190 -15285 -9144 -15247
rect -9190 -15319 -9184 -15285
rect -9150 -15319 -9144 -15285
rect -9190 -15357 -9144 -15319
rect -9190 -15391 -9184 -15357
rect -9150 -15391 -9144 -15357
rect -9190 -15429 -9144 -15391
rect -9190 -15463 -9184 -15429
rect -9150 -15463 -9144 -15429
rect -9190 -15501 -9144 -15463
rect -9190 -15535 -9184 -15501
rect -9150 -15535 -9144 -15501
rect -8172 -15031 -8166 -15010
rect -8132 -15010 -8118 -14997
rect -7158 -14997 -7098 -14718
rect -6136 -14722 -6090 -14717
rect -5120 -14717 -5112 -14714
rect -5078 -14714 -5072 -14683
rect -4100 -14213 -4094 -14184
rect -4060 -14184 -4048 -14179
rect -3086 -14179 -3026 -13899
rect -2066 -13899 -2058 -13894
rect -2024 -13894 -2018 -13865
rect -1046 -13395 -1040 -13366
rect -1006 -13366 -992 -13361
rect -30 -13361 30 -13081
rect -1006 -13395 -1000 -13366
rect -30 -13370 -22 -13361
rect -1046 -13433 -1000 -13395
rect -1046 -13467 -1040 -13433
rect -1006 -13467 -1000 -13433
rect -1046 -13505 -1000 -13467
rect -1046 -13539 -1040 -13505
rect -1006 -13539 -1000 -13505
rect -1046 -13577 -1000 -13539
rect -1046 -13611 -1040 -13577
rect -1006 -13611 -1000 -13577
rect -1046 -13649 -1000 -13611
rect -1046 -13683 -1040 -13649
rect -1006 -13683 -1000 -13649
rect -1046 -13721 -1000 -13683
rect -1046 -13755 -1040 -13721
rect -1006 -13755 -1000 -13721
rect -1046 -13793 -1000 -13755
rect -1046 -13827 -1040 -13793
rect -1006 -13827 -1000 -13793
rect -1046 -13865 -1000 -13827
rect -1046 -13890 -1040 -13865
rect -2024 -13899 -2006 -13894
rect -2794 -13968 -2306 -13962
rect -2794 -14002 -2747 -13968
rect -2713 -14002 -2675 -13968
rect -2641 -14002 -2603 -13968
rect -2569 -14002 -2531 -13968
rect -2497 -14002 -2459 -13968
rect -2425 -14002 -2387 -13968
rect -2353 -14002 -2306 -13968
rect -2794 -14008 -2306 -14002
rect -2582 -14070 -2522 -14008
rect -2794 -14076 -2306 -14070
rect -2794 -14110 -2747 -14076
rect -2713 -14110 -2675 -14076
rect -2641 -14110 -2603 -14076
rect -2569 -14110 -2531 -14076
rect -2497 -14110 -2459 -14076
rect -2425 -14110 -2387 -14076
rect -2353 -14110 -2306 -14076
rect -2794 -14116 -2306 -14110
rect -3086 -14184 -3076 -14179
rect -4060 -14213 -4054 -14184
rect -4100 -14251 -4054 -14213
rect -4100 -14285 -4094 -14251
rect -4060 -14285 -4054 -14251
rect -4100 -14323 -4054 -14285
rect -4100 -14357 -4094 -14323
rect -4060 -14357 -4054 -14323
rect -4100 -14395 -4054 -14357
rect -4100 -14429 -4094 -14395
rect -4060 -14429 -4054 -14395
rect -4100 -14467 -4054 -14429
rect -4100 -14501 -4094 -14467
rect -4060 -14501 -4054 -14467
rect -4100 -14539 -4054 -14501
rect -4100 -14573 -4094 -14539
rect -4060 -14573 -4054 -14539
rect -4100 -14611 -4054 -14573
rect -4100 -14645 -4094 -14611
rect -4060 -14645 -4054 -14611
rect -4100 -14683 -4054 -14645
rect -5078 -14717 -5060 -14714
rect -6866 -14786 -6378 -14780
rect -6866 -14820 -6819 -14786
rect -6785 -14820 -6747 -14786
rect -6713 -14820 -6675 -14786
rect -6641 -14820 -6603 -14786
rect -6569 -14820 -6531 -14786
rect -6497 -14820 -6459 -14786
rect -6425 -14820 -6378 -14786
rect -6866 -14826 -6378 -14820
rect -6658 -14888 -6598 -14826
rect -6866 -14894 -6378 -14888
rect -6866 -14928 -6819 -14894
rect -6785 -14928 -6747 -14894
rect -6713 -14928 -6675 -14894
rect -6641 -14928 -6603 -14894
rect -6569 -14928 -6531 -14894
rect -6497 -14928 -6459 -14894
rect -6425 -14928 -6378 -14894
rect -6866 -14934 -6378 -14928
rect -7158 -15008 -7148 -14997
rect -8132 -15031 -8126 -15010
rect -8172 -15069 -8126 -15031
rect -8172 -15103 -8166 -15069
rect -8132 -15103 -8126 -15069
rect -8172 -15141 -8126 -15103
rect -8172 -15175 -8166 -15141
rect -8132 -15175 -8126 -15141
rect -8172 -15213 -8126 -15175
rect -8172 -15247 -8166 -15213
rect -8132 -15247 -8126 -15213
rect -8172 -15285 -8126 -15247
rect -8172 -15319 -8166 -15285
rect -8132 -15319 -8126 -15285
rect -8172 -15357 -8126 -15319
rect -8172 -15391 -8166 -15357
rect -8132 -15391 -8126 -15357
rect -8172 -15429 -8126 -15391
rect -8172 -15463 -8166 -15429
rect -8132 -15463 -8126 -15429
rect -8172 -15501 -8126 -15463
rect -8172 -15532 -8166 -15501
rect -9190 -15536 -9144 -15535
rect -8178 -15535 -8166 -15532
rect -8132 -15532 -8126 -15501
rect -7154 -15031 -7148 -15008
rect -7114 -15008 -7098 -14997
rect -6140 -14997 -6080 -14722
rect -5848 -14786 -5360 -14780
rect -5848 -14820 -5801 -14786
rect -5767 -14820 -5729 -14786
rect -5695 -14820 -5657 -14786
rect -5623 -14820 -5585 -14786
rect -5551 -14820 -5513 -14786
rect -5479 -14820 -5441 -14786
rect -5407 -14820 -5360 -14786
rect -5848 -14826 -5360 -14820
rect -5656 -14888 -5596 -14826
rect -5848 -14894 -5360 -14888
rect -5848 -14928 -5801 -14894
rect -5767 -14928 -5729 -14894
rect -5695 -14928 -5657 -14894
rect -5623 -14928 -5585 -14894
rect -5551 -14928 -5513 -14894
rect -5479 -14928 -5441 -14894
rect -5407 -14928 -5360 -14894
rect -5848 -14934 -5360 -14928
rect -7114 -15031 -7108 -15008
rect -6140 -15012 -6130 -14997
rect -7154 -15069 -7108 -15031
rect -7154 -15103 -7148 -15069
rect -7114 -15103 -7108 -15069
rect -7154 -15141 -7108 -15103
rect -7154 -15175 -7148 -15141
rect -7114 -15175 -7108 -15141
rect -7154 -15213 -7108 -15175
rect -7154 -15247 -7148 -15213
rect -7114 -15247 -7108 -15213
rect -7154 -15285 -7108 -15247
rect -7154 -15319 -7148 -15285
rect -7114 -15319 -7108 -15285
rect -7154 -15357 -7108 -15319
rect -7154 -15391 -7148 -15357
rect -7114 -15391 -7108 -15357
rect -7154 -15429 -7108 -15391
rect -7154 -15463 -7148 -15429
rect -7114 -15463 -7108 -15429
rect -7154 -15501 -7108 -15463
rect -7154 -15530 -7148 -15501
rect -8132 -15535 -8118 -15532
rect -12328 -15581 -12289 -15547
rect -12255 -15581 -12216 -15547
rect -12328 -15619 -12216 -15581
rect -12328 -15653 -12289 -15619
rect -12255 -15653 -12216 -15619
rect -12328 -15691 -12216 -15653
rect -12328 -15725 -12289 -15691
rect -12255 -15725 -12216 -15691
rect -12328 -15763 -12216 -15725
rect -12328 -15797 -12289 -15763
rect -12255 -15797 -12216 -15763
rect -12328 -15835 -12216 -15797
rect -9198 -15815 -9138 -15536
rect -8902 -15604 -8414 -15598
rect -8902 -15638 -8855 -15604
rect -8821 -15638 -8783 -15604
rect -8749 -15638 -8711 -15604
rect -8677 -15638 -8639 -15604
rect -8605 -15638 -8567 -15604
rect -8533 -15638 -8495 -15604
rect -8461 -15638 -8414 -15604
rect -8902 -15644 -8414 -15638
rect -8694 -15706 -8634 -15644
rect -8902 -15712 -8414 -15706
rect -8902 -15746 -8855 -15712
rect -8821 -15746 -8783 -15712
rect -8749 -15746 -8711 -15712
rect -8677 -15746 -8639 -15712
rect -8605 -15746 -8567 -15712
rect -8533 -15746 -8495 -15712
rect -8461 -15746 -8414 -15712
rect -8902 -15752 -8414 -15746
rect -9198 -15826 -9184 -15815
rect -12328 -15869 -12289 -15835
rect -12255 -15869 -12216 -15835
rect -12328 -15907 -12216 -15869
rect -12328 -15941 -12289 -15907
rect -12255 -15941 -12216 -15907
rect -12328 -15979 -12216 -15941
rect -12328 -16013 -12289 -15979
rect -12255 -16013 -12216 -15979
rect -12328 -16051 -12216 -16013
rect -12328 -16085 -12289 -16051
rect -12255 -16085 -12216 -16051
rect -12328 -16123 -12216 -16085
rect -12328 -16157 -12289 -16123
rect -12255 -16157 -12216 -16123
rect -12328 -16195 -12216 -16157
rect -12328 -16229 -12289 -16195
rect -12255 -16229 -12216 -16195
rect -12328 -16267 -12216 -16229
rect -12328 -16301 -12289 -16267
rect -12255 -16301 -12216 -16267
rect -12328 -16339 -12216 -16301
rect -12328 -16373 -12289 -16339
rect -12255 -16373 -12216 -16339
rect -9190 -15849 -9184 -15826
rect -9150 -15826 -9138 -15815
rect -8178 -15815 -8118 -15535
rect -7158 -15535 -7148 -15530
rect -7114 -15530 -7108 -15501
rect -6136 -15031 -6130 -15012
rect -6096 -15012 -6080 -14997
rect -5120 -14997 -5060 -14717
rect -4100 -14717 -4094 -14683
rect -4060 -14717 -4054 -14683
rect -4100 -14722 -4054 -14717
rect -3082 -14213 -3076 -14184
rect -3042 -14184 -3026 -14179
rect -2066 -14179 -2006 -13899
rect -1050 -13899 -1040 -13890
rect -1006 -13890 -1000 -13865
rect -28 -13395 -22 -13370
rect 12 -13370 30 -13361
rect 12 -13395 18 -13370
rect -28 -13433 18 -13395
rect -28 -13467 -22 -13433
rect 12 -13467 18 -13433
rect -28 -13505 18 -13467
rect -28 -13539 -22 -13505
rect 12 -13539 18 -13505
rect -28 -13577 18 -13539
rect -28 -13611 -22 -13577
rect 12 -13611 18 -13577
rect -28 -13649 18 -13611
rect -28 -13683 -22 -13649
rect 12 -13683 18 -13649
rect -28 -13721 18 -13683
rect -28 -13755 -22 -13721
rect 12 -13755 18 -13721
rect -28 -13793 18 -13755
rect -28 -13827 -22 -13793
rect 12 -13827 18 -13793
rect -28 -13865 18 -13827
rect -1006 -13899 -990 -13890
rect -1776 -13968 -1288 -13962
rect -1776 -14002 -1729 -13968
rect -1695 -14002 -1657 -13968
rect -1623 -14002 -1585 -13968
rect -1551 -14002 -1513 -13968
rect -1479 -14002 -1441 -13968
rect -1407 -14002 -1369 -13968
rect -1335 -14002 -1288 -13968
rect -1776 -14008 -1288 -14002
rect -1570 -14070 -1510 -14008
rect -1776 -14076 -1288 -14070
rect -1776 -14110 -1729 -14076
rect -1695 -14110 -1657 -14076
rect -1623 -14110 -1585 -14076
rect -1551 -14110 -1513 -14076
rect -1479 -14110 -1441 -14076
rect -1407 -14110 -1369 -14076
rect -1335 -14110 -1288 -14076
rect -1776 -14116 -1288 -14110
rect -2066 -14184 -2058 -14179
rect -3042 -14213 -3036 -14184
rect -3082 -14251 -3036 -14213
rect -3082 -14285 -3076 -14251
rect -3042 -14285 -3036 -14251
rect -3082 -14323 -3036 -14285
rect -3082 -14357 -3076 -14323
rect -3042 -14357 -3036 -14323
rect -3082 -14395 -3036 -14357
rect -3082 -14429 -3076 -14395
rect -3042 -14429 -3036 -14395
rect -3082 -14467 -3036 -14429
rect -3082 -14501 -3076 -14467
rect -3042 -14501 -3036 -14467
rect -3082 -14539 -3036 -14501
rect -3082 -14573 -3076 -14539
rect -3042 -14573 -3036 -14539
rect -3082 -14611 -3036 -14573
rect -3082 -14645 -3076 -14611
rect -3042 -14645 -3036 -14611
rect -3082 -14683 -3036 -14645
rect -3082 -14717 -3076 -14683
rect -3042 -14717 -3036 -14683
rect -3082 -14722 -3036 -14717
rect -2064 -14213 -2058 -14184
rect -2024 -14184 -2006 -14179
rect -1050 -14179 -990 -13899
rect -28 -13899 -22 -13865
rect 12 -13894 18 -13865
rect 12 -13899 32 -13894
rect -758 -13968 -270 -13962
rect -758 -14002 -711 -13968
rect -677 -14002 -639 -13968
rect -605 -14002 -567 -13968
rect -533 -14002 -495 -13968
rect -461 -14002 -423 -13968
rect -389 -14002 -351 -13968
rect -317 -14002 -270 -13968
rect -758 -14008 -270 -14002
rect -550 -14070 -490 -14008
rect -758 -14076 -270 -14070
rect -758 -14110 -711 -14076
rect -677 -14110 -639 -14076
rect -605 -14110 -567 -14076
rect -533 -14110 -495 -14076
rect -461 -14110 -423 -14076
rect -389 -14110 -351 -14076
rect -317 -14110 -270 -14076
rect -758 -14116 -270 -14110
rect -1050 -14180 -1040 -14179
rect -2024 -14213 -2018 -14184
rect -2064 -14251 -2018 -14213
rect -2064 -14285 -2058 -14251
rect -2024 -14285 -2018 -14251
rect -2064 -14323 -2018 -14285
rect -2064 -14357 -2058 -14323
rect -2024 -14357 -2018 -14323
rect -2064 -14395 -2018 -14357
rect -2064 -14429 -2058 -14395
rect -2024 -14429 -2018 -14395
rect -2064 -14467 -2018 -14429
rect -2064 -14501 -2058 -14467
rect -2024 -14501 -2018 -14467
rect -2064 -14539 -2018 -14501
rect -2064 -14573 -2058 -14539
rect -2024 -14573 -2018 -14539
rect -2064 -14611 -2018 -14573
rect -2064 -14645 -2058 -14611
rect -2024 -14645 -2018 -14611
rect -2064 -14683 -2018 -14645
rect -2064 -14717 -2058 -14683
rect -2024 -14717 -2018 -14683
rect -2064 -14722 -2018 -14717
rect -1046 -14213 -1040 -14180
rect -1006 -14180 -990 -14179
rect -28 -14179 32 -13899
rect -1006 -14213 -1000 -14180
rect -1046 -14251 -1000 -14213
rect -1046 -14285 -1040 -14251
rect -1006 -14285 -1000 -14251
rect -1046 -14323 -1000 -14285
rect -1046 -14357 -1040 -14323
rect -1006 -14357 -1000 -14323
rect -1046 -14395 -1000 -14357
rect -1046 -14429 -1040 -14395
rect -1006 -14429 -1000 -14395
rect -1046 -14467 -1000 -14429
rect -1046 -14501 -1040 -14467
rect -1006 -14501 -1000 -14467
rect -1046 -14539 -1000 -14501
rect -1046 -14573 -1040 -14539
rect -1006 -14573 -1000 -14539
rect -1046 -14611 -1000 -14573
rect -1046 -14645 -1040 -14611
rect -1006 -14645 -1000 -14611
rect -1046 -14683 -1000 -14645
rect -1046 -14717 -1040 -14683
rect -1006 -14717 -1000 -14683
rect -1046 -14718 -1000 -14717
rect -28 -14213 -22 -14179
rect 12 -14184 32 -14179
rect 12 -14213 18 -14184
rect -28 -14251 18 -14213
rect -28 -14285 -22 -14251
rect 12 -14285 18 -14251
rect -28 -14323 18 -14285
rect -28 -14357 -22 -14323
rect 12 -14357 18 -14323
rect -28 -14395 18 -14357
rect -28 -14429 -22 -14395
rect 12 -14429 18 -14395
rect -28 -14467 18 -14429
rect -28 -14501 -22 -14467
rect 12 -14501 18 -14467
rect -28 -14539 18 -14501
rect -28 -14573 -22 -14539
rect 12 -14573 18 -14539
rect -28 -14611 18 -14573
rect -28 -14645 -22 -14611
rect 12 -14645 18 -14611
rect -28 -14683 18 -14645
rect -28 -14717 -22 -14683
rect 12 -14717 18 -14683
rect -4830 -14786 -4342 -14780
rect -4830 -14820 -4783 -14786
rect -4749 -14820 -4711 -14786
rect -4677 -14820 -4639 -14786
rect -4605 -14820 -4567 -14786
rect -4533 -14820 -4495 -14786
rect -4461 -14820 -4423 -14786
rect -4389 -14820 -4342 -14786
rect -4830 -14826 -4342 -14820
rect -4626 -14888 -4566 -14826
rect -4830 -14894 -4342 -14888
rect -4830 -14928 -4783 -14894
rect -4749 -14928 -4711 -14894
rect -4677 -14928 -4639 -14894
rect -4605 -14928 -4567 -14894
rect -4533 -14928 -4495 -14894
rect -4461 -14928 -4423 -14894
rect -4389 -14928 -4342 -14894
rect -4830 -14934 -4342 -14928
rect -5120 -15004 -5112 -14997
rect -6096 -15031 -6090 -15012
rect -6136 -15069 -6090 -15031
rect -6136 -15103 -6130 -15069
rect -6096 -15103 -6090 -15069
rect -6136 -15141 -6090 -15103
rect -6136 -15175 -6130 -15141
rect -6096 -15175 -6090 -15141
rect -6136 -15213 -6090 -15175
rect -6136 -15247 -6130 -15213
rect -6096 -15247 -6090 -15213
rect -6136 -15285 -6090 -15247
rect -6136 -15319 -6130 -15285
rect -6096 -15319 -6090 -15285
rect -6136 -15357 -6090 -15319
rect -6136 -15391 -6130 -15357
rect -6096 -15391 -6090 -15357
rect -6136 -15429 -6090 -15391
rect -6136 -15463 -6130 -15429
rect -6096 -15463 -6090 -15429
rect -6136 -15501 -6090 -15463
rect -7114 -15535 -7098 -15530
rect -6136 -15534 -6130 -15501
rect -7884 -15604 -7396 -15598
rect -7884 -15638 -7837 -15604
rect -7803 -15638 -7765 -15604
rect -7731 -15638 -7693 -15604
rect -7659 -15638 -7621 -15604
rect -7587 -15638 -7549 -15604
rect -7515 -15638 -7477 -15604
rect -7443 -15638 -7396 -15604
rect -7884 -15644 -7396 -15638
rect -7676 -15706 -7616 -15644
rect -7884 -15712 -7396 -15706
rect -7884 -15746 -7837 -15712
rect -7803 -15746 -7765 -15712
rect -7731 -15746 -7693 -15712
rect -7659 -15746 -7621 -15712
rect -7587 -15746 -7549 -15712
rect -7515 -15746 -7477 -15712
rect -7443 -15746 -7396 -15712
rect -7884 -15752 -7396 -15746
rect -8178 -15822 -8166 -15815
rect -9150 -15849 -9144 -15826
rect -9190 -15887 -9144 -15849
rect -9190 -15921 -9184 -15887
rect -9150 -15921 -9144 -15887
rect -9190 -15959 -9144 -15921
rect -9190 -15993 -9184 -15959
rect -9150 -15993 -9144 -15959
rect -9190 -16031 -9144 -15993
rect -9190 -16065 -9184 -16031
rect -9150 -16065 -9144 -16031
rect -9190 -16103 -9144 -16065
rect -9190 -16137 -9184 -16103
rect -9150 -16137 -9144 -16103
rect -9190 -16175 -9144 -16137
rect -9190 -16209 -9184 -16175
rect -9150 -16209 -9144 -16175
rect -9190 -16247 -9144 -16209
rect -9190 -16281 -9184 -16247
rect -9150 -16281 -9144 -16247
rect -9190 -16319 -9144 -16281
rect -9190 -16353 -9184 -16319
rect -9150 -16353 -9144 -16319
rect -8172 -15849 -8166 -15822
rect -8132 -15822 -8118 -15815
rect -7158 -15815 -7098 -15535
rect -6140 -15535 -6130 -15534
rect -6096 -15534 -6090 -15501
rect -5118 -15031 -5112 -15004
rect -5078 -15004 -5060 -14997
rect -4108 -14997 -4048 -14722
rect -3812 -14786 -3324 -14780
rect -3812 -14820 -3765 -14786
rect -3731 -14820 -3693 -14786
rect -3659 -14820 -3621 -14786
rect -3587 -14820 -3549 -14786
rect -3515 -14820 -3477 -14786
rect -3443 -14820 -3405 -14786
rect -3371 -14820 -3324 -14786
rect -3812 -14826 -3324 -14820
rect -3610 -14888 -3550 -14826
rect -3812 -14894 -3324 -14888
rect -3812 -14928 -3765 -14894
rect -3731 -14928 -3693 -14894
rect -3659 -14928 -3621 -14894
rect -3587 -14928 -3549 -14894
rect -3515 -14928 -3477 -14894
rect -3443 -14928 -3405 -14894
rect -3371 -14928 -3324 -14894
rect -3812 -14934 -3324 -14928
rect -5078 -15031 -5072 -15004
rect -4108 -15012 -4094 -14997
rect -5118 -15069 -5072 -15031
rect -5118 -15103 -5112 -15069
rect -5078 -15103 -5072 -15069
rect -5118 -15141 -5072 -15103
rect -5118 -15175 -5112 -15141
rect -5078 -15175 -5072 -15141
rect -5118 -15213 -5072 -15175
rect -5118 -15247 -5112 -15213
rect -5078 -15247 -5072 -15213
rect -5118 -15285 -5072 -15247
rect -5118 -15319 -5112 -15285
rect -5078 -15319 -5072 -15285
rect -5118 -15357 -5072 -15319
rect -5118 -15391 -5112 -15357
rect -5078 -15391 -5072 -15357
rect -5118 -15429 -5072 -15391
rect -5118 -15463 -5112 -15429
rect -5078 -15463 -5072 -15429
rect -5118 -15501 -5072 -15463
rect -5118 -15526 -5112 -15501
rect -6096 -15535 -6080 -15534
rect -6866 -15604 -6378 -15598
rect -6866 -15638 -6819 -15604
rect -6785 -15638 -6747 -15604
rect -6713 -15638 -6675 -15604
rect -6641 -15638 -6603 -15604
rect -6569 -15638 -6531 -15604
rect -6497 -15638 -6459 -15604
rect -6425 -15638 -6378 -15604
rect -6866 -15644 -6378 -15638
rect -6660 -15706 -6600 -15644
rect -6866 -15712 -6378 -15706
rect -6866 -15746 -6819 -15712
rect -6785 -15746 -6747 -15712
rect -6713 -15746 -6675 -15712
rect -6641 -15746 -6603 -15712
rect -6569 -15746 -6531 -15712
rect -6497 -15746 -6459 -15712
rect -6425 -15746 -6378 -15712
rect -6866 -15752 -6378 -15746
rect -7158 -15820 -7148 -15815
rect -8132 -15849 -8126 -15822
rect -8172 -15887 -8126 -15849
rect -8172 -15921 -8166 -15887
rect -8132 -15921 -8126 -15887
rect -8172 -15959 -8126 -15921
rect -8172 -15993 -8166 -15959
rect -8132 -15993 -8126 -15959
rect -8172 -16031 -8126 -15993
rect -8172 -16065 -8166 -16031
rect -8132 -16065 -8126 -16031
rect -8172 -16103 -8126 -16065
rect -8172 -16137 -8166 -16103
rect -8132 -16137 -8126 -16103
rect -8172 -16175 -8126 -16137
rect -8172 -16209 -8166 -16175
rect -8132 -16209 -8126 -16175
rect -8172 -16247 -8126 -16209
rect -8172 -16281 -8166 -16247
rect -8132 -16281 -8126 -16247
rect -8172 -16319 -8126 -16281
rect -8172 -16352 -8166 -16319
rect -9190 -16356 -9144 -16353
rect -8178 -16353 -8166 -16352
rect -8132 -16352 -8126 -16319
rect -7154 -15849 -7148 -15820
rect -7114 -15820 -7098 -15815
rect -6140 -15815 -6080 -15535
rect -5120 -15535 -5112 -15526
rect -5078 -15526 -5072 -15501
rect -4100 -15031 -4094 -15012
rect -4060 -15012 -4048 -14997
rect -3086 -14997 -3026 -14722
rect -2794 -14786 -2306 -14780
rect -2794 -14820 -2747 -14786
rect -2713 -14820 -2675 -14786
rect -2641 -14820 -2603 -14786
rect -2569 -14820 -2531 -14786
rect -2497 -14820 -2459 -14786
rect -2425 -14820 -2387 -14786
rect -2353 -14820 -2306 -14786
rect -2794 -14826 -2306 -14820
rect -2588 -14888 -2528 -14826
rect -2794 -14894 -2306 -14888
rect -2794 -14928 -2747 -14894
rect -2713 -14928 -2675 -14894
rect -2641 -14928 -2603 -14894
rect -2569 -14928 -2531 -14894
rect -2497 -14928 -2459 -14894
rect -2425 -14928 -2387 -14894
rect -2353 -14928 -2306 -14894
rect -2794 -14934 -2306 -14928
rect -3086 -15012 -3076 -14997
rect -4060 -15031 -4054 -15012
rect -4100 -15069 -4054 -15031
rect -4100 -15103 -4094 -15069
rect -4060 -15103 -4054 -15069
rect -4100 -15141 -4054 -15103
rect -4100 -15175 -4094 -15141
rect -4060 -15175 -4054 -15141
rect -4100 -15213 -4054 -15175
rect -4100 -15247 -4094 -15213
rect -4060 -15247 -4054 -15213
rect -4100 -15285 -4054 -15247
rect -4100 -15319 -4094 -15285
rect -4060 -15319 -4054 -15285
rect -4100 -15357 -4054 -15319
rect -4100 -15391 -4094 -15357
rect -4060 -15391 -4054 -15357
rect -4100 -15429 -4054 -15391
rect -4100 -15463 -4094 -15429
rect -4060 -15463 -4054 -15429
rect -4100 -15501 -4054 -15463
rect -5078 -15535 -5060 -15526
rect -4100 -15534 -4094 -15501
rect -5848 -15604 -5360 -15598
rect -5848 -15638 -5801 -15604
rect -5767 -15638 -5729 -15604
rect -5695 -15638 -5657 -15604
rect -5623 -15638 -5585 -15604
rect -5551 -15638 -5513 -15604
rect -5479 -15638 -5441 -15604
rect -5407 -15638 -5360 -15604
rect -5848 -15644 -5360 -15638
rect -5658 -15706 -5598 -15644
rect -5848 -15712 -5360 -15706
rect -5848 -15746 -5801 -15712
rect -5767 -15746 -5729 -15712
rect -5695 -15746 -5657 -15712
rect -5623 -15746 -5585 -15712
rect -5551 -15746 -5513 -15712
rect -5479 -15746 -5441 -15712
rect -5407 -15746 -5360 -15712
rect -5848 -15752 -5360 -15746
rect -7114 -15849 -7108 -15820
rect -6140 -15824 -6130 -15815
rect -7154 -15887 -7108 -15849
rect -7154 -15921 -7148 -15887
rect -7114 -15921 -7108 -15887
rect -7154 -15959 -7108 -15921
rect -7154 -15993 -7148 -15959
rect -7114 -15993 -7108 -15959
rect -7154 -16031 -7108 -15993
rect -7154 -16065 -7148 -16031
rect -7114 -16065 -7108 -16031
rect -7154 -16103 -7108 -16065
rect -7154 -16137 -7148 -16103
rect -7114 -16137 -7108 -16103
rect -7154 -16175 -7108 -16137
rect -7154 -16209 -7148 -16175
rect -7114 -16209 -7108 -16175
rect -7154 -16247 -7108 -16209
rect -7154 -16281 -7148 -16247
rect -7114 -16281 -7108 -16247
rect -7154 -16319 -7108 -16281
rect -7154 -16350 -7148 -16319
rect -8132 -16353 -8118 -16352
rect -12328 -16411 -12216 -16373
rect -12328 -16445 -12289 -16411
rect -12255 -16445 -12216 -16411
rect -12328 -16483 -12216 -16445
rect -12328 -16517 -12289 -16483
rect -12255 -16517 -12216 -16483
rect -12328 -16555 -12216 -16517
rect -12328 -16589 -12289 -16555
rect -12255 -16589 -12216 -16555
rect -12328 -16627 -12216 -16589
rect -12328 -16661 -12289 -16627
rect -12255 -16661 -12216 -16627
rect -9198 -16633 -9138 -16356
rect -8902 -16422 -8414 -16416
rect -8902 -16456 -8855 -16422
rect -8821 -16456 -8783 -16422
rect -8749 -16456 -8711 -16422
rect -8677 -16456 -8639 -16422
rect -8605 -16456 -8567 -16422
rect -8533 -16456 -8495 -16422
rect -8461 -16456 -8414 -16422
rect -8902 -16462 -8414 -16456
rect -8692 -16524 -8632 -16462
rect -8902 -16530 -8414 -16524
rect -8902 -16564 -8855 -16530
rect -8821 -16564 -8783 -16530
rect -8749 -16564 -8711 -16530
rect -8677 -16564 -8639 -16530
rect -8605 -16564 -8567 -16530
rect -8533 -16564 -8495 -16530
rect -8461 -16564 -8414 -16530
rect -8902 -16570 -8414 -16564
rect -9198 -16646 -9184 -16633
rect -12328 -16699 -12216 -16661
rect -12328 -16733 -12289 -16699
rect -12255 -16733 -12216 -16699
rect -12328 -16771 -12216 -16733
rect -12328 -16805 -12289 -16771
rect -12255 -16805 -12216 -16771
rect -12328 -16843 -12216 -16805
rect -12328 -16877 -12289 -16843
rect -12255 -16877 -12216 -16843
rect -12328 -16915 -12216 -16877
rect -12328 -16949 -12289 -16915
rect -12255 -16949 -12216 -16915
rect -12328 -16987 -12216 -16949
rect -12328 -17021 -12289 -16987
rect -12255 -17021 -12216 -16987
rect -12328 -17059 -12216 -17021
rect -12328 -17093 -12289 -17059
rect -12255 -17093 -12216 -17059
rect -12328 -17131 -12216 -17093
rect -12328 -17165 -12289 -17131
rect -12255 -17165 -12216 -17131
rect -12328 -17203 -12216 -17165
rect -9190 -16667 -9184 -16646
rect -9150 -16646 -9138 -16633
rect -8178 -16633 -8118 -16353
rect -7158 -16353 -7148 -16350
rect -7114 -16350 -7108 -16319
rect -6136 -15849 -6130 -15824
rect -6096 -15824 -6080 -15815
rect -5120 -15815 -5060 -15535
rect -4108 -15535 -4094 -15534
rect -4060 -15534 -4054 -15501
rect -3082 -15031 -3076 -15012
rect -3042 -15012 -3026 -14997
rect -2066 -14997 -2006 -14722
rect -1776 -14786 -1288 -14780
rect -1776 -14820 -1729 -14786
rect -1695 -14820 -1657 -14786
rect -1623 -14820 -1585 -14786
rect -1551 -14820 -1513 -14786
rect -1479 -14820 -1441 -14786
rect -1407 -14820 -1369 -14786
rect -1335 -14820 -1288 -14786
rect -1776 -14826 -1288 -14820
rect -1576 -14888 -1516 -14826
rect -1776 -14894 -1288 -14888
rect -1776 -14928 -1729 -14894
rect -1695 -14928 -1657 -14894
rect -1623 -14928 -1585 -14894
rect -1551 -14928 -1513 -14894
rect -1479 -14928 -1441 -14894
rect -1407 -14928 -1369 -14894
rect -1335 -14928 -1288 -14894
rect -1776 -14934 -1288 -14928
rect -2066 -15012 -2058 -14997
rect -3042 -15031 -3036 -15012
rect -3082 -15069 -3036 -15031
rect -3082 -15103 -3076 -15069
rect -3042 -15103 -3036 -15069
rect -3082 -15141 -3036 -15103
rect -3082 -15175 -3076 -15141
rect -3042 -15175 -3036 -15141
rect -3082 -15213 -3036 -15175
rect -3082 -15247 -3076 -15213
rect -3042 -15247 -3036 -15213
rect -3082 -15285 -3036 -15247
rect -3082 -15319 -3076 -15285
rect -3042 -15319 -3036 -15285
rect -3082 -15357 -3036 -15319
rect -3082 -15391 -3076 -15357
rect -3042 -15391 -3036 -15357
rect -3082 -15429 -3036 -15391
rect -3082 -15463 -3076 -15429
rect -3042 -15463 -3036 -15429
rect -3082 -15501 -3036 -15463
rect -3082 -15534 -3076 -15501
rect -4060 -15535 -4048 -15534
rect -4830 -15604 -4342 -15598
rect -4830 -15638 -4783 -15604
rect -4749 -15638 -4711 -15604
rect -4677 -15638 -4639 -15604
rect -4605 -15638 -4567 -15604
rect -4533 -15638 -4495 -15604
rect -4461 -15638 -4423 -15604
rect -4389 -15638 -4342 -15604
rect -4830 -15644 -4342 -15638
rect -4628 -15706 -4568 -15644
rect -4830 -15712 -4342 -15706
rect -4830 -15746 -4783 -15712
rect -4749 -15746 -4711 -15712
rect -4677 -15746 -4639 -15712
rect -4605 -15746 -4567 -15712
rect -4533 -15746 -4495 -15712
rect -4461 -15746 -4423 -15712
rect -4389 -15746 -4342 -15712
rect -4830 -15752 -4342 -15746
rect -5120 -15816 -5112 -15815
rect -6096 -15849 -6090 -15824
rect -6136 -15887 -6090 -15849
rect -6136 -15921 -6130 -15887
rect -6096 -15921 -6090 -15887
rect -6136 -15959 -6090 -15921
rect -6136 -15993 -6130 -15959
rect -6096 -15993 -6090 -15959
rect -6136 -16031 -6090 -15993
rect -6136 -16065 -6130 -16031
rect -6096 -16065 -6090 -16031
rect -6136 -16103 -6090 -16065
rect -6136 -16137 -6130 -16103
rect -6096 -16137 -6090 -16103
rect -6136 -16175 -6090 -16137
rect -6136 -16209 -6130 -16175
rect -6096 -16209 -6090 -16175
rect -6136 -16247 -6090 -16209
rect -6136 -16281 -6130 -16247
rect -6096 -16281 -6090 -16247
rect -6136 -16319 -6090 -16281
rect -7114 -16353 -7098 -16350
rect -7884 -16422 -7396 -16416
rect -7884 -16456 -7837 -16422
rect -7803 -16456 -7765 -16422
rect -7731 -16456 -7693 -16422
rect -7659 -16456 -7621 -16422
rect -7587 -16456 -7549 -16422
rect -7515 -16456 -7477 -16422
rect -7443 -16456 -7396 -16422
rect -7884 -16462 -7396 -16456
rect -7678 -16524 -7618 -16462
rect -7884 -16530 -7396 -16524
rect -7884 -16564 -7837 -16530
rect -7803 -16564 -7765 -16530
rect -7731 -16564 -7693 -16530
rect -7659 -16564 -7621 -16530
rect -7587 -16564 -7549 -16530
rect -7515 -16564 -7477 -16530
rect -7443 -16564 -7396 -16530
rect -7884 -16570 -7396 -16564
rect -8178 -16642 -8166 -16633
rect -9150 -16667 -9144 -16646
rect -9190 -16705 -9144 -16667
rect -9190 -16739 -9184 -16705
rect -9150 -16739 -9144 -16705
rect -9190 -16777 -9144 -16739
rect -9190 -16811 -9184 -16777
rect -9150 -16811 -9144 -16777
rect -9190 -16849 -9144 -16811
rect -9190 -16883 -9184 -16849
rect -9150 -16883 -9144 -16849
rect -9190 -16921 -9144 -16883
rect -9190 -16955 -9184 -16921
rect -9150 -16955 -9144 -16921
rect -9190 -16993 -9144 -16955
rect -9190 -17027 -9184 -16993
rect -9150 -17027 -9144 -16993
rect -9190 -17065 -9144 -17027
rect -9190 -17099 -9184 -17065
rect -9150 -17099 -9144 -17065
rect -9190 -17137 -9144 -17099
rect -9190 -17168 -9184 -17137
rect -12328 -17237 -12289 -17203
rect -12255 -17237 -12216 -17203
rect -12328 -17275 -12216 -17237
rect -12328 -17309 -12289 -17275
rect -12255 -17309 -12216 -17275
rect -12328 -17347 -12216 -17309
rect -12328 -17381 -12289 -17347
rect -12255 -17381 -12216 -17347
rect -12328 -17419 -12216 -17381
rect -12328 -17453 -12289 -17419
rect -12255 -17453 -12216 -17419
rect -12328 -17491 -12216 -17453
rect -9198 -17171 -9184 -17168
rect -9150 -17168 -9144 -17137
rect -8172 -16667 -8166 -16642
rect -8132 -16642 -8118 -16633
rect -7158 -16633 -7098 -16353
rect -6136 -16353 -6130 -16319
rect -6096 -16353 -6090 -16319
rect -5118 -15849 -5112 -15816
rect -5078 -15816 -5060 -15815
rect -4108 -15815 -4048 -15535
rect -3086 -15535 -3076 -15534
rect -3042 -15534 -3036 -15501
rect -2064 -15031 -2058 -15012
rect -2024 -15012 -2006 -14997
rect -1050 -14997 -990 -14718
rect -28 -14722 18 -14717
rect -758 -14786 -270 -14780
rect -758 -14820 -711 -14786
rect -677 -14820 -639 -14786
rect -605 -14820 -567 -14786
rect -533 -14820 -495 -14786
rect -461 -14820 -423 -14786
rect -389 -14820 -351 -14786
rect -317 -14820 -270 -14786
rect -758 -14826 -270 -14820
rect -556 -14888 -496 -14826
rect -758 -14894 -270 -14888
rect -758 -14928 -711 -14894
rect -677 -14928 -639 -14894
rect -605 -14928 -567 -14894
rect -533 -14928 -495 -14894
rect -461 -14928 -423 -14894
rect -389 -14928 -351 -14894
rect -317 -14928 -270 -14894
rect -758 -14934 -270 -14928
rect -1050 -15008 -1040 -14997
rect -2024 -15031 -2018 -15012
rect -2064 -15069 -2018 -15031
rect -2064 -15103 -2058 -15069
rect -2024 -15103 -2018 -15069
rect -2064 -15141 -2018 -15103
rect -2064 -15175 -2058 -15141
rect -2024 -15175 -2018 -15141
rect -2064 -15213 -2018 -15175
rect -2064 -15247 -2058 -15213
rect -2024 -15247 -2018 -15213
rect -2064 -15285 -2018 -15247
rect -2064 -15319 -2058 -15285
rect -2024 -15319 -2018 -15285
rect -2064 -15357 -2018 -15319
rect -2064 -15391 -2058 -15357
rect -2024 -15391 -2018 -15357
rect -2064 -15429 -2018 -15391
rect -2064 -15463 -2058 -15429
rect -2024 -15463 -2018 -15429
rect -2064 -15501 -2018 -15463
rect -2064 -15534 -2058 -15501
rect -3042 -15535 -3026 -15534
rect -3812 -15604 -3324 -15598
rect -3812 -15638 -3765 -15604
rect -3731 -15638 -3693 -15604
rect -3659 -15638 -3621 -15604
rect -3587 -15638 -3549 -15604
rect -3515 -15638 -3477 -15604
rect -3443 -15638 -3405 -15604
rect -3371 -15638 -3324 -15604
rect -3812 -15644 -3324 -15638
rect -3612 -15706 -3552 -15644
rect -3812 -15712 -3324 -15706
rect -3812 -15746 -3765 -15712
rect -3731 -15746 -3693 -15712
rect -3659 -15746 -3621 -15712
rect -3587 -15746 -3549 -15712
rect -3515 -15746 -3477 -15712
rect -3443 -15746 -3405 -15712
rect -3371 -15746 -3324 -15712
rect -3812 -15752 -3324 -15746
rect -5078 -15849 -5072 -15816
rect -4108 -15824 -4094 -15815
rect -5118 -15887 -5072 -15849
rect -5118 -15921 -5112 -15887
rect -5078 -15921 -5072 -15887
rect -5118 -15959 -5072 -15921
rect -5118 -15993 -5112 -15959
rect -5078 -15993 -5072 -15959
rect -5118 -16031 -5072 -15993
rect -5118 -16065 -5112 -16031
rect -5078 -16065 -5072 -16031
rect -5118 -16103 -5072 -16065
rect -5118 -16137 -5112 -16103
rect -5078 -16137 -5072 -16103
rect -5118 -16175 -5072 -16137
rect -5118 -16209 -5112 -16175
rect -5078 -16209 -5072 -16175
rect -5118 -16247 -5072 -16209
rect -5118 -16281 -5112 -16247
rect -5078 -16281 -5072 -16247
rect -5118 -16319 -5072 -16281
rect -5118 -16346 -5112 -16319
rect -6136 -16354 -6090 -16353
rect -5120 -16353 -5112 -16346
rect -5078 -16346 -5072 -16319
rect -4100 -15849 -4094 -15824
rect -4060 -15824 -4048 -15815
rect -3086 -15815 -3026 -15535
rect -2066 -15535 -2058 -15534
rect -2024 -15534 -2018 -15501
rect -1046 -15031 -1040 -15008
rect -1006 -15008 -990 -14997
rect -28 -14997 32 -14722
rect 1850 -14902 1910 -12508
rect 2110 -13782 2170 -11408
rect 2336 -11412 2340 -11360
rect 2392 -11412 2396 -11360
rect 2110 -13792 2172 -13782
rect 2110 -13844 2116 -13792
rect 2168 -13844 2172 -13792
rect 2110 -13854 2172 -13844
rect 1970 -14004 2042 -14000
rect 1970 -14056 1980 -14004
rect 2032 -14056 2042 -14004
rect 1970 -14060 2042 -14056
rect 1844 -14906 1916 -14902
rect 1844 -14958 1854 -14906
rect 1906 -14958 1916 -14906
rect 1844 -14962 1916 -14958
rect -1006 -15031 -1000 -15008
rect -1046 -15069 -1000 -15031
rect -1046 -15103 -1040 -15069
rect -1006 -15103 -1000 -15069
rect -1046 -15141 -1000 -15103
rect -1046 -15175 -1040 -15141
rect -1006 -15175 -1000 -15141
rect -1046 -15213 -1000 -15175
rect -1046 -15247 -1040 -15213
rect -1006 -15247 -1000 -15213
rect -1046 -15285 -1000 -15247
rect -1046 -15319 -1040 -15285
rect -1006 -15319 -1000 -15285
rect -1046 -15357 -1000 -15319
rect -1046 -15391 -1040 -15357
rect -1006 -15391 -1000 -15357
rect -1046 -15429 -1000 -15391
rect -1046 -15463 -1040 -15429
rect -1006 -15463 -1000 -15429
rect -1046 -15501 -1000 -15463
rect -1046 -15530 -1040 -15501
rect -2024 -15535 -2006 -15534
rect -2794 -15604 -2306 -15598
rect -2794 -15638 -2747 -15604
rect -2713 -15638 -2675 -15604
rect -2641 -15638 -2603 -15604
rect -2569 -15638 -2531 -15604
rect -2497 -15638 -2459 -15604
rect -2425 -15638 -2387 -15604
rect -2353 -15638 -2306 -15604
rect -2794 -15644 -2306 -15638
rect -2590 -15706 -2530 -15644
rect -2794 -15712 -2306 -15706
rect -2794 -15746 -2747 -15712
rect -2713 -15746 -2675 -15712
rect -2641 -15746 -2603 -15712
rect -2569 -15746 -2531 -15712
rect -2497 -15746 -2459 -15712
rect -2425 -15746 -2387 -15712
rect -2353 -15746 -2306 -15712
rect -2794 -15752 -2306 -15746
rect -3086 -15824 -3076 -15815
rect -4060 -15849 -4054 -15824
rect -4100 -15887 -4054 -15849
rect -4100 -15921 -4094 -15887
rect -4060 -15921 -4054 -15887
rect -4100 -15959 -4054 -15921
rect -4100 -15993 -4094 -15959
rect -4060 -15993 -4054 -15959
rect -4100 -16031 -4054 -15993
rect -4100 -16065 -4094 -16031
rect -4060 -16065 -4054 -16031
rect -4100 -16103 -4054 -16065
rect -4100 -16137 -4094 -16103
rect -4060 -16137 -4054 -16103
rect -4100 -16175 -4054 -16137
rect -4100 -16209 -4094 -16175
rect -4060 -16209 -4054 -16175
rect -4100 -16247 -4054 -16209
rect -4100 -16281 -4094 -16247
rect -4060 -16281 -4054 -16247
rect -4100 -16319 -4054 -16281
rect -5078 -16353 -5060 -16346
rect -6866 -16422 -6378 -16416
rect -6866 -16456 -6819 -16422
rect -6785 -16456 -6747 -16422
rect -6713 -16456 -6675 -16422
rect -6641 -16456 -6603 -16422
rect -6569 -16456 -6531 -16422
rect -6497 -16456 -6459 -16422
rect -6425 -16456 -6378 -16422
rect -6866 -16462 -6378 -16456
rect -6658 -16524 -6598 -16462
rect -6866 -16530 -6378 -16524
rect -6866 -16564 -6819 -16530
rect -6785 -16564 -6747 -16530
rect -6713 -16564 -6675 -16530
rect -6641 -16564 -6603 -16530
rect -6569 -16564 -6531 -16530
rect -6497 -16564 -6459 -16530
rect -6425 -16564 -6378 -16530
rect -6866 -16570 -6378 -16564
rect -7158 -16640 -7148 -16633
rect -8132 -16667 -8126 -16642
rect -8172 -16705 -8126 -16667
rect -8172 -16739 -8166 -16705
rect -8132 -16739 -8126 -16705
rect -8172 -16777 -8126 -16739
rect -8172 -16811 -8166 -16777
rect -8132 -16811 -8126 -16777
rect -8172 -16849 -8126 -16811
rect -8172 -16883 -8166 -16849
rect -8132 -16883 -8126 -16849
rect -8172 -16921 -8126 -16883
rect -8172 -16955 -8166 -16921
rect -8132 -16955 -8126 -16921
rect -8172 -16993 -8126 -16955
rect -8172 -17027 -8166 -16993
rect -8132 -17027 -8126 -16993
rect -8172 -17065 -8126 -17027
rect -8172 -17099 -8166 -17065
rect -8132 -17099 -8126 -17065
rect -8172 -17137 -8126 -17099
rect -8172 -17164 -8166 -17137
rect -9150 -17171 -9138 -17168
rect -9198 -17451 -9138 -17171
rect -8178 -17171 -8166 -17164
rect -8132 -17164 -8126 -17137
rect -7154 -16667 -7148 -16640
rect -7114 -16640 -7098 -16633
rect -6140 -16633 -6080 -16354
rect -5848 -16422 -5360 -16416
rect -5848 -16456 -5801 -16422
rect -5767 -16456 -5729 -16422
rect -5695 -16456 -5657 -16422
rect -5623 -16456 -5585 -16422
rect -5551 -16456 -5513 -16422
rect -5479 -16456 -5441 -16422
rect -5407 -16456 -5360 -16422
rect -5848 -16462 -5360 -16456
rect -5656 -16524 -5596 -16462
rect -5848 -16530 -5360 -16524
rect -5848 -16564 -5801 -16530
rect -5767 -16564 -5729 -16530
rect -5695 -16564 -5657 -16530
rect -5623 -16564 -5585 -16530
rect -5551 -16564 -5513 -16530
rect -5479 -16564 -5441 -16530
rect -5407 -16564 -5360 -16530
rect -5848 -16570 -5360 -16564
rect -7114 -16667 -7108 -16640
rect -6140 -16644 -6130 -16633
rect -7154 -16705 -7108 -16667
rect -7154 -16739 -7148 -16705
rect -7114 -16739 -7108 -16705
rect -7154 -16777 -7108 -16739
rect -7154 -16811 -7148 -16777
rect -7114 -16811 -7108 -16777
rect -7154 -16849 -7108 -16811
rect -7154 -16883 -7148 -16849
rect -7114 -16883 -7108 -16849
rect -7154 -16921 -7108 -16883
rect -7154 -16955 -7148 -16921
rect -7114 -16955 -7108 -16921
rect -7154 -16993 -7108 -16955
rect -7154 -17027 -7148 -16993
rect -7114 -17027 -7108 -16993
rect -7154 -17065 -7108 -17027
rect -7154 -17099 -7148 -17065
rect -7114 -17099 -7108 -17065
rect -7154 -17137 -7108 -17099
rect -7154 -17162 -7148 -17137
rect -8132 -17171 -8118 -17164
rect -8902 -17240 -8414 -17234
rect -8902 -17274 -8855 -17240
rect -8821 -17274 -8783 -17240
rect -8749 -17274 -8711 -17240
rect -8677 -17274 -8639 -17240
rect -8605 -17274 -8567 -17240
rect -8533 -17274 -8495 -17240
rect -8461 -17274 -8414 -17240
rect -8902 -17280 -8414 -17274
rect -8690 -17342 -8630 -17280
rect -8902 -17348 -8414 -17342
rect -8902 -17382 -8855 -17348
rect -8821 -17382 -8783 -17348
rect -8749 -17382 -8711 -17348
rect -8677 -17382 -8639 -17348
rect -8605 -17382 -8567 -17348
rect -8533 -17382 -8495 -17348
rect -8461 -17382 -8414 -17348
rect -8902 -17388 -8414 -17382
rect -9198 -17458 -9184 -17451
rect -12328 -17525 -12289 -17491
rect -12255 -17525 -12216 -17491
rect -12328 -17563 -12216 -17525
rect -12328 -17597 -12289 -17563
rect -12255 -17597 -12216 -17563
rect -12328 -17635 -12216 -17597
rect -12328 -17669 -12289 -17635
rect -12255 -17669 -12216 -17635
rect -12328 -17707 -12216 -17669
rect -12328 -17741 -12289 -17707
rect -12255 -17741 -12216 -17707
rect -12328 -17779 -12216 -17741
rect -12328 -17813 -12289 -17779
rect -12255 -17813 -12216 -17779
rect -12328 -17851 -12216 -17813
rect -12328 -17885 -12289 -17851
rect -12255 -17885 -12216 -17851
rect -12328 -17923 -12216 -17885
rect -12328 -17957 -12289 -17923
rect -12255 -17957 -12216 -17923
rect -12328 -17995 -12216 -17957
rect -9190 -17485 -9184 -17458
rect -9150 -17458 -9138 -17451
rect -8178 -17451 -8118 -17171
rect -7158 -17171 -7148 -17162
rect -7114 -17162 -7108 -17137
rect -6136 -16667 -6130 -16644
rect -6096 -16644 -6080 -16633
rect -5120 -16633 -5060 -16353
rect -4100 -16353 -4094 -16319
rect -4060 -16353 -4054 -16319
rect -4100 -16354 -4054 -16353
rect -3082 -15849 -3076 -15824
rect -3042 -15824 -3026 -15815
rect -2066 -15815 -2006 -15535
rect -1050 -15535 -1040 -15530
rect -1006 -15530 -1000 -15501
rect -28 -15031 -22 -14997
rect 12 -15012 32 -14997
rect 12 -15031 18 -15012
rect -28 -15069 18 -15031
rect -28 -15103 -22 -15069
rect 12 -15103 18 -15069
rect -28 -15141 18 -15103
rect -28 -15175 -22 -15141
rect 12 -15175 18 -15141
rect -28 -15213 18 -15175
rect -28 -15247 -22 -15213
rect 12 -15247 18 -15213
rect -28 -15285 18 -15247
rect -28 -15319 -22 -15285
rect 12 -15319 18 -15285
rect -28 -15357 18 -15319
rect -28 -15391 -22 -15357
rect 12 -15391 18 -15357
rect -28 -15429 18 -15391
rect -28 -15463 -22 -15429
rect 12 -15463 18 -15429
rect -28 -15501 18 -15463
rect -1006 -15535 -990 -15530
rect -1776 -15604 -1288 -15598
rect -1776 -15638 -1729 -15604
rect -1695 -15638 -1657 -15604
rect -1623 -15638 -1585 -15604
rect -1551 -15638 -1513 -15604
rect -1479 -15638 -1441 -15604
rect -1407 -15638 -1369 -15604
rect -1335 -15638 -1288 -15604
rect -1776 -15644 -1288 -15638
rect -1578 -15706 -1518 -15644
rect -1776 -15712 -1288 -15706
rect -1776 -15746 -1729 -15712
rect -1695 -15746 -1657 -15712
rect -1623 -15746 -1585 -15712
rect -1551 -15746 -1513 -15712
rect -1479 -15746 -1441 -15712
rect -1407 -15746 -1369 -15712
rect -1335 -15746 -1288 -15712
rect -1776 -15752 -1288 -15746
rect -2066 -15824 -2058 -15815
rect -3042 -15849 -3036 -15824
rect -3082 -15887 -3036 -15849
rect -3082 -15921 -3076 -15887
rect -3042 -15921 -3036 -15887
rect -3082 -15959 -3036 -15921
rect -3082 -15993 -3076 -15959
rect -3042 -15993 -3036 -15959
rect -3082 -16031 -3036 -15993
rect -3082 -16065 -3076 -16031
rect -3042 -16065 -3036 -16031
rect -3082 -16103 -3036 -16065
rect -3082 -16137 -3076 -16103
rect -3042 -16137 -3036 -16103
rect -3082 -16175 -3036 -16137
rect -3082 -16209 -3076 -16175
rect -3042 -16209 -3036 -16175
rect -3082 -16247 -3036 -16209
rect -3082 -16281 -3076 -16247
rect -3042 -16281 -3036 -16247
rect -3082 -16319 -3036 -16281
rect -3082 -16353 -3076 -16319
rect -3042 -16353 -3036 -16319
rect -3082 -16354 -3036 -16353
rect -2064 -15849 -2058 -15824
rect -2024 -15824 -2006 -15815
rect -1050 -15815 -990 -15535
rect -28 -15535 -22 -15501
rect 12 -15534 18 -15501
rect 12 -15535 32 -15534
rect -758 -15604 -270 -15598
rect -758 -15638 -711 -15604
rect -677 -15638 -639 -15604
rect -605 -15638 -567 -15604
rect -533 -15638 -495 -15604
rect -461 -15638 -423 -15604
rect -389 -15638 -351 -15604
rect -317 -15638 -270 -15604
rect -758 -15644 -270 -15638
rect -558 -15706 -498 -15644
rect -758 -15712 -270 -15706
rect -758 -15746 -711 -15712
rect -677 -15746 -639 -15712
rect -605 -15746 -567 -15712
rect -533 -15746 -495 -15712
rect -461 -15746 -423 -15712
rect -389 -15746 -351 -15712
rect -317 -15746 -270 -15712
rect -758 -15752 -270 -15746
rect -1050 -15820 -1040 -15815
rect -2024 -15849 -2018 -15824
rect -2064 -15887 -2018 -15849
rect -2064 -15921 -2058 -15887
rect -2024 -15921 -2018 -15887
rect -2064 -15959 -2018 -15921
rect -2064 -15993 -2058 -15959
rect -2024 -15993 -2018 -15959
rect -2064 -16031 -2018 -15993
rect -2064 -16065 -2058 -16031
rect -2024 -16065 -2018 -16031
rect -2064 -16103 -2018 -16065
rect -2064 -16137 -2058 -16103
rect -2024 -16137 -2018 -16103
rect -2064 -16175 -2018 -16137
rect -2064 -16209 -2058 -16175
rect -2024 -16209 -2018 -16175
rect -2064 -16247 -2018 -16209
rect -2064 -16281 -2058 -16247
rect -2024 -16281 -2018 -16247
rect -2064 -16319 -2018 -16281
rect -2064 -16353 -2058 -16319
rect -2024 -16353 -2018 -16319
rect -1046 -15849 -1040 -15820
rect -1006 -15820 -990 -15815
rect -28 -15815 32 -15535
rect -1006 -15849 -1000 -15820
rect -1046 -15887 -1000 -15849
rect -1046 -15921 -1040 -15887
rect -1006 -15921 -1000 -15887
rect -1046 -15959 -1000 -15921
rect -1046 -15993 -1040 -15959
rect -1006 -15993 -1000 -15959
rect -1046 -16031 -1000 -15993
rect -1046 -16065 -1040 -16031
rect -1006 -16065 -1000 -16031
rect -1046 -16103 -1000 -16065
rect -1046 -16137 -1040 -16103
rect -1006 -16137 -1000 -16103
rect -1046 -16175 -1000 -16137
rect -1046 -16209 -1040 -16175
rect -1006 -16209 -1000 -16175
rect -1046 -16247 -1000 -16209
rect -1046 -16281 -1040 -16247
rect -1006 -16281 -1000 -16247
rect -1046 -16319 -1000 -16281
rect -1046 -16350 -1040 -16319
rect -2064 -16354 -2018 -16353
rect -1050 -16353 -1040 -16350
rect -1006 -16350 -1000 -16319
rect -28 -15849 -22 -15815
rect 12 -15824 32 -15815
rect 12 -15849 18 -15824
rect -28 -15887 18 -15849
rect -28 -15921 -22 -15887
rect 12 -15921 18 -15887
rect -28 -15959 18 -15921
rect -28 -15993 -22 -15959
rect 12 -15993 18 -15959
rect -28 -16031 18 -15993
rect -28 -16065 -22 -16031
rect 12 -16065 18 -16031
rect -28 -16103 18 -16065
rect -28 -16137 -22 -16103
rect 12 -16137 18 -16103
rect -28 -16175 18 -16137
rect -28 -16209 -22 -16175
rect 12 -16209 18 -16175
rect -28 -16247 18 -16209
rect -28 -16281 -22 -16247
rect 12 -16281 18 -16247
rect -28 -16319 18 -16281
rect -1006 -16353 -990 -16350
rect -4830 -16422 -4342 -16416
rect -4830 -16456 -4783 -16422
rect -4749 -16456 -4711 -16422
rect -4677 -16456 -4639 -16422
rect -4605 -16456 -4567 -16422
rect -4533 -16456 -4495 -16422
rect -4461 -16456 -4423 -16422
rect -4389 -16456 -4342 -16422
rect -4830 -16462 -4342 -16456
rect -4626 -16524 -4566 -16462
rect -4830 -16530 -4342 -16524
rect -4830 -16564 -4783 -16530
rect -4749 -16564 -4711 -16530
rect -4677 -16564 -4639 -16530
rect -4605 -16564 -4567 -16530
rect -4533 -16564 -4495 -16530
rect -4461 -16564 -4423 -16530
rect -4389 -16564 -4342 -16530
rect -4830 -16570 -4342 -16564
rect -5120 -16636 -5112 -16633
rect -6096 -16667 -6090 -16644
rect -6136 -16705 -6090 -16667
rect -6136 -16739 -6130 -16705
rect -6096 -16739 -6090 -16705
rect -6136 -16777 -6090 -16739
rect -6136 -16811 -6130 -16777
rect -6096 -16811 -6090 -16777
rect -6136 -16849 -6090 -16811
rect -6136 -16883 -6130 -16849
rect -6096 -16883 -6090 -16849
rect -6136 -16921 -6090 -16883
rect -6136 -16955 -6130 -16921
rect -6096 -16955 -6090 -16921
rect -6136 -16993 -6090 -16955
rect -6136 -17027 -6130 -16993
rect -6096 -17027 -6090 -16993
rect -6136 -17065 -6090 -17027
rect -6136 -17099 -6130 -17065
rect -6096 -17099 -6090 -17065
rect -6136 -17137 -6090 -17099
rect -7114 -17171 -7098 -17162
rect -6136 -17166 -6130 -17137
rect -7884 -17240 -7396 -17234
rect -7884 -17274 -7837 -17240
rect -7803 -17274 -7765 -17240
rect -7731 -17274 -7693 -17240
rect -7659 -17274 -7621 -17240
rect -7587 -17274 -7549 -17240
rect -7515 -17274 -7477 -17240
rect -7443 -17274 -7396 -17240
rect -7884 -17280 -7396 -17274
rect -7676 -17342 -7616 -17280
rect -7884 -17348 -7396 -17342
rect -7884 -17382 -7837 -17348
rect -7803 -17382 -7765 -17348
rect -7731 -17382 -7693 -17348
rect -7659 -17382 -7621 -17348
rect -7587 -17382 -7549 -17348
rect -7515 -17382 -7477 -17348
rect -7443 -17382 -7396 -17348
rect -7884 -17388 -7396 -17382
rect -8178 -17454 -8166 -17451
rect -9150 -17485 -9144 -17458
rect -9190 -17523 -9144 -17485
rect -9190 -17557 -9184 -17523
rect -9150 -17557 -9144 -17523
rect -9190 -17595 -9144 -17557
rect -9190 -17629 -9184 -17595
rect -9150 -17629 -9144 -17595
rect -9190 -17667 -9144 -17629
rect -9190 -17701 -9184 -17667
rect -9150 -17701 -9144 -17667
rect -9190 -17739 -9144 -17701
rect -9190 -17773 -9184 -17739
rect -9150 -17773 -9144 -17739
rect -9190 -17811 -9144 -17773
rect -9190 -17845 -9184 -17811
rect -9150 -17845 -9144 -17811
rect -9190 -17883 -9144 -17845
rect -9190 -17917 -9184 -17883
rect -9150 -17917 -9144 -17883
rect -9190 -17955 -9144 -17917
rect -9190 -17986 -9184 -17955
rect -12328 -18029 -12289 -17995
rect -12255 -18029 -12216 -17995
rect -12328 -18067 -12216 -18029
rect -12328 -18101 -12289 -18067
rect -12255 -18101 -12216 -18067
rect -12328 -18139 -12216 -18101
rect -12328 -18173 -12289 -18139
rect -12255 -18173 -12216 -18139
rect -12328 -18211 -12216 -18173
rect -12328 -18245 -12289 -18211
rect -12255 -18245 -12216 -18211
rect -12328 -18283 -12216 -18245
rect -9198 -17989 -9184 -17986
rect -9150 -17986 -9144 -17955
rect -8172 -17485 -8166 -17454
rect -8132 -17454 -8118 -17451
rect -7158 -17451 -7098 -17171
rect -6140 -17171 -6130 -17166
rect -6096 -17166 -6090 -17137
rect -5118 -16667 -5112 -16636
rect -5078 -16636 -5060 -16633
rect -4108 -16633 -4048 -16354
rect -3812 -16422 -3324 -16416
rect -3812 -16456 -3765 -16422
rect -3731 -16456 -3693 -16422
rect -3659 -16456 -3621 -16422
rect -3587 -16456 -3549 -16422
rect -3515 -16456 -3477 -16422
rect -3443 -16456 -3405 -16422
rect -3371 -16456 -3324 -16422
rect -3812 -16462 -3324 -16456
rect -3610 -16524 -3550 -16462
rect -3812 -16530 -3324 -16524
rect -3812 -16564 -3765 -16530
rect -3731 -16564 -3693 -16530
rect -3659 -16564 -3621 -16530
rect -3587 -16564 -3549 -16530
rect -3515 -16564 -3477 -16530
rect -3443 -16564 -3405 -16530
rect -3371 -16564 -3324 -16530
rect -3812 -16570 -3324 -16564
rect -5078 -16667 -5072 -16636
rect -4108 -16644 -4094 -16633
rect -5118 -16705 -5072 -16667
rect -5118 -16739 -5112 -16705
rect -5078 -16739 -5072 -16705
rect -5118 -16777 -5072 -16739
rect -5118 -16811 -5112 -16777
rect -5078 -16811 -5072 -16777
rect -5118 -16849 -5072 -16811
rect -5118 -16883 -5112 -16849
rect -5078 -16883 -5072 -16849
rect -5118 -16921 -5072 -16883
rect -5118 -16955 -5112 -16921
rect -5078 -16955 -5072 -16921
rect -5118 -16993 -5072 -16955
rect -5118 -17027 -5112 -16993
rect -5078 -17027 -5072 -16993
rect -5118 -17065 -5072 -17027
rect -5118 -17099 -5112 -17065
rect -5078 -17099 -5072 -17065
rect -5118 -17137 -5072 -17099
rect -5118 -17158 -5112 -17137
rect -6096 -17171 -6080 -17166
rect -6866 -17240 -6378 -17234
rect -6866 -17274 -6819 -17240
rect -6785 -17274 -6747 -17240
rect -6713 -17274 -6675 -17240
rect -6641 -17274 -6603 -17240
rect -6569 -17274 -6531 -17240
rect -6497 -17274 -6459 -17240
rect -6425 -17274 -6378 -17240
rect -6866 -17280 -6378 -17274
rect -6656 -17342 -6596 -17280
rect -6866 -17348 -6378 -17342
rect -6866 -17382 -6819 -17348
rect -6785 -17382 -6747 -17348
rect -6713 -17382 -6675 -17348
rect -6641 -17382 -6603 -17348
rect -6569 -17382 -6531 -17348
rect -6497 -17382 -6459 -17348
rect -6425 -17382 -6378 -17348
rect -6866 -17388 -6378 -17382
rect -7158 -17452 -7148 -17451
rect -8132 -17485 -8126 -17454
rect -8172 -17523 -8126 -17485
rect -8172 -17557 -8166 -17523
rect -8132 -17557 -8126 -17523
rect -8172 -17595 -8126 -17557
rect -8172 -17629 -8166 -17595
rect -8132 -17629 -8126 -17595
rect -8172 -17667 -8126 -17629
rect -8172 -17701 -8166 -17667
rect -8132 -17701 -8126 -17667
rect -8172 -17739 -8126 -17701
rect -8172 -17773 -8166 -17739
rect -8132 -17773 -8126 -17739
rect -8172 -17811 -8126 -17773
rect -8172 -17845 -8166 -17811
rect -8132 -17845 -8126 -17811
rect -8172 -17883 -8126 -17845
rect -8172 -17917 -8166 -17883
rect -8132 -17917 -8126 -17883
rect -8172 -17955 -8126 -17917
rect -8172 -17982 -8166 -17955
rect -9150 -17989 -9138 -17986
rect -9198 -18269 -9138 -17989
rect -8178 -17989 -8166 -17982
rect -8132 -17982 -8126 -17955
rect -7154 -17485 -7148 -17452
rect -7114 -17452 -7098 -17451
rect -6140 -17451 -6080 -17171
rect -5120 -17171 -5112 -17158
rect -5078 -17158 -5072 -17137
rect -4100 -16667 -4094 -16644
rect -4060 -16644 -4048 -16633
rect -3086 -16633 -3026 -16354
rect -2794 -16422 -2306 -16416
rect -2794 -16456 -2747 -16422
rect -2713 -16456 -2675 -16422
rect -2641 -16456 -2603 -16422
rect -2569 -16456 -2531 -16422
rect -2497 -16456 -2459 -16422
rect -2425 -16456 -2387 -16422
rect -2353 -16456 -2306 -16422
rect -2794 -16462 -2306 -16456
rect -2588 -16524 -2528 -16462
rect -2794 -16530 -2306 -16524
rect -2794 -16564 -2747 -16530
rect -2713 -16564 -2675 -16530
rect -2641 -16564 -2603 -16530
rect -2569 -16564 -2531 -16530
rect -2497 -16564 -2459 -16530
rect -2425 -16564 -2387 -16530
rect -2353 -16564 -2306 -16530
rect -2794 -16570 -2306 -16564
rect -3086 -16644 -3076 -16633
rect -4060 -16667 -4054 -16644
rect -4100 -16705 -4054 -16667
rect -4100 -16739 -4094 -16705
rect -4060 -16739 -4054 -16705
rect -4100 -16777 -4054 -16739
rect -4100 -16811 -4094 -16777
rect -4060 -16811 -4054 -16777
rect -4100 -16849 -4054 -16811
rect -4100 -16883 -4094 -16849
rect -4060 -16883 -4054 -16849
rect -4100 -16921 -4054 -16883
rect -4100 -16955 -4094 -16921
rect -4060 -16955 -4054 -16921
rect -4100 -16993 -4054 -16955
rect -4100 -17027 -4094 -16993
rect -4060 -17027 -4054 -16993
rect -4100 -17065 -4054 -17027
rect -4100 -17099 -4094 -17065
rect -4060 -17099 -4054 -17065
rect -4100 -17137 -4054 -17099
rect -5078 -17171 -5060 -17158
rect -4100 -17166 -4094 -17137
rect -5848 -17240 -5360 -17234
rect -5848 -17274 -5801 -17240
rect -5767 -17274 -5729 -17240
rect -5695 -17274 -5657 -17240
rect -5623 -17274 -5585 -17240
rect -5551 -17274 -5513 -17240
rect -5479 -17274 -5441 -17240
rect -5407 -17274 -5360 -17240
rect -5848 -17280 -5360 -17274
rect -5654 -17342 -5594 -17280
rect -5848 -17348 -5360 -17342
rect -5848 -17382 -5801 -17348
rect -5767 -17382 -5729 -17348
rect -5695 -17382 -5657 -17348
rect -5623 -17382 -5585 -17348
rect -5551 -17382 -5513 -17348
rect -5479 -17382 -5441 -17348
rect -5407 -17382 -5360 -17348
rect -5848 -17388 -5360 -17382
rect -5120 -17448 -5060 -17171
rect -4108 -17171 -4094 -17166
rect -4060 -17166 -4054 -17137
rect -3082 -16667 -3076 -16644
rect -3042 -16644 -3026 -16633
rect -2066 -16633 -2006 -16354
rect -1776 -16422 -1288 -16416
rect -1776 -16456 -1729 -16422
rect -1695 -16456 -1657 -16422
rect -1623 -16456 -1585 -16422
rect -1551 -16456 -1513 -16422
rect -1479 -16456 -1441 -16422
rect -1407 -16456 -1369 -16422
rect -1335 -16456 -1288 -16422
rect -1776 -16462 -1288 -16456
rect -1576 -16524 -1516 -16462
rect -1776 -16530 -1288 -16524
rect -1776 -16564 -1729 -16530
rect -1695 -16564 -1657 -16530
rect -1623 -16564 -1585 -16530
rect -1551 -16564 -1513 -16530
rect -1479 -16564 -1441 -16530
rect -1407 -16564 -1369 -16530
rect -1335 -16564 -1288 -16530
rect -1776 -16570 -1288 -16564
rect -2066 -16644 -2058 -16633
rect -3042 -16667 -3036 -16644
rect -3082 -16705 -3036 -16667
rect -3082 -16739 -3076 -16705
rect -3042 -16739 -3036 -16705
rect -3082 -16777 -3036 -16739
rect -3082 -16811 -3076 -16777
rect -3042 -16811 -3036 -16777
rect -3082 -16849 -3036 -16811
rect -3082 -16883 -3076 -16849
rect -3042 -16883 -3036 -16849
rect -3082 -16921 -3036 -16883
rect -3082 -16955 -3076 -16921
rect -3042 -16955 -3036 -16921
rect -3082 -16993 -3036 -16955
rect -3082 -17027 -3076 -16993
rect -3042 -17027 -3036 -16993
rect -3082 -17065 -3036 -17027
rect -3082 -17099 -3076 -17065
rect -3042 -17099 -3036 -17065
rect -3082 -17137 -3036 -17099
rect -3082 -17166 -3076 -17137
rect -4060 -17171 -4048 -17166
rect -4830 -17240 -4342 -17234
rect -4830 -17274 -4783 -17240
rect -4749 -17274 -4711 -17240
rect -4677 -17274 -4639 -17240
rect -4605 -17274 -4567 -17240
rect -4533 -17274 -4495 -17240
rect -4461 -17274 -4423 -17240
rect -4389 -17274 -4342 -17240
rect -4830 -17280 -4342 -17274
rect -4624 -17342 -4564 -17280
rect -4830 -17348 -4342 -17342
rect -4830 -17382 -4783 -17348
rect -4749 -17382 -4711 -17348
rect -4677 -17382 -4639 -17348
rect -4605 -17382 -4567 -17348
rect -4533 -17382 -4495 -17348
rect -4461 -17382 -4423 -17348
rect -4389 -17382 -4342 -17348
rect -4830 -17388 -4342 -17382
rect -7114 -17485 -7108 -17452
rect -6140 -17456 -6130 -17451
rect -7154 -17523 -7108 -17485
rect -7154 -17557 -7148 -17523
rect -7114 -17557 -7108 -17523
rect -7154 -17595 -7108 -17557
rect -7154 -17629 -7148 -17595
rect -7114 -17629 -7108 -17595
rect -7154 -17667 -7108 -17629
rect -7154 -17701 -7148 -17667
rect -7114 -17701 -7108 -17667
rect -7154 -17739 -7108 -17701
rect -7154 -17773 -7148 -17739
rect -7114 -17773 -7108 -17739
rect -7154 -17811 -7108 -17773
rect -7154 -17845 -7148 -17811
rect -7114 -17845 -7108 -17811
rect -7154 -17883 -7108 -17845
rect -7154 -17917 -7148 -17883
rect -7114 -17917 -7108 -17883
rect -7154 -17955 -7108 -17917
rect -7154 -17980 -7148 -17955
rect -8132 -17989 -8118 -17982
rect -8902 -18058 -8414 -18052
rect -8902 -18092 -8855 -18058
rect -8821 -18092 -8783 -18058
rect -8749 -18092 -8711 -18058
rect -8677 -18092 -8639 -18058
rect -8605 -18092 -8567 -18058
rect -8533 -18092 -8495 -18058
rect -8461 -18092 -8414 -18058
rect -8902 -18098 -8414 -18092
rect -8688 -18160 -8628 -18098
rect -8902 -18166 -8414 -18160
rect -8902 -18200 -8855 -18166
rect -8821 -18200 -8783 -18166
rect -8749 -18200 -8711 -18166
rect -8677 -18200 -8639 -18166
rect -8605 -18200 -8567 -18166
rect -8533 -18200 -8495 -18166
rect -8461 -18200 -8414 -18166
rect -8902 -18206 -8414 -18200
rect -9198 -18276 -9184 -18269
rect -12328 -18317 -12289 -18283
rect -12255 -18317 -12216 -18283
rect -12328 -18355 -12216 -18317
rect -12328 -18389 -12289 -18355
rect -12255 -18389 -12216 -18355
rect -12328 -18427 -12216 -18389
rect -12328 -18461 -12289 -18427
rect -12255 -18461 -12216 -18427
rect -12328 -18499 -12216 -18461
rect -12328 -18533 -12289 -18499
rect -12255 -18533 -12216 -18499
rect -12328 -18571 -12216 -18533
rect -12328 -18605 -12289 -18571
rect -12255 -18605 -12216 -18571
rect -12328 -18643 -12216 -18605
rect -12328 -18677 -12289 -18643
rect -12255 -18677 -12216 -18643
rect -12328 -18715 -12216 -18677
rect -12328 -18749 -12289 -18715
rect -12255 -18749 -12216 -18715
rect -12328 -18787 -12216 -18749
rect -12328 -18821 -12289 -18787
rect -12255 -18821 -12216 -18787
rect -12328 -18859 -12216 -18821
rect -9190 -18303 -9184 -18276
rect -9150 -18276 -9138 -18269
rect -8178 -18269 -8118 -17989
rect -7158 -17989 -7148 -17980
rect -7114 -17980 -7108 -17955
rect -6136 -17485 -6130 -17456
rect -6096 -17456 -6080 -17451
rect -5118 -17451 -5072 -17448
rect -6096 -17485 -6090 -17456
rect -6136 -17523 -6090 -17485
rect -6136 -17557 -6130 -17523
rect -6096 -17557 -6090 -17523
rect -6136 -17595 -6090 -17557
rect -6136 -17629 -6130 -17595
rect -6096 -17629 -6090 -17595
rect -6136 -17667 -6090 -17629
rect -6136 -17701 -6130 -17667
rect -6096 -17701 -6090 -17667
rect -6136 -17739 -6090 -17701
rect -6136 -17773 -6130 -17739
rect -6096 -17773 -6090 -17739
rect -6136 -17811 -6090 -17773
rect -6136 -17845 -6130 -17811
rect -6096 -17845 -6090 -17811
rect -6136 -17883 -6090 -17845
rect -6136 -17917 -6130 -17883
rect -6096 -17917 -6090 -17883
rect -6136 -17955 -6090 -17917
rect -7114 -17989 -7098 -17980
rect -6136 -17984 -6130 -17955
rect -7884 -18058 -7396 -18052
rect -7884 -18092 -7837 -18058
rect -7803 -18092 -7765 -18058
rect -7731 -18092 -7693 -18058
rect -7659 -18092 -7621 -18058
rect -7587 -18092 -7549 -18058
rect -7515 -18092 -7477 -18058
rect -7443 -18092 -7396 -18058
rect -7884 -18098 -7396 -18092
rect -7674 -18160 -7614 -18098
rect -7884 -18166 -7396 -18160
rect -7884 -18200 -7837 -18166
rect -7803 -18200 -7765 -18166
rect -7731 -18200 -7693 -18166
rect -7659 -18200 -7621 -18166
rect -7587 -18200 -7549 -18166
rect -7515 -18200 -7477 -18166
rect -7443 -18200 -7396 -18166
rect -7884 -18206 -7396 -18200
rect -8178 -18272 -8166 -18269
rect -9150 -18303 -9144 -18276
rect -9190 -18341 -9144 -18303
rect -9190 -18375 -9184 -18341
rect -9150 -18375 -9144 -18341
rect -9190 -18413 -9144 -18375
rect -9190 -18447 -9184 -18413
rect -9150 -18447 -9144 -18413
rect -9190 -18485 -9144 -18447
rect -9190 -18519 -9184 -18485
rect -9150 -18519 -9144 -18485
rect -9190 -18557 -9144 -18519
rect -9190 -18591 -9184 -18557
rect -9150 -18591 -9144 -18557
rect -9190 -18629 -9144 -18591
rect -9190 -18663 -9184 -18629
rect -9150 -18663 -9144 -18629
rect -9190 -18701 -9144 -18663
rect -9190 -18735 -9184 -18701
rect -9150 -18735 -9144 -18701
rect -9190 -18773 -9144 -18735
rect -9190 -18807 -9184 -18773
rect -9150 -18807 -9144 -18773
rect -9190 -18838 -9144 -18807
rect -8172 -18303 -8166 -18272
rect -8132 -18272 -8118 -18269
rect -7158 -18269 -7098 -17989
rect -6140 -17989 -6130 -17984
rect -6096 -17984 -6090 -17955
rect -5118 -17485 -5112 -17451
rect -5078 -17485 -5072 -17451
rect -4108 -17451 -4048 -17171
rect -3086 -17171 -3076 -17166
rect -3042 -17166 -3036 -17137
rect -2064 -16667 -2058 -16644
rect -2024 -16644 -2006 -16633
rect -1050 -16633 -990 -16353
rect -28 -16353 -22 -16319
rect 12 -16353 18 -16319
rect -28 -16354 18 -16353
rect -758 -16422 -270 -16416
rect -758 -16456 -711 -16422
rect -677 -16456 -639 -16422
rect -605 -16456 -567 -16422
rect -533 -16456 -495 -16422
rect -461 -16456 -423 -16422
rect -389 -16456 -351 -16422
rect -317 -16456 -270 -16422
rect -758 -16462 -270 -16456
rect -556 -16524 -496 -16462
rect -758 -16530 -270 -16524
rect -758 -16564 -711 -16530
rect -677 -16564 -639 -16530
rect -605 -16564 -567 -16530
rect -533 -16564 -495 -16530
rect -461 -16564 -423 -16530
rect -389 -16564 -351 -16530
rect -317 -16564 -270 -16530
rect -758 -16570 -270 -16564
rect -1050 -16640 -1040 -16633
rect -2024 -16667 -2018 -16644
rect -2064 -16705 -2018 -16667
rect -2064 -16739 -2058 -16705
rect -2024 -16739 -2018 -16705
rect -2064 -16777 -2018 -16739
rect -2064 -16811 -2058 -16777
rect -2024 -16811 -2018 -16777
rect -2064 -16849 -2018 -16811
rect -2064 -16883 -2058 -16849
rect -2024 -16883 -2018 -16849
rect -2064 -16921 -2018 -16883
rect -2064 -16955 -2058 -16921
rect -2024 -16955 -2018 -16921
rect -2064 -16993 -2018 -16955
rect -2064 -17027 -2058 -16993
rect -2024 -17027 -2018 -16993
rect -2064 -17065 -2018 -17027
rect -2064 -17099 -2058 -17065
rect -2024 -17099 -2018 -17065
rect -2064 -17137 -2018 -17099
rect -2064 -17166 -2058 -17137
rect -3042 -17171 -3026 -17166
rect -3812 -17240 -3324 -17234
rect -3812 -17274 -3765 -17240
rect -3731 -17274 -3693 -17240
rect -3659 -17274 -3621 -17240
rect -3587 -17274 -3549 -17240
rect -3515 -17274 -3477 -17240
rect -3443 -17274 -3405 -17240
rect -3371 -17274 -3324 -17240
rect -3812 -17280 -3324 -17274
rect -3608 -17342 -3548 -17280
rect -3812 -17348 -3324 -17342
rect -3812 -17382 -3765 -17348
rect -3731 -17382 -3693 -17348
rect -3659 -17382 -3621 -17348
rect -3587 -17382 -3549 -17348
rect -3515 -17382 -3477 -17348
rect -3443 -17382 -3405 -17348
rect -3371 -17382 -3324 -17348
rect -3812 -17388 -3324 -17382
rect -4108 -17456 -4094 -17451
rect -5118 -17523 -5072 -17485
rect -5118 -17557 -5112 -17523
rect -5078 -17557 -5072 -17523
rect -5118 -17595 -5072 -17557
rect -5118 -17629 -5112 -17595
rect -5078 -17629 -5072 -17595
rect -5118 -17667 -5072 -17629
rect -5118 -17701 -5112 -17667
rect -5078 -17701 -5072 -17667
rect -5118 -17739 -5072 -17701
rect -5118 -17773 -5112 -17739
rect -5078 -17773 -5072 -17739
rect -5118 -17811 -5072 -17773
rect -5118 -17845 -5112 -17811
rect -5078 -17845 -5072 -17811
rect -5118 -17883 -5072 -17845
rect -5118 -17917 -5112 -17883
rect -5078 -17917 -5072 -17883
rect -5118 -17955 -5072 -17917
rect -5118 -17976 -5112 -17955
rect -6096 -17989 -6080 -17984
rect -6866 -18058 -6378 -18052
rect -6866 -18092 -6819 -18058
rect -6785 -18092 -6747 -18058
rect -6713 -18092 -6675 -18058
rect -6641 -18092 -6603 -18058
rect -6569 -18092 -6531 -18058
rect -6497 -18092 -6459 -18058
rect -6425 -18092 -6378 -18058
rect -6866 -18098 -6378 -18092
rect -6654 -18160 -6594 -18098
rect -6866 -18166 -6378 -18160
rect -6866 -18200 -6819 -18166
rect -6785 -18200 -6747 -18166
rect -6713 -18200 -6675 -18166
rect -6641 -18200 -6603 -18166
rect -6569 -18200 -6531 -18166
rect -6497 -18200 -6459 -18166
rect -6425 -18200 -6378 -18166
rect -6866 -18206 -6378 -18200
rect -7158 -18270 -7148 -18269
rect -8132 -18303 -8126 -18272
rect -8172 -18341 -8126 -18303
rect -8172 -18375 -8166 -18341
rect -8132 -18375 -8126 -18341
rect -8172 -18413 -8126 -18375
rect -8172 -18447 -8166 -18413
rect -8132 -18447 -8126 -18413
rect -8172 -18485 -8126 -18447
rect -8172 -18519 -8166 -18485
rect -8132 -18519 -8126 -18485
rect -8172 -18557 -8126 -18519
rect -8172 -18591 -8166 -18557
rect -8132 -18591 -8126 -18557
rect -8172 -18629 -8126 -18591
rect -8172 -18663 -8166 -18629
rect -8132 -18663 -8126 -18629
rect -8172 -18701 -8126 -18663
rect -8172 -18735 -8166 -18701
rect -8132 -18735 -8126 -18701
rect -8172 -18773 -8126 -18735
rect -8172 -18807 -8166 -18773
rect -8132 -18807 -8126 -18773
rect -7154 -18303 -7148 -18270
rect -7114 -18270 -7098 -18269
rect -6140 -18269 -6080 -17989
rect -5120 -17989 -5112 -17976
rect -5078 -17976 -5072 -17955
rect -4100 -17485 -4094 -17456
rect -4060 -17456 -4048 -17451
rect -3086 -17451 -3026 -17171
rect -2066 -17171 -2058 -17166
rect -2024 -17166 -2018 -17137
rect -1046 -16667 -1040 -16640
rect -1006 -16640 -990 -16633
rect -28 -16633 32 -16354
rect -1006 -16667 -1000 -16640
rect -1046 -16705 -1000 -16667
rect -1046 -16739 -1040 -16705
rect -1006 -16739 -1000 -16705
rect -1046 -16777 -1000 -16739
rect -1046 -16811 -1040 -16777
rect -1006 -16811 -1000 -16777
rect -1046 -16849 -1000 -16811
rect -1046 -16883 -1040 -16849
rect -1006 -16883 -1000 -16849
rect -1046 -16921 -1000 -16883
rect -1046 -16955 -1040 -16921
rect -1006 -16955 -1000 -16921
rect -1046 -16993 -1000 -16955
rect -1046 -17027 -1040 -16993
rect -1006 -17027 -1000 -16993
rect -1046 -17065 -1000 -17027
rect -1046 -17099 -1040 -17065
rect -1006 -17099 -1000 -17065
rect -1046 -17137 -1000 -17099
rect -1046 -17162 -1040 -17137
rect -2024 -17171 -2006 -17166
rect -2794 -17240 -2306 -17234
rect -2794 -17274 -2747 -17240
rect -2713 -17274 -2675 -17240
rect -2641 -17274 -2603 -17240
rect -2569 -17274 -2531 -17240
rect -2497 -17274 -2459 -17240
rect -2425 -17274 -2387 -17240
rect -2353 -17274 -2306 -17240
rect -2794 -17280 -2306 -17274
rect -2586 -17342 -2526 -17280
rect -2794 -17348 -2306 -17342
rect -2794 -17382 -2747 -17348
rect -2713 -17382 -2675 -17348
rect -2641 -17382 -2603 -17348
rect -2569 -17382 -2531 -17348
rect -2497 -17382 -2459 -17348
rect -2425 -17382 -2387 -17348
rect -2353 -17382 -2306 -17348
rect -2794 -17388 -2306 -17382
rect -3086 -17456 -3076 -17451
rect -4060 -17485 -4054 -17456
rect -4100 -17523 -4054 -17485
rect -4100 -17557 -4094 -17523
rect -4060 -17557 -4054 -17523
rect -4100 -17595 -4054 -17557
rect -4100 -17629 -4094 -17595
rect -4060 -17629 -4054 -17595
rect -4100 -17667 -4054 -17629
rect -4100 -17701 -4094 -17667
rect -4060 -17701 -4054 -17667
rect -4100 -17739 -4054 -17701
rect -4100 -17773 -4094 -17739
rect -4060 -17773 -4054 -17739
rect -4100 -17811 -4054 -17773
rect -4100 -17845 -4094 -17811
rect -4060 -17845 -4054 -17811
rect -4100 -17883 -4054 -17845
rect -4100 -17917 -4094 -17883
rect -4060 -17917 -4054 -17883
rect -4100 -17955 -4054 -17917
rect -5078 -17989 -5060 -17976
rect -4100 -17984 -4094 -17955
rect -5848 -18058 -5360 -18052
rect -5848 -18092 -5801 -18058
rect -5767 -18092 -5729 -18058
rect -5695 -18092 -5657 -18058
rect -5623 -18092 -5585 -18058
rect -5551 -18092 -5513 -18058
rect -5479 -18092 -5441 -18058
rect -5407 -18092 -5360 -18058
rect -5848 -18098 -5360 -18092
rect -5652 -18160 -5592 -18098
rect -5848 -18166 -5360 -18160
rect -5848 -18200 -5801 -18166
rect -5767 -18200 -5729 -18166
rect -5695 -18200 -5657 -18166
rect -5623 -18200 -5585 -18166
rect -5551 -18200 -5513 -18166
rect -5479 -18200 -5441 -18166
rect -5407 -18200 -5360 -18166
rect -5848 -18206 -5360 -18200
rect -5120 -18266 -5060 -17989
rect -4108 -17989 -4094 -17984
rect -4060 -17984 -4054 -17955
rect -3082 -17485 -3076 -17456
rect -3042 -17456 -3026 -17451
rect -2066 -17451 -2006 -17171
rect -1050 -17171 -1040 -17162
rect -1006 -17162 -1000 -17137
rect -28 -16667 -22 -16633
rect 12 -16644 32 -16633
rect 12 -16667 18 -16644
rect -28 -16705 18 -16667
rect -28 -16739 -22 -16705
rect 12 -16739 18 -16705
rect -28 -16777 18 -16739
rect -28 -16811 -22 -16777
rect 12 -16811 18 -16777
rect -28 -16849 18 -16811
rect -28 -16883 -22 -16849
rect 12 -16883 18 -16849
rect -28 -16921 18 -16883
rect -28 -16955 -22 -16921
rect 12 -16955 18 -16921
rect -28 -16993 18 -16955
rect -28 -17027 -22 -16993
rect 12 -17027 18 -16993
rect -28 -17065 18 -17027
rect -28 -17099 -22 -17065
rect 12 -17099 18 -17065
rect -28 -17137 18 -17099
rect -1006 -17171 -990 -17162
rect -1776 -17240 -1288 -17234
rect -1776 -17274 -1729 -17240
rect -1695 -17274 -1657 -17240
rect -1623 -17274 -1585 -17240
rect -1551 -17274 -1513 -17240
rect -1479 -17274 -1441 -17240
rect -1407 -17274 -1369 -17240
rect -1335 -17274 -1288 -17240
rect -1776 -17280 -1288 -17274
rect -1574 -17342 -1514 -17280
rect -1776 -17348 -1288 -17342
rect -1776 -17382 -1729 -17348
rect -1695 -17382 -1657 -17348
rect -1623 -17382 -1585 -17348
rect -1551 -17382 -1513 -17348
rect -1479 -17382 -1441 -17348
rect -1407 -17382 -1369 -17348
rect -1335 -17382 -1288 -17348
rect -1776 -17388 -1288 -17382
rect -2066 -17456 -2058 -17451
rect -3042 -17485 -3036 -17456
rect -3082 -17523 -3036 -17485
rect -3082 -17557 -3076 -17523
rect -3042 -17557 -3036 -17523
rect -3082 -17595 -3036 -17557
rect -3082 -17629 -3076 -17595
rect -3042 -17629 -3036 -17595
rect -3082 -17667 -3036 -17629
rect -3082 -17701 -3076 -17667
rect -3042 -17701 -3036 -17667
rect -3082 -17739 -3036 -17701
rect -3082 -17773 -3076 -17739
rect -3042 -17773 -3036 -17739
rect -3082 -17811 -3036 -17773
rect -3082 -17845 -3076 -17811
rect -3042 -17845 -3036 -17811
rect -3082 -17883 -3036 -17845
rect -3082 -17917 -3076 -17883
rect -3042 -17917 -3036 -17883
rect -3082 -17955 -3036 -17917
rect -3082 -17984 -3076 -17955
rect -4060 -17989 -4048 -17984
rect -4830 -18058 -4342 -18052
rect -4830 -18092 -4783 -18058
rect -4749 -18092 -4711 -18058
rect -4677 -18092 -4639 -18058
rect -4605 -18092 -4567 -18058
rect -4533 -18092 -4495 -18058
rect -4461 -18092 -4423 -18058
rect -4389 -18092 -4342 -18058
rect -4830 -18098 -4342 -18092
rect -4622 -18160 -4562 -18098
rect -4830 -18166 -4342 -18160
rect -4830 -18200 -4783 -18166
rect -4749 -18200 -4711 -18166
rect -4677 -18200 -4639 -18166
rect -4605 -18200 -4567 -18166
rect -4533 -18200 -4495 -18166
rect -4461 -18200 -4423 -18166
rect -4389 -18200 -4342 -18166
rect -4830 -18206 -4342 -18200
rect -7114 -18303 -7108 -18270
rect -6140 -18274 -6130 -18269
rect -7154 -18341 -7108 -18303
rect -7154 -18375 -7148 -18341
rect -7114 -18375 -7108 -18341
rect -7154 -18413 -7108 -18375
rect -7154 -18447 -7148 -18413
rect -7114 -18447 -7108 -18413
rect -7154 -18485 -7108 -18447
rect -7154 -18519 -7148 -18485
rect -7114 -18519 -7108 -18485
rect -7154 -18557 -7108 -18519
rect -7154 -18591 -7148 -18557
rect -7114 -18591 -7108 -18557
rect -7154 -18629 -7108 -18591
rect -7154 -18663 -7148 -18629
rect -7114 -18663 -7108 -18629
rect -7154 -18701 -7108 -18663
rect -7154 -18735 -7148 -18701
rect -7114 -18735 -7108 -18701
rect -7154 -18773 -7108 -18735
rect -7154 -18780 -7148 -18773
rect -8172 -18838 -8126 -18807
rect -7164 -18807 -7148 -18780
rect -7114 -18780 -7108 -18773
rect -6136 -18303 -6130 -18274
rect -6096 -18274 -6080 -18269
rect -5118 -18269 -5072 -18266
rect -6096 -18303 -6090 -18274
rect -6136 -18341 -6090 -18303
rect -6136 -18375 -6130 -18341
rect -6096 -18375 -6090 -18341
rect -6136 -18413 -6090 -18375
rect -6136 -18447 -6130 -18413
rect -6096 -18447 -6090 -18413
rect -6136 -18485 -6090 -18447
rect -6136 -18519 -6130 -18485
rect -6096 -18519 -6090 -18485
rect -6136 -18557 -6090 -18519
rect -6136 -18591 -6130 -18557
rect -6096 -18591 -6090 -18557
rect -6136 -18629 -6090 -18591
rect -6136 -18663 -6130 -18629
rect -6096 -18663 -6090 -18629
rect -6136 -18701 -6090 -18663
rect -6136 -18735 -6130 -18701
rect -6096 -18735 -6090 -18701
rect -6136 -18773 -6090 -18735
rect -7114 -18807 -7104 -18780
rect -12328 -18893 -12289 -18859
rect -12255 -18893 -12216 -18859
rect -12328 -18931 -12216 -18893
rect -8902 -18876 -8414 -18870
rect -8902 -18910 -8855 -18876
rect -8821 -18910 -8783 -18876
rect -8749 -18910 -8711 -18876
rect -8677 -18910 -8639 -18876
rect -8605 -18910 -8567 -18876
rect -8533 -18910 -8495 -18876
rect -8461 -18910 -8414 -18876
rect -8902 -18916 -8414 -18910
rect -7884 -18876 -7396 -18870
rect -7884 -18910 -7837 -18876
rect -7803 -18910 -7765 -18876
rect -7731 -18910 -7693 -18876
rect -7659 -18910 -7621 -18876
rect -7587 -18910 -7549 -18876
rect -7515 -18910 -7477 -18876
rect -7443 -18910 -7396 -18876
rect -7884 -18916 -7672 -18910
rect -7612 -18916 -7396 -18910
rect -12328 -18965 -12289 -18931
rect -12255 -18965 -12216 -18931
rect -12328 -19003 -12216 -18965
rect -12328 -19037 -12289 -19003
rect -12255 -19037 -12216 -19003
rect -12328 -19075 -12216 -19037
rect -7164 -19000 -7104 -18807
rect -6136 -18807 -6130 -18773
rect -6096 -18807 -6090 -18773
rect -5118 -18303 -5112 -18269
rect -5078 -18303 -5072 -18269
rect -4108 -18269 -4048 -17989
rect -3086 -17989 -3076 -17984
rect -3042 -17984 -3036 -17955
rect -2064 -17485 -2058 -17456
rect -2024 -17456 -2006 -17451
rect -1050 -17451 -990 -17171
rect -28 -17171 -22 -17137
rect 12 -17166 18 -17137
rect 12 -17171 32 -17166
rect -758 -17240 -270 -17234
rect -758 -17274 -711 -17240
rect -677 -17274 -639 -17240
rect -605 -17274 -567 -17240
rect -533 -17274 -495 -17240
rect -461 -17274 -423 -17240
rect -389 -17274 -351 -17240
rect -317 -17274 -270 -17240
rect -758 -17280 -270 -17274
rect -554 -17342 -494 -17280
rect -758 -17348 -270 -17342
rect -758 -17382 -711 -17348
rect -677 -17382 -639 -17348
rect -605 -17382 -567 -17348
rect -533 -17382 -495 -17348
rect -461 -17382 -423 -17348
rect -389 -17382 -351 -17348
rect -317 -17382 -270 -17348
rect -758 -17388 -270 -17382
rect -1050 -17452 -1040 -17451
rect -2024 -17485 -2018 -17456
rect -2064 -17523 -2018 -17485
rect -2064 -17557 -2058 -17523
rect -2024 -17557 -2018 -17523
rect -2064 -17595 -2018 -17557
rect -2064 -17629 -2058 -17595
rect -2024 -17629 -2018 -17595
rect -2064 -17667 -2018 -17629
rect -2064 -17701 -2058 -17667
rect -2024 -17701 -2018 -17667
rect -2064 -17739 -2018 -17701
rect -2064 -17773 -2058 -17739
rect -2024 -17773 -2018 -17739
rect -2064 -17811 -2018 -17773
rect -2064 -17845 -2058 -17811
rect -2024 -17845 -2018 -17811
rect -2064 -17883 -2018 -17845
rect -2064 -17917 -2058 -17883
rect -2024 -17917 -2018 -17883
rect -2064 -17955 -2018 -17917
rect -2064 -17984 -2058 -17955
rect -3042 -17989 -3026 -17984
rect -3812 -18058 -3324 -18052
rect -3812 -18092 -3765 -18058
rect -3731 -18092 -3693 -18058
rect -3659 -18092 -3621 -18058
rect -3587 -18092 -3549 -18058
rect -3515 -18092 -3477 -18058
rect -3443 -18092 -3405 -18058
rect -3371 -18092 -3324 -18058
rect -3812 -18098 -3324 -18092
rect -3606 -18160 -3546 -18098
rect -3812 -18166 -3324 -18160
rect -3812 -18200 -3765 -18166
rect -3731 -18200 -3693 -18166
rect -3659 -18200 -3621 -18166
rect -3587 -18200 -3549 -18166
rect -3515 -18200 -3477 -18166
rect -3443 -18200 -3405 -18166
rect -3371 -18200 -3324 -18166
rect -3812 -18206 -3324 -18200
rect -4108 -18274 -4094 -18269
rect -5118 -18341 -5072 -18303
rect -5118 -18375 -5112 -18341
rect -5078 -18375 -5072 -18341
rect -5118 -18413 -5072 -18375
rect -5118 -18447 -5112 -18413
rect -5078 -18447 -5072 -18413
rect -5118 -18485 -5072 -18447
rect -5118 -18519 -5112 -18485
rect -5078 -18519 -5072 -18485
rect -5118 -18557 -5072 -18519
rect -5118 -18591 -5112 -18557
rect -5078 -18591 -5072 -18557
rect -5118 -18629 -5072 -18591
rect -5118 -18663 -5112 -18629
rect -5078 -18663 -5072 -18629
rect -5118 -18701 -5072 -18663
rect -5118 -18735 -5112 -18701
rect -5078 -18735 -5072 -18701
rect -5118 -18773 -5072 -18735
rect -5118 -18778 -5112 -18773
rect -6136 -18838 -6090 -18807
rect -5126 -18807 -5112 -18778
rect -5078 -18778 -5072 -18773
rect -4100 -18303 -4094 -18274
rect -4060 -18274 -4048 -18269
rect -3086 -18269 -3026 -17989
rect -2066 -17989 -2058 -17984
rect -2024 -17984 -2018 -17955
rect -1046 -17485 -1040 -17452
rect -1006 -17452 -990 -17451
rect -28 -17451 32 -17171
rect -1006 -17485 -1000 -17452
rect -1046 -17523 -1000 -17485
rect -1046 -17557 -1040 -17523
rect -1006 -17557 -1000 -17523
rect -1046 -17595 -1000 -17557
rect -1046 -17629 -1040 -17595
rect -1006 -17629 -1000 -17595
rect -1046 -17667 -1000 -17629
rect -1046 -17701 -1040 -17667
rect -1006 -17701 -1000 -17667
rect -1046 -17739 -1000 -17701
rect -1046 -17773 -1040 -17739
rect -1006 -17773 -1000 -17739
rect -1046 -17811 -1000 -17773
rect -1046 -17845 -1040 -17811
rect -1006 -17845 -1000 -17811
rect -1046 -17883 -1000 -17845
rect -1046 -17917 -1040 -17883
rect -1006 -17917 -1000 -17883
rect -1046 -17955 -1000 -17917
rect -1046 -17980 -1040 -17955
rect -2024 -17989 -2006 -17984
rect -2794 -18058 -2306 -18052
rect -2794 -18092 -2747 -18058
rect -2713 -18092 -2675 -18058
rect -2641 -18092 -2603 -18058
rect -2569 -18092 -2531 -18058
rect -2497 -18092 -2459 -18058
rect -2425 -18092 -2387 -18058
rect -2353 -18092 -2306 -18058
rect -2794 -18098 -2306 -18092
rect -2584 -18160 -2524 -18098
rect -2794 -18166 -2306 -18160
rect -2794 -18200 -2747 -18166
rect -2713 -18200 -2675 -18166
rect -2641 -18200 -2603 -18166
rect -2569 -18200 -2531 -18166
rect -2497 -18200 -2459 -18166
rect -2425 -18200 -2387 -18166
rect -2353 -18200 -2306 -18166
rect -2794 -18206 -2306 -18200
rect -3086 -18274 -3076 -18269
rect -4060 -18303 -4054 -18274
rect -4100 -18341 -4054 -18303
rect -4100 -18375 -4094 -18341
rect -4060 -18375 -4054 -18341
rect -4100 -18413 -4054 -18375
rect -4100 -18447 -4094 -18413
rect -4060 -18447 -4054 -18413
rect -4100 -18485 -4054 -18447
rect -4100 -18519 -4094 -18485
rect -4060 -18519 -4054 -18485
rect -4100 -18557 -4054 -18519
rect -4100 -18591 -4094 -18557
rect -4060 -18591 -4054 -18557
rect -4100 -18629 -4054 -18591
rect -4100 -18663 -4094 -18629
rect -4060 -18663 -4054 -18629
rect -4100 -18701 -4054 -18663
rect -4100 -18735 -4094 -18701
rect -4060 -18735 -4054 -18701
rect -4100 -18773 -4054 -18735
rect -5078 -18807 -5066 -18778
rect -6866 -18876 -6378 -18870
rect -6866 -18910 -6819 -18876
rect -6785 -18910 -6747 -18876
rect -6713 -18910 -6675 -18876
rect -6641 -18910 -6603 -18876
rect -6569 -18910 -6531 -18876
rect -6497 -18910 -6459 -18876
rect -6425 -18910 -6378 -18876
rect -6866 -18916 -6378 -18910
rect -5848 -18876 -5360 -18870
rect -5848 -18910 -5801 -18876
rect -5767 -18910 -5729 -18876
rect -5695 -18910 -5657 -18876
rect -5623 -18910 -5585 -18876
rect -5551 -18910 -5513 -18876
rect -5479 -18910 -5441 -18876
rect -5407 -18910 -5360 -18876
rect -5848 -18916 -5360 -18910
rect -5126 -19000 -5066 -18807
rect -4100 -18807 -4094 -18773
rect -4060 -18807 -4054 -18773
rect -3082 -18303 -3076 -18274
rect -3042 -18274 -3026 -18269
rect -2066 -18269 -2006 -17989
rect -1050 -17989 -1040 -17980
rect -1006 -17980 -1000 -17955
rect -28 -17485 -22 -17451
rect 12 -17456 32 -17451
rect 12 -17485 18 -17456
rect -28 -17523 18 -17485
rect -28 -17557 -22 -17523
rect 12 -17557 18 -17523
rect -28 -17595 18 -17557
rect -28 -17629 -22 -17595
rect 12 -17629 18 -17595
rect -28 -17667 18 -17629
rect -28 -17701 -22 -17667
rect 12 -17701 18 -17667
rect -28 -17739 18 -17701
rect -28 -17773 -22 -17739
rect 12 -17773 18 -17739
rect -28 -17811 18 -17773
rect -28 -17845 -22 -17811
rect 12 -17845 18 -17811
rect -28 -17883 18 -17845
rect -28 -17917 -22 -17883
rect 12 -17917 18 -17883
rect -28 -17955 18 -17917
rect -1006 -17989 -990 -17980
rect -1776 -18058 -1288 -18052
rect -1776 -18092 -1729 -18058
rect -1695 -18092 -1657 -18058
rect -1623 -18092 -1585 -18058
rect -1551 -18092 -1513 -18058
rect -1479 -18092 -1441 -18058
rect -1407 -18092 -1369 -18058
rect -1335 -18092 -1288 -18058
rect -1776 -18098 -1288 -18092
rect -1572 -18160 -1512 -18098
rect -1776 -18166 -1288 -18160
rect -1776 -18200 -1729 -18166
rect -1695 -18200 -1657 -18166
rect -1623 -18200 -1585 -18166
rect -1551 -18200 -1513 -18166
rect -1479 -18200 -1441 -18166
rect -1407 -18200 -1369 -18166
rect -1335 -18200 -1288 -18166
rect -1776 -18206 -1288 -18200
rect -2066 -18274 -2058 -18269
rect -3042 -18303 -3036 -18274
rect -3082 -18341 -3036 -18303
rect -3082 -18375 -3076 -18341
rect -3042 -18375 -3036 -18341
rect -3082 -18413 -3036 -18375
rect -3082 -18447 -3076 -18413
rect -3042 -18447 -3036 -18413
rect -3082 -18485 -3036 -18447
rect -3082 -18519 -3076 -18485
rect -3042 -18519 -3036 -18485
rect -3082 -18557 -3036 -18519
rect -3082 -18591 -3076 -18557
rect -3042 -18591 -3036 -18557
rect -3082 -18629 -3036 -18591
rect -3082 -18663 -3076 -18629
rect -3042 -18663 -3036 -18629
rect -3082 -18701 -3036 -18663
rect -3082 -18735 -3076 -18701
rect -3042 -18735 -3036 -18701
rect -3082 -18773 -3036 -18735
rect -3082 -18782 -3076 -18773
rect -4100 -18838 -4054 -18807
rect -3090 -18807 -3076 -18782
rect -3042 -18782 -3036 -18773
rect -2064 -18303 -2058 -18274
rect -2024 -18274 -2006 -18269
rect -1050 -18269 -990 -17989
rect -28 -17989 -22 -17955
rect 12 -17984 18 -17955
rect 12 -17989 32 -17984
rect -758 -18058 -270 -18052
rect -758 -18092 -711 -18058
rect -677 -18092 -639 -18058
rect -605 -18092 -567 -18058
rect -533 -18092 -495 -18058
rect -461 -18092 -423 -18058
rect -389 -18092 -351 -18058
rect -317 -18092 -270 -18058
rect -758 -18098 -270 -18092
rect -552 -18160 -492 -18098
rect -758 -18166 -270 -18160
rect -758 -18200 -711 -18166
rect -677 -18200 -639 -18166
rect -605 -18200 -567 -18166
rect -533 -18200 -495 -18166
rect -461 -18200 -423 -18166
rect -389 -18200 -351 -18166
rect -317 -18200 -270 -18166
rect -758 -18206 -270 -18200
rect -1050 -18270 -1040 -18269
rect -2024 -18303 -2018 -18274
rect -2064 -18341 -2018 -18303
rect -2064 -18375 -2058 -18341
rect -2024 -18375 -2018 -18341
rect -2064 -18413 -2018 -18375
rect -2064 -18447 -2058 -18413
rect -2024 -18447 -2018 -18413
rect -2064 -18485 -2018 -18447
rect -2064 -18519 -2058 -18485
rect -2024 -18519 -2018 -18485
rect -2064 -18557 -2018 -18519
rect -2064 -18591 -2058 -18557
rect -2024 -18591 -2018 -18557
rect -2064 -18629 -2018 -18591
rect -2064 -18663 -2058 -18629
rect -2024 -18663 -2018 -18629
rect -2064 -18701 -2018 -18663
rect -2064 -18735 -2058 -18701
rect -2024 -18735 -2018 -18701
rect -2064 -18773 -2018 -18735
rect -3042 -18807 -3030 -18782
rect -4830 -18876 -4342 -18870
rect -4830 -18910 -4783 -18876
rect -4749 -18910 -4711 -18876
rect -4677 -18910 -4639 -18876
rect -4605 -18910 -4567 -18876
rect -4533 -18910 -4495 -18876
rect -4461 -18910 -4423 -18876
rect -4389 -18910 -4342 -18876
rect -4830 -18916 -4342 -18910
rect -3812 -18876 -3324 -18870
rect -3812 -18910 -3765 -18876
rect -3731 -18910 -3693 -18876
rect -3659 -18910 -3621 -18876
rect -3587 -18910 -3549 -18876
rect -3515 -18910 -3477 -18876
rect -3443 -18910 -3405 -18876
rect -3371 -18910 -3324 -18876
rect -3812 -18916 -3324 -18910
rect -3090 -19000 -3030 -18807
rect -2064 -18807 -2058 -18773
rect -2024 -18807 -2018 -18773
rect -1046 -18303 -1040 -18270
rect -1006 -18270 -990 -18269
rect -28 -18269 32 -17989
rect -1006 -18303 -1000 -18270
rect -1046 -18341 -1000 -18303
rect -1046 -18375 -1040 -18341
rect -1006 -18375 -1000 -18341
rect -1046 -18413 -1000 -18375
rect -1046 -18447 -1040 -18413
rect -1006 -18447 -1000 -18413
rect -1046 -18485 -1000 -18447
rect -1046 -18519 -1040 -18485
rect -1006 -18519 -1000 -18485
rect -1046 -18557 -1000 -18519
rect -1046 -18591 -1040 -18557
rect -1006 -18591 -1000 -18557
rect -1046 -18629 -1000 -18591
rect -1046 -18663 -1040 -18629
rect -1006 -18663 -1000 -18629
rect -1046 -18701 -1000 -18663
rect -1046 -18735 -1040 -18701
rect -1006 -18735 -1000 -18701
rect -1046 -18773 -1000 -18735
rect -28 -18303 -22 -18269
rect 12 -18274 32 -18269
rect 12 -18303 18 -18274
rect -28 -18341 18 -18303
rect -28 -18375 -22 -18341
rect 12 -18375 18 -18341
rect -28 -18413 18 -18375
rect -28 -18447 -22 -18413
rect 12 -18447 18 -18413
rect -28 -18485 18 -18447
rect -28 -18519 -22 -18485
rect 12 -18519 18 -18485
rect -28 -18557 18 -18519
rect -28 -18591 -22 -18557
rect 12 -18591 18 -18557
rect -28 -18629 18 -18591
rect -28 -18663 -22 -18629
rect 12 -18663 18 -18629
rect -28 -18701 18 -18663
rect -28 -18735 -22 -18701
rect 12 -18735 18 -18701
rect -28 -18772 18 -18735
rect -1046 -18784 -1040 -18773
rect -2064 -18838 -2018 -18807
rect -1054 -18807 -1040 -18784
rect -1006 -18784 -1000 -18773
rect -34 -18773 26 -18772
rect -1006 -18807 -994 -18784
rect -2794 -18876 -2306 -18870
rect -2794 -18910 -2747 -18876
rect -2713 -18910 -2675 -18876
rect -2641 -18910 -2603 -18876
rect -2569 -18910 -2531 -18876
rect -2497 -18910 -2459 -18876
rect -2425 -18910 -2387 -18876
rect -2353 -18910 -2306 -18876
rect -2794 -18916 -2306 -18910
rect -1776 -18876 -1288 -18870
rect -1776 -18910 -1729 -18876
rect -1695 -18910 -1657 -18876
rect -1623 -18910 -1585 -18876
rect -1551 -18910 -1513 -18876
rect -1479 -18910 -1441 -18876
rect -1407 -18910 -1369 -18876
rect -1335 -18910 -1288 -18876
rect -1776 -18916 -1288 -18910
rect -1054 -19000 -994 -18807
rect -34 -18807 -22 -18773
rect 12 -18807 26 -18773
rect -758 -18876 -270 -18870
rect -758 -18910 -711 -18876
rect -677 -18910 -639 -18876
rect -605 -18910 -567 -18876
rect -533 -18910 -495 -18876
rect -461 -18910 -423 -18876
rect -389 -18910 -351 -18876
rect -317 -18910 -270 -18876
rect -758 -18916 -270 -18910
rect -540 -19000 -480 -18916
rect -34 -19000 26 -18807
rect 952 -18862 1012 -18852
rect -7164 -19060 26 -19000
rect 690 -18892 750 -18866
rect 690 -18944 694 -18892
rect 746 -18944 750 -18892
rect -12328 -19109 -12289 -19075
rect -12255 -19109 -12216 -19075
rect -12328 -19147 -12216 -19109
rect -12328 -19181 -12289 -19147
rect -12255 -19181 -12216 -19147
rect -12328 -19219 -12216 -19181
rect -12328 -19253 -12289 -19219
rect -12255 -19253 -12216 -19219
rect -12328 -19291 -12216 -19253
rect -12328 -19325 -12289 -19291
rect -12255 -19325 -12216 -19291
rect -12328 -19363 -12216 -19325
rect -12328 -19397 -12289 -19363
rect -12255 -19397 -12216 -19363
rect -12328 -19435 -12216 -19397
rect -12328 -19469 -12289 -19435
rect -12255 -19469 -12216 -19435
rect -12328 -19507 -12216 -19469
rect -12328 -19541 -12289 -19507
rect -12255 -19541 -12216 -19507
rect -12328 -19579 -12216 -19541
rect -12328 -19613 -12289 -19579
rect -12255 -19613 -12216 -19579
rect -12328 -19651 -12216 -19613
rect -12328 -19685 -12289 -19651
rect -12255 -19685 -12216 -19651
rect -12328 -19723 -12216 -19685
rect -12328 -19757 -12289 -19723
rect -12255 -19757 -12216 -19723
rect -12328 -19795 -12216 -19757
rect -12328 -19829 -12289 -19795
rect -12255 -19829 -12216 -19795
rect -12328 -19867 -12216 -19829
rect -12328 -19901 -12289 -19867
rect -12255 -19901 -12216 -19867
rect -12328 -19939 -12216 -19901
rect -12328 -19973 -12289 -19939
rect -12255 -19973 -12216 -19939
rect -12328 -20011 -12216 -19973
rect -12328 -20045 -12289 -20011
rect -12255 -20045 -12216 -20011
rect -12328 -20083 -12216 -20045
rect -12328 -20117 -12289 -20083
rect -12255 -20117 -12216 -20083
rect -12328 -20155 -12216 -20117
rect -12328 -20189 -12289 -20155
rect -12255 -20189 -12216 -20155
rect -12328 -20227 -12216 -20189
rect -2982 -20164 -2910 -20160
rect -2982 -20216 -2972 -20164
rect -2920 -20216 -2910 -20164
rect -2982 -20220 -2910 -20216
rect -12328 -20261 -12289 -20227
rect -12255 -20261 -12216 -20227
rect -12328 -20299 -12216 -20261
rect -12328 -20333 -12289 -20299
rect -12255 -20333 -12216 -20299
rect -12328 -20371 -12216 -20333
rect -12328 -20405 -12289 -20371
rect -12255 -20405 -12216 -20371
rect -12328 -20443 -12216 -20405
rect -12328 -20477 -12289 -20443
rect -12255 -20477 -12216 -20443
rect -12328 -20515 -12216 -20477
rect -12328 -20549 -12289 -20515
rect -12255 -20549 -12216 -20515
rect -12328 -20587 -12216 -20549
rect -12328 -20621 -12289 -20587
rect -12255 -20621 -12216 -20587
rect -12328 -20659 -12216 -20621
rect -12328 -20693 -12289 -20659
rect -12255 -20693 -12216 -20659
rect -12328 -20731 -12216 -20693
rect -12328 -20765 -12289 -20731
rect -12255 -20765 -12216 -20731
rect -12328 -20803 -12216 -20765
rect -12328 -20837 -12289 -20803
rect -12255 -20837 -12216 -20803
rect -12328 -20875 -12216 -20837
rect -12328 -20909 -12289 -20875
rect -12255 -20909 -12216 -20875
rect -12328 -20947 -12216 -20909
rect -12328 -20981 -12289 -20947
rect -12255 -20981 -12216 -20947
rect -12328 -21019 -12216 -20981
rect -12328 -21053 -12289 -21019
rect -12255 -21053 -12216 -21019
rect -12328 -21091 -12216 -21053
rect -12328 -21125 -12289 -21091
rect -12255 -21125 -12216 -21091
rect -12328 -21163 -12216 -21125
rect -12328 -21197 -12289 -21163
rect -12255 -21197 -12216 -21163
rect -12328 -21235 -12216 -21197
rect -12328 -21269 -12289 -21235
rect -12255 -21269 -12216 -21235
rect -12328 -21307 -12216 -21269
rect -12328 -21341 -12289 -21307
rect -12255 -21341 -12216 -21307
rect -12328 -21379 -12216 -21341
rect -12328 -21413 -12289 -21379
rect -12255 -21413 -12216 -21379
rect -12328 -21451 -12216 -21413
rect -12328 -21485 -12289 -21451
rect -12255 -21485 -12216 -21451
rect -12328 -21523 -12216 -21485
rect -12328 -21557 -12289 -21523
rect -12255 -21557 -12216 -21523
rect -12328 -21595 -12216 -21557
rect -12328 -21629 -12289 -21595
rect -12255 -21629 -12216 -21595
rect -12328 -21667 -12216 -21629
rect -12328 -21701 -12289 -21667
rect -12255 -21701 -12216 -21667
rect -12328 -21739 -12216 -21701
rect -12328 -21773 -12289 -21739
rect -12255 -21773 -12216 -21739
rect -12328 -21811 -12216 -21773
rect -12328 -21845 -12289 -21811
rect -12255 -21845 -12216 -21811
rect -9416 -21614 -8338 -21554
rect -9416 -21812 -9356 -21614
rect -8902 -21703 -8842 -21614
rect -9123 -21709 -8635 -21703
rect -9123 -21743 -9076 -21709
rect -9042 -21743 -9004 -21709
rect -8970 -21743 -8932 -21709
rect -8898 -21743 -8860 -21709
rect -8826 -21743 -8788 -21709
rect -8754 -21743 -8716 -21709
rect -8682 -21743 -8635 -21709
rect -9123 -21749 -8635 -21743
rect -9416 -21838 -9405 -21812
rect -12328 -21883 -12216 -21845
rect -12328 -21917 -12289 -21883
rect -12255 -21917 -12216 -21883
rect -12328 -21955 -12216 -21917
rect -12328 -21989 -12289 -21955
rect -12255 -21989 -12216 -21955
rect -12328 -22027 -12216 -21989
rect -12328 -22061 -12289 -22027
rect -12255 -22061 -12216 -22027
rect -12328 -22099 -12216 -22061
rect -12328 -22133 -12289 -22099
rect -12255 -22133 -12216 -22099
rect -12328 -22171 -12216 -22133
rect -12328 -22205 -12289 -22171
rect -12255 -22205 -12216 -22171
rect -12328 -22243 -12216 -22205
rect -12328 -22277 -12289 -22243
rect -12255 -22277 -12216 -22243
rect -12328 -22315 -12216 -22277
rect -12328 -22349 -12289 -22315
rect -12255 -22349 -12216 -22315
rect -12328 -22387 -12216 -22349
rect -9411 -21846 -9405 -21838
rect -9371 -21838 -9356 -21812
rect -8398 -21812 -8338 -21614
rect -7392 -21604 -7320 -21600
rect -7392 -21656 -7382 -21604
rect -7330 -21656 -7320 -21604
rect -7392 -21660 -7320 -21656
rect -6878 -21614 -5796 -21554
rect -2976 -21556 -2916 -20220
rect -8105 -21709 -7617 -21703
rect -8105 -21743 -8058 -21709
rect -8024 -21743 -7986 -21709
rect -7952 -21743 -7914 -21709
rect -7880 -21743 -7842 -21709
rect -7808 -21743 -7770 -21709
rect -7736 -21743 -7698 -21709
rect -7664 -21743 -7617 -21709
rect -8105 -21749 -7617 -21743
rect -9371 -21846 -9365 -21838
rect -8398 -21842 -8387 -21812
rect -9411 -21884 -9365 -21846
rect -9411 -21918 -9405 -21884
rect -9371 -21918 -9365 -21884
rect -9411 -21956 -9365 -21918
rect -9411 -21990 -9405 -21956
rect -9371 -21990 -9365 -21956
rect -9411 -22028 -9365 -21990
rect -9411 -22062 -9405 -22028
rect -9371 -22062 -9365 -22028
rect -9411 -22100 -9365 -22062
rect -9411 -22134 -9405 -22100
rect -9371 -22134 -9365 -22100
rect -9411 -22172 -9365 -22134
rect -9411 -22206 -9405 -22172
rect -9371 -22206 -9365 -22172
rect -9411 -22244 -9365 -22206
rect -9411 -22278 -9405 -22244
rect -9371 -22278 -9365 -22244
rect -9411 -22316 -9365 -22278
rect -9411 -22350 -9405 -22316
rect -9371 -22350 -9365 -22316
rect -8393 -21846 -8387 -21842
rect -8353 -21842 -8338 -21812
rect -7386 -21812 -7326 -21660
rect -6878 -21703 -6818 -21614
rect -7087 -21709 -6599 -21703
rect -7087 -21743 -7040 -21709
rect -7006 -21743 -6968 -21709
rect -6934 -21743 -6896 -21709
rect -6862 -21743 -6824 -21709
rect -6790 -21743 -6752 -21709
rect -6718 -21743 -6680 -21709
rect -6646 -21743 -6599 -21709
rect -7087 -21749 -6599 -21743
rect -8353 -21846 -8347 -21842
rect -8393 -21884 -8347 -21846
rect -8393 -21918 -8387 -21884
rect -8353 -21918 -8347 -21884
rect -8393 -21956 -8347 -21918
rect -8393 -21990 -8387 -21956
rect -8353 -21990 -8347 -21956
rect -8393 -22028 -8347 -21990
rect -8393 -22062 -8387 -22028
rect -8353 -22062 -8347 -22028
rect -8393 -22100 -8347 -22062
rect -8393 -22134 -8387 -22100
rect -8353 -22134 -8347 -22100
rect -8393 -22172 -8347 -22134
rect -8393 -22206 -8387 -22172
rect -8353 -22206 -8347 -22172
rect -8393 -22244 -8347 -22206
rect -8393 -22278 -8387 -22244
rect -8353 -22278 -8347 -22244
rect -8393 -22316 -8347 -22278
rect -8393 -22324 -8387 -22316
rect -9411 -22381 -9365 -22350
rect -8400 -22350 -8387 -22324
rect -8353 -22324 -8347 -22316
rect -7386 -21846 -7369 -21812
rect -7335 -21846 -7326 -21812
rect -7386 -21884 -7326 -21846
rect -6362 -21812 -6302 -21614
rect -5856 -21703 -5796 -21614
rect -5352 -21604 -5280 -21600
rect -5352 -21656 -5342 -21604
rect -5290 -21656 -5280 -21604
rect -5352 -21660 -5280 -21656
rect -4326 -21616 -2916 -21556
rect -6069 -21709 -5581 -21703
rect -6069 -21743 -6022 -21709
rect -5988 -21743 -5950 -21709
rect -5916 -21743 -5878 -21709
rect -5844 -21743 -5806 -21709
rect -5772 -21743 -5734 -21709
rect -5700 -21743 -5662 -21709
rect -5628 -21743 -5581 -21709
rect -6069 -21749 -5581 -21743
rect -6362 -21846 -6351 -21812
rect -6317 -21846 -6302 -21812
rect -5346 -21812 -5286 -21660
rect -5051 -21709 -4563 -21703
rect -5051 -21743 -5004 -21709
rect -4970 -21743 -4932 -21709
rect -4898 -21743 -4860 -21709
rect -4826 -21743 -4788 -21709
rect -4754 -21743 -4716 -21709
rect -4682 -21743 -4644 -21709
rect -4610 -21743 -4563 -21709
rect -5051 -21749 -4563 -21743
rect -5346 -21838 -5333 -21812
rect -6362 -21850 -6302 -21846
rect -5339 -21846 -5333 -21838
rect -5299 -21838 -5286 -21812
rect -4326 -21812 -4266 -21616
rect -3818 -21703 -3758 -21616
rect -4033 -21709 -3545 -21703
rect -4033 -21743 -3986 -21709
rect -3952 -21743 -3914 -21709
rect -3880 -21743 -3842 -21709
rect -3808 -21743 -3770 -21709
rect -3736 -21743 -3698 -21709
rect -3664 -21743 -3626 -21709
rect -3592 -21743 -3545 -21709
rect -4033 -21749 -3545 -21743
rect -5299 -21846 -5293 -21838
rect -4326 -21846 -4315 -21812
rect -4281 -21846 -4266 -21812
rect -3310 -21812 -3250 -21616
rect -3310 -21840 -3297 -21812
rect -3303 -21846 -3297 -21840
rect -3263 -21840 -3250 -21812
rect -3263 -21846 -3257 -21840
rect -7386 -21918 -7369 -21884
rect -7335 -21918 -7326 -21884
rect -7386 -21956 -7326 -21918
rect -7386 -21990 -7369 -21956
rect -7335 -21990 -7326 -21956
rect -7386 -22028 -7326 -21990
rect -7386 -22062 -7369 -22028
rect -7335 -22062 -7326 -22028
rect -7386 -22100 -7326 -22062
rect -7386 -22134 -7369 -22100
rect -7335 -22134 -7326 -22100
rect -7386 -22172 -7326 -22134
rect -7386 -22206 -7369 -22172
rect -7335 -22206 -7326 -22172
rect -7386 -22244 -7326 -22206
rect -7386 -22278 -7369 -22244
rect -7335 -22278 -7326 -22244
rect -7386 -22316 -7326 -22278
rect -8353 -22350 -8340 -22324
rect -12328 -22421 -12289 -22387
rect -12255 -22421 -12216 -22387
rect -12328 -22459 -12216 -22421
rect -9123 -22419 -8635 -22413
rect -9123 -22453 -9076 -22419
rect -9042 -22453 -9004 -22419
rect -8970 -22453 -8932 -22419
rect -8898 -22453 -8860 -22419
rect -8826 -22453 -8788 -22419
rect -8754 -22453 -8716 -22419
rect -8682 -22453 -8635 -22419
rect -9123 -22459 -8635 -22453
rect -12328 -22493 -12289 -22459
rect -12255 -22493 -12216 -22459
rect -12328 -22531 -12216 -22493
rect -8400 -22504 -8340 -22350
rect -7386 -22350 -7369 -22316
rect -7335 -22350 -7326 -22316
rect -6357 -21884 -6311 -21850
rect -6357 -21918 -6351 -21884
rect -6317 -21918 -6311 -21884
rect -6357 -21956 -6311 -21918
rect -6357 -21990 -6351 -21956
rect -6317 -21990 -6311 -21956
rect -6357 -22028 -6311 -21990
rect -6357 -22062 -6351 -22028
rect -6317 -22062 -6311 -22028
rect -6357 -22100 -6311 -22062
rect -6357 -22134 -6351 -22100
rect -6317 -22134 -6311 -22100
rect -6357 -22172 -6311 -22134
rect -6357 -22206 -6351 -22172
rect -6317 -22206 -6311 -22172
rect -6357 -22244 -6311 -22206
rect -6357 -22278 -6351 -22244
rect -6317 -22278 -6311 -22244
rect -6357 -22316 -6311 -22278
rect -6357 -22328 -6351 -22316
rect -8105 -22419 -7617 -22413
rect -8105 -22453 -8058 -22419
rect -8024 -22453 -7986 -22419
rect -7952 -22453 -7914 -22419
rect -7880 -22453 -7842 -22419
rect -7808 -22453 -7770 -22419
rect -7736 -22453 -7698 -22419
rect -7664 -22453 -7617 -22419
rect -8105 -22459 -7617 -22453
rect -12328 -22565 -12289 -22531
rect -12255 -22565 -12216 -22531
rect -9544 -22508 -9472 -22504
rect -9544 -22560 -9534 -22508
rect -9482 -22560 -9472 -22508
rect -9544 -22564 -9472 -22560
rect -8406 -22508 -8334 -22504
rect -8406 -22560 -8396 -22508
rect -8344 -22560 -8334 -22508
rect -8406 -22564 -8334 -22560
rect -12328 -22603 -12216 -22565
rect -12328 -22637 -12289 -22603
rect -12255 -22637 -12216 -22603
rect -12328 -22675 -12216 -22637
rect -12328 -22709 -12289 -22675
rect -12255 -22709 -12216 -22675
rect -12328 -22747 -12216 -22709
rect -12328 -22781 -12289 -22747
rect -12255 -22781 -12216 -22747
rect -12328 -22819 -12216 -22781
rect -12328 -22853 -12289 -22819
rect -12255 -22853 -12216 -22819
rect -12328 -22891 -12216 -22853
rect -12328 -22925 -12289 -22891
rect -12255 -22925 -12216 -22891
rect -12328 -22963 -12216 -22925
rect -12328 -22997 -12289 -22963
rect -12255 -22997 -12216 -22963
rect -12328 -23035 -12216 -22997
rect -12328 -23069 -12289 -23035
rect -12255 -23069 -12216 -23035
rect -12328 -23107 -12216 -23069
rect -12328 -23141 -12289 -23107
rect -12255 -23141 -12216 -23107
rect -12328 -23179 -12216 -23141
rect -12328 -23213 -12289 -23179
rect -12255 -23213 -12216 -23179
rect -12328 -23251 -12216 -23213
rect -12328 -23285 -12289 -23251
rect -12255 -23285 -12216 -23251
rect -12328 -23323 -12216 -23285
rect -12328 -23357 -12289 -23323
rect -12255 -23357 -12216 -23323
rect -12328 -23395 -12216 -23357
rect -12328 -23429 -12289 -23395
rect -12255 -23429 -12216 -23395
rect -12328 -23467 -12216 -23429
rect -12328 -23501 -12289 -23467
rect -12255 -23501 -12216 -23467
rect -12328 -23539 -12216 -23501
rect -12328 -23573 -12289 -23539
rect -12255 -23573 -12216 -23539
rect -12328 -23611 -12216 -23573
rect -12328 -23645 -12289 -23611
rect -12255 -23645 -12216 -23611
rect -12328 -23683 -12216 -23645
rect -12328 -23717 -12289 -23683
rect -12255 -23717 -12216 -23683
rect -12328 -23755 -12216 -23717
rect -12328 -23789 -12289 -23755
rect -12255 -23789 -12216 -23755
rect -12328 -23827 -12216 -23789
rect -12328 -23861 -12289 -23827
rect -12255 -23861 -12216 -23827
rect -12328 -23899 -12216 -23861
rect -12328 -23933 -12289 -23899
rect -12255 -23933 -12216 -23899
rect -12328 -23971 -12216 -23933
rect -12328 -24005 -12289 -23971
rect -12255 -24005 -12216 -23971
rect -12328 -24043 -12216 -24005
rect -12328 -24077 -12289 -24043
rect -12255 -24077 -12216 -24043
rect -12328 -24115 -12216 -24077
rect -12328 -24149 -12289 -24115
rect -12255 -24149 -12216 -24115
rect -12328 -24187 -12216 -24149
rect -12328 -24221 -12289 -24187
rect -12255 -24221 -12216 -24187
rect -12328 -24259 -12216 -24221
rect -12328 -24293 -12289 -24259
rect -12255 -24293 -12216 -24259
rect -12328 -24331 -12216 -24293
rect -12328 -24365 -12289 -24331
rect -12255 -24365 -12216 -24331
rect -12328 -24403 -12216 -24365
rect -12328 -24437 -12289 -24403
rect -12255 -24437 -12216 -24403
rect -12328 -24475 -12216 -24437
rect -12328 -24509 -12289 -24475
rect -12255 -24509 -12216 -24475
rect -12328 -24547 -12216 -24509
rect -12328 -24581 -12289 -24547
rect -12255 -24581 -12216 -24547
rect -12328 -24619 -12216 -24581
rect -12328 -24653 -12289 -24619
rect -12255 -24653 -12216 -24619
rect -12328 -24691 -12216 -24653
rect -12328 -24725 -12289 -24691
rect -12255 -24725 -12216 -24691
rect -12328 -24763 -12216 -24725
rect -12328 -24797 -12289 -24763
rect -12255 -24797 -12216 -24763
rect -12328 -24835 -12216 -24797
rect -12328 -24869 -12289 -24835
rect -12255 -24869 -12216 -24835
rect -12328 -24907 -12216 -24869
rect -12328 -24941 -12289 -24907
rect -12255 -24941 -12216 -24907
rect -9538 -24926 -9478 -22564
rect -9418 -22780 -8342 -22720
rect -9418 -22925 -9358 -22780
rect -8908 -22816 -8848 -22780
rect -9124 -22822 -8636 -22816
rect -9124 -22856 -9077 -22822
rect -9043 -22856 -9005 -22822
rect -8971 -22856 -8933 -22822
rect -8899 -22856 -8861 -22822
rect -8827 -22856 -8789 -22822
rect -8755 -22856 -8717 -22822
rect -8683 -22856 -8636 -22822
rect -9124 -22862 -8636 -22856
rect -9418 -22959 -9406 -22925
rect -9372 -22959 -9358 -22925
rect -8402 -22925 -8342 -22780
rect -7890 -22816 -7830 -22459
rect -7386 -22600 -7326 -22350
rect -6364 -22350 -6351 -22328
rect -6317 -22328 -6311 -22316
rect -5339 -21884 -5293 -21846
rect -5339 -21918 -5333 -21884
rect -5299 -21918 -5293 -21884
rect -5339 -21956 -5293 -21918
rect -5339 -21990 -5333 -21956
rect -5299 -21990 -5293 -21956
rect -5339 -22028 -5293 -21990
rect -5339 -22062 -5333 -22028
rect -5299 -22062 -5293 -22028
rect -5339 -22100 -5293 -22062
rect -5339 -22134 -5333 -22100
rect -5299 -22134 -5293 -22100
rect -5339 -22172 -5293 -22134
rect -5339 -22206 -5333 -22172
rect -5299 -22206 -5293 -22172
rect -5339 -22244 -5293 -22206
rect -5339 -22278 -5333 -22244
rect -5299 -22278 -5293 -22244
rect -5339 -22316 -5293 -22278
rect -6317 -22350 -6304 -22328
rect -5339 -22330 -5333 -22316
rect -7087 -22419 -6599 -22413
rect -7087 -22453 -7040 -22419
rect -7006 -22453 -6968 -22419
rect -6934 -22453 -6896 -22419
rect -6862 -22453 -6824 -22419
rect -6790 -22453 -6752 -22419
rect -6718 -22453 -6680 -22419
rect -6646 -22453 -6599 -22419
rect -7087 -22459 -6599 -22453
rect -7392 -22604 -7320 -22600
rect -7392 -22656 -7382 -22604
rect -7330 -22656 -7320 -22604
rect -7392 -22660 -7320 -22656
rect -8106 -22822 -7618 -22816
rect -8106 -22856 -8059 -22822
rect -8025 -22856 -7987 -22822
rect -7953 -22856 -7915 -22822
rect -7881 -22856 -7843 -22822
rect -7809 -22856 -7771 -22822
rect -7737 -22856 -7699 -22822
rect -7665 -22856 -7618 -22822
rect -8106 -22862 -7618 -22856
rect -8402 -22952 -8388 -22925
rect -9418 -22966 -9358 -22959
rect -8394 -22959 -8388 -22952
rect -8354 -22952 -8342 -22925
rect -7386 -22925 -7326 -22660
rect -6870 -22816 -6810 -22459
rect -6364 -22716 -6304 -22350
rect -5346 -22350 -5333 -22330
rect -5299 -22330 -5293 -22316
rect -4321 -21884 -4275 -21846
rect -4321 -21918 -4315 -21884
rect -4281 -21918 -4275 -21884
rect -4321 -21956 -4275 -21918
rect -4321 -21990 -4315 -21956
rect -4281 -21990 -4275 -21956
rect -4321 -22028 -4275 -21990
rect -4321 -22062 -4315 -22028
rect -4281 -22062 -4275 -22028
rect -4321 -22100 -4275 -22062
rect -4321 -22134 -4315 -22100
rect -4281 -22134 -4275 -22100
rect -4321 -22172 -4275 -22134
rect -4321 -22206 -4315 -22172
rect -4281 -22206 -4275 -22172
rect -4321 -22244 -4275 -22206
rect -4321 -22278 -4315 -22244
rect -4281 -22278 -4275 -22244
rect -4321 -22316 -4275 -22278
rect -4321 -22324 -4315 -22316
rect -5299 -22350 -5286 -22330
rect -6069 -22419 -5581 -22413
rect -6069 -22453 -6022 -22419
rect -5988 -22453 -5950 -22419
rect -5916 -22453 -5878 -22419
rect -5844 -22453 -5806 -22419
rect -5772 -22453 -5734 -22419
rect -5700 -22453 -5662 -22419
rect -5628 -22453 -5581 -22419
rect -6069 -22459 -5581 -22453
rect -6370 -22720 -6298 -22716
rect -6370 -22772 -6360 -22720
rect -6308 -22772 -6298 -22720
rect -6370 -22776 -6298 -22772
rect -5862 -22816 -5802 -22459
rect -5346 -22600 -5286 -22350
rect -4326 -22350 -4315 -22324
rect -4281 -22324 -4275 -22316
rect -3303 -21884 -3257 -21846
rect -3303 -21918 -3297 -21884
rect -3263 -21918 -3257 -21884
rect -3303 -21956 -3257 -21918
rect -3303 -21990 -3297 -21956
rect -3263 -21990 -3257 -21956
rect -3303 -22028 -3257 -21990
rect -3303 -22062 -3297 -22028
rect -3263 -22062 -3257 -22028
rect -3303 -22100 -3257 -22062
rect -3303 -22134 -3297 -22100
rect -3263 -22134 -3257 -22100
rect -3303 -22172 -3257 -22134
rect -3303 -22206 -3297 -22172
rect -3263 -22206 -3257 -22172
rect -3303 -22244 -3257 -22206
rect -3303 -22278 -3297 -22244
rect -3263 -22278 -3257 -22244
rect -3303 -22316 -3257 -22278
rect -4281 -22350 -4266 -22324
rect -5051 -22419 -4563 -22413
rect -5051 -22453 -5004 -22419
rect -4970 -22453 -4932 -22419
rect -4898 -22453 -4860 -22419
rect -4826 -22453 -4788 -22419
rect -4754 -22453 -4716 -22419
rect -4682 -22453 -4644 -22419
rect -4610 -22453 -4563 -22419
rect -5051 -22459 -4563 -22453
rect -5352 -22604 -5280 -22600
rect -5352 -22656 -5342 -22604
rect -5290 -22656 -5280 -22604
rect -5352 -22660 -5280 -22656
rect -7088 -22822 -6600 -22816
rect -7088 -22856 -7041 -22822
rect -7007 -22856 -6969 -22822
rect -6935 -22856 -6897 -22822
rect -6863 -22856 -6825 -22822
rect -6791 -22856 -6753 -22822
rect -6719 -22856 -6681 -22822
rect -6647 -22856 -6600 -22822
rect -7088 -22862 -6600 -22856
rect -6070 -22822 -5582 -22816
rect -6070 -22856 -6023 -22822
rect -5989 -22856 -5951 -22822
rect -5917 -22856 -5879 -22822
rect -5845 -22856 -5807 -22822
rect -5773 -22856 -5735 -22822
rect -5701 -22856 -5663 -22822
rect -5629 -22856 -5582 -22822
rect -6070 -22862 -5582 -22856
rect -7386 -22952 -7370 -22925
rect -8354 -22959 -8348 -22952
rect -9412 -22997 -9366 -22966
rect -9412 -23031 -9406 -22997
rect -9372 -23031 -9366 -22997
rect -9412 -23069 -9366 -23031
rect -9412 -23103 -9406 -23069
rect -9372 -23103 -9366 -23069
rect -9412 -23141 -9366 -23103
rect -9412 -23175 -9406 -23141
rect -9372 -23175 -9366 -23141
rect -9412 -23213 -9366 -23175
rect -9412 -23247 -9406 -23213
rect -9372 -23247 -9366 -23213
rect -9412 -23285 -9366 -23247
rect -9412 -23319 -9406 -23285
rect -9372 -23319 -9366 -23285
rect -9412 -23357 -9366 -23319
rect -9412 -23391 -9406 -23357
rect -9372 -23391 -9366 -23357
rect -9412 -23429 -9366 -23391
rect -9412 -23463 -9406 -23429
rect -9372 -23463 -9366 -23429
rect -8394 -22997 -8348 -22959
rect -8394 -23031 -8388 -22997
rect -8354 -23031 -8348 -22997
rect -8394 -23069 -8348 -23031
rect -8394 -23103 -8388 -23069
rect -8354 -23103 -8348 -23069
rect -8394 -23141 -8348 -23103
rect -8394 -23175 -8388 -23141
rect -8354 -23175 -8348 -23141
rect -8394 -23213 -8348 -23175
rect -8394 -23247 -8388 -23213
rect -8354 -23247 -8348 -23213
rect -8394 -23285 -8348 -23247
rect -8394 -23319 -8388 -23285
rect -8354 -23319 -8348 -23285
rect -8394 -23357 -8348 -23319
rect -8394 -23391 -8388 -23357
rect -8354 -23391 -8348 -23357
rect -8394 -23429 -8348 -23391
rect -8394 -23436 -8388 -23429
rect -9412 -23494 -9366 -23463
rect -8402 -23463 -8388 -23436
rect -8354 -23436 -8348 -23429
rect -7376 -22959 -7370 -22952
rect -7336 -22952 -7326 -22925
rect -6358 -22925 -6312 -22894
rect -7336 -22959 -7330 -22952
rect -7376 -22997 -7330 -22959
rect -7376 -23031 -7370 -22997
rect -7336 -23031 -7330 -22997
rect -7376 -23069 -7330 -23031
rect -7376 -23103 -7370 -23069
rect -7336 -23103 -7330 -23069
rect -7376 -23141 -7330 -23103
rect -7376 -23175 -7370 -23141
rect -7336 -23175 -7330 -23141
rect -7376 -23213 -7330 -23175
rect -7376 -23247 -7370 -23213
rect -7336 -23247 -7330 -23213
rect -7376 -23285 -7330 -23247
rect -7376 -23319 -7370 -23285
rect -7336 -23319 -7330 -23285
rect -7376 -23357 -7330 -23319
rect -7376 -23391 -7370 -23357
rect -7336 -23391 -7330 -23357
rect -7376 -23429 -7330 -23391
rect -8354 -23463 -8342 -23436
rect -7376 -23440 -7370 -23429
rect -9124 -23532 -8636 -23526
rect -9124 -23566 -9077 -23532
rect -9043 -23566 -9005 -23532
rect -8971 -23566 -8933 -23532
rect -8899 -23566 -8861 -23532
rect -8827 -23566 -8789 -23532
rect -8755 -23566 -8717 -23532
rect -8683 -23566 -8636 -23532
rect -9124 -23572 -8636 -23566
rect -8402 -23724 -8342 -23463
rect -7384 -23463 -7370 -23440
rect -7336 -23440 -7330 -23429
rect -6358 -22959 -6352 -22925
rect -6318 -22959 -6312 -22925
rect -5346 -22925 -5286 -22660
rect -4840 -22816 -4780 -22459
rect -4326 -22504 -4266 -22350
rect -3303 -22350 -3297 -22316
rect -3263 -22350 -3257 -22316
rect -3303 -22381 -3257 -22350
rect -4033 -22419 -3545 -22413
rect -4033 -22453 -3986 -22419
rect -3952 -22453 -3914 -22419
rect -3880 -22453 -3842 -22419
rect -3808 -22453 -3770 -22419
rect -3736 -22453 -3698 -22419
rect -3664 -22453 -3626 -22419
rect -3592 -22453 -3545 -22419
rect -4033 -22459 -3545 -22453
rect -4332 -22508 -4260 -22504
rect -4332 -22560 -4322 -22508
rect -4270 -22560 -4260 -22508
rect -4332 -22564 -4260 -22560
rect -2846 -22610 -2786 -19060
rect -820 -19128 -748 -19124
rect -820 -19180 -810 -19128
rect -758 -19180 -748 -19128
rect -820 -19184 -748 -19180
rect 92 -19128 164 -19124
rect 92 -19180 102 -19128
rect 154 -19180 164 -19128
rect 92 -19184 164 -19180
rect -1690 -19238 -1618 -19234
rect -1690 -19290 -1680 -19238
rect -1628 -19290 -1618 -19238
rect -1690 -19294 -1618 -19290
rect -2604 -19346 -2532 -19342
rect -2604 -19398 -2594 -19346
rect -2542 -19398 -2532 -19346
rect -2604 -19402 -2532 -19398
rect -2598 -20896 -2538 -19402
rect -2474 -19454 -2402 -19450
rect -2474 -19506 -2464 -19454
rect -2412 -19506 -2402 -19454
rect -2474 -19510 -2402 -19506
rect -2468 -20774 -2408 -19510
rect -2242 -19550 -2154 -19544
rect -2242 -19584 -2215 -19550
rect -2181 -19584 -2154 -19550
rect -2242 -19590 -2154 -19584
rect -2024 -19550 -1936 -19544
rect -2024 -19584 -1997 -19550
rect -1963 -19584 -1936 -19550
rect -2024 -19590 -1936 -19584
rect -1806 -19550 -1718 -19544
rect -1806 -19584 -1779 -19550
rect -1745 -19584 -1718 -19550
rect -1806 -19590 -1718 -19584
rect -2330 -19669 -2284 -19622
rect -2330 -19703 -2324 -19669
rect -2290 -19703 -2284 -19669
rect -2330 -19741 -2284 -19703
rect -2330 -19775 -2324 -19741
rect -2290 -19775 -2284 -19741
rect -2330 -19780 -2284 -19775
rect -2112 -19669 -2066 -19622
rect -2112 -19703 -2106 -19669
rect -2072 -19703 -2066 -19669
rect -2112 -19741 -2066 -19703
rect -2112 -19775 -2106 -19741
rect -2072 -19775 -2066 -19741
rect -2338 -19960 -2278 -19780
rect -2112 -19788 -2066 -19775
rect -1894 -19669 -1848 -19622
rect -1684 -19650 -1624 -19294
rect -926 -19346 -854 -19342
rect -926 -19398 -916 -19346
rect -864 -19398 -854 -19346
rect -926 -19402 -854 -19398
rect -1144 -19454 -1072 -19450
rect -1144 -19506 -1134 -19454
rect -1082 -19506 -1072 -19454
rect -1144 -19510 -1072 -19506
rect -1138 -19544 -1078 -19510
rect -920 -19544 -860 -19402
rect -1588 -19550 -1500 -19544
rect -1588 -19584 -1561 -19550
rect -1527 -19584 -1500 -19550
rect -1588 -19590 -1500 -19584
rect -1370 -19550 -1282 -19544
rect -1370 -19584 -1343 -19550
rect -1309 -19584 -1282 -19550
rect -1370 -19590 -1282 -19584
rect -1152 -19550 -1064 -19544
rect -1152 -19584 -1125 -19550
rect -1091 -19584 -1064 -19550
rect -1152 -19590 -1064 -19584
rect -934 -19550 -846 -19544
rect -934 -19584 -907 -19550
rect -873 -19584 -846 -19550
rect -934 -19590 -846 -19584
rect -1894 -19703 -1888 -19669
rect -1854 -19703 -1848 -19669
rect -1894 -19741 -1848 -19703
rect -1894 -19775 -1888 -19741
rect -1854 -19775 -1848 -19741
rect -2242 -19860 -2154 -19854
rect -2242 -19894 -2215 -19860
rect -2181 -19894 -2154 -19860
rect -2242 -19900 -2154 -19894
rect -2230 -19960 -2170 -19900
rect -2118 -19960 -2058 -19788
rect -1894 -19798 -1848 -19775
rect -1676 -19669 -1630 -19650
rect -1676 -19703 -1670 -19669
rect -1636 -19703 -1630 -19669
rect -1676 -19741 -1630 -19703
rect -1676 -19775 -1670 -19741
rect -1636 -19775 -1630 -19741
rect -2024 -19860 -1936 -19854
rect -2024 -19894 -1997 -19860
rect -1963 -19894 -1936 -19860
rect -2024 -19900 -1936 -19894
rect -2010 -19950 -1950 -19900
rect -2338 -20020 -2058 -19960
rect -2016 -19954 -1944 -19950
rect -2016 -20006 -2006 -19954
rect -1954 -20006 -1944 -19954
rect -2016 -20010 -1944 -20006
rect -2118 -20278 -2058 -20020
rect -1902 -20050 -1842 -19798
rect -1676 -19822 -1630 -19775
rect -1458 -19669 -1412 -19622
rect -1458 -19703 -1452 -19669
rect -1418 -19703 -1412 -19669
rect -1458 -19741 -1412 -19703
rect -1458 -19775 -1452 -19741
rect -1418 -19775 -1412 -19741
rect -1240 -19669 -1194 -19622
rect -1240 -19703 -1234 -19669
rect -1200 -19703 -1194 -19669
rect -1240 -19741 -1194 -19703
rect -1240 -19774 -1234 -19741
rect -1458 -19784 -1412 -19775
rect -1248 -19775 -1234 -19774
rect -1200 -19774 -1194 -19741
rect -1022 -19669 -976 -19622
rect -1022 -19703 -1016 -19669
rect -982 -19703 -976 -19669
rect -814 -19669 -754 -19184
rect -28 -19238 44 -19234
rect -28 -19290 -18 -19238
rect 34 -19290 44 -19238
rect -28 -19294 44 -19290
rect -708 -19346 -636 -19342
rect -708 -19398 -698 -19346
rect -646 -19398 -636 -19346
rect -708 -19402 -636 -19398
rect -702 -19544 -642 -19402
rect -490 -19454 -418 -19450
rect -490 -19506 -480 -19454
rect -428 -19506 -418 -19454
rect -490 -19510 -418 -19506
rect -484 -19544 -424 -19510
rect -716 -19550 -628 -19544
rect -716 -19584 -689 -19550
rect -655 -19584 -628 -19550
rect -716 -19590 -628 -19584
rect -498 -19550 -410 -19544
rect -498 -19584 -471 -19550
rect -437 -19584 -410 -19550
rect -498 -19590 -410 -19584
rect -280 -19550 -192 -19544
rect -280 -19584 -253 -19550
rect -219 -19584 -192 -19550
rect -280 -19590 -192 -19584
rect -814 -19680 -798 -19669
rect -1022 -19741 -976 -19703
rect -1200 -19775 -1188 -19774
rect -1806 -19860 -1718 -19854
rect -1806 -19894 -1779 -19860
rect -1745 -19894 -1718 -19860
rect -1806 -19900 -1718 -19894
rect -1588 -19860 -1500 -19854
rect -1588 -19894 -1561 -19860
rect -1527 -19894 -1500 -19860
rect -1588 -19900 -1500 -19894
rect -1908 -20054 -1836 -20050
rect -1908 -20106 -1898 -20054
rect -1846 -20106 -1836 -20054
rect -1908 -20110 -1836 -20106
rect -1906 -20164 -1834 -20160
rect -1906 -20216 -1896 -20164
rect -1844 -20216 -1834 -20164
rect -1906 -20220 -1834 -20216
rect -2336 -20338 -2058 -20278
rect -2336 -20492 -2276 -20338
rect -2226 -20376 -2166 -20338
rect -2242 -20382 -2154 -20376
rect -2242 -20416 -2215 -20382
rect -2181 -20416 -2154 -20382
rect -2242 -20422 -2154 -20416
rect -2330 -20501 -2284 -20492
rect -2330 -20535 -2324 -20501
rect -2290 -20535 -2284 -20501
rect -2330 -20573 -2284 -20535
rect -2330 -20607 -2324 -20573
rect -2290 -20607 -2284 -20573
rect -2330 -20654 -2284 -20607
rect -2118 -20501 -2058 -20338
rect -2024 -20382 -1936 -20376
rect -2024 -20416 -1997 -20382
rect -1963 -20416 -1936 -20382
rect -2024 -20422 -1936 -20416
rect -2118 -20535 -2106 -20501
rect -2072 -20535 -2058 -20501
rect -1900 -20501 -1840 -20220
rect -1792 -20270 -1732 -19900
rect -1572 -20270 -1512 -19900
rect -1464 -20050 -1404 -19784
rect -1370 -19860 -1282 -19854
rect -1370 -19894 -1343 -19860
rect -1309 -19894 -1282 -19860
rect -1370 -19900 -1282 -19894
rect -1354 -19950 -1294 -19900
rect -1360 -19954 -1288 -19950
rect -1360 -20006 -1350 -19954
rect -1298 -20006 -1288 -19954
rect -1360 -20010 -1288 -20006
rect -1470 -20054 -1398 -20050
rect -1470 -20106 -1460 -20054
rect -1408 -20106 -1398 -20054
rect -1470 -20110 -1398 -20106
rect -1472 -20164 -1400 -20160
rect -1472 -20216 -1462 -20164
rect -1410 -20216 -1400 -20164
rect -1472 -20220 -1400 -20216
rect -1798 -20274 -1726 -20270
rect -1798 -20326 -1788 -20274
rect -1736 -20326 -1726 -20274
rect -1798 -20330 -1726 -20326
rect -1578 -20274 -1506 -20270
rect -1578 -20326 -1568 -20274
rect -1516 -20326 -1506 -20274
rect -1578 -20330 -1506 -20326
rect -1792 -20376 -1732 -20330
rect -1572 -20376 -1512 -20330
rect -1806 -20382 -1718 -20376
rect -1806 -20416 -1779 -20382
rect -1745 -20416 -1718 -20382
rect -1806 -20422 -1718 -20416
rect -1588 -20382 -1500 -20376
rect -1588 -20416 -1561 -20382
rect -1527 -20416 -1500 -20382
rect -1588 -20422 -1500 -20416
rect -1900 -20502 -1888 -20501
rect -2118 -20573 -2058 -20535
rect -2118 -20607 -2106 -20573
rect -2072 -20607 -2058 -20573
rect -2242 -20692 -2154 -20686
rect -2242 -20726 -2215 -20692
rect -2181 -20726 -2154 -20692
rect -2242 -20732 -2154 -20726
rect -2474 -20778 -2402 -20774
rect -2474 -20830 -2464 -20778
rect -2412 -20830 -2402 -20778
rect -2474 -20834 -2402 -20830
rect -2604 -20900 -2532 -20896
rect -2604 -20952 -2594 -20900
rect -2542 -20952 -2532 -20900
rect -2604 -20956 -2532 -20952
rect -2118 -21020 -2058 -20607
rect -1894 -20535 -1888 -20502
rect -1854 -20502 -1840 -20501
rect -1676 -20501 -1630 -20454
rect -1466 -20496 -1406 -20220
rect -1370 -20382 -1282 -20376
rect -1370 -20416 -1343 -20382
rect -1309 -20416 -1282 -20382
rect -1370 -20422 -1282 -20416
rect -1854 -20535 -1848 -20502
rect -1894 -20573 -1848 -20535
rect -1894 -20607 -1888 -20573
rect -1854 -20607 -1848 -20573
rect -1676 -20535 -1670 -20501
rect -1636 -20535 -1630 -20501
rect -1676 -20573 -1630 -20535
rect -1676 -20602 -1670 -20573
rect -1894 -20654 -1848 -20607
rect -1680 -20607 -1670 -20602
rect -1636 -20602 -1630 -20573
rect -1458 -20501 -1412 -20496
rect -1458 -20535 -1452 -20501
rect -1418 -20535 -1412 -20501
rect -1458 -20573 -1412 -20535
rect -1636 -20607 -1620 -20602
rect -2024 -20692 -1936 -20686
rect -2024 -20726 -1997 -20692
rect -1963 -20726 -1936 -20692
rect -2024 -20732 -1936 -20726
rect -1806 -20692 -1718 -20686
rect -1806 -20726 -1779 -20692
rect -1745 -20726 -1718 -20692
rect -1806 -20732 -1718 -20726
rect -2010 -20774 -1950 -20732
rect -2016 -20778 -1944 -20774
rect -2016 -20830 -2006 -20778
rect -1954 -20830 -1944 -20778
rect -2016 -20834 -1944 -20830
rect -1792 -20896 -1732 -20732
rect -1798 -20900 -1726 -20896
rect -1798 -20952 -1788 -20900
rect -1736 -20952 -1726 -20900
rect -1798 -20956 -1726 -20952
rect -2124 -21024 -2052 -21020
rect -2124 -21076 -2114 -21024
rect -2062 -21076 -2052 -21024
rect -2124 -21080 -2052 -21076
rect -1680 -21146 -1620 -20607
rect -1458 -20607 -1452 -20573
rect -1418 -20607 -1412 -20573
rect -1458 -20654 -1412 -20607
rect -1248 -20501 -1188 -19775
rect -1022 -19775 -1016 -19741
rect -982 -19775 -976 -19741
rect -1022 -19776 -976 -19775
rect -804 -19703 -798 -19680
rect -764 -19680 -754 -19669
rect -586 -19669 -540 -19622
rect -764 -19703 -758 -19680
rect -804 -19741 -758 -19703
rect -804 -19775 -798 -19741
rect -764 -19775 -758 -19741
rect -1152 -19860 -1064 -19854
rect -1152 -19894 -1125 -19860
rect -1091 -19894 -1064 -19860
rect -1152 -19900 -1064 -19894
rect -1028 -20050 -968 -19776
rect -804 -19822 -758 -19775
rect -586 -19703 -580 -19669
rect -546 -19703 -540 -19669
rect -586 -19741 -540 -19703
rect -586 -19775 -580 -19741
rect -546 -19775 -540 -19741
rect -586 -19784 -540 -19775
rect -368 -19669 -322 -19622
rect -368 -19703 -362 -19669
rect -328 -19703 -322 -19669
rect -368 -19741 -322 -19703
rect -368 -19775 -362 -19741
rect -328 -19775 -322 -19741
rect -150 -19669 -104 -19622
rect -150 -19703 -144 -19669
rect -110 -19703 -104 -19669
rect -150 -19741 -104 -19703
rect -150 -19774 -144 -19741
rect -934 -19860 -846 -19854
rect -934 -19894 -907 -19860
rect -873 -19894 -846 -19860
rect -934 -19900 -846 -19894
rect -716 -19860 -628 -19854
rect -716 -19894 -689 -19860
rect -655 -19894 -628 -19860
rect -716 -19900 -628 -19894
rect -592 -20050 -532 -19784
rect -368 -19792 -322 -19775
rect -156 -19775 -144 -19774
rect -110 -19774 -104 -19741
rect -22 -19728 38 -19294
rect -110 -19775 -96 -19774
rect -498 -19860 -410 -19854
rect -498 -19894 -471 -19860
rect -437 -19894 -410 -19860
rect -498 -19900 -410 -19894
rect -490 -19954 -418 -19950
rect -490 -20006 -480 -19954
rect -428 -20006 -418 -19954
rect -490 -20010 -418 -20006
rect -374 -19952 -314 -19792
rect -280 -19860 -192 -19854
rect -280 -19894 -253 -19860
rect -219 -19894 -192 -19860
rect -280 -19900 -192 -19894
rect -266 -19952 -206 -19900
rect -156 -19952 -96 -19775
rect -1138 -20110 -532 -20050
rect -1138 -20160 -1078 -20110
rect -1144 -20164 -1072 -20160
rect -1144 -20216 -1134 -20164
rect -1082 -20216 -1072 -20164
rect -1144 -20220 -1072 -20216
rect -1034 -20164 -962 -20160
rect -1034 -20216 -1024 -20164
rect -972 -20216 -962 -20164
rect -1034 -20220 -962 -20216
rect -598 -20164 -526 -20160
rect -598 -20216 -588 -20164
rect -536 -20216 -526 -20164
rect -598 -20220 -526 -20216
rect -1152 -20382 -1064 -20376
rect -1152 -20416 -1125 -20382
rect -1091 -20416 -1064 -20382
rect -1152 -20422 -1064 -20416
rect -1028 -20484 -968 -20220
rect -924 -20274 -852 -20270
rect -924 -20326 -914 -20274
rect -862 -20326 -852 -20274
rect -924 -20330 -852 -20326
rect -708 -20274 -636 -20270
rect -708 -20326 -698 -20274
rect -646 -20326 -636 -20274
rect -708 -20330 -636 -20326
rect -918 -20376 -858 -20330
rect -702 -20376 -642 -20330
rect -934 -20382 -846 -20376
rect -934 -20416 -907 -20382
rect -873 -20416 -846 -20382
rect -934 -20422 -846 -20416
rect -716 -20382 -628 -20376
rect -716 -20416 -689 -20382
rect -655 -20416 -628 -20382
rect -716 -20422 -628 -20416
rect -1248 -20535 -1234 -20501
rect -1200 -20535 -1188 -20501
rect -1248 -20573 -1188 -20535
rect -1248 -20607 -1234 -20573
rect -1200 -20607 -1188 -20573
rect -1588 -20692 -1500 -20686
rect -1588 -20726 -1561 -20692
rect -1527 -20726 -1500 -20692
rect -1588 -20732 -1500 -20726
rect -1370 -20692 -1282 -20686
rect -1370 -20726 -1343 -20692
rect -1309 -20726 -1282 -20692
rect -1370 -20732 -1282 -20726
rect -1574 -20896 -1514 -20732
rect -1354 -20774 -1294 -20732
rect -1360 -20778 -1288 -20774
rect -1360 -20830 -1350 -20778
rect -1298 -20830 -1288 -20778
rect -1360 -20834 -1288 -20830
rect -1580 -20900 -1508 -20896
rect -1580 -20952 -1570 -20900
rect -1518 -20952 -1508 -20900
rect -1580 -20956 -1508 -20952
rect -1686 -21150 -1614 -21146
rect -1686 -21202 -1676 -21150
rect -1624 -21202 -1614 -21150
rect -1686 -21206 -1614 -21202
rect -1344 -21260 -1296 -20834
rect -1248 -21020 -1188 -20607
rect -1022 -20501 -976 -20484
rect -1022 -20535 -1016 -20501
rect -982 -20535 -976 -20501
rect -1022 -20573 -976 -20535
rect -1022 -20607 -1016 -20573
rect -982 -20607 -976 -20573
rect -1022 -20654 -976 -20607
rect -804 -20501 -758 -20454
rect -592 -20498 -532 -20220
rect -484 -20376 -424 -20010
rect -374 -20012 -96 -19952
rect -22 -19780 -18 -19728
rect 34 -19780 38 -19728
rect -374 -20070 -314 -20012
rect -380 -20074 -308 -20070
rect -380 -20126 -370 -20074
rect -318 -20126 -308 -20074
rect -380 -20130 -308 -20126
rect -374 -20268 -314 -20130
rect -374 -20328 -96 -20268
rect -498 -20382 -410 -20376
rect -498 -20416 -471 -20382
rect -437 -20416 -410 -20382
rect -498 -20422 -410 -20416
rect -374 -20484 -314 -20328
rect -266 -20376 -206 -20328
rect -280 -20382 -192 -20376
rect -280 -20416 -253 -20382
rect -219 -20416 -192 -20382
rect -280 -20422 -192 -20416
rect -804 -20535 -798 -20501
rect -764 -20535 -758 -20501
rect -804 -20573 -758 -20535
rect -804 -20607 -798 -20573
rect -764 -20607 -758 -20573
rect -804 -20620 -758 -20607
rect -586 -20501 -540 -20498
rect -586 -20535 -580 -20501
rect -546 -20535 -540 -20501
rect -586 -20573 -540 -20535
rect -586 -20607 -580 -20573
rect -546 -20607 -540 -20573
rect -1152 -20692 -1064 -20686
rect -1152 -20726 -1125 -20692
rect -1091 -20726 -1064 -20692
rect -1152 -20732 -1064 -20726
rect -934 -20692 -846 -20686
rect -934 -20726 -907 -20692
rect -873 -20726 -846 -20692
rect -934 -20732 -846 -20726
rect -1138 -20894 -1078 -20732
rect -810 -20774 -750 -20620
rect -586 -20654 -540 -20607
rect -368 -20501 -322 -20484
rect -156 -20486 -96 -20328
rect -368 -20535 -362 -20501
rect -328 -20535 -322 -20501
rect -368 -20573 -322 -20535
rect -368 -20607 -362 -20573
rect -328 -20607 -322 -20573
rect -368 -20612 -322 -20607
rect -150 -20501 -104 -20486
rect -150 -20535 -144 -20501
rect -110 -20535 -104 -20501
rect -150 -20573 -104 -20535
rect -150 -20607 -144 -20573
rect -110 -20607 -104 -20573
rect -716 -20692 -628 -20686
rect -716 -20726 -689 -20692
rect -655 -20726 -628 -20692
rect -716 -20732 -628 -20726
rect -498 -20692 -410 -20686
rect -498 -20726 -471 -20692
rect -437 -20726 -410 -20692
rect -498 -20732 -410 -20726
rect -816 -20778 -744 -20774
rect -816 -20830 -806 -20778
rect -754 -20830 -744 -20778
rect -816 -20834 -744 -20830
rect -482 -20894 -422 -20732
rect -1144 -20898 -1072 -20894
rect -1144 -20950 -1134 -20898
rect -1082 -20950 -1072 -20898
rect -1144 -20954 -1072 -20950
rect -488 -20898 -416 -20894
rect -488 -20950 -478 -20898
rect -426 -20950 -416 -20898
rect -488 -20954 -416 -20950
rect -376 -21020 -316 -20612
rect -150 -20654 -104 -20607
rect -280 -20692 -192 -20686
rect -280 -20726 -253 -20692
rect -219 -20726 -192 -20692
rect -280 -20732 -192 -20726
rect -22 -20774 38 -19780
rect -28 -20778 44 -20774
rect -28 -20830 -18 -20778
rect 34 -20830 44 -20778
rect -28 -20834 44 -20830
rect -1254 -21024 -1182 -21020
rect -1254 -21076 -1244 -21024
rect -1192 -21076 -1182 -21024
rect -1254 -21080 -1182 -21076
rect -382 -21024 -310 -21020
rect -382 -21076 -372 -21024
rect -320 -21076 -310 -21024
rect -382 -21080 -310 -21076
rect 98 -21146 158 -19184
rect 214 -19954 286 -19950
rect 214 -20006 224 -19954
rect 276 -20006 286 -19954
rect 214 -20010 286 -20006
rect 220 -20200 280 -20010
rect 220 -20252 224 -20200
rect 276 -20252 280 -20200
rect 220 -20264 280 -20252
rect 92 -21150 164 -21146
rect 92 -21202 102 -21150
rect 154 -21202 164 -21150
rect 92 -21206 164 -21202
rect -1352 -21312 -1346 -21260
rect -1294 -21312 -1288 -21260
rect 690 -21340 750 -18944
rect -2538 -21400 750 -21340
rect 952 -18914 956 -18862
rect 1008 -18914 1012 -18862
rect -2676 -21584 -2604 -21580
rect -2676 -21636 -2666 -21584
rect -2614 -21636 -2604 -21584
rect -2676 -21640 -2604 -21636
rect -4328 -22670 -2786 -22610
rect -5052 -22822 -4564 -22816
rect -5052 -22856 -5005 -22822
rect -4971 -22856 -4933 -22822
rect -4899 -22856 -4861 -22822
rect -4827 -22856 -4789 -22822
rect -4755 -22856 -4717 -22822
rect -4683 -22856 -4645 -22822
rect -4611 -22856 -4564 -22822
rect -5052 -22862 -4564 -22856
rect -5346 -22940 -5334 -22925
rect -6358 -22997 -6312 -22959
rect -6358 -23031 -6352 -22997
rect -6318 -23031 -6312 -22997
rect -6358 -23069 -6312 -23031
rect -6358 -23103 -6352 -23069
rect -6318 -23103 -6312 -23069
rect -6358 -23141 -6312 -23103
rect -6358 -23175 -6352 -23141
rect -6318 -23175 -6312 -23141
rect -6358 -23213 -6312 -23175
rect -6358 -23247 -6352 -23213
rect -6318 -23247 -6312 -23213
rect -6358 -23285 -6312 -23247
rect -6358 -23319 -6352 -23285
rect -6318 -23319 -6312 -23285
rect -6358 -23357 -6312 -23319
rect -6358 -23391 -6352 -23357
rect -6318 -23391 -6312 -23357
rect -6358 -23429 -6312 -23391
rect -6358 -23430 -6352 -23429
rect -7336 -23463 -7324 -23440
rect -8106 -23532 -7618 -23526
rect -8106 -23566 -8059 -23532
rect -8025 -23566 -7987 -23532
rect -7953 -23566 -7915 -23532
rect -7881 -23566 -7843 -23532
rect -7809 -23566 -7771 -23532
rect -7737 -23566 -7699 -23532
rect -7665 -23566 -7618 -23532
rect -8106 -23572 -7618 -23566
rect -8260 -23620 -8188 -23616
rect -8260 -23672 -8250 -23620
rect -8198 -23672 -8188 -23620
rect -8260 -23676 -8188 -23672
rect -8408 -23728 -8336 -23724
rect -8408 -23780 -8398 -23728
rect -8346 -23780 -8336 -23728
rect -8408 -23784 -8336 -23780
rect -8254 -23826 -8194 -23676
rect -9418 -23886 -8194 -23826
rect -9418 -24036 -9358 -23886
rect -8902 -23927 -8842 -23886
rect -9123 -23933 -8635 -23927
rect -9123 -23967 -9076 -23933
rect -9042 -23967 -9004 -23933
rect -8970 -23967 -8932 -23933
rect -8898 -23967 -8860 -23933
rect -8826 -23967 -8788 -23933
rect -8754 -23967 -8716 -23933
rect -8682 -23967 -8635 -23933
rect -9123 -23973 -8635 -23967
rect -9418 -24058 -9405 -24036
rect -9411 -24070 -9405 -24058
rect -9371 -24058 -9358 -24036
rect -8400 -24036 -8340 -23886
rect -7884 -23927 -7824 -23572
rect -7384 -23836 -7324 -23463
rect -6368 -23463 -6352 -23430
rect -6318 -23430 -6312 -23429
rect -5340 -22959 -5334 -22940
rect -5300 -22940 -5286 -22925
rect -4328 -22906 -4268 -22670
rect -3818 -22816 -3758 -22670
rect -4034 -22822 -3546 -22816
rect -4034 -22856 -3987 -22822
rect -3953 -22856 -3915 -22822
rect -3881 -22856 -3843 -22822
rect -3809 -22856 -3771 -22822
rect -3737 -22856 -3699 -22822
rect -3665 -22856 -3627 -22822
rect -3593 -22856 -3546 -22822
rect -4034 -22862 -3546 -22856
rect -3312 -22906 -3252 -22670
rect -3208 -22720 -3136 -22716
rect -3208 -22772 -3198 -22720
rect -3146 -22772 -3136 -22720
rect -3208 -22776 -3136 -22772
rect -4328 -22925 -4266 -22906
rect -5300 -22959 -5294 -22940
rect -4328 -22952 -4316 -22925
rect -4326 -22954 -4316 -22952
rect -5340 -22997 -5294 -22959
rect -5340 -23031 -5334 -22997
rect -5300 -23031 -5294 -22997
rect -5340 -23069 -5294 -23031
rect -5340 -23103 -5334 -23069
rect -5300 -23103 -5294 -23069
rect -5340 -23141 -5294 -23103
rect -5340 -23175 -5334 -23141
rect -5300 -23175 -5294 -23141
rect -5340 -23213 -5294 -23175
rect -5340 -23247 -5334 -23213
rect -5300 -23247 -5294 -23213
rect -5340 -23285 -5294 -23247
rect -5340 -23319 -5334 -23285
rect -5300 -23319 -5294 -23285
rect -5340 -23357 -5294 -23319
rect -5340 -23391 -5334 -23357
rect -5300 -23391 -5294 -23357
rect -5340 -23429 -5294 -23391
rect -6318 -23463 -6308 -23430
rect -5340 -23448 -5334 -23429
rect -7088 -23532 -6600 -23526
rect -7088 -23566 -7041 -23532
rect -7007 -23566 -6969 -23532
rect -6935 -23566 -6897 -23532
rect -6863 -23566 -6825 -23532
rect -6791 -23566 -6753 -23532
rect -6719 -23566 -6681 -23532
rect -6647 -23566 -6600 -23532
rect -7088 -23572 -6600 -23566
rect -7390 -23840 -7318 -23836
rect -7390 -23892 -7380 -23840
rect -7328 -23892 -7318 -23840
rect -7390 -23896 -7318 -23892
rect -8105 -23933 -7617 -23927
rect -8105 -23967 -8058 -23933
rect -8024 -23967 -7986 -23933
rect -7952 -23967 -7914 -23933
rect -7880 -23967 -7842 -23933
rect -7808 -23967 -7770 -23933
rect -7736 -23967 -7698 -23933
rect -7664 -23967 -7617 -23933
rect -8105 -23973 -7617 -23967
rect -8400 -24058 -8387 -24036
rect -9371 -24070 -9365 -24058
rect -9411 -24108 -9365 -24070
rect -9411 -24142 -9405 -24108
rect -9371 -24142 -9365 -24108
rect -9411 -24180 -9365 -24142
rect -9411 -24214 -9405 -24180
rect -9371 -24214 -9365 -24180
rect -9411 -24252 -9365 -24214
rect -9411 -24286 -9405 -24252
rect -9371 -24286 -9365 -24252
rect -9411 -24324 -9365 -24286
rect -9411 -24358 -9405 -24324
rect -9371 -24358 -9365 -24324
rect -9411 -24396 -9365 -24358
rect -9411 -24430 -9405 -24396
rect -9371 -24430 -9365 -24396
rect -9411 -24468 -9365 -24430
rect -9411 -24502 -9405 -24468
rect -9371 -24502 -9365 -24468
rect -9411 -24540 -9365 -24502
rect -9411 -24574 -9405 -24540
rect -9371 -24574 -9365 -24540
rect -9411 -24605 -9365 -24574
rect -8393 -24070 -8387 -24058
rect -8353 -24058 -8340 -24036
rect -7384 -24036 -7324 -23896
rect -6870 -23927 -6810 -23572
rect -6368 -23616 -6308 -23463
rect -5344 -23463 -5334 -23448
rect -5300 -23448 -5294 -23429
rect -4322 -22959 -4316 -22954
rect -4282 -22954 -4266 -22925
rect -3312 -22925 -3250 -22906
rect -3312 -22936 -3298 -22925
rect -3310 -22938 -3298 -22936
rect -4282 -22959 -4276 -22954
rect -4322 -22997 -4276 -22959
rect -4322 -23031 -4316 -22997
rect -4282 -23031 -4276 -22997
rect -4322 -23069 -4276 -23031
rect -4322 -23103 -4316 -23069
rect -4282 -23103 -4276 -23069
rect -4322 -23141 -4276 -23103
rect -4322 -23175 -4316 -23141
rect -4282 -23175 -4276 -23141
rect -4322 -23213 -4276 -23175
rect -4322 -23247 -4316 -23213
rect -4282 -23247 -4276 -23213
rect -4322 -23285 -4276 -23247
rect -4322 -23319 -4316 -23285
rect -4282 -23319 -4276 -23285
rect -4322 -23357 -4276 -23319
rect -4322 -23391 -4316 -23357
rect -4282 -23391 -4276 -23357
rect -4322 -23429 -4276 -23391
rect -4322 -23444 -4316 -23429
rect -5300 -23463 -5284 -23448
rect -6070 -23532 -5582 -23526
rect -6070 -23566 -6023 -23532
rect -5989 -23566 -5951 -23532
rect -5917 -23566 -5879 -23532
rect -5845 -23566 -5807 -23532
rect -5773 -23566 -5735 -23532
rect -5701 -23566 -5663 -23532
rect -5629 -23566 -5582 -23532
rect -6070 -23572 -5582 -23566
rect -6374 -23620 -6302 -23616
rect -6374 -23672 -6364 -23620
rect -6312 -23672 -6302 -23620
rect -6374 -23676 -6302 -23672
rect -6372 -23728 -6300 -23724
rect -6372 -23780 -6362 -23728
rect -6310 -23780 -6300 -23728
rect -6372 -23784 -6300 -23780
rect -7087 -23933 -6599 -23927
rect -7087 -23967 -7040 -23933
rect -7006 -23967 -6968 -23933
rect -6934 -23967 -6896 -23933
rect -6862 -23967 -6824 -23933
rect -6790 -23967 -6752 -23933
rect -6718 -23967 -6680 -23933
rect -6646 -23967 -6599 -23933
rect -7087 -23973 -6599 -23967
rect -7384 -24046 -7369 -24036
rect -8353 -24070 -8347 -24058
rect -8393 -24108 -8347 -24070
rect -8393 -24142 -8387 -24108
rect -8353 -24142 -8347 -24108
rect -8393 -24180 -8347 -24142
rect -8393 -24214 -8387 -24180
rect -8353 -24214 -8347 -24180
rect -8393 -24252 -8347 -24214
rect -8393 -24286 -8387 -24252
rect -8353 -24286 -8347 -24252
rect -8393 -24324 -8347 -24286
rect -8393 -24358 -8387 -24324
rect -8353 -24358 -8347 -24324
rect -8393 -24396 -8347 -24358
rect -8393 -24430 -8387 -24396
rect -8353 -24430 -8347 -24396
rect -8393 -24468 -8347 -24430
rect -8393 -24502 -8387 -24468
rect -8353 -24502 -8347 -24468
rect -8393 -24540 -8347 -24502
rect -8393 -24574 -8387 -24540
rect -8353 -24574 -8347 -24540
rect -7375 -24070 -7369 -24046
rect -7335 -24046 -7324 -24036
rect -6366 -24036 -6306 -23784
rect -5842 -23927 -5782 -23572
rect -5344 -23830 -5284 -23463
rect -4330 -23463 -4316 -23444
rect -4282 -23444 -4276 -23429
rect -3304 -22959 -3298 -22938
rect -3264 -22938 -3250 -22925
rect -3264 -22959 -3258 -22938
rect -3304 -22997 -3258 -22959
rect -3304 -23031 -3298 -22997
rect -3264 -23031 -3258 -22997
rect -3304 -23069 -3258 -23031
rect -3304 -23103 -3298 -23069
rect -3264 -23103 -3258 -23069
rect -3304 -23141 -3258 -23103
rect -3304 -23175 -3298 -23141
rect -3264 -23175 -3258 -23141
rect -3304 -23213 -3258 -23175
rect -3304 -23247 -3298 -23213
rect -3264 -23247 -3258 -23213
rect -3304 -23285 -3258 -23247
rect -3304 -23319 -3298 -23285
rect -3264 -23319 -3258 -23285
rect -3304 -23357 -3258 -23319
rect -3304 -23391 -3298 -23357
rect -3264 -23391 -3258 -23357
rect -3304 -23429 -3258 -23391
rect -4282 -23463 -4270 -23444
rect -5052 -23532 -4564 -23526
rect -5052 -23566 -5005 -23532
rect -4971 -23566 -4933 -23532
rect -4899 -23566 -4861 -23532
rect -4827 -23566 -4789 -23532
rect -4755 -23566 -4717 -23532
rect -4683 -23566 -4645 -23532
rect -4611 -23566 -4564 -23532
rect -5052 -23572 -4564 -23566
rect -5346 -23840 -5284 -23830
rect -5346 -23892 -5342 -23840
rect -5290 -23892 -5284 -23840
rect -5346 -23902 -5284 -23892
rect -6069 -23933 -5581 -23927
rect -6069 -23967 -6022 -23933
rect -5988 -23967 -5950 -23933
rect -5916 -23967 -5878 -23933
rect -5844 -23967 -5806 -23933
rect -5772 -23967 -5734 -23933
rect -5700 -23967 -5662 -23933
rect -5628 -23967 -5581 -23933
rect -6069 -23973 -5581 -23967
rect -7335 -24070 -7329 -24046
rect -6366 -24060 -6351 -24036
rect -7375 -24108 -7329 -24070
rect -7375 -24142 -7369 -24108
rect -7335 -24142 -7329 -24108
rect -7375 -24180 -7329 -24142
rect -7375 -24214 -7369 -24180
rect -7335 -24214 -7329 -24180
rect -7375 -24252 -7329 -24214
rect -7375 -24286 -7369 -24252
rect -7335 -24286 -7329 -24252
rect -7375 -24324 -7329 -24286
rect -7375 -24358 -7369 -24324
rect -7335 -24358 -7329 -24324
rect -7375 -24396 -7329 -24358
rect -7375 -24430 -7369 -24396
rect -7335 -24430 -7329 -24396
rect -7375 -24468 -7329 -24430
rect -7375 -24502 -7369 -24468
rect -7335 -24502 -7329 -24468
rect -7375 -24540 -7329 -24502
rect -7375 -24556 -7369 -24540
rect -8393 -24605 -8347 -24574
rect -7382 -24574 -7369 -24556
rect -7335 -24556 -7329 -24540
rect -6357 -24070 -6351 -24060
rect -6317 -24060 -6306 -24036
rect -5344 -24036 -5284 -23902
rect -4832 -23927 -4772 -23572
rect -4504 -23620 -4432 -23616
rect -4504 -23672 -4494 -23620
rect -4442 -23672 -4432 -23620
rect -4504 -23676 -4432 -23672
rect -4498 -23826 -4438 -23676
rect -4330 -23724 -4270 -23463
rect -3304 -23463 -3298 -23429
rect -3264 -23463 -3258 -23429
rect -3304 -23494 -3258 -23463
rect -4034 -23532 -3546 -23526
rect -4034 -23566 -3987 -23532
rect -3953 -23566 -3915 -23532
rect -3881 -23566 -3843 -23532
rect -3809 -23566 -3771 -23532
rect -3737 -23566 -3699 -23532
rect -3665 -23566 -3627 -23532
rect -3593 -23566 -3546 -23532
rect -4034 -23572 -3546 -23566
rect -4336 -23728 -4264 -23724
rect -4336 -23780 -4326 -23728
rect -4274 -23780 -4264 -23728
rect -4336 -23784 -4264 -23780
rect -4498 -23886 -3254 -23826
rect -5051 -23933 -4563 -23927
rect -5051 -23967 -5004 -23933
rect -4970 -23967 -4932 -23933
rect -4898 -23967 -4860 -23933
rect -4826 -23967 -4788 -23933
rect -4754 -23967 -4716 -23933
rect -4682 -23967 -4644 -23933
rect -4610 -23967 -4563 -23933
rect -5051 -23973 -4563 -23967
rect -5344 -24054 -5333 -24036
rect -6317 -24070 -6311 -24060
rect -6357 -24108 -6311 -24070
rect -6357 -24142 -6351 -24108
rect -6317 -24142 -6311 -24108
rect -6357 -24180 -6311 -24142
rect -6357 -24214 -6351 -24180
rect -6317 -24214 -6311 -24180
rect -6357 -24252 -6311 -24214
rect -6357 -24286 -6351 -24252
rect -6317 -24286 -6311 -24252
rect -6357 -24324 -6311 -24286
rect -6357 -24358 -6351 -24324
rect -6317 -24358 -6311 -24324
rect -6357 -24396 -6311 -24358
rect -6357 -24430 -6351 -24396
rect -6317 -24430 -6311 -24396
rect -6357 -24468 -6311 -24430
rect -6357 -24502 -6351 -24468
rect -6317 -24502 -6311 -24468
rect -6357 -24540 -6311 -24502
rect -7335 -24574 -7322 -24556
rect -9123 -24643 -8635 -24637
rect -9123 -24677 -9076 -24643
rect -9042 -24677 -9004 -24643
rect -8970 -24677 -8932 -24643
rect -8898 -24677 -8860 -24643
rect -8826 -24677 -8788 -24643
rect -8754 -24677 -8716 -24643
rect -8682 -24677 -8635 -24643
rect -9123 -24683 -8635 -24677
rect -8105 -24643 -7617 -24637
rect -8105 -24677 -8058 -24643
rect -8024 -24677 -7986 -24643
rect -7952 -24677 -7914 -24643
rect -7880 -24677 -7842 -24643
rect -7808 -24677 -7770 -24643
rect -7736 -24677 -7698 -24643
rect -7664 -24677 -7617 -24643
rect -8105 -24683 -7617 -24677
rect -8406 -24824 -8334 -24820
rect -8406 -24876 -8396 -24824
rect -8344 -24876 -8334 -24824
rect -8406 -24880 -8334 -24876
rect -12328 -24979 -12216 -24941
rect -12328 -25013 -12289 -24979
rect -12255 -25013 -12216 -24979
rect -9544 -24930 -9472 -24926
rect -9544 -24982 -9534 -24930
rect -9482 -24982 -9472 -24930
rect -9544 -24986 -9472 -24982
rect -12328 -25051 -12216 -25013
rect -12328 -25085 -12289 -25051
rect -12255 -25085 -12216 -25051
rect -12328 -25123 -12216 -25085
rect -9124 -25046 -8636 -25040
rect -9124 -25080 -9077 -25046
rect -9043 -25080 -9005 -25046
rect -8971 -25080 -8933 -25046
rect -8899 -25080 -8861 -25046
rect -8827 -25080 -8789 -25046
rect -8755 -25080 -8717 -25046
rect -8683 -25080 -8636 -25046
rect -9124 -25086 -8636 -25080
rect -12328 -25157 -12289 -25123
rect -12255 -25157 -12216 -25123
rect -12328 -25195 -12216 -25157
rect -12328 -25229 -12289 -25195
rect -12255 -25229 -12216 -25195
rect -12328 -25267 -12216 -25229
rect -12328 -25301 -12289 -25267
rect -12255 -25301 -12216 -25267
rect -12328 -25339 -12216 -25301
rect -12328 -25373 -12289 -25339
rect -12255 -25373 -12216 -25339
rect -12328 -25411 -12216 -25373
rect -12328 -25445 -12289 -25411
rect -12255 -25445 -12216 -25411
rect -12328 -25483 -12216 -25445
rect -12328 -25517 -12289 -25483
rect -12255 -25517 -12216 -25483
rect -12328 -25555 -12216 -25517
rect -12328 -25589 -12289 -25555
rect -12255 -25589 -12216 -25555
rect -12328 -25627 -12216 -25589
rect -12328 -25661 -12289 -25627
rect -12255 -25661 -12216 -25627
rect -12328 -25699 -12216 -25661
rect -9412 -25149 -9366 -25118
rect -9412 -25183 -9406 -25149
rect -9372 -25183 -9366 -25149
rect -8400 -25149 -8340 -24880
rect -7876 -25040 -7816 -24683
rect -7382 -24718 -7322 -24574
rect -6357 -24574 -6351 -24540
rect -6317 -24574 -6311 -24540
rect -5339 -24070 -5333 -24054
rect -5299 -24054 -5284 -24036
rect -4328 -24036 -4268 -23886
rect -3810 -23927 -3750 -23886
rect -4033 -23933 -3545 -23927
rect -4033 -23967 -3986 -23933
rect -3952 -23967 -3914 -23933
rect -3880 -23967 -3842 -23933
rect -3808 -23967 -3770 -23933
rect -3736 -23967 -3698 -23933
rect -3664 -23967 -3626 -23933
rect -3592 -23967 -3545 -23933
rect -4033 -23973 -3545 -23967
rect -5299 -24070 -5293 -24054
rect -4328 -24058 -4315 -24036
rect -5339 -24108 -5293 -24070
rect -5339 -24142 -5333 -24108
rect -5299 -24142 -5293 -24108
rect -5339 -24180 -5293 -24142
rect -5339 -24214 -5333 -24180
rect -5299 -24214 -5293 -24180
rect -5339 -24252 -5293 -24214
rect -5339 -24286 -5333 -24252
rect -5299 -24286 -5293 -24252
rect -5339 -24324 -5293 -24286
rect -5339 -24358 -5333 -24324
rect -5299 -24358 -5293 -24324
rect -5339 -24396 -5293 -24358
rect -5339 -24430 -5333 -24396
rect -5299 -24430 -5293 -24396
rect -5339 -24468 -5293 -24430
rect -5339 -24502 -5333 -24468
rect -5299 -24502 -5293 -24468
rect -5339 -24540 -5293 -24502
rect -5339 -24560 -5333 -24540
rect -6357 -24605 -6311 -24574
rect -5348 -24574 -5333 -24560
rect -5299 -24560 -5293 -24540
rect -4321 -24070 -4315 -24058
rect -4281 -24058 -4268 -24036
rect -3314 -24036 -3254 -23886
rect -3314 -24052 -3297 -24036
rect -4281 -24070 -4275 -24058
rect -4321 -24108 -4275 -24070
rect -4321 -24142 -4315 -24108
rect -4281 -24142 -4275 -24108
rect -4321 -24180 -4275 -24142
rect -4321 -24214 -4315 -24180
rect -4281 -24214 -4275 -24180
rect -4321 -24252 -4275 -24214
rect -4321 -24286 -4315 -24252
rect -4281 -24286 -4275 -24252
rect -4321 -24324 -4275 -24286
rect -4321 -24358 -4315 -24324
rect -4281 -24358 -4275 -24324
rect -4321 -24396 -4275 -24358
rect -4321 -24430 -4315 -24396
rect -4281 -24430 -4275 -24396
rect -4321 -24468 -4275 -24430
rect -4321 -24502 -4315 -24468
rect -4281 -24502 -4275 -24468
rect -4321 -24540 -4275 -24502
rect -5299 -24574 -5288 -24560
rect -7087 -24643 -6599 -24637
rect -7087 -24677 -7040 -24643
rect -7006 -24677 -6968 -24643
rect -6934 -24677 -6896 -24643
rect -6862 -24677 -6824 -24643
rect -6790 -24677 -6752 -24643
rect -6718 -24677 -6680 -24643
rect -6646 -24677 -6599 -24643
rect -7087 -24683 -6599 -24677
rect -6069 -24643 -5581 -24637
rect -6069 -24677 -6022 -24643
rect -5988 -24677 -5950 -24643
rect -5916 -24677 -5878 -24643
rect -5844 -24677 -5806 -24643
rect -5772 -24677 -5734 -24643
rect -5700 -24677 -5662 -24643
rect -5628 -24677 -5581 -24643
rect -6069 -24683 -5581 -24677
rect -7388 -24722 -7316 -24718
rect -7388 -24774 -7378 -24722
rect -7326 -24774 -7316 -24722
rect -7388 -24778 -7316 -24774
rect -8106 -25046 -7618 -25040
rect -8106 -25080 -8059 -25046
rect -8025 -25080 -7987 -25046
rect -7953 -25080 -7915 -25046
rect -7881 -25080 -7843 -25046
rect -7809 -25080 -7771 -25046
rect -7737 -25080 -7699 -25046
rect -7665 -25080 -7618 -25046
rect -8106 -25086 -7618 -25080
rect -8400 -25174 -8388 -25149
rect -9412 -25221 -9366 -25183
rect -9412 -25255 -9406 -25221
rect -9372 -25255 -9366 -25221
rect -9412 -25293 -9366 -25255
rect -9412 -25327 -9406 -25293
rect -9372 -25327 -9366 -25293
rect -9412 -25365 -9366 -25327
rect -9412 -25399 -9406 -25365
rect -9372 -25399 -9366 -25365
rect -9412 -25437 -9366 -25399
rect -9412 -25471 -9406 -25437
rect -9372 -25471 -9366 -25437
rect -9412 -25509 -9366 -25471
rect -9412 -25543 -9406 -25509
rect -9372 -25543 -9366 -25509
rect -9412 -25581 -9366 -25543
rect -9412 -25615 -9406 -25581
rect -9372 -25615 -9366 -25581
rect -9412 -25653 -9366 -25615
rect -9412 -25666 -9406 -25653
rect -12328 -25733 -12289 -25699
rect -12255 -25733 -12216 -25699
rect -12328 -25771 -12216 -25733
rect -12328 -25805 -12289 -25771
rect -12255 -25805 -12216 -25771
rect -12328 -25843 -12216 -25805
rect -12328 -25877 -12289 -25843
rect -12255 -25877 -12216 -25843
rect -12328 -25915 -12216 -25877
rect -12328 -25949 -12289 -25915
rect -12255 -25949 -12216 -25915
rect -9418 -25687 -9406 -25666
rect -9372 -25666 -9366 -25653
rect -8394 -25183 -8388 -25174
rect -8354 -25174 -8340 -25149
rect -7382 -25149 -7322 -24778
rect -6876 -25040 -6816 -24683
rect -6372 -24930 -6300 -24926
rect -6372 -24982 -6362 -24930
rect -6310 -24982 -6300 -24930
rect -6372 -24986 -6300 -24982
rect -7088 -25046 -6600 -25040
rect -7088 -25080 -7041 -25046
rect -7007 -25080 -6969 -25046
rect -6935 -25080 -6897 -25046
rect -6863 -25080 -6825 -25046
rect -6791 -25080 -6753 -25046
rect -6719 -25080 -6681 -25046
rect -6647 -25080 -6600 -25046
rect -7088 -25086 -6600 -25080
rect -8354 -25183 -8348 -25174
rect -8394 -25221 -8348 -25183
rect -8394 -25255 -8388 -25221
rect -8354 -25255 -8348 -25221
rect -8394 -25293 -8348 -25255
rect -8394 -25327 -8388 -25293
rect -8354 -25327 -8348 -25293
rect -8394 -25365 -8348 -25327
rect -8394 -25399 -8388 -25365
rect -8354 -25399 -8348 -25365
rect -8394 -25437 -8348 -25399
rect -8394 -25471 -8388 -25437
rect -8354 -25471 -8348 -25437
rect -8394 -25509 -8348 -25471
rect -8394 -25543 -8388 -25509
rect -8354 -25543 -8348 -25509
rect -8394 -25581 -8348 -25543
rect -8394 -25615 -8388 -25581
rect -8354 -25615 -8348 -25581
rect -8394 -25653 -8348 -25615
rect -9372 -25687 -9358 -25666
rect -8394 -25672 -8388 -25653
rect -9418 -25870 -9358 -25687
rect -8402 -25687 -8388 -25672
rect -8354 -25672 -8348 -25653
rect -7382 -25183 -7370 -25149
rect -7336 -25183 -7322 -25149
rect -6366 -25149 -6306 -24986
rect -5852 -25040 -5792 -24683
rect -5348 -24712 -5288 -24574
rect -4321 -24574 -4315 -24540
rect -4281 -24574 -4275 -24540
rect -4321 -24605 -4275 -24574
rect -3303 -24070 -3297 -24052
rect -3263 -24052 -3254 -24036
rect -3263 -24070 -3257 -24052
rect -3303 -24108 -3257 -24070
rect -3303 -24142 -3297 -24108
rect -3263 -24142 -3257 -24108
rect -3303 -24180 -3257 -24142
rect -3303 -24214 -3297 -24180
rect -3263 -24214 -3257 -24180
rect -3303 -24252 -3257 -24214
rect -3303 -24286 -3297 -24252
rect -3263 -24286 -3257 -24252
rect -3303 -24324 -3257 -24286
rect -3303 -24358 -3297 -24324
rect -3263 -24358 -3257 -24324
rect -3303 -24396 -3257 -24358
rect -3303 -24430 -3297 -24396
rect -3263 -24430 -3257 -24396
rect -3303 -24468 -3257 -24430
rect -3303 -24502 -3297 -24468
rect -3263 -24502 -3257 -24468
rect -3303 -24540 -3257 -24502
rect -3303 -24574 -3297 -24540
rect -3263 -24574 -3257 -24540
rect -3303 -24605 -3257 -24574
rect -5051 -24643 -4563 -24637
rect -5051 -24677 -5004 -24643
rect -4970 -24677 -4932 -24643
rect -4898 -24677 -4860 -24643
rect -4826 -24677 -4788 -24643
rect -4754 -24677 -4716 -24643
rect -4682 -24677 -4644 -24643
rect -4610 -24677 -4563 -24643
rect -5051 -24683 -4563 -24677
rect -4033 -24643 -3545 -24637
rect -4033 -24677 -3986 -24643
rect -3952 -24677 -3914 -24643
rect -3880 -24677 -3842 -24643
rect -3808 -24677 -3770 -24643
rect -3736 -24677 -3698 -24643
rect -3664 -24677 -3626 -24643
rect -3592 -24677 -3545 -24643
rect -4033 -24683 -3545 -24677
rect -5352 -24722 -5288 -24712
rect -5352 -24774 -5348 -24722
rect -5296 -24774 -5288 -24722
rect -5352 -24784 -5288 -24774
rect -6070 -25046 -5582 -25040
rect -6070 -25080 -6023 -25046
rect -5989 -25080 -5951 -25046
rect -5917 -25080 -5879 -25046
rect -5845 -25080 -5807 -25046
rect -5773 -25080 -5735 -25046
rect -5701 -25080 -5663 -25046
rect -5629 -25080 -5582 -25046
rect -6070 -25086 -5582 -25080
rect -6366 -25182 -6352 -25149
rect -7382 -25221 -7322 -25183
rect -7382 -25255 -7370 -25221
rect -7336 -25255 -7322 -25221
rect -7382 -25293 -7322 -25255
rect -7382 -25327 -7370 -25293
rect -7336 -25327 -7322 -25293
rect -7382 -25365 -7322 -25327
rect -7382 -25399 -7370 -25365
rect -7336 -25399 -7322 -25365
rect -7382 -25437 -7322 -25399
rect -7382 -25471 -7370 -25437
rect -7336 -25471 -7322 -25437
rect -7382 -25509 -7322 -25471
rect -7382 -25543 -7370 -25509
rect -7336 -25543 -7322 -25509
rect -7382 -25581 -7322 -25543
rect -7382 -25615 -7370 -25581
rect -7336 -25615 -7322 -25581
rect -7382 -25653 -7322 -25615
rect -8354 -25687 -8342 -25672
rect -9124 -25756 -8636 -25750
rect -9124 -25790 -9077 -25756
rect -9043 -25790 -9005 -25756
rect -8971 -25790 -8933 -25756
rect -8899 -25790 -8861 -25756
rect -8827 -25790 -8789 -25756
rect -8755 -25790 -8717 -25756
rect -8683 -25790 -8636 -25756
rect -9124 -25796 -8636 -25790
rect -8910 -25870 -8850 -25796
rect -8402 -25870 -8342 -25687
rect -7382 -25687 -7370 -25653
rect -7336 -25687 -7322 -25653
rect -8106 -25756 -7618 -25750
rect -8106 -25790 -8059 -25756
rect -8025 -25790 -7987 -25756
rect -7953 -25790 -7915 -25756
rect -7881 -25790 -7843 -25756
rect -7809 -25790 -7771 -25756
rect -7737 -25790 -7699 -25756
rect -7665 -25790 -7618 -25756
rect -8106 -25796 -7618 -25790
rect -7896 -25870 -7836 -25796
rect -9418 -25874 -7830 -25870
rect -9418 -25926 -7892 -25874
rect -7840 -25926 -7830 -25874
rect -9418 -25930 -7830 -25926
rect -12328 -25987 -12216 -25949
rect -12328 -26021 -12289 -25987
rect -12255 -26021 -12216 -25987
rect -12328 -26059 -12216 -26021
rect -12328 -26093 -12289 -26059
rect -12255 -26093 -12216 -26059
rect -12328 -26131 -12216 -26093
rect -12328 -26165 -12289 -26131
rect -12255 -26165 -12216 -26131
rect -12328 -26203 -12216 -26165
rect -12328 -26237 -12289 -26203
rect -12255 -26237 -12216 -26203
rect -12328 -26275 -12216 -26237
rect -12328 -26309 -12289 -26275
rect -12255 -26309 -12216 -26275
rect -12328 -26816 -12216 -26309
rect -7382 -26430 -7322 -25687
rect -6358 -25183 -6352 -25182
rect -6318 -25182 -6306 -25149
rect -5348 -25149 -5288 -24784
rect -4836 -25040 -4776 -24683
rect -3202 -24820 -3142 -22776
rect -2670 -23620 -2610 -21640
rect -2538 -22614 -2478 -21400
rect -2122 -21484 -2062 -21474
rect 952 -21480 1012 -18914
rect -2122 -21534 -2118 -21484
rect -2124 -21536 -2118 -21534
rect -2066 -21536 -2062 -21484
rect -2124 -21575 -2062 -21536
rect -938 -21484 -866 -21480
rect -938 -21536 -928 -21484
rect -876 -21536 -866 -21484
rect -938 -21540 -866 -21536
rect 256 -21484 328 -21480
rect 256 -21536 266 -21484
rect 318 -21536 328 -21484
rect 256 -21540 328 -21536
rect 946 -21484 1018 -21480
rect 946 -21536 956 -21484
rect 1008 -21536 1018 -21484
rect 946 -21540 1018 -21536
rect -2427 -21637 -2062 -21575
rect -2427 -21792 -2365 -21637
rect -2275 -21702 -2213 -21637
rect -2308 -21708 -2180 -21702
rect -2308 -21742 -2261 -21708
rect -2227 -21742 -2180 -21708
rect -2308 -21748 -2180 -21742
rect -2427 -21811 -2362 -21792
rect -2427 -21825 -2410 -21811
rect -2416 -21845 -2410 -21825
rect -2376 -21824 -2362 -21811
rect -2124 -21811 -2062 -21637
rect -1684 -21584 -1612 -21580
rect -1684 -21636 -1674 -21584
rect -1622 -21636 -1612 -21584
rect -1684 -21640 -1612 -21636
rect -1386 -21584 -1314 -21580
rect -1386 -21636 -1376 -21584
rect -1324 -21636 -1314 -21584
rect -1386 -21640 -1314 -21636
rect -1678 -21702 -1618 -21640
rect -1380 -21702 -1320 -21640
rect -2010 -21708 -1882 -21702
rect -2010 -21742 -1963 -21708
rect -1929 -21742 -1882 -21708
rect -2010 -21748 -1882 -21742
rect -1712 -21708 -1584 -21702
rect -1712 -21742 -1665 -21708
rect -1631 -21742 -1584 -21708
rect -1712 -21748 -1584 -21742
rect -1414 -21708 -1286 -21702
rect -1414 -21742 -1367 -21708
rect -1333 -21742 -1286 -21708
rect -1414 -21748 -1286 -21742
rect -1116 -21708 -988 -21702
rect -1116 -21742 -1069 -21708
rect -1035 -21742 -988 -21708
rect -1116 -21748 -988 -21742
rect -2376 -21825 -2365 -21824
rect -2376 -21845 -2370 -21825
rect -2124 -21832 -2112 -21811
rect -2122 -21844 -2112 -21832
rect -2416 -21883 -2370 -21845
rect -2416 -21917 -2410 -21883
rect -2376 -21917 -2370 -21883
rect -2416 -21955 -2370 -21917
rect -2416 -21989 -2410 -21955
rect -2376 -21989 -2370 -21955
rect -2416 -22027 -2370 -21989
rect -2416 -22061 -2410 -22027
rect -2376 -22061 -2370 -22027
rect -2416 -22099 -2370 -22061
rect -2416 -22133 -2410 -22099
rect -2376 -22133 -2370 -22099
rect -2416 -22171 -2370 -22133
rect -2416 -22205 -2410 -22171
rect -2376 -22205 -2370 -22171
rect -2416 -22243 -2370 -22205
rect -2416 -22277 -2410 -22243
rect -2376 -22277 -2370 -22243
rect -2416 -22315 -2370 -22277
rect -2416 -22349 -2410 -22315
rect -2376 -22349 -2370 -22315
rect -2416 -22380 -2370 -22349
rect -2118 -21845 -2112 -21844
rect -2078 -21844 -2062 -21811
rect -1814 -21811 -1780 -21792
rect -2078 -21845 -2072 -21844
rect -2118 -21883 -2072 -21845
rect -2118 -21917 -2112 -21883
rect -2078 -21917 -2072 -21883
rect -2118 -21955 -2072 -21917
rect -2118 -21989 -2112 -21955
rect -2078 -21989 -2072 -21955
rect -2118 -22027 -2072 -21989
rect -2118 -22061 -2112 -22027
rect -2078 -22061 -2072 -22027
rect -2118 -22099 -2072 -22061
rect -2118 -22133 -2112 -22099
rect -2078 -22133 -2072 -22099
rect -2118 -22171 -2072 -22133
rect -2118 -22205 -2112 -22171
rect -2078 -22205 -2072 -22171
rect -2118 -22243 -2072 -22205
rect -2118 -22277 -2112 -22243
rect -2078 -22277 -2072 -22243
rect -2118 -22315 -2072 -22277
rect -2118 -22349 -2112 -22315
rect -2078 -22349 -2072 -22315
rect -1820 -21845 -1814 -21832
rect -1522 -21811 -1476 -21780
rect -1780 -21845 -1774 -21832
rect -1820 -21883 -1774 -21845
rect -1820 -21917 -1814 -21883
rect -1780 -21917 -1774 -21883
rect -1820 -21955 -1774 -21917
rect -1820 -21989 -1814 -21955
rect -1780 -21989 -1774 -21955
rect -1820 -22027 -1774 -21989
rect -1820 -22061 -1814 -22027
rect -1780 -22061 -1774 -22027
rect -1820 -22099 -1774 -22061
rect -1820 -22133 -1814 -22099
rect -1780 -22133 -1774 -22099
rect -1820 -22171 -1774 -22133
rect -1820 -22205 -1814 -22171
rect -1780 -22205 -1774 -22171
rect -1820 -22243 -1774 -22205
rect -1820 -22277 -1814 -22243
rect -1780 -22277 -1774 -22243
rect -1820 -22315 -1774 -22277
rect -1522 -21845 -1516 -21811
rect -1482 -21845 -1476 -21811
rect -1522 -21883 -1476 -21845
rect -1522 -21917 -1516 -21883
rect -1482 -21917 -1476 -21883
rect -1522 -21955 -1476 -21917
rect -1522 -21989 -1516 -21955
rect -1482 -21989 -1476 -21955
rect -1522 -22027 -1476 -21989
rect -1522 -22061 -1516 -22027
rect -1482 -22061 -1476 -22027
rect -1522 -22099 -1476 -22061
rect -1522 -22133 -1516 -22099
rect -1482 -22133 -1476 -22099
rect -1522 -22171 -1476 -22133
rect -1522 -22205 -1516 -22171
rect -1482 -22205 -1476 -22171
rect -1522 -22243 -1476 -22205
rect -1522 -22277 -1516 -22243
rect -1482 -22277 -1476 -22243
rect -1522 -22312 -1476 -22277
rect -1224 -21811 -1178 -21786
rect -1224 -21845 -1218 -21811
rect -1184 -21845 -1178 -21811
rect -1224 -21883 -1178 -21845
rect -932 -21811 -872 -21540
rect -490 -21584 -418 -21580
rect -490 -21636 -480 -21584
rect -428 -21636 -418 -21584
rect -490 -21640 -418 -21636
rect -194 -21584 -122 -21580
rect -194 -21636 -184 -21584
rect -132 -21636 -122 -21584
rect -194 -21640 -122 -21636
rect -484 -21702 -424 -21640
rect -188 -21702 -128 -21640
rect -818 -21708 -690 -21702
rect -818 -21742 -771 -21708
rect -737 -21742 -690 -21708
rect -818 -21748 -690 -21742
rect -520 -21708 -392 -21702
rect -520 -21742 -473 -21708
rect -439 -21742 -392 -21708
rect -520 -21748 -392 -21742
rect -222 -21708 -94 -21702
rect -222 -21742 -175 -21708
rect -141 -21742 -94 -21708
rect -222 -21748 -94 -21742
rect 76 -21708 204 -21702
rect 76 -21742 123 -21708
rect 157 -21742 204 -21708
rect 76 -21748 204 -21742
rect -932 -21845 -920 -21811
rect -886 -21845 -872 -21811
rect -932 -21852 -872 -21845
rect -622 -21811 -588 -21792
rect -1224 -21917 -1218 -21883
rect -1184 -21917 -1178 -21883
rect -1224 -21955 -1178 -21917
rect -1224 -21989 -1218 -21955
rect -1184 -21989 -1178 -21955
rect -1224 -22027 -1178 -21989
rect -1224 -22061 -1218 -22027
rect -1184 -22061 -1178 -22027
rect -1224 -22099 -1178 -22061
rect -1224 -22133 -1218 -22099
rect -1184 -22133 -1178 -22099
rect -1224 -22171 -1178 -22133
rect -1224 -22205 -1218 -22171
rect -1184 -22205 -1178 -22171
rect -1224 -22243 -1178 -22205
rect -1224 -22277 -1218 -22243
rect -1184 -22277 -1178 -22243
rect -1820 -22319 -1814 -22315
rect -2118 -22380 -2072 -22349
rect -1829 -22349 -1814 -22319
rect -1780 -22319 -1774 -22315
rect -1530 -22315 -1470 -22312
rect -1780 -22349 -1771 -22319
rect -1530 -22332 -1516 -22315
rect -2308 -22418 -2180 -22412
rect -2308 -22452 -2261 -22418
rect -2227 -22452 -2180 -22418
rect -1998 -22452 -1963 -22418
rect -1929 -22452 -1894 -22418
rect -2308 -22458 -2180 -22452
rect -2548 -22618 -2476 -22614
rect -2548 -22670 -2538 -22618
rect -2486 -22670 -2476 -22618
rect -2548 -22674 -2476 -22670
rect -2126 -22618 -2066 -22608
rect -2126 -22670 -2122 -22618
rect -2070 -22664 -2066 -22618
rect -2070 -22670 -2064 -22664
rect -2126 -22704 -2064 -22670
rect -2422 -22764 -2064 -22704
rect -1974 -22722 -1914 -22452
rect -1829 -22483 -1771 -22349
rect -1532 -22349 -1516 -22332
rect -1482 -22349 -1470 -22315
rect -1532 -22368 -1470 -22349
rect -1224 -22315 -1178 -22277
rect -1224 -22349 -1218 -22315
rect -1184 -22349 -1178 -22315
rect -1224 -22354 -1178 -22349
rect -926 -21883 -880 -21852
rect -622 -21878 -588 -21845
rect -330 -21811 -284 -21780
rect -330 -21845 -324 -21811
rect -290 -21845 -284 -21811
rect -926 -21917 -920 -21883
rect -886 -21917 -880 -21883
rect -926 -21955 -880 -21917
rect -926 -21989 -920 -21955
rect -886 -21989 -880 -21955
rect -926 -22027 -880 -21989
rect -926 -22061 -920 -22027
rect -886 -22061 -880 -22027
rect -926 -22099 -880 -22061
rect -926 -22133 -920 -22099
rect -886 -22133 -880 -22099
rect -926 -22171 -880 -22133
rect -926 -22205 -920 -22171
rect -886 -22205 -880 -22171
rect -926 -22243 -880 -22205
rect -926 -22277 -920 -22243
rect -886 -22277 -880 -22243
rect -926 -22315 -880 -22277
rect -926 -22349 -920 -22315
rect -886 -22349 -880 -22315
rect -628 -21883 -582 -21878
rect -628 -21917 -622 -21883
rect -588 -21917 -582 -21883
rect -628 -21955 -582 -21917
rect -628 -21989 -622 -21955
rect -588 -21989 -582 -21955
rect -628 -22027 -582 -21989
rect -628 -22061 -622 -22027
rect -588 -22061 -582 -22027
rect -628 -22099 -582 -22061
rect -628 -22133 -622 -22099
rect -588 -22133 -582 -22099
rect -628 -22171 -582 -22133
rect -628 -22205 -622 -22171
rect -588 -22205 -582 -22171
rect -628 -22243 -582 -22205
rect -628 -22277 -622 -22243
rect -588 -22277 -582 -22243
rect -628 -22315 -582 -22277
rect -330 -21883 -284 -21845
rect -26 -21811 8 -21792
rect -26 -21878 8 -21845
rect 262 -21811 322 -21540
rect 374 -21708 502 -21702
rect 374 -21742 421 -21708
rect 455 -21742 502 -21708
rect 374 -21748 502 -21742
rect 672 -21708 800 -21702
rect 672 -21742 719 -21708
rect 753 -21742 800 -21708
rect 672 -21748 800 -21742
rect 262 -21845 272 -21811
rect 306 -21845 322 -21811
rect 262 -21848 322 -21845
rect 564 -21811 610 -21780
rect 564 -21845 570 -21811
rect 604 -21845 610 -21811
rect -330 -21917 -324 -21883
rect -290 -21917 -284 -21883
rect -330 -21955 -284 -21917
rect -330 -21989 -324 -21955
rect -290 -21989 -284 -21955
rect -330 -22027 -284 -21989
rect -330 -22061 -324 -22027
rect -290 -22061 -284 -22027
rect -330 -22099 -284 -22061
rect -330 -22133 -324 -22099
rect -290 -22133 -284 -22099
rect -330 -22171 -284 -22133
rect -330 -22205 -324 -22171
rect -290 -22205 -284 -22171
rect -330 -22243 -284 -22205
rect -330 -22277 -324 -22243
rect -290 -22277 -284 -22243
rect -330 -22310 -284 -22277
rect -32 -21883 14 -21878
rect -32 -21917 -26 -21883
rect 8 -21917 14 -21883
rect -32 -21955 14 -21917
rect -32 -21989 -26 -21955
rect 8 -21989 14 -21955
rect -32 -22027 14 -21989
rect -32 -22061 -26 -22027
rect 8 -22061 14 -22027
rect -32 -22099 14 -22061
rect -32 -22133 -26 -22099
rect 8 -22133 14 -22099
rect -32 -22171 14 -22133
rect -32 -22205 -26 -22171
rect 8 -22205 14 -22171
rect -32 -22243 14 -22205
rect -32 -22277 -26 -22243
rect 8 -22277 14 -22243
rect -628 -22345 -622 -22315
rect -1230 -22361 -1170 -22354
rect -1712 -22418 -1584 -22412
rect -1712 -22452 -1665 -22418
rect -1631 -22452 -1584 -22418
rect -1712 -22458 -1584 -22452
rect -1835 -22486 -1765 -22483
rect -1835 -22538 -1826 -22486
rect -1774 -22538 -1765 -22486
rect -1835 -22541 -1765 -22538
rect -2422 -22923 -2362 -22764
rect -2274 -22814 -2214 -22764
rect -2308 -22820 -2180 -22814
rect -2308 -22854 -2261 -22820
rect -2227 -22854 -2180 -22820
rect -2308 -22860 -2180 -22854
rect -2422 -22952 -2410 -22923
rect -2416 -22957 -2410 -22952
rect -2376 -22952 -2362 -22923
rect -2126 -22923 -2064 -22764
rect -1980 -22726 -1908 -22722
rect -1980 -22778 -1970 -22726
rect -1918 -22778 -1908 -22726
rect -1980 -22782 -1908 -22778
rect -2010 -22820 -1882 -22814
rect -2010 -22854 -1963 -22820
rect -1929 -22854 -1882 -22820
rect -2010 -22860 -1882 -22854
rect -2126 -22942 -2112 -22923
rect -2376 -22957 -2370 -22952
rect -2124 -22954 -2112 -22942
rect -2416 -22995 -2370 -22957
rect -2416 -23029 -2410 -22995
rect -2376 -23029 -2370 -22995
rect -2416 -23067 -2370 -23029
rect -2416 -23101 -2410 -23067
rect -2376 -23101 -2370 -23067
rect -2416 -23139 -2370 -23101
rect -2416 -23173 -2410 -23139
rect -2376 -23173 -2370 -23139
rect -2416 -23211 -2370 -23173
rect -2416 -23245 -2410 -23211
rect -2376 -23245 -2370 -23211
rect -2416 -23283 -2370 -23245
rect -2416 -23317 -2410 -23283
rect -2376 -23317 -2370 -23283
rect -2416 -23355 -2370 -23317
rect -2416 -23389 -2410 -23355
rect -2376 -23389 -2370 -23355
rect -2416 -23427 -2370 -23389
rect -2416 -23461 -2410 -23427
rect -2376 -23461 -2370 -23427
rect -2118 -22957 -2112 -22954
rect -2078 -22954 -2064 -22923
rect -1829 -22923 -1771 -22541
rect -1532 -22614 -1472 -22368
rect -1414 -22418 -1286 -22412
rect -1414 -22452 -1367 -22418
rect -1333 -22452 -1286 -22418
rect -1414 -22458 -1286 -22452
rect -1230 -22483 -1167 -22361
rect -926 -22380 -880 -22349
rect -634 -22349 -622 -22345
rect -588 -22345 -582 -22315
rect -338 -22315 -278 -22310
rect -338 -22326 -324 -22315
rect -588 -22349 -576 -22345
rect -1116 -22418 -988 -22412
rect -1116 -22452 -1069 -22418
rect -1035 -22452 -988 -22418
rect -1116 -22458 -988 -22452
rect -818 -22418 -690 -22412
rect -818 -22452 -771 -22418
rect -737 -22452 -690 -22418
rect -818 -22458 -690 -22452
rect -1231 -22486 -1161 -22483
rect -1231 -22538 -1222 -22486
rect -1170 -22538 -1161 -22486
rect -1231 -22541 -1161 -22538
rect -1538 -22618 -1466 -22614
rect -1538 -22670 -1528 -22618
rect -1476 -22670 -1466 -22618
rect -1538 -22674 -1466 -22670
rect -1682 -22726 -1610 -22722
rect -1682 -22778 -1672 -22726
rect -1620 -22778 -1610 -22726
rect -1682 -22782 -1610 -22778
rect -1382 -22726 -1310 -22722
rect -1382 -22778 -1372 -22726
rect -1320 -22778 -1310 -22726
rect -1382 -22782 -1310 -22778
rect -1676 -22814 -1616 -22782
rect -1376 -22814 -1316 -22782
rect -1704 -22820 -1584 -22814
rect -1704 -22854 -1665 -22820
rect -1631 -22854 -1584 -22820
rect -1704 -22860 -1584 -22854
rect -1414 -22820 -1286 -22814
rect -1414 -22854 -1367 -22820
rect -1333 -22854 -1286 -22820
rect -1414 -22860 -1286 -22854
rect -1829 -22935 -1814 -22923
rect -2078 -22957 -2072 -22954
rect -2118 -22995 -2072 -22957
rect -2118 -23029 -2112 -22995
rect -2078 -23029 -2072 -22995
rect -1780 -22935 -1771 -22923
rect -1522 -22923 -1476 -22892
rect -1230 -22917 -1167 -22541
rect -1082 -22722 -1022 -22458
rect -940 -22618 -868 -22614
rect -940 -22670 -930 -22618
rect -878 -22670 -868 -22618
rect -940 -22674 -868 -22670
rect -1088 -22726 -1016 -22722
rect -1088 -22778 -1078 -22726
rect -1026 -22778 -1016 -22726
rect -1088 -22782 -1016 -22778
rect -1116 -22820 -988 -22814
rect -1116 -22854 -1069 -22820
rect -1035 -22854 -988 -22820
rect -1116 -22860 -988 -22854
rect -1814 -22995 -1780 -22957
rect -2118 -23067 -2072 -23029
rect -2118 -23101 -2112 -23067
rect -2078 -23101 -2072 -23067
rect -2118 -23139 -2072 -23101
rect -2118 -23173 -2112 -23139
rect -2078 -23173 -2072 -23139
rect -2118 -23211 -2072 -23173
rect -2118 -23245 -2112 -23211
rect -2078 -23245 -2072 -23211
rect -2118 -23283 -2072 -23245
rect -2118 -23317 -2112 -23283
rect -2078 -23317 -2072 -23283
rect -2118 -23355 -2072 -23317
rect -2118 -23389 -2112 -23355
rect -2078 -23389 -2072 -23355
rect -2118 -23427 -2072 -23389
rect -2118 -23440 -2112 -23427
rect -2416 -23492 -2370 -23461
rect -2126 -23461 -2112 -23440
rect -2078 -23440 -2072 -23427
rect -1820 -23029 -1814 -23002
rect -1522 -22957 -1516 -22923
rect -1482 -22957 -1476 -22923
rect -1522 -22995 -1476 -22957
rect -1218 -22923 -1184 -22917
rect -934 -22923 -874 -22674
rect -786 -22722 -726 -22458
rect -634 -22483 -576 -22349
rect -340 -22349 -324 -22326
rect -290 -22349 -278 -22315
rect -32 -22315 14 -22277
rect -32 -22317 -26 -22315
rect -37 -22338 -26 -22317
rect -340 -22368 -278 -22349
rect -38 -22349 -26 -22338
rect 8 -22317 14 -22315
rect 266 -21883 312 -21848
rect 266 -21917 272 -21883
rect 306 -21917 312 -21883
rect 266 -21955 312 -21917
rect 266 -21989 272 -21955
rect 306 -21989 312 -21955
rect 266 -22027 312 -21989
rect 266 -22061 272 -22027
rect 306 -22061 312 -22027
rect 266 -22099 312 -22061
rect 266 -22133 272 -22099
rect 306 -22133 312 -22099
rect 266 -22171 312 -22133
rect 266 -22205 272 -22171
rect 306 -22205 312 -22171
rect 266 -22243 312 -22205
rect 266 -22277 272 -22243
rect 306 -22277 312 -22243
rect 266 -22315 312 -22277
rect 8 -22338 21 -22317
rect 8 -22349 22 -22338
rect -520 -22418 -392 -22412
rect -520 -22452 -473 -22418
rect -439 -22452 -392 -22418
rect -520 -22458 -392 -22452
rect -640 -22486 -570 -22483
rect -640 -22538 -631 -22486
rect -579 -22538 -570 -22486
rect -640 -22541 -570 -22538
rect -792 -22726 -720 -22722
rect -792 -22778 -782 -22726
rect -730 -22778 -720 -22726
rect -792 -22782 -720 -22778
rect -818 -22820 -690 -22814
rect -818 -22854 -771 -22820
rect -737 -22854 -690 -22820
rect -818 -22860 -690 -22854
rect -934 -22954 -920 -22923
rect -1218 -22962 -1184 -22957
rect -926 -22957 -920 -22954
rect -886 -22954 -874 -22923
rect -634 -22904 -576 -22541
rect -340 -22614 -280 -22368
rect -222 -22418 -94 -22412
rect -222 -22452 -175 -22418
rect -141 -22452 -94 -22418
rect -222 -22458 -94 -22452
rect -38 -22486 22 -22349
rect 266 -22349 272 -22315
rect 306 -22349 312 -22315
rect 564 -21883 610 -21845
rect 564 -21917 570 -21883
rect 604 -21917 610 -21883
rect 564 -21955 610 -21917
rect 564 -21989 570 -21955
rect 604 -21989 610 -21955
rect 564 -22027 610 -21989
rect 564 -22061 570 -22027
rect 604 -22061 610 -22027
rect 564 -22099 610 -22061
rect 564 -22133 570 -22099
rect 604 -22133 610 -22099
rect 564 -22171 610 -22133
rect 564 -22205 570 -22171
rect 604 -22205 610 -22171
rect 564 -22243 610 -22205
rect 564 -22277 570 -22243
rect 604 -22277 610 -22243
rect 564 -22315 610 -22277
rect 564 -22323 570 -22315
rect 559 -22330 570 -22323
rect 266 -22380 312 -22349
rect 556 -22349 570 -22330
rect 604 -22323 610 -22315
rect 862 -21811 908 -21780
rect 862 -21845 868 -21811
rect 902 -21845 908 -21811
rect 862 -21883 908 -21845
rect 862 -21917 868 -21883
rect 902 -21917 908 -21883
rect 862 -21955 908 -21917
rect 862 -21989 868 -21955
rect 902 -21989 908 -21955
rect 862 -22027 908 -21989
rect 862 -22061 868 -22027
rect 902 -22061 908 -22027
rect 862 -22099 908 -22061
rect 862 -22133 868 -22099
rect 902 -22133 908 -22099
rect 862 -22171 908 -22133
rect 862 -22205 868 -22171
rect 902 -22205 908 -22171
rect 862 -22243 908 -22205
rect 862 -22277 868 -22243
rect 902 -22277 908 -22243
rect 862 -22315 908 -22277
rect 604 -22349 617 -22323
rect 862 -22328 868 -22315
rect 76 -22418 204 -22412
rect 76 -22452 123 -22418
rect 157 -22452 204 -22418
rect 76 -22458 204 -22452
rect 374 -22418 502 -22412
rect 374 -22452 421 -22418
rect 455 -22452 502 -22418
rect 374 -22458 502 -22452
rect -38 -22538 -34 -22486
rect 18 -22538 22 -22486
rect -346 -22618 -274 -22614
rect -346 -22670 -336 -22618
rect -284 -22670 -274 -22618
rect -346 -22674 -274 -22670
rect -492 -22726 -420 -22722
rect -492 -22778 -482 -22726
rect -430 -22778 -420 -22726
rect -492 -22782 -420 -22778
rect -190 -22726 -118 -22722
rect -190 -22778 -180 -22726
rect -128 -22778 -118 -22726
rect -190 -22782 -118 -22778
rect -486 -22814 -426 -22782
rect -184 -22814 -124 -22782
rect -520 -22820 -392 -22814
rect -520 -22854 -473 -22820
rect -439 -22854 -392 -22820
rect -520 -22860 -392 -22854
rect -222 -22820 -94 -22814
rect -222 -22854 -175 -22820
rect -141 -22854 -94 -22820
rect -222 -22860 -94 -22854
rect -634 -22923 -572 -22904
rect -634 -22933 -622 -22923
rect -886 -22957 -880 -22954
rect -1780 -23029 -1774 -23002
rect -1820 -23067 -1774 -23029
rect -1820 -23101 -1814 -23067
rect -1780 -23101 -1774 -23067
rect -1820 -23139 -1774 -23101
rect -1820 -23173 -1814 -23139
rect -1780 -23173 -1774 -23139
rect -1820 -23211 -1774 -23173
rect -1820 -23245 -1814 -23211
rect -1780 -23245 -1774 -23211
rect -1820 -23283 -1774 -23245
rect -1820 -23317 -1814 -23283
rect -1780 -23317 -1774 -23283
rect -1820 -23355 -1774 -23317
rect -1820 -23389 -1814 -23355
rect -1780 -23389 -1774 -23355
rect -1820 -23427 -1774 -23389
rect -1820 -23440 -1814 -23427
rect -2078 -23461 -2066 -23440
rect -2308 -23530 -2180 -23524
rect -2308 -23564 -2261 -23530
rect -2227 -23564 -2180 -23530
rect -2308 -23570 -2180 -23564
rect -2676 -23624 -2604 -23620
rect -2676 -23676 -2666 -23624
rect -2614 -23676 -2604 -23624
rect -2676 -23680 -2604 -23676
rect -4338 -24824 -4266 -24820
rect -4338 -24876 -4328 -24824
rect -4276 -24876 -4266 -24824
rect -4338 -24880 -4266 -24876
rect -3208 -24824 -3136 -24820
rect -3208 -24876 -3198 -24824
rect -3146 -24876 -3136 -24824
rect -3208 -24880 -3136 -24876
rect -5052 -25046 -4564 -25040
rect -5052 -25080 -5005 -25046
rect -4971 -25080 -4933 -25046
rect -4899 -25080 -4861 -25046
rect -4827 -25080 -4789 -25046
rect -4755 -25080 -4717 -25046
rect -4683 -25080 -4645 -25046
rect -4611 -25080 -4564 -25046
rect -5052 -25086 -4564 -25080
rect -6318 -25183 -6312 -25182
rect -6358 -25221 -6312 -25183
rect -6358 -25255 -6352 -25221
rect -6318 -25255 -6312 -25221
rect -6358 -25293 -6312 -25255
rect -6358 -25327 -6352 -25293
rect -6318 -25327 -6312 -25293
rect -6358 -25365 -6312 -25327
rect -6358 -25399 -6352 -25365
rect -6318 -25399 -6312 -25365
rect -6358 -25437 -6312 -25399
rect -6358 -25471 -6352 -25437
rect -6318 -25471 -6312 -25437
rect -6358 -25509 -6312 -25471
rect -6358 -25543 -6352 -25509
rect -6318 -25543 -6312 -25509
rect -6358 -25581 -6312 -25543
rect -6358 -25615 -6352 -25581
rect -6318 -25615 -6312 -25581
rect -6358 -25653 -6312 -25615
rect -6358 -25687 -6352 -25653
rect -6318 -25687 -6312 -25653
rect -6358 -25718 -6312 -25687
rect -5348 -25183 -5334 -25149
rect -5300 -25183 -5288 -25149
rect -4332 -25149 -4272 -24880
rect -4034 -25046 -3546 -25040
rect -4034 -25080 -3987 -25046
rect -3953 -25080 -3915 -25046
rect -3881 -25080 -3843 -25046
rect -3809 -25080 -3771 -25046
rect -3737 -25080 -3699 -25046
rect -3665 -25080 -3627 -25046
rect -3593 -25080 -3546 -25046
rect -4034 -25086 -3546 -25080
rect -4332 -25170 -4316 -25149
rect -5348 -25221 -5288 -25183
rect -5348 -25255 -5334 -25221
rect -5300 -25255 -5288 -25221
rect -5348 -25293 -5288 -25255
rect -5348 -25327 -5334 -25293
rect -5300 -25327 -5288 -25293
rect -5348 -25365 -5288 -25327
rect -5348 -25399 -5334 -25365
rect -5300 -25399 -5288 -25365
rect -5348 -25437 -5288 -25399
rect -5348 -25471 -5334 -25437
rect -5300 -25471 -5288 -25437
rect -5348 -25509 -5288 -25471
rect -5348 -25543 -5334 -25509
rect -5300 -25543 -5288 -25509
rect -5348 -25581 -5288 -25543
rect -5348 -25615 -5334 -25581
rect -5300 -25615 -5288 -25581
rect -5348 -25653 -5288 -25615
rect -4322 -25183 -4316 -25170
rect -4282 -25170 -4272 -25149
rect -3304 -25149 -3258 -25118
rect -4282 -25183 -4276 -25170
rect -4322 -25221 -4276 -25183
rect -4322 -25255 -4316 -25221
rect -4282 -25255 -4276 -25221
rect -4322 -25293 -4276 -25255
rect -4322 -25327 -4316 -25293
rect -4282 -25327 -4276 -25293
rect -4322 -25365 -4276 -25327
rect -4322 -25399 -4316 -25365
rect -4282 -25399 -4276 -25365
rect -4322 -25437 -4276 -25399
rect -4322 -25471 -4316 -25437
rect -4282 -25471 -4276 -25437
rect -4322 -25509 -4276 -25471
rect -4322 -25543 -4316 -25509
rect -4282 -25543 -4276 -25509
rect -4322 -25581 -4276 -25543
rect -4322 -25615 -4316 -25581
rect -4282 -25615 -4276 -25581
rect -4322 -25650 -4276 -25615
rect -3304 -25183 -3298 -25149
rect -3264 -25183 -3258 -25149
rect -3304 -25221 -3258 -25183
rect -3304 -25255 -3298 -25221
rect -3264 -25255 -3258 -25221
rect -3304 -25293 -3258 -25255
rect -3304 -25327 -3298 -25293
rect -3264 -25327 -3258 -25293
rect -3304 -25365 -3258 -25327
rect -3304 -25399 -3298 -25365
rect -3264 -25399 -3258 -25365
rect -3304 -25437 -3258 -25399
rect -3304 -25471 -3298 -25437
rect -3264 -25471 -3258 -25437
rect -3304 -25509 -3258 -25471
rect -3304 -25543 -3298 -25509
rect -3264 -25543 -3258 -25509
rect -3304 -25581 -3258 -25543
rect -3304 -25615 -3298 -25581
rect -3264 -25615 -3258 -25581
rect -5348 -25687 -5334 -25653
rect -5300 -25687 -5288 -25653
rect -7088 -25756 -6600 -25750
rect -7088 -25790 -7041 -25756
rect -7007 -25790 -6969 -25756
rect -6935 -25790 -6897 -25756
rect -6863 -25790 -6825 -25756
rect -6791 -25790 -6753 -25756
rect -6719 -25790 -6681 -25756
rect -6647 -25790 -6600 -25756
rect -7088 -25796 -6600 -25790
rect -6070 -25756 -5582 -25750
rect -6070 -25790 -6023 -25756
rect -5989 -25790 -5951 -25756
rect -5917 -25790 -5879 -25756
rect -5845 -25790 -5807 -25756
rect -5773 -25790 -5735 -25756
rect -5701 -25790 -5663 -25756
rect -5629 -25790 -5582 -25756
rect -6070 -25796 -5582 -25790
rect -6870 -25870 -6810 -25796
rect -5846 -25870 -5786 -25796
rect -6876 -25874 -6804 -25870
rect -6876 -25926 -6866 -25874
rect -6814 -25926 -6804 -25874
rect -6876 -25930 -6804 -25926
rect -5852 -25874 -5780 -25870
rect -5852 -25926 -5842 -25874
rect -5790 -25926 -5780 -25874
rect -5852 -25930 -5780 -25926
rect -5348 -26430 -5288 -25687
rect -4328 -25653 -4268 -25650
rect -4328 -25687 -4316 -25653
rect -4282 -25687 -4268 -25653
rect -3304 -25653 -3258 -25615
rect -3304 -25666 -3298 -25653
rect -5052 -25756 -4564 -25750
rect -5052 -25790 -5005 -25756
rect -4971 -25790 -4933 -25756
rect -4899 -25790 -4861 -25756
rect -4827 -25790 -4789 -25756
rect -4755 -25790 -4717 -25756
rect -4683 -25790 -4645 -25756
rect -4611 -25790 -4564 -25756
rect -5052 -25796 -4564 -25790
rect -4946 -25870 -4886 -25864
rect -4844 -25870 -4784 -25796
rect -4328 -25870 -4268 -25687
rect -3312 -25687 -3298 -25666
rect -3264 -25666 -3258 -25653
rect -3264 -25687 -3252 -25666
rect -4034 -25756 -3546 -25750
rect -4034 -25790 -3987 -25756
rect -3953 -25790 -3915 -25756
rect -3881 -25790 -3843 -25756
rect -3809 -25790 -3771 -25756
rect -3737 -25790 -3699 -25756
rect -3665 -25790 -3627 -25756
rect -3593 -25790 -3546 -25756
rect -4034 -25796 -3546 -25790
rect -3820 -25870 -3760 -25796
rect -3312 -25870 -3252 -25687
rect -2670 -25840 -2610 -23680
rect -2310 -23932 -2182 -23926
rect -2310 -23966 -2263 -23932
rect -2229 -23966 -2182 -23932
rect -2310 -23972 -2182 -23966
rect -2418 -24035 -2372 -24004
rect -2418 -24069 -2412 -24035
rect -2378 -24069 -2372 -24035
rect -2126 -24035 -2066 -23461
rect -1828 -23461 -1814 -23440
rect -1780 -23440 -1774 -23427
rect -1522 -23029 -1516 -22995
rect -1482 -23029 -1476 -22995
rect -1522 -23067 -1476 -23029
rect -1522 -23101 -1516 -23067
rect -1482 -23101 -1476 -23067
rect -1522 -23139 -1476 -23101
rect -1522 -23173 -1516 -23139
rect -1482 -23173 -1476 -23139
rect -1522 -23211 -1476 -23173
rect -1522 -23245 -1516 -23211
rect -1482 -23245 -1476 -23211
rect -1522 -23283 -1476 -23245
rect -1522 -23317 -1516 -23283
rect -1482 -23317 -1476 -23283
rect -1522 -23355 -1476 -23317
rect -1522 -23389 -1516 -23355
rect -1482 -23389 -1476 -23355
rect -1522 -23427 -1476 -23389
rect -1522 -23440 -1516 -23427
rect -1780 -23461 -1768 -23440
rect -1972 -23524 -1924 -23522
rect -2010 -23530 -1882 -23524
rect -2010 -23564 -1963 -23530
rect -1929 -23564 -1882 -23530
rect -2010 -23570 -1882 -23564
rect -1976 -23620 -1916 -23570
rect -1982 -23624 -1910 -23620
rect -1982 -23676 -1972 -23624
rect -1920 -23676 -1910 -23624
rect -1982 -23680 -1910 -23676
rect -1976 -23926 -1916 -23680
rect -2012 -23932 -1884 -23926
rect -2012 -23966 -1965 -23932
rect -1931 -23966 -1884 -23932
rect -2012 -23972 -1884 -23966
rect -2126 -24054 -2114 -24035
rect -2418 -24107 -2372 -24069
rect -2418 -24141 -2412 -24107
rect -2378 -24141 -2372 -24107
rect -2418 -24179 -2372 -24141
rect -2418 -24213 -2412 -24179
rect -2378 -24213 -2372 -24179
rect -2418 -24251 -2372 -24213
rect -2418 -24285 -2412 -24251
rect -2378 -24285 -2372 -24251
rect -2418 -24323 -2372 -24285
rect -2418 -24357 -2412 -24323
rect -2378 -24357 -2372 -24323
rect -2418 -24395 -2372 -24357
rect -2418 -24429 -2412 -24395
rect -2378 -24429 -2372 -24395
rect -2418 -24467 -2372 -24429
rect -2418 -24501 -2412 -24467
rect -2378 -24501 -2372 -24467
rect -2418 -24539 -2372 -24501
rect -2418 -24544 -2412 -24539
rect -2424 -24573 -2412 -24544
rect -2378 -24544 -2372 -24539
rect -2120 -24069 -2114 -24054
rect -2080 -24054 -2066 -24035
rect -1828 -24035 -1768 -23461
rect -1530 -23461 -1516 -23440
rect -1482 -23440 -1476 -23427
rect -1224 -22995 -1178 -22962
rect -1224 -23029 -1218 -22995
rect -1184 -23029 -1178 -22995
rect -1224 -23067 -1178 -23029
rect -1224 -23101 -1218 -23067
rect -1184 -23101 -1178 -23067
rect -1224 -23139 -1178 -23101
rect -1224 -23173 -1218 -23139
rect -1184 -23173 -1178 -23139
rect -1224 -23211 -1178 -23173
rect -1224 -23245 -1218 -23211
rect -1184 -23245 -1178 -23211
rect -1224 -23283 -1178 -23245
rect -1224 -23317 -1218 -23283
rect -1184 -23317 -1178 -23283
rect -1224 -23355 -1178 -23317
rect -1224 -23389 -1218 -23355
rect -1184 -23389 -1178 -23355
rect -1224 -23427 -1178 -23389
rect -1482 -23461 -1470 -23440
rect -1712 -23530 -1584 -23524
rect -1712 -23564 -1665 -23530
rect -1631 -23564 -1584 -23530
rect -1712 -23570 -1584 -23564
rect -1530 -23728 -1470 -23461
rect -1224 -23461 -1218 -23427
rect -1184 -23461 -1178 -23427
rect -1224 -23480 -1178 -23461
rect -926 -22995 -880 -22957
rect -926 -23029 -920 -22995
rect -886 -23029 -880 -22995
rect -926 -23067 -880 -23029
rect -926 -23101 -920 -23067
rect -886 -23101 -880 -23067
rect -926 -23139 -880 -23101
rect -926 -23173 -920 -23139
rect -886 -23173 -880 -23139
rect -926 -23211 -880 -23173
rect -926 -23245 -920 -23211
rect -886 -23245 -880 -23211
rect -926 -23283 -880 -23245
rect -926 -23317 -920 -23283
rect -886 -23317 -880 -23283
rect -926 -23355 -880 -23317
rect -926 -23389 -920 -23355
rect -886 -23389 -880 -23355
rect -926 -23427 -880 -23389
rect -628 -22957 -622 -22933
rect -588 -22932 -572 -22923
rect -330 -22923 -284 -22892
rect -588 -22933 -576 -22932
rect -588 -22957 -582 -22933
rect -628 -22995 -582 -22957
rect -628 -23029 -622 -22995
rect -588 -23029 -582 -22995
rect -628 -23067 -582 -23029
rect -628 -23101 -622 -23067
rect -588 -23101 -582 -23067
rect -628 -23139 -582 -23101
rect -628 -23173 -622 -23139
rect -588 -23173 -582 -23139
rect -628 -23211 -582 -23173
rect -628 -23245 -622 -23211
rect -588 -23245 -582 -23211
rect -628 -23283 -582 -23245
rect -628 -23317 -622 -23283
rect -588 -23317 -582 -23283
rect -628 -23355 -582 -23317
rect -628 -23389 -622 -23355
rect -588 -23389 -582 -23355
rect -628 -23396 -582 -23389
rect -330 -22957 -324 -22923
rect -290 -22957 -284 -22923
rect -38 -22923 22 -22538
rect 106 -22722 166 -22458
rect 252 -22618 324 -22614
rect 252 -22670 262 -22618
rect 314 -22670 324 -22618
rect 252 -22674 324 -22670
rect 100 -22726 172 -22722
rect 100 -22778 110 -22726
rect 162 -22778 172 -22726
rect 100 -22782 172 -22778
rect 76 -22820 204 -22814
rect 76 -22854 123 -22820
rect 157 -22854 204 -22820
rect 76 -22860 204 -22854
rect -38 -22924 -26 -22923
rect -330 -22995 -284 -22957
rect 8 -22924 22 -22923
rect 258 -22923 318 -22674
rect 410 -22722 470 -22458
rect 556 -22486 617 -22349
rect 854 -22349 868 -22328
rect 902 -22328 908 -22315
rect 902 -22349 914 -22328
rect 672 -22418 800 -22412
rect 672 -22452 719 -22418
rect 753 -22452 800 -22418
rect 672 -22458 800 -22452
rect 710 -22486 770 -22458
rect 854 -22486 914 -22349
rect 556 -22492 562 -22486
rect 558 -22538 562 -22492
rect 614 -22538 914 -22486
rect 558 -22546 914 -22538
rect 558 -22698 618 -22546
rect 404 -22726 476 -22722
rect 404 -22778 414 -22726
rect 466 -22778 476 -22726
rect 404 -22782 476 -22778
rect 558 -22758 916 -22698
rect 374 -22820 502 -22814
rect 374 -22854 421 -22820
rect 455 -22854 502 -22820
rect 374 -22860 502 -22854
rect 258 -22954 272 -22923
rect -26 -22974 8 -22957
rect 266 -22957 272 -22954
rect 306 -22954 318 -22923
rect 558 -22923 618 -22758
rect 706 -22814 766 -22758
rect 672 -22820 800 -22814
rect 672 -22854 719 -22820
rect 753 -22854 800 -22820
rect 672 -22860 800 -22854
rect 558 -22936 570 -22923
rect 306 -22957 312 -22954
rect -330 -23029 -324 -22995
rect -290 -23029 -284 -22995
rect -330 -23067 -284 -23029
rect -330 -23101 -324 -23067
rect -290 -23101 -284 -23067
rect -330 -23139 -284 -23101
rect -330 -23173 -324 -23139
rect -290 -23173 -284 -23139
rect -330 -23211 -284 -23173
rect -330 -23245 -324 -23211
rect -290 -23245 -284 -23211
rect -330 -23283 -284 -23245
rect -330 -23317 -324 -23283
rect -290 -23317 -284 -23283
rect -330 -23355 -284 -23317
rect -330 -23389 -324 -23355
rect -290 -23389 -284 -23355
rect -926 -23461 -920 -23427
rect -886 -23461 -880 -23427
rect -1414 -23530 -1286 -23524
rect -1414 -23564 -1367 -23530
rect -1333 -23564 -1286 -23530
rect -1414 -23570 -1286 -23564
rect -1536 -23732 -1464 -23728
rect -1536 -23784 -1526 -23732
rect -1474 -23784 -1464 -23732
rect -1536 -23788 -1464 -23784
rect -1714 -23932 -1586 -23926
rect -1714 -23966 -1667 -23932
rect -1633 -23966 -1586 -23932
rect -1714 -23972 -1586 -23966
rect -1828 -24054 -1816 -24035
rect -2080 -24069 -2074 -24054
rect -2120 -24107 -2074 -24069
rect -2120 -24141 -2114 -24107
rect -2080 -24141 -2074 -24107
rect -2120 -24179 -2074 -24141
rect -2120 -24213 -2114 -24179
rect -2080 -24213 -2074 -24179
rect -2120 -24251 -2074 -24213
rect -2120 -24285 -2114 -24251
rect -2080 -24285 -2074 -24251
rect -2120 -24323 -2074 -24285
rect -2120 -24357 -2114 -24323
rect -2080 -24357 -2074 -24323
rect -2120 -24395 -2074 -24357
rect -2120 -24429 -2114 -24395
rect -2080 -24429 -2074 -24395
rect -2120 -24467 -2074 -24429
rect -2120 -24501 -2114 -24467
rect -2080 -24501 -2074 -24467
rect -2120 -24539 -2074 -24501
rect -1822 -24069 -1816 -24054
rect -1782 -24054 -1768 -24035
rect -1530 -24035 -1470 -23788
rect -1416 -23932 -1288 -23926
rect -1416 -23966 -1369 -23932
rect -1335 -23966 -1288 -23932
rect -1416 -23972 -1288 -23966
rect -1230 -24016 -1170 -23480
rect -926 -23492 -880 -23461
rect -622 -23427 -588 -23396
rect -330 -23424 -284 -23389
rect -32 -22995 14 -22974
rect -32 -23029 -26 -22995
rect 8 -23029 14 -22995
rect -32 -23067 14 -23029
rect -32 -23101 -26 -23067
rect 8 -23101 14 -23067
rect -32 -23139 14 -23101
rect -32 -23173 -26 -23139
rect 8 -23173 14 -23139
rect -32 -23211 14 -23173
rect -32 -23245 -26 -23211
rect 8 -23245 14 -23211
rect -32 -23283 14 -23245
rect -32 -23317 -26 -23283
rect 8 -23317 14 -23283
rect -32 -23355 14 -23317
rect -32 -23389 -26 -23355
rect 8 -23389 14 -23355
rect -32 -23416 14 -23389
rect 266 -22995 312 -22957
rect 266 -23029 272 -22995
rect 306 -23029 312 -22995
rect 266 -23067 312 -23029
rect 266 -23101 272 -23067
rect 306 -23101 312 -23067
rect 266 -23139 312 -23101
rect 266 -23173 272 -23139
rect 306 -23173 312 -23139
rect 266 -23211 312 -23173
rect 266 -23245 272 -23211
rect 306 -23245 312 -23211
rect 266 -23283 312 -23245
rect 266 -23317 272 -23283
rect 306 -23317 312 -23283
rect 266 -23355 312 -23317
rect 266 -23389 272 -23355
rect 306 -23389 312 -23355
rect -336 -23427 -276 -23424
rect -336 -23438 -324 -23427
rect -622 -23474 -588 -23461
rect -338 -23461 -324 -23438
rect -290 -23461 -276 -23427
rect -1116 -23530 -988 -23524
rect -1116 -23564 -1069 -23530
rect -1035 -23564 -988 -23530
rect -1116 -23570 -988 -23564
rect -818 -23530 -690 -23524
rect -818 -23564 -771 -23530
rect -737 -23564 -690 -23530
rect -818 -23570 -690 -23564
rect -1080 -23620 -1020 -23570
rect -786 -23620 -726 -23570
rect -1086 -23624 -1014 -23620
rect -1086 -23676 -1076 -23624
rect -1024 -23676 -1014 -23624
rect -1086 -23680 -1014 -23676
rect -792 -23624 -720 -23620
rect -792 -23676 -782 -23624
rect -730 -23676 -720 -23624
rect -792 -23680 -720 -23676
rect -1076 -23926 -1020 -23680
rect -786 -23926 -730 -23680
rect -1118 -23932 -990 -23926
rect -1118 -23966 -1071 -23932
rect -1037 -23966 -990 -23932
rect -1118 -23972 -990 -23966
rect -820 -23932 -692 -23926
rect -820 -23966 -773 -23932
rect -739 -23966 -692 -23932
rect -820 -23972 -692 -23966
rect -1530 -24054 -1518 -24035
rect -1782 -24069 -1776 -24054
rect -1822 -24107 -1776 -24069
rect -1822 -24141 -1816 -24107
rect -1782 -24141 -1776 -24107
rect -1822 -24179 -1776 -24141
rect -1822 -24213 -1816 -24179
rect -1782 -24213 -1776 -24179
rect -1822 -24251 -1776 -24213
rect -1822 -24285 -1816 -24251
rect -1782 -24285 -1776 -24251
rect -1822 -24323 -1776 -24285
rect -1822 -24357 -1816 -24323
rect -1782 -24357 -1776 -24323
rect -1822 -24395 -1776 -24357
rect -1822 -24429 -1816 -24395
rect -1782 -24429 -1776 -24395
rect -1822 -24467 -1776 -24429
rect -1822 -24501 -1816 -24467
rect -1782 -24501 -1776 -24467
rect -1822 -24534 -1776 -24501
rect -1524 -24069 -1518 -24054
rect -1484 -24054 -1470 -24035
rect -1220 -24035 -1186 -24016
rect -1484 -24069 -1478 -24054
rect -1524 -24107 -1478 -24069
rect -1524 -24141 -1518 -24107
rect -1484 -24141 -1478 -24107
rect -1524 -24179 -1478 -24141
rect -1524 -24213 -1518 -24179
rect -1484 -24213 -1478 -24179
rect -1524 -24251 -1478 -24213
rect -1524 -24285 -1518 -24251
rect -1484 -24285 -1478 -24251
rect -1524 -24323 -1478 -24285
rect -1524 -24357 -1518 -24323
rect -1484 -24357 -1478 -24323
rect -1524 -24395 -1478 -24357
rect -1524 -24429 -1518 -24395
rect -1484 -24429 -1478 -24395
rect -1524 -24467 -1478 -24429
rect -1524 -24501 -1518 -24467
rect -1484 -24501 -1478 -24467
rect -1524 -24534 -1478 -24501
rect -1226 -24069 -1220 -24056
rect -928 -24035 -882 -24004
rect -636 -24010 -576 -23474
rect -338 -23480 -276 -23461
rect -26 -23427 8 -23416
rect -26 -23480 8 -23461
rect 266 -23427 312 -23389
rect 564 -22957 570 -22936
rect 604 -22936 618 -22923
rect 856 -22923 916 -22758
rect 604 -22957 610 -22936
rect 856 -22940 868 -22923
rect 564 -22995 610 -22957
rect 564 -23029 570 -22995
rect 604 -23029 610 -22995
rect 564 -23067 610 -23029
rect 564 -23101 570 -23067
rect 604 -23101 610 -23067
rect 564 -23139 610 -23101
rect 564 -23173 570 -23139
rect 604 -23173 610 -23139
rect 564 -23211 610 -23173
rect 564 -23245 570 -23211
rect 604 -23245 610 -23211
rect 564 -23283 610 -23245
rect 564 -23317 570 -23283
rect 604 -23317 610 -23283
rect 564 -23355 610 -23317
rect 564 -23389 570 -23355
rect 604 -23389 610 -23355
rect 564 -23402 610 -23389
rect 862 -22957 868 -22940
rect 902 -22940 916 -22923
rect 902 -22957 908 -22940
rect 862 -22995 908 -22957
rect 862 -23029 868 -22995
rect 902 -23029 908 -22995
rect 862 -23067 908 -23029
rect 862 -23101 868 -23067
rect 902 -23101 908 -23067
rect 862 -23139 908 -23101
rect 862 -23173 868 -23139
rect 902 -23173 908 -23139
rect 862 -23211 908 -23173
rect 862 -23245 868 -23211
rect 902 -23245 908 -23211
rect 862 -23283 908 -23245
rect 862 -23317 868 -23283
rect 902 -23317 908 -23283
rect 862 -23355 908 -23317
rect 862 -23389 868 -23355
rect 902 -23389 908 -23355
rect 266 -23461 272 -23427
rect 306 -23461 312 -23427
rect 570 -23427 604 -23402
rect -512 -23530 -392 -23524
rect -512 -23564 -473 -23530
rect -439 -23564 -392 -23530
rect -512 -23570 -392 -23564
rect -336 -23728 -276 -23480
rect -222 -23530 -96 -23524
rect -222 -23564 -175 -23530
rect -141 -23564 -96 -23530
rect -222 -23570 -96 -23564
rect -342 -23732 -270 -23728
rect -342 -23784 -332 -23732
rect -280 -23784 -270 -23732
rect -342 -23788 -270 -23784
rect -522 -23932 -394 -23926
rect -522 -23966 -475 -23932
rect -441 -23966 -394 -23932
rect -522 -23972 -394 -23966
rect -336 -24016 -276 -23788
rect -224 -23932 -96 -23926
rect -224 -23966 -177 -23932
rect -143 -23966 -96 -23932
rect -224 -23972 -96 -23966
rect -1186 -24069 -1180 -24056
rect -1226 -24107 -1180 -24069
rect -1226 -24141 -1220 -24107
rect -1186 -24141 -1180 -24107
rect -1226 -24179 -1180 -24141
rect -1226 -24213 -1220 -24179
rect -1186 -24213 -1180 -24179
rect -1226 -24251 -1180 -24213
rect -1226 -24285 -1220 -24251
rect -1186 -24285 -1180 -24251
rect -1226 -24323 -1180 -24285
rect -1226 -24357 -1220 -24323
rect -1186 -24357 -1180 -24323
rect -1226 -24395 -1180 -24357
rect -1226 -24429 -1220 -24395
rect -1186 -24429 -1180 -24395
rect -1226 -24467 -1180 -24429
rect -1226 -24501 -1220 -24467
rect -1186 -24501 -1180 -24467
rect -1226 -24532 -1180 -24501
rect -928 -24069 -922 -24035
rect -888 -24069 -882 -24035
rect -624 -24035 -590 -24016
rect -928 -24107 -882 -24069
rect -928 -24141 -922 -24107
rect -888 -24141 -882 -24107
rect -928 -24179 -882 -24141
rect -928 -24213 -922 -24179
rect -888 -24213 -882 -24179
rect -928 -24251 -882 -24213
rect -928 -24285 -922 -24251
rect -888 -24285 -882 -24251
rect -928 -24323 -882 -24285
rect -928 -24357 -922 -24323
rect -888 -24357 -882 -24323
rect -928 -24395 -882 -24357
rect -928 -24429 -922 -24395
rect -888 -24429 -882 -24395
rect -928 -24467 -882 -24429
rect -928 -24501 -922 -24467
rect -888 -24501 -882 -24467
rect -1816 -24538 -1782 -24534
rect -2378 -24573 -2364 -24544
rect -2120 -24546 -2114 -24539
rect -2424 -24740 -2364 -24573
rect -2128 -24573 -2114 -24546
rect -2080 -24542 -2074 -24539
rect -1828 -24539 -1768 -24538
rect -2080 -24573 -2060 -24542
rect -2128 -24592 -2060 -24573
rect -1828 -24573 -1816 -24539
rect -1782 -24573 -1768 -24539
rect -2310 -24642 -2182 -24636
rect -2310 -24676 -2263 -24642
rect -2229 -24676 -2182 -24642
rect -2310 -24682 -2182 -24676
rect -2278 -24740 -2218 -24682
rect -2128 -24740 -2068 -24592
rect -2012 -24642 -1884 -24636
rect -2012 -24676 -1965 -24642
rect -1931 -24676 -1884 -24642
rect -2012 -24682 -1884 -24676
rect -1828 -24712 -1768 -24573
rect -1518 -24539 -1484 -24534
rect -1518 -24592 -1484 -24573
rect -1234 -24539 -1174 -24532
rect -1234 -24573 -1220 -24539
rect -1186 -24573 -1174 -24539
rect -928 -24539 -882 -24501
rect -928 -24544 -922 -24539
rect -1714 -24642 -1586 -24636
rect -1714 -24676 -1667 -24642
rect -1633 -24676 -1586 -24642
rect -1714 -24682 -1586 -24676
rect -1416 -24642 -1288 -24636
rect -1416 -24676 -1369 -24642
rect -1335 -24676 -1288 -24642
rect -1416 -24682 -1288 -24676
rect -2424 -24800 -2068 -24740
rect -1834 -24716 -1762 -24712
rect -1834 -24768 -1824 -24716
rect -1772 -24768 -1762 -24716
rect -1834 -24772 -1762 -24768
rect -2426 -24810 -2364 -24800
rect -2426 -24862 -2422 -24810
rect -2370 -24860 -2364 -24810
rect -2370 -24862 -2366 -24860
rect -2426 -24872 -2366 -24862
rect -1984 -24918 -1912 -24914
rect -1984 -24970 -1974 -24918
rect -1922 -24970 -1912 -24918
rect -1984 -24974 -1912 -24970
rect -1978 -25036 -1918 -24974
rect -2310 -25042 -2182 -25036
rect -2310 -25076 -2263 -25042
rect -2229 -25076 -2182 -25042
rect -2310 -25082 -2182 -25076
rect -2012 -25042 -1884 -25036
rect -2012 -25076 -1965 -25042
rect -1931 -25076 -1884 -25042
rect -2012 -25082 -1884 -25076
rect -2418 -25145 -2372 -25114
rect -2418 -25179 -2412 -25145
rect -2378 -25179 -2372 -25145
rect -2418 -25217 -2372 -25179
rect -2418 -25251 -2412 -25217
rect -2378 -25251 -2372 -25217
rect -2418 -25289 -2372 -25251
rect -2418 -25323 -2412 -25289
rect -2378 -25323 -2372 -25289
rect -2418 -25361 -2372 -25323
rect -2418 -25395 -2412 -25361
rect -2378 -25395 -2372 -25361
rect -2418 -25433 -2372 -25395
rect -2418 -25467 -2412 -25433
rect -2378 -25467 -2372 -25433
rect -2418 -25505 -2372 -25467
rect -2418 -25539 -2412 -25505
rect -2378 -25539 -2372 -25505
rect -2418 -25577 -2372 -25539
rect -2418 -25611 -2412 -25577
rect -2378 -25611 -2372 -25577
rect -2418 -25649 -2372 -25611
rect -2418 -25650 -2412 -25649
rect -2426 -25683 -2412 -25650
rect -2378 -25650 -2372 -25649
rect -2120 -25145 -2074 -25114
rect -2120 -25179 -2114 -25145
rect -2080 -25179 -2074 -25145
rect -1828 -25145 -1768 -24772
rect -1680 -24914 -1620 -24682
rect -1540 -24810 -1468 -24806
rect -1540 -24862 -1530 -24810
rect -1478 -24862 -1468 -24810
rect -1540 -24866 -1468 -24862
rect -1686 -24918 -1614 -24914
rect -1686 -24970 -1676 -24918
rect -1624 -24970 -1614 -24918
rect -1686 -24974 -1614 -24970
rect -1714 -25042 -1586 -25036
rect -1714 -25076 -1667 -25042
rect -1633 -25076 -1586 -25042
rect -1714 -25082 -1586 -25076
rect -1828 -25170 -1816 -25145
rect -2120 -25217 -2074 -25179
rect -2120 -25251 -2114 -25217
rect -2080 -25251 -2074 -25217
rect -2120 -25289 -2074 -25251
rect -2120 -25323 -2114 -25289
rect -2080 -25323 -2074 -25289
rect -2120 -25361 -2074 -25323
rect -2120 -25395 -2114 -25361
rect -2080 -25395 -2074 -25361
rect -2120 -25433 -2074 -25395
rect -2120 -25467 -2114 -25433
rect -2080 -25467 -2074 -25433
rect -2120 -25505 -2074 -25467
rect -2120 -25539 -2114 -25505
rect -2080 -25539 -2074 -25505
rect -2120 -25577 -2074 -25539
rect -2120 -25611 -2114 -25577
rect -2080 -25611 -2074 -25577
rect -2120 -25649 -2074 -25611
rect -2378 -25683 -2366 -25650
rect -2120 -25654 -2114 -25649
rect -2426 -25840 -2366 -25683
rect -2126 -25683 -2114 -25654
rect -2080 -25654 -2074 -25649
rect -1822 -25179 -1816 -25170
rect -1782 -25170 -1768 -25145
rect -1534 -25126 -1474 -24866
rect -1384 -24914 -1324 -24682
rect -1234 -24712 -1174 -24573
rect -936 -24573 -922 -24544
rect -888 -24544 -882 -24539
rect -630 -24069 -624 -24044
rect -338 -24035 -276 -24016
rect -590 -24069 -584 -24044
rect -338 -24054 -326 -24035
rect -630 -24107 -584 -24069
rect -630 -24141 -624 -24107
rect -590 -24141 -584 -24107
rect -630 -24179 -584 -24141
rect -630 -24213 -624 -24179
rect -590 -24213 -584 -24179
rect -630 -24251 -584 -24213
rect -630 -24285 -624 -24251
rect -590 -24285 -584 -24251
rect -630 -24323 -584 -24285
rect -630 -24357 -624 -24323
rect -590 -24357 -584 -24323
rect -630 -24395 -584 -24357
rect -630 -24429 -624 -24395
rect -590 -24429 -584 -24395
rect -630 -24467 -584 -24429
rect -630 -24501 -624 -24467
rect -590 -24501 -584 -24467
rect -630 -24539 -584 -24501
rect -888 -24550 -876 -24544
rect -888 -24573 -870 -24550
rect -630 -24562 -624 -24539
rect -936 -24592 -870 -24573
rect -634 -24573 -624 -24562
rect -590 -24562 -584 -24539
rect -332 -24069 -326 -24054
rect -292 -24054 -276 -24035
rect -42 -24035 18 -23480
rect 266 -23492 312 -23461
rect 554 -23461 570 -23436
rect 862 -23427 908 -23389
rect 604 -23461 614 -23436
rect 862 -23440 868 -23427
rect 76 -23530 204 -23524
rect 76 -23564 123 -23530
rect 157 -23564 204 -23530
rect 76 -23570 204 -23564
rect 374 -23530 502 -23524
rect 374 -23564 421 -23530
rect 455 -23564 502 -23530
rect 374 -23570 502 -23564
rect 108 -23620 168 -23570
rect 410 -23620 470 -23570
rect 102 -23624 174 -23620
rect 102 -23676 112 -23624
rect 164 -23676 174 -23624
rect 102 -23680 174 -23676
rect 404 -23624 476 -23620
rect 404 -23676 414 -23624
rect 466 -23676 476 -23624
rect 404 -23680 476 -23676
rect 112 -23926 168 -23680
rect 414 -23926 470 -23680
rect 74 -23932 202 -23926
rect 74 -23966 121 -23932
rect 155 -23966 202 -23932
rect 74 -23972 202 -23966
rect 372 -23932 500 -23926
rect 372 -23966 419 -23932
rect 453 -23966 500 -23932
rect 372 -23972 500 -23966
rect -42 -24044 -28 -24035
rect -292 -24069 -286 -24054
rect -332 -24107 -286 -24069
rect -332 -24141 -326 -24107
rect -292 -24141 -286 -24107
rect -332 -24179 -286 -24141
rect -332 -24213 -326 -24179
rect -292 -24213 -286 -24179
rect -332 -24251 -286 -24213
rect -332 -24285 -326 -24251
rect -292 -24285 -286 -24251
rect -332 -24323 -286 -24285
rect -332 -24357 -326 -24323
rect -292 -24357 -286 -24323
rect -332 -24395 -286 -24357
rect -332 -24429 -326 -24395
rect -292 -24429 -286 -24395
rect -332 -24467 -286 -24429
rect -332 -24501 -326 -24467
rect -292 -24501 -286 -24467
rect -332 -24539 -286 -24501
rect -34 -24069 -28 -24044
rect 6 -24044 18 -24035
rect 264 -24035 310 -24004
rect 6 -24069 12 -24044
rect -34 -24107 12 -24069
rect -34 -24141 -28 -24107
rect 6 -24141 12 -24107
rect -34 -24179 12 -24141
rect -34 -24213 -28 -24179
rect 6 -24213 12 -24179
rect -34 -24251 12 -24213
rect -34 -24285 -28 -24251
rect 6 -24285 12 -24251
rect -34 -24323 12 -24285
rect -34 -24357 -28 -24323
rect 6 -24357 12 -24323
rect -34 -24395 12 -24357
rect -34 -24429 -28 -24395
rect 6 -24429 12 -24395
rect -34 -24467 12 -24429
rect -34 -24501 -28 -24467
rect 6 -24501 12 -24467
rect -34 -24502 12 -24501
rect 264 -24069 270 -24035
rect 304 -24069 310 -24035
rect 264 -24107 310 -24069
rect 264 -24141 270 -24107
rect 304 -24141 310 -24107
rect 264 -24179 310 -24141
rect 264 -24213 270 -24179
rect 304 -24213 310 -24179
rect 264 -24251 310 -24213
rect 264 -24285 270 -24251
rect 304 -24285 310 -24251
rect 264 -24323 310 -24285
rect 264 -24357 270 -24323
rect 304 -24357 310 -24323
rect 264 -24395 310 -24357
rect 264 -24429 270 -24395
rect 304 -24429 310 -24395
rect 264 -24467 310 -24429
rect 264 -24501 270 -24467
rect 304 -24501 310 -24467
rect -28 -24538 6 -24502
rect -590 -24573 -574 -24562
rect -1118 -24642 -990 -24636
rect -1118 -24676 -1071 -24642
rect -1037 -24676 -990 -24642
rect -1118 -24682 -990 -24676
rect -1240 -24716 -1168 -24712
rect -1240 -24768 -1230 -24716
rect -1178 -24768 -1168 -24716
rect -1240 -24772 -1168 -24768
rect -1390 -24918 -1318 -24914
rect -1390 -24970 -1380 -24918
rect -1328 -24970 -1318 -24918
rect -1390 -24974 -1318 -24970
rect -1416 -25042 -1288 -25036
rect -1416 -25076 -1369 -25042
rect -1335 -25076 -1288 -25042
rect -1416 -25082 -1288 -25076
rect -1534 -25145 -1466 -25126
rect -1534 -25160 -1518 -25145
rect -1782 -25179 -1776 -25170
rect -1822 -25217 -1776 -25179
rect -1526 -25179 -1518 -25160
rect -1484 -25179 -1466 -25145
rect -1234 -25145 -1174 -24772
rect -936 -24806 -876 -24592
rect -820 -24642 -692 -24636
rect -820 -24676 -773 -24642
rect -739 -24676 -692 -24642
rect -820 -24682 -692 -24676
rect -634 -24712 -574 -24573
rect -332 -24573 -326 -24539
rect -292 -24573 -286 -24539
rect -332 -24604 -286 -24573
rect -40 -24539 20 -24538
rect -40 -24573 -28 -24539
rect 6 -24573 20 -24539
rect 264 -24539 310 -24501
rect 264 -24542 270 -24539
rect -522 -24642 -394 -24636
rect -522 -24676 -475 -24642
rect -441 -24676 -394 -24642
rect -522 -24682 -394 -24676
rect -224 -24642 -96 -24636
rect -224 -24676 -177 -24642
rect -143 -24676 -96 -24642
rect -224 -24682 -96 -24676
rect -640 -24716 -568 -24712
rect -640 -24768 -630 -24716
rect -578 -24768 -568 -24716
rect -640 -24772 -568 -24768
rect -942 -24810 -870 -24806
rect -942 -24862 -932 -24810
rect -880 -24862 -870 -24810
rect -942 -24866 -870 -24862
rect -1086 -24918 -1014 -24914
rect -1086 -24970 -1076 -24918
rect -1024 -24970 -1014 -24918
rect -1086 -24974 -1014 -24970
rect -790 -24918 -718 -24914
rect -790 -24970 -780 -24918
rect -728 -24970 -718 -24918
rect -790 -24974 -718 -24970
rect -1080 -25042 -1020 -24974
rect -784 -25042 -724 -24974
rect -1106 -25076 -1071 -25042
rect -1037 -25076 -1002 -25042
rect -808 -25076 -773 -25042
rect -739 -25076 -704 -25042
rect -1234 -25160 -1220 -25145
rect -1526 -25184 -1466 -25179
rect -1226 -25179 -1220 -25170
rect -1186 -25160 -1174 -25145
rect -922 -25145 -888 -25126
rect -1186 -25179 -1180 -25170
rect -1822 -25251 -1816 -25217
rect -1782 -25251 -1776 -25217
rect -1822 -25289 -1776 -25251
rect -1822 -25323 -1816 -25289
rect -1782 -25323 -1776 -25289
rect -1822 -25361 -1776 -25323
rect -1822 -25395 -1816 -25361
rect -1782 -25395 -1776 -25361
rect -1822 -25433 -1776 -25395
rect -1822 -25467 -1816 -25433
rect -1782 -25467 -1776 -25433
rect -1822 -25505 -1776 -25467
rect -1822 -25539 -1816 -25505
rect -1782 -25539 -1776 -25505
rect -1822 -25577 -1776 -25539
rect -1822 -25611 -1816 -25577
rect -1782 -25611 -1776 -25577
rect -1822 -25649 -1776 -25611
rect -1822 -25654 -1816 -25649
rect -2080 -25683 -2066 -25654
rect -2310 -25752 -2182 -25746
rect -2310 -25786 -2263 -25752
rect -2229 -25786 -2182 -25752
rect -2310 -25792 -2218 -25786
rect -2216 -25792 -2182 -25786
rect -2278 -25840 -2218 -25792
rect -2126 -25840 -2066 -25683
rect -1782 -25654 -1776 -25649
rect -1524 -25217 -1478 -25184
rect -1524 -25251 -1518 -25217
rect -1484 -25251 -1478 -25217
rect -1524 -25289 -1478 -25251
rect -1524 -25323 -1518 -25289
rect -1484 -25323 -1478 -25289
rect -1524 -25361 -1478 -25323
rect -1524 -25395 -1518 -25361
rect -1484 -25395 -1478 -25361
rect -1524 -25433 -1478 -25395
rect -1524 -25467 -1518 -25433
rect -1484 -25467 -1478 -25433
rect -1524 -25505 -1478 -25467
rect -1524 -25539 -1518 -25505
rect -1484 -25539 -1478 -25505
rect -1524 -25577 -1478 -25539
rect -1524 -25611 -1518 -25577
rect -1484 -25611 -1478 -25577
rect -1524 -25649 -1478 -25611
rect -1524 -25654 -1518 -25649
rect -1816 -25702 -1782 -25683
rect -1484 -25654 -1478 -25649
rect -1226 -25217 -1180 -25179
rect -1226 -25251 -1220 -25217
rect -1186 -25251 -1180 -25217
rect -1226 -25289 -1180 -25251
rect -1226 -25323 -1220 -25289
rect -1186 -25323 -1180 -25289
rect -1226 -25361 -1180 -25323
rect -1226 -25395 -1220 -25361
rect -1186 -25395 -1180 -25361
rect -1226 -25433 -1180 -25395
rect -1226 -25467 -1220 -25433
rect -1186 -25467 -1180 -25433
rect -1226 -25505 -1180 -25467
rect -1226 -25539 -1220 -25505
rect -1186 -25539 -1180 -25505
rect -1226 -25577 -1180 -25539
rect -1226 -25611 -1220 -25577
rect -1186 -25611 -1180 -25577
rect -1226 -25649 -1180 -25611
rect -1226 -25654 -1220 -25649
rect -1518 -25702 -1484 -25683
rect -1186 -25654 -1180 -25649
rect -928 -25179 -922 -25170
rect -634 -25145 -574 -24772
rect -486 -24914 -426 -24682
rect -344 -24810 -272 -24806
rect -344 -24862 -334 -24810
rect -282 -24862 -272 -24810
rect -344 -24866 -272 -24862
rect -492 -24918 -420 -24914
rect -492 -24970 -482 -24918
rect -430 -24970 -420 -24918
rect -492 -24974 -420 -24970
rect -522 -25042 -394 -25036
rect -522 -25076 -475 -25042
rect -441 -25076 -394 -25042
rect -522 -25082 -394 -25076
rect -634 -25158 -624 -25145
rect -888 -25179 -882 -25170
rect -928 -25217 -882 -25179
rect -928 -25251 -922 -25217
rect -888 -25251 -882 -25217
rect -928 -25289 -882 -25251
rect -928 -25323 -922 -25289
rect -888 -25323 -882 -25289
rect -928 -25361 -882 -25323
rect -928 -25395 -922 -25361
rect -888 -25395 -882 -25361
rect -928 -25433 -882 -25395
rect -928 -25467 -922 -25433
rect -888 -25467 -882 -25433
rect -928 -25505 -882 -25467
rect -928 -25539 -922 -25505
rect -888 -25539 -882 -25505
rect -928 -25577 -882 -25539
rect -928 -25611 -922 -25577
rect -888 -25611 -882 -25577
rect -928 -25649 -882 -25611
rect -630 -25179 -624 -25170
rect -590 -25158 -574 -25145
rect -338 -25126 -278 -24866
rect -190 -24914 -130 -24682
rect -40 -24712 20 -24573
rect 262 -24573 270 -24542
rect 304 -24542 310 -24539
rect 554 -24016 614 -23461
rect 856 -23461 868 -23440
rect 902 -23440 908 -23427
rect 902 -23461 916 -23440
rect 856 -23480 916 -23461
rect 672 -23530 800 -23524
rect 672 -23564 719 -23530
rect 753 -23564 800 -23530
rect 672 -23570 708 -23564
rect 768 -23570 800 -23564
rect 952 -23732 1012 -21540
rect 952 -23784 956 -23732
rect 1008 -23784 1012 -23732
rect 670 -23932 798 -23926
rect 670 -23966 717 -23932
rect 751 -23966 798 -23932
rect 670 -23972 798 -23966
rect 554 -24035 618 -24016
rect 554 -24069 568 -24035
rect 602 -24052 618 -24035
rect 852 -24035 912 -24016
rect 852 -24048 866 -24035
rect 602 -24069 614 -24052
rect 554 -24107 614 -24069
rect 554 -24141 568 -24107
rect 602 -24141 614 -24107
rect 554 -24179 614 -24141
rect 554 -24213 568 -24179
rect 602 -24213 614 -24179
rect 554 -24251 614 -24213
rect 554 -24285 568 -24251
rect 602 -24285 614 -24251
rect 554 -24323 614 -24285
rect 554 -24357 568 -24323
rect 602 -24357 614 -24323
rect 554 -24395 614 -24357
rect 554 -24429 568 -24395
rect 602 -24429 614 -24395
rect 554 -24467 614 -24429
rect 554 -24501 568 -24467
rect 602 -24501 614 -24467
rect 554 -24539 614 -24501
rect 304 -24573 322 -24542
rect 74 -24642 202 -24636
rect 74 -24676 121 -24642
rect 155 -24676 202 -24642
rect 74 -24682 202 -24676
rect -46 -24716 26 -24712
rect -46 -24768 -36 -24716
rect 16 -24768 26 -24716
rect -46 -24772 26 -24768
rect -196 -24918 -124 -24914
rect -196 -24970 -186 -24918
rect -134 -24970 -124 -24918
rect -196 -24974 -124 -24970
rect -224 -25042 -96 -25036
rect -224 -25076 -177 -25042
rect -143 -25076 -96 -25042
rect -224 -25082 -96 -25076
rect -338 -25145 -274 -25126
rect -338 -25164 -326 -25145
rect -590 -25179 -584 -25170
rect -630 -25217 -584 -25179
rect -334 -25179 -326 -25164
rect -292 -25179 -274 -25145
rect -40 -25145 20 -24772
rect 262 -24806 322 -24573
rect 554 -24573 568 -24539
rect 602 -24573 614 -24539
rect 860 -24069 866 -24048
rect 900 -24048 912 -24035
rect 900 -24069 906 -24048
rect 860 -24107 906 -24069
rect 860 -24141 866 -24107
rect 900 -24141 906 -24107
rect 860 -24179 906 -24141
rect 860 -24213 866 -24179
rect 900 -24213 906 -24179
rect 860 -24251 906 -24213
rect 860 -24285 866 -24251
rect 900 -24285 906 -24251
rect 860 -24323 906 -24285
rect 860 -24357 866 -24323
rect 900 -24357 906 -24323
rect 860 -24395 906 -24357
rect 860 -24429 866 -24395
rect 900 -24429 906 -24395
rect 860 -24467 906 -24429
rect 860 -24501 866 -24467
rect 900 -24501 906 -24467
rect 860 -24539 906 -24501
rect 860 -24540 866 -24539
rect 852 -24562 866 -24540
rect 372 -24642 500 -24636
rect 372 -24676 419 -24642
rect 453 -24676 500 -24642
rect 372 -24682 500 -24676
rect 554 -24712 614 -24573
rect 850 -24573 866 -24562
rect 900 -24540 906 -24539
rect 900 -24573 912 -24540
rect 850 -24592 912 -24573
rect 670 -24642 798 -24636
rect 670 -24676 717 -24642
rect 751 -24676 798 -24642
rect 670 -24682 762 -24676
rect 764 -24682 798 -24676
rect 548 -24716 620 -24712
rect 702 -24716 762 -24682
rect 852 -24716 912 -24592
rect 548 -24768 558 -24716
rect 610 -24768 912 -24716
rect 548 -24772 912 -24768
rect 554 -24776 912 -24772
rect 256 -24810 328 -24806
rect 256 -24862 266 -24810
rect 318 -24862 328 -24810
rect 256 -24866 328 -24862
rect 100 -24918 172 -24914
rect 100 -24970 110 -24918
rect 162 -24970 172 -24918
rect 100 -24974 172 -24970
rect 404 -24918 476 -24914
rect 404 -24970 414 -24918
rect 466 -24970 476 -24918
rect 404 -24974 476 -24970
rect 554 -24938 614 -24776
rect 106 -25036 166 -24974
rect 410 -25036 470 -24974
rect 554 -24998 914 -24938
rect 74 -25042 202 -25036
rect 74 -25076 121 -25042
rect 155 -25076 202 -25042
rect 74 -25082 202 -25076
rect 372 -25042 500 -25036
rect 372 -25076 419 -25042
rect 453 -25076 500 -25042
rect 372 -25082 500 -25076
rect -40 -25152 -28 -25145
rect -334 -25186 -274 -25179
rect -34 -25179 -28 -25152
rect 6 -25152 20 -25145
rect 264 -25145 310 -25114
rect 6 -25179 12 -25152
rect -630 -25251 -624 -25217
rect -590 -25251 -584 -25217
rect -630 -25289 -584 -25251
rect -630 -25323 -624 -25289
rect -590 -25323 -584 -25289
rect -630 -25361 -584 -25323
rect -630 -25395 -624 -25361
rect -590 -25395 -584 -25361
rect -630 -25433 -584 -25395
rect -630 -25467 -624 -25433
rect -590 -25467 -584 -25433
rect -630 -25505 -584 -25467
rect -630 -25539 -624 -25505
rect -590 -25539 -584 -25505
rect -630 -25577 -584 -25539
rect -630 -25611 -624 -25577
rect -590 -25611 -584 -25577
rect -630 -25638 -584 -25611
rect -332 -25217 -286 -25186
rect -332 -25251 -326 -25217
rect -292 -25251 -286 -25217
rect -332 -25289 -286 -25251
rect -332 -25323 -326 -25289
rect -292 -25323 -286 -25289
rect -332 -25361 -286 -25323
rect -332 -25395 -326 -25361
rect -292 -25395 -286 -25361
rect -332 -25433 -286 -25395
rect -332 -25467 -326 -25433
rect -292 -25467 -286 -25433
rect -332 -25505 -286 -25467
rect -332 -25539 -326 -25505
rect -292 -25539 -286 -25505
rect -332 -25577 -286 -25539
rect -332 -25611 -326 -25577
rect -292 -25611 -286 -25577
rect -332 -25638 -286 -25611
rect -34 -25217 12 -25179
rect -34 -25251 -28 -25217
rect 6 -25251 12 -25217
rect -34 -25289 12 -25251
rect -34 -25323 -28 -25289
rect 6 -25323 12 -25289
rect -34 -25361 12 -25323
rect -34 -25395 -28 -25361
rect 6 -25395 12 -25361
rect -34 -25433 12 -25395
rect -34 -25467 -28 -25433
rect 6 -25467 12 -25433
rect -34 -25505 12 -25467
rect -34 -25539 -28 -25505
rect 6 -25539 12 -25505
rect -34 -25577 12 -25539
rect -34 -25611 -28 -25577
rect 6 -25611 12 -25577
rect -34 -25638 12 -25611
rect 264 -25179 270 -25145
rect 304 -25179 310 -25145
rect 264 -25217 310 -25179
rect 554 -25145 614 -24998
rect 704 -25036 764 -24998
rect 670 -25042 798 -25036
rect 670 -25076 717 -25042
rect 751 -25076 798 -25042
rect 670 -25082 798 -25076
rect 554 -25179 568 -25145
rect 602 -25179 614 -25145
rect 854 -25145 914 -24998
rect 854 -25152 866 -25145
rect 554 -25182 614 -25179
rect 860 -25179 866 -25152
rect 900 -25152 914 -25145
rect 900 -25179 906 -25152
rect 264 -25251 270 -25217
rect 304 -25251 310 -25217
rect 264 -25289 310 -25251
rect 264 -25323 270 -25289
rect 304 -25323 310 -25289
rect 264 -25361 310 -25323
rect 264 -25395 270 -25361
rect 304 -25395 310 -25361
rect 264 -25433 310 -25395
rect 264 -25467 270 -25433
rect 304 -25467 310 -25433
rect 264 -25505 310 -25467
rect 264 -25539 270 -25505
rect 304 -25539 310 -25505
rect 264 -25577 310 -25539
rect 264 -25611 270 -25577
rect 304 -25611 310 -25577
rect -928 -25662 -922 -25649
rect -936 -25664 -922 -25662
rect -1220 -25702 -1186 -25683
rect -938 -25683 -922 -25664
rect -888 -25662 -882 -25649
rect -624 -25649 -590 -25638
rect -888 -25683 -876 -25662
rect -938 -25702 -876 -25683
rect -624 -25702 -590 -25683
rect -326 -25649 -292 -25638
rect -326 -25702 -292 -25683
rect -28 -25649 6 -25638
rect 264 -25649 310 -25611
rect 264 -25654 270 -25649
rect -28 -25702 6 -25683
rect 256 -25683 270 -25654
rect 304 -25654 310 -25649
rect 562 -25217 608 -25182
rect 562 -25251 568 -25217
rect 602 -25251 608 -25217
rect 562 -25289 608 -25251
rect 562 -25323 568 -25289
rect 602 -25323 608 -25289
rect 562 -25361 608 -25323
rect 562 -25395 568 -25361
rect 602 -25395 608 -25361
rect 562 -25433 608 -25395
rect 562 -25467 568 -25433
rect 602 -25467 608 -25433
rect 562 -25505 608 -25467
rect 562 -25539 568 -25505
rect 602 -25539 608 -25505
rect 562 -25577 608 -25539
rect 562 -25611 568 -25577
rect 602 -25611 608 -25577
rect 562 -25649 608 -25611
rect 304 -25666 316 -25654
rect 304 -25683 318 -25666
rect 256 -25702 318 -25683
rect -2012 -25752 -1884 -25746
rect -1118 -25752 -990 -25746
rect -2012 -25786 -1965 -25752
rect -1931 -25786 -1884 -25752
rect -1702 -25758 -1667 -25752
rect -2012 -25792 -1884 -25786
rect -1714 -25786 -1667 -25758
rect -1633 -25758 -1598 -25752
rect -1404 -25758 -1369 -25752
rect -1633 -25786 -1586 -25758
rect -1714 -25792 -1586 -25786
rect -1416 -25786 -1369 -25758
rect -1335 -25758 -1300 -25752
rect -1335 -25786 -1288 -25758
rect -1416 -25792 -1288 -25786
rect -1118 -25786 -1071 -25752
rect -1037 -25786 -990 -25752
rect -1118 -25792 -990 -25786
rect -1680 -25840 -1620 -25792
rect -1382 -25840 -1322 -25792
rect -4946 -25874 -3252 -25870
rect -4946 -25926 -4942 -25874
rect -4890 -25926 -3252 -25874
rect -2676 -25844 -2604 -25840
rect -2676 -25896 -2666 -25844
rect -2614 -25896 -2604 -25844
rect -2676 -25900 -2604 -25896
rect -2426 -25900 -2066 -25840
rect -1686 -25844 -1614 -25840
rect -1686 -25896 -1676 -25844
rect -1624 -25896 -1614 -25844
rect -1686 -25900 -1614 -25896
rect -1388 -25844 -1316 -25840
rect -1388 -25896 -1378 -25844
rect -1326 -25896 -1316 -25844
rect -1388 -25900 -1316 -25896
rect -4946 -25930 -3252 -25926
rect -4946 -25936 -4886 -25930
rect -2126 -25940 -2066 -25900
rect -938 -25940 -878 -25702
rect -820 -25752 -692 -25746
rect -486 -25752 -426 -25750
rect 74 -25752 202 -25746
rect -820 -25786 -773 -25752
rect -739 -25786 -692 -25752
rect -510 -25780 -475 -25752
rect -820 -25792 -692 -25786
rect -522 -25786 -475 -25780
rect -441 -25780 -406 -25752
rect -212 -25780 -177 -25752
rect -441 -25786 -394 -25780
rect -522 -25792 -394 -25786
rect -224 -25786 -177 -25780
rect -143 -25780 -108 -25752
rect -143 -25786 -96 -25780
rect -224 -25792 -96 -25786
rect 74 -25786 121 -25752
rect 155 -25786 202 -25752
rect 74 -25792 202 -25786
rect -486 -25840 -426 -25792
rect -184 -25840 -124 -25792
rect -492 -25844 -420 -25840
rect -492 -25896 -482 -25844
rect -430 -25896 -420 -25844
rect -492 -25900 -420 -25896
rect -190 -25844 -118 -25840
rect -190 -25896 -180 -25844
rect -128 -25896 -118 -25844
rect -190 -25900 -118 -25896
rect 258 -25940 318 -25702
rect 562 -25683 568 -25649
rect 602 -25683 608 -25649
rect 562 -25714 608 -25683
rect 860 -25217 906 -25179
rect 860 -25251 866 -25217
rect 900 -25251 906 -25217
rect 860 -25289 906 -25251
rect 860 -25323 866 -25289
rect 900 -25323 906 -25289
rect 860 -25361 906 -25323
rect 860 -25395 866 -25361
rect 900 -25395 906 -25361
rect 860 -25433 906 -25395
rect 860 -25467 866 -25433
rect 900 -25467 906 -25433
rect 860 -25505 906 -25467
rect 860 -25539 866 -25505
rect 900 -25539 906 -25505
rect 860 -25577 906 -25539
rect 860 -25611 866 -25577
rect 900 -25611 906 -25577
rect 860 -25649 906 -25611
rect 860 -25683 866 -25649
rect 900 -25683 906 -25649
rect 860 -25714 906 -25683
rect 372 -25752 500 -25746
rect 372 -25786 419 -25752
rect 453 -25786 500 -25752
rect 372 -25792 500 -25786
rect 670 -25752 798 -25746
rect 670 -25786 717 -25752
rect 751 -25786 798 -25752
rect 670 -25792 798 -25786
rect 952 -25940 1012 -23784
rect 1076 -22726 1136 -22716
rect 1076 -22778 1080 -22726
rect 1132 -22778 1136 -22726
rect 1076 -24914 1136 -22778
rect 1976 -23544 2036 -14060
rect 1970 -23548 2042 -23544
rect 1970 -23600 1980 -23548
rect 2032 -23600 2042 -23548
rect 1970 -23604 2042 -23600
rect 2110 -23762 2170 -13854
rect 2336 -15116 2396 -11412
rect 3070 -11594 22482 -11534
rect 3070 -11640 3130 -11594
rect 2864 -11646 3352 -11640
rect 2864 -11680 2911 -11646
rect 2945 -11680 2983 -11646
rect 3017 -11680 3055 -11646
rect 3089 -11680 3127 -11646
rect 3161 -11680 3199 -11646
rect 3233 -11680 3271 -11646
rect 3305 -11680 3352 -11646
rect 2864 -11686 3352 -11680
rect 2576 -11749 2622 -11718
rect 2576 -11783 2582 -11749
rect 2616 -11783 2622 -11749
rect 2576 -11821 2622 -11783
rect 2576 -11855 2582 -11821
rect 2616 -11855 2622 -11821
rect 2576 -11893 2622 -11855
rect 2576 -11927 2582 -11893
rect 2616 -11927 2622 -11893
rect 2576 -11965 2622 -11927
rect 2576 -11999 2582 -11965
rect 2616 -11999 2622 -11965
rect 2576 -12037 2622 -11999
rect 2576 -12071 2582 -12037
rect 2616 -12071 2622 -12037
rect 2576 -12109 2622 -12071
rect 2576 -12143 2582 -12109
rect 2616 -12143 2622 -12109
rect 2576 -12181 2622 -12143
rect 2576 -12215 2582 -12181
rect 2616 -12215 2622 -12181
rect 2576 -12253 2622 -12215
rect 2576 -12272 2582 -12253
rect 2568 -12287 2582 -12272
rect 2616 -12272 2622 -12253
rect 3586 -11749 3646 -11594
rect 4098 -11640 4158 -11594
rect 5106 -11640 5166 -11594
rect 3882 -11646 4370 -11640
rect 3882 -11680 3929 -11646
rect 3963 -11680 4001 -11646
rect 4035 -11680 4073 -11646
rect 4107 -11680 4145 -11646
rect 4179 -11680 4217 -11646
rect 4251 -11680 4289 -11646
rect 4323 -11680 4370 -11646
rect 3882 -11686 4370 -11680
rect 4900 -11646 5388 -11640
rect 4900 -11680 4947 -11646
rect 4981 -11680 5019 -11646
rect 5053 -11680 5091 -11646
rect 5125 -11680 5163 -11646
rect 5197 -11680 5235 -11646
rect 5269 -11680 5307 -11646
rect 5341 -11680 5388 -11646
rect 4900 -11686 5388 -11680
rect 3586 -11783 3600 -11749
rect 3634 -11783 3646 -11749
rect 3586 -11821 3646 -11783
rect 3586 -11855 3600 -11821
rect 3634 -11855 3646 -11821
rect 3586 -11893 3646 -11855
rect 3586 -11927 3600 -11893
rect 3634 -11927 3646 -11893
rect 3586 -11965 3646 -11927
rect 3586 -11999 3600 -11965
rect 3634 -11999 3646 -11965
rect 3586 -12037 3646 -11999
rect 3586 -12071 3600 -12037
rect 3634 -12071 3646 -12037
rect 3586 -12109 3646 -12071
rect 3586 -12143 3600 -12109
rect 3634 -12143 3646 -12109
rect 3586 -12181 3646 -12143
rect 3586 -12215 3600 -12181
rect 3634 -12215 3646 -12181
rect 3586 -12253 3646 -12215
rect 2616 -12287 2628 -12272
rect 2568 -12448 2628 -12287
rect 3586 -12287 3600 -12253
rect 3634 -12287 3646 -12253
rect 4612 -11749 4658 -11718
rect 4612 -11783 4618 -11749
rect 4652 -11783 4658 -11749
rect 4612 -11821 4658 -11783
rect 4612 -11855 4618 -11821
rect 4652 -11855 4658 -11821
rect 4612 -11893 4658 -11855
rect 4612 -11927 4618 -11893
rect 4652 -11927 4658 -11893
rect 4612 -11965 4658 -11927
rect 4612 -11999 4618 -11965
rect 4652 -11999 4658 -11965
rect 4612 -12037 4658 -11999
rect 4612 -12071 4618 -12037
rect 4652 -12071 4658 -12037
rect 4612 -12109 4658 -12071
rect 4612 -12143 4618 -12109
rect 4652 -12143 4658 -12109
rect 4612 -12181 4658 -12143
rect 4612 -12215 4618 -12181
rect 4652 -12215 4658 -12181
rect 4612 -12253 4658 -12215
rect 4612 -12268 4618 -12253
rect 2864 -12356 3352 -12350
rect 2864 -12390 2911 -12356
rect 2945 -12390 2983 -12356
rect 3017 -12390 3055 -12356
rect 3089 -12390 3127 -12356
rect 3161 -12390 3199 -12356
rect 3233 -12390 3271 -12356
rect 3305 -12390 3352 -12356
rect 2864 -12396 3352 -12390
rect 2562 -12452 2634 -12448
rect 2562 -12504 2572 -12452
rect 2624 -12504 2634 -12452
rect 2562 -12508 2634 -12504
rect 2568 -12983 2628 -12508
rect 3076 -12874 3136 -12396
rect 3586 -12546 3646 -12287
rect 4604 -12287 4618 -12268
rect 4652 -12268 4658 -12253
rect 5624 -11749 5684 -11594
rect 6116 -11640 6176 -11594
rect 7128 -11640 7188 -11594
rect 5918 -11646 6406 -11640
rect 5918 -11680 5965 -11646
rect 5999 -11680 6037 -11646
rect 6071 -11680 6109 -11646
rect 6143 -11680 6181 -11646
rect 6215 -11680 6253 -11646
rect 6287 -11680 6325 -11646
rect 6359 -11680 6406 -11646
rect 5918 -11686 6406 -11680
rect 6936 -11646 7424 -11640
rect 6936 -11680 6983 -11646
rect 7017 -11680 7055 -11646
rect 7089 -11680 7127 -11646
rect 7161 -11680 7199 -11646
rect 7233 -11680 7271 -11646
rect 7305 -11680 7343 -11646
rect 7377 -11680 7424 -11646
rect 6936 -11686 7424 -11680
rect 5624 -11783 5636 -11749
rect 5670 -11783 5684 -11749
rect 5624 -11821 5684 -11783
rect 5624 -11855 5636 -11821
rect 5670 -11855 5684 -11821
rect 5624 -11893 5684 -11855
rect 5624 -11927 5636 -11893
rect 5670 -11927 5684 -11893
rect 5624 -11965 5684 -11927
rect 5624 -11999 5636 -11965
rect 5670 -11999 5684 -11965
rect 5624 -12037 5684 -11999
rect 5624 -12071 5636 -12037
rect 5670 -12071 5684 -12037
rect 5624 -12109 5684 -12071
rect 5624 -12143 5636 -12109
rect 5670 -12143 5684 -12109
rect 5624 -12181 5684 -12143
rect 5624 -12215 5636 -12181
rect 5670 -12215 5684 -12181
rect 5624 -12253 5684 -12215
rect 4652 -12287 4664 -12268
rect 3882 -12356 4370 -12350
rect 3882 -12390 3929 -12356
rect 3963 -12390 4001 -12356
rect 4035 -12390 4073 -12356
rect 4107 -12390 4145 -12356
rect 4179 -12390 4217 -12356
rect 4251 -12390 4289 -12356
rect 4323 -12390 4370 -12356
rect 3882 -12396 4370 -12390
rect 3580 -12550 3652 -12546
rect 3580 -12602 3590 -12550
rect 3642 -12602 3652 -12550
rect 3580 -12606 3652 -12602
rect 2864 -12880 3352 -12874
rect 2864 -12914 2911 -12880
rect 2945 -12914 2983 -12880
rect 3017 -12914 3055 -12880
rect 3089 -12914 3127 -12880
rect 3161 -12914 3199 -12880
rect 3233 -12914 3271 -12880
rect 3305 -12914 3352 -12880
rect 2864 -12920 3352 -12914
rect 2568 -12998 2582 -12983
rect 2576 -13017 2582 -12998
rect 2616 -12998 2628 -12983
rect 3586 -12983 3646 -12606
rect 4078 -12874 4138 -12396
rect 4604 -12448 4664 -12287
rect 5624 -12287 5636 -12253
rect 5670 -12287 5684 -12253
rect 6648 -11749 6694 -11718
rect 6648 -11783 6654 -11749
rect 6688 -11783 6694 -11749
rect 6648 -11821 6694 -11783
rect 6648 -11855 6654 -11821
rect 6688 -11855 6694 -11821
rect 6648 -11893 6694 -11855
rect 6648 -11927 6654 -11893
rect 6688 -11927 6694 -11893
rect 6648 -11965 6694 -11927
rect 6648 -11999 6654 -11965
rect 6688 -11999 6694 -11965
rect 6648 -12037 6694 -11999
rect 6648 -12071 6654 -12037
rect 6688 -12071 6694 -12037
rect 6648 -12109 6694 -12071
rect 6648 -12143 6654 -12109
rect 6688 -12143 6694 -12109
rect 6648 -12181 6694 -12143
rect 6648 -12215 6654 -12181
rect 6688 -12215 6694 -12181
rect 6648 -12253 6694 -12215
rect 6648 -12276 6654 -12253
rect 5100 -12350 5160 -12348
rect 4900 -12356 5388 -12350
rect 4900 -12390 4947 -12356
rect 4981 -12390 5019 -12356
rect 5053 -12390 5091 -12356
rect 5125 -12390 5163 -12356
rect 5197 -12390 5235 -12356
rect 5269 -12390 5307 -12356
rect 5341 -12390 5388 -12356
rect 4900 -12396 5388 -12390
rect 4598 -12452 4670 -12448
rect 4598 -12504 4608 -12452
rect 4660 -12504 4670 -12452
rect 4598 -12508 4670 -12504
rect 3882 -12880 4370 -12874
rect 3882 -12914 3929 -12880
rect 3963 -12914 4001 -12880
rect 4035 -12914 4073 -12880
rect 4107 -12914 4145 -12880
rect 4179 -12914 4217 -12880
rect 4251 -12914 4289 -12880
rect 4323 -12914 4370 -12880
rect 3882 -12920 4370 -12914
rect 2616 -13017 2622 -12998
rect 3586 -13012 3600 -12983
rect 2576 -13055 2622 -13017
rect 2576 -13089 2582 -13055
rect 2616 -13089 2622 -13055
rect 2576 -13127 2622 -13089
rect 2576 -13161 2582 -13127
rect 2616 -13161 2622 -13127
rect 2576 -13199 2622 -13161
rect 2576 -13233 2582 -13199
rect 2616 -13233 2622 -13199
rect 2576 -13271 2622 -13233
rect 2576 -13305 2582 -13271
rect 2616 -13305 2622 -13271
rect 2576 -13343 2622 -13305
rect 2576 -13377 2582 -13343
rect 2616 -13377 2622 -13343
rect 2576 -13415 2622 -13377
rect 2576 -13449 2582 -13415
rect 2616 -13449 2622 -13415
rect 2576 -13487 2622 -13449
rect 2576 -13521 2582 -13487
rect 2616 -13521 2622 -13487
rect 2576 -13552 2622 -13521
rect 3594 -13017 3600 -13012
rect 3634 -13012 3646 -12983
rect 4604 -12983 4664 -12508
rect 5100 -12874 5160 -12396
rect 5624 -12546 5684 -12287
rect 6638 -12287 6654 -12276
rect 6688 -12276 6694 -12253
rect 7658 -11749 7718 -11594
rect 8176 -11640 8236 -11594
rect 9164 -11640 9224 -11594
rect 7954 -11646 8442 -11640
rect 7954 -11680 8001 -11646
rect 8035 -11680 8073 -11646
rect 8107 -11680 8145 -11646
rect 8179 -11680 8217 -11646
rect 8251 -11680 8289 -11646
rect 8323 -11680 8361 -11646
rect 8395 -11680 8442 -11646
rect 7954 -11686 8442 -11680
rect 8972 -11646 9460 -11640
rect 8972 -11680 9019 -11646
rect 9053 -11680 9091 -11646
rect 9125 -11680 9163 -11646
rect 9197 -11680 9235 -11646
rect 9269 -11680 9307 -11646
rect 9341 -11680 9379 -11646
rect 9413 -11680 9460 -11646
rect 8972 -11686 9460 -11680
rect 7658 -11783 7672 -11749
rect 7706 -11783 7718 -11749
rect 7658 -11821 7718 -11783
rect 7658 -11855 7672 -11821
rect 7706 -11855 7718 -11821
rect 7658 -11893 7718 -11855
rect 7658 -11927 7672 -11893
rect 7706 -11927 7718 -11893
rect 7658 -11965 7718 -11927
rect 7658 -11999 7672 -11965
rect 7706 -11999 7718 -11965
rect 7658 -12037 7718 -11999
rect 7658 -12071 7672 -12037
rect 7706 -12071 7718 -12037
rect 7658 -12109 7718 -12071
rect 7658 -12143 7672 -12109
rect 7706 -12143 7718 -12109
rect 7658 -12181 7718 -12143
rect 7658 -12215 7672 -12181
rect 7706 -12215 7718 -12181
rect 7658 -12253 7718 -12215
rect 6688 -12287 6698 -12276
rect 5918 -12356 6406 -12350
rect 5918 -12390 5965 -12356
rect 5999 -12390 6037 -12356
rect 6071 -12390 6109 -12356
rect 6143 -12390 6181 -12356
rect 6215 -12390 6253 -12356
rect 6287 -12390 6325 -12356
rect 6359 -12390 6406 -12356
rect 5918 -12396 6406 -12390
rect 6638 -12448 6698 -12287
rect 7658 -12287 7672 -12253
rect 7706 -12287 7718 -12253
rect 8684 -11749 8730 -11718
rect 8684 -11783 8690 -11749
rect 8724 -11783 8730 -11749
rect 8684 -11821 8730 -11783
rect 8684 -11855 8690 -11821
rect 8724 -11855 8730 -11821
rect 8684 -11893 8730 -11855
rect 8684 -11927 8690 -11893
rect 8724 -11927 8730 -11893
rect 8684 -11965 8730 -11927
rect 8684 -11999 8690 -11965
rect 8724 -11999 8730 -11965
rect 8684 -12037 8730 -11999
rect 8684 -12071 8690 -12037
rect 8724 -12071 8730 -12037
rect 8684 -12109 8730 -12071
rect 8684 -12143 8690 -12109
rect 8724 -12143 8730 -12109
rect 8684 -12181 8730 -12143
rect 8684 -12215 8690 -12181
rect 8724 -12215 8730 -12181
rect 8684 -12253 8730 -12215
rect 8684 -12262 8690 -12253
rect 6936 -12356 7424 -12350
rect 6936 -12390 6983 -12356
rect 7017 -12390 7055 -12356
rect 7089 -12390 7127 -12356
rect 7161 -12390 7199 -12356
rect 7233 -12390 7271 -12356
rect 7305 -12390 7343 -12356
rect 7377 -12390 7424 -12356
rect 6936 -12396 7424 -12390
rect 6632 -12452 6704 -12448
rect 6632 -12504 6642 -12452
rect 6694 -12504 6704 -12452
rect 6632 -12508 6704 -12504
rect 7658 -12546 7718 -12287
rect 8678 -12287 8690 -12262
rect 8724 -12262 8730 -12253
rect 9692 -11749 9752 -11594
rect 10208 -11640 10268 -11594
rect 11210 -11640 11270 -11594
rect 9990 -11646 10478 -11640
rect 9990 -11680 10037 -11646
rect 10071 -11680 10109 -11646
rect 10143 -11680 10181 -11646
rect 10215 -11680 10253 -11646
rect 10287 -11680 10325 -11646
rect 10359 -11680 10397 -11646
rect 10431 -11680 10478 -11646
rect 9990 -11686 10478 -11680
rect 11008 -11646 11496 -11640
rect 11008 -11680 11055 -11646
rect 11089 -11680 11127 -11646
rect 11161 -11680 11199 -11646
rect 11233 -11680 11271 -11646
rect 11305 -11680 11343 -11646
rect 11377 -11680 11415 -11646
rect 11449 -11680 11496 -11646
rect 11008 -11686 11496 -11680
rect 9692 -11783 9708 -11749
rect 9742 -11783 9752 -11749
rect 9692 -11821 9752 -11783
rect 9692 -11855 9708 -11821
rect 9742 -11855 9752 -11821
rect 9692 -11893 9752 -11855
rect 9692 -11927 9708 -11893
rect 9742 -11927 9752 -11893
rect 9692 -11965 9752 -11927
rect 9692 -11999 9708 -11965
rect 9742 -11999 9752 -11965
rect 9692 -12037 9752 -11999
rect 9692 -12071 9708 -12037
rect 9742 -12071 9752 -12037
rect 9692 -12109 9752 -12071
rect 9692 -12143 9708 -12109
rect 9742 -12143 9752 -12109
rect 9692 -12181 9752 -12143
rect 9692 -12215 9708 -12181
rect 9742 -12215 9752 -12181
rect 9692 -12253 9752 -12215
rect 8724 -12287 8738 -12262
rect 7954 -12356 8442 -12350
rect 7954 -12390 8001 -12356
rect 8035 -12390 8073 -12356
rect 8107 -12390 8145 -12356
rect 8179 -12390 8217 -12356
rect 8251 -12390 8289 -12356
rect 8323 -12390 8361 -12356
rect 8395 -12390 8442 -12356
rect 7954 -12396 8442 -12390
rect 8678 -12448 8738 -12287
rect 9692 -12287 9708 -12253
rect 9742 -12287 9752 -12253
rect 10720 -11749 10766 -11718
rect 10720 -11783 10726 -11749
rect 10760 -11783 10766 -11749
rect 10720 -11821 10766 -11783
rect 10720 -11855 10726 -11821
rect 10760 -11855 10766 -11821
rect 10720 -11893 10766 -11855
rect 10720 -11927 10726 -11893
rect 10760 -11927 10766 -11893
rect 10720 -11965 10766 -11927
rect 10720 -11999 10726 -11965
rect 10760 -11999 10766 -11965
rect 10720 -12037 10766 -11999
rect 10720 -12071 10726 -12037
rect 10760 -12071 10766 -12037
rect 10720 -12109 10766 -12071
rect 10720 -12143 10726 -12109
rect 10760 -12143 10766 -12109
rect 10720 -12181 10766 -12143
rect 10720 -12215 10726 -12181
rect 10760 -12215 10766 -12181
rect 10720 -12253 10766 -12215
rect 10720 -12266 10726 -12253
rect 8972 -12356 9460 -12350
rect 8972 -12390 9019 -12356
rect 9053 -12390 9091 -12356
rect 9125 -12390 9163 -12356
rect 9197 -12390 9235 -12356
rect 9269 -12390 9307 -12356
rect 9341 -12390 9379 -12356
rect 9413 -12390 9460 -12356
rect 8972 -12396 9460 -12390
rect 8672 -12452 8744 -12448
rect 8672 -12504 8682 -12452
rect 8734 -12504 8744 -12452
rect 8672 -12508 8744 -12504
rect 9692 -12546 9752 -12287
rect 10714 -12287 10726 -12266
rect 10760 -12266 10766 -12253
rect 11732 -11749 11792 -11594
rect 12238 -11640 12298 -11594
rect 13256 -11640 13316 -11594
rect 12026 -11646 12514 -11640
rect 12026 -11680 12073 -11646
rect 12107 -11680 12145 -11646
rect 12179 -11680 12217 -11646
rect 12251 -11680 12289 -11646
rect 12323 -11680 12361 -11646
rect 12395 -11680 12433 -11646
rect 12467 -11680 12514 -11646
rect 12026 -11686 12514 -11680
rect 13044 -11646 13532 -11640
rect 13044 -11680 13091 -11646
rect 13125 -11680 13163 -11646
rect 13197 -11680 13235 -11646
rect 13269 -11680 13307 -11646
rect 13341 -11680 13379 -11646
rect 13413 -11680 13451 -11646
rect 13485 -11680 13532 -11646
rect 13044 -11686 13532 -11680
rect 12238 -11688 12298 -11686
rect 11732 -11783 11744 -11749
rect 11778 -11783 11792 -11749
rect 11732 -11821 11792 -11783
rect 11732 -11855 11744 -11821
rect 11778 -11855 11792 -11821
rect 11732 -11893 11792 -11855
rect 11732 -11927 11744 -11893
rect 11778 -11927 11792 -11893
rect 11732 -11965 11792 -11927
rect 11732 -11999 11744 -11965
rect 11778 -11999 11792 -11965
rect 11732 -12037 11792 -11999
rect 11732 -12071 11744 -12037
rect 11778 -12071 11792 -12037
rect 11732 -12109 11792 -12071
rect 11732 -12143 11744 -12109
rect 11778 -12143 11792 -12109
rect 11732 -12181 11792 -12143
rect 11732 -12215 11744 -12181
rect 11778 -12215 11792 -12181
rect 11732 -12253 11792 -12215
rect 10760 -12287 10774 -12266
rect 9990 -12356 10478 -12350
rect 9990 -12390 10037 -12356
rect 10071 -12390 10109 -12356
rect 10143 -12390 10181 -12356
rect 10215 -12390 10253 -12356
rect 10287 -12390 10325 -12356
rect 10359 -12390 10397 -12356
rect 10431 -12390 10478 -12356
rect 9990 -12396 10478 -12390
rect 10714 -12448 10774 -12287
rect 11732 -12287 11744 -12253
rect 11778 -12287 11792 -12253
rect 12756 -11749 12802 -11718
rect 12756 -11783 12762 -11749
rect 12796 -11783 12802 -11749
rect 12756 -11821 12802 -11783
rect 12756 -11855 12762 -11821
rect 12796 -11855 12802 -11821
rect 12756 -11893 12802 -11855
rect 12756 -11927 12762 -11893
rect 12796 -11927 12802 -11893
rect 12756 -11965 12802 -11927
rect 12756 -11999 12762 -11965
rect 12796 -11999 12802 -11965
rect 12756 -12037 12802 -11999
rect 12756 -12071 12762 -12037
rect 12796 -12071 12802 -12037
rect 12756 -12109 12802 -12071
rect 12756 -12143 12762 -12109
rect 12796 -12143 12802 -12109
rect 12756 -12181 12802 -12143
rect 12756 -12215 12762 -12181
rect 12796 -12215 12802 -12181
rect 12756 -12253 12802 -12215
rect 12756 -12266 12762 -12253
rect 11008 -12356 11496 -12350
rect 11008 -12390 11055 -12356
rect 11089 -12390 11127 -12356
rect 11161 -12390 11199 -12356
rect 11233 -12390 11271 -12356
rect 11305 -12390 11343 -12356
rect 11377 -12390 11415 -12356
rect 11449 -12390 11496 -12356
rect 11008 -12396 11496 -12390
rect 10708 -12452 10780 -12448
rect 10708 -12504 10718 -12452
rect 10770 -12504 10780 -12452
rect 10708 -12508 10780 -12504
rect 11732 -12546 11792 -12287
rect 12748 -12287 12762 -12266
rect 12796 -12266 12802 -12253
rect 13766 -11749 13826 -11594
rect 14274 -11640 14334 -11594
rect 15294 -11640 15354 -11594
rect 14062 -11646 14550 -11640
rect 14062 -11680 14109 -11646
rect 14143 -11680 14181 -11646
rect 14215 -11680 14253 -11646
rect 14287 -11680 14325 -11646
rect 14359 -11680 14397 -11646
rect 14431 -11680 14469 -11646
rect 14503 -11680 14550 -11646
rect 14062 -11686 14550 -11680
rect 15080 -11646 15568 -11640
rect 15080 -11680 15127 -11646
rect 15161 -11680 15199 -11646
rect 15233 -11680 15271 -11646
rect 15305 -11680 15343 -11646
rect 15377 -11680 15415 -11646
rect 15449 -11680 15487 -11646
rect 15521 -11680 15568 -11646
rect 15080 -11686 15568 -11680
rect 13766 -11783 13780 -11749
rect 13814 -11783 13826 -11749
rect 13766 -11821 13826 -11783
rect 13766 -11855 13780 -11821
rect 13814 -11855 13826 -11821
rect 13766 -11893 13826 -11855
rect 13766 -11927 13780 -11893
rect 13814 -11927 13826 -11893
rect 13766 -11965 13826 -11927
rect 13766 -11999 13780 -11965
rect 13814 -11999 13826 -11965
rect 13766 -12037 13826 -11999
rect 13766 -12071 13780 -12037
rect 13814 -12071 13826 -12037
rect 13766 -12109 13826 -12071
rect 13766 -12143 13780 -12109
rect 13814 -12143 13826 -12109
rect 13766 -12181 13826 -12143
rect 13766 -12215 13780 -12181
rect 13814 -12215 13826 -12181
rect 13766 -12253 13826 -12215
rect 12796 -12287 12808 -12266
rect 12026 -12356 12514 -12350
rect 12026 -12390 12073 -12356
rect 12107 -12390 12145 -12356
rect 12179 -12390 12217 -12356
rect 12251 -12390 12289 -12356
rect 12323 -12390 12361 -12356
rect 12395 -12390 12433 -12356
rect 12467 -12390 12514 -12356
rect 12026 -12396 12514 -12390
rect 12748 -12448 12808 -12287
rect 13766 -12287 13780 -12253
rect 13814 -12287 13826 -12253
rect 14792 -11749 14838 -11718
rect 14792 -11783 14798 -11749
rect 14832 -11783 14838 -11749
rect 14792 -11821 14838 -11783
rect 14792 -11855 14798 -11821
rect 14832 -11855 14838 -11821
rect 14792 -11893 14838 -11855
rect 14792 -11927 14798 -11893
rect 14832 -11927 14838 -11893
rect 14792 -11965 14838 -11927
rect 14792 -11999 14798 -11965
rect 14832 -11999 14838 -11965
rect 14792 -12037 14838 -11999
rect 14792 -12071 14798 -12037
rect 14832 -12071 14838 -12037
rect 14792 -12109 14838 -12071
rect 14792 -12143 14798 -12109
rect 14832 -12143 14838 -12109
rect 14792 -12181 14838 -12143
rect 14792 -12215 14798 -12181
rect 14832 -12215 14838 -12181
rect 14792 -12253 14838 -12215
rect 14792 -12260 14798 -12253
rect 13044 -12356 13532 -12350
rect 13044 -12390 13091 -12356
rect 13125 -12390 13163 -12356
rect 13197 -12390 13235 -12356
rect 13269 -12390 13307 -12356
rect 13341 -12390 13379 -12356
rect 13413 -12390 13451 -12356
rect 13485 -12390 13532 -12356
rect 13044 -12396 13532 -12390
rect 12742 -12452 12814 -12448
rect 12742 -12504 12752 -12452
rect 12804 -12504 12814 -12452
rect 12742 -12508 12814 -12504
rect 13766 -12546 13826 -12287
rect 14784 -12287 14798 -12260
rect 14832 -12260 14838 -12253
rect 15804 -11749 15864 -11594
rect 16302 -11640 16362 -11594
rect 17330 -11640 17390 -11594
rect 16098 -11646 16586 -11640
rect 16098 -11680 16145 -11646
rect 16179 -11680 16217 -11646
rect 16251 -11680 16289 -11646
rect 16323 -11680 16361 -11646
rect 16395 -11680 16433 -11646
rect 16467 -11680 16505 -11646
rect 16539 -11680 16586 -11646
rect 16098 -11686 16586 -11680
rect 17116 -11646 17604 -11640
rect 17116 -11680 17163 -11646
rect 17197 -11680 17235 -11646
rect 17269 -11680 17307 -11646
rect 17341 -11680 17379 -11646
rect 17413 -11680 17451 -11646
rect 17485 -11680 17523 -11646
rect 17557 -11680 17604 -11646
rect 17116 -11686 17604 -11680
rect 15804 -11783 15816 -11749
rect 15850 -11783 15864 -11749
rect 15804 -11821 15864 -11783
rect 15804 -11855 15816 -11821
rect 15850 -11855 15864 -11821
rect 15804 -11893 15864 -11855
rect 15804 -11927 15816 -11893
rect 15850 -11927 15864 -11893
rect 15804 -11965 15864 -11927
rect 15804 -11999 15816 -11965
rect 15850 -11999 15864 -11965
rect 15804 -12037 15864 -11999
rect 15804 -12071 15816 -12037
rect 15850 -12071 15864 -12037
rect 15804 -12109 15864 -12071
rect 15804 -12143 15816 -12109
rect 15850 -12143 15864 -12109
rect 15804 -12181 15864 -12143
rect 15804 -12215 15816 -12181
rect 15850 -12215 15864 -12181
rect 15804 -12253 15864 -12215
rect 14832 -12287 14844 -12260
rect 14062 -12356 14550 -12350
rect 14062 -12390 14109 -12356
rect 14143 -12390 14181 -12356
rect 14215 -12390 14253 -12356
rect 14287 -12390 14325 -12356
rect 14359 -12390 14397 -12356
rect 14431 -12390 14469 -12356
rect 14503 -12390 14550 -12356
rect 14062 -12396 14550 -12390
rect 14784 -12448 14844 -12287
rect 15804 -12287 15816 -12253
rect 15850 -12287 15864 -12253
rect 16828 -11749 16874 -11718
rect 16828 -11783 16834 -11749
rect 16868 -11783 16874 -11749
rect 16828 -11821 16874 -11783
rect 16828 -11855 16834 -11821
rect 16868 -11855 16874 -11821
rect 16828 -11893 16874 -11855
rect 16828 -11927 16834 -11893
rect 16868 -11927 16874 -11893
rect 16828 -11965 16874 -11927
rect 16828 -11999 16834 -11965
rect 16868 -11999 16874 -11965
rect 16828 -12037 16874 -11999
rect 16828 -12071 16834 -12037
rect 16868 -12071 16874 -12037
rect 16828 -12109 16874 -12071
rect 16828 -12143 16834 -12109
rect 16868 -12143 16874 -12109
rect 16828 -12181 16874 -12143
rect 16828 -12215 16834 -12181
rect 16868 -12215 16874 -12181
rect 16828 -12253 16874 -12215
rect 16828 -12258 16834 -12253
rect 15080 -12356 15568 -12350
rect 15080 -12390 15127 -12356
rect 15161 -12390 15199 -12356
rect 15233 -12390 15271 -12356
rect 15305 -12390 15343 -12356
rect 15377 -12390 15415 -12356
rect 15449 -12390 15487 -12356
rect 15521 -12390 15568 -12356
rect 15080 -12396 15568 -12390
rect 14778 -12452 14850 -12448
rect 14778 -12504 14788 -12452
rect 14840 -12504 14850 -12452
rect 14778 -12508 14850 -12504
rect 15804 -12546 15864 -12287
rect 16820 -12287 16834 -12258
rect 16868 -12258 16874 -12253
rect 17836 -11749 17896 -11594
rect 18332 -11640 18392 -11594
rect 19362 -11640 19422 -11594
rect 18134 -11646 18622 -11640
rect 18134 -11680 18181 -11646
rect 18215 -11680 18253 -11646
rect 18287 -11680 18325 -11646
rect 18359 -11680 18397 -11646
rect 18431 -11680 18469 -11646
rect 18503 -11680 18541 -11646
rect 18575 -11680 18622 -11646
rect 18134 -11686 18622 -11680
rect 19152 -11646 19640 -11640
rect 19152 -11680 19199 -11646
rect 19233 -11680 19271 -11646
rect 19305 -11680 19343 -11646
rect 19377 -11680 19415 -11646
rect 19449 -11680 19487 -11646
rect 19521 -11680 19559 -11646
rect 19593 -11680 19640 -11646
rect 19152 -11686 19640 -11680
rect 17836 -11783 17852 -11749
rect 17886 -11783 17896 -11749
rect 17836 -11821 17896 -11783
rect 17836 -11855 17852 -11821
rect 17886 -11855 17896 -11821
rect 17836 -11893 17896 -11855
rect 17836 -11927 17852 -11893
rect 17886 -11927 17896 -11893
rect 17836 -11965 17896 -11927
rect 17836 -11999 17852 -11965
rect 17886 -11999 17896 -11965
rect 17836 -12037 17896 -11999
rect 17836 -12071 17852 -12037
rect 17886 -12071 17896 -12037
rect 17836 -12109 17896 -12071
rect 17836 -12143 17852 -12109
rect 17886 -12143 17896 -12109
rect 17836 -12181 17896 -12143
rect 17836 -12215 17852 -12181
rect 17886 -12215 17896 -12181
rect 17836 -12253 17896 -12215
rect 18864 -11749 18910 -11718
rect 18864 -11783 18870 -11749
rect 18904 -11783 18910 -11749
rect 18864 -11821 18910 -11783
rect 18864 -11855 18870 -11821
rect 18904 -11855 18910 -11821
rect 18864 -11893 18910 -11855
rect 18864 -11927 18870 -11893
rect 18904 -11927 18910 -11893
rect 18864 -11965 18910 -11927
rect 18864 -11999 18870 -11965
rect 18904 -11999 18910 -11965
rect 18864 -12037 18910 -11999
rect 18864 -12071 18870 -12037
rect 18904 -12071 18910 -12037
rect 18864 -12109 18910 -12071
rect 18864 -12143 18870 -12109
rect 18904 -12143 18910 -12109
rect 18864 -12181 18910 -12143
rect 18864 -12215 18870 -12181
rect 18904 -12215 18910 -12181
rect 18864 -12252 18910 -12215
rect 19874 -11749 19934 -11594
rect 20410 -11640 20470 -11594
rect 21384 -11640 21444 -11594
rect 20170 -11646 20658 -11640
rect 20170 -11680 20217 -11646
rect 20251 -11680 20289 -11646
rect 20323 -11680 20361 -11646
rect 20395 -11680 20433 -11646
rect 20467 -11680 20505 -11646
rect 20539 -11680 20577 -11646
rect 20611 -11680 20658 -11646
rect 20170 -11686 20658 -11680
rect 21188 -11646 21676 -11640
rect 21188 -11680 21235 -11646
rect 21269 -11680 21307 -11646
rect 21341 -11680 21379 -11646
rect 21413 -11680 21451 -11646
rect 21485 -11680 21523 -11646
rect 21557 -11680 21595 -11646
rect 21629 -11680 21676 -11646
rect 21188 -11686 21676 -11680
rect 19874 -11783 19888 -11749
rect 19922 -11783 19934 -11749
rect 19874 -11821 19934 -11783
rect 19874 -11855 19888 -11821
rect 19922 -11855 19934 -11821
rect 19874 -11893 19934 -11855
rect 19874 -11927 19888 -11893
rect 19922 -11927 19934 -11893
rect 19874 -11965 19934 -11927
rect 19874 -11999 19888 -11965
rect 19922 -11999 19934 -11965
rect 19874 -12037 19934 -11999
rect 19874 -12071 19888 -12037
rect 19922 -12071 19934 -12037
rect 19874 -12109 19934 -12071
rect 19874 -12143 19888 -12109
rect 19922 -12143 19934 -12109
rect 19874 -12181 19934 -12143
rect 19874 -12215 19888 -12181
rect 19922 -12215 19934 -12181
rect 16868 -12287 16880 -12258
rect 16098 -12356 16586 -12350
rect 16098 -12390 16145 -12356
rect 16179 -12390 16217 -12356
rect 16251 -12390 16289 -12356
rect 16323 -12390 16361 -12356
rect 16395 -12390 16433 -12356
rect 16467 -12390 16505 -12356
rect 16539 -12390 16586 -12356
rect 16098 -12396 16586 -12390
rect 16820 -12448 16880 -12287
rect 17836 -12287 17852 -12253
rect 17886 -12287 17896 -12253
rect 17116 -12356 17604 -12350
rect 17116 -12390 17163 -12356
rect 17197 -12390 17235 -12356
rect 17269 -12390 17307 -12356
rect 17341 -12390 17379 -12356
rect 17413 -12390 17451 -12356
rect 17485 -12390 17523 -12356
rect 17557 -12390 17604 -12356
rect 17116 -12396 17604 -12390
rect 16814 -12452 16886 -12448
rect 16814 -12504 16824 -12452
rect 16876 -12504 16886 -12452
rect 16814 -12508 16886 -12504
rect 17836 -12546 17896 -12287
rect 18856 -12253 18916 -12252
rect 18856 -12287 18870 -12253
rect 18904 -12287 18916 -12253
rect 18134 -12356 18622 -12350
rect 18134 -12390 18181 -12356
rect 18215 -12390 18253 -12356
rect 18287 -12390 18325 -12356
rect 18359 -12390 18397 -12356
rect 18431 -12390 18469 -12356
rect 18503 -12390 18541 -12356
rect 18575 -12390 18622 -12356
rect 18134 -12396 18622 -12390
rect 18856 -12448 18916 -12287
rect 19874 -12253 19934 -12215
rect 19874 -12287 19888 -12253
rect 19922 -12287 19934 -12253
rect 20900 -11749 20946 -11718
rect 20900 -11783 20906 -11749
rect 20940 -11783 20946 -11749
rect 20900 -11821 20946 -11783
rect 20900 -11855 20906 -11821
rect 20940 -11855 20946 -11821
rect 20900 -11893 20946 -11855
rect 20900 -11927 20906 -11893
rect 20940 -11927 20946 -11893
rect 20900 -11965 20946 -11927
rect 20900 -11999 20906 -11965
rect 20940 -11999 20946 -11965
rect 20900 -12037 20946 -11999
rect 20900 -12071 20906 -12037
rect 20940 -12071 20946 -12037
rect 20900 -12109 20946 -12071
rect 20900 -12143 20906 -12109
rect 20940 -12143 20946 -12109
rect 20900 -12181 20946 -12143
rect 20900 -12215 20906 -12181
rect 20940 -12215 20946 -12181
rect 20900 -12253 20946 -12215
rect 20900 -12260 20906 -12253
rect 19152 -12356 19640 -12350
rect 19152 -12390 19199 -12356
rect 19233 -12390 19271 -12356
rect 19305 -12390 19343 -12356
rect 19377 -12390 19415 -12356
rect 19449 -12390 19487 -12356
rect 19521 -12390 19559 -12356
rect 19593 -12390 19640 -12356
rect 19152 -12396 19640 -12390
rect 18850 -12452 18922 -12448
rect 18850 -12504 18860 -12452
rect 18912 -12504 18922 -12452
rect 18850 -12508 18922 -12504
rect 19874 -12546 19934 -12287
rect 20894 -12287 20906 -12260
rect 20940 -12260 20946 -12253
rect 21912 -11749 21972 -11594
rect 22422 -11640 22482 -11594
rect 22206 -11646 22694 -11640
rect 22206 -11680 22253 -11646
rect 22287 -11680 22325 -11646
rect 22359 -11680 22397 -11646
rect 22431 -11680 22469 -11646
rect 22503 -11680 22541 -11646
rect 22575 -11680 22613 -11646
rect 22647 -11680 22694 -11646
rect 22206 -11686 22694 -11680
rect 21912 -11783 21924 -11749
rect 21958 -11783 21972 -11749
rect 21912 -11821 21972 -11783
rect 21912 -11855 21924 -11821
rect 21958 -11855 21972 -11821
rect 21912 -11893 21972 -11855
rect 21912 -11927 21924 -11893
rect 21958 -11927 21972 -11893
rect 21912 -11965 21972 -11927
rect 21912 -11999 21924 -11965
rect 21958 -11999 21972 -11965
rect 21912 -12037 21972 -11999
rect 21912 -12071 21924 -12037
rect 21958 -12071 21972 -12037
rect 21912 -12109 21972 -12071
rect 21912 -12143 21924 -12109
rect 21958 -12143 21972 -12109
rect 21912 -12181 21972 -12143
rect 21912 -12215 21924 -12181
rect 21958 -12215 21972 -12181
rect 21912 -12253 21972 -12215
rect 22936 -11749 22982 -11718
rect 22936 -11783 22942 -11749
rect 22976 -11783 22982 -11749
rect 22936 -11821 22982 -11783
rect 22936 -11855 22942 -11821
rect 22976 -11855 22982 -11821
rect 22936 -11893 22982 -11855
rect 22936 -11927 22942 -11893
rect 22976 -11927 22982 -11893
rect 22936 -11965 22982 -11927
rect 22936 -11999 22942 -11965
rect 22976 -11999 22982 -11965
rect 22936 -12037 22982 -11999
rect 22936 -12071 22942 -12037
rect 22976 -12071 22982 -12037
rect 22936 -12109 22982 -12071
rect 22936 -12143 22942 -12109
rect 22976 -12143 22982 -12109
rect 22936 -12181 22982 -12143
rect 22936 -12215 22942 -12181
rect 22976 -12215 22982 -12181
rect 22936 -12252 22982 -12215
rect 24816 -12091 24928 -11284
rect 24816 -12125 24855 -12091
rect 24889 -12125 24928 -12091
rect 24816 -12163 24928 -12125
rect 24816 -12197 24855 -12163
rect 24889 -12197 24928 -12163
rect 24816 -12235 24928 -12197
rect 20940 -12287 20954 -12260
rect 20170 -12356 20658 -12350
rect 20170 -12390 20217 -12356
rect 20251 -12390 20289 -12356
rect 20323 -12390 20361 -12356
rect 20395 -12390 20433 -12356
rect 20467 -12390 20505 -12356
rect 20539 -12390 20577 -12356
rect 20611 -12390 20658 -12356
rect 20170 -12396 20658 -12390
rect 5618 -12550 5690 -12546
rect 5618 -12602 5628 -12550
rect 5680 -12602 5690 -12550
rect 5618 -12606 5690 -12602
rect 7652 -12550 7724 -12546
rect 7652 -12602 7662 -12550
rect 7714 -12602 7724 -12550
rect 7652 -12606 7724 -12602
rect 9686 -12550 9758 -12546
rect 9686 -12602 9696 -12550
rect 9748 -12602 9758 -12550
rect 9686 -12606 9758 -12602
rect 11726 -12550 11798 -12546
rect 11726 -12602 11736 -12550
rect 11788 -12602 11798 -12550
rect 11726 -12606 11798 -12602
rect 13760 -12550 13832 -12546
rect 13760 -12602 13770 -12550
rect 13822 -12602 13832 -12550
rect 13760 -12606 13832 -12602
rect 15798 -12550 15870 -12546
rect 15798 -12602 15808 -12550
rect 15860 -12602 15870 -12550
rect 15798 -12606 15870 -12602
rect 17830 -12550 17902 -12546
rect 17830 -12602 17840 -12550
rect 17892 -12602 17902 -12550
rect 17830 -12606 17902 -12602
rect 19868 -12550 19940 -12546
rect 19868 -12602 19878 -12550
rect 19930 -12602 19940 -12550
rect 19868 -12606 19940 -12602
rect 12218 -12660 12278 -12652
rect 12218 -12720 14326 -12660
rect 11726 -12762 11798 -12758
rect 9190 -12838 10260 -12778
rect 11726 -12814 11736 -12762
rect 11788 -12814 11798 -12762
rect 11726 -12818 11798 -12814
rect 9190 -12874 9250 -12838
rect 4900 -12880 5388 -12874
rect 4900 -12914 4947 -12880
rect 4981 -12914 5019 -12880
rect 5053 -12914 5091 -12880
rect 5125 -12914 5163 -12880
rect 5197 -12914 5235 -12880
rect 5269 -12914 5307 -12880
rect 5341 -12914 5388 -12880
rect 4900 -12920 5388 -12914
rect 5918 -12880 6406 -12874
rect 5918 -12914 5965 -12880
rect 5999 -12914 6037 -12880
rect 6071 -12914 6109 -12880
rect 6143 -12914 6181 -12880
rect 6215 -12914 6253 -12880
rect 6287 -12914 6325 -12880
rect 6359 -12914 6406 -12880
rect 5918 -12920 6406 -12914
rect 6936 -12880 7424 -12874
rect 6936 -12914 6983 -12880
rect 7017 -12914 7055 -12880
rect 7089 -12914 7127 -12880
rect 7161 -12914 7199 -12880
rect 7233 -12914 7271 -12880
rect 7305 -12914 7343 -12880
rect 7377 -12914 7424 -12880
rect 6936 -12920 7424 -12914
rect 7954 -12880 8162 -12874
rect 8222 -12880 8442 -12874
rect 7954 -12914 8001 -12880
rect 8035 -12914 8073 -12880
rect 8107 -12914 8145 -12880
rect 8179 -12914 8217 -12880
rect 8251 -12914 8289 -12880
rect 8323 -12914 8361 -12880
rect 8395 -12914 8442 -12880
rect 7954 -12920 8442 -12914
rect 8972 -12880 9460 -12874
rect 8972 -12914 9019 -12880
rect 9053 -12914 9091 -12880
rect 9125 -12914 9163 -12880
rect 9197 -12914 9235 -12880
rect 9269 -12914 9307 -12880
rect 9341 -12914 9379 -12880
rect 9413 -12914 9460 -12880
rect 8972 -12920 9460 -12914
rect 4604 -12996 4618 -12983
rect 3634 -13017 3640 -13012
rect 3594 -13055 3640 -13017
rect 3594 -13089 3600 -13055
rect 3634 -13089 3640 -13055
rect 3594 -13127 3640 -13089
rect 3594 -13161 3600 -13127
rect 3634 -13161 3640 -13127
rect 3594 -13199 3640 -13161
rect 3594 -13233 3600 -13199
rect 3634 -13233 3640 -13199
rect 3594 -13271 3640 -13233
rect 3594 -13305 3600 -13271
rect 3634 -13305 3640 -13271
rect 3594 -13343 3640 -13305
rect 3594 -13377 3600 -13343
rect 3634 -13377 3640 -13343
rect 3594 -13415 3640 -13377
rect 3594 -13449 3600 -13415
rect 3634 -13449 3640 -13415
rect 3594 -13487 3640 -13449
rect 3594 -13521 3600 -13487
rect 3634 -13521 3640 -13487
rect 3594 -13552 3640 -13521
rect 4612 -13017 4618 -12996
rect 4652 -12996 4664 -12983
rect 5630 -12983 5676 -12952
rect 4652 -13017 4658 -12996
rect 4612 -13055 4658 -13017
rect 4612 -13089 4618 -13055
rect 4652 -13089 4658 -13055
rect 4612 -13127 4658 -13089
rect 4612 -13161 4618 -13127
rect 4652 -13161 4658 -13127
rect 4612 -13199 4658 -13161
rect 4612 -13233 4618 -13199
rect 4652 -13233 4658 -13199
rect 4612 -13271 4658 -13233
rect 4612 -13305 4618 -13271
rect 4652 -13305 4658 -13271
rect 4612 -13343 4658 -13305
rect 4612 -13377 4618 -13343
rect 4652 -13377 4658 -13343
rect 4612 -13415 4658 -13377
rect 4612 -13449 4618 -13415
rect 4652 -13449 4658 -13415
rect 4612 -13487 4658 -13449
rect 4612 -13521 4618 -13487
rect 4652 -13521 4658 -13487
rect 5630 -13017 5636 -12983
rect 5670 -13017 5676 -12983
rect 5630 -13055 5676 -13017
rect 5630 -13089 5636 -13055
rect 5670 -13089 5676 -13055
rect 5630 -13127 5676 -13089
rect 5630 -13161 5636 -13127
rect 5670 -13161 5676 -13127
rect 5630 -13199 5676 -13161
rect 5630 -13233 5636 -13199
rect 5670 -13233 5676 -13199
rect 5630 -13271 5676 -13233
rect 5630 -13305 5636 -13271
rect 5670 -13305 5676 -13271
rect 5630 -13343 5676 -13305
rect 5630 -13377 5636 -13343
rect 5670 -13377 5676 -13343
rect 5630 -13415 5676 -13377
rect 5630 -13449 5636 -13415
rect 5670 -13449 5676 -13415
rect 5630 -13487 5676 -13449
rect 5630 -13512 5636 -13487
rect 4612 -13552 4658 -13521
rect 5624 -13521 5636 -13512
rect 5670 -13512 5676 -13487
rect 6648 -12983 6694 -12952
rect 6648 -13017 6654 -12983
rect 6688 -13017 6694 -12983
rect 7656 -12983 7716 -12964
rect 7656 -12998 7672 -12983
rect 6648 -13055 6694 -13017
rect 6648 -13089 6654 -13055
rect 6688 -13089 6694 -13055
rect 6648 -13127 6694 -13089
rect 6648 -13161 6654 -13127
rect 6688 -13161 6694 -13127
rect 6648 -13199 6694 -13161
rect 6648 -13233 6654 -13199
rect 6688 -13233 6694 -13199
rect 6648 -13271 6694 -13233
rect 6648 -13305 6654 -13271
rect 6688 -13305 6694 -13271
rect 6648 -13343 6694 -13305
rect 6648 -13377 6654 -13343
rect 6688 -13377 6694 -13343
rect 6648 -13415 6694 -13377
rect 6648 -13449 6654 -13415
rect 6688 -13449 6694 -13415
rect 6648 -13487 6694 -13449
rect 7666 -13017 7672 -12998
rect 7706 -12998 7716 -12983
rect 8684 -12983 8730 -12952
rect 7706 -13017 7712 -12998
rect 7666 -13055 7712 -13017
rect 7666 -13089 7672 -13055
rect 7706 -13089 7712 -13055
rect 7666 -13127 7712 -13089
rect 7666 -13161 7672 -13127
rect 7706 -13161 7712 -13127
rect 7666 -13199 7712 -13161
rect 7666 -13233 7672 -13199
rect 7706 -13233 7712 -13199
rect 7666 -13271 7712 -13233
rect 7666 -13305 7672 -13271
rect 7706 -13305 7712 -13271
rect 7666 -13343 7712 -13305
rect 7666 -13377 7672 -13343
rect 7706 -13377 7712 -13343
rect 7666 -13415 7712 -13377
rect 7666 -13449 7672 -13415
rect 7706 -13449 7712 -13415
rect 7666 -13464 7712 -13449
rect 8684 -13017 8690 -12983
rect 8724 -13017 8730 -12983
rect 9696 -12983 9756 -12838
rect 10200 -12874 10260 -12838
rect 9990 -12880 10478 -12874
rect 9990 -12914 10037 -12880
rect 10071 -12914 10109 -12880
rect 10143 -12914 10181 -12880
rect 10215 -12914 10253 -12880
rect 10287 -12914 10325 -12880
rect 10359 -12914 10397 -12880
rect 10431 -12914 10478 -12880
rect 9990 -12920 10478 -12914
rect 11008 -12880 11496 -12874
rect 11008 -12914 11055 -12880
rect 11089 -12914 11127 -12880
rect 11161 -12914 11199 -12880
rect 11233 -12914 11271 -12880
rect 11305 -12914 11343 -12880
rect 11377 -12914 11415 -12880
rect 11449 -12914 11496 -12880
rect 11008 -12920 11496 -12914
rect 9696 -13014 9708 -12983
rect 8684 -13055 8730 -13017
rect 8684 -13089 8690 -13055
rect 8724 -13089 8730 -13055
rect 8684 -13127 8730 -13089
rect 8684 -13161 8690 -13127
rect 8724 -13161 8730 -13127
rect 8684 -13199 8730 -13161
rect 8684 -13233 8690 -13199
rect 8724 -13233 8730 -13199
rect 8684 -13271 8730 -13233
rect 8684 -13305 8690 -13271
rect 8724 -13305 8730 -13271
rect 8684 -13343 8730 -13305
rect 8684 -13377 8690 -13343
rect 8724 -13377 8730 -13343
rect 8684 -13415 8730 -13377
rect 8684 -13449 8690 -13415
rect 8724 -13449 8730 -13415
rect 6648 -13492 6654 -13487
rect 5670 -13521 5684 -13512
rect 2864 -13590 3352 -13584
rect 2864 -13624 2911 -13590
rect 2945 -13624 2983 -13590
rect 3017 -13624 3055 -13590
rect 3089 -13624 3127 -13590
rect 3161 -13624 3199 -13590
rect 3233 -13624 3271 -13590
rect 3305 -13624 3352 -13590
rect 2864 -13630 3352 -13624
rect 3882 -13590 4370 -13584
rect 3882 -13624 3929 -13590
rect 3963 -13624 4001 -13590
rect 4035 -13624 4073 -13590
rect 4107 -13624 4145 -13590
rect 4179 -13624 4217 -13590
rect 4251 -13624 4289 -13590
rect 4323 -13624 4370 -13590
rect 3882 -13630 4370 -13624
rect 4900 -13590 5388 -13584
rect 4900 -13624 4947 -13590
rect 4981 -13624 5019 -13590
rect 5053 -13624 5091 -13590
rect 5125 -13624 5163 -13590
rect 5197 -13624 5235 -13590
rect 5269 -13624 5307 -13590
rect 5341 -13624 5388 -13590
rect 4900 -13630 5388 -13624
rect 5624 -13682 5684 -13521
rect 6642 -13521 6654 -13492
rect 6688 -13492 6694 -13487
rect 7656 -13480 7716 -13464
rect 7656 -13487 7720 -13480
rect 8684 -13484 8730 -13449
rect 9702 -13017 9708 -13014
rect 9742 -13014 9756 -12983
rect 10720 -12983 10766 -12952
rect 9742 -13017 9748 -13014
rect 9702 -13055 9748 -13017
rect 9702 -13089 9708 -13055
rect 9742 -13089 9748 -13055
rect 9702 -13127 9748 -13089
rect 9702 -13161 9708 -13127
rect 9742 -13161 9748 -13127
rect 9702 -13199 9748 -13161
rect 9702 -13233 9708 -13199
rect 9742 -13233 9748 -13199
rect 9702 -13271 9748 -13233
rect 9702 -13305 9708 -13271
rect 9742 -13305 9748 -13271
rect 9702 -13343 9748 -13305
rect 9702 -13377 9708 -13343
rect 9742 -13377 9748 -13343
rect 9702 -13415 9748 -13377
rect 9702 -13449 9708 -13415
rect 9742 -13449 9748 -13415
rect 6688 -13521 6702 -13492
rect 5918 -13590 6406 -13584
rect 5918 -13624 5965 -13590
rect 5999 -13624 6037 -13590
rect 6071 -13624 6109 -13590
rect 6143 -13624 6181 -13590
rect 6215 -13624 6253 -13590
rect 6287 -13624 6325 -13590
rect 6359 -13624 6406 -13590
rect 5918 -13630 6406 -13624
rect 6272 -13678 6332 -13630
rect 6642 -13678 6702 -13521
rect 7656 -13521 7672 -13487
rect 7706 -13521 7720 -13487
rect 7656 -13540 7720 -13521
rect 8676 -13487 8736 -13484
rect 8676 -13521 8690 -13487
rect 8724 -13521 8736 -13487
rect 9702 -13487 9748 -13449
rect 10720 -13017 10726 -12983
rect 10760 -13017 10766 -12983
rect 11732 -12983 11792 -12818
rect 12218 -12874 12278 -12720
rect 13252 -12874 13312 -12720
rect 13758 -12762 13830 -12758
rect 13758 -12814 13768 -12762
rect 13820 -12814 13830 -12762
rect 13758 -12818 13830 -12814
rect 12026 -12880 12514 -12874
rect 12026 -12914 12073 -12880
rect 12107 -12914 12145 -12880
rect 12179 -12914 12217 -12880
rect 12251 -12914 12289 -12880
rect 12323 -12914 12361 -12880
rect 12395 -12914 12433 -12880
rect 12467 -12914 12514 -12880
rect 12026 -12920 12514 -12914
rect 13044 -12880 13532 -12874
rect 13044 -12914 13091 -12880
rect 13125 -12914 13163 -12880
rect 13197 -12914 13235 -12880
rect 13269 -12914 13307 -12880
rect 13341 -12914 13379 -12880
rect 13413 -12914 13451 -12880
rect 13485 -12914 13532 -12880
rect 13044 -12920 13532 -12914
rect 11732 -12998 11744 -12983
rect 10720 -13055 10766 -13017
rect 10720 -13089 10726 -13055
rect 10760 -13089 10766 -13055
rect 10720 -13127 10766 -13089
rect 10720 -13161 10726 -13127
rect 10760 -13161 10766 -13127
rect 10720 -13199 10766 -13161
rect 10720 -13233 10726 -13199
rect 10760 -13233 10766 -13199
rect 10720 -13271 10766 -13233
rect 10720 -13305 10726 -13271
rect 10760 -13305 10766 -13271
rect 10720 -13343 10766 -13305
rect 10720 -13377 10726 -13343
rect 10760 -13377 10766 -13343
rect 10720 -13415 10766 -13377
rect 10720 -13449 10726 -13415
rect 10760 -13449 10766 -13415
rect 10720 -13464 10766 -13449
rect 11738 -13017 11744 -12998
rect 11778 -12998 11792 -12983
rect 12756 -12983 12802 -12952
rect 11778 -13017 11784 -12998
rect 11738 -13055 11784 -13017
rect 11738 -13089 11744 -13055
rect 11778 -13089 11784 -13055
rect 11738 -13127 11784 -13089
rect 11738 -13161 11744 -13127
rect 11778 -13161 11784 -13127
rect 11738 -13199 11784 -13161
rect 11738 -13233 11744 -13199
rect 11778 -13233 11784 -13199
rect 11738 -13271 11784 -13233
rect 11738 -13305 11744 -13271
rect 11778 -13305 11784 -13271
rect 11738 -13343 11784 -13305
rect 11738 -13377 11744 -13343
rect 11778 -13377 11784 -13343
rect 11738 -13415 11784 -13377
rect 11738 -13449 11744 -13415
rect 11778 -13449 11784 -13415
rect 9702 -13490 9708 -13487
rect 9696 -13504 9708 -13490
rect 6936 -13590 7424 -13584
rect 6936 -13624 6983 -13590
rect 7017 -13624 7055 -13590
rect 7089 -13624 7127 -13590
rect 7161 -13624 7199 -13590
rect 7233 -13624 7271 -13590
rect 7305 -13624 7343 -13590
rect 7377 -13624 7424 -13590
rect 6936 -13630 7424 -13624
rect 7144 -13678 7204 -13630
rect 7656 -13678 7716 -13540
rect 7954 -13590 8442 -13584
rect 7954 -13624 8001 -13590
rect 8035 -13624 8073 -13590
rect 8107 -13624 8145 -13590
rect 8179 -13624 8217 -13590
rect 8251 -13624 8289 -13590
rect 8323 -13624 8361 -13590
rect 8395 -13624 8442 -13590
rect 7954 -13630 8442 -13624
rect 8184 -13678 8244 -13630
rect 8676 -13678 8736 -13521
rect 9694 -13521 9708 -13504
rect 9742 -13490 9748 -13487
rect 10708 -13487 10768 -13464
rect 11738 -13478 11784 -13449
rect 12756 -13017 12762 -12983
rect 12796 -13017 12802 -12983
rect 13764 -12983 13824 -12818
rect 14266 -12874 14326 -12720
rect 15290 -12808 16372 -12748
rect 15290 -12874 15350 -12808
rect 14062 -12880 14550 -12874
rect 14062 -12914 14109 -12880
rect 14143 -12914 14181 -12880
rect 14215 -12914 14253 -12880
rect 14287 -12914 14325 -12880
rect 14359 -12914 14397 -12880
rect 14431 -12914 14469 -12880
rect 14503 -12914 14550 -12880
rect 14062 -12920 14550 -12914
rect 15080 -12880 15568 -12874
rect 15080 -12914 15127 -12880
rect 15161 -12914 15199 -12880
rect 15233 -12914 15271 -12880
rect 15305 -12914 15343 -12880
rect 15377 -12914 15415 -12880
rect 15449 -12914 15487 -12880
rect 15521 -12914 15568 -12880
rect 15080 -12920 15568 -12914
rect 13764 -12998 13780 -12983
rect 12756 -13055 12802 -13017
rect 12756 -13089 12762 -13055
rect 12796 -13089 12802 -13055
rect 12756 -13127 12802 -13089
rect 12756 -13161 12762 -13127
rect 12796 -13161 12802 -13127
rect 12756 -13199 12802 -13161
rect 12756 -13233 12762 -13199
rect 12796 -13233 12802 -13199
rect 12756 -13271 12802 -13233
rect 12756 -13305 12762 -13271
rect 12796 -13305 12802 -13271
rect 12756 -13343 12802 -13305
rect 12756 -13377 12762 -13343
rect 12796 -13377 12802 -13343
rect 12756 -13415 12802 -13377
rect 12756 -13449 12762 -13415
rect 12796 -13449 12802 -13415
rect 12756 -13474 12802 -13449
rect 13774 -13017 13780 -12998
rect 13814 -12998 13824 -12983
rect 14792 -12983 14838 -12952
rect 13814 -13017 13820 -12998
rect 13774 -13055 13820 -13017
rect 13774 -13089 13780 -13055
rect 13814 -13089 13820 -13055
rect 13774 -13127 13820 -13089
rect 13774 -13161 13780 -13127
rect 13814 -13161 13820 -13127
rect 13774 -13199 13820 -13161
rect 13774 -13233 13780 -13199
rect 13814 -13233 13820 -13199
rect 13774 -13271 13820 -13233
rect 13774 -13305 13780 -13271
rect 13814 -13305 13820 -13271
rect 13774 -13343 13820 -13305
rect 13774 -13377 13780 -13343
rect 13814 -13377 13820 -13343
rect 13774 -13415 13820 -13377
rect 13774 -13449 13780 -13415
rect 13814 -13449 13820 -13415
rect 11732 -13482 11792 -13478
rect 9742 -13521 9756 -13490
rect 9694 -13540 9756 -13521
rect 10708 -13521 10726 -13487
rect 10760 -13521 10768 -13487
rect 8972 -13590 9460 -13584
rect 8972 -13624 9019 -13590
rect 9053 -13624 9091 -13590
rect 9125 -13624 9163 -13590
rect 9197 -13624 9235 -13590
rect 9269 -13624 9307 -13590
rect 9341 -13624 9379 -13590
rect 9413 -13624 9460 -13590
rect 8972 -13630 9460 -13624
rect 6266 -13682 6338 -13678
rect 5624 -13742 6196 -13682
rect 6266 -13734 6276 -13682
rect 6328 -13734 6338 -13682
rect 6266 -13738 6338 -13734
rect 6636 -13682 6708 -13678
rect 6636 -13734 6646 -13682
rect 6698 -13734 6708 -13682
rect 6636 -13738 6708 -13734
rect 7138 -13682 7210 -13678
rect 7138 -13734 7148 -13682
rect 7200 -13734 7210 -13682
rect 7138 -13738 7210 -13734
rect 7650 -13682 7722 -13678
rect 7650 -13734 7660 -13682
rect 7712 -13734 7722 -13682
rect 7650 -13738 7722 -13734
rect 8178 -13682 8250 -13678
rect 8178 -13734 8188 -13682
rect 8240 -13734 8250 -13682
rect 8178 -13738 8250 -13734
rect 8670 -13682 8742 -13678
rect 8670 -13734 8680 -13682
rect 8732 -13734 8742 -13682
rect 8670 -13738 8742 -13734
rect 4090 -13792 4162 -13788
rect 4090 -13844 4100 -13792
rect 4152 -13844 4162 -13792
rect 4090 -13848 4162 -13844
rect 5112 -13792 5184 -13788
rect 5112 -13844 5122 -13792
rect 5174 -13844 5184 -13792
rect 5112 -13848 5184 -13844
rect 2566 -14004 2638 -14000
rect 2566 -14056 2576 -14004
rect 2628 -14056 2638 -14004
rect 2566 -14060 2638 -14056
rect 3064 -14004 3136 -14000
rect 3064 -14056 3074 -14004
rect 3126 -14056 3136 -14004
rect 3064 -14060 3136 -14056
rect 3576 -14004 3648 -14000
rect 3576 -14056 3586 -14004
rect 3638 -14056 3648 -14004
rect 3576 -14060 3648 -14056
rect 2572 -14215 2632 -14060
rect 3070 -14106 3130 -14060
rect 2864 -14112 3352 -14106
rect 2864 -14146 2911 -14112
rect 2945 -14146 2983 -14112
rect 3017 -14146 3055 -14112
rect 3089 -14146 3127 -14112
rect 3161 -14146 3199 -14112
rect 3233 -14146 3271 -14112
rect 3305 -14146 3352 -14112
rect 2864 -14152 3352 -14146
rect 2572 -14236 2582 -14215
rect 2576 -14249 2582 -14236
rect 2616 -14236 2632 -14215
rect 3582 -14215 3642 -14060
rect 4096 -14106 4156 -13848
rect 5118 -14106 5178 -13848
rect 6136 -13886 6196 -13742
rect 6136 -13896 6198 -13886
rect 6136 -13948 6142 -13896
rect 6194 -13948 6198 -13896
rect 6136 -13958 6198 -13948
rect 5618 -14004 5690 -14000
rect 5618 -14056 5628 -14004
rect 5680 -14056 5690 -14004
rect 5618 -14060 5690 -14056
rect 3882 -14112 4370 -14106
rect 3882 -14146 3929 -14112
rect 3963 -14146 4001 -14112
rect 4035 -14146 4073 -14112
rect 4107 -14146 4145 -14112
rect 4179 -14146 4217 -14112
rect 4251 -14146 4289 -14112
rect 4323 -14146 4370 -14112
rect 3882 -14152 4370 -14146
rect 4900 -14112 5388 -14106
rect 4900 -14146 4947 -14112
rect 4981 -14146 5019 -14112
rect 5053 -14146 5091 -14112
rect 5125 -14146 5163 -14112
rect 5197 -14146 5235 -14112
rect 5269 -14146 5307 -14112
rect 5341 -14146 5388 -14112
rect 4900 -14152 5388 -14146
rect 2616 -14249 2622 -14236
rect 3582 -14242 3600 -14215
rect 2576 -14287 2622 -14249
rect 2576 -14321 2582 -14287
rect 2616 -14321 2622 -14287
rect 2576 -14359 2622 -14321
rect 2576 -14393 2582 -14359
rect 2616 -14393 2622 -14359
rect 2576 -14431 2622 -14393
rect 2576 -14465 2582 -14431
rect 2616 -14465 2622 -14431
rect 2576 -14503 2622 -14465
rect 2576 -14537 2582 -14503
rect 2616 -14537 2622 -14503
rect 2576 -14575 2622 -14537
rect 2576 -14609 2582 -14575
rect 2616 -14609 2622 -14575
rect 2576 -14647 2622 -14609
rect 2576 -14681 2582 -14647
rect 2616 -14681 2622 -14647
rect 2576 -14719 2622 -14681
rect 2576 -14753 2582 -14719
rect 2616 -14753 2622 -14719
rect 2576 -14784 2622 -14753
rect 3594 -14249 3600 -14242
rect 3634 -14242 3642 -14215
rect 4612 -14215 4658 -14184
rect 3634 -14249 3640 -14242
rect 3594 -14287 3640 -14249
rect 3594 -14321 3600 -14287
rect 3634 -14321 3640 -14287
rect 3594 -14359 3640 -14321
rect 3594 -14393 3600 -14359
rect 3634 -14393 3640 -14359
rect 3594 -14431 3640 -14393
rect 3594 -14465 3600 -14431
rect 3634 -14465 3640 -14431
rect 3594 -14503 3640 -14465
rect 3594 -14537 3600 -14503
rect 3634 -14537 3640 -14503
rect 3594 -14575 3640 -14537
rect 3594 -14609 3600 -14575
rect 3634 -14609 3640 -14575
rect 3594 -14647 3640 -14609
rect 3594 -14681 3600 -14647
rect 3634 -14681 3640 -14647
rect 3594 -14719 3640 -14681
rect 4612 -14249 4618 -14215
rect 4652 -14249 4658 -14215
rect 5624 -14215 5684 -14060
rect 6136 -14106 6196 -13958
rect 5918 -14112 6406 -14106
rect 5918 -14146 5965 -14112
rect 5999 -14146 6037 -14112
rect 6071 -14146 6109 -14112
rect 6143 -14146 6181 -14112
rect 6215 -14146 6253 -14112
rect 6287 -14146 6325 -14112
rect 6359 -14146 6406 -14112
rect 5918 -14152 6406 -14146
rect 5624 -14248 5636 -14215
rect 4612 -14287 4658 -14249
rect 4612 -14321 4618 -14287
rect 4652 -14321 4658 -14287
rect 4612 -14359 4658 -14321
rect 4612 -14393 4618 -14359
rect 4652 -14393 4658 -14359
rect 4612 -14431 4658 -14393
rect 4612 -14465 4618 -14431
rect 4652 -14465 4658 -14431
rect 4612 -14503 4658 -14465
rect 4612 -14537 4618 -14503
rect 4652 -14537 4658 -14503
rect 4612 -14575 4658 -14537
rect 4612 -14609 4618 -14575
rect 4652 -14609 4658 -14575
rect 4612 -14647 4658 -14609
rect 4612 -14681 4618 -14647
rect 4652 -14681 4658 -14647
rect 4612 -14714 4658 -14681
rect 3594 -14753 3600 -14719
rect 3634 -14753 3640 -14719
rect 3594 -14784 3640 -14753
rect 4598 -14719 4658 -14714
rect 4598 -14753 4618 -14719
rect 4652 -14753 4658 -14719
rect 2864 -14822 3352 -14816
rect 2864 -14856 2911 -14822
rect 2945 -14856 2983 -14822
rect 3017 -14856 3055 -14822
rect 3089 -14856 3127 -14822
rect 3161 -14856 3199 -14822
rect 3233 -14856 3271 -14822
rect 3305 -14856 3352 -14822
rect 2864 -14862 3352 -14856
rect 3882 -14822 4370 -14816
rect 3882 -14856 3929 -14822
rect 3963 -14856 4001 -14822
rect 4035 -14856 4073 -14822
rect 4107 -14856 4145 -14822
rect 4179 -14856 4217 -14822
rect 4251 -14856 4289 -14822
rect 4323 -14856 4370 -14822
rect 3882 -14862 4370 -14856
rect 4080 -14906 4152 -14902
rect 4080 -14958 4090 -14906
rect 4142 -14958 4152 -14906
rect 4080 -14962 4152 -14958
rect 2330 -15120 2402 -15116
rect 2330 -15172 2340 -15120
rect 2392 -15172 2402 -15120
rect 2330 -15176 2402 -15172
rect 2336 -16358 2396 -15176
rect 2568 -15272 3646 -15212
rect 2568 -15449 2628 -15272
rect 3076 -15340 3136 -15272
rect 2862 -15346 3350 -15340
rect 2862 -15380 2909 -15346
rect 2943 -15380 2981 -15346
rect 3015 -15380 3053 -15346
rect 3087 -15380 3125 -15346
rect 3159 -15380 3197 -15346
rect 3231 -15380 3269 -15346
rect 3303 -15380 3350 -15346
rect 2862 -15386 3350 -15380
rect 2568 -15456 2580 -15449
rect 2574 -15483 2580 -15456
rect 2614 -15456 2628 -15449
rect 3586 -15449 3646 -15272
rect 4086 -15340 4146 -14962
rect 4598 -14994 4658 -14753
rect 5630 -14249 5636 -14248
rect 5670 -14248 5684 -14215
rect 6642 -14215 6702 -13738
rect 7132 -13896 7204 -13892
rect 7132 -13948 7142 -13896
rect 7194 -13948 7204 -13896
rect 7132 -13952 7204 -13948
rect 8152 -13896 8224 -13892
rect 8152 -13948 8162 -13896
rect 8214 -13948 8224 -13896
rect 8152 -13952 8224 -13948
rect 7138 -14106 7198 -13952
rect 7652 -14004 7724 -14000
rect 7652 -14056 7662 -14004
rect 7714 -14056 7724 -14004
rect 7652 -14060 7724 -14056
rect 6936 -14112 7424 -14106
rect 6936 -14146 6983 -14112
rect 7017 -14146 7055 -14112
rect 7089 -14146 7127 -14112
rect 7161 -14146 7199 -14112
rect 7233 -14146 7271 -14112
rect 7305 -14146 7343 -14112
rect 7377 -14146 7424 -14112
rect 6936 -14152 7424 -14146
rect 5670 -14249 5676 -14248
rect 5630 -14287 5676 -14249
rect 6642 -14249 6654 -14215
rect 6688 -14249 6702 -14215
rect 7658 -14215 7718 -14060
rect 8158 -14106 8218 -13952
rect 7954 -14112 8442 -14106
rect 7954 -14146 8001 -14112
rect 8035 -14146 8073 -14112
rect 8107 -14146 8145 -14112
rect 8179 -14146 8217 -14112
rect 8251 -14146 8289 -14112
rect 8323 -14146 8361 -14112
rect 8395 -14146 8442 -14112
rect 7954 -14152 8442 -14146
rect 7658 -14230 7672 -14215
rect 6642 -14260 6702 -14249
rect 7666 -14249 7672 -14230
rect 7706 -14230 7718 -14215
rect 8676 -14215 8736 -13738
rect 9190 -13788 9250 -13630
rect 9694 -13788 9754 -13540
rect 9990 -13590 10478 -13584
rect 9990 -13624 10037 -13590
rect 10071 -13624 10109 -13590
rect 10143 -13624 10181 -13590
rect 10215 -13624 10253 -13590
rect 10287 -13624 10325 -13590
rect 10359 -13624 10397 -13590
rect 10431 -13624 10478 -13590
rect 9990 -13630 10478 -13624
rect 10210 -13788 10270 -13630
rect 10708 -13678 10768 -13521
rect 11730 -13487 11792 -13482
rect 11730 -13521 11744 -13487
rect 11778 -13521 11792 -13487
rect 11730 -13540 11792 -13521
rect 12744 -13487 12804 -13474
rect 12744 -13521 12762 -13487
rect 12796 -13521 12804 -13487
rect 13774 -13487 13820 -13449
rect 14792 -13017 14798 -12983
rect 14832 -13017 14838 -12983
rect 15802 -12983 15862 -12808
rect 16312 -12874 16372 -12808
rect 17328 -12808 17900 -12748
rect 17328 -12874 17388 -12808
rect 16098 -12880 16586 -12874
rect 16098 -12914 16145 -12880
rect 16179 -12914 16217 -12880
rect 16251 -12914 16289 -12880
rect 16323 -12914 16361 -12880
rect 16395 -12914 16433 -12880
rect 16467 -12914 16505 -12880
rect 16539 -12914 16586 -12880
rect 16098 -12920 16586 -12914
rect 17116 -12880 17604 -12874
rect 17116 -12914 17163 -12880
rect 17197 -12914 17235 -12880
rect 17269 -12914 17307 -12880
rect 17341 -12914 17379 -12880
rect 17413 -12914 17451 -12880
rect 17485 -12914 17523 -12880
rect 17557 -12914 17604 -12880
rect 17116 -12920 17604 -12914
rect 15802 -13004 15816 -12983
rect 14792 -13055 14838 -13017
rect 14792 -13089 14798 -13055
rect 14832 -13089 14838 -13055
rect 14792 -13127 14838 -13089
rect 14792 -13161 14798 -13127
rect 14832 -13161 14838 -13127
rect 14792 -13199 14838 -13161
rect 14792 -13233 14798 -13199
rect 14832 -13233 14838 -13199
rect 14792 -13271 14838 -13233
rect 14792 -13305 14798 -13271
rect 14832 -13305 14838 -13271
rect 14792 -13343 14838 -13305
rect 14792 -13377 14798 -13343
rect 14832 -13377 14838 -13343
rect 14792 -13415 14838 -13377
rect 14792 -13449 14798 -13415
rect 14832 -13449 14838 -13415
rect 14792 -13480 14838 -13449
rect 15810 -13017 15816 -13004
rect 15850 -13004 15862 -12983
rect 16828 -12983 16874 -12952
rect 15850 -13017 15856 -13004
rect 15810 -13055 15856 -13017
rect 15810 -13089 15816 -13055
rect 15850 -13089 15856 -13055
rect 15810 -13127 15856 -13089
rect 15810 -13161 15816 -13127
rect 15850 -13161 15856 -13127
rect 15810 -13199 15856 -13161
rect 15810 -13233 15816 -13199
rect 15850 -13233 15856 -13199
rect 15810 -13271 15856 -13233
rect 15810 -13305 15816 -13271
rect 15850 -13305 15856 -13271
rect 15810 -13343 15856 -13305
rect 15810 -13377 15816 -13343
rect 15850 -13377 15856 -13343
rect 15810 -13415 15856 -13377
rect 15810 -13449 15816 -13415
rect 15850 -13449 15856 -13415
rect 15810 -13474 15856 -13449
rect 16828 -13017 16834 -12983
rect 16868 -13017 16874 -12983
rect 17840 -12983 17900 -12808
rect 18134 -12880 18622 -12874
rect 18134 -12914 18181 -12880
rect 18215 -12914 18253 -12880
rect 18287 -12914 18325 -12880
rect 18359 -12914 18397 -12880
rect 18431 -12914 18469 -12880
rect 18503 -12914 18541 -12880
rect 18575 -12914 18622 -12880
rect 18134 -12920 18622 -12914
rect 19152 -12880 19640 -12874
rect 19152 -12914 19199 -12880
rect 19233 -12914 19271 -12880
rect 19305 -12914 19343 -12880
rect 19377 -12914 19415 -12880
rect 19449 -12914 19487 -12880
rect 19521 -12914 19559 -12880
rect 19593 -12914 19640 -12880
rect 19152 -12920 19640 -12914
rect 17840 -12990 17852 -12983
rect 16828 -13055 16874 -13017
rect 16828 -13089 16834 -13055
rect 16868 -13089 16874 -13055
rect 16828 -13127 16874 -13089
rect 16828 -13161 16834 -13127
rect 16868 -13161 16874 -13127
rect 16828 -13199 16874 -13161
rect 16828 -13233 16834 -13199
rect 16868 -13233 16874 -13199
rect 16828 -13271 16874 -13233
rect 16828 -13305 16834 -13271
rect 16868 -13305 16874 -13271
rect 16828 -13343 16874 -13305
rect 16828 -13377 16834 -13343
rect 16868 -13377 16874 -13343
rect 16828 -13415 16874 -13377
rect 16828 -13449 16834 -13415
rect 16868 -13449 16874 -13415
rect 13774 -13514 13780 -13487
rect 11008 -13590 11496 -13584
rect 11008 -13624 11055 -13590
rect 11089 -13624 11127 -13590
rect 11161 -13624 11199 -13590
rect 11233 -13624 11271 -13590
rect 11305 -13624 11343 -13590
rect 11377 -13624 11415 -13590
rect 11449 -13624 11496 -13590
rect 11008 -13630 11496 -13624
rect 10702 -13682 10774 -13678
rect 10702 -13734 10712 -13682
rect 10764 -13734 10774 -13682
rect 10702 -13738 10774 -13734
rect 9184 -13792 9256 -13788
rect 9184 -13844 9194 -13792
rect 9246 -13844 9256 -13792
rect 9184 -13848 9256 -13844
rect 9688 -13792 9760 -13788
rect 9688 -13844 9698 -13792
rect 9750 -13844 9760 -13792
rect 9688 -13848 9760 -13844
rect 10204 -13792 10276 -13788
rect 10204 -13844 10214 -13792
rect 10266 -13844 10276 -13792
rect 10204 -13848 10276 -13844
rect 9190 -14106 9250 -13848
rect 9686 -14004 9758 -14000
rect 9686 -14056 9696 -14004
rect 9748 -14056 9758 -14004
rect 9686 -14060 9758 -14056
rect 8972 -14112 9460 -14106
rect 8972 -14146 9019 -14112
rect 9053 -14146 9091 -14112
rect 9125 -14146 9163 -14112
rect 9197 -14146 9235 -14112
rect 9269 -14146 9307 -14112
rect 9341 -14146 9379 -14112
rect 9413 -14146 9460 -14112
rect 8972 -14152 9460 -14146
rect 7706 -14249 7712 -14230
rect 8676 -14238 8690 -14215
rect 5630 -14321 5636 -14287
rect 5670 -14321 5676 -14287
rect 5630 -14359 5676 -14321
rect 5630 -14393 5636 -14359
rect 5670 -14393 5676 -14359
rect 5630 -14431 5676 -14393
rect 5630 -14465 5636 -14431
rect 5670 -14465 5676 -14431
rect 5630 -14503 5676 -14465
rect 5630 -14537 5636 -14503
rect 5670 -14537 5676 -14503
rect 5630 -14575 5676 -14537
rect 5630 -14609 5636 -14575
rect 5670 -14609 5676 -14575
rect 5630 -14647 5676 -14609
rect 5630 -14681 5636 -14647
rect 5670 -14681 5676 -14647
rect 5630 -14719 5676 -14681
rect 6648 -14287 6694 -14260
rect 6648 -14321 6654 -14287
rect 6688 -14321 6694 -14287
rect 6648 -14359 6694 -14321
rect 6648 -14393 6654 -14359
rect 6688 -14393 6694 -14359
rect 6648 -14431 6694 -14393
rect 6648 -14465 6654 -14431
rect 6688 -14465 6694 -14431
rect 6648 -14503 6694 -14465
rect 6648 -14537 6654 -14503
rect 6688 -14537 6694 -14503
rect 6648 -14575 6694 -14537
rect 6648 -14609 6654 -14575
rect 6688 -14609 6694 -14575
rect 6648 -14647 6694 -14609
rect 6648 -14681 6654 -14647
rect 6688 -14681 6694 -14647
rect 6648 -14708 6694 -14681
rect 5630 -14753 5636 -14719
rect 5670 -14753 5676 -14719
rect 5630 -14784 5676 -14753
rect 6634 -14719 6694 -14708
rect 6634 -14753 6654 -14719
rect 6688 -14753 6694 -14719
rect 4900 -14822 5388 -14816
rect 4900 -14856 4947 -14822
rect 4981 -14856 5019 -14822
rect 5053 -14856 5091 -14822
rect 5125 -14856 5163 -14822
rect 5197 -14856 5235 -14822
rect 5269 -14856 5307 -14822
rect 5341 -14856 5388 -14822
rect 4900 -14862 5388 -14856
rect 5918 -14822 6120 -14816
rect 6122 -14822 6406 -14816
rect 5918 -14856 5965 -14822
rect 5999 -14856 6037 -14822
rect 6071 -14856 6109 -14822
rect 6143 -14856 6181 -14822
rect 6215 -14856 6253 -14822
rect 6287 -14856 6325 -14822
rect 6359 -14856 6406 -14822
rect 5918 -14862 6120 -14856
rect 6122 -14862 6406 -14856
rect 6122 -14890 6182 -14862
rect 5096 -14894 5168 -14890
rect 5096 -14946 5106 -14894
rect 5158 -14946 5168 -14894
rect 5096 -14950 5168 -14946
rect 6116 -14894 6188 -14890
rect 6116 -14946 6126 -14894
rect 6178 -14946 6188 -14894
rect 6116 -14950 6188 -14946
rect 4592 -14998 4664 -14994
rect 4592 -15050 4602 -14998
rect 4654 -15050 4664 -14998
rect 4592 -15054 4664 -15050
rect 4598 -15232 4670 -15228
rect 4598 -15284 4608 -15232
rect 4660 -15284 4670 -15232
rect 4598 -15288 4670 -15284
rect 3880 -15346 4368 -15340
rect 3880 -15380 3927 -15346
rect 3961 -15380 3999 -15346
rect 4033 -15380 4071 -15346
rect 4105 -15380 4143 -15346
rect 4177 -15380 4215 -15346
rect 4249 -15380 4287 -15346
rect 4321 -15380 4368 -15346
rect 3880 -15386 4368 -15380
rect 2614 -15483 2620 -15456
rect 3586 -15462 3598 -15449
rect 2574 -15521 2620 -15483
rect 2574 -15555 2580 -15521
rect 2614 -15555 2620 -15521
rect 2574 -15593 2620 -15555
rect 2574 -15627 2580 -15593
rect 2614 -15627 2620 -15593
rect 2574 -15665 2620 -15627
rect 2574 -15699 2580 -15665
rect 2614 -15699 2620 -15665
rect 2574 -15737 2620 -15699
rect 2574 -15771 2580 -15737
rect 2614 -15771 2620 -15737
rect 2574 -15809 2620 -15771
rect 2574 -15843 2580 -15809
rect 2614 -15843 2620 -15809
rect 2574 -15881 2620 -15843
rect 2574 -15915 2580 -15881
rect 2614 -15915 2620 -15881
rect 2574 -15953 2620 -15915
rect 2574 -15987 2580 -15953
rect 2614 -15987 2620 -15953
rect 3592 -15483 3598 -15462
rect 3632 -15462 3646 -15449
rect 4604 -15449 4664 -15288
rect 5102 -15340 5162 -14950
rect 5616 -14998 5688 -14994
rect 5616 -15050 5626 -14998
rect 5678 -15050 5688 -14998
rect 5616 -15054 5688 -15050
rect 4898 -15346 5386 -15340
rect 4898 -15380 4945 -15346
rect 4979 -15380 5017 -15346
rect 5051 -15380 5089 -15346
rect 5123 -15380 5161 -15346
rect 5195 -15380 5233 -15346
rect 5267 -15380 5305 -15346
rect 5339 -15380 5386 -15346
rect 4898 -15386 5386 -15380
rect 4604 -15456 4616 -15449
rect 3632 -15483 3638 -15462
rect 3592 -15521 3638 -15483
rect 3592 -15555 3598 -15521
rect 3632 -15555 3638 -15521
rect 3592 -15593 3638 -15555
rect 3592 -15627 3598 -15593
rect 3632 -15627 3638 -15593
rect 3592 -15665 3638 -15627
rect 3592 -15699 3598 -15665
rect 3632 -15699 3638 -15665
rect 3592 -15737 3638 -15699
rect 3592 -15771 3598 -15737
rect 3632 -15771 3638 -15737
rect 3592 -15809 3638 -15771
rect 3592 -15843 3598 -15809
rect 3632 -15843 3638 -15809
rect 3592 -15881 3638 -15843
rect 3592 -15915 3598 -15881
rect 3632 -15915 3638 -15881
rect 3592 -15953 3638 -15915
rect 3592 -15962 3598 -15953
rect 2574 -16018 2620 -15987
rect 3586 -15987 3598 -15962
rect 3632 -15962 3638 -15953
rect 4610 -15483 4616 -15456
rect 4650 -15456 4664 -15449
rect 5622 -15449 5682 -15054
rect 6122 -15340 6182 -14950
rect 6634 -14994 6694 -14753
rect 7666 -14287 7712 -14249
rect 7666 -14321 7672 -14287
rect 7706 -14321 7712 -14287
rect 7666 -14359 7712 -14321
rect 7666 -14393 7672 -14359
rect 7706 -14393 7712 -14359
rect 7666 -14431 7712 -14393
rect 7666 -14465 7672 -14431
rect 7706 -14465 7712 -14431
rect 7666 -14503 7712 -14465
rect 7666 -14537 7672 -14503
rect 7706 -14537 7712 -14503
rect 7666 -14575 7712 -14537
rect 7666 -14609 7672 -14575
rect 7706 -14609 7712 -14575
rect 7666 -14647 7712 -14609
rect 7666 -14681 7672 -14647
rect 7706 -14681 7712 -14647
rect 7666 -14719 7712 -14681
rect 7666 -14753 7672 -14719
rect 7706 -14753 7712 -14719
rect 8684 -14249 8690 -14238
rect 8724 -14238 8736 -14215
rect 9692 -14215 9752 -14060
rect 10210 -14106 10270 -13848
rect 9990 -14112 10478 -14106
rect 9990 -14146 10037 -14112
rect 10071 -14146 10109 -14112
rect 10143 -14146 10181 -14112
rect 10215 -14146 10253 -14112
rect 10287 -14146 10325 -14112
rect 10359 -14146 10397 -14112
rect 10431 -14146 10478 -14112
rect 9990 -14152 10478 -14146
rect 8724 -14249 8730 -14238
rect 8684 -14287 8730 -14249
rect 9692 -14249 9708 -14215
rect 9742 -14249 9752 -14215
rect 9692 -14258 9752 -14249
rect 10708 -14215 10768 -13738
rect 11230 -13788 11290 -13630
rect 11730 -13676 11790 -13540
rect 12026 -13590 12514 -13584
rect 12026 -13624 12073 -13590
rect 12107 -13624 12145 -13590
rect 12179 -13624 12217 -13590
rect 12251 -13624 12289 -13590
rect 12323 -13624 12361 -13590
rect 12395 -13624 12433 -13590
rect 12467 -13624 12514 -13590
rect 12026 -13630 12514 -13624
rect 11730 -13736 11908 -13676
rect 11224 -13792 11296 -13788
rect 11224 -13844 11234 -13792
rect 11286 -13844 11296 -13792
rect 11224 -13848 11296 -13844
rect 11726 -13792 11798 -13788
rect 11726 -13844 11736 -13792
rect 11788 -13844 11798 -13792
rect 11726 -13848 11798 -13844
rect 11230 -14106 11290 -13848
rect 11008 -14112 11496 -14106
rect 11008 -14146 11055 -14112
rect 11089 -14146 11127 -14112
rect 11161 -14146 11199 -14112
rect 11233 -14146 11271 -14112
rect 11305 -14146 11343 -14112
rect 11377 -14146 11415 -14112
rect 11449 -14146 11496 -14112
rect 11008 -14152 11496 -14146
rect 11732 -14196 11792 -13848
rect 11848 -14004 11908 -13736
rect 12226 -13792 12298 -13788
rect 12226 -13844 12236 -13792
rect 12288 -13844 12298 -13792
rect 12226 -13848 12298 -13844
rect 11848 -14056 11852 -14004
rect 11904 -14056 11908 -14004
rect 11848 -14066 11908 -14056
rect 12232 -14106 12292 -13848
rect 12372 -13892 12432 -13630
rect 12744 -13678 12804 -13521
rect 13766 -13521 13780 -13514
rect 13814 -13514 13820 -13487
rect 14780 -13487 14840 -13480
rect 13814 -13521 13826 -13514
rect 13044 -13590 13532 -13584
rect 13044 -13624 13091 -13590
rect 13125 -13624 13163 -13590
rect 13197 -13624 13235 -13590
rect 13269 -13624 13307 -13590
rect 13341 -13624 13379 -13590
rect 13413 -13624 13451 -13590
rect 13485 -13624 13532 -13590
rect 13044 -13630 13532 -13624
rect 12738 -13682 12810 -13678
rect 12738 -13734 12748 -13682
rect 12800 -13734 12810 -13682
rect 12738 -13738 12810 -13734
rect 12366 -13896 12438 -13892
rect 12366 -13948 12376 -13896
rect 12428 -13948 12438 -13896
rect 12366 -13952 12438 -13948
rect 12026 -14112 12514 -14106
rect 12026 -14146 12073 -14112
rect 12107 -14146 12145 -14112
rect 12179 -14146 12217 -14112
rect 12251 -14146 12289 -14112
rect 12323 -14146 12361 -14112
rect 12395 -14146 12433 -14112
rect 12467 -14146 12514 -14112
rect 12026 -14152 12514 -14146
rect 10708 -14249 10726 -14215
rect 10760 -14249 10768 -14215
rect 11728 -14215 11792 -14196
rect 11728 -14248 11744 -14215
rect 10708 -14252 10768 -14249
rect 11738 -14249 11744 -14248
rect 11778 -14240 11792 -14215
rect 12744 -14215 12804 -13738
rect 13252 -13792 13324 -13788
rect 13252 -13844 13262 -13792
rect 13314 -13844 13324 -13792
rect 13252 -13848 13324 -13844
rect 13258 -14106 13318 -13848
rect 13380 -13892 13440 -13630
rect 13766 -13676 13826 -13521
rect 14780 -13521 14798 -13487
rect 14832 -13521 14840 -13487
rect 14062 -13590 14550 -13584
rect 14062 -13624 14109 -13590
rect 14143 -13624 14181 -13590
rect 14215 -13624 14253 -13590
rect 14287 -13624 14325 -13590
rect 14359 -13624 14397 -13590
rect 14431 -13624 14469 -13590
rect 14503 -13624 14550 -13590
rect 14062 -13630 14550 -13624
rect 13572 -13736 13826 -13676
rect 13374 -13896 13446 -13892
rect 13374 -13948 13384 -13896
rect 13436 -13948 13446 -13896
rect 13374 -13952 13446 -13948
rect 13572 -14006 13632 -13736
rect 13762 -13792 13834 -13788
rect 13762 -13844 13772 -13792
rect 13824 -13844 13834 -13792
rect 13762 -13848 13834 -13844
rect 14270 -13792 14342 -13788
rect 14270 -13844 14280 -13792
rect 14332 -13844 14342 -13792
rect 14270 -13848 14342 -13844
rect 13572 -14058 13576 -14006
rect 13628 -14058 13632 -14006
rect 13572 -14068 13632 -14058
rect 13044 -14112 13532 -14106
rect 13044 -14146 13091 -14112
rect 13125 -14146 13163 -14112
rect 13197 -14146 13235 -14112
rect 13269 -14146 13307 -14112
rect 13341 -14146 13379 -14112
rect 13413 -14146 13451 -14112
rect 13485 -14146 13532 -14112
rect 13044 -14152 13532 -14146
rect 13768 -14196 13828 -13848
rect 14276 -14106 14336 -13848
rect 14422 -13892 14482 -13630
rect 14780 -13678 14840 -13521
rect 15806 -13487 15866 -13474
rect 15806 -13521 15816 -13487
rect 15850 -13521 15866 -13487
rect 16828 -13487 16874 -13449
rect 17846 -13017 17852 -12990
rect 17886 -12990 17900 -12983
rect 18864 -12983 18910 -12952
rect 17886 -13017 17892 -12990
rect 17846 -13055 17892 -13017
rect 17846 -13089 17852 -13055
rect 17886 -13089 17892 -13055
rect 17846 -13127 17892 -13089
rect 17846 -13161 17852 -13127
rect 17886 -13161 17892 -13127
rect 17846 -13199 17892 -13161
rect 17846 -13233 17852 -13199
rect 17886 -13233 17892 -13199
rect 17846 -13271 17892 -13233
rect 17846 -13305 17852 -13271
rect 17886 -13305 17892 -13271
rect 17846 -13343 17892 -13305
rect 17846 -13377 17852 -13343
rect 17886 -13377 17892 -13343
rect 17846 -13415 17892 -13377
rect 17846 -13449 17852 -13415
rect 17886 -13449 17892 -13415
rect 17846 -13484 17892 -13449
rect 18864 -13017 18870 -12983
rect 18904 -13017 18910 -12983
rect 19874 -12983 19934 -12606
rect 20378 -12874 20438 -12396
rect 20894 -12448 20954 -12287
rect 21912 -12287 21924 -12253
rect 21958 -12287 21972 -12253
rect 21188 -12356 21676 -12350
rect 21188 -12390 21235 -12356
rect 21269 -12390 21307 -12356
rect 21341 -12390 21379 -12356
rect 21413 -12390 21451 -12356
rect 21485 -12390 21523 -12356
rect 21557 -12390 21595 -12356
rect 21629 -12390 21676 -12356
rect 21188 -12396 21676 -12390
rect 20888 -12452 20960 -12448
rect 20888 -12504 20898 -12452
rect 20950 -12504 20960 -12452
rect 20888 -12508 20960 -12504
rect 20170 -12880 20658 -12874
rect 20170 -12914 20217 -12880
rect 20251 -12914 20289 -12880
rect 20323 -12914 20361 -12880
rect 20395 -12914 20433 -12880
rect 20467 -12914 20505 -12880
rect 20539 -12914 20577 -12880
rect 20611 -12914 20658 -12880
rect 20170 -12920 20658 -12914
rect 19874 -13004 19888 -12983
rect 18864 -13055 18910 -13017
rect 18864 -13089 18870 -13055
rect 18904 -13089 18910 -13055
rect 18864 -13127 18910 -13089
rect 18864 -13161 18870 -13127
rect 18904 -13161 18910 -13127
rect 18864 -13199 18910 -13161
rect 18864 -13233 18870 -13199
rect 18904 -13233 18910 -13199
rect 18864 -13271 18910 -13233
rect 18864 -13305 18870 -13271
rect 18904 -13305 18910 -13271
rect 18864 -13343 18910 -13305
rect 18864 -13377 18870 -13343
rect 18904 -13377 18910 -13343
rect 18864 -13415 18910 -13377
rect 18864 -13449 18870 -13415
rect 18904 -13449 18910 -13415
rect 16828 -13490 16834 -13487
rect 15080 -13590 15568 -13584
rect 15080 -13624 15127 -13590
rect 15161 -13624 15199 -13590
rect 15233 -13624 15271 -13590
rect 15305 -13624 15343 -13590
rect 15377 -13624 15415 -13590
rect 15449 -13624 15487 -13590
rect 15521 -13624 15568 -13590
rect 15080 -13630 15568 -13624
rect 14774 -13682 14846 -13678
rect 14774 -13734 14784 -13682
rect 14836 -13734 14846 -13682
rect 14774 -13738 14846 -13734
rect 14416 -13896 14488 -13892
rect 14416 -13948 14426 -13896
rect 14478 -13948 14488 -13896
rect 14416 -13952 14488 -13948
rect 14062 -14112 14550 -14106
rect 14062 -14146 14109 -14112
rect 14143 -14146 14181 -14112
rect 14215 -14146 14253 -14112
rect 14287 -14146 14325 -14112
rect 14359 -14146 14397 -14112
rect 14431 -14146 14469 -14112
rect 14503 -14146 14550 -14112
rect 14062 -14152 14550 -14146
rect 11778 -14248 11788 -14240
rect 12744 -14244 12762 -14215
rect 11778 -14249 11784 -14248
rect 8684 -14321 8690 -14287
rect 8724 -14321 8730 -14287
rect 8684 -14359 8730 -14321
rect 8684 -14393 8690 -14359
rect 8724 -14393 8730 -14359
rect 8684 -14431 8730 -14393
rect 8684 -14465 8690 -14431
rect 8724 -14465 8730 -14431
rect 8684 -14503 8730 -14465
rect 8684 -14537 8690 -14503
rect 8724 -14537 8730 -14503
rect 8684 -14575 8730 -14537
rect 8684 -14609 8690 -14575
rect 8724 -14609 8730 -14575
rect 8684 -14647 8730 -14609
rect 8684 -14681 8690 -14647
rect 8724 -14681 8730 -14647
rect 8684 -14719 8730 -14681
rect 8684 -14730 8690 -14719
rect 7666 -14784 7712 -14753
rect 8676 -14753 8690 -14730
rect 8724 -14730 8730 -14719
rect 9702 -14287 9748 -14258
rect 9702 -14321 9708 -14287
rect 9742 -14321 9748 -14287
rect 9702 -14359 9748 -14321
rect 9702 -14393 9708 -14359
rect 9742 -14393 9748 -14359
rect 9702 -14431 9748 -14393
rect 9702 -14465 9708 -14431
rect 9742 -14465 9748 -14431
rect 9702 -14503 9748 -14465
rect 9702 -14537 9708 -14503
rect 9742 -14537 9748 -14503
rect 9702 -14575 9748 -14537
rect 9702 -14609 9708 -14575
rect 9742 -14609 9748 -14575
rect 9702 -14647 9748 -14609
rect 9702 -14681 9708 -14647
rect 9742 -14681 9748 -14647
rect 9702 -14719 9748 -14681
rect 8724 -14753 8736 -14730
rect 6936 -14822 7424 -14816
rect 6936 -14856 6983 -14822
rect 7017 -14856 7055 -14822
rect 7089 -14856 7127 -14822
rect 7161 -14856 7199 -14822
rect 7233 -14856 7271 -14822
rect 7305 -14856 7343 -14822
rect 7377 -14856 7424 -14822
rect 6936 -14862 7132 -14856
rect 7134 -14862 7424 -14856
rect 7954 -14822 8442 -14816
rect 7954 -14856 8001 -14822
rect 8035 -14856 8073 -14822
rect 8107 -14856 8145 -14822
rect 8179 -14856 8217 -14822
rect 8251 -14856 8289 -14822
rect 8323 -14856 8361 -14822
rect 8395 -14856 8442 -14822
rect 7954 -14862 8442 -14856
rect 7134 -14890 7194 -14862
rect 8160 -14890 8220 -14862
rect 7128 -14894 7200 -14890
rect 7128 -14946 7138 -14894
rect 7190 -14946 7200 -14894
rect 7128 -14950 7200 -14946
rect 8154 -14894 8226 -14890
rect 8154 -14946 8164 -14894
rect 8216 -14946 8226 -14894
rect 8154 -14950 8226 -14946
rect 6628 -14998 6700 -14994
rect 6628 -15050 6638 -14998
rect 6690 -15050 6700 -14998
rect 6628 -15054 6700 -15050
rect 6634 -15232 6706 -15228
rect 6634 -15284 6644 -15232
rect 6696 -15284 6706 -15232
rect 6634 -15288 6706 -15284
rect 5916 -15346 6120 -15340
rect 6122 -15346 6404 -15340
rect 5916 -15380 5963 -15346
rect 5997 -15380 6035 -15346
rect 6069 -15380 6107 -15346
rect 6141 -15380 6179 -15346
rect 6213 -15380 6251 -15346
rect 6285 -15380 6323 -15346
rect 6357 -15380 6404 -15346
rect 5916 -15386 6404 -15380
rect 4650 -15483 4656 -15456
rect 5622 -15462 5634 -15449
rect 4610 -15521 4656 -15483
rect 4610 -15555 4616 -15521
rect 4650 -15555 4656 -15521
rect 4610 -15593 4656 -15555
rect 4610 -15627 4616 -15593
rect 4650 -15627 4656 -15593
rect 4610 -15665 4656 -15627
rect 4610 -15699 4616 -15665
rect 4650 -15699 4656 -15665
rect 4610 -15737 4656 -15699
rect 4610 -15771 4616 -15737
rect 4650 -15771 4656 -15737
rect 4610 -15809 4656 -15771
rect 4610 -15843 4616 -15809
rect 4650 -15843 4656 -15809
rect 4610 -15881 4656 -15843
rect 4610 -15915 4616 -15881
rect 4650 -15915 4656 -15881
rect 4610 -15953 4656 -15915
rect 3632 -15987 3646 -15962
rect 2862 -16056 3350 -16050
rect 2862 -16090 2909 -16056
rect 2943 -16090 2981 -16056
rect 3015 -16090 3053 -16056
rect 3087 -16090 3125 -16056
rect 3159 -16090 3197 -16056
rect 3231 -16090 3269 -16056
rect 3303 -16090 3350 -16056
rect 2862 -16096 3350 -16090
rect 3586 -16158 3646 -15987
rect 4610 -15987 4616 -15953
rect 4650 -15987 4656 -15953
rect 5628 -15483 5634 -15462
rect 5668 -15462 5682 -15449
rect 6640 -15449 6700 -15288
rect 7134 -15340 7194 -14950
rect 7648 -14998 7720 -14994
rect 7648 -15050 7658 -14998
rect 7710 -15050 7720 -14998
rect 7648 -15054 7720 -15050
rect 6934 -15346 7132 -15340
rect 7134 -15346 7422 -15340
rect 6934 -15380 6981 -15346
rect 7015 -15380 7053 -15346
rect 7087 -15380 7125 -15346
rect 7159 -15380 7197 -15346
rect 7231 -15380 7269 -15346
rect 7303 -15380 7341 -15346
rect 7375 -15380 7422 -15346
rect 6934 -15386 7422 -15380
rect 6640 -15460 6652 -15449
rect 5668 -15483 5674 -15462
rect 5628 -15521 5674 -15483
rect 5628 -15555 5634 -15521
rect 5668 -15555 5674 -15521
rect 5628 -15593 5674 -15555
rect 5628 -15627 5634 -15593
rect 5668 -15627 5674 -15593
rect 5628 -15665 5674 -15627
rect 5628 -15699 5634 -15665
rect 5668 -15699 5674 -15665
rect 5628 -15737 5674 -15699
rect 5628 -15771 5634 -15737
rect 5668 -15771 5674 -15737
rect 5628 -15809 5674 -15771
rect 5628 -15843 5634 -15809
rect 5668 -15843 5674 -15809
rect 5628 -15881 5674 -15843
rect 5628 -15915 5634 -15881
rect 5668 -15915 5674 -15881
rect 5628 -15953 5674 -15915
rect 5628 -15966 5634 -15953
rect 4610 -16018 4656 -15987
rect 5620 -15987 5634 -15966
rect 5668 -15966 5674 -15953
rect 6646 -15483 6652 -15460
rect 6686 -15460 6700 -15449
rect 7654 -15449 7714 -15054
rect 8160 -15340 8220 -14950
rect 8676 -14994 8736 -14753
rect 9702 -14753 9708 -14719
rect 9742 -14753 9748 -14719
rect 10720 -14287 10766 -14252
rect 10720 -14321 10726 -14287
rect 10760 -14321 10766 -14287
rect 10720 -14359 10766 -14321
rect 10720 -14393 10726 -14359
rect 10760 -14393 10766 -14359
rect 10720 -14431 10766 -14393
rect 10720 -14465 10726 -14431
rect 10760 -14465 10766 -14431
rect 10720 -14503 10766 -14465
rect 10720 -14537 10726 -14503
rect 10760 -14537 10766 -14503
rect 10720 -14575 10766 -14537
rect 10720 -14609 10726 -14575
rect 10760 -14609 10766 -14575
rect 10720 -14647 10766 -14609
rect 10720 -14681 10726 -14647
rect 10760 -14681 10766 -14647
rect 11738 -14287 11784 -14249
rect 11738 -14321 11744 -14287
rect 11778 -14321 11784 -14287
rect 11738 -14359 11784 -14321
rect 11738 -14393 11744 -14359
rect 11778 -14393 11784 -14359
rect 11738 -14431 11784 -14393
rect 11738 -14465 11744 -14431
rect 11778 -14465 11784 -14431
rect 11738 -14503 11784 -14465
rect 11738 -14537 11744 -14503
rect 11778 -14537 11784 -14503
rect 11738 -14575 11784 -14537
rect 11738 -14609 11744 -14575
rect 11778 -14609 11784 -14575
rect 11738 -14647 11784 -14609
rect 11738 -14648 11744 -14647
rect 10720 -14719 10766 -14681
rect 10720 -14730 10726 -14719
rect 9702 -14784 9748 -14753
rect 10712 -14753 10726 -14730
rect 10760 -14730 10766 -14719
rect 11778 -14648 11784 -14647
rect 12756 -14249 12762 -14244
rect 12796 -14244 12804 -14215
rect 13764 -14215 13830 -14196
rect 13764 -14236 13780 -14215
rect 12796 -14249 12802 -14244
rect 12756 -14287 12802 -14249
rect 12756 -14321 12762 -14287
rect 12796 -14321 12802 -14287
rect 12756 -14359 12802 -14321
rect 12756 -14393 12762 -14359
rect 12796 -14393 12802 -14359
rect 12756 -14431 12802 -14393
rect 12756 -14465 12762 -14431
rect 12796 -14465 12802 -14431
rect 12756 -14503 12802 -14465
rect 12756 -14537 12762 -14503
rect 12796 -14537 12802 -14503
rect 12756 -14575 12802 -14537
rect 12756 -14609 12762 -14575
rect 12796 -14609 12802 -14575
rect 12756 -14647 12802 -14609
rect 11744 -14719 11778 -14681
rect 10760 -14753 10772 -14730
rect 8972 -14822 9460 -14816
rect 8972 -14856 9019 -14822
rect 9053 -14856 9091 -14822
rect 9125 -14856 9163 -14822
rect 9197 -14856 9235 -14822
rect 9269 -14856 9307 -14822
rect 9341 -14856 9379 -14822
rect 9413 -14856 9460 -14822
rect 8972 -14862 9460 -14856
rect 9990 -14822 10478 -14816
rect 9990 -14856 10037 -14822
rect 10071 -14856 10109 -14822
rect 10143 -14856 10181 -14822
rect 10215 -14856 10253 -14822
rect 10287 -14856 10325 -14822
rect 10359 -14856 10397 -14822
rect 10431 -14856 10478 -14822
rect 9990 -14862 10478 -14856
rect 10712 -14994 10772 -14753
rect 11730 -14753 11744 -14724
rect 12756 -14681 12762 -14647
rect 12796 -14681 12802 -14647
rect 13774 -14249 13780 -14236
rect 13814 -14234 13830 -14215
rect 14780 -14215 14840 -13738
rect 15284 -13788 15344 -13630
rect 15806 -13788 15866 -13521
rect 16818 -13521 16834 -13490
rect 16868 -13490 16874 -13487
rect 17838 -13486 17898 -13484
rect 17838 -13487 17900 -13486
rect 16868 -13521 16878 -13490
rect 16296 -13584 16356 -13582
rect 16098 -13590 16586 -13584
rect 16098 -13624 16145 -13590
rect 16179 -13624 16217 -13590
rect 16251 -13624 16289 -13590
rect 16323 -13624 16361 -13590
rect 16395 -13624 16433 -13590
rect 16467 -13624 16505 -13590
rect 16539 -13624 16586 -13590
rect 16098 -13630 16586 -13624
rect 16296 -13788 16356 -13630
rect 16818 -13678 16878 -13521
rect 17838 -13521 17852 -13487
rect 17886 -13521 17900 -13487
rect 18864 -13487 18910 -13449
rect 18864 -13504 18870 -13487
rect 17838 -13540 17900 -13521
rect 17328 -13584 17388 -13582
rect 17116 -13590 17604 -13584
rect 17116 -13624 17163 -13590
rect 17197 -13624 17235 -13590
rect 17269 -13624 17307 -13590
rect 17341 -13624 17379 -13590
rect 17413 -13624 17451 -13590
rect 17485 -13624 17523 -13590
rect 17557 -13624 17604 -13590
rect 17116 -13630 17604 -13624
rect 16812 -13682 16884 -13678
rect 16812 -13734 16822 -13682
rect 16874 -13734 16884 -13682
rect 16812 -13738 16884 -13734
rect 15278 -13792 15350 -13788
rect 15278 -13844 15288 -13792
rect 15340 -13844 15350 -13792
rect 15278 -13848 15350 -13844
rect 15800 -13792 15872 -13788
rect 15800 -13844 15810 -13792
rect 15862 -13844 15872 -13792
rect 15800 -13848 15872 -13844
rect 16290 -13792 16362 -13788
rect 16290 -13844 16300 -13792
rect 16352 -13844 16362 -13792
rect 16290 -13848 16362 -13844
rect 15284 -14106 15344 -13848
rect 15800 -14004 15872 -14000
rect 15800 -14056 15810 -14004
rect 15862 -14056 15872 -14004
rect 15800 -14060 15872 -14056
rect 15080 -14112 15568 -14106
rect 15080 -14146 15127 -14112
rect 15161 -14146 15199 -14112
rect 15233 -14146 15271 -14112
rect 15305 -14146 15343 -14112
rect 15377 -14146 15415 -14112
rect 15449 -14146 15487 -14112
rect 15521 -14146 15568 -14112
rect 15080 -14152 15568 -14146
rect 13814 -14236 13828 -14234
rect 13814 -14249 13820 -14236
rect 14780 -14242 14798 -14215
rect 13774 -14287 13820 -14249
rect 13774 -14321 13780 -14287
rect 13814 -14321 13820 -14287
rect 13774 -14359 13820 -14321
rect 13774 -14393 13780 -14359
rect 13814 -14393 13820 -14359
rect 13774 -14431 13820 -14393
rect 13774 -14465 13780 -14431
rect 13814 -14465 13820 -14431
rect 13774 -14503 13820 -14465
rect 13774 -14537 13780 -14503
rect 13814 -14537 13820 -14503
rect 13774 -14575 13820 -14537
rect 13774 -14609 13780 -14575
rect 13814 -14609 13820 -14575
rect 13774 -14647 13820 -14609
rect 13774 -14658 13780 -14647
rect 12756 -14719 12802 -14681
rect 12756 -14724 12762 -14719
rect 11778 -14753 11790 -14724
rect 11008 -14822 11176 -14816
rect 11008 -14856 11055 -14822
rect 11089 -14856 11127 -14822
rect 11161 -14856 11199 -14822
rect 11233 -14856 11271 -14822
rect 11305 -14856 11343 -14822
rect 11377 -14856 11415 -14822
rect 11449 -14856 11484 -14822
rect 11008 -14862 11176 -14856
rect 11212 -14922 11272 -14856
rect 11730 -14922 11790 -14753
rect 12750 -14753 12762 -14724
rect 12796 -14724 12802 -14719
rect 13814 -14658 13820 -14647
rect 14792 -14249 14798 -14242
rect 14832 -14242 14840 -14215
rect 15806 -14215 15866 -14060
rect 16296 -14106 16356 -13848
rect 16098 -14112 16586 -14106
rect 16098 -14146 16145 -14112
rect 16179 -14146 16217 -14112
rect 16251 -14146 16289 -14112
rect 16323 -14146 16361 -14112
rect 16395 -14146 16433 -14112
rect 16467 -14146 16505 -14112
rect 16539 -14146 16586 -14112
rect 16098 -14152 16586 -14146
rect 15806 -14238 15816 -14215
rect 14832 -14249 14838 -14242
rect 14792 -14287 14838 -14249
rect 14792 -14321 14798 -14287
rect 14832 -14321 14838 -14287
rect 14792 -14359 14838 -14321
rect 14792 -14393 14798 -14359
rect 14832 -14393 14838 -14359
rect 14792 -14431 14838 -14393
rect 14792 -14465 14798 -14431
rect 14832 -14465 14838 -14431
rect 14792 -14503 14838 -14465
rect 14792 -14537 14798 -14503
rect 14832 -14537 14838 -14503
rect 14792 -14575 14838 -14537
rect 14792 -14609 14798 -14575
rect 14832 -14609 14838 -14575
rect 14792 -14647 14838 -14609
rect 13780 -14719 13814 -14681
rect 14792 -14681 14798 -14647
rect 14832 -14681 14838 -14647
rect 14792 -14718 14838 -14681
rect 15810 -14249 15816 -14238
rect 15850 -14238 15866 -14215
rect 16818 -14215 16878 -13738
rect 17328 -13788 17388 -13630
rect 17840 -13788 17900 -13540
rect 18856 -13521 18870 -13504
rect 18904 -13504 18910 -13487
rect 19882 -13017 19888 -13004
rect 19922 -13004 19934 -12983
rect 20894 -12983 20954 -12508
rect 21404 -12874 21464 -12396
rect 21912 -12546 21972 -12287
rect 22924 -12253 22984 -12252
rect 22924 -12287 22942 -12253
rect 22976 -12287 22984 -12253
rect 22206 -12356 22694 -12350
rect 22206 -12390 22253 -12356
rect 22287 -12390 22325 -12356
rect 22359 -12390 22397 -12356
rect 22431 -12390 22469 -12356
rect 22503 -12390 22541 -12356
rect 22575 -12390 22613 -12356
rect 22647 -12390 22694 -12356
rect 22206 -12396 22694 -12390
rect 21906 -12550 21978 -12546
rect 21906 -12602 21916 -12550
rect 21968 -12602 21978 -12550
rect 21906 -12606 21978 -12602
rect 21188 -12880 21676 -12874
rect 21188 -12914 21235 -12880
rect 21269 -12914 21307 -12880
rect 21341 -12914 21379 -12880
rect 21413 -12914 21451 -12880
rect 21485 -12914 21523 -12880
rect 21557 -12914 21595 -12880
rect 21629 -12914 21676 -12880
rect 21188 -12920 21676 -12914
rect 20894 -12996 20906 -12983
rect 19922 -13017 19928 -13004
rect 19882 -13055 19928 -13017
rect 19882 -13089 19888 -13055
rect 19922 -13089 19928 -13055
rect 19882 -13127 19928 -13089
rect 19882 -13161 19888 -13127
rect 19922 -13161 19928 -13127
rect 19882 -13199 19928 -13161
rect 19882 -13233 19888 -13199
rect 19922 -13233 19928 -13199
rect 19882 -13271 19928 -13233
rect 19882 -13305 19888 -13271
rect 19922 -13305 19928 -13271
rect 19882 -13343 19928 -13305
rect 19882 -13377 19888 -13343
rect 19922 -13377 19928 -13343
rect 19882 -13415 19928 -13377
rect 19882 -13449 19888 -13415
rect 19922 -13449 19928 -13415
rect 19882 -13487 19928 -13449
rect 18904 -13521 18916 -13504
rect 18134 -13590 18622 -13584
rect 18134 -13624 18181 -13590
rect 18215 -13624 18253 -13590
rect 18287 -13624 18325 -13590
rect 18359 -13624 18397 -13590
rect 18431 -13624 18469 -13590
rect 18503 -13624 18541 -13590
rect 18575 -13624 18622 -13590
rect 18134 -13630 18622 -13624
rect 18342 -13682 18402 -13630
rect 18856 -13678 18916 -13521
rect 19882 -13521 19888 -13487
rect 19922 -13521 19928 -13487
rect 19882 -13552 19928 -13521
rect 20900 -13017 20906 -12996
rect 20940 -12996 20954 -12983
rect 21912 -12983 21972 -12606
rect 22426 -12874 22486 -12396
rect 22924 -12448 22984 -12287
rect 24816 -12269 24855 -12235
rect 24889 -12269 24928 -12235
rect 24816 -12307 24928 -12269
rect 24816 -12341 24855 -12307
rect 24889 -12341 24928 -12307
rect 24816 -12379 24928 -12341
rect 24816 -12413 24855 -12379
rect 24889 -12413 24928 -12379
rect 22918 -12452 22990 -12448
rect 22918 -12504 22928 -12452
rect 22980 -12504 22990 -12452
rect 22918 -12508 22990 -12504
rect 24816 -12451 24928 -12413
rect 24816 -12485 24855 -12451
rect 24889 -12485 24928 -12451
rect 22206 -12880 22694 -12874
rect 22206 -12914 22253 -12880
rect 22287 -12914 22325 -12880
rect 22359 -12914 22397 -12880
rect 22431 -12914 22469 -12880
rect 22503 -12914 22541 -12880
rect 22575 -12914 22613 -12880
rect 22647 -12914 22694 -12880
rect 22206 -12920 22694 -12914
rect 21912 -12992 21924 -12983
rect 20940 -13017 20946 -12996
rect 20900 -13055 20946 -13017
rect 20900 -13089 20906 -13055
rect 20940 -13089 20946 -13055
rect 20900 -13127 20946 -13089
rect 20900 -13161 20906 -13127
rect 20940 -13161 20946 -13127
rect 20900 -13199 20946 -13161
rect 20900 -13233 20906 -13199
rect 20940 -13233 20946 -13199
rect 20900 -13271 20946 -13233
rect 20900 -13305 20906 -13271
rect 20940 -13305 20946 -13271
rect 20900 -13343 20946 -13305
rect 20900 -13377 20906 -13343
rect 20940 -13377 20946 -13343
rect 20900 -13415 20946 -13377
rect 20900 -13449 20906 -13415
rect 20940 -13449 20946 -13415
rect 20900 -13487 20946 -13449
rect 20900 -13521 20906 -13487
rect 20940 -13521 20946 -13487
rect 20900 -13552 20946 -13521
rect 21918 -13017 21924 -12992
rect 21958 -12992 21972 -12983
rect 22924 -12983 22984 -12508
rect 24816 -12523 24928 -12485
rect 23642 -12550 23714 -12546
rect 23642 -12602 23652 -12550
rect 23704 -12602 23714 -12550
rect 23642 -12606 23714 -12602
rect 24816 -12557 24855 -12523
rect 24889 -12557 24928 -12523
rect 24816 -12595 24928 -12557
rect 22924 -12990 22942 -12983
rect 21958 -13017 21964 -12992
rect 21918 -13055 21964 -13017
rect 21918 -13089 21924 -13055
rect 21958 -13089 21964 -13055
rect 21918 -13127 21964 -13089
rect 21918 -13161 21924 -13127
rect 21958 -13161 21964 -13127
rect 21918 -13199 21964 -13161
rect 21918 -13233 21924 -13199
rect 21958 -13233 21964 -13199
rect 21918 -13271 21964 -13233
rect 21918 -13305 21924 -13271
rect 21958 -13305 21964 -13271
rect 21918 -13343 21964 -13305
rect 21918 -13377 21924 -13343
rect 21958 -13377 21964 -13343
rect 21918 -13415 21964 -13377
rect 21918 -13449 21924 -13415
rect 21958 -13449 21964 -13415
rect 21918 -13487 21964 -13449
rect 21918 -13521 21924 -13487
rect 21958 -13521 21964 -13487
rect 21918 -13552 21964 -13521
rect 22936 -13017 22942 -12990
rect 22976 -12990 22984 -12983
rect 22976 -13017 22982 -12990
rect 22936 -13055 22982 -13017
rect 22936 -13089 22942 -13055
rect 22976 -13089 22982 -13055
rect 22936 -13127 22982 -13089
rect 22936 -13161 22942 -13127
rect 22976 -13161 22982 -13127
rect 22936 -13199 22982 -13161
rect 22936 -13233 22942 -13199
rect 22976 -13233 22982 -13199
rect 22936 -13271 22982 -13233
rect 22936 -13305 22942 -13271
rect 22976 -13305 22982 -13271
rect 22936 -13343 22982 -13305
rect 22936 -13377 22942 -13343
rect 22976 -13377 22982 -13343
rect 22936 -13415 22982 -13377
rect 22936 -13449 22942 -13415
rect 22976 -13449 22982 -13415
rect 22936 -13487 22982 -13449
rect 22936 -13521 22942 -13487
rect 22976 -13521 22982 -13487
rect 22936 -13552 22982 -13521
rect 19152 -13590 19640 -13584
rect 19152 -13624 19199 -13590
rect 19233 -13624 19271 -13590
rect 19305 -13624 19343 -13590
rect 19377 -13624 19415 -13590
rect 19449 -13624 19487 -13590
rect 19521 -13624 19559 -13590
rect 19593 -13624 19640 -13590
rect 19152 -13630 19640 -13624
rect 20170 -13590 20658 -13584
rect 20170 -13624 20217 -13590
rect 20251 -13624 20289 -13590
rect 20323 -13624 20361 -13590
rect 20395 -13624 20433 -13590
rect 20467 -13624 20505 -13590
rect 20539 -13624 20577 -13590
rect 20611 -13624 20658 -13590
rect 20170 -13630 20658 -13624
rect 21188 -13590 21676 -13584
rect 21188 -13624 21235 -13590
rect 21269 -13624 21307 -13590
rect 21341 -13624 21379 -13590
rect 21413 -13624 21451 -13590
rect 21485 -13624 21523 -13590
rect 21557 -13624 21595 -13590
rect 21629 -13624 21676 -13590
rect 21188 -13630 21676 -13624
rect 22206 -13590 22694 -13584
rect 22206 -13624 22253 -13590
rect 22287 -13624 22325 -13590
rect 22359 -13624 22397 -13590
rect 22431 -13624 22469 -13590
rect 22503 -13624 22541 -13590
rect 22575 -13624 22613 -13590
rect 22647 -13624 22694 -13590
rect 22206 -13630 22694 -13624
rect 19364 -13678 19424 -13630
rect 18342 -13734 18346 -13682
rect 18398 -13734 18402 -13682
rect 18342 -13744 18402 -13734
rect 18850 -13682 18922 -13678
rect 18850 -13734 18860 -13682
rect 18912 -13734 18922 -13682
rect 18850 -13738 18922 -13734
rect 19358 -13682 19430 -13678
rect 19358 -13734 19368 -13682
rect 19420 -13734 19430 -13682
rect 19358 -13738 19430 -13734
rect 17322 -13792 17394 -13788
rect 17322 -13844 17332 -13792
rect 17384 -13844 17394 -13792
rect 17322 -13848 17394 -13844
rect 17834 -13792 17906 -13788
rect 17834 -13844 17844 -13792
rect 17896 -13844 17906 -13792
rect 17834 -13848 17906 -13844
rect 17308 -13896 17380 -13892
rect 17308 -13948 17318 -13896
rect 17370 -13948 17380 -13896
rect 17308 -13952 17380 -13948
rect 18346 -13896 18418 -13892
rect 18346 -13948 18356 -13896
rect 18408 -13948 18418 -13896
rect 18346 -13952 18418 -13948
rect 17314 -14106 17374 -13952
rect 17832 -14004 17904 -14000
rect 17832 -14056 17842 -14004
rect 17894 -14056 17904 -14004
rect 17832 -14060 17904 -14056
rect 17116 -14112 17604 -14106
rect 17116 -14146 17163 -14112
rect 17197 -14146 17235 -14112
rect 17269 -14146 17307 -14112
rect 17341 -14146 17379 -14112
rect 17413 -14146 17451 -14112
rect 17485 -14146 17523 -14112
rect 17557 -14146 17604 -14112
rect 17116 -14152 17604 -14146
rect 15850 -14249 15856 -14238
rect 15810 -14287 15856 -14249
rect 15810 -14321 15816 -14287
rect 15850 -14321 15856 -14287
rect 15810 -14359 15856 -14321
rect 15810 -14393 15816 -14359
rect 15850 -14393 15856 -14359
rect 15810 -14431 15856 -14393
rect 15810 -14465 15816 -14431
rect 15850 -14465 15856 -14431
rect 15810 -14503 15856 -14465
rect 15810 -14537 15816 -14503
rect 15850 -14537 15856 -14503
rect 15810 -14575 15856 -14537
rect 15810 -14609 15816 -14575
rect 15850 -14609 15856 -14575
rect 15810 -14647 15856 -14609
rect 15810 -14681 15816 -14647
rect 15850 -14681 15856 -14647
rect 12796 -14753 12810 -14724
rect 12424 -14822 12514 -14816
rect 12038 -14856 12073 -14822
rect 12107 -14856 12145 -14822
rect 12179 -14856 12217 -14822
rect 12251 -14856 12289 -14822
rect 12323 -14856 12361 -14822
rect 12395 -14856 12433 -14822
rect 12467 -14856 12514 -14822
rect 12232 -14922 12292 -14856
rect 12424 -14862 12514 -14856
rect 11212 -14982 12292 -14922
rect 12750 -14994 12810 -14753
rect 13780 -14754 13814 -14753
rect 14780 -14719 14840 -14718
rect 14780 -14753 14798 -14719
rect 14832 -14753 14840 -14719
rect 13044 -14822 13236 -14816
rect 13044 -14856 13091 -14822
rect 13125 -14856 13163 -14822
rect 13197 -14856 13235 -14822
rect 13269 -14856 13307 -14822
rect 13341 -14856 13379 -14822
rect 13413 -14856 13451 -14822
rect 13485 -14856 13520 -14822
rect 13044 -14862 13236 -14856
rect 13256 -14918 13316 -14856
rect 13768 -14918 13828 -14754
rect 14062 -14822 14550 -14816
rect 14074 -14856 14109 -14822
rect 14143 -14856 14181 -14822
rect 14215 -14856 14253 -14822
rect 14287 -14856 14325 -14822
rect 14359 -14856 14397 -14822
rect 14431 -14856 14469 -14822
rect 14503 -14856 14550 -14822
rect 14062 -14862 14550 -14856
rect 14258 -14918 14318 -14862
rect 13256 -14978 14318 -14918
rect 14780 -14994 14840 -14753
rect 15810 -14719 15856 -14681
rect 15810 -14753 15816 -14719
rect 15850 -14753 15856 -14719
rect 15810 -14784 15856 -14753
rect 16818 -14249 16834 -14215
rect 16868 -14249 16878 -14215
rect 17838 -14215 17898 -14060
rect 18352 -14106 18412 -13952
rect 18134 -14112 18622 -14106
rect 18134 -14146 18181 -14112
rect 18215 -14146 18253 -14112
rect 18287 -14146 18325 -14112
rect 18359 -14146 18397 -14112
rect 18431 -14146 18469 -14112
rect 18503 -14146 18541 -14112
rect 18575 -14146 18622 -14112
rect 18134 -14152 18622 -14146
rect 17838 -14238 17852 -14215
rect 16818 -14287 16878 -14249
rect 16818 -14321 16834 -14287
rect 16868 -14321 16878 -14287
rect 16818 -14359 16878 -14321
rect 16818 -14393 16834 -14359
rect 16868 -14393 16878 -14359
rect 16818 -14431 16878 -14393
rect 16818 -14465 16834 -14431
rect 16868 -14465 16878 -14431
rect 16818 -14503 16878 -14465
rect 16818 -14537 16834 -14503
rect 16868 -14537 16878 -14503
rect 16818 -14575 16878 -14537
rect 16818 -14609 16834 -14575
rect 16868 -14609 16878 -14575
rect 16818 -14647 16878 -14609
rect 16818 -14681 16834 -14647
rect 16868 -14681 16878 -14647
rect 16818 -14719 16878 -14681
rect 16818 -14753 16834 -14719
rect 16868 -14753 16878 -14719
rect 15080 -14822 15568 -14816
rect 15080 -14856 15127 -14822
rect 15161 -14856 15199 -14822
rect 15233 -14856 15271 -14822
rect 15305 -14856 15343 -14822
rect 15377 -14856 15415 -14822
rect 15449 -14856 15487 -14822
rect 15521 -14856 15568 -14822
rect 15080 -14862 15568 -14856
rect 16098 -14822 16586 -14816
rect 16098 -14856 16145 -14822
rect 16179 -14856 16217 -14822
rect 16251 -14856 16289 -14822
rect 16323 -14856 16361 -14822
rect 16395 -14856 16433 -14822
rect 16467 -14856 16505 -14822
rect 16539 -14856 16586 -14822
rect 16098 -14862 16586 -14856
rect 15304 -14964 16366 -14904
rect 8670 -14998 8742 -14994
rect 8670 -15050 8680 -14998
rect 8732 -15050 8742 -14998
rect 8670 -15054 8742 -15050
rect 10706 -14998 10778 -14994
rect 10706 -15050 10716 -14998
rect 10768 -15050 10778 -14998
rect 10706 -15054 10778 -15050
rect 12744 -14998 12816 -14994
rect 12744 -15050 12754 -14998
rect 12806 -15050 12816 -14998
rect 12744 -15054 12816 -15050
rect 14774 -14998 14846 -14994
rect 14774 -15050 14784 -14998
rect 14836 -15050 14846 -14998
rect 14774 -15054 14846 -15050
rect 9690 -15120 9762 -15116
rect 9690 -15172 9700 -15120
rect 9752 -15172 9762 -15120
rect 9690 -15176 9762 -15172
rect 11724 -15120 11796 -15116
rect 11724 -15172 11734 -15120
rect 11786 -15172 11796 -15120
rect 11724 -15176 11796 -15172
rect 13754 -15120 13826 -15116
rect 13754 -15172 13764 -15120
rect 13816 -15172 13826 -15120
rect 13754 -15176 13826 -15172
rect 7952 -15346 8440 -15340
rect 7952 -15380 7999 -15346
rect 8033 -15380 8071 -15346
rect 8105 -15380 8143 -15346
rect 8177 -15380 8215 -15346
rect 8249 -15380 8287 -15346
rect 8321 -15380 8359 -15346
rect 8393 -15380 8440 -15346
rect 7952 -15386 8440 -15380
rect 8970 -15346 9458 -15340
rect 8970 -15380 9017 -15346
rect 9051 -15380 9089 -15346
rect 9123 -15380 9161 -15346
rect 9195 -15380 9233 -15346
rect 9267 -15380 9305 -15346
rect 9339 -15380 9377 -15346
rect 9411 -15380 9458 -15346
rect 8970 -15386 9458 -15380
rect 6686 -15483 6692 -15460
rect 7654 -15474 7670 -15449
rect 6646 -15521 6692 -15483
rect 6646 -15555 6652 -15521
rect 6686 -15555 6692 -15521
rect 6646 -15593 6692 -15555
rect 6646 -15627 6652 -15593
rect 6686 -15627 6692 -15593
rect 6646 -15665 6692 -15627
rect 6646 -15699 6652 -15665
rect 6686 -15699 6692 -15665
rect 6646 -15737 6692 -15699
rect 6646 -15771 6652 -15737
rect 6686 -15771 6692 -15737
rect 6646 -15809 6692 -15771
rect 6646 -15843 6652 -15809
rect 6686 -15843 6692 -15809
rect 6646 -15881 6692 -15843
rect 6646 -15915 6652 -15881
rect 6686 -15915 6692 -15881
rect 6646 -15953 6692 -15915
rect 5668 -15987 5680 -15966
rect 3880 -16056 4368 -16050
rect 3880 -16090 3927 -16056
rect 3961 -16090 3999 -16056
rect 4033 -16090 4071 -16056
rect 4105 -16090 4143 -16056
rect 4177 -16090 4215 -16056
rect 4249 -16090 4287 -16056
rect 4321 -16090 4368 -16056
rect 3880 -16096 4368 -16090
rect 4898 -16056 5386 -16050
rect 4898 -16090 4945 -16056
rect 4979 -16090 5017 -16056
rect 5051 -16090 5089 -16056
rect 5123 -16090 5161 -16056
rect 5195 -16090 5233 -16056
rect 5267 -16090 5305 -16056
rect 5339 -16090 5386 -16056
rect 4898 -16096 5386 -16090
rect 2442 -16162 2514 -16158
rect 2442 -16214 2452 -16162
rect 2504 -16214 2514 -16162
rect 2442 -16218 2514 -16214
rect 3580 -16162 3652 -16158
rect 3580 -16214 3590 -16162
rect 3642 -16214 3652 -16162
rect 3580 -16218 3652 -16214
rect 2330 -16362 2402 -16358
rect 2330 -16414 2340 -16362
rect 2392 -16414 2402 -16362
rect 2330 -16418 2402 -16414
rect 2224 -16464 2296 -16460
rect 2224 -16516 2234 -16464
rect 2286 -16516 2296 -16464
rect 2224 -16520 2296 -16516
rect 2230 -19950 2290 -16520
rect 2336 -17594 2396 -16418
rect 2330 -17598 2402 -17594
rect 2330 -17650 2340 -17598
rect 2392 -17650 2402 -17598
rect 2330 -17654 2402 -17650
rect 2224 -19954 2296 -19950
rect 2224 -20006 2234 -19954
rect 2286 -20006 2296 -19954
rect 2224 -20010 2296 -20006
rect 2230 -21254 2290 -20010
rect 2336 -20196 2396 -17654
rect 2448 -18932 2508 -16218
rect 3578 -16362 3650 -16358
rect 3578 -16414 3588 -16362
rect 3640 -16414 3650 -16362
rect 3578 -16418 3650 -16414
rect 3584 -16462 3644 -16418
rect 2568 -16522 3644 -16462
rect 2568 -16524 3132 -16522
rect 2568 -16683 2628 -16524
rect 3072 -16574 3132 -16524
rect 2862 -16580 3350 -16574
rect 2862 -16614 2909 -16580
rect 2943 -16614 2981 -16580
rect 3015 -16614 3053 -16580
rect 3087 -16614 3125 -16580
rect 3159 -16614 3197 -16580
rect 3231 -16614 3269 -16580
rect 3303 -16614 3350 -16580
rect 2862 -16620 3350 -16614
rect 2568 -16696 2580 -16683
rect 2574 -16717 2580 -16696
rect 2614 -16696 2628 -16683
rect 3584 -16683 3644 -16522
rect 4088 -16574 4148 -16096
rect 4596 -16242 4668 -16238
rect 4596 -16294 4606 -16242
rect 4658 -16294 4668 -16242
rect 4596 -16298 4668 -16294
rect 3880 -16580 4368 -16574
rect 3880 -16614 3927 -16580
rect 3961 -16614 3999 -16580
rect 4033 -16614 4071 -16580
rect 4105 -16614 4143 -16580
rect 4177 -16614 4215 -16580
rect 4249 -16614 4287 -16580
rect 4321 -16614 4368 -16580
rect 3880 -16620 4368 -16614
rect 2614 -16717 2620 -16696
rect 3584 -16700 3598 -16683
rect 2574 -16755 2620 -16717
rect 2574 -16789 2580 -16755
rect 2614 -16789 2620 -16755
rect 2574 -16827 2620 -16789
rect 2574 -16861 2580 -16827
rect 2614 -16861 2620 -16827
rect 2574 -16899 2620 -16861
rect 2574 -16933 2580 -16899
rect 2614 -16933 2620 -16899
rect 2574 -16971 2620 -16933
rect 2574 -17005 2580 -16971
rect 2614 -17005 2620 -16971
rect 2574 -17043 2620 -17005
rect 2574 -17077 2580 -17043
rect 2614 -17077 2620 -17043
rect 2574 -17115 2620 -17077
rect 2574 -17149 2580 -17115
rect 2614 -17149 2620 -17115
rect 2574 -17187 2620 -17149
rect 2574 -17221 2580 -17187
rect 2614 -17221 2620 -17187
rect 2574 -17252 2620 -17221
rect 3592 -16717 3598 -16700
rect 3632 -16700 3644 -16683
rect 4602 -16683 4662 -16298
rect 5116 -16352 5176 -16096
rect 5620 -16134 5680 -15987
rect 6646 -15987 6652 -15953
rect 6686 -15987 6692 -15953
rect 7664 -15483 7670 -15474
rect 7704 -15474 7714 -15449
rect 8682 -15449 8728 -15418
rect 7704 -15483 7710 -15474
rect 7664 -15521 7710 -15483
rect 7664 -15555 7670 -15521
rect 7704 -15555 7710 -15521
rect 7664 -15593 7710 -15555
rect 7664 -15627 7670 -15593
rect 7704 -15627 7710 -15593
rect 7664 -15665 7710 -15627
rect 7664 -15699 7670 -15665
rect 7704 -15699 7710 -15665
rect 7664 -15737 7710 -15699
rect 7664 -15771 7670 -15737
rect 7704 -15771 7710 -15737
rect 7664 -15809 7710 -15771
rect 7664 -15843 7670 -15809
rect 7704 -15843 7710 -15809
rect 7664 -15881 7710 -15843
rect 7664 -15915 7670 -15881
rect 7704 -15915 7710 -15881
rect 7664 -15953 7710 -15915
rect 7664 -15956 7670 -15953
rect 6646 -16018 6692 -15987
rect 7656 -15987 7670 -15956
rect 7704 -15956 7710 -15953
rect 8682 -15483 8688 -15449
rect 8722 -15483 8728 -15449
rect 8682 -15521 8728 -15483
rect 9696 -15449 9756 -15176
rect 9988 -15346 10476 -15340
rect 9988 -15380 10035 -15346
rect 10069 -15380 10107 -15346
rect 10141 -15380 10179 -15346
rect 10213 -15380 10251 -15346
rect 10285 -15380 10323 -15346
rect 10357 -15380 10395 -15346
rect 10429 -15380 10476 -15346
rect 9988 -15386 10476 -15380
rect 11006 -15346 11494 -15340
rect 11006 -15380 11053 -15346
rect 11087 -15380 11125 -15346
rect 11159 -15380 11197 -15346
rect 11231 -15380 11269 -15346
rect 11303 -15380 11341 -15346
rect 11375 -15380 11413 -15346
rect 11447 -15380 11494 -15346
rect 11006 -15386 11494 -15380
rect 9696 -15483 9706 -15449
rect 9740 -15483 9756 -15449
rect 9696 -15486 9756 -15483
rect 10718 -15449 10764 -15418
rect 10718 -15483 10724 -15449
rect 10758 -15483 10764 -15449
rect 11730 -15449 11790 -15176
rect 12024 -15346 12512 -15340
rect 12024 -15380 12071 -15346
rect 12105 -15380 12143 -15346
rect 12177 -15380 12215 -15346
rect 12249 -15380 12287 -15346
rect 12321 -15380 12359 -15346
rect 12393 -15380 12431 -15346
rect 12465 -15380 12512 -15346
rect 12024 -15386 12512 -15380
rect 13042 -15346 13530 -15340
rect 13042 -15380 13089 -15346
rect 13123 -15380 13161 -15346
rect 13195 -15380 13233 -15346
rect 13267 -15380 13305 -15346
rect 13339 -15380 13377 -15346
rect 13411 -15380 13449 -15346
rect 13483 -15380 13530 -15346
rect 13042 -15386 13530 -15380
rect 11730 -15480 11742 -15449
rect 8682 -15555 8688 -15521
rect 8722 -15555 8728 -15521
rect 8682 -15593 8728 -15555
rect 8682 -15627 8688 -15593
rect 8722 -15627 8728 -15593
rect 8682 -15665 8728 -15627
rect 8682 -15699 8688 -15665
rect 8722 -15699 8728 -15665
rect 8682 -15737 8728 -15699
rect 8682 -15771 8688 -15737
rect 8722 -15771 8728 -15737
rect 8682 -15809 8728 -15771
rect 8682 -15843 8688 -15809
rect 8722 -15843 8728 -15809
rect 8682 -15881 8728 -15843
rect 8682 -15915 8688 -15881
rect 8722 -15915 8728 -15881
rect 8682 -15953 8728 -15915
rect 7704 -15987 7716 -15956
rect 8682 -15970 8688 -15953
rect 5916 -16056 6404 -16050
rect 5916 -16090 5963 -16056
rect 5997 -16090 6035 -16056
rect 6069 -16090 6107 -16056
rect 6141 -16090 6179 -16056
rect 6213 -16090 6251 -16056
rect 6285 -16090 6323 -16056
rect 6357 -16090 6404 -16056
rect 5916 -16096 6404 -16090
rect 6934 -16056 7422 -16050
rect 6934 -16090 6981 -16056
rect 7015 -16090 7053 -16056
rect 7087 -16090 7125 -16056
rect 7159 -16090 7197 -16056
rect 7231 -16090 7269 -16056
rect 7303 -16090 7341 -16056
rect 7375 -16090 7422 -16056
rect 6934 -16096 7422 -16090
rect 5614 -16138 5686 -16134
rect 5614 -16190 5624 -16138
rect 5676 -16190 5686 -16138
rect 5614 -16194 5686 -16190
rect 5110 -16356 5182 -16352
rect 5110 -16408 5120 -16356
rect 5172 -16408 5182 -16356
rect 5110 -16412 5182 -16408
rect 5116 -16574 5176 -16412
rect 4898 -16580 5386 -16574
rect 4898 -16614 4945 -16580
rect 4979 -16614 5017 -16580
rect 5051 -16614 5089 -16580
rect 5123 -16614 5161 -16580
rect 5195 -16614 5233 -16580
rect 5267 -16614 5305 -16580
rect 5339 -16614 5386 -16580
rect 4898 -16620 5386 -16614
rect 3632 -16717 3638 -16700
rect 4602 -16706 4616 -16683
rect 3592 -16755 3638 -16717
rect 3592 -16789 3598 -16755
rect 3632 -16789 3638 -16755
rect 3592 -16827 3638 -16789
rect 3592 -16861 3598 -16827
rect 3632 -16861 3638 -16827
rect 3592 -16899 3638 -16861
rect 3592 -16933 3598 -16899
rect 3632 -16933 3638 -16899
rect 3592 -16971 3638 -16933
rect 3592 -17005 3598 -16971
rect 3632 -17005 3638 -16971
rect 3592 -17043 3638 -17005
rect 3592 -17077 3598 -17043
rect 3632 -17077 3638 -17043
rect 3592 -17115 3638 -17077
rect 3592 -17149 3598 -17115
rect 3632 -17149 3638 -17115
rect 3592 -17187 3638 -17149
rect 4610 -16717 4616 -16706
rect 4650 -16706 4662 -16683
rect 5620 -16683 5680 -16194
rect 6118 -16346 6178 -16096
rect 6636 -16242 6708 -16238
rect 6636 -16294 6646 -16242
rect 6698 -16294 6708 -16242
rect 6636 -16298 6708 -16294
rect 6118 -16356 6180 -16346
rect 6118 -16408 6124 -16356
rect 6176 -16408 6180 -16356
rect 6118 -16418 6180 -16408
rect 6118 -16574 6178 -16418
rect 5916 -16580 6404 -16574
rect 5916 -16614 5963 -16580
rect 5997 -16614 6035 -16580
rect 6069 -16614 6107 -16580
rect 6141 -16614 6179 -16580
rect 6213 -16614 6251 -16580
rect 6285 -16614 6323 -16580
rect 6357 -16614 6404 -16580
rect 5916 -16620 6404 -16614
rect 4650 -16717 4656 -16706
rect 5620 -16708 5634 -16683
rect 4610 -16755 4656 -16717
rect 4610 -16789 4616 -16755
rect 4650 -16789 4656 -16755
rect 4610 -16827 4656 -16789
rect 4610 -16861 4616 -16827
rect 4650 -16861 4656 -16827
rect 4610 -16899 4656 -16861
rect 4610 -16933 4616 -16899
rect 4650 -16933 4656 -16899
rect 4610 -16971 4656 -16933
rect 4610 -17005 4616 -16971
rect 4650 -17005 4656 -16971
rect 4610 -17043 4656 -17005
rect 4610 -17077 4616 -17043
rect 4650 -17077 4656 -17043
rect 4610 -17115 4656 -17077
rect 4610 -17149 4616 -17115
rect 4650 -17149 4656 -17115
rect 4610 -17182 4656 -17149
rect 5628 -16717 5634 -16708
rect 5668 -16708 5680 -16683
rect 6642 -16683 6702 -16298
rect 7134 -16346 7194 -16096
rect 7656 -16134 7716 -15987
rect 8674 -15987 8688 -15970
rect 8722 -15970 8728 -15953
rect 9700 -15521 9746 -15486
rect 9700 -15555 9706 -15521
rect 9740 -15555 9746 -15521
rect 9700 -15593 9746 -15555
rect 9700 -15627 9706 -15593
rect 9740 -15627 9746 -15593
rect 9700 -15665 9746 -15627
rect 9700 -15699 9706 -15665
rect 9740 -15699 9746 -15665
rect 9700 -15737 9746 -15699
rect 9700 -15771 9706 -15737
rect 9740 -15771 9746 -15737
rect 9700 -15809 9746 -15771
rect 9700 -15843 9706 -15809
rect 9740 -15843 9746 -15809
rect 9700 -15881 9746 -15843
rect 9700 -15915 9706 -15881
rect 9740 -15915 9746 -15881
rect 9700 -15953 9746 -15915
rect 8722 -15987 8734 -15970
rect 7952 -16056 8440 -16050
rect 7952 -16090 7999 -16056
rect 8033 -16090 8071 -16056
rect 8105 -16090 8143 -16056
rect 8177 -16090 8215 -16056
rect 8249 -16090 8287 -16056
rect 8321 -16090 8359 -16056
rect 8393 -16090 8440 -16056
rect 7952 -16096 8440 -16090
rect 7650 -16138 7722 -16134
rect 7650 -16190 7660 -16138
rect 7712 -16190 7722 -16138
rect 7650 -16194 7722 -16190
rect 7132 -16356 7194 -16346
rect 7132 -16408 7136 -16356
rect 7188 -16408 7194 -16356
rect 7132 -16418 7194 -16408
rect 7134 -16574 7194 -16418
rect 6934 -16580 7422 -16574
rect 6934 -16614 6981 -16580
rect 7015 -16614 7053 -16580
rect 7087 -16614 7125 -16580
rect 7159 -16614 7197 -16580
rect 7231 -16614 7269 -16580
rect 7303 -16614 7341 -16580
rect 7375 -16614 7422 -16580
rect 6934 -16620 7422 -16614
rect 6642 -16706 6652 -16683
rect 5668 -16717 5674 -16708
rect 5628 -16755 5674 -16717
rect 5628 -16789 5634 -16755
rect 5668 -16789 5674 -16755
rect 5628 -16827 5674 -16789
rect 5628 -16861 5634 -16827
rect 5668 -16861 5674 -16827
rect 5628 -16899 5674 -16861
rect 5628 -16933 5634 -16899
rect 5668 -16933 5674 -16899
rect 5628 -16971 5674 -16933
rect 5628 -17005 5634 -16971
rect 5668 -17005 5674 -16971
rect 5628 -17043 5674 -17005
rect 5628 -17077 5634 -17043
rect 5668 -17077 5674 -17043
rect 5628 -17115 5674 -17077
rect 5628 -17149 5634 -17115
rect 5668 -17149 5674 -17115
rect 3592 -17221 3598 -17187
rect 3632 -17221 3638 -17187
rect 3592 -17252 3638 -17221
rect 4604 -17187 4664 -17182
rect 4604 -17221 4616 -17187
rect 4650 -17221 4664 -17187
rect 5628 -17187 5674 -17149
rect 5628 -17192 5634 -17187
rect 2862 -17290 3350 -17284
rect 2862 -17324 2909 -17290
rect 2943 -17324 2981 -17290
rect 3015 -17324 3053 -17290
rect 3087 -17324 3125 -17290
rect 3159 -17324 3197 -17290
rect 3231 -17324 3269 -17290
rect 3303 -17324 3350 -17290
rect 2862 -17330 3350 -17324
rect 3880 -17290 4368 -17284
rect 3880 -17324 3927 -17290
rect 3961 -17324 3999 -17290
rect 4033 -17324 4071 -17290
rect 4105 -17324 4143 -17290
rect 4177 -17324 4215 -17290
rect 4249 -17324 4287 -17290
rect 4321 -17324 4368 -17290
rect 3880 -17330 4368 -17324
rect 3578 -17394 3650 -17390
rect 3578 -17446 3588 -17394
rect 3640 -17446 3650 -17394
rect 3578 -17450 3650 -17446
rect 2862 -17812 3350 -17806
rect 2862 -17846 2909 -17812
rect 2943 -17846 2981 -17812
rect 3015 -17846 3053 -17812
rect 3087 -17846 3125 -17812
rect 3159 -17846 3197 -17812
rect 3231 -17846 3269 -17812
rect 3303 -17846 3350 -17812
rect 2862 -17852 3350 -17846
rect 2574 -17915 2620 -17884
rect 2574 -17949 2580 -17915
rect 2614 -17949 2620 -17915
rect 3584 -17915 3644 -17450
rect 4090 -17492 4150 -17330
rect 4084 -17496 4156 -17492
rect 4084 -17548 4094 -17496
rect 4146 -17548 4156 -17496
rect 4084 -17552 4156 -17548
rect 4604 -17694 4664 -17221
rect 5622 -17221 5634 -17192
rect 5668 -17192 5674 -17187
rect 6646 -16717 6652 -16706
rect 6686 -16706 6702 -16683
rect 7656 -16683 7716 -16194
rect 8152 -16356 8212 -16096
rect 8674 -16238 8734 -15987
rect 9700 -15987 9706 -15953
rect 9740 -15987 9746 -15953
rect 10718 -15521 10764 -15483
rect 10718 -15555 10724 -15521
rect 10758 -15555 10764 -15521
rect 10718 -15593 10764 -15555
rect 10718 -15627 10724 -15593
rect 10758 -15627 10764 -15593
rect 10718 -15665 10764 -15627
rect 10718 -15699 10724 -15665
rect 10758 -15699 10764 -15665
rect 10718 -15737 10764 -15699
rect 10718 -15771 10724 -15737
rect 10758 -15771 10764 -15737
rect 10718 -15809 10764 -15771
rect 10718 -15843 10724 -15809
rect 10758 -15843 10764 -15809
rect 10718 -15881 10764 -15843
rect 10718 -15915 10724 -15881
rect 10758 -15915 10764 -15881
rect 10718 -15953 10764 -15915
rect 10718 -15976 10724 -15953
rect 9700 -16018 9746 -15987
rect 10708 -15987 10724 -15976
rect 10758 -15976 10764 -15953
rect 11736 -15483 11742 -15480
rect 11776 -15480 11790 -15449
rect 12754 -15449 12800 -15418
rect 11776 -15483 11782 -15480
rect 11736 -15521 11782 -15483
rect 11736 -15555 11742 -15521
rect 11776 -15555 11782 -15521
rect 11736 -15593 11782 -15555
rect 11736 -15627 11742 -15593
rect 11776 -15627 11782 -15593
rect 11736 -15665 11782 -15627
rect 11736 -15699 11742 -15665
rect 11776 -15699 11782 -15665
rect 11736 -15737 11782 -15699
rect 11736 -15771 11742 -15737
rect 11776 -15771 11782 -15737
rect 11736 -15809 11782 -15771
rect 11736 -15843 11742 -15809
rect 11776 -15843 11782 -15809
rect 11736 -15881 11782 -15843
rect 11736 -15915 11742 -15881
rect 11776 -15915 11782 -15881
rect 11736 -15953 11782 -15915
rect 10758 -15987 10768 -15976
rect 8970 -16056 9458 -16050
rect 8970 -16090 9017 -16056
rect 9051 -16090 9089 -16056
rect 9123 -16090 9161 -16056
rect 9195 -16090 9233 -16056
rect 9267 -16090 9305 -16056
rect 9339 -16090 9377 -16056
rect 9411 -16090 9458 -16056
rect 8970 -16096 9458 -16090
rect 9988 -16056 10476 -16050
rect 9988 -16090 10035 -16056
rect 10069 -16090 10107 -16056
rect 10141 -16090 10179 -16056
rect 10213 -16090 10251 -16056
rect 10285 -16090 10323 -16056
rect 10357 -16090 10395 -16056
rect 10429 -16090 10476 -16056
rect 9988 -16096 10476 -16090
rect 8668 -16242 8740 -16238
rect 8668 -16294 8678 -16242
rect 8730 -16294 8740 -16242
rect 8668 -16298 8740 -16294
rect 9164 -16294 9224 -16096
rect 10206 -16294 10266 -16096
rect 10708 -16238 10768 -15987
rect 11736 -15987 11742 -15953
rect 11776 -15987 11782 -15953
rect 12754 -15483 12760 -15449
rect 12794 -15483 12800 -15449
rect 13760 -15449 13820 -15176
rect 15304 -15340 15364 -14964
rect 15794 -14998 15866 -14994
rect 15794 -15050 15804 -14998
rect 15856 -15050 15866 -14998
rect 15794 -15054 15866 -15050
rect 14060 -15346 14548 -15340
rect 14060 -15380 14107 -15346
rect 14141 -15380 14179 -15346
rect 14213 -15380 14251 -15346
rect 14285 -15380 14323 -15346
rect 14357 -15380 14395 -15346
rect 14429 -15380 14467 -15346
rect 14501 -15380 14548 -15346
rect 14060 -15386 14548 -15380
rect 15078 -15346 15566 -15340
rect 15078 -15380 15125 -15346
rect 15159 -15380 15197 -15346
rect 15231 -15380 15269 -15346
rect 15303 -15380 15341 -15346
rect 15375 -15380 15413 -15346
rect 15447 -15380 15485 -15346
rect 15519 -15380 15566 -15346
rect 15078 -15386 15566 -15380
rect 13760 -15474 13778 -15449
rect 12754 -15521 12800 -15483
rect 12754 -15555 12760 -15521
rect 12794 -15555 12800 -15521
rect 12754 -15593 12800 -15555
rect 12754 -15627 12760 -15593
rect 12794 -15627 12800 -15593
rect 12754 -15665 12800 -15627
rect 12754 -15699 12760 -15665
rect 12794 -15699 12800 -15665
rect 12754 -15737 12800 -15699
rect 12754 -15771 12760 -15737
rect 12794 -15771 12800 -15737
rect 12754 -15809 12800 -15771
rect 12754 -15843 12760 -15809
rect 12794 -15843 12800 -15809
rect 12754 -15881 12800 -15843
rect 12754 -15915 12760 -15881
rect 12794 -15915 12800 -15881
rect 12754 -15953 12800 -15915
rect 12754 -15964 12760 -15953
rect 11736 -16018 11782 -15987
rect 12748 -15987 12760 -15964
rect 12794 -15964 12800 -15953
rect 13772 -15483 13778 -15474
rect 13812 -15474 13820 -15449
rect 14790 -15449 14836 -15418
rect 13812 -15483 13818 -15474
rect 13772 -15521 13818 -15483
rect 13772 -15555 13778 -15521
rect 13812 -15555 13818 -15521
rect 13772 -15593 13818 -15555
rect 13772 -15627 13778 -15593
rect 13812 -15627 13818 -15593
rect 13772 -15665 13818 -15627
rect 13772 -15699 13778 -15665
rect 13812 -15699 13818 -15665
rect 13772 -15737 13818 -15699
rect 13772 -15771 13778 -15737
rect 13812 -15771 13818 -15737
rect 13772 -15809 13818 -15771
rect 13772 -15843 13778 -15809
rect 13812 -15843 13818 -15809
rect 13772 -15881 13818 -15843
rect 13772 -15915 13778 -15881
rect 13812 -15915 13818 -15881
rect 13772 -15953 13818 -15915
rect 12794 -15987 12808 -15964
rect 11006 -16056 11494 -16050
rect 11006 -16090 11053 -16056
rect 11087 -16090 11125 -16056
rect 11159 -16090 11197 -16056
rect 11231 -16090 11269 -16056
rect 11303 -16090 11341 -16056
rect 11375 -16090 11413 -16056
rect 11447 -16090 11494 -16056
rect 11006 -16096 11494 -16090
rect 12024 -16056 12512 -16050
rect 12024 -16090 12071 -16056
rect 12105 -16090 12143 -16056
rect 12177 -16090 12215 -16056
rect 12249 -16090 12287 -16056
rect 12321 -16090 12359 -16056
rect 12393 -16090 12431 -16056
rect 12465 -16090 12512 -16056
rect 12024 -16096 12512 -16090
rect 8152 -16408 8156 -16356
rect 8208 -16408 8212 -16356
rect 8152 -16574 8212 -16408
rect 8668 -16354 8740 -16350
rect 8668 -16406 8678 -16354
rect 8730 -16406 8740 -16354
rect 8668 -16410 8740 -16406
rect 9164 -16354 10266 -16294
rect 10702 -16242 10774 -16238
rect 10702 -16294 10712 -16242
rect 10764 -16294 10774 -16242
rect 10702 -16298 10774 -16294
rect 7952 -16580 8440 -16574
rect 7952 -16614 7999 -16580
rect 8033 -16614 8071 -16580
rect 8105 -16614 8143 -16580
rect 8177 -16614 8215 -16580
rect 8249 -16614 8287 -16580
rect 8321 -16614 8359 -16580
rect 8393 -16614 8440 -16580
rect 7952 -16620 8440 -16614
rect 6686 -16717 6692 -16706
rect 7656 -16712 7670 -16683
rect 6646 -16755 6692 -16717
rect 6646 -16789 6652 -16755
rect 6686 -16789 6692 -16755
rect 6646 -16827 6692 -16789
rect 6646 -16861 6652 -16827
rect 6686 -16861 6692 -16827
rect 6646 -16899 6692 -16861
rect 6646 -16933 6652 -16899
rect 6686 -16933 6692 -16899
rect 6646 -16971 6692 -16933
rect 6646 -17005 6652 -16971
rect 6686 -17005 6692 -16971
rect 6646 -17043 6692 -17005
rect 6646 -17077 6652 -17043
rect 6686 -17077 6692 -17043
rect 6646 -17115 6692 -17077
rect 6646 -17149 6652 -17115
rect 6686 -17149 6692 -17115
rect 6646 -17187 6692 -17149
rect 5668 -17221 5682 -17192
rect 4898 -17290 5386 -17284
rect 4898 -17324 4945 -17290
rect 4979 -17324 5017 -17290
rect 5051 -17324 5089 -17290
rect 5123 -17324 5161 -17290
rect 5195 -17324 5233 -17290
rect 5267 -17324 5305 -17290
rect 5339 -17324 5386 -17290
rect 4898 -17330 5386 -17324
rect 5622 -17390 5682 -17221
rect 6646 -17221 6652 -17187
rect 6686 -17221 6692 -17187
rect 7664 -16717 7670 -16712
rect 7704 -16712 7716 -16683
rect 8674 -16683 8734 -16410
rect 9164 -16574 9224 -16354
rect 9686 -16464 9758 -16460
rect 9686 -16516 9696 -16464
rect 9748 -16516 9758 -16464
rect 9686 -16520 9758 -16516
rect 8970 -16580 9458 -16574
rect 8970 -16614 9017 -16580
rect 9051 -16614 9089 -16580
rect 9123 -16614 9161 -16580
rect 9195 -16614 9233 -16580
rect 9267 -16614 9305 -16580
rect 9339 -16614 9377 -16580
rect 9411 -16614 9458 -16580
rect 8970 -16620 9458 -16614
rect 7704 -16717 7710 -16712
rect 7664 -16755 7710 -16717
rect 8674 -16717 8688 -16683
rect 8722 -16717 8734 -16683
rect 9692 -16683 9752 -16520
rect 10206 -16574 10266 -16354
rect 10704 -16354 10776 -16350
rect 10704 -16406 10714 -16354
rect 10766 -16406 10776 -16354
rect 10704 -16410 10776 -16406
rect 9988 -16580 10476 -16574
rect 9988 -16614 10035 -16580
rect 10069 -16614 10107 -16580
rect 10141 -16614 10179 -16580
rect 10213 -16614 10251 -16580
rect 10285 -16614 10323 -16580
rect 10357 -16614 10395 -16580
rect 10429 -16614 10476 -16580
rect 9988 -16620 10476 -16614
rect 9692 -16710 9706 -16683
rect 8674 -16722 8734 -16717
rect 9700 -16717 9706 -16710
rect 9740 -16710 9752 -16683
rect 10710 -16683 10770 -16410
rect 11206 -16574 11266 -16096
rect 11720 -16464 11792 -16460
rect 11720 -16516 11730 -16464
rect 11782 -16516 11792 -16464
rect 11720 -16520 11792 -16516
rect 11006 -16580 11494 -16574
rect 11006 -16614 11053 -16580
rect 11087 -16614 11125 -16580
rect 11159 -16614 11197 -16580
rect 11231 -16614 11269 -16580
rect 11303 -16614 11341 -16580
rect 11375 -16614 11413 -16580
rect 11447 -16614 11494 -16580
rect 11006 -16620 11494 -16614
rect 9740 -16717 9746 -16710
rect 7664 -16789 7670 -16755
rect 7704 -16789 7710 -16755
rect 7664 -16827 7710 -16789
rect 7664 -16861 7670 -16827
rect 7704 -16861 7710 -16827
rect 7664 -16899 7710 -16861
rect 7664 -16933 7670 -16899
rect 7704 -16933 7710 -16899
rect 7664 -16971 7710 -16933
rect 7664 -17005 7670 -16971
rect 7704 -17005 7710 -16971
rect 7664 -17043 7710 -17005
rect 7664 -17077 7670 -17043
rect 7704 -17077 7710 -17043
rect 7664 -17115 7710 -17077
rect 7664 -17149 7670 -17115
rect 7704 -17149 7710 -17115
rect 7664 -17187 7710 -17149
rect 7664 -17190 7670 -17187
rect 6646 -17252 6692 -17221
rect 7658 -17221 7670 -17190
rect 7704 -17190 7710 -17187
rect 8682 -16755 8728 -16722
rect 8682 -16789 8688 -16755
rect 8722 -16789 8728 -16755
rect 8682 -16827 8728 -16789
rect 8682 -16861 8688 -16827
rect 8722 -16861 8728 -16827
rect 8682 -16899 8728 -16861
rect 8682 -16933 8688 -16899
rect 8722 -16933 8728 -16899
rect 8682 -16971 8728 -16933
rect 8682 -17005 8688 -16971
rect 8722 -17005 8728 -16971
rect 8682 -17043 8728 -17005
rect 8682 -17077 8688 -17043
rect 8722 -17077 8728 -17043
rect 8682 -17115 8728 -17077
rect 8682 -17149 8688 -17115
rect 8722 -17149 8728 -17115
rect 8682 -17187 8728 -17149
rect 7704 -17221 7718 -17190
rect 5916 -17290 6404 -17284
rect 5916 -17324 5963 -17290
rect 5997 -17324 6035 -17290
rect 6069 -17324 6107 -17290
rect 6141 -17324 6179 -17290
rect 6213 -17324 6251 -17290
rect 6285 -17324 6323 -17290
rect 6357 -17324 6404 -17290
rect 5916 -17330 6404 -17324
rect 6934 -17290 7422 -17284
rect 6934 -17324 6981 -17290
rect 7015 -17324 7053 -17290
rect 7087 -17324 7125 -17290
rect 7159 -17324 7197 -17290
rect 7231 -17324 7269 -17290
rect 7303 -17324 7341 -17290
rect 7375 -17324 7422 -17290
rect 6934 -17330 7422 -17324
rect 5616 -17394 5688 -17390
rect 5616 -17446 5626 -17394
rect 5678 -17446 5688 -17394
rect 5616 -17450 5688 -17446
rect 5614 -17598 5686 -17594
rect 5614 -17650 5624 -17598
rect 5676 -17650 5686 -17598
rect 6128 -17600 6188 -17330
rect 7150 -17600 7210 -17330
rect 7658 -17390 7718 -17221
rect 8682 -17221 8688 -17187
rect 8722 -17221 8728 -17187
rect 8682 -17252 8728 -17221
rect 9700 -16755 9746 -16717
rect 10710 -16717 10724 -16683
rect 10758 -16717 10770 -16683
rect 11726 -16683 11786 -16520
rect 12240 -16574 12300 -16096
rect 12748 -16238 12808 -15987
rect 13772 -15987 13778 -15953
rect 13812 -15987 13818 -15953
rect 14790 -15483 14796 -15449
rect 14830 -15483 14836 -15449
rect 15800 -15449 15860 -15054
rect 16306 -15170 16366 -14964
rect 16818 -14994 16878 -14753
rect 17846 -14249 17852 -14238
rect 17886 -14238 17898 -14215
rect 18856 -14215 18916 -13738
rect 20378 -13792 20450 -13788
rect 20378 -13844 20388 -13792
rect 20440 -13844 20450 -13792
rect 20378 -13848 20450 -13844
rect 21398 -13792 21470 -13788
rect 21398 -13844 21408 -13792
rect 21460 -13844 21470 -13792
rect 21398 -13848 21470 -13844
rect 19346 -13896 19418 -13892
rect 19346 -13948 19356 -13896
rect 19408 -13948 19418 -13896
rect 19346 -13952 19418 -13948
rect 19352 -14106 19412 -13952
rect 19864 -14004 19936 -14000
rect 19864 -14056 19874 -14004
rect 19926 -14056 19936 -14004
rect 19864 -14060 19936 -14056
rect 19152 -14112 19640 -14106
rect 19152 -14146 19199 -14112
rect 19233 -14146 19271 -14112
rect 19305 -14146 19343 -14112
rect 19377 -14146 19415 -14112
rect 19449 -14146 19487 -14112
rect 19521 -14146 19559 -14112
rect 19593 -14146 19640 -14112
rect 19152 -14152 19640 -14146
rect 19352 -14164 19412 -14152
rect 17886 -14249 17892 -14238
rect 17846 -14287 17892 -14249
rect 18856 -14249 18870 -14215
rect 18904 -14249 18916 -14215
rect 19870 -14215 19930 -14060
rect 20384 -14106 20444 -13848
rect 21404 -14106 21464 -13848
rect 21906 -14004 21978 -14000
rect 21906 -14056 21916 -14004
rect 21968 -14056 21978 -14004
rect 21906 -14060 21978 -14056
rect 22410 -14004 22482 -14000
rect 22410 -14056 22420 -14004
rect 22472 -14056 22482 -14004
rect 22410 -14060 22482 -14056
rect 22920 -14004 22992 -14000
rect 22920 -14056 22930 -14004
rect 22982 -14056 22992 -14004
rect 22920 -14060 22992 -14056
rect 20170 -14112 20658 -14106
rect 20170 -14146 20217 -14112
rect 20251 -14146 20289 -14112
rect 20323 -14146 20361 -14112
rect 20395 -14146 20433 -14112
rect 20467 -14146 20505 -14112
rect 20539 -14146 20577 -14112
rect 20611 -14146 20658 -14112
rect 20170 -14152 20658 -14146
rect 21188 -14112 21676 -14106
rect 21188 -14146 21235 -14112
rect 21269 -14146 21307 -14112
rect 21341 -14146 21379 -14112
rect 21413 -14146 21451 -14112
rect 21485 -14146 21523 -14112
rect 21557 -14146 21595 -14112
rect 21629 -14146 21676 -14112
rect 21188 -14152 21676 -14146
rect 19870 -14242 19888 -14215
rect 18856 -14254 18916 -14249
rect 19882 -14249 19888 -14242
rect 19922 -14242 19930 -14215
rect 20900 -14215 20946 -14184
rect 19922 -14249 19928 -14242
rect 17846 -14321 17852 -14287
rect 17886 -14321 17892 -14287
rect 17846 -14359 17892 -14321
rect 17846 -14393 17852 -14359
rect 17886 -14393 17892 -14359
rect 17846 -14431 17892 -14393
rect 17846 -14465 17852 -14431
rect 17886 -14465 17892 -14431
rect 17846 -14503 17892 -14465
rect 17846 -14537 17852 -14503
rect 17886 -14537 17892 -14503
rect 17846 -14575 17892 -14537
rect 17846 -14609 17852 -14575
rect 17886 -14609 17892 -14575
rect 17846 -14647 17892 -14609
rect 17846 -14681 17852 -14647
rect 17886 -14681 17892 -14647
rect 17846 -14719 17892 -14681
rect 17846 -14753 17852 -14719
rect 17886 -14753 17892 -14719
rect 18864 -14287 18910 -14254
rect 18864 -14321 18870 -14287
rect 18904 -14321 18910 -14287
rect 18864 -14359 18910 -14321
rect 18864 -14393 18870 -14359
rect 18904 -14393 18910 -14359
rect 18864 -14431 18910 -14393
rect 18864 -14465 18870 -14431
rect 18904 -14465 18910 -14431
rect 18864 -14503 18910 -14465
rect 18864 -14537 18870 -14503
rect 18904 -14537 18910 -14503
rect 18864 -14575 18910 -14537
rect 18864 -14609 18870 -14575
rect 18904 -14609 18910 -14575
rect 18864 -14647 18910 -14609
rect 18864 -14681 18870 -14647
rect 18904 -14681 18910 -14647
rect 18864 -14719 18910 -14681
rect 18864 -14724 18870 -14719
rect 17846 -14784 17892 -14753
rect 18854 -14753 18870 -14724
rect 18904 -14724 18910 -14719
rect 19882 -14287 19928 -14249
rect 19882 -14321 19888 -14287
rect 19922 -14321 19928 -14287
rect 19882 -14359 19928 -14321
rect 19882 -14393 19888 -14359
rect 19922 -14393 19928 -14359
rect 19882 -14431 19928 -14393
rect 19882 -14465 19888 -14431
rect 19922 -14465 19928 -14431
rect 19882 -14503 19928 -14465
rect 19882 -14537 19888 -14503
rect 19922 -14537 19928 -14503
rect 19882 -14575 19928 -14537
rect 19882 -14609 19888 -14575
rect 19922 -14609 19928 -14575
rect 19882 -14647 19928 -14609
rect 19882 -14681 19888 -14647
rect 19922 -14681 19928 -14647
rect 19882 -14719 19928 -14681
rect 20900 -14249 20906 -14215
rect 20940 -14249 20946 -14215
rect 20900 -14287 20946 -14249
rect 21912 -14215 21972 -14060
rect 22416 -14106 22476 -14060
rect 22206 -14112 22694 -14106
rect 22206 -14146 22253 -14112
rect 22287 -14146 22325 -14112
rect 22359 -14146 22397 -14112
rect 22431 -14146 22469 -14112
rect 22503 -14146 22541 -14112
rect 22575 -14146 22613 -14112
rect 22647 -14146 22694 -14112
rect 22206 -14152 22694 -14146
rect 21912 -14249 21924 -14215
rect 21958 -14249 21972 -14215
rect 22926 -14215 22986 -14060
rect 22926 -14232 22942 -14215
rect 21912 -14252 21972 -14249
rect 22936 -14249 22942 -14232
rect 22976 -14232 22986 -14215
rect 22976 -14249 22982 -14232
rect 20900 -14321 20906 -14287
rect 20940 -14321 20946 -14287
rect 20900 -14359 20946 -14321
rect 20900 -14393 20906 -14359
rect 20940 -14393 20946 -14359
rect 20900 -14431 20946 -14393
rect 20900 -14465 20906 -14431
rect 20940 -14465 20946 -14431
rect 20900 -14503 20946 -14465
rect 20900 -14537 20906 -14503
rect 20940 -14537 20946 -14503
rect 20900 -14575 20946 -14537
rect 20900 -14609 20906 -14575
rect 20940 -14609 20946 -14575
rect 20900 -14647 20946 -14609
rect 20900 -14681 20906 -14647
rect 20940 -14681 20946 -14647
rect 20900 -14714 20946 -14681
rect 21918 -14287 21964 -14252
rect 21918 -14321 21924 -14287
rect 21958 -14321 21964 -14287
rect 21918 -14359 21964 -14321
rect 21918 -14393 21924 -14359
rect 21958 -14393 21964 -14359
rect 21918 -14431 21964 -14393
rect 21918 -14465 21924 -14431
rect 21958 -14465 21964 -14431
rect 21918 -14503 21964 -14465
rect 21918 -14537 21924 -14503
rect 21958 -14537 21964 -14503
rect 21918 -14575 21964 -14537
rect 21918 -14609 21924 -14575
rect 21958 -14609 21964 -14575
rect 21918 -14647 21964 -14609
rect 21918 -14681 21924 -14647
rect 21958 -14681 21964 -14647
rect 18904 -14753 18914 -14724
rect 17116 -14822 17604 -14816
rect 17116 -14856 17163 -14822
rect 17197 -14856 17235 -14822
rect 17269 -14856 17379 -14822
rect 17413 -14856 17451 -14822
rect 17485 -14856 17523 -14822
rect 17557 -14856 17604 -14822
rect 17116 -14862 17604 -14856
rect 18134 -14822 18622 -14816
rect 18134 -14856 18181 -14822
rect 18215 -14856 18253 -14822
rect 18287 -14856 18469 -14822
rect 18503 -14856 18541 -14822
rect 18575 -14856 18622 -14822
rect 18134 -14862 18622 -14856
rect 17318 -14890 17378 -14862
rect 18352 -14890 18412 -14862
rect 17310 -14894 17382 -14890
rect 17310 -14946 17320 -14894
rect 17372 -14946 17382 -14894
rect 17310 -14950 17382 -14946
rect 18346 -14894 18418 -14890
rect 18346 -14946 18356 -14894
rect 18408 -14946 18418 -14894
rect 18346 -14950 18418 -14946
rect 16812 -14998 16884 -14994
rect 16812 -15050 16822 -14998
rect 16874 -15050 16884 -14998
rect 16812 -15054 16884 -15050
rect 17318 -15170 17378 -14950
rect 17832 -14998 17904 -14994
rect 17832 -15050 17842 -14998
rect 17894 -15050 17904 -14998
rect 17832 -15054 17904 -15050
rect 16306 -15230 17378 -15170
rect 16306 -15340 16366 -15230
rect 17318 -15340 17378 -15230
rect 16096 -15346 16584 -15340
rect 16096 -15380 16143 -15346
rect 16177 -15380 16215 -15346
rect 16249 -15380 16287 -15346
rect 16321 -15380 16359 -15346
rect 16393 -15380 16431 -15346
rect 16465 -15380 16503 -15346
rect 16537 -15380 16584 -15346
rect 16096 -15386 16584 -15380
rect 17114 -15346 17602 -15340
rect 17114 -15380 17161 -15346
rect 17195 -15380 17233 -15346
rect 17267 -15380 17305 -15346
rect 17339 -15380 17377 -15346
rect 17411 -15380 17449 -15346
rect 17483 -15380 17521 -15346
rect 17555 -15380 17602 -15346
rect 17114 -15386 17602 -15380
rect 15800 -15478 15814 -15449
rect 14790 -15521 14836 -15483
rect 14790 -15555 14796 -15521
rect 14830 -15555 14836 -15521
rect 14790 -15593 14836 -15555
rect 14790 -15627 14796 -15593
rect 14830 -15627 14836 -15593
rect 14790 -15665 14836 -15627
rect 14790 -15699 14796 -15665
rect 14830 -15699 14836 -15665
rect 14790 -15737 14836 -15699
rect 14790 -15771 14796 -15737
rect 14830 -15771 14836 -15737
rect 14790 -15809 14836 -15771
rect 14790 -15843 14796 -15809
rect 14830 -15843 14836 -15809
rect 14790 -15881 14836 -15843
rect 14790 -15915 14796 -15881
rect 14830 -15915 14836 -15881
rect 14790 -15953 14836 -15915
rect 14790 -15954 14796 -15953
rect 13772 -16018 13818 -15987
rect 14782 -15987 14796 -15954
rect 14830 -15954 14836 -15953
rect 15808 -15483 15814 -15478
rect 15848 -15478 15860 -15449
rect 16826 -15449 16872 -15418
rect 15848 -15483 15854 -15478
rect 15808 -15521 15854 -15483
rect 15808 -15555 15814 -15521
rect 15848 -15555 15854 -15521
rect 15808 -15593 15854 -15555
rect 15808 -15627 15814 -15593
rect 15848 -15627 15854 -15593
rect 15808 -15665 15854 -15627
rect 15808 -15699 15814 -15665
rect 15848 -15699 15854 -15665
rect 15808 -15737 15854 -15699
rect 15808 -15771 15814 -15737
rect 15848 -15771 15854 -15737
rect 15808 -15809 15854 -15771
rect 15808 -15843 15814 -15809
rect 15848 -15843 15854 -15809
rect 15808 -15881 15854 -15843
rect 15808 -15915 15814 -15881
rect 15848 -15915 15854 -15881
rect 15808 -15953 15854 -15915
rect 14830 -15987 14842 -15954
rect 15808 -15974 15814 -15953
rect 13042 -16056 13530 -16050
rect 13042 -16090 13089 -16056
rect 13123 -16090 13161 -16056
rect 13195 -16090 13233 -16056
rect 13267 -16090 13305 -16056
rect 13339 -16090 13377 -16056
rect 13411 -16090 13449 -16056
rect 13483 -16090 13530 -16056
rect 13042 -16096 13530 -16090
rect 14060 -16056 14548 -16050
rect 14060 -16090 14107 -16056
rect 14141 -16090 14179 -16056
rect 14213 -16090 14251 -16056
rect 14285 -16090 14323 -16056
rect 14357 -16090 14395 -16056
rect 14429 -16090 14467 -16056
rect 14501 -16090 14548 -16056
rect 14060 -16096 14548 -16090
rect 12742 -16242 12814 -16238
rect 12742 -16294 12752 -16242
rect 12804 -16294 12814 -16242
rect 12742 -16298 12814 -16294
rect 13262 -16294 13322 -16096
rect 14270 -16294 14330 -16096
rect 14782 -16238 14842 -15987
rect 15800 -15987 15814 -15974
rect 15848 -15974 15854 -15953
rect 16826 -15483 16832 -15449
rect 16866 -15483 16872 -15449
rect 16826 -15521 16872 -15483
rect 17838 -15449 17898 -15054
rect 18352 -15178 18412 -14950
rect 18854 -14994 18914 -14753
rect 19882 -14753 19888 -14719
rect 19922 -14753 19928 -14719
rect 19882 -14784 19928 -14753
rect 20890 -14719 20950 -14714
rect 20890 -14753 20906 -14719
rect 20940 -14753 20950 -14719
rect 19152 -14822 19640 -14816
rect 19152 -14856 19199 -14822
rect 19233 -14856 19271 -14822
rect 19305 -14856 19343 -14822
rect 19377 -14856 19415 -14822
rect 19449 -14856 19487 -14822
rect 19521 -14856 19559 -14822
rect 19593 -14856 19640 -14822
rect 19152 -14862 19640 -14856
rect 20170 -14822 20658 -14816
rect 20170 -14856 20217 -14822
rect 20251 -14856 20289 -14822
rect 20323 -14856 20361 -14822
rect 20395 -14856 20433 -14822
rect 20467 -14856 20505 -14822
rect 20539 -14856 20577 -14822
rect 20611 -14856 20658 -14822
rect 20170 -14862 20658 -14856
rect 19368 -14890 19428 -14862
rect 19362 -14894 19434 -14890
rect 19362 -14946 19372 -14894
rect 19424 -14946 19434 -14894
rect 19362 -14950 19434 -14946
rect 20890 -14994 20950 -14753
rect 21918 -14719 21964 -14681
rect 21918 -14753 21924 -14719
rect 21958 -14753 21964 -14719
rect 21918 -14784 21964 -14753
rect 22936 -14287 22982 -14249
rect 22936 -14321 22942 -14287
rect 22976 -14321 22982 -14287
rect 22936 -14359 22982 -14321
rect 22936 -14393 22942 -14359
rect 22976 -14393 22982 -14359
rect 22936 -14431 22982 -14393
rect 22936 -14465 22942 -14431
rect 22976 -14465 22982 -14431
rect 22936 -14503 22982 -14465
rect 22936 -14537 22942 -14503
rect 22976 -14537 22982 -14503
rect 22936 -14575 22982 -14537
rect 22936 -14609 22942 -14575
rect 22976 -14609 22982 -14575
rect 22936 -14647 22982 -14609
rect 22936 -14681 22942 -14647
rect 22976 -14681 22982 -14647
rect 22936 -14719 22982 -14681
rect 22936 -14753 22942 -14719
rect 22976 -14753 22982 -14719
rect 22936 -14784 22982 -14753
rect 21188 -14822 21676 -14816
rect 21188 -14856 21235 -14822
rect 21269 -14856 21307 -14822
rect 21341 -14856 21379 -14822
rect 21413 -14856 21451 -14822
rect 21485 -14856 21523 -14822
rect 21557 -14856 21595 -14822
rect 21629 -14856 21676 -14822
rect 21188 -14862 21676 -14856
rect 22206 -14822 22694 -14816
rect 22206 -14856 22253 -14822
rect 22287 -14856 22325 -14822
rect 22359 -14856 22397 -14822
rect 22431 -14856 22469 -14822
rect 22503 -14856 22541 -14822
rect 22575 -14856 22613 -14822
rect 22647 -14856 22694 -14822
rect 22206 -14862 22694 -14856
rect 18848 -14998 18920 -14994
rect 18848 -15050 18858 -14998
rect 18910 -15050 18920 -14998
rect 18848 -15054 18920 -15050
rect 20884 -14998 20956 -14994
rect 20884 -15050 20894 -14998
rect 20946 -15050 20956 -14998
rect 20884 -15054 20956 -15050
rect 18352 -15238 21440 -15178
rect 18352 -15340 18412 -15238
rect 21380 -15340 21440 -15238
rect 22418 -15264 22986 -15204
rect 22418 -15340 22478 -15264
rect 18132 -15346 18620 -15340
rect 18132 -15380 18179 -15346
rect 18213 -15380 18251 -15346
rect 18285 -15380 18323 -15346
rect 18357 -15380 18395 -15346
rect 18429 -15380 18467 -15346
rect 18501 -15380 18539 -15346
rect 18573 -15380 18620 -15346
rect 18132 -15386 18620 -15380
rect 19150 -15346 19638 -15340
rect 19150 -15380 19197 -15346
rect 19231 -15380 19269 -15346
rect 19303 -15380 19341 -15346
rect 19375 -15380 19413 -15346
rect 19447 -15380 19485 -15346
rect 19519 -15380 19557 -15346
rect 19591 -15380 19638 -15346
rect 19150 -15386 19638 -15380
rect 20168 -15346 20656 -15340
rect 20168 -15380 20215 -15346
rect 20249 -15380 20287 -15346
rect 20321 -15380 20359 -15346
rect 20393 -15380 20431 -15346
rect 20465 -15380 20503 -15346
rect 20537 -15380 20575 -15346
rect 20609 -15380 20656 -15346
rect 20168 -15386 20656 -15380
rect 21186 -15346 21674 -15340
rect 21186 -15380 21233 -15346
rect 21267 -15380 21305 -15346
rect 21339 -15380 21377 -15346
rect 21411 -15380 21449 -15346
rect 21483 -15380 21521 -15346
rect 21555 -15380 21593 -15346
rect 21627 -15380 21674 -15346
rect 21186 -15386 21674 -15380
rect 22204 -15346 22692 -15340
rect 22204 -15380 22251 -15346
rect 22285 -15380 22323 -15346
rect 22357 -15380 22395 -15346
rect 22429 -15380 22467 -15346
rect 22501 -15380 22539 -15346
rect 22573 -15380 22611 -15346
rect 22645 -15380 22692 -15346
rect 22204 -15386 22692 -15380
rect 17838 -15483 17850 -15449
rect 17884 -15483 17898 -15449
rect 17838 -15488 17898 -15483
rect 18862 -15449 18908 -15418
rect 18862 -15483 18868 -15449
rect 18902 -15483 18908 -15449
rect 16826 -15555 16832 -15521
rect 16866 -15555 16872 -15521
rect 16826 -15593 16872 -15555
rect 16826 -15627 16832 -15593
rect 16866 -15627 16872 -15593
rect 16826 -15665 16872 -15627
rect 16826 -15699 16832 -15665
rect 16866 -15699 16872 -15665
rect 16826 -15737 16872 -15699
rect 16826 -15771 16832 -15737
rect 16866 -15771 16872 -15737
rect 16826 -15809 16872 -15771
rect 16826 -15843 16832 -15809
rect 16866 -15843 16872 -15809
rect 16826 -15881 16872 -15843
rect 16826 -15915 16832 -15881
rect 16866 -15915 16872 -15881
rect 16826 -15953 16872 -15915
rect 16826 -15970 16832 -15953
rect 15848 -15987 15860 -15974
rect 15078 -16056 15566 -16050
rect 15078 -16090 15125 -16056
rect 15159 -16090 15197 -16056
rect 15231 -16090 15269 -16056
rect 15303 -16090 15341 -16056
rect 15375 -16090 15413 -16056
rect 15447 -16090 15485 -16056
rect 15519 -16090 15566 -16056
rect 15078 -16096 15566 -16090
rect 12740 -16354 12812 -16350
rect 12740 -16406 12750 -16354
rect 12802 -16406 12812 -16354
rect 12740 -16410 12812 -16406
rect 13262 -16354 14330 -16294
rect 14776 -16242 14848 -16238
rect 14776 -16294 14786 -16242
rect 14838 -16294 14848 -16242
rect 14776 -16298 14848 -16294
rect 14972 -16246 15044 -16242
rect 14972 -16298 14982 -16246
rect 15034 -16298 15044 -16246
rect 14972 -16302 15044 -16298
rect 12024 -16580 12512 -16574
rect 12024 -16614 12071 -16580
rect 12105 -16614 12143 -16580
rect 12177 -16614 12215 -16580
rect 12249 -16614 12287 -16580
rect 12321 -16614 12359 -16580
rect 12393 -16614 12431 -16580
rect 12465 -16614 12512 -16580
rect 12024 -16620 12512 -16614
rect 11726 -16712 11742 -16683
rect 10710 -16732 10770 -16717
rect 11736 -16717 11742 -16712
rect 11776 -16712 11786 -16683
rect 12746 -16683 12806 -16410
rect 13262 -16574 13322 -16354
rect 13760 -16464 13832 -16460
rect 13760 -16516 13770 -16464
rect 13822 -16516 13832 -16464
rect 13760 -16520 13832 -16516
rect 13042 -16580 13530 -16574
rect 13042 -16614 13089 -16580
rect 13123 -16614 13161 -16580
rect 13195 -16614 13233 -16580
rect 13267 -16614 13305 -16580
rect 13339 -16614 13377 -16580
rect 13411 -16614 13449 -16580
rect 13483 -16614 13530 -16580
rect 13042 -16620 13530 -16614
rect 11776 -16717 11782 -16712
rect 12746 -16714 12760 -16683
rect 9700 -16789 9706 -16755
rect 9740 -16789 9746 -16755
rect 9700 -16827 9746 -16789
rect 9700 -16861 9706 -16827
rect 9740 -16861 9746 -16827
rect 9700 -16899 9746 -16861
rect 9700 -16933 9706 -16899
rect 9740 -16933 9746 -16899
rect 9700 -16971 9746 -16933
rect 9700 -17005 9706 -16971
rect 9740 -17005 9746 -16971
rect 9700 -17043 9746 -17005
rect 9700 -17077 9706 -17043
rect 9740 -17077 9746 -17043
rect 9700 -17115 9746 -17077
rect 9700 -17149 9706 -17115
rect 9740 -17149 9746 -17115
rect 9700 -17187 9746 -17149
rect 9700 -17221 9706 -17187
rect 9740 -17221 9746 -17187
rect 9700 -17252 9746 -17221
rect 10718 -16755 10764 -16732
rect 10718 -16789 10724 -16755
rect 10758 -16789 10764 -16755
rect 10718 -16827 10764 -16789
rect 10718 -16861 10724 -16827
rect 10758 -16861 10764 -16827
rect 10718 -16899 10764 -16861
rect 10718 -16933 10724 -16899
rect 10758 -16933 10764 -16899
rect 10718 -16971 10764 -16933
rect 10718 -17005 10724 -16971
rect 10758 -17005 10764 -16971
rect 10718 -17043 10764 -17005
rect 10718 -17077 10724 -17043
rect 10758 -17077 10764 -17043
rect 10718 -17115 10764 -17077
rect 10718 -17149 10724 -17115
rect 10758 -17149 10764 -17115
rect 10718 -17187 10764 -17149
rect 10718 -17221 10724 -17187
rect 10758 -17221 10764 -17187
rect 10718 -17252 10764 -17221
rect 11736 -16755 11782 -16717
rect 11736 -16789 11742 -16755
rect 11776 -16789 11782 -16755
rect 11736 -16827 11782 -16789
rect 11736 -16861 11742 -16827
rect 11776 -16861 11782 -16827
rect 11736 -16899 11782 -16861
rect 11736 -16933 11742 -16899
rect 11776 -16933 11782 -16899
rect 11736 -16971 11782 -16933
rect 11736 -17005 11742 -16971
rect 11776 -17005 11782 -16971
rect 11736 -17043 11782 -17005
rect 11736 -17077 11742 -17043
rect 11776 -17077 11782 -17043
rect 11736 -17115 11782 -17077
rect 11736 -17149 11742 -17115
rect 11776 -17149 11782 -17115
rect 11736 -17187 11782 -17149
rect 11736 -17221 11742 -17187
rect 11776 -17221 11782 -17187
rect 11736 -17252 11782 -17221
rect 12754 -16717 12760 -16714
rect 12794 -16714 12806 -16683
rect 13766 -16683 13826 -16520
rect 14270 -16574 14330 -16354
rect 14776 -16354 14848 -16350
rect 14776 -16406 14786 -16354
rect 14838 -16406 14848 -16354
rect 14776 -16410 14848 -16406
rect 14060 -16580 14548 -16574
rect 14060 -16614 14107 -16580
rect 14141 -16614 14179 -16580
rect 14213 -16614 14251 -16580
rect 14285 -16614 14323 -16580
rect 14357 -16614 14395 -16580
rect 14429 -16614 14467 -16580
rect 14501 -16614 14548 -16580
rect 14060 -16620 14548 -16614
rect 13766 -16702 13778 -16683
rect 12794 -16717 12800 -16714
rect 12754 -16755 12800 -16717
rect 12754 -16789 12760 -16755
rect 12794 -16789 12800 -16755
rect 12754 -16827 12800 -16789
rect 12754 -16861 12760 -16827
rect 12794 -16861 12800 -16827
rect 12754 -16899 12800 -16861
rect 12754 -16933 12760 -16899
rect 12794 -16933 12800 -16899
rect 12754 -16971 12800 -16933
rect 12754 -17005 12760 -16971
rect 12794 -17005 12800 -16971
rect 12754 -17043 12800 -17005
rect 12754 -17077 12760 -17043
rect 12794 -17077 12800 -17043
rect 12754 -17115 12800 -17077
rect 12754 -17149 12760 -17115
rect 12794 -17149 12800 -17115
rect 12754 -17187 12800 -17149
rect 12754 -17221 12760 -17187
rect 12794 -17221 12800 -17187
rect 13772 -16717 13778 -16702
rect 13812 -16702 13826 -16683
rect 14782 -16683 14842 -16410
rect 14978 -16460 15038 -16302
rect 15272 -16458 15332 -16096
rect 15800 -16134 15860 -15987
rect 16816 -15987 16832 -15970
rect 16866 -15970 16872 -15953
rect 17844 -15521 17890 -15488
rect 17844 -15555 17850 -15521
rect 17884 -15555 17890 -15521
rect 17844 -15593 17890 -15555
rect 17844 -15627 17850 -15593
rect 17884 -15627 17890 -15593
rect 17844 -15665 17890 -15627
rect 17844 -15699 17850 -15665
rect 17884 -15699 17890 -15665
rect 17844 -15737 17890 -15699
rect 17844 -15771 17850 -15737
rect 17884 -15771 17890 -15737
rect 17844 -15809 17890 -15771
rect 17844 -15843 17850 -15809
rect 17884 -15843 17890 -15809
rect 17844 -15881 17890 -15843
rect 17844 -15915 17850 -15881
rect 17884 -15915 17890 -15881
rect 17844 -15953 17890 -15915
rect 18862 -15521 18908 -15483
rect 18862 -15555 18868 -15521
rect 18902 -15555 18908 -15521
rect 18862 -15593 18908 -15555
rect 18862 -15627 18868 -15593
rect 18902 -15627 18908 -15593
rect 18862 -15665 18908 -15627
rect 18862 -15699 18868 -15665
rect 18902 -15699 18908 -15665
rect 18862 -15737 18908 -15699
rect 18862 -15771 18868 -15737
rect 18902 -15771 18908 -15737
rect 18862 -15809 18908 -15771
rect 18862 -15843 18868 -15809
rect 18902 -15843 18908 -15809
rect 18862 -15881 18908 -15843
rect 18862 -15915 18868 -15881
rect 18902 -15915 18908 -15881
rect 18862 -15950 18908 -15915
rect 19880 -15449 19926 -15418
rect 19880 -15483 19886 -15449
rect 19920 -15483 19926 -15449
rect 19880 -15521 19926 -15483
rect 19880 -15555 19886 -15521
rect 19920 -15555 19926 -15521
rect 19880 -15593 19926 -15555
rect 19880 -15627 19886 -15593
rect 19920 -15627 19926 -15593
rect 19880 -15665 19926 -15627
rect 19880 -15699 19886 -15665
rect 19920 -15699 19926 -15665
rect 19880 -15737 19926 -15699
rect 19880 -15771 19886 -15737
rect 19920 -15771 19926 -15737
rect 19880 -15809 19926 -15771
rect 19880 -15843 19886 -15809
rect 19920 -15843 19926 -15809
rect 19880 -15881 19926 -15843
rect 19880 -15915 19886 -15881
rect 19920 -15915 19926 -15881
rect 17844 -15960 17850 -15953
rect 16866 -15987 16876 -15970
rect 16096 -16056 16584 -16050
rect 16096 -16090 16143 -16056
rect 16177 -16090 16215 -16056
rect 16249 -16090 16287 -16056
rect 16321 -16090 16359 -16056
rect 16393 -16090 16431 -16056
rect 16465 -16090 16503 -16056
rect 16537 -16090 16584 -16056
rect 16096 -16096 16584 -16090
rect 15794 -16138 15866 -16134
rect 15794 -16190 15804 -16138
rect 15856 -16190 15866 -16138
rect 15794 -16194 15866 -16190
rect 14972 -16464 15044 -16460
rect 14972 -16516 14982 -16464
rect 15034 -16516 15044 -16464
rect 14972 -16520 15044 -16516
rect 15266 -16462 15338 -16458
rect 15266 -16514 15276 -16462
rect 15328 -16514 15338 -16462
rect 15266 -16518 15338 -16514
rect 15272 -16574 15332 -16518
rect 15078 -16580 15566 -16574
rect 15078 -16614 15125 -16580
rect 15159 -16614 15197 -16580
rect 15231 -16614 15269 -16580
rect 15303 -16614 15341 -16580
rect 15375 -16614 15413 -16580
rect 15447 -16614 15485 -16580
rect 15519 -16614 15566 -16580
rect 15078 -16620 15566 -16614
rect 13812 -16717 13818 -16702
rect 14782 -16708 14796 -16683
rect 13772 -16755 13818 -16717
rect 13772 -16789 13778 -16755
rect 13812 -16789 13818 -16755
rect 13772 -16827 13818 -16789
rect 13772 -16861 13778 -16827
rect 13812 -16861 13818 -16827
rect 13772 -16899 13818 -16861
rect 13772 -16933 13778 -16899
rect 13812 -16933 13818 -16899
rect 13772 -16971 13818 -16933
rect 13772 -17005 13778 -16971
rect 13812 -17005 13818 -16971
rect 13772 -17043 13818 -17005
rect 13772 -17077 13778 -17043
rect 13812 -17077 13818 -17043
rect 13772 -17115 13818 -17077
rect 13772 -17149 13778 -17115
rect 13812 -17149 13818 -17115
rect 13772 -17187 13818 -17149
rect 13772 -17194 13778 -17187
rect 12754 -17252 12800 -17221
rect 13766 -17221 13778 -17194
rect 13812 -17194 13818 -17187
rect 14790 -16717 14796 -16708
rect 14830 -16708 14842 -16683
rect 15800 -16683 15860 -16194
rect 16302 -16452 16362 -16096
rect 16816 -16350 16876 -15987
rect 17836 -15987 17850 -15960
rect 17884 -15960 17890 -15953
rect 18854 -15953 18914 -15950
rect 17884 -15987 17896 -15960
rect 17114 -16056 17602 -16050
rect 17114 -16090 17161 -16056
rect 17195 -16090 17233 -16056
rect 17267 -16090 17305 -16056
rect 17339 -16090 17377 -16056
rect 17411 -16090 17449 -16056
rect 17483 -16090 17521 -16056
rect 17555 -16090 17602 -16056
rect 17114 -16096 17602 -16090
rect 16810 -16354 16882 -16350
rect 16810 -16406 16820 -16354
rect 16872 -16406 16882 -16354
rect 16810 -16410 16882 -16406
rect 16300 -16462 16362 -16452
rect 16300 -16514 16304 -16462
rect 16356 -16514 16362 -16462
rect 16300 -16524 16362 -16514
rect 16812 -16468 16884 -16464
rect 16812 -16520 16822 -16468
rect 16874 -16520 16884 -16468
rect 16812 -16524 16884 -16520
rect 16302 -16574 16362 -16524
rect 16096 -16580 16584 -16574
rect 16096 -16614 16143 -16580
rect 16177 -16614 16215 -16580
rect 16249 -16614 16287 -16580
rect 16321 -16614 16359 -16580
rect 16393 -16614 16431 -16580
rect 16465 -16614 16503 -16580
rect 16537 -16614 16584 -16580
rect 16096 -16620 16584 -16614
rect 15800 -16708 15814 -16683
rect 14830 -16717 14836 -16708
rect 14790 -16755 14836 -16717
rect 14790 -16789 14796 -16755
rect 14830 -16789 14836 -16755
rect 14790 -16827 14836 -16789
rect 14790 -16861 14796 -16827
rect 14830 -16861 14836 -16827
rect 14790 -16899 14836 -16861
rect 14790 -16933 14796 -16899
rect 14830 -16933 14836 -16899
rect 14790 -16971 14836 -16933
rect 14790 -17005 14796 -16971
rect 14830 -17005 14836 -16971
rect 14790 -17043 14836 -17005
rect 14790 -17077 14796 -17043
rect 14830 -17077 14836 -17043
rect 14790 -17115 14836 -17077
rect 14790 -17149 14796 -17115
rect 14830 -17149 14836 -17115
rect 14790 -17187 14836 -17149
rect 13812 -17221 13826 -17194
rect 7952 -17290 8440 -17284
rect 7952 -17324 7999 -17290
rect 8033 -17324 8071 -17290
rect 8105 -17324 8143 -17290
rect 8177 -17324 8215 -17290
rect 8249 -17324 8287 -17290
rect 8321 -17324 8359 -17290
rect 8393 -17324 8440 -17290
rect 7952 -17330 8440 -17324
rect 8970 -17290 9458 -17284
rect 8970 -17324 9017 -17290
rect 9051 -17324 9089 -17290
rect 9123 -17324 9161 -17290
rect 9195 -17324 9233 -17290
rect 9267 -17324 9305 -17290
rect 9339 -17324 9377 -17290
rect 9411 -17324 9458 -17290
rect 8970 -17330 9458 -17324
rect 9988 -17290 10476 -17284
rect 9988 -17324 10035 -17290
rect 10069 -17324 10107 -17290
rect 10141 -17324 10179 -17290
rect 10213 -17324 10251 -17290
rect 10285 -17324 10323 -17290
rect 10357 -17324 10395 -17290
rect 10429 -17324 10476 -17290
rect 9988 -17330 10476 -17324
rect 11006 -17290 11494 -17284
rect 11006 -17324 11053 -17290
rect 11087 -17324 11125 -17290
rect 11159 -17324 11197 -17290
rect 11231 -17324 11269 -17290
rect 11303 -17324 11341 -17290
rect 11375 -17324 11413 -17290
rect 11447 -17324 11494 -17290
rect 11006 -17330 11494 -17324
rect 12024 -17290 12512 -17284
rect 12024 -17324 12071 -17290
rect 12105 -17324 12143 -17290
rect 12177 -17324 12215 -17290
rect 12249 -17324 12287 -17290
rect 12321 -17324 12359 -17290
rect 12393 -17324 12431 -17290
rect 12465 -17324 12512 -17290
rect 12024 -17330 12238 -17324
rect 12240 -17330 12512 -17324
rect 13042 -17290 13530 -17284
rect 13042 -17324 13089 -17290
rect 13123 -17324 13161 -17290
rect 13195 -17324 13233 -17290
rect 13267 -17324 13305 -17290
rect 13339 -17324 13377 -17290
rect 13411 -17324 13449 -17290
rect 13483 -17324 13530 -17290
rect 13042 -17330 13264 -17324
rect 13268 -17330 13530 -17324
rect 7652 -17394 7724 -17390
rect 7652 -17446 7662 -17394
rect 7714 -17446 7724 -17394
rect 7652 -17450 7724 -17446
rect 5614 -17654 5686 -17650
rect 6122 -17604 6194 -17600
rect 4598 -17698 4670 -17694
rect 4598 -17750 4608 -17698
rect 4660 -17750 4670 -17698
rect 4598 -17754 4670 -17750
rect 3880 -17812 4368 -17806
rect 3880 -17846 3927 -17812
rect 3961 -17846 3999 -17812
rect 4033 -17846 4071 -17812
rect 4105 -17846 4143 -17812
rect 4177 -17846 4215 -17812
rect 4249 -17846 4287 -17812
rect 4321 -17846 4368 -17812
rect 3880 -17852 4368 -17846
rect 3584 -17934 3598 -17915
rect 2574 -17987 2620 -17949
rect 2574 -18021 2580 -17987
rect 2614 -18021 2620 -17987
rect 2574 -18059 2620 -18021
rect 2574 -18093 2580 -18059
rect 2614 -18093 2620 -18059
rect 2574 -18131 2620 -18093
rect 2574 -18165 2580 -18131
rect 2614 -18165 2620 -18131
rect 2574 -18203 2620 -18165
rect 2574 -18237 2580 -18203
rect 2614 -18237 2620 -18203
rect 2574 -18275 2620 -18237
rect 2574 -18309 2580 -18275
rect 2614 -18309 2620 -18275
rect 2574 -18347 2620 -18309
rect 2574 -18381 2580 -18347
rect 2614 -18381 2620 -18347
rect 2574 -18419 2620 -18381
rect 2574 -18426 2580 -18419
rect 2564 -18453 2580 -18426
rect 2614 -18426 2620 -18419
rect 3592 -17949 3598 -17934
rect 3632 -17934 3644 -17915
rect 4604 -17915 4664 -17754
rect 4898 -17812 5386 -17806
rect 4898 -17846 4945 -17812
rect 4979 -17846 5017 -17812
rect 5051 -17846 5089 -17812
rect 5123 -17846 5161 -17812
rect 5195 -17846 5233 -17812
rect 5267 -17846 5305 -17812
rect 5339 -17846 5386 -17812
rect 4898 -17852 5386 -17846
rect 3632 -17949 3638 -17934
rect 4604 -17936 4616 -17915
rect 3592 -17987 3638 -17949
rect 3592 -18021 3598 -17987
rect 3632 -18021 3638 -17987
rect 3592 -18059 3638 -18021
rect 3592 -18093 3598 -18059
rect 3632 -18093 3638 -18059
rect 3592 -18131 3638 -18093
rect 3592 -18165 3598 -18131
rect 3632 -18165 3638 -18131
rect 3592 -18203 3638 -18165
rect 3592 -18237 3598 -18203
rect 3632 -18237 3638 -18203
rect 3592 -18275 3638 -18237
rect 3592 -18309 3598 -18275
rect 3632 -18309 3638 -18275
rect 3592 -18347 3638 -18309
rect 3592 -18381 3598 -18347
rect 3632 -18381 3638 -18347
rect 3592 -18419 3638 -18381
rect 2614 -18453 2624 -18426
rect 3592 -18430 3598 -18419
rect 2564 -18634 2624 -18453
rect 3582 -18453 3598 -18430
rect 3632 -18430 3638 -18419
rect 4610 -17949 4616 -17936
rect 4650 -17936 4664 -17915
rect 5620 -17915 5680 -17654
rect 6122 -17656 6132 -17604
rect 6184 -17656 6194 -17604
rect 6122 -17660 6194 -17656
rect 7144 -17604 7216 -17600
rect 7144 -17656 7154 -17604
rect 7206 -17656 7216 -17604
rect 7144 -17660 7216 -17656
rect 6632 -17698 6704 -17694
rect 6632 -17750 6642 -17698
rect 6694 -17750 6704 -17698
rect 6632 -17754 6704 -17750
rect 5916 -17812 6404 -17806
rect 5916 -17846 5963 -17812
rect 5997 -17846 6035 -17812
rect 6069 -17846 6107 -17812
rect 6141 -17846 6179 -17812
rect 6213 -17846 6251 -17812
rect 6285 -17846 6323 -17812
rect 6357 -17846 6404 -17812
rect 5916 -17852 6404 -17846
rect 4650 -17949 4656 -17936
rect 5620 -17948 5634 -17915
rect 4610 -17987 4656 -17949
rect 4610 -18021 4616 -17987
rect 4650 -18021 4656 -17987
rect 4610 -18059 4656 -18021
rect 4610 -18093 4616 -18059
rect 4650 -18093 4656 -18059
rect 4610 -18131 4656 -18093
rect 4610 -18165 4616 -18131
rect 4650 -18165 4656 -18131
rect 4610 -18203 4656 -18165
rect 4610 -18237 4616 -18203
rect 4650 -18237 4656 -18203
rect 4610 -18275 4656 -18237
rect 4610 -18309 4616 -18275
rect 4650 -18309 4656 -18275
rect 4610 -18347 4656 -18309
rect 4610 -18381 4616 -18347
rect 4650 -18381 4656 -18347
rect 4610 -18419 4656 -18381
rect 3632 -18453 3642 -18430
rect 2862 -18522 3350 -18516
rect 2862 -18556 2909 -18522
rect 2943 -18556 2981 -18522
rect 3015 -18556 3053 -18522
rect 3087 -18556 3125 -18522
rect 3159 -18556 3197 -18522
rect 3231 -18556 3269 -18522
rect 3303 -18556 3350 -18522
rect 2862 -18562 3350 -18556
rect 3076 -18634 3136 -18562
rect 3582 -18634 3642 -18453
rect 4610 -18453 4616 -18419
rect 4650 -18453 4656 -18419
rect 4610 -18484 4656 -18453
rect 5628 -17949 5634 -17948
rect 5668 -17948 5680 -17915
rect 6638 -17915 6698 -17754
rect 7150 -17806 7210 -17660
rect 6934 -17812 7422 -17806
rect 6934 -17846 6981 -17812
rect 7015 -17846 7053 -17812
rect 7087 -17846 7125 -17812
rect 7159 -17846 7197 -17812
rect 7231 -17846 7269 -17812
rect 7303 -17846 7341 -17812
rect 7375 -17846 7422 -17812
rect 6934 -17852 7422 -17846
rect 6638 -17940 6652 -17915
rect 5668 -17949 5674 -17948
rect 5628 -17987 5674 -17949
rect 5628 -18021 5634 -17987
rect 5668 -18021 5674 -17987
rect 5628 -18059 5674 -18021
rect 5628 -18093 5634 -18059
rect 5668 -18093 5674 -18059
rect 5628 -18131 5674 -18093
rect 5628 -18165 5634 -18131
rect 5668 -18165 5674 -18131
rect 5628 -18203 5674 -18165
rect 5628 -18237 5634 -18203
rect 5668 -18237 5674 -18203
rect 5628 -18275 5674 -18237
rect 5628 -18309 5634 -18275
rect 5668 -18309 5674 -18275
rect 5628 -18347 5674 -18309
rect 5628 -18381 5634 -18347
rect 5668 -18381 5674 -18347
rect 5628 -18419 5674 -18381
rect 5628 -18453 5634 -18419
rect 5668 -18453 5674 -18419
rect 6646 -17949 6652 -17940
rect 6686 -17940 6698 -17915
rect 7658 -17915 7718 -17450
rect 8164 -17600 8224 -17330
rect 9182 -17492 9242 -17330
rect 10202 -17380 10262 -17330
rect 11202 -17380 11262 -17330
rect 12240 -17380 12300 -17330
rect 13268 -17380 13328 -17330
rect 9684 -17394 9756 -17390
rect 9684 -17446 9694 -17394
rect 9746 -17446 9756 -17394
rect 10202 -17440 13328 -17380
rect 9684 -17450 9756 -17446
rect 9176 -17496 9248 -17492
rect 9176 -17548 9186 -17496
rect 9238 -17548 9248 -17496
rect 9176 -17552 9248 -17548
rect 8158 -17604 8230 -17600
rect 8158 -17656 8168 -17604
rect 8220 -17656 8230 -17604
rect 8158 -17660 8230 -17656
rect 9176 -17604 9248 -17600
rect 9176 -17656 9186 -17604
rect 9238 -17656 9248 -17604
rect 9176 -17660 9248 -17656
rect 8164 -17806 8224 -17660
rect 8668 -17698 8740 -17694
rect 8668 -17750 8678 -17698
rect 8730 -17750 8740 -17698
rect 8668 -17754 8740 -17750
rect 7952 -17812 8440 -17806
rect 7952 -17846 7999 -17812
rect 8033 -17846 8071 -17812
rect 8105 -17846 8143 -17812
rect 8177 -17846 8215 -17812
rect 8249 -17846 8287 -17812
rect 8321 -17846 8359 -17812
rect 8393 -17846 8440 -17812
rect 7952 -17852 8440 -17846
rect 6686 -17949 6692 -17940
rect 6646 -17987 6692 -17949
rect 6646 -18021 6652 -17987
rect 6686 -18021 6692 -17987
rect 6646 -18059 6692 -18021
rect 6646 -18093 6652 -18059
rect 6686 -18093 6692 -18059
rect 6646 -18131 6692 -18093
rect 6646 -18165 6652 -18131
rect 6686 -18165 6692 -18131
rect 6646 -18203 6692 -18165
rect 6646 -18237 6652 -18203
rect 6686 -18237 6692 -18203
rect 6646 -18275 6692 -18237
rect 6646 -18309 6652 -18275
rect 6686 -18309 6692 -18275
rect 6646 -18347 6692 -18309
rect 6646 -18381 6652 -18347
rect 6686 -18381 6692 -18347
rect 6646 -18419 6692 -18381
rect 6646 -18436 6652 -18419
rect 5628 -18484 5674 -18453
rect 6638 -18453 6652 -18436
rect 6686 -18436 6692 -18419
rect 7658 -17949 7670 -17915
rect 7704 -17949 7718 -17915
rect 8674 -17915 8734 -17754
rect 9182 -17806 9242 -17660
rect 8970 -17812 9458 -17806
rect 8970 -17846 9017 -17812
rect 9051 -17846 9089 -17812
rect 9123 -17846 9161 -17812
rect 9195 -17846 9233 -17812
rect 9267 -17846 9305 -17812
rect 9339 -17846 9377 -17812
rect 9411 -17846 9458 -17812
rect 8970 -17852 9458 -17846
rect 8674 -17932 8688 -17915
rect 7658 -17987 7718 -17949
rect 7658 -18021 7670 -17987
rect 7704 -18021 7718 -17987
rect 7658 -18059 7718 -18021
rect 7658 -18093 7670 -18059
rect 7704 -18093 7718 -18059
rect 7658 -18131 7718 -18093
rect 7658 -18165 7670 -18131
rect 7704 -18165 7718 -18131
rect 7658 -18203 7718 -18165
rect 7658 -18237 7670 -18203
rect 7704 -18237 7718 -18203
rect 7658 -18275 7718 -18237
rect 7658 -18309 7670 -18275
rect 7704 -18309 7718 -18275
rect 7658 -18347 7718 -18309
rect 7658 -18381 7670 -18347
rect 7704 -18381 7718 -18347
rect 7658 -18419 7718 -18381
rect 6686 -18453 6698 -18436
rect 3880 -18522 4368 -18516
rect 3880 -18556 3927 -18522
rect 3961 -18556 3999 -18522
rect 4033 -18556 4071 -18522
rect 4105 -18556 4143 -18522
rect 4177 -18556 4215 -18522
rect 4249 -18556 4287 -18522
rect 4321 -18556 4368 -18522
rect 3880 -18562 4368 -18556
rect 4898 -18522 5386 -18516
rect 4898 -18556 4945 -18522
rect 4979 -18556 5017 -18522
rect 5051 -18556 5089 -18522
rect 5123 -18556 5161 -18522
rect 5195 -18556 5233 -18522
rect 5267 -18556 5305 -18522
rect 5339 -18556 5386 -18522
rect 4898 -18562 5386 -18556
rect 5916 -18522 6404 -18516
rect 5916 -18556 5963 -18522
rect 5997 -18556 6035 -18522
rect 6069 -18556 6107 -18522
rect 6141 -18556 6179 -18522
rect 6213 -18556 6251 -18522
rect 6285 -18556 6323 -18522
rect 6357 -18556 6404 -18522
rect 5916 -18562 6404 -18556
rect 4086 -18618 4146 -18562
rect 2564 -18694 3642 -18634
rect 4080 -18622 4152 -18618
rect 4080 -18674 4090 -18622
rect 4142 -18674 4152 -18622
rect 4080 -18678 4152 -18674
rect 4990 -18622 5062 -18618
rect 4990 -18674 5000 -18622
rect 5052 -18674 5062 -18622
rect 4990 -18678 5062 -18674
rect 4080 -18838 4152 -18834
rect 4080 -18890 4090 -18838
rect 4142 -18890 4152 -18838
rect 4080 -18894 4152 -18890
rect 4086 -18900 4148 -18894
rect 2448 -18942 2510 -18932
rect 2448 -18994 2454 -18942
rect 2506 -18994 2510 -18942
rect 2448 -19004 2510 -18994
rect 2330 -20200 2402 -20196
rect 2330 -20252 2340 -20200
rect 2392 -20252 2402 -20200
rect 2330 -20256 2402 -20252
rect 2230 -21260 2294 -21254
rect 2230 -21312 2242 -21260
rect 2230 -21318 2294 -21312
rect 2230 -22440 2290 -21318
rect 2336 -22314 2396 -20256
rect 2448 -21182 2508 -19004
rect 4088 -19040 4148 -18900
rect 4996 -19040 5056 -18678
rect 5124 -18838 5184 -18562
rect 5992 -18622 6064 -18618
rect 5992 -18674 6002 -18622
rect 6054 -18674 6064 -18622
rect 5992 -18678 6064 -18674
rect 5124 -18890 5128 -18838
rect 5180 -18890 5184 -18838
rect 5124 -18900 5184 -18890
rect 5998 -19040 6058 -18678
rect 6138 -18834 6198 -18562
rect 6638 -18720 6698 -18453
rect 7658 -18453 7670 -18419
rect 7704 -18453 7718 -18419
rect 6934 -18522 7422 -18516
rect 6934 -18556 6981 -18522
rect 7015 -18556 7053 -18522
rect 7087 -18556 7125 -18522
rect 7159 -18556 7197 -18522
rect 7231 -18556 7269 -18522
rect 7303 -18556 7341 -18522
rect 7375 -18556 7422 -18522
rect 6934 -18562 7126 -18556
rect 7150 -18562 7422 -18556
rect 7150 -18618 7210 -18562
rect 7144 -18622 7216 -18618
rect 7144 -18674 7154 -18622
rect 7206 -18674 7216 -18622
rect 7144 -18678 7216 -18674
rect 6632 -18724 6704 -18720
rect 6632 -18776 6642 -18724
rect 6694 -18776 6704 -18724
rect 6632 -18780 6704 -18776
rect 6132 -18838 6204 -18834
rect 6132 -18890 6142 -18838
rect 6194 -18890 6204 -18838
rect 6132 -18894 6204 -18890
rect 7150 -19040 7210 -18678
rect 2862 -19046 3350 -19040
rect 2862 -19080 2909 -19046
rect 2943 -19080 2981 -19046
rect 3015 -19080 3053 -19046
rect 3087 -19080 3125 -19046
rect 3159 -19080 3197 -19046
rect 3231 -19080 3269 -19046
rect 3303 -19080 3350 -19046
rect 2862 -19086 3350 -19080
rect 3880 -19046 4368 -19040
rect 3880 -19080 3927 -19046
rect 3961 -19080 3999 -19046
rect 4033 -19080 4071 -19046
rect 4105 -19080 4143 -19046
rect 4177 -19080 4215 -19046
rect 4249 -19080 4287 -19046
rect 4321 -19080 4368 -19046
rect 3880 -19086 4368 -19080
rect 4898 -19046 5386 -19040
rect 4898 -19080 4945 -19046
rect 4979 -19080 5017 -19046
rect 5051 -19080 5089 -19046
rect 5123 -19080 5161 -19046
rect 5195 -19080 5233 -19046
rect 5267 -19080 5305 -19046
rect 5339 -19080 5386 -19046
rect 4898 -19086 5386 -19080
rect 5916 -19046 6404 -19040
rect 5916 -19080 5963 -19046
rect 5997 -19080 6035 -19046
rect 6069 -19080 6107 -19046
rect 6141 -19080 6179 -19046
rect 6213 -19080 6251 -19046
rect 6285 -19080 6323 -19046
rect 6357 -19080 6404 -19046
rect 5916 -19086 6404 -19080
rect 6934 -19046 7422 -19040
rect 6934 -19080 6981 -19046
rect 7015 -19080 7053 -19046
rect 7087 -19080 7125 -19046
rect 7159 -19080 7197 -19046
rect 7231 -19080 7269 -19046
rect 7303 -19080 7341 -19046
rect 7375 -19080 7422 -19046
rect 6934 -19086 7422 -19080
rect 2574 -19149 2620 -19118
rect 2574 -19183 2580 -19149
rect 2614 -19183 2620 -19149
rect 2574 -19221 2620 -19183
rect 2574 -19255 2580 -19221
rect 2614 -19255 2620 -19221
rect 2574 -19293 2620 -19255
rect 2574 -19327 2580 -19293
rect 2614 -19327 2620 -19293
rect 2574 -19365 2620 -19327
rect 2574 -19399 2580 -19365
rect 2614 -19399 2620 -19365
rect 2574 -19437 2620 -19399
rect 2574 -19471 2580 -19437
rect 2614 -19471 2620 -19437
rect 2574 -19509 2620 -19471
rect 2574 -19543 2580 -19509
rect 2614 -19543 2620 -19509
rect 2574 -19581 2620 -19543
rect 2574 -19615 2580 -19581
rect 2614 -19615 2620 -19581
rect 2574 -19653 2620 -19615
rect 2574 -19668 2580 -19653
rect 2568 -19687 2580 -19668
rect 2614 -19668 2620 -19653
rect 3592 -19149 3638 -19118
rect 3592 -19183 3598 -19149
rect 3632 -19183 3638 -19149
rect 3592 -19221 3638 -19183
rect 3592 -19255 3598 -19221
rect 3632 -19255 3638 -19221
rect 3592 -19293 3638 -19255
rect 3592 -19327 3598 -19293
rect 3632 -19327 3638 -19293
rect 3592 -19365 3638 -19327
rect 3592 -19399 3598 -19365
rect 3632 -19399 3638 -19365
rect 3592 -19437 3638 -19399
rect 3592 -19471 3598 -19437
rect 3632 -19471 3638 -19437
rect 3592 -19509 3638 -19471
rect 3592 -19543 3598 -19509
rect 3632 -19543 3638 -19509
rect 3592 -19581 3638 -19543
rect 3592 -19615 3598 -19581
rect 3632 -19615 3638 -19581
rect 3592 -19653 3638 -19615
rect 3592 -19668 3598 -19653
rect 2614 -19687 2628 -19668
rect 2568 -19836 2628 -19687
rect 3586 -19687 3598 -19668
rect 3632 -19668 3638 -19653
rect 4610 -19149 4656 -19118
rect 4610 -19183 4616 -19149
rect 4650 -19183 4656 -19149
rect 4610 -19221 4656 -19183
rect 4610 -19255 4616 -19221
rect 4650 -19255 4656 -19221
rect 4610 -19293 4656 -19255
rect 4610 -19327 4616 -19293
rect 4650 -19327 4656 -19293
rect 4610 -19365 4656 -19327
rect 4610 -19399 4616 -19365
rect 4650 -19399 4656 -19365
rect 4610 -19437 4656 -19399
rect 4610 -19471 4616 -19437
rect 4650 -19471 4656 -19437
rect 4610 -19509 4656 -19471
rect 4610 -19543 4616 -19509
rect 4650 -19543 4656 -19509
rect 4610 -19581 4656 -19543
rect 4610 -19615 4616 -19581
rect 4650 -19615 4656 -19581
rect 4610 -19653 4656 -19615
rect 5628 -19149 5674 -19118
rect 5628 -19183 5634 -19149
rect 5668 -19183 5674 -19149
rect 5628 -19221 5674 -19183
rect 5628 -19255 5634 -19221
rect 5668 -19255 5674 -19221
rect 5628 -19293 5674 -19255
rect 5628 -19327 5634 -19293
rect 5668 -19327 5674 -19293
rect 5628 -19365 5674 -19327
rect 5628 -19399 5634 -19365
rect 5668 -19399 5674 -19365
rect 5628 -19437 5674 -19399
rect 5628 -19471 5634 -19437
rect 5668 -19471 5674 -19437
rect 5628 -19509 5674 -19471
rect 5628 -19543 5634 -19509
rect 5668 -19543 5674 -19509
rect 5628 -19581 5674 -19543
rect 5628 -19615 5634 -19581
rect 5668 -19615 5674 -19581
rect 5628 -19648 5674 -19615
rect 6646 -19149 6692 -19118
rect 6646 -19183 6652 -19149
rect 6686 -19183 6692 -19149
rect 6646 -19221 6692 -19183
rect 7658 -19149 7718 -18453
rect 8682 -17949 8688 -17932
rect 8722 -17932 8734 -17915
rect 9690 -17915 9750 -17450
rect 10196 -17604 10268 -17600
rect 10196 -17656 10206 -17604
rect 10258 -17656 10268 -17604
rect 10196 -17660 10268 -17656
rect 13268 -17616 13328 -17440
rect 13766 -17506 13826 -17221
rect 14790 -17221 14796 -17187
rect 14830 -17221 14836 -17187
rect 14790 -17252 14836 -17221
rect 15808 -16717 15814 -16708
rect 15848 -16708 15860 -16683
rect 16818 -16683 16878 -16524
rect 17326 -16574 17386 -16096
rect 17836 -16134 17896 -15987
rect 18854 -15987 18868 -15953
rect 18902 -15987 18914 -15953
rect 19880 -15953 19926 -15915
rect 19880 -15962 19886 -15953
rect 18132 -16056 18620 -16050
rect 18132 -16090 18179 -16056
rect 18213 -16090 18251 -16056
rect 18285 -16090 18323 -16056
rect 18357 -16090 18395 -16056
rect 18429 -16090 18467 -16056
rect 18501 -16090 18539 -16056
rect 18573 -16090 18620 -16056
rect 18132 -16096 18620 -16090
rect 17830 -16138 17902 -16134
rect 17830 -16190 17840 -16138
rect 17892 -16190 17902 -16138
rect 17830 -16194 17902 -16190
rect 17114 -16580 17602 -16574
rect 17114 -16614 17161 -16580
rect 17195 -16614 17233 -16580
rect 17267 -16614 17305 -16580
rect 17339 -16614 17377 -16580
rect 17411 -16614 17449 -16580
rect 17483 -16614 17521 -16580
rect 17555 -16614 17602 -16580
rect 17114 -16620 17602 -16614
rect 16818 -16694 16832 -16683
rect 15848 -16717 15854 -16708
rect 15808 -16755 15854 -16717
rect 15808 -16789 15814 -16755
rect 15848 -16789 15854 -16755
rect 15808 -16827 15854 -16789
rect 15808 -16861 15814 -16827
rect 15848 -16861 15854 -16827
rect 15808 -16899 15854 -16861
rect 15808 -16933 15814 -16899
rect 15848 -16933 15854 -16899
rect 15808 -16971 15854 -16933
rect 15808 -17005 15814 -16971
rect 15848 -17005 15854 -16971
rect 15808 -17043 15854 -17005
rect 15808 -17077 15814 -17043
rect 15848 -17077 15854 -17043
rect 15808 -17115 15854 -17077
rect 15808 -17149 15814 -17115
rect 15848 -17149 15854 -17115
rect 15808 -17187 15854 -17149
rect 15808 -17221 15814 -17187
rect 15848 -17221 15854 -17187
rect 16826 -16717 16832 -16694
rect 16866 -16694 16878 -16683
rect 17836 -16683 17896 -16194
rect 18352 -16574 18412 -16096
rect 18854 -16350 18914 -15987
rect 19870 -15987 19886 -15962
rect 19920 -15962 19926 -15953
rect 20898 -15449 20944 -15418
rect 20898 -15483 20904 -15449
rect 20938 -15483 20944 -15449
rect 20898 -15521 20944 -15483
rect 20898 -15555 20904 -15521
rect 20938 -15555 20944 -15521
rect 20898 -15593 20944 -15555
rect 20898 -15627 20904 -15593
rect 20938 -15627 20944 -15593
rect 20898 -15665 20944 -15627
rect 20898 -15699 20904 -15665
rect 20938 -15699 20944 -15665
rect 20898 -15737 20944 -15699
rect 20898 -15771 20904 -15737
rect 20938 -15771 20944 -15737
rect 20898 -15809 20944 -15771
rect 20898 -15843 20904 -15809
rect 20938 -15843 20944 -15809
rect 20898 -15881 20944 -15843
rect 20898 -15915 20904 -15881
rect 20938 -15915 20944 -15881
rect 20898 -15953 20944 -15915
rect 20898 -15962 20904 -15953
rect 19920 -15987 19930 -15962
rect 19150 -16056 19638 -16050
rect 19150 -16090 19197 -16056
rect 19231 -16090 19269 -16056
rect 19303 -16090 19341 -16056
rect 19375 -16090 19413 -16056
rect 19447 -16090 19485 -16056
rect 19519 -16090 19557 -16056
rect 19591 -16090 19638 -16056
rect 19150 -16096 19638 -16090
rect 18848 -16354 18920 -16350
rect 18848 -16406 18858 -16354
rect 18910 -16406 18920 -16354
rect 18848 -16410 18920 -16406
rect 19360 -16400 19420 -16096
rect 19870 -16242 19930 -15987
rect 20894 -15987 20904 -15962
rect 20938 -15962 20944 -15953
rect 21916 -15449 21962 -15418
rect 21916 -15483 21922 -15449
rect 21956 -15483 21962 -15449
rect 22926 -15449 22986 -15264
rect 23028 -15232 23100 -15228
rect 23028 -15284 23038 -15232
rect 23090 -15284 23100 -15232
rect 23028 -15288 23100 -15284
rect 22926 -15458 22940 -15449
rect 21916 -15521 21962 -15483
rect 21916 -15555 21922 -15521
rect 21956 -15555 21962 -15521
rect 21916 -15593 21962 -15555
rect 21916 -15627 21922 -15593
rect 21956 -15627 21962 -15593
rect 21916 -15665 21962 -15627
rect 21916 -15699 21922 -15665
rect 21956 -15699 21962 -15665
rect 21916 -15737 21962 -15699
rect 21916 -15771 21922 -15737
rect 21956 -15771 21962 -15737
rect 21916 -15809 21962 -15771
rect 21916 -15843 21922 -15809
rect 21956 -15843 21962 -15809
rect 21916 -15881 21962 -15843
rect 21916 -15915 21922 -15881
rect 21956 -15915 21962 -15881
rect 21916 -15953 21962 -15915
rect 22934 -15483 22940 -15458
rect 22974 -15458 22986 -15449
rect 22974 -15483 22980 -15458
rect 22934 -15521 22980 -15483
rect 22934 -15555 22940 -15521
rect 22974 -15555 22980 -15521
rect 22934 -15593 22980 -15555
rect 22934 -15627 22940 -15593
rect 22974 -15627 22980 -15593
rect 22934 -15665 22980 -15627
rect 22934 -15699 22940 -15665
rect 22974 -15699 22980 -15665
rect 22934 -15737 22980 -15699
rect 22934 -15771 22940 -15737
rect 22974 -15771 22980 -15737
rect 22934 -15809 22980 -15771
rect 22934 -15843 22940 -15809
rect 22974 -15843 22980 -15809
rect 22934 -15881 22980 -15843
rect 22934 -15915 22940 -15881
rect 22974 -15915 22980 -15881
rect 22934 -15948 22980 -15915
rect 21916 -15956 21922 -15953
rect 20938 -15987 20954 -15962
rect 20168 -16056 20656 -16050
rect 20168 -16090 20215 -16056
rect 20249 -16090 20287 -16056
rect 20321 -16090 20359 -16056
rect 20393 -16090 20431 -16056
rect 20465 -16090 20503 -16056
rect 20537 -16090 20575 -16056
rect 20609 -16090 20656 -16056
rect 20168 -16096 20656 -16090
rect 20376 -16240 20436 -16096
rect 19864 -16246 19936 -16242
rect 19864 -16298 19874 -16246
rect 19926 -16298 19936 -16246
rect 19864 -16302 19936 -16298
rect 20374 -16250 20436 -16240
rect 20374 -16302 20378 -16250
rect 20430 -16302 20436 -16250
rect 20374 -16312 20436 -16302
rect 20376 -16400 20436 -16312
rect 20894 -16350 20954 -15987
rect 21910 -15987 21922 -15956
rect 21956 -15956 21962 -15953
rect 22928 -15953 22988 -15948
rect 21956 -15987 21970 -15956
rect 21186 -16056 21674 -16050
rect 21186 -16090 21233 -16056
rect 21267 -16090 21305 -16056
rect 21339 -16090 21377 -16056
rect 21411 -16090 21449 -16056
rect 21483 -16090 21521 -16056
rect 21555 -16090 21593 -16056
rect 21627 -16090 21674 -16056
rect 21186 -16096 21674 -16090
rect 19360 -16460 20436 -16400
rect 20888 -16354 20960 -16350
rect 20888 -16406 20898 -16354
rect 20950 -16406 20960 -16354
rect 20888 -16410 20960 -16406
rect 18848 -16468 18920 -16464
rect 18848 -16520 18858 -16468
rect 18910 -16520 18920 -16468
rect 18848 -16524 18920 -16520
rect 18132 -16580 18620 -16574
rect 18132 -16614 18179 -16580
rect 18213 -16614 18251 -16580
rect 18285 -16614 18323 -16580
rect 18357 -16614 18395 -16580
rect 18429 -16614 18467 -16580
rect 18501 -16614 18539 -16580
rect 18573 -16614 18620 -16580
rect 18132 -16620 18620 -16614
rect 16866 -16717 16872 -16694
rect 17836 -16704 17850 -16683
rect 16826 -16755 16872 -16717
rect 16826 -16789 16832 -16755
rect 16866 -16789 16872 -16755
rect 16826 -16827 16872 -16789
rect 16826 -16861 16832 -16827
rect 16866 -16861 16872 -16827
rect 16826 -16899 16872 -16861
rect 16826 -16933 16832 -16899
rect 16866 -16933 16872 -16899
rect 16826 -16971 16872 -16933
rect 16826 -17005 16832 -16971
rect 16866 -17005 16872 -16971
rect 16826 -17043 16872 -17005
rect 16826 -17077 16832 -17043
rect 16866 -17077 16872 -17043
rect 16826 -17115 16872 -17077
rect 16826 -17149 16832 -17115
rect 16866 -17149 16872 -17115
rect 16826 -17187 16872 -17149
rect 16826 -17200 16832 -17187
rect 15808 -17252 15854 -17221
rect 16818 -17221 16832 -17200
rect 16866 -17200 16872 -17187
rect 17844 -16717 17850 -16704
rect 17884 -16704 17896 -16683
rect 18854 -16683 18914 -16524
rect 19360 -16574 19420 -16460
rect 20376 -16574 20436 -16460
rect 20886 -16468 20958 -16464
rect 20886 -16520 20896 -16468
rect 20948 -16520 20958 -16468
rect 20886 -16524 20958 -16520
rect 19150 -16580 19638 -16574
rect 19150 -16614 19197 -16580
rect 19231 -16614 19269 -16580
rect 19303 -16614 19341 -16580
rect 19375 -16614 19413 -16580
rect 19447 -16614 19485 -16580
rect 19519 -16614 19557 -16580
rect 19591 -16614 19638 -16580
rect 19150 -16620 19638 -16614
rect 20168 -16580 20656 -16574
rect 20168 -16614 20215 -16580
rect 20249 -16614 20287 -16580
rect 20321 -16614 20359 -16580
rect 20393 -16614 20431 -16580
rect 20465 -16614 20503 -16580
rect 20537 -16614 20575 -16580
rect 20609 -16614 20656 -16580
rect 20168 -16620 20656 -16614
rect 17884 -16717 17890 -16704
rect 18854 -16706 18868 -16683
rect 17844 -16755 17890 -16717
rect 17844 -16789 17850 -16755
rect 17884 -16789 17890 -16755
rect 17844 -16827 17890 -16789
rect 17844 -16861 17850 -16827
rect 17884 -16861 17890 -16827
rect 17844 -16899 17890 -16861
rect 17844 -16933 17850 -16899
rect 17884 -16933 17890 -16899
rect 17844 -16971 17890 -16933
rect 17844 -17005 17850 -16971
rect 17884 -17005 17890 -16971
rect 17844 -17043 17890 -17005
rect 17844 -17077 17850 -17043
rect 17884 -17077 17890 -17043
rect 17844 -17115 17890 -17077
rect 17844 -17149 17850 -17115
rect 17884 -17149 17890 -17115
rect 17844 -17187 17890 -17149
rect 16866 -17221 16878 -17200
rect 17844 -17206 17850 -17187
rect 14060 -17290 14548 -17284
rect 14060 -17324 14107 -17290
rect 14141 -17324 14179 -17290
rect 14213 -17324 14251 -17290
rect 14285 -17324 14323 -17290
rect 14357 -17324 14395 -17290
rect 14429 -17324 14467 -17290
rect 14501 -17324 14548 -17290
rect 14060 -17330 14548 -17324
rect 15078 -17290 15566 -17284
rect 15078 -17324 15125 -17290
rect 15159 -17324 15197 -17290
rect 15231 -17324 15269 -17290
rect 15303 -17324 15341 -17290
rect 15375 -17324 15413 -17290
rect 15447 -17324 15485 -17290
rect 15519 -17324 15566 -17290
rect 15078 -17330 15566 -17324
rect 16096 -17290 16584 -17284
rect 16096 -17324 16143 -17290
rect 16177 -17324 16215 -17290
rect 16249 -17324 16287 -17290
rect 16321 -17324 16359 -17290
rect 16393 -17324 16431 -17290
rect 16465 -17324 16503 -17290
rect 16537 -17324 16584 -17290
rect 16096 -17330 16584 -17324
rect 14272 -17382 14332 -17330
rect 14272 -17434 14276 -17382
rect 14328 -17434 14332 -17382
rect 13760 -17510 13832 -17506
rect 13760 -17562 13770 -17510
rect 13822 -17562 13832 -17510
rect 13760 -17566 13832 -17562
rect 14272 -17616 14332 -17434
rect 10202 -17806 10262 -17660
rect 13268 -17676 14332 -17616
rect 15796 -17708 15868 -17704
rect 15796 -17760 15806 -17708
rect 15858 -17760 15868 -17708
rect 15796 -17764 15868 -17760
rect 9988 -17812 10476 -17806
rect 9988 -17846 10035 -17812
rect 10069 -17846 10107 -17812
rect 10141 -17846 10179 -17812
rect 10213 -17846 10251 -17812
rect 10285 -17846 10323 -17812
rect 10357 -17846 10395 -17812
rect 10429 -17846 10476 -17812
rect 9988 -17852 10476 -17846
rect 11006 -17812 11494 -17806
rect 11006 -17846 11053 -17812
rect 11087 -17846 11125 -17812
rect 11159 -17846 11197 -17812
rect 11231 -17846 11269 -17812
rect 11303 -17846 11341 -17812
rect 11375 -17846 11413 -17812
rect 11447 -17846 11494 -17812
rect 11006 -17852 11494 -17846
rect 12024 -17812 12512 -17806
rect 12024 -17846 12071 -17812
rect 12105 -17846 12143 -17812
rect 12177 -17846 12215 -17812
rect 12249 -17846 12287 -17812
rect 12321 -17846 12359 -17812
rect 12393 -17846 12431 -17812
rect 12465 -17846 12512 -17812
rect 12024 -17852 12512 -17846
rect 13042 -17812 13530 -17806
rect 13042 -17846 13089 -17812
rect 13123 -17846 13161 -17812
rect 13195 -17846 13233 -17812
rect 13267 -17846 13305 -17812
rect 13339 -17846 13377 -17812
rect 13411 -17846 13449 -17812
rect 13483 -17846 13530 -17812
rect 13042 -17852 13530 -17846
rect 14060 -17812 14548 -17806
rect 14060 -17846 14107 -17812
rect 14141 -17846 14179 -17812
rect 14213 -17846 14251 -17812
rect 14285 -17846 14323 -17812
rect 14357 -17846 14395 -17812
rect 14429 -17846 14467 -17812
rect 14501 -17846 14548 -17812
rect 14060 -17852 14548 -17846
rect 15078 -17812 15566 -17806
rect 15078 -17846 15125 -17812
rect 15159 -17846 15197 -17812
rect 15231 -17846 15269 -17812
rect 15303 -17846 15341 -17812
rect 15375 -17846 15413 -17812
rect 15447 -17846 15485 -17812
rect 15519 -17846 15566 -17812
rect 15078 -17852 15566 -17846
rect 8722 -17949 8728 -17932
rect 9690 -17934 9706 -17915
rect 8682 -17987 8728 -17949
rect 8682 -18021 8688 -17987
rect 8722 -18021 8728 -17987
rect 8682 -18059 8728 -18021
rect 8682 -18093 8688 -18059
rect 8722 -18093 8728 -18059
rect 8682 -18131 8728 -18093
rect 8682 -18165 8688 -18131
rect 8722 -18165 8728 -18131
rect 8682 -18203 8728 -18165
rect 8682 -18237 8688 -18203
rect 8722 -18237 8728 -18203
rect 8682 -18275 8728 -18237
rect 8682 -18309 8688 -18275
rect 8722 -18309 8728 -18275
rect 8682 -18347 8728 -18309
rect 8682 -18381 8688 -18347
rect 8722 -18381 8728 -18347
rect 8682 -18419 8728 -18381
rect 8682 -18453 8688 -18419
rect 8722 -18453 8728 -18419
rect 8682 -18484 8728 -18453
rect 9700 -17949 9706 -17934
rect 9740 -17934 9750 -17915
rect 10718 -17915 10764 -17884
rect 9740 -17949 9746 -17934
rect 9700 -17987 9746 -17949
rect 9700 -18021 9706 -17987
rect 9740 -18021 9746 -17987
rect 9700 -18059 9746 -18021
rect 9700 -18093 9706 -18059
rect 9740 -18093 9746 -18059
rect 9700 -18131 9746 -18093
rect 9700 -18165 9706 -18131
rect 9740 -18165 9746 -18131
rect 9700 -18203 9746 -18165
rect 9700 -18237 9706 -18203
rect 9740 -18237 9746 -18203
rect 9700 -18275 9746 -18237
rect 9700 -18309 9706 -18275
rect 9740 -18309 9746 -18275
rect 9700 -18347 9746 -18309
rect 9700 -18381 9706 -18347
rect 9740 -18381 9746 -18347
rect 9700 -18419 9746 -18381
rect 9700 -18453 9706 -18419
rect 9740 -18453 9746 -18419
rect 10718 -17949 10724 -17915
rect 10758 -17949 10764 -17915
rect 10718 -17987 10764 -17949
rect 10718 -18021 10724 -17987
rect 10758 -18021 10764 -17987
rect 10718 -18059 10764 -18021
rect 10718 -18093 10724 -18059
rect 10758 -18093 10764 -18059
rect 10718 -18131 10764 -18093
rect 10718 -18165 10724 -18131
rect 10758 -18165 10764 -18131
rect 10718 -18203 10764 -18165
rect 10718 -18237 10724 -18203
rect 10758 -18237 10764 -18203
rect 10718 -18275 10764 -18237
rect 10718 -18309 10724 -18275
rect 10758 -18309 10764 -18275
rect 10718 -18347 10764 -18309
rect 10718 -18381 10724 -18347
rect 10758 -18381 10764 -18347
rect 10718 -18419 10764 -18381
rect 10718 -18430 10724 -18419
rect 9700 -18484 9746 -18453
rect 10710 -18453 10724 -18430
rect 10758 -18430 10764 -18419
rect 11736 -17915 11782 -17884
rect 11736 -17949 11742 -17915
rect 11776 -17949 11782 -17915
rect 11736 -17987 11782 -17949
rect 11736 -18021 11742 -17987
rect 11776 -18021 11782 -17987
rect 11736 -18059 11782 -18021
rect 11736 -18093 11742 -18059
rect 11776 -18093 11782 -18059
rect 11736 -18131 11782 -18093
rect 11736 -18165 11742 -18131
rect 11776 -18165 11782 -18131
rect 11736 -18203 11782 -18165
rect 11736 -18237 11742 -18203
rect 11776 -18237 11782 -18203
rect 11736 -18275 11782 -18237
rect 11736 -18309 11742 -18275
rect 11776 -18309 11782 -18275
rect 11736 -18347 11782 -18309
rect 11736 -18381 11742 -18347
rect 11776 -18381 11782 -18347
rect 11736 -18419 11782 -18381
rect 10758 -18453 10770 -18430
rect 11736 -18434 11742 -18419
rect 7952 -18522 8440 -18516
rect 7952 -18556 7999 -18522
rect 8033 -18556 8071 -18522
rect 8105 -18556 8143 -18522
rect 8177 -18556 8215 -18522
rect 8249 -18556 8287 -18522
rect 8321 -18556 8359 -18522
rect 8393 -18556 8440 -18522
rect 7952 -18562 8220 -18556
rect 8224 -18562 8440 -18556
rect 8970 -18522 9458 -18516
rect 8970 -18556 9017 -18522
rect 9051 -18556 9089 -18522
rect 9123 -18556 9161 -18522
rect 9195 -18556 9233 -18522
rect 9267 -18556 9305 -18522
rect 9339 -18556 9377 -18522
rect 9411 -18556 9458 -18522
rect 8970 -18562 9458 -18556
rect 9988 -18522 10476 -18516
rect 9988 -18556 10035 -18522
rect 10069 -18556 10107 -18522
rect 10141 -18556 10179 -18522
rect 10213 -18556 10251 -18522
rect 10285 -18556 10323 -18522
rect 10357 -18556 10395 -18522
rect 10429 -18556 10476 -18522
rect 9988 -18562 10476 -18556
rect 8160 -18618 8220 -18562
rect 9166 -18618 9226 -18562
rect 10210 -18618 10270 -18562
rect 10710 -18612 10770 -18453
rect 11730 -18453 11742 -18434
rect 11776 -18434 11782 -18419
rect 12754 -17915 12800 -17884
rect 12754 -17949 12760 -17915
rect 12794 -17949 12800 -17915
rect 12754 -17987 12800 -17949
rect 12754 -18021 12760 -17987
rect 12794 -18021 12800 -17987
rect 12754 -18059 12800 -18021
rect 12754 -18093 12760 -18059
rect 12794 -18093 12800 -18059
rect 12754 -18131 12800 -18093
rect 12754 -18165 12760 -18131
rect 12794 -18165 12800 -18131
rect 12754 -18203 12800 -18165
rect 12754 -18237 12760 -18203
rect 12794 -18237 12800 -18203
rect 12754 -18275 12800 -18237
rect 12754 -18309 12760 -18275
rect 12794 -18309 12800 -18275
rect 12754 -18347 12800 -18309
rect 12754 -18381 12760 -18347
rect 12794 -18381 12800 -18347
rect 12754 -18419 12800 -18381
rect 11776 -18453 11790 -18434
rect 12754 -18440 12760 -18419
rect 11006 -18522 11494 -18516
rect 11006 -18556 11053 -18522
rect 11087 -18556 11125 -18522
rect 11159 -18556 11197 -18522
rect 11231 -18556 11269 -18522
rect 11303 -18556 11341 -18522
rect 11375 -18556 11413 -18522
rect 11447 -18556 11494 -18522
rect 11006 -18562 11494 -18556
rect 10704 -18616 10776 -18612
rect 8154 -18622 8226 -18618
rect 8154 -18674 8164 -18622
rect 8216 -18674 8226 -18622
rect 8154 -18678 8226 -18674
rect 9160 -18622 9232 -18618
rect 9160 -18674 9170 -18622
rect 9222 -18674 9232 -18622
rect 9160 -18678 9232 -18674
rect 10204 -18622 10276 -18618
rect 10204 -18674 10214 -18622
rect 10266 -18674 10276 -18622
rect 10704 -18668 10714 -18616
rect 10766 -18668 10776 -18616
rect 10704 -18672 10776 -18668
rect 10204 -18678 10276 -18674
rect 8160 -19040 8220 -18678
rect 9158 -18838 9230 -18834
rect 9158 -18890 9168 -18838
rect 9220 -18890 9230 -18838
rect 9158 -18894 9230 -18890
rect 10198 -18838 10270 -18834
rect 10198 -18890 10208 -18838
rect 10260 -18890 10270 -18838
rect 10198 -18894 10270 -18890
rect 9164 -19040 9224 -18894
rect 9682 -18942 9754 -18938
rect 9682 -18994 9692 -18942
rect 9744 -18994 9754 -18942
rect 9682 -18998 9754 -18994
rect 7952 -19046 8440 -19040
rect 7952 -19080 7999 -19046
rect 8033 -19080 8071 -19046
rect 8105 -19080 8143 -19046
rect 8177 -19080 8215 -19046
rect 8249 -19080 8287 -19046
rect 8321 -19080 8359 -19046
rect 8393 -19080 8440 -19046
rect 7952 -19086 8440 -19080
rect 8970 -19046 9458 -19040
rect 8970 -19080 9017 -19046
rect 9051 -19080 9089 -19046
rect 9123 -19080 9161 -19046
rect 9195 -19080 9233 -19046
rect 9267 -19080 9305 -19046
rect 9339 -19080 9377 -19046
rect 9411 -19080 9458 -19046
rect 8970 -19086 9458 -19080
rect 7658 -19183 7670 -19149
rect 7704 -19183 7718 -19149
rect 7658 -19212 7718 -19183
rect 8682 -19149 8728 -19118
rect 8682 -19183 8688 -19149
rect 8722 -19183 8728 -19149
rect 6646 -19255 6652 -19221
rect 6686 -19255 6692 -19221
rect 6646 -19293 6692 -19255
rect 6646 -19327 6652 -19293
rect 6686 -19327 6692 -19293
rect 6646 -19365 6692 -19327
rect 6646 -19399 6652 -19365
rect 6686 -19399 6692 -19365
rect 6646 -19437 6692 -19399
rect 6646 -19471 6652 -19437
rect 6686 -19471 6692 -19437
rect 6646 -19509 6692 -19471
rect 6646 -19543 6652 -19509
rect 6686 -19543 6692 -19509
rect 6646 -19581 6692 -19543
rect 6646 -19615 6652 -19581
rect 6686 -19615 6692 -19581
rect 4610 -19656 4616 -19653
rect 3632 -19687 3646 -19668
rect 2862 -19756 3350 -19750
rect 2862 -19790 2909 -19756
rect 2943 -19790 2981 -19756
rect 3015 -19790 3053 -19756
rect 3087 -19790 3125 -19756
rect 3159 -19790 3197 -19756
rect 3231 -19790 3269 -19756
rect 3303 -19790 3350 -19756
rect 2862 -19796 3350 -19790
rect 3066 -19836 3126 -19796
rect 3586 -19836 3646 -19687
rect 4602 -19687 4616 -19656
rect 4650 -19656 4656 -19653
rect 5620 -19653 5680 -19648
rect 4650 -19687 4662 -19656
rect 3880 -19756 4368 -19750
rect 3880 -19790 3927 -19756
rect 3961 -19790 3999 -19756
rect 4033 -19790 4071 -19756
rect 4105 -19790 4143 -19756
rect 4177 -19790 4215 -19756
rect 4249 -19790 4287 -19756
rect 4321 -19790 4368 -19756
rect 3880 -19796 4368 -19790
rect 2568 -19896 3646 -19836
rect 3586 -19950 3646 -19896
rect 4078 -19850 4150 -19846
rect 4078 -19902 4088 -19850
rect 4140 -19902 4150 -19850
rect 4078 -19906 4150 -19902
rect 3580 -19954 3652 -19950
rect 3580 -20006 3590 -19954
rect 3642 -20006 3652 -19954
rect 3580 -20010 3652 -20006
rect 3576 -20164 3648 -20160
rect 3576 -20216 3586 -20164
rect 3638 -20216 3648 -20164
rect 3576 -20220 3648 -20216
rect 2862 -20280 3350 -20274
rect 2862 -20314 2909 -20280
rect 2943 -20314 2981 -20280
rect 3015 -20314 3053 -20280
rect 3087 -20314 3125 -20280
rect 3159 -20314 3197 -20280
rect 3231 -20314 3269 -20280
rect 3303 -20314 3350 -20280
rect 2862 -20320 3350 -20314
rect 2574 -20383 2620 -20352
rect 2574 -20417 2580 -20383
rect 2614 -20417 2620 -20383
rect 2574 -20455 2620 -20417
rect 3582 -20383 3642 -20220
rect 4084 -20274 4144 -19906
rect 4602 -20062 4662 -19687
rect 5620 -19687 5634 -19653
rect 5668 -19687 5680 -19653
rect 6646 -19653 6692 -19615
rect 6646 -19660 6652 -19653
rect 4898 -19756 5386 -19750
rect 4898 -19790 4945 -19756
rect 4979 -19790 5017 -19756
rect 5051 -19790 5089 -19756
rect 5123 -19790 5161 -19756
rect 5195 -19790 5233 -19756
rect 5267 -19790 5305 -19756
rect 5339 -19790 5386 -19756
rect 4898 -19796 5386 -19790
rect 5092 -19846 5152 -19796
rect 5086 -19850 5158 -19846
rect 5086 -19902 5096 -19850
rect 5148 -19902 5158 -19850
rect 5086 -19906 5158 -19902
rect 4596 -20066 4668 -20062
rect 4596 -20118 4606 -20066
rect 4658 -20118 4668 -20066
rect 4596 -20122 4668 -20118
rect 5620 -20160 5680 -19687
rect 6640 -19687 6652 -19660
rect 6686 -19660 6692 -19653
rect 7664 -19221 7710 -19212
rect 7664 -19255 7670 -19221
rect 7704 -19255 7710 -19221
rect 7664 -19293 7710 -19255
rect 7664 -19327 7670 -19293
rect 7704 -19327 7710 -19293
rect 7664 -19365 7710 -19327
rect 7664 -19399 7670 -19365
rect 7704 -19399 7710 -19365
rect 7664 -19437 7710 -19399
rect 7664 -19471 7670 -19437
rect 7704 -19471 7710 -19437
rect 7664 -19509 7710 -19471
rect 7664 -19543 7670 -19509
rect 7704 -19543 7710 -19509
rect 7664 -19581 7710 -19543
rect 7664 -19615 7670 -19581
rect 7704 -19615 7710 -19581
rect 7664 -19653 7710 -19615
rect 7664 -19660 7670 -19653
rect 6686 -19687 6700 -19660
rect 5916 -19756 6404 -19750
rect 5916 -19790 5963 -19756
rect 5997 -19790 6035 -19756
rect 6069 -19790 6107 -19756
rect 6141 -19790 6179 -19756
rect 6213 -19790 6251 -19756
rect 6285 -19790 6323 -19756
rect 6357 -19790 6404 -19756
rect 5916 -19796 6404 -19790
rect 6106 -19846 6166 -19796
rect 6100 -19850 6172 -19846
rect 6100 -19902 6110 -19850
rect 6162 -19902 6172 -19850
rect 6100 -19906 6172 -19902
rect 6640 -20062 6700 -19687
rect 7660 -19687 7670 -19660
rect 7704 -19660 7710 -19653
rect 8682 -19221 8728 -19183
rect 9688 -19149 9748 -18998
rect 10204 -19040 10264 -18894
rect 9988 -19046 10476 -19040
rect 9988 -19080 10035 -19046
rect 10069 -19080 10107 -19046
rect 10141 -19080 10179 -19046
rect 10213 -19080 10251 -19046
rect 10285 -19080 10323 -19046
rect 10357 -19080 10395 -19046
rect 10429 -19080 10476 -19046
rect 9988 -19086 10476 -19080
rect 9688 -19183 9706 -19149
rect 9740 -19183 9748 -19149
rect 10710 -19149 10770 -18672
rect 11218 -18834 11278 -18562
rect 11212 -18838 11284 -18834
rect 11212 -18890 11222 -18838
rect 11274 -18890 11284 -18838
rect 11212 -18894 11284 -18890
rect 11218 -19040 11278 -18894
rect 11730 -18938 11790 -18453
rect 12746 -18453 12760 -18440
rect 12794 -18440 12800 -18419
rect 13772 -17915 13818 -17884
rect 13772 -17949 13778 -17915
rect 13812 -17949 13818 -17915
rect 13772 -17987 13818 -17949
rect 13772 -18021 13778 -17987
rect 13812 -18021 13818 -17987
rect 13772 -18059 13818 -18021
rect 13772 -18093 13778 -18059
rect 13812 -18093 13818 -18059
rect 13772 -18131 13818 -18093
rect 13772 -18165 13778 -18131
rect 13812 -18165 13818 -18131
rect 13772 -18203 13818 -18165
rect 13772 -18237 13778 -18203
rect 13812 -18237 13818 -18203
rect 13772 -18275 13818 -18237
rect 13772 -18309 13778 -18275
rect 13812 -18309 13818 -18275
rect 13772 -18347 13818 -18309
rect 13772 -18381 13778 -18347
rect 13812 -18381 13818 -18347
rect 13772 -18419 13818 -18381
rect 13772 -18438 13778 -18419
rect 12794 -18453 12806 -18440
rect 12024 -18522 12512 -18516
rect 12024 -18556 12071 -18522
rect 12105 -18556 12143 -18522
rect 12177 -18556 12215 -18522
rect 12249 -18556 12287 -18522
rect 12321 -18556 12359 -18522
rect 12393 -18556 12431 -18522
rect 12465 -18556 12512 -18522
rect 12024 -18562 12512 -18556
rect 12226 -18834 12286 -18562
rect 12746 -18612 12806 -18453
rect 13768 -18453 13778 -18438
rect 13812 -18438 13818 -18419
rect 14790 -17915 14836 -17884
rect 14790 -17949 14796 -17915
rect 14830 -17949 14836 -17915
rect 14790 -17987 14836 -17949
rect 14790 -18021 14796 -17987
rect 14830 -18021 14836 -17987
rect 14790 -18059 14836 -18021
rect 14790 -18093 14796 -18059
rect 14830 -18093 14836 -18059
rect 14790 -18131 14836 -18093
rect 14790 -18165 14796 -18131
rect 14830 -18165 14836 -18131
rect 14790 -18203 14836 -18165
rect 14790 -18237 14796 -18203
rect 14830 -18237 14836 -18203
rect 14790 -18275 14836 -18237
rect 14790 -18309 14796 -18275
rect 14830 -18309 14836 -18275
rect 14790 -18347 14836 -18309
rect 14790 -18381 14796 -18347
rect 14830 -18381 14836 -18347
rect 14790 -18419 14836 -18381
rect 13812 -18453 13828 -18438
rect 14790 -18440 14796 -18419
rect 13042 -18522 13530 -18516
rect 13042 -18556 13089 -18522
rect 13123 -18556 13161 -18522
rect 13195 -18556 13233 -18522
rect 13267 -18556 13305 -18522
rect 13339 -18556 13377 -18522
rect 13411 -18556 13449 -18522
rect 13483 -18556 13530 -18522
rect 13042 -18562 13530 -18556
rect 12740 -18616 12812 -18612
rect 12740 -18668 12750 -18616
rect 12802 -18668 12812 -18616
rect 12740 -18672 12812 -18668
rect 13270 -18834 13330 -18562
rect 12220 -18838 12292 -18834
rect 12220 -18890 12230 -18838
rect 12282 -18890 12292 -18838
rect 12220 -18894 12292 -18890
rect 13264 -18838 13336 -18834
rect 13264 -18890 13274 -18838
rect 13326 -18890 13336 -18838
rect 13264 -18894 13336 -18890
rect 11724 -18942 11796 -18938
rect 11724 -18994 11734 -18942
rect 11786 -18994 11796 -18942
rect 11724 -18998 11796 -18994
rect 11006 -19046 11494 -19040
rect 11006 -19080 11053 -19046
rect 11087 -19080 11125 -19046
rect 11159 -19080 11197 -19046
rect 11231 -19080 11269 -19046
rect 11303 -19080 11341 -19046
rect 11375 -19080 11413 -19046
rect 11447 -19080 11494 -19046
rect 11006 -19086 11494 -19080
rect 10710 -19166 10724 -19149
rect 9688 -19194 9748 -19183
rect 10718 -19183 10724 -19166
rect 10758 -19166 10770 -19149
rect 11730 -19149 11790 -18998
rect 12226 -19040 12286 -18894
rect 13270 -19040 13330 -18894
rect 13768 -18938 13828 -18453
rect 14782 -18453 14796 -18440
rect 14830 -18440 14836 -18419
rect 15802 -17915 15862 -17764
rect 16096 -17812 16584 -17806
rect 16096 -17846 16143 -17812
rect 16177 -17846 16215 -17812
rect 16249 -17846 16287 -17812
rect 16321 -17846 16359 -17812
rect 16393 -17846 16431 -17812
rect 16465 -17846 16503 -17812
rect 16537 -17846 16584 -17812
rect 16096 -17852 16584 -17846
rect 15802 -17949 15814 -17915
rect 15848 -17949 15862 -17915
rect 16818 -17915 16878 -17221
rect 17838 -17221 17850 -17206
rect 17884 -17206 17890 -17187
rect 18862 -16717 18868 -16706
rect 18902 -16706 18914 -16683
rect 19880 -16683 19926 -16652
rect 18902 -16717 18908 -16706
rect 18862 -16755 18908 -16717
rect 18862 -16789 18868 -16755
rect 18902 -16789 18908 -16755
rect 18862 -16827 18908 -16789
rect 18862 -16861 18868 -16827
rect 18902 -16861 18908 -16827
rect 18862 -16899 18908 -16861
rect 18862 -16933 18868 -16899
rect 18902 -16933 18908 -16899
rect 18862 -16971 18908 -16933
rect 18862 -17005 18868 -16971
rect 18902 -17005 18908 -16971
rect 18862 -17043 18908 -17005
rect 18862 -17077 18868 -17043
rect 18902 -17077 18908 -17043
rect 18862 -17115 18908 -17077
rect 18862 -17149 18868 -17115
rect 18902 -17149 18908 -17115
rect 18862 -17187 18908 -17149
rect 19880 -16717 19886 -16683
rect 19920 -16717 19926 -16683
rect 20892 -16683 20952 -16524
rect 21394 -16574 21454 -16096
rect 21910 -16134 21970 -15987
rect 22928 -15987 22940 -15953
rect 22974 -15987 22988 -15953
rect 22204 -16056 22692 -16050
rect 22204 -16090 22251 -16056
rect 22285 -16090 22323 -16056
rect 22357 -16090 22395 -16056
rect 22429 -16090 22467 -16056
rect 22501 -16090 22539 -16056
rect 22573 -16090 22611 -16056
rect 22645 -16090 22692 -16056
rect 22204 -16096 22692 -16090
rect 22928 -16116 22988 -15987
rect 22922 -16120 22994 -16116
rect 21904 -16138 21976 -16134
rect 21904 -16190 21914 -16138
rect 21966 -16190 21976 -16138
rect 22922 -16172 22932 -16120
rect 22984 -16172 22994 -16120
rect 22922 -16176 22994 -16172
rect 21904 -16194 21976 -16190
rect 21910 -16412 21970 -16194
rect 21910 -16472 22984 -16412
rect 23034 -16464 23094 -15288
rect 23522 -16250 23594 -16246
rect 23522 -16302 23532 -16250
rect 23584 -16302 23594 -16250
rect 23522 -16306 23594 -16302
rect 23272 -16354 23344 -16350
rect 23272 -16406 23282 -16354
rect 23334 -16406 23344 -16354
rect 23272 -16410 23344 -16406
rect 21186 -16580 21674 -16574
rect 21186 -16614 21233 -16580
rect 21267 -16614 21305 -16580
rect 21339 -16614 21377 -16580
rect 21411 -16614 21449 -16580
rect 21483 -16614 21521 -16580
rect 21555 -16614 21593 -16580
rect 21627 -16614 21674 -16580
rect 21186 -16620 21674 -16614
rect 20892 -16706 20904 -16683
rect 19880 -16755 19926 -16717
rect 19880 -16789 19886 -16755
rect 19920 -16789 19926 -16755
rect 19880 -16827 19926 -16789
rect 19880 -16861 19886 -16827
rect 19920 -16861 19926 -16827
rect 19880 -16899 19926 -16861
rect 19880 -16933 19886 -16899
rect 19920 -16933 19926 -16899
rect 19880 -16971 19926 -16933
rect 19880 -17005 19886 -16971
rect 19920 -17005 19926 -16971
rect 19880 -17043 19926 -17005
rect 19880 -17077 19886 -17043
rect 19920 -17077 19926 -17043
rect 19880 -17115 19926 -17077
rect 19880 -17149 19886 -17115
rect 19920 -17149 19926 -17115
rect 19880 -17182 19926 -17149
rect 20898 -16717 20904 -16706
rect 20938 -16706 20952 -16683
rect 21910 -16683 21970 -16472
rect 22414 -16574 22474 -16472
rect 22204 -16580 22692 -16574
rect 22204 -16614 22251 -16580
rect 22285 -16614 22323 -16580
rect 22357 -16614 22395 -16580
rect 22429 -16614 22467 -16580
rect 22501 -16614 22539 -16580
rect 22573 -16614 22611 -16580
rect 22645 -16614 22692 -16580
rect 22204 -16620 22692 -16614
rect 21910 -16698 21922 -16683
rect 20938 -16717 20944 -16706
rect 20898 -16755 20944 -16717
rect 20898 -16789 20904 -16755
rect 20938 -16789 20944 -16755
rect 20898 -16827 20944 -16789
rect 20898 -16861 20904 -16827
rect 20938 -16861 20944 -16827
rect 20898 -16899 20944 -16861
rect 20898 -16933 20904 -16899
rect 20938 -16933 20944 -16899
rect 20898 -16971 20944 -16933
rect 20898 -17005 20904 -16971
rect 20938 -17005 20944 -16971
rect 20898 -17043 20944 -17005
rect 20898 -17077 20904 -17043
rect 20938 -17077 20944 -17043
rect 20898 -17115 20944 -17077
rect 20898 -17149 20904 -17115
rect 20938 -17149 20944 -17115
rect 17884 -17221 17898 -17206
rect 17114 -17290 17602 -17284
rect 17114 -17324 17161 -17290
rect 17195 -17324 17233 -17290
rect 17267 -17324 17305 -17290
rect 17339 -17324 17377 -17290
rect 17411 -17324 17449 -17290
rect 17483 -17324 17521 -17290
rect 17555 -17324 17602 -17290
rect 17114 -17330 17602 -17324
rect 17314 -17600 17374 -17330
rect 17308 -17604 17380 -17600
rect 17308 -17656 17318 -17604
rect 17370 -17656 17380 -17604
rect 17308 -17660 17380 -17656
rect 17314 -17806 17374 -17660
rect 17114 -17812 17602 -17806
rect 17114 -17846 17161 -17812
rect 17195 -17846 17233 -17812
rect 17267 -17846 17305 -17812
rect 17339 -17846 17377 -17812
rect 17411 -17846 17449 -17812
rect 17483 -17846 17521 -17812
rect 17555 -17846 17602 -17812
rect 17114 -17852 17602 -17846
rect 16818 -17936 16832 -17915
rect 15802 -17987 15862 -17949
rect 15802 -18021 15814 -17987
rect 15848 -18021 15862 -17987
rect 15802 -18059 15862 -18021
rect 15802 -18093 15814 -18059
rect 15848 -18093 15862 -18059
rect 15802 -18131 15862 -18093
rect 15802 -18165 15814 -18131
rect 15848 -18165 15862 -18131
rect 15802 -18203 15862 -18165
rect 15802 -18237 15814 -18203
rect 15848 -18237 15862 -18203
rect 15802 -18275 15862 -18237
rect 15802 -18309 15814 -18275
rect 15848 -18309 15862 -18275
rect 15802 -18347 15862 -18309
rect 15802 -18381 15814 -18347
rect 15848 -18381 15862 -18347
rect 15802 -18419 15862 -18381
rect 14830 -18453 14842 -18440
rect 14060 -18522 14548 -18516
rect 14060 -18556 14107 -18522
rect 14141 -18556 14179 -18522
rect 14213 -18556 14251 -18522
rect 14285 -18556 14323 -18522
rect 14357 -18556 14395 -18522
rect 14429 -18556 14467 -18522
rect 14501 -18556 14548 -18522
rect 14060 -18562 14548 -18556
rect 14260 -18834 14320 -18562
rect 14782 -18612 14842 -18453
rect 15802 -18453 15814 -18419
rect 15848 -18453 15862 -18419
rect 16826 -17949 16832 -17936
rect 16866 -17936 16878 -17915
rect 17838 -17915 17898 -17221
rect 18862 -17221 18868 -17187
rect 18902 -17221 18908 -17187
rect 18862 -17252 18908 -17221
rect 19872 -17187 19932 -17182
rect 19872 -17221 19886 -17187
rect 19920 -17221 19932 -17187
rect 18344 -17284 18404 -17282
rect 18132 -17290 18620 -17284
rect 18132 -17324 18179 -17290
rect 18213 -17324 18251 -17290
rect 18285 -17324 18323 -17290
rect 18357 -17324 18395 -17290
rect 18429 -17324 18467 -17290
rect 18501 -17324 18539 -17290
rect 18573 -17324 18620 -17290
rect 18132 -17330 18620 -17324
rect 19150 -17290 19638 -17284
rect 19150 -17324 19197 -17290
rect 19231 -17324 19269 -17290
rect 19303 -17324 19341 -17290
rect 19375 -17324 19413 -17290
rect 19447 -17324 19485 -17290
rect 19519 -17324 19557 -17290
rect 19591 -17324 19638 -17290
rect 19150 -17330 19638 -17324
rect 18344 -17600 18404 -17330
rect 19366 -17378 19426 -17330
rect 19498 -17378 19570 -17374
rect 19360 -17382 19432 -17378
rect 19360 -17434 19370 -17382
rect 19422 -17434 19432 -17382
rect 19498 -17430 19508 -17378
rect 19560 -17430 19570 -17378
rect 19498 -17434 19570 -17430
rect 19360 -17438 19432 -17434
rect 19504 -17600 19564 -17434
rect 19872 -17600 19932 -17221
rect 20898 -17187 20944 -17149
rect 20898 -17221 20904 -17187
rect 20938 -17221 20944 -17187
rect 21916 -16717 21922 -16698
rect 21956 -16698 21970 -16683
rect 22924 -16683 22984 -16472
rect 23028 -16468 23100 -16464
rect 23028 -16520 23038 -16468
rect 23090 -16520 23100 -16468
rect 23028 -16524 23100 -16520
rect 22924 -16688 22940 -16683
rect 21956 -16717 21962 -16698
rect 21916 -16755 21962 -16717
rect 21916 -16789 21922 -16755
rect 21956 -16789 21962 -16755
rect 21916 -16827 21962 -16789
rect 21916 -16861 21922 -16827
rect 21956 -16861 21962 -16827
rect 21916 -16899 21962 -16861
rect 21916 -16933 21922 -16899
rect 21956 -16933 21962 -16899
rect 21916 -16971 21962 -16933
rect 21916 -17005 21922 -16971
rect 21956 -17005 21962 -16971
rect 21916 -17043 21962 -17005
rect 21916 -17077 21922 -17043
rect 21956 -17077 21962 -17043
rect 21916 -17115 21962 -17077
rect 21916 -17149 21922 -17115
rect 21956 -17149 21962 -17115
rect 21916 -17187 21962 -17149
rect 21916 -17200 21922 -17187
rect 20898 -17252 20944 -17221
rect 21910 -17221 21922 -17200
rect 21956 -17200 21962 -17187
rect 22934 -16717 22940 -16688
rect 22974 -16688 22984 -16683
rect 22974 -16717 22980 -16688
rect 22934 -16755 22980 -16717
rect 22934 -16789 22940 -16755
rect 22974 -16789 22980 -16755
rect 22934 -16827 22980 -16789
rect 22934 -16861 22940 -16827
rect 22974 -16861 22980 -16827
rect 22934 -16899 22980 -16861
rect 22934 -16933 22940 -16899
rect 22974 -16933 22980 -16899
rect 22934 -16971 22980 -16933
rect 22934 -17005 22940 -16971
rect 22974 -17005 22980 -16971
rect 22934 -17043 22980 -17005
rect 22934 -17077 22940 -17043
rect 22974 -17077 22980 -17043
rect 22934 -17115 22980 -17077
rect 22934 -17149 22940 -17115
rect 22974 -17149 22980 -17115
rect 22934 -17187 22980 -17149
rect 21956 -17221 21970 -17200
rect 20168 -17290 20656 -17284
rect 20168 -17324 20215 -17290
rect 20249 -17324 20287 -17290
rect 20321 -17324 20359 -17290
rect 20393 -17324 20431 -17290
rect 20465 -17324 20503 -17290
rect 20537 -17324 20575 -17290
rect 20609 -17324 20656 -17290
rect 20168 -17330 20656 -17324
rect 21186 -17290 21674 -17284
rect 21186 -17324 21233 -17290
rect 21267 -17324 21305 -17290
rect 21339 -17324 21521 -17290
rect 21555 -17324 21593 -17290
rect 21627 -17324 21674 -17290
rect 21186 -17330 21674 -17324
rect 21392 -17374 21452 -17330
rect 20380 -17378 20452 -17374
rect 20380 -17430 20390 -17378
rect 20442 -17430 20452 -17378
rect 20380 -17434 20452 -17430
rect 21386 -17378 21458 -17374
rect 21910 -17378 21970 -17221
rect 22934 -17221 22940 -17187
rect 22974 -17221 22980 -17187
rect 22934 -17252 22980 -17221
rect 22204 -17290 22692 -17284
rect 22204 -17324 22251 -17290
rect 22285 -17324 22323 -17290
rect 22357 -17324 22395 -17290
rect 22429 -17324 22467 -17290
rect 22501 -17324 22539 -17290
rect 22573 -17324 22611 -17290
rect 22645 -17324 22692 -17290
rect 22204 -17330 22692 -17324
rect 21386 -17430 21396 -17378
rect 21448 -17430 21458 -17378
rect 21386 -17434 21458 -17430
rect 21904 -17382 21976 -17378
rect 21904 -17434 21914 -17382
rect 21966 -17434 21976 -17382
rect 18338 -17604 18410 -17600
rect 18338 -17656 18348 -17604
rect 18400 -17656 18410 -17604
rect 18338 -17660 18410 -17656
rect 19498 -17604 19570 -17600
rect 19498 -17656 19508 -17604
rect 19560 -17656 19570 -17604
rect 19498 -17660 19570 -17656
rect 19866 -17604 19938 -17600
rect 19866 -17656 19876 -17604
rect 19928 -17656 19938 -17604
rect 19866 -17660 19938 -17656
rect 18344 -17806 18404 -17660
rect 19504 -17806 19564 -17660
rect 19872 -17704 19932 -17660
rect 19866 -17708 19938 -17704
rect 19866 -17760 19876 -17708
rect 19928 -17760 19938 -17708
rect 19866 -17764 19938 -17760
rect 20386 -17806 20446 -17434
rect 21904 -17438 21976 -17434
rect 21904 -17510 21976 -17506
rect 21904 -17562 21914 -17510
rect 21966 -17562 21976 -17510
rect 21904 -17566 21976 -17562
rect 20882 -17706 20954 -17702
rect 20882 -17758 20892 -17706
rect 20944 -17758 20954 -17706
rect 20882 -17762 20954 -17758
rect 18132 -17812 18620 -17806
rect 18132 -17846 18179 -17812
rect 18213 -17846 18251 -17812
rect 18285 -17846 18323 -17812
rect 18357 -17846 18395 -17812
rect 18429 -17846 18467 -17812
rect 18501 -17846 18539 -17812
rect 18573 -17846 18620 -17812
rect 18132 -17852 18620 -17846
rect 19150 -17812 19638 -17806
rect 19150 -17846 19197 -17812
rect 19231 -17846 19269 -17812
rect 19303 -17846 19341 -17812
rect 19375 -17846 19413 -17812
rect 19447 -17846 19485 -17812
rect 19519 -17846 19557 -17812
rect 19591 -17846 19638 -17812
rect 19150 -17852 19638 -17846
rect 20168 -17812 20656 -17806
rect 20168 -17846 20215 -17812
rect 20249 -17846 20287 -17812
rect 20321 -17846 20359 -17812
rect 20393 -17846 20431 -17812
rect 20465 -17846 20503 -17812
rect 20537 -17846 20575 -17812
rect 20609 -17846 20656 -17812
rect 20168 -17852 20656 -17846
rect 20386 -17854 20446 -17852
rect 16866 -17949 16872 -17936
rect 17838 -17942 17850 -17915
rect 16826 -17987 16872 -17949
rect 16826 -18021 16832 -17987
rect 16866 -18021 16872 -17987
rect 16826 -18059 16872 -18021
rect 16826 -18093 16832 -18059
rect 16866 -18093 16872 -18059
rect 16826 -18131 16872 -18093
rect 16826 -18165 16832 -18131
rect 16866 -18165 16872 -18131
rect 16826 -18203 16872 -18165
rect 16826 -18237 16832 -18203
rect 16866 -18237 16872 -18203
rect 16826 -18275 16872 -18237
rect 16826 -18309 16832 -18275
rect 16866 -18309 16872 -18275
rect 16826 -18347 16872 -18309
rect 16826 -18381 16832 -18347
rect 16866 -18381 16872 -18347
rect 16826 -18419 16872 -18381
rect 16826 -18440 16832 -18419
rect 15078 -18522 15566 -18516
rect 15078 -18556 15125 -18522
rect 15159 -18556 15197 -18522
rect 15231 -18556 15269 -18522
rect 15303 -18556 15341 -18522
rect 15375 -18556 15413 -18522
rect 15447 -18556 15485 -18522
rect 15519 -18556 15566 -18522
rect 15078 -18562 15566 -18556
rect 14776 -18616 14848 -18612
rect 14776 -18668 14786 -18616
rect 14838 -18668 14848 -18616
rect 14776 -18672 14848 -18668
rect 15278 -18834 15338 -18562
rect 14254 -18838 14326 -18834
rect 14254 -18890 14264 -18838
rect 14316 -18890 14326 -18838
rect 14254 -18894 14326 -18890
rect 15272 -18838 15344 -18834
rect 15272 -18890 15282 -18838
rect 15334 -18890 15344 -18838
rect 15272 -18894 15344 -18890
rect 13762 -18942 13834 -18938
rect 13762 -18994 13772 -18942
rect 13824 -18994 13834 -18942
rect 13762 -18998 13834 -18994
rect 12024 -19046 12512 -19040
rect 12024 -19080 12071 -19046
rect 12105 -19080 12143 -19046
rect 12177 -19080 12215 -19046
rect 12249 -19080 12287 -19046
rect 12321 -19080 12359 -19046
rect 12393 -19080 12431 -19046
rect 12465 -19080 12512 -19046
rect 12024 -19086 12512 -19080
rect 13042 -19046 13530 -19040
rect 13042 -19080 13089 -19046
rect 13123 -19080 13161 -19046
rect 13195 -19080 13233 -19046
rect 13267 -19080 13305 -19046
rect 13339 -19080 13377 -19046
rect 13411 -19080 13449 -19046
rect 13483 -19080 13530 -19046
rect 13042 -19086 13530 -19080
rect 10758 -19183 10764 -19166
rect 11730 -19168 11742 -19149
rect 8682 -19255 8688 -19221
rect 8722 -19255 8728 -19221
rect 8682 -19293 8728 -19255
rect 8682 -19327 8688 -19293
rect 8722 -19327 8728 -19293
rect 8682 -19365 8728 -19327
rect 8682 -19399 8688 -19365
rect 8722 -19399 8728 -19365
rect 8682 -19437 8728 -19399
rect 8682 -19471 8688 -19437
rect 8722 -19471 8728 -19437
rect 8682 -19509 8728 -19471
rect 8682 -19543 8688 -19509
rect 8722 -19543 8728 -19509
rect 8682 -19581 8728 -19543
rect 8682 -19615 8688 -19581
rect 8722 -19615 8728 -19581
rect 8682 -19653 8728 -19615
rect 7704 -19687 7720 -19660
rect 8682 -19662 8688 -19653
rect 6934 -19756 7422 -19750
rect 6934 -19790 6981 -19756
rect 7015 -19790 7053 -19756
rect 7087 -19790 7125 -19756
rect 7159 -19790 7197 -19756
rect 7231 -19790 7269 -19756
rect 7303 -19790 7341 -19756
rect 7375 -19790 7422 -19756
rect 6934 -19796 7422 -19790
rect 7144 -19846 7204 -19796
rect 7138 -19850 7210 -19846
rect 7138 -19902 7148 -19850
rect 7200 -19902 7210 -19850
rect 7138 -19906 7210 -19902
rect 6634 -20066 6706 -20062
rect 6634 -20118 6644 -20066
rect 6696 -20118 6706 -20066
rect 6634 -20122 6706 -20118
rect 5614 -20164 5686 -20160
rect 5614 -20216 5624 -20164
rect 5676 -20216 5686 -20164
rect 5614 -20220 5686 -20216
rect 7144 -20274 7204 -19906
rect 7660 -20160 7720 -19687
rect 8678 -19687 8688 -19662
rect 8722 -19662 8728 -19653
rect 9700 -19221 9746 -19194
rect 9700 -19255 9706 -19221
rect 9740 -19255 9746 -19221
rect 9700 -19293 9746 -19255
rect 9700 -19327 9706 -19293
rect 9740 -19327 9746 -19293
rect 9700 -19365 9746 -19327
rect 9700 -19399 9706 -19365
rect 9740 -19399 9746 -19365
rect 9700 -19437 9746 -19399
rect 9700 -19471 9706 -19437
rect 9740 -19471 9746 -19437
rect 9700 -19509 9746 -19471
rect 9700 -19543 9706 -19509
rect 9740 -19543 9746 -19509
rect 9700 -19581 9746 -19543
rect 9700 -19615 9706 -19581
rect 9740 -19615 9746 -19581
rect 9700 -19653 9746 -19615
rect 10718 -19221 10764 -19183
rect 10718 -19255 10724 -19221
rect 10758 -19255 10764 -19221
rect 10718 -19293 10764 -19255
rect 10718 -19327 10724 -19293
rect 10758 -19327 10764 -19293
rect 10718 -19365 10764 -19327
rect 10718 -19399 10724 -19365
rect 10758 -19399 10764 -19365
rect 10718 -19437 10764 -19399
rect 10718 -19471 10724 -19437
rect 10758 -19471 10764 -19437
rect 10718 -19509 10764 -19471
rect 10718 -19543 10724 -19509
rect 10758 -19543 10764 -19509
rect 10718 -19581 10764 -19543
rect 10718 -19615 10724 -19581
rect 10758 -19615 10764 -19581
rect 10718 -19648 10764 -19615
rect 11736 -19183 11742 -19168
rect 11776 -19168 11790 -19149
rect 12754 -19149 12800 -19118
rect 11776 -19183 11782 -19168
rect 11736 -19221 11782 -19183
rect 11736 -19255 11742 -19221
rect 11776 -19255 11782 -19221
rect 11736 -19293 11782 -19255
rect 11736 -19327 11742 -19293
rect 11776 -19327 11782 -19293
rect 11736 -19365 11782 -19327
rect 11736 -19399 11742 -19365
rect 11776 -19399 11782 -19365
rect 11736 -19437 11782 -19399
rect 11736 -19471 11742 -19437
rect 11776 -19471 11782 -19437
rect 11736 -19509 11782 -19471
rect 11736 -19543 11742 -19509
rect 11776 -19543 11782 -19509
rect 11736 -19581 11782 -19543
rect 11736 -19615 11742 -19581
rect 11776 -19615 11782 -19581
rect 8722 -19687 8738 -19662
rect 7952 -19756 8440 -19750
rect 7952 -19790 7999 -19756
rect 8033 -19790 8071 -19756
rect 8105 -19790 8143 -19756
rect 8177 -19790 8215 -19756
rect 8249 -19790 8287 -19756
rect 8321 -19790 8359 -19756
rect 8393 -19790 8440 -19756
rect 7952 -19796 8222 -19790
rect 8230 -19796 8440 -19790
rect 8162 -19846 8222 -19796
rect 8678 -19840 8738 -19687
rect 9700 -19687 9706 -19653
rect 9740 -19687 9746 -19653
rect 9700 -19718 9746 -19687
rect 10714 -19653 10774 -19648
rect 10714 -19687 10724 -19653
rect 10758 -19687 10774 -19653
rect 8970 -19756 9458 -19750
rect 8970 -19790 9017 -19756
rect 9051 -19790 9089 -19756
rect 9123 -19790 9161 -19756
rect 9195 -19790 9233 -19756
rect 9267 -19790 9305 -19756
rect 9339 -19790 9377 -19756
rect 9411 -19790 9458 -19756
rect 8970 -19796 9458 -19790
rect 9988 -19756 10476 -19750
rect 9988 -19790 10035 -19756
rect 10069 -19790 10107 -19756
rect 10141 -19790 10179 -19756
rect 10213 -19790 10251 -19756
rect 10285 -19790 10323 -19756
rect 10357 -19790 10395 -19756
rect 10429 -19790 10476 -19756
rect 9988 -19796 10476 -19790
rect 8672 -19844 8744 -19840
rect 8156 -19850 8228 -19846
rect 8156 -19902 8166 -19850
rect 8218 -19902 8228 -19850
rect 8672 -19896 8682 -19844
rect 8734 -19896 8744 -19844
rect 8672 -19900 8744 -19896
rect 10714 -19844 10774 -19687
rect 11736 -19653 11782 -19615
rect 11736 -19687 11742 -19653
rect 11776 -19687 11782 -19653
rect 12754 -19183 12760 -19149
rect 12794 -19183 12800 -19149
rect 13768 -19149 13828 -18998
rect 14260 -19040 14320 -18894
rect 15802 -18938 15862 -18453
rect 16820 -18453 16832 -18440
rect 16866 -18440 16872 -18419
rect 17844 -17949 17850 -17942
rect 17884 -17942 17898 -17915
rect 18862 -17915 18908 -17884
rect 17884 -17949 17890 -17942
rect 17844 -17987 17890 -17949
rect 17844 -18021 17850 -17987
rect 17884 -18021 17890 -17987
rect 17844 -18059 17890 -18021
rect 17844 -18093 17850 -18059
rect 17884 -18093 17890 -18059
rect 17844 -18131 17890 -18093
rect 17844 -18165 17850 -18131
rect 17884 -18165 17890 -18131
rect 17844 -18203 17890 -18165
rect 17844 -18237 17850 -18203
rect 17884 -18237 17890 -18203
rect 17844 -18275 17890 -18237
rect 17844 -18309 17850 -18275
rect 17884 -18309 17890 -18275
rect 17844 -18347 17890 -18309
rect 17844 -18381 17850 -18347
rect 17884 -18381 17890 -18347
rect 17844 -18419 17890 -18381
rect 17844 -18428 17850 -18419
rect 16866 -18453 16880 -18440
rect 16096 -18522 16584 -18516
rect 16096 -18556 16143 -18522
rect 16177 -18556 16215 -18522
rect 16249 -18556 16287 -18522
rect 16321 -18556 16359 -18522
rect 16393 -18556 16431 -18522
rect 16465 -18556 16503 -18522
rect 16537 -18556 16584 -18522
rect 16096 -18562 16584 -18556
rect 16312 -18834 16372 -18562
rect 16820 -18612 16880 -18453
rect 17836 -18453 17850 -18428
rect 17884 -18428 17890 -18419
rect 18862 -17949 18868 -17915
rect 18902 -17949 18908 -17915
rect 18862 -17987 18908 -17949
rect 18862 -18021 18868 -17987
rect 18902 -18021 18908 -17987
rect 18862 -18059 18908 -18021
rect 18862 -18093 18868 -18059
rect 18902 -18093 18908 -18059
rect 18862 -18131 18908 -18093
rect 18862 -18165 18868 -18131
rect 18902 -18165 18908 -18131
rect 18862 -18203 18908 -18165
rect 18862 -18237 18868 -18203
rect 18902 -18237 18908 -18203
rect 18862 -18275 18908 -18237
rect 18862 -18309 18868 -18275
rect 18902 -18309 18908 -18275
rect 18862 -18347 18908 -18309
rect 18862 -18381 18868 -18347
rect 18902 -18381 18908 -18347
rect 18862 -18419 18908 -18381
rect 17884 -18453 17896 -18428
rect 18862 -18432 18868 -18419
rect 17114 -18522 17602 -18516
rect 17114 -18556 17161 -18522
rect 17195 -18556 17233 -18522
rect 17267 -18556 17305 -18522
rect 17339 -18556 17377 -18522
rect 17411 -18556 17449 -18522
rect 17483 -18556 17521 -18522
rect 17555 -18556 17602 -18522
rect 17114 -18562 17602 -18556
rect 16814 -18616 16886 -18612
rect 16814 -18668 16824 -18616
rect 16876 -18668 16886 -18616
rect 16814 -18672 16886 -18668
rect 16806 -18724 16878 -18720
rect 16806 -18776 16816 -18724
rect 16868 -18776 16878 -18724
rect 16806 -18780 16878 -18776
rect 16306 -18838 16378 -18834
rect 16306 -18890 16316 -18838
rect 16368 -18890 16378 -18838
rect 16306 -18894 16378 -18890
rect 15796 -18942 15868 -18938
rect 15796 -18994 15806 -18942
rect 15858 -18994 15868 -18942
rect 15796 -18998 15868 -18994
rect 16308 -18946 16380 -18942
rect 16308 -18998 16318 -18946
rect 16370 -18998 16380 -18946
rect 16308 -19002 16380 -18998
rect 16314 -19040 16374 -19002
rect 14060 -19046 14548 -19040
rect 14060 -19080 14107 -19046
rect 14141 -19080 14179 -19046
rect 14213 -19080 14251 -19046
rect 14285 -19080 14323 -19046
rect 14357 -19080 14395 -19046
rect 14429 -19080 14467 -19046
rect 14501 -19080 14548 -19046
rect 14060 -19086 14548 -19080
rect 15078 -19046 15566 -19040
rect 15078 -19080 15125 -19046
rect 15159 -19080 15197 -19046
rect 15231 -19080 15269 -19046
rect 15303 -19080 15341 -19046
rect 15375 -19080 15413 -19046
rect 15447 -19080 15485 -19046
rect 15519 -19080 15566 -19046
rect 15078 -19086 15566 -19080
rect 16096 -19046 16584 -19040
rect 16096 -19080 16143 -19046
rect 16177 -19080 16215 -19046
rect 16249 -19080 16287 -19046
rect 16321 -19080 16359 -19046
rect 16393 -19080 16431 -19046
rect 16465 -19080 16503 -19046
rect 16537 -19080 16584 -19046
rect 16096 -19086 16584 -19080
rect 13768 -19166 13778 -19149
rect 12754 -19221 12800 -19183
rect 12754 -19255 12760 -19221
rect 12794 -19255 12800 -19221
rect 12754 -19293 12800 -19255
rect 12754 -19327 12760 -19293
rect 12794 -19327 12800 -19293
rect 12754 -19365 12800 -19327
rect 12754 -19399 12760 -19365
rect 12794 -19399 12800 -19365
rect 12754 -19437 12800 -19399
rect 12754 -19471 12760 -19437
rect 12794 -19471 12800 -19437
rect 12754 -19509 12800 -19471
rect 12754 -19543 12760 -19509
rect 12794 -19543 12800 -19509
rect 12754 -19581 12800 -19543
rect 12754 -19615 12760 -19581
rect 12794 -19615 12800 -19581
rect 12754 -19653 12800 -19615
rect 12754 -19656 12760 -19653
rect 11736 -19718 11782 -19687
rect 12746 -19687 12760 -19656
rect 12794 -19656 12800 -19653
rect 13772 -19183 13778 -19166
rect 13812 -19166 13828 -19149
rect 14790 -19149 14836 -19118
rect 13812 -19183 13818 -19166
rect 13772 -19221 13818 -19183
rect 13772 -19255 13778 -19221
rect 13812 -19255 13818 -19221
rect 13772 -19293 13818 -19255
rect 13772 -19327 13778 -19293
rect 13812 -19327 13818 -19293
rect 13772 -19365 13818 -19327
rect 13772 -19399 13778 -19365
rect 13812 -19399 13818 -19365
rect 13772 -19437 13818 -19399
rect 13772 -19471 13778 -19437
rect 13812 -19471 13818 -19437
rect 13772 -19509 13818 -19471
rect 13772 -19543 13778 -19509
rect 13812 -19543 13818 -19509
rect 13772 -19581 13818 -19543
rect 13772 -19615 13778 -19581
rect 13812 -19615 13818 -19581
rect 13772 -19653 13818 -19615
rect 14790 -19183 14796 -19149
rect 14830 -19183 14836 -19149
rect 14790 -19221 14836 -19183
rect 14790 -19255 14796 -19221
rect 14830 -19255 14836 -19221
rect 14790 -19293 14836 -19255
rect 14790 -19327 14796 -19293
rect 14830 -19327 14836 -19293
rect 14790 -19365 14836 -19327
rect 14790 -19399 14796 -19365
rect 14830 -19399 14836 -19365
rect 14790 -19437 14836 -19399
rect 14790 -19471 14796 -19437
rect 14830 -19471 14836 -19437
rect 14790 -19509 14836 -19471
rect 14790 -19543 14796 -19509
rect 14830 -19543 14836 -19509
rect 14790 -19581 14836 -19543
rect 14790 -19615 14796 -19581
rect 14830 -19615 14836 -19581
rect 14790 -19644 14836 -19615
rect 15808 -19149 15854 -19118
rect 15808 -19183 15814 -19149
rect 15848 -19183 15854 -19149
rect 16812 -19149 16872 -18780
rect 17336 -18942 17396 -18562
rect 17836 -18936 17896 -18453
rect 18856 -18453 18868 -18432
rect 18902 -18432 18908 -18419
rect 19880 -17915 19926 -17884
rect 19880 -17949 19886 -17915
rect 19920 -17949 19926 -17915
rect 20888 -17915 20948 -17762
rect 21186 -17812 21674 -17806
rect 21186 -17846 21233 -17812
rect 21267 -17846 21305 -17812
rect 21339 -17846 21377 -17812
rect 21411 -17846 21449 -17812
rect 21483 -17846 21521 -17812
rect 21555 -17846 21593 -17812
rect 21627 -17846 21674 -17812
rect 21186 -17852 21674 -17846
rect 20888 -17946 20904 -17915
rect 19880 -17987 19926 -17949
rect 19880 -18021 19886 -17987
rect 19920 -18021 19926 -17987
rect 19880 -18059 19926 -18021
rect 19880 -18093 19886 -18059
rect 19920 -18093 19926 -18059
rect 19880 -18131 19926 -18093
rect 19880 -18165 19886 -18131
rect 19920 -18165 19926 -18131
rect 19880 -18203 19926 -18165
rect 19880 -18237 19886 -18203
rect 19920 -18237 19926 -18203
rect 19880 -18275 19926 -18237
rect 19880 -18309 19886 -18275
rect 19920 -18309 19926 -18275
rect 19880 -18347 19926 -18309
rect 19880 -18381 19886 -18347
rect 19920 -18381 19926 -18347
rect 19880 -18419 19926 -18381
rect 19880 -18428 19886 -18419
rect 18902 -18453 18916 -18432
rect 18132 -18522 18620 -18516
rect 18132 -18556 18179 -18522
rect 18213 -18556 18251 -18522
rect 18285 -18556 18323 -18522
rect 18357 -18556 18395 -18522
rect 18429 -18556 18467 -18522
rect 18501 -18556 18539 -18522
rect 18573 -18556 18620 -18522
rect 18132 -18562 18620 -18556
rect 17830 -18940 17902 -18936
rect 17330 -18946 17402 -18942
rect 17330 -18998 17340 -18946
rect 17392 -18998 17402 -18946
rect 17830 -18992 17840 -18940
rect 17892 -18992 17902 -18940
rect 17830 -18996 17902 -18992
rect 17330 -19002 17402 -18998
rect 17336 -19040 17396 -19002
rect 17114 -19046 17602 -19040
rect 17114 -19080 17161 -19046
rect 17195 -19080 17233 -19046
rect 17267 -19080 17305 -19046
rect 17339 -19080 17377 -19046
rect 17411 -19080 17449 -19046
rect 17483 -19080 17521 -19046
rect 17555 -19080 17602 -19046
rect 17114 -19086 17602 -19080
rect 16812 -19166 16832 -19149
rect 15808 -19221 15854 -19183
rect 15808 -19255 15814 -19221
rect 15848 -19255 15854 -19221
rect 15808 -19293 15854 -19255
rect 15808 -19327 15814 -19293
rect 15848 -19327 15854 -19293
rect 15808 -19365 15854 -19327
rect 15808 -19399 15814 -19365
rect 15848 -19399 15854 -19365
rect 15808 -19437 15854 -19399
rect 15808 -19471 15814 -19437
rect 15848 -19471 15854 -19437
rect 15808 -19509 15854 -19471
rect 15808 -19543 15814 -19509
rect 15848 -19543 15854 -19509
rect 15808 -19581 15854 -19543
rect 15808 -19615 15814 -19581
rect 15848 -19615 15854 -19581
rect 12794 -19687 12806 -19656
rect 11006 -19756 11494 -19750
rect 11006 -19790 11053 -19756
rect 11087 -19790 11125 -19756
rect 11159 -19790 11197 -19756
rect 11231 -19790 11269 -19756
rect 11303 -19790 11341 -19756
rect 11375 -19790 11413 -19756
rect 11447 -19790 11494 -19756
rect 11006 -19796 11494 -19790
rect 12024 -19756 12512 -19750
rect 12024 -19790 12071 -19756
rect 12105 -19790 12143 -19756
rect 12177 -19790 12215 -19756
rect 12249 -19790 12287 -19756
rect 12321 -19790 12359 -19756
rect 12393 -19790 12431 -19756
rect 12465 -19790 12512 -19756
rect 12024 -19796 12512 -19790
rect 12746 -19840 12806 -19687
rect 13772 -19687 13778 -19653
rect 13812 -19687 13818 -19653
rect 13772 -19718 13818 -19687
rect 14780 -19653 14840 -19644
rect 14780 -19687 14796 -19653
rect 14830 -19687 14840 -19653
rect 15808 -19653 15854 -19615
rect 15808 -19664 15814 -19653
rect 13042 -19756 13530 -19750
rect 13042 -19790 13089 -19756
rect 13123 -19790 13161 -19756
rect 13195 -19790 13233 -19756
rect 13267 -19790 13305 -19756
rect 13339 -19790 13377 -19756
rect 13411 -19790 13449 -19756
rect 13483 -19790 13530 -19756
rect 13042 -19796 13530 -19790
rect 14060 -19756 14548 -19750
rect 14060 -19790 14107 -19756
rect 14141 -19790 14179 -19756
rect 14213 -19790 14251 -19756
rect 14285 -19790 14323 -19756
rect 14357 -19790 14395 -19756
rect 14429 -19790 14467 -19756
rect 14501 -19790 14548 -19756
rect 14060 -19796 14548 -19790
rect 14780 -19840 14840 -19687
rect 15802 -19687 15814 -19664
rect 15848 -19664 15854 -19653
rect 16826 -19183 16832 -19166
rect 16866 -19183 16872 -19149
rect 16826 -19221 16872 -19183
rect 16826 -19255 16832 -19221
rect 16866 -19255 16872 -19221
rect 17836 -19149 17896 -18996
rect 18314 -19040 18374 -18562
rect 18856 -18612 18916 -18453
rect 19870 -18453 19886 -18428
rect 19920 -18428 19926 -18419
rect 20898 -17949 20904 -17946
rect 20938 -17946 20948 -17915
rect 21910 -17915 21970 -17566
rect 22204 -17812 22692 -17806
rect 22204 -17846 22251 -17812
rect 22285 -17846 22323 -17812
rect 22357 -17846 22395 -17812
rect 22429 -17846 22467 -17812
rect 22501 -17846 22539 -17812
rect 22573 -17846 22611 -17812
rect 22645 -17846 22692 -17812
rect 22204 -17852 22692 -17846
rect 20938 -17949 20944 -17946
rect 21910 -17948 21922 -17915
rect 20898 -17987 20944 -17949
rect 20898 -18021 20904 -17987
rect 20938 -18021 20944 -17987
rect 20898 -18059 20944 -18021
rect 20898 -18093 20904 -18059
rect 20938 -18093 20944 -18059
rect 20898 -18131 20944 -18093
rect 20898 -18165 20904 -18131
rect 20938 -18165 20944 -18131
rect 20898 -18203 20944 -18165
rect 20898 -18237 20904 -18203
rect 20938 -18237 20944 -18203
rect 20898 -18275 20944 -18237
rect 20898 -18309 20904 -18275
rect 20938 -18309 20944 -18275
rect 20898 -18347 20944 -18309
rect 20898 -18381 20904 -18347
rect 20938 -18381 20944 -18347
rect 20898 -18419 20944 -18381
rect 19920 -18453 19930 -18428
rect 20898 -18444 20904 -18419
rect 19150 -18522 19638 -18516
rect 19150 -18556 19197 -18522
rect 19231 -18556 19269 -18522
rect 19303 -18556 19341 -18522
rect 19375 -18556 19413 -18522
rect 19447 -18556 19485 -18522
rect 19519 -18556 19557 -18522
rect 19591 -18556 19638 -18522
rect 19150 -18562 19638 -18556
rect 18850 -18616 18922 -18612
rect 18850 -18668 18860 -18616
rect 18912 -18668 18922 -18616
rect 18850 -18672 18922 -18668
rect 18846 -18724 18918 -18720
rect 18846 -18776 18856 -18724
rect 18908 -18776 18918 -18724
rect 18846 -18780 18918 -18776
rect 18132 -19046 18620 -19040
rect 18132 -19080 18179 -19046
rect 18213 -19080 18251 -19046
rect 18285 -19080 18323 -19046
rect 18357 -19080 18395 -19046
rect 18429 -19080 18467 -19046
rect 18501 -19080 18539 -19046
rect 18573 -19080 18620 -19046
rect 18132 -19086 18620 -19080
rect 17836 -19183 17850 -19149
rect 17884 -19183 17896 -19149
rect 17836 -19221 17896 -19183
rect 18852 -19149 18912 -18780
rect 19338 -18838 19410 -18834
rect 19338 -18890 19348 -18838
rect 19400 -18890 19410 -18838
rect 19338 -18894 19410 -18890
rect 19344 -19040 19404 -18894
rect 19870 -18936 19930 -18453
rect 20894 -18453 20904 -18444
rect 20938 -18444 20944 -18419
rect 21916 -17949 21922 -17948
rect 21956 -17948 21970 -17915
rect 22934 -17915 22980 -17884
rect 21956 -17949 21962 -17948
rect 21916 -17987 21962 -17949
rect 21916 -18021 21922 -17987
rect 21956 -18021 21962 -17987
rect 21916 -18059 21962 -18021
rect 21916 -18093 21922 -18059
rect 21956 -18093 21962 -18059
rect 21916 -18131 21962 -18093
rect 21916 -18165 21922 -18131
rect 21956 -18165 21962 -18131
rect 21916 -18203 21962 -18165
rect 21916 -18237 21922 -18203
rect 21956 -18237 21962 -18203
rect 21916 -18275 21962 -18237
rect 21916 -18309 21922 -18275
rect 21956 -18309 21962 -18275
rect 21916 -18347 21962 -18309
rect 21916 -18381 21922 -18347
rect 21956 -18381 21962 -18347
rect 21916 -18419 21962 -18381
rect 21916 -18444 21922 -18419
rect 20938 -18453 20954 -18444
rect 20168 -18522 20656 -18516
rect 20168 -18556 20215 -18522
rect 20249 -18556 20287 -18522
rect 20321 -18556 20359 -18522
rect 20393 -18556 20431 -18522
rect 20465 -18556 20503 -18522
rect 20537 -18556 20575 -18522
rect 20609 -18556 20656 -18522
rect 20168 -18562 20656 -18556
rect 20894 -18612 20954 -18453
rect 21910 -18453 21922 -18444
rect 21956 -18444 21962 -18419
rect 22934 -17949 22940 -17915
rect 22974 -17949 22980 -17915
rect 22934 -17987 22980 -17949
rect 22934 -18021 22940 -17987
rect 22974 -18021 22980 -17987
rect 22934 -18059 22980 -18021
rect 22934 -18093 22940 -18059
rect 22974 -18093 22980 -18059
rect 22934 -18131 22980 -18093
rect 22934 -18165 22940 -18131
rect 22974 -18165 22980 -18131
rect 22934 -18203 22980 -18165
rect 22934 -18237 22940 -18203
rect 22974 -18237 22980 -18203
rect 22934 -18275 22980 -18237
rect 22934 -18309 22940 -18275
rect 22974 -18309 22980 -18275
rect 22934 -18347 22980 -18309
rect 22934 -18381 22940 -18347
rect 22974 -18381 22980 -18347
rect 22934 -18419 22980 -18381
rect 22934 -18438 22940 -18419
rect 21956 -18453 21970 -18444
rect 21186 -18522 21674 -18516
rect 21186 -18556 21233 -18522
rect 21267 -18556 21305 -18522
rect 21339 -18556 21377 -18522
rect 21411 -18556 21449 -18522
rect 21483 -18556 21521 -18522
rect 21555 -18556 21593 -18522
rect 21627 -18556 21674 -18522
rect 21186 -18562 21674 -18556
rect 20888 -18616 20960 -18612
rect 20888 -18668 20898 -18616
rect 20950 -18668 20960 -18616
rect 20888 -18672 20960 -18668
rect 20884 -18724 20956 -18720
rect 20884 -18776 20894 -18724
rect 20946 -18776 20956 -18724
rect 20884 -18780 20956 -18776
rect 20376 -18838 20448 -18834
rect 20376 -18890 20386 -18838
rect 20438 -18890 20448 -18838
rect 20376 -18894 20448 -18890
rect 19864 -18940 19936 -18936
rect 19864 -18992 19874 -18940
rect 19926 -18992 19936 -18940
rect 19864 -18996 19936 -18992
rect 20382 -19040 20442 -18894
rect 19150 -19046 19638 -19040
rect 19150 -19080 19197 -19046
rect 19231 -19080 19269 -19046
rect 19303 -19080 19341 -19046
rect 19375 -19080 19413 -19046
rect 19447 -19080 19485 -19046
rect 19519 -19080 19557 -19046
rect 19591 -19080 19638 -19046
rect 19150 -19086 19638 -19080
rect 20168 -19046 20656 -19040
rect 20168 -19080 20215 -19046
rect 20249 -19080 20287 -19046
rect 20321 -19080 20359 -19046
rect 20393 -19080 20431 -19046
rect 20465 -19080 20503 -19046
rect 20537 -19080 20575 -19046
rect 20609 -19080 20656 -19046
rect 20168 -19086 20656 -19080
rect 18852 -19183 18868 -19149
rect 18902 -19183 18912 -19149
rect 18852 -19196 18912 -19183
rect 19880 -19149 19926 -19118
rect 19880 -19183 19886 -19149
rect 19920 -19183 19926 -19149
rect 20890 -19149 20950 -18780
rect 21408 -18834 21468 -18562
rect 21910 -18654 21970 -18453
rect 22924 -18453 22940 -18438
rect 22974 -18438 22980 -18419
rect 22974 -18453 22984 -18438
rect 22204 -18522 22692 -18516
rect 22204 -18556 22251 -18522
rect 22285 -18556 22323 -18522
rect 22357 -18556 22395 -18522
rect 22429 -18556 22467 -18522
rect 22501 -18556 22539 -18522
rect 22573 -18556 22611 -18522
rect 22645 -18556 22692 -18522
rect 22204 -18562 22692 -18556
rect 22418 -18654 22478 -18562
rect 22924 -18654 22984 -18453
rect 21910 -18714 22984 -18654
rect 21402 -18838 21474 -18834
rect 21402 -18890 21412 -18838
rect 21464 -18890 21474 -18838
rect 21402 -18894 21474 -18890
rect 21906 -18940 21978 -18936
rect 21906 -18992 21916 -18940
rect 21968 -18992 21978 -18940
rect 21906 -18996 21978 -18992
rect 21186 -19046 21674 -19040
rect 21186 -19080 21233 -19046
rect 21267 -19080 21305 -19046
rect 21339 -19080 21377 -19046
rect 21411 -19080 21449 -19046
rect 21483 -19080 21521 -19046
rect 21555 -19080 21593 -19046
rect 21627 -19080 21674 -19046
rect 21186 -19086 21674 -19080
rect 20890 -19182 20904 -19149
rect 17836 -19224 17850 -19221
rect 16826 -19293 16872 -19255
rect 16826 -19327 16832 -19293
rect 16866 -19327 16872 -19293
rect 16826 -19365 16872 -19327
rect 16826 -19399 16832 -19365
rect 16866 -19399 16872 -19365
rect 16826 -19437 16872 -19399
rect 16826 -19471 16832 -19437
rect 16866 -19471 16872 -19437
rect 16826 -19509 16872 -19471
rect 16826 -19543 16832 -19509
rect 16866 -19543 16872 -19509
rect 16826 -19581 16872 -19543
rect 16826 -19615 16832 -19581
rect 16866 -19615 16872 -19581
rect 16826 -19653 16872 -19615
rect 15848 -19687 15862 -19664
rect 15078 -19756 15566 -19750
rect 15078 -19790 15125 -19756
rect 15159 -19790 15197 -19756
rect 15231 -19790 15269 -19756
rect 15303 -19790 15341 -19756
rect 15375 -19790 15413 -19756
rect 15447 -19790 15485 -19756
rect 15519 -19790 15566 -19756
rect 15078 -19796 15566 -19790
rect 10714 -19896 10718 -19844
rect 10770 -19896 10774 -19844
rect 8156 -19906 8228 -19902
rect 7654 -20164 7726 -20160
rect 7654 -20216 7664 -20164
rect 7716 -20216 7726 -20164
rect 7654 -20220 7726 -20216
rect 3880 -20280 4368 -20274
rect 3880 -20314 3927 -20280
rect 3961 -20314 3999 -20280
rect 4033 -20314 4071 -20280
rect 4105 -20314 4143 -20280
rect 4177 -20314 4215 -20280
rect 4249 -20314 4287 -20280
rect 4321 -20314 4368 -20280
rect 3880 -20320 4368 -20314
rect 4898 -20280 5386 -20274
rect 4898 -20314 4945 -20280
rect 4979 -20314 5017 -20280
rect 5051 -20314 5089 -20280
rect 5123 -20314 5161 -20280
rect 5195 -20314 5233 -20280
rect 5267 -20314 5305 -20280
rect 5339 -20314 5386 -20280
rect 4898 -20320 5386 -20314
rect 5916 -20280 6404 -20274
rect 5916 -20314 5963 -20280
rect 5997 -20314 6035 -20280
rect 6069 -20314 6107 -20280
rect 6141 -20314 6179 -20280
rect 6213 -20314 6251 -20280
rect 6285 -20314 6323 -20280
rect 6357 -20314 6404 -20280
rect 5916 -20320 6404 -20314
rect 6934 -20280 7422 -20274
rect 6934 -20314 6981 -20280
rect 7015 -20314 7053 -20280
rect 7087 -20314 7125 -20280
rect 7159 -20314 7197 -20280
rect 7231 -20314 7269 -20280
rect 7303 -20314 7341 -20280
rect 7375 -20314 7422 -20280
rect 6934 -20320 7422 -20314
rect 3582 -20417 3598 -20383
rect 3632 -20417 3642 -20383
rect 3582 -20418 3642 -20417
rect 4610 -20383 4656 -20352
rect 4610 -20417 4616 -20383
rect 4650 -20417 4656 -20383
rect 2574 -20489 2580 -20455
rect 2614 -20489 2620 -20455
rect 2574 -20527 2620 -20489
rect 2574 -20561 2580 -20527
rect 2614 -20561 2620 -20527
rect 2574 -20599 2620 -20561
rect 2574 -20633 2580 -20599
rect 2614 -20633 2620 -20599
rect 2574 -20671 2620 -20633
rect 2574 -20705 2580 -20671
rect 2614 -20705 2620 -20671
rect 2574 -20743 2620 -20705
rect 2574 -20777 2580 -20743
rect 2614 -20777 2620 -20743
rect 2574 -20815 2620 -20777
rect 2574 -20849 2580 -20815
rect 2614 -20849 2620 -20815
rect 2574 -20887 2620 -20849
rect 2574 -20906 2580 -20887
rect 2564 -20921 2580 -20906
rect 2614 -20906 2620 -20887
rect 3592 -20455 3638 -20418
rect 3592 -20489 3598 -20455
rect 3632 -20489 3638 -20455
rect 3592 -20527 3638 -20489
rect 3592 -20561 3598 -20527
rect 3632 -20561 3638 -20527
rect 3592 -20599 3638 -20561
rect 3592 -20633 3598 -20599
rect 3632 -20633 3638 -20599
rect 3592 -20671 3638 -20633
rect 3592 -20705 3598 -20671
rect 3632 -20705 3638 -20671
rect 3592 -20743 3638 -20705
rect 3592 -20777 3598 -20743
rect 3632 -20777 3638 -20743
rect 3592 -20815 3638 -20777
rect 3592 -20849 3598 -20815
rect 3632 -20849 3638 -20815
rect 3592 -20887 3638 -20849
rect 2614 -20921 2624 -20906
rect 3592 -20910 3598 -20887
rect 2564 -21072 2624 -20921
rect 3588 -20921 3598 -20910
rect 3632 -20910 3638 -20887
rect 4610 -20455 4656 -20417
rect 4610 -20489 4616 -20455
rect 4650 -20489 4656 -20455
rect 4610 -20527 4656 -20489
rect 4610 -20561 4616 -20527
rect 4650 -20561 4656 -20527
rect 4610 -20599 4656 -20561
rect 4610 -20633 4616 -20599
rect 4650 -20633 4656 -20599
rect 4610 -20671 4656 -20633
rect 4610 -20705 4616 -20671
rect 4650 -20705 4656 -20671
rect 4610 -20743 4656 -20705
rect 4610 -20777 4616 -20743
rect 4650 -20777 4656 -20743
rect 4610 -20815 4656 -20777
rect 4610 -20849 4616 -20815
rect 4650 -20849 4656 -20815
rect 4610 -20887 4656 -20849
rect 4610 -20894 4616 -20887
rect 3632 -20921 3648 -20910
rect 2862 -20990 3350 -20984
rect 2862 -21024 2909 -20990
rect 2943 -21024 2981 -20990
rect 3015 -21024 3053 -20990
rect 3087 -21024 3125 -20990
rect 3159 -21024 3197 -20990
rect 3231 -21024 3269 -20990
rect 3303 -21024 3350 -20990
rect 2862 -21030 3350 -21024
rect 3084 -21072 3144 -21030
rect 3588 -21072 3648 -20921
rect 4602 -20921 4616 -20894
rect 4650 -20894 4656 -20887
rect 5628 -20383 5674 -20352
rect 5628 -20417 5634 -20383
rect 5668 -20417 5674 -20383
rect 5628 -20455 5674 -20417
rect 5628 -20489 5634 -20455
rect 5668 -20489 5674 -20455
rect 5628 -20527 5674 -20489
rect 5628 -20561 5634 -20527
rect 5668 -20561 5674 -20527
rect 5628 -20599 5674 -20561
rect 5628 -20633 5634 -20599
rect 5668 -20633 5674 -20599
rect 5628 -20671 5674 -20633
rect 5628 -20705 5634 -20671
rect 5668 -20705 5674 -20671
rect 5628 -20743 5674 -20705
rect 5628 -20777 5634 -20743
rect 5668 -20777 5674 -20743
rect 5628 -20815 5674 -20777
rect 5628 -20849 5634 -20815
rect 5668 -20849 5674 -20815
rect 5628 -20887 5674 -20849
rect 4650 -20921 4662 -20894
rect 5628 -20910 5634 -20887
rect 3880 -20990 4368 -20984
rect 3880 -21024 3927 -20990
rect 3961 -21024 3999 -20990
rect 4033 -21024 4071 -20990
rect 4105 -21024 4143 -20990
rect 4177 -21024 4215 -20990
rect 4249 -21024 4287 -20990
rect 4321 -21024 4368 -20990
rect 3880 -21030 4368 -21024
rect 2564 -21132 3648 -21072
rect 2442 -21186 2514 -21182
rect 2442 -21238 2452 -21186
rect 2504 -21238 2514 -21186
rect 2442 -21242 2514 -21238
rect 3588 -21278 3648 -21132
rect 2564 -21338 3648 -21278
rect 2564 -21615 2624 -21338
rect 3076 -21506 3136 -21338
rect 3588 -21398 3648 -21338
rect 3582 -21402 3654 -21398
rect 3582 -21454 3592 -21402
rect 3644 -21454 3654 -21402
rect 3582 -21458 3654 -21454
rect 2862 -21512 3350 -21506
rect 2862 -21546 2909 -21512
rect 2943 -21546 2981 -21512
rect 3015 -21546 3053 -21512
rect 3087 -21546 3125 -21512
rect 3159 -21546 3197 -21512
rect 3231 -21546 3269 -21512
rect 3303 -21546 3350 -21512
rect 2862 -21552 3350 -21546
rect 2564 -21632 2580 -21615
rect 2574 -21649 2580 -21632
rect 2614 -21632 2624 -21615
rect 3588 -21615 3648 -21458
rect 4080 -21506 4140 -21030
rect 4602 -21084 4662 -20921
rect 5620 -20921 5634 -20910
rect 5668 -20910 5674 -20887
rect 6646 -20383 6692 -20352
rect 6646 -20417 6652 -20383
rect 6686 -20417 6692 -20383
rect 7660 -20383 7720 -20220
rect 8162 -20274 8222 -19906
rect 7952 -20280 8440 -20274
rect 7952 -20314 7999 -20280
rect 8033 -20314 8071 -20280
rect 8105 -20314 8143 -20280
rect 8177 -20314 8215 -20280
rect 8249 -20314 8287 -20280
rect 8321 -20314 8359 -20280
rect 8393 -20314 8440 -20280
rect 7952 -20320 8440 -20314
rect 7660 -20394 7670 -20383
rect 6646 -20455 6692 -20417
rect 6646 -20489 6652 -20455
rect 6686 -20489 6692 -20455
rect 6646 -20527 6692 -20489
rect 6646 -20561 6652 -20527
rect 6686 -20561 6692 -20527
rect 6646 -20599 6692 -20561
rect 6646 -20633 6652 -20599
rect 6686 -20633 6692 -20599
rect 6646 -20671 6692 -20633
rect 6646 -20705 6652 -20671
rect 6686 -20705 6692 -20671
rect 6646 -20743 6692 -20705
rect 6646 -20777 6652 -20743
rect 6686 -20777 6692 -20743
rect 6646 -20815 6692 -20777
rect 6646 -20849 6652 -20815
rect 6686 -20849 6692 -20815
rect 6646 -20887 6692 -20849
rect 7664 -20417 7670 -20394
rect 7704 -20394 7720 -20383
rect 8678 -20383 8738 -19900
rect 10714 -19906 10774 -19896
rect 12740 -19844 12812 -19840
rect 12740 -19896 12750 -19844
rect 12802 -19896 12812 -19844
rect 12740 -19900 12812 -19896
rect 14774 -19844 14846 -19840
rect 14774 -19896 14784 -19844
rect 14836 -19896 14846 -19844
rect 14774 -19900 14846 -19896
rect 11724 -19954 11796 -19950
rect 11724 -20006 11734 -19954
rect 11786 -20006 11796 -19954
rect 11724 -20010 11796 -20006
rect 13760 -19954 13832 -19950
rect 13760 -20006 13770 -19954
rect 13822 -20006 13832 -19954
rect 13760 -20010 13832 -20006
rect 10706 -20066 10778 -20062
rect 10706 -20118 10716 -20066
rect 10768 -20118 10778 -20066
rect 10706 -20122 10778 -20118
rect 9690 -20164 9762 -20160
rect 9690 -20216 9700 -20164
rect 9752 -20216 9762 -20164
rect 9690 -20220 9762 -20216
rect 8970 -20280 9458 -20274
rect 8970 -20314 9017 -20280
rect 9051 -20314 9089 -20280
rect 9123 -20314 9161 -20280
rect 9195 -20314 9233 -20280
rect 9267 -20314 9305 -20280
rect 9339 -20314 9377 -20280
rect 9411 -20314 9458 -20280
rect 8970 -20320 9458 -20314
rect 7704 -20417 7710 -20394
rect 8678 -20406 8688 -20383
rect 7664 -20455 7710 -20417
rect 7664 -20489 7670 -20455
rect 7704 -20489 7710 -20455
rect 7664 -20527 7710 -20489
rect 7664 -20561 7670 -20527
rect 7704 -20561 7710 -20527
rect 7664 -20599 7710 -20561
rect 7664 -20633 7670 -20599
rect 7704 -20633 7710 -20599
rect 7664 -20671 7710 -20633
rect 7664 -20705 7670 -20671
rect 7704 -20705 7710 -20671
rect 7664 -20743 7710 -20705
rect 7664 -20777 7670 -20743
rect 7704 -20777 7710 -20743
rect 7664 -20815 7710 -20777
rect 7664 -20849 7670 -20815
rect 7704 -20849 7710 -20815
rect 7664 -20876 7710 -20849
rect 8682 -20417 8688 -20406
rect 8722 -20406 8738 -20383
rect 9696 -20383 9756 -20220
rect 9988 -20280 10476 -20274
rect 9988 -20314 10035 -20280
rect 10069 -20314 10107 -20280
rect 10141 -20314 10179 -20280
rect 10213 -20314 10251 -20280
rect 10285 -20314 10323 -20280
rect 10357 -20314 10395 -20280
rect 10429 -20314 10476 -20280
rect 9988 -20320 10476 -20314
rect 9696 -20400 9706 -20383
rect 8722 -20417 8728 -20406
rect 8682 -20455 8728 -20417
rect 8682 -20489 8688 -20455
rect 8722 -20489 8728 -20455
rect 8682 -20527 8728 -20489
rect 8682 -20561 8688 -20527
rect 8722 -20561 8728 -20527
rect 8682 -20599 8728 -20561
rect 8682 -20633 8688 -20599
rect 8722 -20633 8728 -20599
rect 8682 -20671 8728 -20633
rect 8682 -20705 8688 -20671
rect 8722 -20705 8728 -20671
rect 8682 -20743 8728 -20705
rect 8682 -20777 8688 -20743
rect 8722 -20777 8728 -20743
rect 8682 -20815 8728 -20777
rect 8682 -20849 8688 -20815
rect 8722 -20849 8728 -20815
rect 6646 -20898 6652 -20887
rect 5668 -20921 5680 -20910
rect 4898 -20990 5386 -20984
rect 4898 -21024 4945 -20990
rect 4979 -21024 5017 -20990
rect 5051 -21024 5089 -20990
rect 5123 -21024 5161 -20990
rect 5195 -21024 5233 -20990
rect 5267 -21024 5305 -20990
rect 5339 -21024 5386 -20990
rect 4898 -21030 5386 -21024
rect 4596 -21088 4668 -21084
rect 4596 -21140 4606 -21088
rect 4658 -21140 4668 -21088
rect 4596 -21144 4668 -21140
rect 4600 -21282 4672 -21278
rect 4600 -21334 4610 -21282
rect 4662 -21334 4672 -21282
rect 4600 -21338 4672 -21334
rect 3880 -21512 4368 -21506
rect 3880 -21546 3927 -21512
rect 3961 -21546 3999 -21512
rect 4033 -21546 4071 -21512
rect 4105 -21546 4143 -21512
rect 4177 -21546 4215 -21512
rect 4249 -21546 4287 -21512
rect 4321 -21546 4368 -21512
rect 3880 -21552 4368 -21546
rect 2614 -21649 2620 -21632
rect 3588 -21636 3598 -21615
rect 2574 -21687 2620 -21649
rect 2574 -21721 2580 -21687
rect 2614 -21721 2620 -21687
rect 2574 -21759 2620 -21721
rect 2574 -21793 2580 -21759
rect 2614 -21793 2620 -21759
rect 2574 -21831 2620 -21793
rect 2574 -21865 2580 -21831
rect 2614 -21865 2620 -21831
rect 2574 -21903 2620 -21865
rect 2574 -21937 2580 -21903
rect 2614 -21937 2620 -21903
rect 2574 -21975 2620 -21937
rect 2574 -22009 2580 -21975
rect 2614 -22009 2620 -21975
rect 2574 -22047 2620 -22009
rect 2574 -22081 2580 -22047
rect 2614 -22081 2620 -22047
rect 2574 -22119 2620 -22081
rect 2574 -22153 2580 -22119
rect 2614 -22153 2620 -22119
rect 2574 -22184 2620 -22153
rect 3592 -21649 3598 -21636
rect 3632 -21636 3648 -21615
rect 4606 -21615 4666 -21338
rect 5100 -21342 5160 -21030
rect 5620 -21182 5680 -20921
rect 6638 -20921 6652 -20898
rect 6686 -20898 6692 -20887
rect 7656 -20887 7716 -20876
rect 6686 -20921 6698 -20898
rect 5916 -20990 6404 -20984
rect 5916 -21024 5963 -20990
rect 5997 -21024 6035 -20990
rect 6069 -21024 6107 -20990
rect 6141 -21024 6179 -20990
rect 6213 -21024 6251 -20990
rect 6285 -21024 6323 -20990
rect 6357 -21024 6404 -20990
rect 5916 -21030 6404 -21024
rect 5614 -21186 5686 -21182
rect 5614 -21238 5624 -21186
rect 5676 -21238 5686 -21186
rect 5614 -21242 5686 -21238
rect 6134 -21342 6194 -21030
rect 6638 -21084 6698 -20921
rect 7656 -20921 7670 -20887
rect 7704 -20921 7716 -20887
rect 8682 -20887 8728 -20849
rect 8682 -20900 8688 -20887
rect 6934 -20990 7422 -20984
rect 6934 -21024 6981 -20990
rect 7015 -21024 7053 -20990
rect 7087 -21024 7125 -20990
rect 7159 -21024 7197 -20990
rect 7231 -21024 7269 -20990
rect 7303 -21024 7341 -20990
rect 7375 -21024 7422 -20990
rect 6934 -21030 7422 -21024
rect 6632 -21088 6704 -21084
rect 6632 -21140 6642 -21088
rect 6694 -21140 6704 -21088
rect 6632 -21144 6704 -21140
rect 7144 -21182 7204 -21030
rect 7138 -21186 7210 -21182
rect 7138 -21238 7148 -21186
rect 7200 -21238 7210 -21186
rect 7138 -21242 7210 -21238
rect 6636 -21282 6708 -21278
rect 6636 -21334 6646 -21282
rect 6698 -21334 6708 -21282
rect 6636 -21338 6708 -21334
rect 5100 -21402 6194 -21342
rect 5100 -21506 5160 -21402
rect 6134 -21506 6194 -21402
rect 4898 -21512 5386 -21506
rect 4898 -21546 4945 -21512
rect 4979 -21546 5017 -21512
rect 5051 -21546 5089 -21512
rect 5123 -21546 5161 -21512
rect 5195 -21546 5233 -21512
rect 5267 -21546 5305 -21512
rect 5339 -21546 5386 -21512
rect 4898 -21552 5386 -21546
rect 5916 -21512 6404 -21506
rect 5916 -21546 5963 -21512
rect 5997 -21546 6035 -21512
rect 6069 -21546 6107 -21512
rect 6141 -21546 6179 -21512
rect 6213 -21546 6251 -21512
rect 6285 -21546 6323 -21512
rect 6357 -21546 6404 -21512
rect 5916 -21552 6404 -21546
rect 3632 -21649 3638 -21636
rect 4606 -21640 4616 -21615
rect 3592 -21687 3638 -21649
rect 3592 -21721 3598 -21687
rect 3632 -21721 3638 -21687
rect 3592 -21759 3638 -21721
rect 3592 -21793 3598 -21759
rect 3632 -21793 3638 -21759
rect 3592 -21831 3638 -21793
rect 3592 -21865 3598 -21831
rect 3632 -21865 3638 -21831
rect 3592 -21903 3638 -21865
rect 3592 -21937 3598 -21903
rect 3632 -21937 3638 -21903
rect 3592 -21975 3638 -21937
rect 3592 -22009 3598 -21975
rect 3632 -22009 3638 -21975
rect 3592 -22047 3638 -22009
rect 3592 -22081 3598 -22047
rect 3632 -22081 3638 -22047
rect 3592 -22119 3638 -22081
rect 3592 -22153 3598 -22119
rect 3632 -22153 3638 -22119
rect 3592 -22184 3638 -22153
rect 4610 -21649 4616 -21640
rect 4650 -21640 4666 -21615
rect 5628 -21615 5674 -21584
rect 4650 -21649 4656 -21640
rect 4610 -21687 4656 -21649
rect 4610 -21721 4616 -21687
rect 4650 -21721 4656 -21687
rect 4610 -21759 4656 -21721
rect 4610 -21793 4616 -21759
rect 4650 -21793 4656 -21759
rect 4610 -21831 4656 -21793
rect 4610 -21865 4616 -21831
rect 4650 -21865 4656 -21831
rect 4610 -21903 4656 -21865
rect 4610 -21937 4616 -21903
rect 4650 -21937 4656 -21903
rect 4610 -21975 4656 -21937
rect 4610 -22009 4616 -21975
rect 4650 -22009 4656 -21975
rect 4610 -22047 4656 -22009
rect 4610 -22081 4616 -22047
rect 4650 -22081 4656 -22047
rect 4610 -22119 4656 -22081
rect 4610 -22153 4616 -22119
rect 4650 -22153 4656 -22119
rect 5628 -21649 5634 -21615
rect 5668 -21649 5674 -21615
rect 6642 -21615 6702 -21338
rect 7144 -21506 7204 -21242
rect 7656 -21398 7716 -20921
rect 8676 -20921 8688 -20900
rect 8722 -20900 8728 -20887
rect 9700 -20417 9706 -20400
rect 9740 -20400 9756 -20383
rect 10712 -20383 10772 -20122
rect 11006 -20280 11494 -20274
rect 11006 -20314 11053 -20280
rect 11087 -20314 11125 -20280
rect 11159 -20314 11197 -20280
rect 11231 -20314 11269 -20280
rect 11303 -20314 11341 -20280
rect 11375 -20314 11413 -20280
rect 11447 -20314 11494 -20280
rect 11006 -20320 11494 -20314
rect 10712 -20390 10724 -20383
rect 9740 -20417 9746 -20400
rect 9700 -20455 9746 -20417
rect 9700 -20489 9706 -20455
rect 9740 -20489 9746 -20455
rect 9700 -20527 9746 -20489
rect 9700 -20561 9706 -20527
rect 9740 -20561 9746 -20527
rect 9700 -20599 9746 -20561
rect 9700 -20633 9706 -20599
rect 9740 -20633 9746 -20599
rect 9700 -20671 9746 -20633
rect 9700 -20705 9706 -20671
rect 9740 -20705 9746 -20671
rect 9700 -20743 9746 -20705
rect 9700 -20777 9706 -20743
rect 9740 -20777 9746 -20743
rect 9700 -20815 9746 -20777
rect 9700 -20849 9706 -20815
rect 9740 -20849 9746 -20815
rect 9700 -20887 9746 -20849
rect 10718 -20417 10724 -20390
rect 10758 -20390 10772 -20383
rect 11730 -20383 11790 -20010
rect 12024 -20280 12512 -20274
rect 12024 -20314 12071 -20280
rect 12105 -20314 12143 -20280
rect 12177 -20314 12215 -20280
rect 12249 -20314 12287 -20280
rect 12321 -20314 12359 -20280
rect 12393 -20314 12431 -20280
rect 12465 -20314 12512 -20280
rect 12024 -20320 12512 -20314
rect 13042 -20280 13530 -20274
rect 13042 -20314 13089 -20280
rect 13123 -20314 13161 -20280
rect 13195 -20314 13233 -20280
rect 13267 -20314 13305 -20280
rect 13339 -20314 13377 -20280
rect 13411 -20314 13449 -20280
rect 13483 -20314 13530 -20280
rect 13042 -20320 13530 -20314
rect 10758 -20417 10764 -20390
rect 11730 -20396 11742 -20383
rect 10718 -20455 10764 -20417
rect 10718 -20489 10724 -20455
rect 10758 -20489 10764 -20455
rect 10718 -20527 10764 -20489
rect 10718 -20561 10724 -20527
rect 10758 -20561 10764 -20527
rect 10718 -20599 10764 -20561
rect 10718 -20633 10724 -20599
rect 10758 -20633 10764 -20599
rect 10718 -20671 10764 -20633
rect 10718 -20705 10724 -20671
rect 10758 -20705 10764 -20671
rect 10718 -20743 10764 -20705
rect 10718 -20777 10724 -20743
rect 10758 -20777 10764 -20743
rect 10718 -20815 10764 -20777
rect 10718 -20849 10724 -20815
rect 10758 -20849 10764 -20815
rect 10718 -20884 10764 -20849
rect 11736 -20417 11742 -20396
rect 11776 -20396 11790 -20383
rect 12754 -20383 12800 -20352
rect 11776 -20417 11782 -20396
rect 11736 -20455 11782 -20417
rect 11736 -20489 11742 -20455
rect 11776 -20489 11782 -20455
rect 11736 -20527 11782 -20489
rect 11736 -20561 11742 -20527
rect 11776 -20561 11782 -20527
rect 11736 -20599 11782 -20561
rect 11736 -20633 11742 -20599
rect 11776 -20633 11782 -20599
rect 11736 -20671 11782 -20633
rect 11736 -20705 11742 -20671
rect 11776 -20705 11782 -20671
rect 11736 -20743 11782 -20705
rect 11736 -20777 11742 -20743
rect 11776 -20777 11782 -20743
rect 11736 -20815 11782 -20777
rect 11736 -20849 11742 -20815
rect 11776 -20849 11782 -20815
rect 8722 -20921 8736 -20900
rect 9700 -20906 9706 -20887
rect 7952 -20990 8440 -20984
rect 7952 -21024 7999 -20990
rect 8033 -21024 8071 -20990
rect 8105 -21024 8143 -20990
rect 8177 -21024 8215 -20990
rect 8249 -21024 8287 -20990
rect 8321 -21024 8359 -20990
rect 8393 -21024 8440 -20990
rect 7952 -21030 8440 -21024
rect 8166 -21186 8226 -21030
rect 8676 -21084 8736 -20921
rect 9690 -20921 9706 -20906
rect 9740 -20906 9746 -20887
rect 10708 -20887 10768 -20884
rect 9740 -20921 9750 -20906
rect 8970 -20990 9458 -20984
rect 8970 -21024 9017 -20990
rect 9051 -21024 9089 -20990
rect 9123 -21024 9161 -20990
rect 9195 -21024 9233 -20990
rect 9267 -21024 9305 -20990
rect 9339 -21024 9377 -20990
rect 9411 -21024 9458 -20990
rect 8970 -21030 9458 -21024
rect 8670 -21088 8742 -21084
rect 8670 -21140 8680 -21088
rect 8732 -21140 8742 -21088
rect 8670 -21144 8742 -21140
rect 9190 -21176 9250 -21030
rect 8166 -21238 8170 -21186
rect 8222 -21238 8226 -21186
rect 7650 -21402 7722 -21398
rect 7650 -21454 7660 -21402
rect 7712 -21454 7722 -21402
rect 7650 -21458 7722 -21454
rect 6934 -21512 7422 -21506
rect 6934 -21546 6981 -21512
rect 7015 -21546 7053 -21512
rect 7087 -21546 7125 -21512
rect 7159 -21546 7197 -21512
rect 7231 -21546 7269 -21512
rect 7303 -21546 7341 -21512
rect 7375 -21546 7422 -21512
rect 6934 -21552 7422 -21546
rect 6642 -21648 6652 -21615
rect 5628 -21687 5674 -21649
rect 5628 -21721 5634 -21687
rect 5668 -21721 5674 -21687
rect 5628 -21759 5674 -21721
rect 5628 -21793 5634 -21759
rect 5668 -21793 5674 -21759
rect 5628 -21831 5674 -21793
rect 5628 -21865 5634 -21831
rect 5668 -21865 5674 -21831
rect 5628 -21903 5674 -21865
rect 5628 -21937 5634 -21903
rect 5668 -21937 5674 -21903
rect 5628 -21975 5674 -21937
rect 5628 -22009 5634 -21975
rect 5668 -22009 5674 -21975
rect 5628 -22047 5674 -22009
rect 5628 -22081 5634 -22047
rect 5668 -22081 5674 -22047
rect 5628 -22119 5674 -22081
rect 5628 -22130 5634 -22119
rect 4610 -22184 4656 -22153
rect 5620 -22153 5634 -22130
rect 5668 -22130 5674 -22119
rect 6646 -21649 6652 -21648
rect 6686 -21648 6702 -21615
rect 7656 -21615 7716 -21458
rect 8166 -21506 8226 -21238
rect 9188 -21186 9250 -21176
rect 9188 -21238 9192 -21186
rect 9244 -21238 9250 -21186
rect 9188 -21248 9250 -21238
rect 8664 -21282 8736 -21278
rect 8664 -21334 8674 -21282
rect 8726 -21334 8736 -21282
rect 8664 -21338 8736 -21334
rect 7952 -21512 8440 -21506
rect 7952 -21546 7999 -21512
rect 8033 -21546 8071 -21512
rect 8105 -21546 8143 -21512
rect 8177 -21546 8215 -21512
rect 8249 -21546 8287 -21512
rect 8321 -21546 8359 -21512
rect 8393 -21546 8440 -21512
rect 7952 -21552 8440 -21546
rect 7656 -21636 7670 -21615
rect 6686 -21649 6692 -21648
rect 6646 -21687 6692 -21649
rect 6646 -21721 6652 -21687
rect 6686 -21721 6692 -21687
rect 6646 -21759 6692 -21721
rect 6646 -21793 6652 -21759
rect 6686 -21793 6692 -21759
rect 6646 -21831 6692 -21793
rect 6646 -21865 6652 -21831
rect 6686 -21865 6692 -21831
rect 6646 -21903 6692 -21865
rect 6646 -21937 6652 -21903
rect 6686 -21937 6692 -21903
rect 6646 -21975 6692 -21937
rect 6646 -22009 6652 -21975
rect 6686 -22009 6692 -21975
rect 6646 -22047 6692 -22009
rect 6646 -22081 6652 -22047
rect 6686 -22081 6692 -22047
rect 6646 -22119 6692 -22081
rect 7664 -21649 7670 -21636
rect 7704 -21636 7716 -21615
rect 8670 -21615 8730 -21338
rect 9190 -21506 9250 -21248
rect 9690 -21398 9750 -20921
rect 10708 -20921 10724 -20887
rect 10758 -20921 10768 -20887
rect 9988 -20990 10476 -20984
rect 9988 -21024 10035 -20990
rect 10069 -21024 10107 -20990
rect 10141 -21024 10179 -20990
rect 10213 -21024 10251 -20990
rect 10285 -21024 10323 -20990
rect 10357 -21024 10395 -20990
rect 10429 -21024 10476 -20990
rect 9988 -21030 10252 -21024
rect 10264 -21030 10476 -21024
rect 10192 -21182 10252 -21030
rect 10538 -21068 10598 -21058
rect 10708 -21064 10768 -20921
rect 11736 -20887 11782 -20849
rect 12754 -20417 12760 -20383
rect 12794 -20417 12800 -20383
rect 13766 -20383 13826 -20010
rect 15308 -20048 15368 -19796
rect 15802 -19838 15862 -19687
rect 16826 -19687 16832 -19653
rect 16866 -19687 16872 -19653
rect 17844 -19255 17850 -19224
rect 17884 -19224 17896 -19221
rect 18862 -19221 18908 -19196
rect 17884 -19255 17890 -19224
rect 17844 -19293 17890 -19255
rect 17844 -19327 17850 -19293
rect 17884 -19327 17890 -19293
rect 17844 -19365 17890 -19327
rect 17844 -19399 17850 -19365
rect 17884 -19399 17890 -19365
rect 17844 -19437 17890 -19399
rect 17844 -19471 17850 -19437
rect 17884 -19471 17890 -19437
rect 17844 -19509 17890 -19471
rect 17844 -19543 17850 -19509
rect 17884 -19543 17890 -19509
rect 17844 -19581 17890 -19543
rect 17844 -19615 17850 -19581
rect 17884 -19615 17890 -19581
rect 17844 -19653 17890 -19615
rect 17844 -19664 17850 -19653
rect 16826 -19718 16872 -19687
rect 17836 -19687 17850 -19664
rect 17884 -19664 17890 -19653
rect 18862 -19255 18868 -19221
rect 18902 -19255 18908 -19221
rect 18862 -19293 18908 -19255
rect 18862 -19327 18868 -19293
rect 18902 -19327 18908 -19293
rect 18862 -19365 18908 -19327
rect 18862 -19399 18868 -19365
rect 18902 -19399 18908 -19365
rect 18862 -19437 18908 -19399
rect 18862 -19471 18868 -19437
rect 18902 -19471 18908 -19437
rect 18862 -19509 18908 -19471
rect 18862 -19543 18868 -19509
rect 18902 -19543 18908 -19509
rect 18862 -19581 18908 -19543
rect 18862 -19615 18868 -19581
rect 18902 -19615 18908 -19581
rect 18862 -19653 18908 -19615
rect 17884 -19687 17896 -19664
rect 16096 -19756 16584 -19750
rect 16096 -19790 16143 -19756
rect 16177 -19790 16215 -19756
rect 16249 -19790 16287 -19756
rect 16321 -19790 16359 -19756
rect 16393 -19790 16431 -19756
rect 16465 -19790 16503 -19756
rect 16537 -19790 16584 -19756
rect 16096 -19796 16584 -19790
rect 17114 -19756 17602 -19750
rect 17114 -19790 17161 -19756
rect 17195 -19790 17233 -19756
rect 17267 -19790 17305 -19756
rect 17339 -19790 17377 -19756
rect 17411 -19790 17449 -19756
rect 17483 -19790 17521 -19756
rect 17555 -19790 17602 -19756
rect 17114 -19796 17602 -19790
rect 15796 -19842 15868 -19838
rect 15796 -19894 15806 -19842
rect 15858 -19894 15868 -19842
rect 15796 -19898 15868 -19894
rect 16150 -19842 16222 -19838
rect 16150 -19894 16160 -19842
rect 16212 -19894 16222 -19842
rect 16150 -19898 16222 -19894
rect 15792 -19954 15864 -19950
rect 15792 -20006 15802 -19954
rect 15854 -20006 15864 -19954
rect 15792 -20010 15864 -20006
rect 15302 -20052 15374 -20048
rect 15302 -20104 15312 -20052
rect 15364 -20104 15374 -20052
rect 15302 -20108 15374 -20104
rect 14060 -20280 14548 -20274
rect 14060 -20314 14107 -20280
rect 14141 -20314 14179 -20280
rect 14213 -20314 14251 -20280
rect 14285 -20314 14323 -20280
rect 14357 -20314 14395 -20280
rect 14429 -20314 14467 -20280
rect 14501 -20314 14548 -20280
rect 14060 -20320 14548 -20314
rect 15078 -20280 15566 -20274
rect 15078 -20314 15125 -20280
rect 15159 -20314 15197 -20280
rect 15231 -20314 15269 -20280
rect 15303 -20314 15341 -20280
rect 15375 -20314 15413 -20280
rect 15447 -20314 15485 -20280
rect 15519 -20314 15566 -20280
rect 15078 -20320 15566 -20314
rect 13766 -20402 13778 -20383
rect 12754 -20455 12800 -20417
rect 12754 -20489 12760 -20455
rect 12794 -20489 12800 -20455
rect 12754 -20527 12800 -20489
rect 12754 -20561 12760 -20527
rect 12794 -20561 12800 -20527
rect 12754 -20599 12800 -20561
rect 12754 -20633 12760 -20599
rect 12794 -20633 12800 -20599
rect 12754 -20671 12800 -20633
rect 12754 -20705 12760 -20671
rect 12794 -20705 12800 -20671
rect 12754 -20743 12800 -20705
rect 12754 -20777 12760 -20743
rect 12794 -20777 12800 -20743
rect 12754 -20815 12800 -20777
rect 12754 -20849 12760 -20815
rect 12794 -20849 12800 -20815
rect 12754 -20870 12800 -20849
rect 13772 -20417 13778 -20402
rect 13812 -20402 13826 -20383
rect 14790 -20383 14836 -20352
rect 13812 -20417 13818 -20402
rect 13772 -20455 13818 -20417
rect 13772 -20489 13778 -20455
rect 13812 -20489 13818 -20455
rect 13772 -20527 13818 -20489
rect 13772 -20561 13778 -20527
rect 13812 -20561 13818 -20527
rect 13772 -20599 13818 -20561
rect 13772 -20633 13778 -20599
rect 13812 -20633 13818 -20599
rect 13772 -20671 13818 -20633
rect 13772 -20705 13778 -20671
rect 13812 -20705 13818 -20671
rect 13772 -20743 13818 -20705
rect 13772 -20777 13778 -20743
rect 13812 -20777 13818 -20743
rect 13772 -20815 13818 -20777
rect 13772 -20849 13778 -20815
rect 13812 -20849 13818 -20815
rect 11736 -20921 11742 -20887
rect 11776 -20921 11782 -20887
rect 11736 -20952 11782 -20921
rect 12750 -20887 12810 -20870
rect 12750 -20921 12760 -20887
rect 12794 -20921 12810 -20887
rect 11006 -20990 11494 -20984
rect 11006 -21024 11053 -20990
rect 11087 -21024 11125 -20990
rect 11159 -21024 11197 -20990
rect 11231 -21024 11269 -20990
rect 11303 -21024 11341 -20990
rect 11375 -21024 11413 -20990
rect 11447 -21024 11494 -20990
rect 11006 -21030 11494 -21024
rect 12024 -20990 12512 -20984
rect 12024 -21024 12071 -20990
rect 12105 -21024 12143 -20990
rect 12177 -21024 12215 -20990
rect 12249 -21024 12287 -20990
rect 12321 -21024 12359 -20990
rect 12393 -21024 12431 -20990
rect 12465 -21024 12512 -20990
rect 12024 -21030 12512 -21024
rect 10538 -21120 10542 -21068
rect 10594 -21120 10598 -21068
rect 10186 -21186 10258 -21182
rect 10186 -21238 10196 -21186
rect 10248 -21238 10258 -21186
rect 10186 -21242 10258 -21238
rect 9684 -21402 9756 -21398
rect 9684 -21454 9694 -21402
rect 9746 -21454 9756 -21402
rect 9684 -21458 9756 -21454
rect 8970 -21512 9458 -21506
rect 8970 -21546 9017 -21512
rect 9051 -21546 9089 -21512
rect 9123 -21546 9161 -21512
rect 9195 -21546 9233 -21512
rect 9267 -21546 9305 -21512
rect 9339 -21546 9377 -21512
rect 9411 -21546 9458 -21512
rect 8970 -21552 9458 -21546
rect 7704 -21649 7710 -21636
rect 7664 -21687 7710 -21649
rect 8670 -21649 8688 -21615
rect 8722 -21649 8730 -21615
rect 9690 -21615 9750 -21458
rect 10192 -21506 10252 -21242
rect 10538 -21278 10598 -21120
rect 10702 -21068 10774 -21064
rect 10702 -21120 10712 -21068
rect 10764 -21120 10774 -21068
rect 10702 -21124 10774 -21120
rect 10708 -21276 10780 -21272
rect 10532 -21282 10604 -21278
rect 10532 -21334 10542 -21282
rect 10594 -21334 10604 -21282
rect 10708 -21328 10718 -21276
rect 10770 -21328 10780 -21276
rect 10708 -21332 10780 -21328
rect 10532 -21338 10604 -21334
rect 9988 -21512 10252 -21506
rect 10264 -21512 10476 -21506
rect 9988 -21546 10035 -21512
rect 10069 -21546 10107 -21512
rect 10141 -21546 10179 -21512
rect 10213 -21546 10251 -21512
rect 10285 -21546 10323 -21512
rect 10357 -21546 10395 -21512
rect 10429 -21546 10476 -21512
rect 9988 -21552 10476 -21546
rect 9690 -21636 9706 -21615
rect 8670 -21656 8730 -21649
rect 9700 -21649 9706 -21636
rect 9740 -21636 9750 -21615
rect 10714 -21615 10774 -21332
rect 11230 -21334 11290 -21030
rect 12244 -21170 12304 -21030
rect 12750 -21064 12810 -20921
rect 13772 -20887 13818 -20849
rect 14790 -20417 14796 -20383
rect 14830 -20417 14836 -20383
rect 15798 -20383 15858 -20010
rect 16156 -20160 16216 -19898
rect 16346 -20048 16406 -19796
rect 17322 -20048 17382 -19796
rect 16340 -20052 16412 -20048
rect 16340 -20104 16350 -20052
rect 16402 -20104 16412 -20052
rect 16340 -20108 16412 -20104
rect 17316 -20052 17388 -20048
rect 17316 -20104 17326 -20052
rect 17378 -20104 17388 -20052
rect 17316 -20108 17388 -20104
rect 17836 -20160 17896 -19687
rect 18862 -19687 18868 -19653
rect 18902 -19687 18908 -19653
rect 19880 -19221 19926 -19183
rect 19880 -19255 19886 -19221
rect 19920 -19255 19926 -19221
rect 19880 -19293 19926 -19255
rect 19880 -19327 19886 -19293
rect 19920 -19327 19926 -19293
rect 19880 -19365 19926 -19327
rect 19880 -19399 19886 -19365
rect 19920 -19399 19926 -19365
rect 19880 -19437 19926 -19399
rect 19880 -19471 19886 -19437
rect 19920 -19471 19926 -19437
rect 19880 -19509 19926 -19471
rect 19880 -19543 19886 -19509
rect 19920 -19543 19926 -19509
rect 19880 -19581 19926 -19543
rect 19880 -19615 19886 -19581
rect 19920 -19615 19926 -19581
rect 19880 -19653 19926 -19615
rect 19880 -19662 19886 -19653
rect 18862 -19718 18908 -19687
rect 19874 -19687 19886 -19662
rect 19920 -19662 19926 -19653
rect 20898 -19183 20904 -19182
rect 20938 -19182 20950 -19149
rect 21912 -19149 21972 -18996
rect 22204 -19046 22692 -19040
rect 22204 -19080 22251 -19046
rect 22285 -19080 22323 -19046
rect 22357 -19080 22395 -19046
rect 22429 -19080 22467 -19046
rect 22501 -19080 22539 -19046
rect 22573 -19080 22611 -19046
rect 22645 -19080 22692 -19046
rect 22204 -19086 22692 -19080
rect 21912 -19164 21922 -19149
rect 20938 -19183 20944 -19182
rect 20898 -19221 20944 -19183
rect 20898 -19255 20904 -19221
rect 20938 -19255 20944 -19221
rect 20898 -19293 20944 -19255
rect 20898 -19327 20904 -19293
rect 20938 -19327 20944 -19293
rect 20898 -19365 20944 -19327
rect 20898 -19399 20904 -19365
rect 20938 -19399 20944 -19365
rect 20898 -19437 20944 -19399
rect 20898 -19471 20904 -19437
rect 20938 -19471 20944 -19437
rect 20898 -19509 20944 -19471
rect 20898 -19543 20904 -19509
rect 20938 -19543 20944 -19509
rect 20898 -19581 20944 -19543
rect 20898 -19615 20904 -19581
rect 20938 -19615 20944 -19581
rect 20898 -19653 20944 -19615
rect 20898 -19656 20904 -19653
rect 19920 -19687 19934 -19662
rect 18132 -19756 18620 -19750
rect 18132 -19790 18179 -19756
rect 18213 -19790 18251 -19756
rect 18285 -19790 18323 -19756
rect 18357 -19790 18395 -19756
rect 18429 -19790 18467 -19756
rect 18501 -19790 18539 -19756
rect 18573 -19790 18620 -19756
rect 18132 -19796 18620 -19790
rect 19150 -19756 19638 -19750
rect 19150 -19790 19197 -19756
rect 19231 -19790 19269 -19756
rect 19303 -19790 19341 -19756
rect 19375 -19790 19413 -19756
rect 19447 -19790 19485 -19756
rect 19519 -19790 19557 -19756
rect 19591 -19790 19638 -19756
rect 19150 -19796 19638 -19790
rect 18338 -20048 18398 -19796
rect 19874 -19838 19934 -19687
rect 20892 -19687 20904 -19656
rect 20938 -19656 20944 -19653
rect 21916 -19183 21922 -19164
rect 21956 -19164 21972 -19149
rect 22934 -19149 22980 -19118
rect 21956 -19183 21962 -19164
rect 21916 -19221 21962 -19183
rect 21916 -19255 21922 -19221
rect 21956 -19255 21962 -19221
rect 21916 -19293 21962 -19255
rect 21916 -19327 21922 -19293
rect 21956 -19327 21962 -19293
rect 21916 -19365 21962 -19327
rect 21916 -19399 21922 -19365
rect 21956 -19399 21962 -19365
rect 21916 -19437 21962 -19399
rect 21916 -19471 21922 -19437
rect 21956 -19471 21962 -19437
rect 21916 -19509 21962 -19471
rect 21916 -19543 21922 -19509
rect 21956 -19543 21962 -19509
rect 21916 -19581 21962 -19543
rect 21916 -19615 21922 -19581
rect 21956 -19615 21962 -19581
rect 21916 -19653 21962 -19615
rect 20938 -19687 20952 -19656
rect 21916 -19662 21922 -19653
rect 20168 -19756 20656 -19750
rect 20168 -19790 20215 -19756
rect 20249 -19790 20287 -19756
rect 20321 -19790 20359 -19756
rect 20393 -19790 20431 -19756
rect 20465 -19790 20503 -19756
rect 20537 -19790 20575 -19756
rect 20609 -19790 20656 -19756
rect 20168 -19796 20656 -19790
rect 19868 -19842 19940 -19838
rect 19868 -19894 19878 -19842
rect 19930 -19894 19940 -19842
rect 19868 -19898 19940 -19894
rect 18332 -20052 18404 -20048
rect 18332 -20104 18342 -20052
rect 18394 -20104 18404 -20052
rect 18332 -20108 18404 -20104
rect 20358 -20052 20430 -20048
rect 20358 -20104 20368 -20052
rect 20420 -20104 20430 -20052
rect 20358 -20108 20430 -20104
rect 16156 -20212 16160 -20160
rect 16212 -20212 16216 -20160
rect 16156 -20222 16216 -20212
rect 17830 -20164 17902 -20160
rect 17830 -20216 17840 -20164
rect 17892 -20216 17902 -20164
rect 17830 -20220 17902 -20216
rect 19866 -20164 19938 -20160
rect 19866 -20216 19876 -20164
rect 19928 -20216 19938 -20164
rect 19866 -20220 19938 -20216
rect 16096 -20280 16584 -20274
rect 16096 -20314 16143 -20280
rect 16177 -20314 16215 -20280
rect 16249 -20314 16287 -20280
rect 16321 -20314 16359 -20280
rect 16393 -20314 16431 -20280
rect 16465 -20314 16503 -20280
rect 16537 -20314 16584 -20280
rect 16096 -20320 16584 -20314
rect 17114 -20280 17602 -20274
rect 17114 -20314 17161 -20280
rect 17195 -20314 17233 -20280
rect 17267 -20314 17305 -20280
rect 17339 -20314 17377 -20280
rect 17411 -20314 17449 -20280
rect 17483 -20314 17521 -20280
rect 17555 -20314 17602 -20280
rect 17114 -20320 17602 -20314
rect 15798 -20406 15814 -20383
rect 14790 -20455 14836 -20417
rect 14790 -20489 14796 -20455
rect 14830 -20489 14836 -20455
rect 14790 -20527 14836 -20489
rect 14790 -20561 14796 -20527
rect 14830 -20561 14836 -20527
rect 14790 -20599 14836 -20561
rect 14790 -20633 14796 -20599
rect 14830 -20633 14836 -20599
rect 14790 -20671 14836 -20633
rect 14790 -20705 14796 -20671
rect 14830 -20705 14836 -20671
rect 14790 -20743 14836 -20705
rect 14790 -20777 14796 -20743
rect 14830 -20777 14836 -20743
rect 14790 -20815 14836 -20777
rect 14790 -20849 14796 -20815
rect 14830 -20849 14836 -20815
rect 14790 -20870 14836 -20849
rect 15808 -20417 15814 -20406
rect 15848 -20406 15858 -20383
rect 16826 -20383 16872 -20352
rect 15848 -20417 15854 -20406
rect 15808 -20455 15854 -20417
rect 15808 -20489 15814 -20455
rect 15848 -20489 15854 -20455
rect 15808 -20527 15854 -20489
rect 15808 -20561 15814 -20527
rect 15848 -20561 15854 -20527
rect 15808 -20599 15854 -20561
rect 15808 -20633 15814 -20599
rect 15848 -20633 15854 -20599
rect 15808 -20671 15854 -20633
rect 15808 -20705 15814 -20671
rect 15848 -20705 15854 -20671
rect 15808 -20743 15854 -20705
rect 15808 -20777 15814 -20743
rect 15848 -20777 15854 -20743
rect 15808 -20815 15854 -20777
rect 15808 -20849 15814 -20815
rect 15848 -20849 15854 -20815
rect 13772 -20921 13778 -20887
rect 13812 -20921 13818 -20887
rect 13772 -20952 13818 -20921
rect 14782 -20887 14842 -20870
rect 14782 -20921 14796 -20887
rect 14830 -20921 14842 -20887
rect 13042 -20990 13530 -20984
rect 13042 -21024 13089 -20990
rect 13123 -21024 13161 -20990
rect 13195 -21024 13233 -20990
rect 13267 -21024 13305 -20990
rect 13339 -21024 13377 -20990
rect 13411 -21024 13449 -20990
rect 13483 -21024 13530 -20990
rect 13042 -21030 13530 -21024
rect 14060 -20990 14548 -20984
rect 14060 -21024 14107 -20990
rect 14141 -21024 14179 -20990
rect 14213 -21024 14251 -20990
rect 14285 -21024 14323 -20990
rect 14357 -21024 14395 -20990
rect 14429 -21024 14467 -20990
rect 14501 -21024 14548 -20990
rect 14060 -21030 14548 -21024
rect 12744 -21068 12816 -21064
rect 12744 -21120 12754 -21068
rect 12806 -21120 12816 -21068
rect 12744 -21124 12816 -21120
rect 13266 -21170 13326 -21030
rect 14280 -21170 14340 -21030
rect 14782 -21064 14842 -20921
rect 15808 -20887 15854 -20849
rect 15808 -20921 15814 -20887
rect 15848 -20921 15854 -20887
rect 16826 -20417 16832 -20383
rect 16866 -20417 16872 -20383
rect 17836 -20383 17896 -20220
rect 18132 -20280 18620 -20274
rect 18132 -20314 18179 -20280
rect 18213 -20314 18251 -20280
rect 18285 -20314 18323 -20280
rect 18357 -20314 18395 -20280
rect 18429 -20314 18467 -20280
rect 18501 -20314 18539 -20280
rect 18573 -20314 18620 -20280
rect 18132 -20320 18620 -20314
rect 19150 -20280 19638 -20274
rect 19150 -20314 19197 -20280
rect 19231 -20314 19269 -20280
rect 19303 -20314 19341 -20280
rect 19375 -20314 19413 -20280
rect 19447 -20314 19485 -20280
rect 19519 -20314 19557 -20280
rect 19591 -20314 19638 -20280
rect 19150 -20320 19638 -20314
rect 17836 -20402 17850 -20383
rect 16826 -20455 16872 -20417
rect 16826 -20489 16832 -20455
rect 16866 -20489 16872 -20455
rect 16826 -20527 16872 -20489
rect 16826 -20561 16832 -20527
rect 16866 -20561 16872 -20527
rect 16826 -20599 16872 -20561
rect 16826 -20633 16832 -20599
rect 16866 -20633 16872 -20599
rect 16826 -20671 16872 -20633
rect 16826 -20705 16832 -20671
rect 16866 -20705 16872 -20671
rect 16826 -20743 16872 -20705
rect 16826 -20777 16832 -20743
rect 16866 -20777 16872 -20743
rect 16826 -20815 16872 -20777
rect 16826 -20849 16832 -20815
rect 16866 -20849 16872 -20815
rect 16826 -20887 16872 -20849
rect 16826 -20904 16832 -20887
rect 15808 -20952 15854 -20921
rect 16822 -20921 16832 -20904
rect 16866 -20904 16872 -20887
rect 17844 -20417 17850 -20402
rect 17884 -20402 17896 -20383
rect 18862 -20383 18908 -20352
rect 17884 -20417 17890 -20402
rect 17844 -20455 17890 -20417
rect 17844 -20489 17850 -20455
rect 17884 -20489 17890 -20455
rect 17844 -20527 17890 -20489
rect 17844 -20561 17850 -20527
rect 17884 -20561 17890 -20527
rect 17844 -20599 17890 -20561
rect 17844 -20633 17850 -20599
rect 17884 -20633 17890 -20599
rect 17844 -20671 17890 -20633
rect 17844 -20705 17850 -20671
rect 17884 -20705 17890 -20671
rect 17844 -20743 17890 -20705
rect 17844 -20777 17850 -20743
rect 17884 -20777 17890 -20743
rect 17844 -20815 17890 -20777
rect 17844 -20849 17850 -20815
rect 17884 -20849 17890 -20815
rect 17844 -20887 17890 -20849
rect 17844 -20888 17850 -20887
rect 16866 -20921 16882 -20904
rect 15078 -20990 15566 -20984
rect 15078 -21024 15125 -20990
rect 15159 -21024 15197 -20990
rect 15231 -21024 15269 -20990
rect 15303 -21024 15341 -20990
rect 15375 -21024 15413 -20990
rect 15447 -21024 15485 -20990
rect 15519 -21024 15566 -20990
rect 15078 -21030 15566 -21024
rect 16096 -20990 16584 -20984
rect 16096 -21024 16143 -20990
rect 16177 -21024 16215 -20990
rect 16249 -21024 16287 -20990
rect 16321 -21024 16359 -20990
rect 16393 -21024 16431 -20990
rect 16465 -21024 16503 -20990
rect 16537 -21024 16584 -20990
rect 16096 -21030 16584 -21024
rect 14776 -21068 14848 -21064
rect 14776 -21120 14786 -21068
rect 14838 -21120 14848 -21068
rect 14776 -21124 14848 -21120
rect 15282 -21070 15342 -21030
rect 16308 -21070 16368 -21030
rect 16822 -21064 16882 -20921
rect 17840 -20921 17850 -20888
rect 17884 -20888 17890 -20887
rect 18862 -20417 18868 -20383
rect 18902 -20417 18908 -20383
rect 18862 -20455 18908 -20417
rect 19872 -20383 19932 -20220
rect 20364 -20274 20424 -20108
rect 20168 -20280 20656 -20274
rect 20168 -20314 20215 -20280
rect 20249 -20314 20287 -20280
rect 20321 -20314 20359 -20280
rect 20393 -20314 20431 -20280
rect 20465 -20314 20503 -20280
rect 20537 -20314 20575 -20280
rect 20609 -20314 20656 -20280
rect 20168 -20320 20656 -20314
rect 19872 -20417 19886 -20383
rect 19920 -20417 19932 -20383
rect 20892 -20383 20952 -19687
rect 21908 -19687 21922 -19662
rect 21956 -19662 21962 -19653
rect 22934 -19183 22940 -19149
rect 22974 -19183 22980 -19149
rect 22934 -19221 22980 -19183
rect 22934 -19255 22940 -19221
rect 22974 -19255 22980 -19221
rect 22934 -19293 22980 -19255
rect 22934 -19327 22940 -19293
rect 22974 -19327 22980 -19293
rect 22934 -19365 22980 -19327
rect 22934 -19399 22940 -19365
rect 22974 -19399 22980 -19365
rect 22934 -19437 22980 -19399
rect 22934 -19471 22940 -19437
rect 22974 -19471 22980 -19437
rect 22934 -19509 22980 -19471
rect 22934 -19543 22940 -19509
rect 22974 -19543 22980 -19509
rect 22934 -19581 22980 -19543
rect 22934 -19615 22940 -19581
rect 22974 -19615 22980 -19581
rect 22934 -19653 22980 -19615
rect 21956 -19687 21968 -19662
rect 22934 -19676 22940 -19653
rect 21186 -19756 21674 -19750
rect 21186 -19790 21233 -19756
rect 21267 -19790 21305 -19756
rect 21339 -19790 21377 -19756
rect 21411 -19790 21449 -19756
rect 21483 -19790 21521 -19756
rect 21555 -19790 21593 -19756
rect 21627 -19790 21674 -19756
rect 21186 -19796 21674 -19790
rect 21394 -20048 21454 -19796
rect 21908 -19888 21968 -19687
rect 22924 -19687 22940 -19676
rect 22974 -19676 22980 -19653
rect 22974 -19687 22984 -19676
rect 22204 -19756 22692 -19750
rect 22204 -19790 22251 -19756
rect 22285 -19790 22323 -19756
rect 22357 -19790 22395 -19756
rect 22429 -19790 22467 -19756
rect 22501 -19790 22539 -19756
rect 22573 -19790 22611 -19756
rect 22645 -19790 22692 -19756
rect 22204 -19796 22692 -19790
rect 22414 -19888 22474 -19796
rect 22924 -19888 22984 -19687
rect 21908 -19948 22984 -19888
rect 21388 -20052 21460 -20048
rect 21388 -20104 21398 -20052
rect 21450 -20104 21460 -20052
rect 21388 -20108 21460 -20104
rect 21908 -20160 21968 -19948
rect 21902 -20164 21974 -20160
rect 21902 -20216 21912 -20164
rect 21964 -20216 21974 -20164
rect 21902 -20220 21974 -20216
rect 21186 -20280 21674 -20274
rect 21186 -20314 21233 -20280
rect 21267 -20314 21305 -20280
rect 21339 -20314 21377 -20280
rect 21411 -20314 21449 -20280
rect 21483 -20314 21521 -20280
rect 21555 -20314 21593 -20280
rect 21627 -20314 21674 -20280
rect 21186 -20320 21674 -20314
rect 22204 -20280 22692 -20274
rect 22204 -20314 22251 -20280
rect 22285 -20314 22323 -20280
rect 22357 -20314 22395 -20280
rect 22429 -20314 22467 -20280
rect 22501 -20314 22539 -20280
rect 22573 -20314 22611 -20280
rect 22645 -20314 22692 -20280
rect 22204 -20320 22692 -20314
rect 20892 -20406 20904 -20383
rect 19872 -20422 19932 -20417
rect 20898 -20417 20904 -20406
rect 20938 -20406 20952 -20383
rect 21916 -20383 21962 -20352
rect 20938 -20417 20944 -20406
rect 18862 -20489 18868 -20455
rect 18902 -20489 18908 -20455
rect 18862 -20527 18908 -20489
rect 18862 -20561 18868 -20527
rect 18902 -20561 18908 -20527
rect 18862 -20599 18908 -20561
rect 18862 -20633 18868 -20599
rect 18902 -20633 18908 -20599
rect 18862 -20671 18908 -20633
rect 18862 -20705 18868 -20671
rect 18902 -20705 18908 -20671
rect 18862 -20743 18908 -20705
rect 18862 -20777 18868 -20743
rect 18902 -20777 18908 -20743
rect 18862 -20815 18908 -20777
rect 18862 -20849 18868 -20815
rect 18902 -20849 18908 -20815
rect 18862 -20887 18908 -20849
rect 17884 -20921 17900 -20888
rect 18862 -20896 18868 -20887
rect 17114 -20990 17602 -20984
rect 17114 -21024 17161 -20990
rect 17195 -21024 17233 -20990
rect 17267 -21024 17305 -20990
rect 17339 -21024 17377 -20990
rect 17411 -21024 17449 -20990
rect 17483 -21024 17521 -20990
rect 17555 -21024 17602 -20990
rect 17114 -21030 17602 -21024
rect 15282 -21130 16368 -21070
rect 16816 -21068 16888 -21064
rect 16816 -21120 16826 -21068
rect 16878 -21120 16888 -21068
rect 16816 -21124 16888 -21120
rect 15282 -21170 15342 -21130
rect 12244 -21230 15342 -21170
rect 15794 -21166 15866 -21162
rect 15794 -21218 15804 -21166
rect 15856 -21218 15866 -21166
rect 15794 -21222 15866 -21218
rect 12244 -21334 12304 -21230
rect 12736 -21276 12808 -21272
rect 12736 -21328 12746 -21276
rect 12798 -21328 12808 -21276
rect 12736 -21332 12808 -21328
rect 11230 -21394 12304 -21334
rect 11230 -21506 11290 -21394
rect 12244 -21506 12304 -21394
rect 11006 -21512 11494 -21506
rect 11006 -21546 11053 -21512
rect 11087 -21546 11125 -21512
rect 11159 -21546 11197 -21512
rect 11231 -21546 11269 -21512
rect 11303 -21546 11341 -21512
rect 11375 -21546 11413 -21512
rect 11447 -21546 11494 -21512
rect 11006 -21552 11494 -21546
rect 12024 -21512 12512 -21506
rect 12024 -21546 12071 -21512
rect 12105 -21546 12143 -21512
rect 12177 -21546 12215 -21512
rect 12249 -21546 12287 -21512
rect 12321 -21546 12359 -21512
rect 12393 -21546 12431 -21512
rect 12465 -21546 12512 -21512
rect 12024 -21552 12512 -21546
rect 9740 -21649 9746 -21636
rect 10714 -21640 10724 -21615
rect 7664 -21721 7670 -21687
rect 7704 -21721 7710 -21687
rect 7664 -21759 7710 -21721
rect 7664 -21793 7670 -21759
rect 7704 -21793 7710 -21759
rect 7664 -21831 7710 -21793
rect 7664 -21865 7670 -21831
rect 7704 -21865 7710 -21831
rect 7664 -21903 7710 -21865
rect 7664 -21937 7670 -21903
rect 7704 -21937 7710 -21903
rect 7664 -21975 7710 -21937
rect 7664 -22009 7670 -21975
rect 7704 -22009 7710 -21975
rect 7664 -22047 7710 -22009
rect 7664 -22081 7670 -22047
rect 7704 -22081 7710 -22047
rect 7664 -22118 7710 -22081
rect 8682 -21687 8728 -21656
rect 8682 -21721 8688 -21687
rect 8722 -21721 8728 -21687
rect 8682 -21759 8728 -21721
rect 8682 -21793 8688 -21759
rect 8722 -21793 8728 -21759
rect 8682 -21831 8728 -21793
rect 8682 -21865 8688 -21831
rect 8722 -21865 8728 -21831
rect 8682 -21903 8728 -21865
rect 8682 -21937 8688 -21903
rect 8722 -21937 8728 -21903
rect 8682 -21975 8728 -21937
rect 8682 -22009 8688 -21975
rect 8722 -22009 8728 -21975
rect 8682 -22047 8728 -22009
rect 8682 -22081 8688 -22047
rect 8722 -22081 8728 -22047
rect 5668 -22153 5680 -22130
rect 2862 -22222 3350 -22216
rect 2862 -22256 2909 -22222
rect 2943 -22256 2981 -22222
rect 3015 -22256 3053 -22222
rect 3087 -22256 3125 -22222
rect 3159 -22256 3197 -22222
rect 3231 -22256 3269 -22222
rect 3303 -22256 3350 -22222
rect 2862 -22262 3350 -22256
rect 3880 -22222 4368 -22216
rect 3880 -22256 3927 -22222
rect 3961 -22256 3999 -22222
rect 4033 -22256 4071 -22222
rect 4105 -22256 4143 -22222
rect 4177 -22256 4215 -22222
rect 4249 -22256 4287 -22222
rect 4321 -22256 4368 -22222
rect 3880 -22262 4368 -22256
rect 4898 -22222 5386 -22216
rect 4898 -22256 4945 -22222
rect 4979 -22256 5017 -22222
rect 5051 -22256 5089 -22222
rect 5123 -22256 5161 -22222
rect 5195 -22256 5233 -22222
rect 5267 -22256 5305 -22222
rect 5339 -22256 5386 -22222
rect 4898 -22262 5386 -22256
rect 2330 -22318 2402 -22314
rect 2330 -22370 2340 -22318
rect 2392 -22370 2402 -22318
rect 2330 -22374 2402 -22370
rect 5620 -22440 5680 -22153
rect 6646 -22153 6652 -22119
rect 6686 -22153 6692 -22119
rect 6646 -22184 6692 -22153
rect 7658 -22119 7718 -22118
rect 7658 -22153 7670 -22119
rect 7704 -22153 7718 -22119
rect 5916 -22222 6404 -22216
rect 5916 -22256 5963 -22222
rect 5997 -22256 6035 -22222
rect 6069 -22256 6107 -22222
rect 6141 -22256 6179 -22222
rect 6213 -22256 6251 -22222
rect 6285 -22256 6323 -22222
rect 6357 -22256 6404 -22222
rect 5916 -22262 6256 -22256
rect 6316 -22262 6404 -22256
rect 6934 -22222 7422 -22216
rect 6934 -22256 6981 -22222
rect 7015 -22256 7053 -22222
rect 7087 -22256 7125 -22222
rect 7159 -22256 7197 -22222
rect 7231 -22256 7269 -22222
rect 7303 -22256 7341 -22222
rect 7375 -22256 7422 -22222
rect 6934 -22262 7422 -22256
rect 6140 -22428 6200 -22262
rect 6134 -22432 6206 -22428
rect 2224 -22444 2296 -22440
rect 2224 -22496 2234 -22444
rect 2286 -22496 2296 -22444
rect 2224 -22500 2296 -22496
rect 5614 -22444 5686 -22440
rect 5614 -22496 5624 -22444
rect 5676 -22496 5686 -22444
rect 6134 -22484 6144 -22432
rect 6196 -22484 6206 -22432
rect 6134 -22488 6206 -22484
rect 5614 -22500 5686 -22496
rect 4596 -22554 4668 -22550
rect 4596 -22606 4606 -22554
rect 4658 -22606 4668 -22554
rect 4596 -22610 4668 -22606
rect 6632 -22554 6704 -22550
rect 6632 -22606 6642 -22554
rect 6694 -22606 6704 -22554
rect 6632 -22610 6704 -22606
rect 2862 -22746 3350 -22740
rect 2862 -22780 2909 -22746
rect 2943 -22780 2981 -22746
rect 3015 -22780 3053 -22746
rect 3087 -22780 3125 -22746
rect 3159 -22780 3197 -22746
rect 3231 -22780 3269 -22746
rect 3303 -22780 3350 -22746
rect 2862 -22786 3350 -22780
rect 3880 -22746 4368 -22740
rect 3880 -22780 3927 -22746
rect 3961 -22780 3999 -22746
rect 4033 -22780 4071 -22746
rect 4105 -22780 4143 -22746
rect 4177 -22780 4215 -22746
rect 4249 -22780 4287 -22746
rect 4321 -22780 4368 -22746
rect 3880 -22786 4368 -22780
rect 2574 -22849 2620 -22818
rect 2574 -22883 2580 -22849
rect 2614 -22883 2620 -22849
rect 2574 -22921 2620 -22883
rect 2574 -22955 2580 -22921
rect 2614 -22955 2620 -22921
rect 2574 -22993 2620 -22955
rect 2574 -23027 2580 -22993
rect 2614 -23027 2620 -22993
rect 2574 -23065 2620 -23027
rect 2574 -23099 2580 -23065
rect 2614 -23099 2620 -23065
rect 2574 -23137 2620 -23099
rect 2574 -23171 2580 -23137
rect 2614 -23171 2620 -23137
rect 2574 -23209 2620 -23171
rect 2574 -23243 2580 -23209
rect 2614 -23243 2620 -23209
rect 2574 -23281 2620 -23243
rect 2574 -23315 2580 -23281
rect 2614 -23315 2620 -23281
rect 2574 -23353 2620 -23315
rect 3592 -22849 3638 -22818
rect 3592 -22883 3598 -22849
rect 3632 -22883 3638 -22849
rect 3592 -22921 3638 -22883
rect 4602 -22849 4662 -22610
rect 6250 -22648 6322 -22644
rect 6250 -22700 6260 -22648
rect 6312 -22700 6322 -22648
rect 6250 -22704 6322 -22700
rect 6256 -22740 6316 -22704
rect 4898 -22746 5386 -22740
rect 4898 -22780 4945 -22746
rect 4979 -22780 5017 -22746
rect 5051 -22780 5089 -22746
rect 5123 -22780 5161 -22746
rect 5195 -22780 5233 -22746
rect 5267 -22780 5305 -22746
rect 5339 -22780 5386 -22746
rect 4898 -22786 5386 -22780
rect 5916 -22746 6404 -22740
rect 5916 -22780 5963 -22746
rect 5997 -22780 6035 -22746
rect 6069 -22780 6107 -22746
rect 6141 -22780 6179 -22746
rect 6213 -22780 6251 -22746
rect 6285 -22780 6323 -22746
rect 6357 -22780 6404 -22746
rect 5916 -22786 6404 -22780
rect 4602 -22883 4616 -22849
rect 4650 -22883 4662 -22849
rect 4602 -22890 4662 -22883
rect 5628 -22849 5674 -22818
rect 5628 -22883 5634 -22849
rect 5668 -22883 5674 -22849
rect 6638 -22849 6698 -22610
rect 7140 -22644 7200 -22262
rect 7658 -22550 7718 -22153
rect 8682 -22119 8728 -22081
rect 9700 -21687 9746 -21649
rect 9700 -21721 9706 -21687
rect 9740 -21721 9746 -21687
rect 9700 -21759 9746 -21721
rect 9700 -21793 9706 -21759
rect 9740 -21793 9746 -21759
rect 9700 -21831 9746 -21793
rect 9700 -21865 9706 -21831
rect 9740 -21865 9746 -21831
rect 9700 -21903 9746 -21865
rect 9700 -21937 9706 -21903
rect 9740 -21937 9746 -21903
rect 9700 -21975 9746 -21937
rect 9700 -22009 9706 -21975
rect 9740 -22009 9746 -21975
rect 9700 -22047 9746 -22009
rect 9700 -22081 9706 -22047
rect 9740 -22081 9746 -22047
rect 9700 -22106 9746 -22081
rect 10718 -21649 10724 -21640
rect 10758 -21640 10774 -21615
rect 11736 -21615 11782 -21584
rect 10758 -21649 10764 -21640
rect 10718 -21687 10764 -21649
rect 10718 -21721 10724 -21687
rect 10758 -21721 10764 -21687
rect 10718 -21759 10764 -21721
rect 10718 -21793 10724 -21759
rect 10758 -21793 10764 -21759
rect 10718 -21831 10764 -21793
rect 10718 -21865 10724 -21831
rect 10758 -21865 10764 -21831
rect 10718 -21903 10764 -21865
rect 10718 -21937 10724 -21903
rect 10758 -21937 10764 -21903
rect 10718 -21975 10764 -21937
rect 10718 -22009 10724 -21975
rect 10758 -22009 10764 -21975
rect 10718 -22047 10764 -22009
rect 10718 -22081 10724 -22047
rect 10758 -22081 10764 -22047
rect 8682 -22153 8688 -22119
rect 8722 -22153 8728 -22119
rect 8682 -22184 8728 -22153
rect 9694 -22119 9754 -22106
rect 9694 -22153 9706 -22119
rect 9740 -22153 9754 -22119
rect 7952 -22222 8440 -22216
rect 7952 -22256 7999 -22222
rect 8033 -22256 8071 -22222
rect 8105 -22256 8143 -22222
rect 8177 -22256 8215 -22222
rect 8249 -22256 8287 -22222
rect 8321 -22256 8359 -22222
rect 8393 -22256 8440 -22222
rect 7952 -22262 8440 -22256
rect 8970 -22222 9458 -22216
rect 8970 -22256 9017 -22222
rect 9051 -22256 9089 -22222
rect 9123 -22256 9161 -22222
rect 9195 -22256 9233 -22222
rect 9267 -22256 9305 -22222
rect 9339 -22256 9377 -22222
rect 9411 -22256 9458 -22222
rect 8970 -22262 9458 -22256
rect 7652 -22554 7724 -22550
rect 7652 -22606 7662 -22554
rect 7714 -22606 7724 -22554
rect 7652 -22610 7724 -22606
rect 8162 -22644 8222 -22262
rect 9694 -22550 9754 -22153
rect 10718 -22119 10764 -22081
rect 10718 -22153 10724 -22119
rect 10758 -22153 10764 -22119
rect 11736 -21649 11742 -21615
rect 11776 -21649 11782 -21615
rect 12742 -21615 12802 -21332
rect 13266 -21506 13326 -21230
rect 14280 -21506 14340 -21230
rect 14780 -21276 14852 -21272
rect 14780 -21328 14790 -21276
rect 14842 -21328 14852 -21276
rect 14780 -21332 14852 -21328
rect 13042 -21512 13530 -21506
rect 13042 -21546 13089 -21512
rect 13123 -21546 13161 -21512
rect 13195 -21546 13233 -21512
rect 13267 -21546 13305 -21512
rect 13339 -21546 13377 -21512
rect 13411 -21546 13449 -21512
rect 13483 -21546 13530 -21512
rect 13042 -21552 13530 -21546
rect 14060 -21512 14548 -21506
rect 14060 -21546 14107 -21512
rect 14141 -21546 14179 -21512
rect 14213 -21546 14251 -21512
rect 14285 -21546 14323 -21512
rect 14357 -21546 14395 -21512
rect 14429 -21546 14467 -21512
rect 14501 -21546 14548 -21512
rect 14060 -21552 14548 -21546
rect 12742 -21640 12760 -21615
rect 11736 -21687 11782 -21649
rect 11736 -21721 11742 -21687
rect 11776 -21721 11782 -21687
rect 11736 -21759 11782 -21721
rect 11736 -21793 11742 -21759
rect 11776 -21793 11782 -21759
rect 11736 -21831 11782 -21793
rect 11736 -21865 11742 -21831
rect 11776 -21865 11782 -21831
rect 11736 -21903 11782 -21865
rect 11736 -21937 11742 -21903
rect 11776 -21937 11782 -21903
rect 11736 -21975 11782 -21937
rect 11736 -22009 11742 -21975
rect 11776 -22009 11782 -21975
rect 11736 -22047 11782 -22009
rect 11736 -22081 11742 -22047
rect 11776 -22081 11782 -22047
rect 11736 -22119 11782 -22081
rect 11736 -22120 11742 -22119
rect 10718 -22184 10764 -22153
rect 11724 -22153 11742 -22120
rect 11776 -22120 11782 -22119
rect 12754 -21649 12760 -21640
rect 12794 -21640 12802 -21615
rect 13772 -21615 13818 -21584
rect 12794 -21649 12800 -21640
rect 12754 -21687 12800 -21649
rect 12754 -21721 12760 -21687
rect 12794 -21721 12800 -21687
rect 12754 -21759 12800 -21721
rect 12754 -21793 12760 -21759
rect 12794 -21793 12800 -21759
rect 12754 -21831 12800 -21793
rect 12754 -21865 12760 -21831
rect 12794 -21865 12800 -21831
rect 12754 -21903 12800 -21865
rect 12754 -21937 12760 -21903
rect 12794 -21937 12800 -21903
rect 12754 -21975 12800 -21937
rect 12754 -22009 12760 -21975
rect 12794 -22009 12800 -21975
rect 12754 -22047 12800 -22009
rect 12754 -22081 12760 -22047
rect 12794 -22081 12800 -22047
rect 12754 -22119 12800 -22081
rect 11776 -22153 11784 -22120
rect 9988 -22222 10476 -22216
rect 9988 -22256 10035 -22222
rect 10069 -22256 10107 -22222
rect 10141 -22256 10179 -22222
rect 10213 -22256 10251 -22222
rect 10285 -22256 10323 -22222
rect 10357 -22256 10395 -22222
rect 10429 -22256 10476 -22222
rect 9988 -22262 10476 -22256
rect 11006 -22222 11494 -22216
rect 11006 -22256 11053 -22222
rect 11087 -22256 11125 -22222
rect 11159 -22256 11197 -22222
rect 11231 -22256 11269 -22222
rect 11303 -22256 11341 -22222
rect 11375 -22256 11413 -22222
rect 11447 -22256 11494 -22222
rect 11006 -22262 11494 -22256
rect 8668 -22554 8740 -22550
rect 8668 -22606 8678 -22554
rect 8730 -22606 8740 -22554
rect 8668 -22610 8740 -22606
rect 9688 -22554 9760 -22550
rect 9688 -22606 9698 -22554
rect 9750 -22606 9760 -22554
rect 9688 -22610 9760 -22606
rect 7134 -22648 7206 -22644
rect 7134 -22700 7144 -22648
rect 7196 -22700 7206 -22648
rect 7134 -22704 7206 -22700
rect 8156 -22648 8228 -22644
rect 8156 -22700 8166 -22648
rect 8218 -22700 8228 -22648
rect 8156 -22704 8228 -22700
rect 7140 -22740 7200 -22704
rect 8162 -22740 8222 -22704
rect 6934 -22746 7422 -22740
rect 6934 -22780 6981 -22746
rect 7015 -22780 7053 -22746
rect 7087 -22780 7125 -22746
rect 7159 -22780 7197 -22746
rect 7231 -22780 7269 -22746
rect 7303 -22780 7341 -22746
rect 7375 -22780 7422 -22746
rect 6934 -22786 7422 -22780
rect 7952 -22746 8440 -22740
rect 7952 -22780 7999 -22746
rect 8033 -22780 8071 -22746
rect 8105 -22780 8143 -22746
rect 8177 -22780 8215 -22746
rect 8249 -22780 8287 -22746
rect 8321 -22780 8359 -22746
rect 8393 -22780 8440 -22746
rect 7952 -22786 8440 -22780
rect 6638 -22880 6652 -22849
rect 3592 -22955 3598 -22921
rect 3632 -22955 3638 -22921
rect 3592 -22993 3638 -22955
rect 3592 -23027 3598 -22993
rect 3632 -23027 3638 -22993
rect 3592 -23065 3638 -23027
rect 3592 -23099 3598 -23065
rect 3632 -23099 3638 -23065
rect 3592 -23137 3638 -23099
rect 3592 -23171 3598 -23137
rect 3632 -23171 3638 -23137
rect 3592 -23209 3638 -23171
rect 3592 -23243 3598 -23209
rect 3632 -23243 3638 -23209
rect 3592 -23281 3638 -23243
rect 3592 -23315 3598 -23281
rect 3632 -23315 3638 -23281
rect 3592 -23352 3638 -23315
rect 4610 -22921 4656 -22890
rect 4610 -22955 4616 -22921
rect 4650 -22955 4656 -22921
rect 4610 -22993 4656 -22955
rect 4610 -23027 4616 -22993
rect 4650 -23027 4656 -22993
rect 4610 -23065 4656 -23027
rect 4610 -23099 4616 -23065
rect 4650 -23099 4656 -23065
rect 4610 -23137 4656 -23099
rect 4610 -23171 4616 -23137
rect 4650 -23171 4656 -23137
rect 4610 -23209 4656 -23171
rect 4610 -23243 4616 -23209
rect 4650 -23243 4656 -23209
rect 4610 -23281 4656 -23243
rect 4610 -23315 4616 -23281
rect 4650 -23315 4656 -23281
rect 2574 -23380 2580 -23353
rect 2568 -23387 2580 -23380
rect 2614 -23380 2620 -23353
rect 3580 -23353 3640 -23352
rect 2614 -23387 2628 -23380
rect 2568 -23544 2628 -23387
rect 3580 -23387 3598 -23353
rect 3632 -23387 3640 -23353
rect 2862 -23456 3350 -23450
rect 2862 -23490 2909 -23456
rect 2943 -23490 2981 -23456
rect 3015 -23490 3053 -23456
rect 3087 -23490 3125 -23456
rect 3159 -23490 3197 -23456
rect 3231 -23490 3269 -23456
rect 3303 -23490 3350 -23456
rect 2862 -23496 3350 -23490
rect 3082 -23544 3142 -23496
rect 3580 -23544 3640 -23387
rect 4610 -23353 4656 -23315
rect 4610 -23387 4616 -23353
rect 4650 -23387 4656 -23353
rect 5628 -22921 5674 -22883
rect 5628 -22955 5634 -22921
rect 5668 -22955 5674 -22921
rect 5628 -22993 5674 -22955
rect 5628 -23027 5634 -22993
rect 5668 -23027 5674 -22993
rect 5628 -23065 5674 -23027
rect 5628 -23099 5634 -23065
rect 5668 -23099 5674 -23065
rect 5628 -23137 5674 -23099
rect 5628 -23171 5634 -23137
rect 5668 -23171 5674 -23137
rect 5628 -23209 5674 -23171
rect 5628 -23243 5634 -23209
rect 5668 -23243 5674 -23209
rect 5628 -23281 5674 -23243
rect 5628 -23315 5634 -23281
rect 5668 -23315 5674 -23281
rect 5628 -23353 5674 -23315
rect 6646 -22883 6652 -22880
rect 6686 -22880 6698 -22849
rect 7664 -22849 7710 -22818
rect 6686 -22883 6692 -22880
rect 6646 -22921 6692 -22883
rect 6646 -22955 6652 -22921
rect 6686 -22955 6692 -22921
rect 6646 -22993 6692 -22955
rect 6646 -23027 6652 -22993
rect 6686 -23027 6692 -22993
rect 6646 -23065 6692 -23027
rect 6646 -23099 6652 -23065
rect 6686 -23099 6692 -23065
rect 6646 -23137 6692 -23099
rect 6646 -23171 6652 -23137
rect 6686 -23171 6692 -23137
rect 6646 -23209 6692 -23171
rect 6646 -23243 6652 -23209
rect 6686 -23243 6692 -23209
rect 6646 -23281 6692 -23243
rect 6646 -23315 6652 -23281
rect 6686 -23315 6692 -23281
rect 6646 -23344 6692 -23315
rect 7664 -22883 7670 -22849
rect 7704 -22883 7710 -22849
rect 7664 -22921 7710 -22883
rect 7664 -22955 7670 -22921
rect 7704 -22955 7710 -22921
rect 7664 -22993 7710 -22955
rect 7664 -23027 7670 -22993
rect 7704 -23027 7710 -22993
rect 7664 -23065 7710 -23027
rect 7664 -23099 7670 -23065
rect 7704 -23099 7710 -23065
rect 7664 -23137 7710 -23099
rect 7664 -23171 7670 -23137
rect 7704 -23171 7710 -23137
rect 7664 -23209 7710 -23171
rect 7664 -23243 7670 -23209
rect 7704 -23243 7710 -23209
rect 7664 -23281 7710 -23243
rect 7664 -23315 7670 -23281
rect 7704 -23315 7710 -23281
rect 5628 -23362 5634 -23353
rect 4610 -23418 4656 -23387
rect 5622 -23387 5634 -23362
rect 5668 -23362 5674 -23353
rect 6636 -23353 6696 -23344
rect 5668 -23387 5682 -23362
rect 3880 -23456 4368 -23450
rect 3880 -23490 3927 -23456
rect 3961 -23490 3999 -23456
rect 4033 -23490 4071 -23456
rect 4105 -23490 4143 -23456
rect 4177 -23490 4215 -23456
rect 4249 -23490 4287 -23456
rect 4321 -23490 4368 -23456
rect 3880 -23496 4368 -23490
rect 4898 -23456 5386 -23450
rect 4898 -23490 4945 -23456
rect 4979 -23490 5017 -23456
rect 5051 -23490 5089 -23456
rect 5123 -23490 5161 -23456
rect 5195 -23490 5233 -23456
rect 5267 -23490 5305 -23456
rect 5339 -23490 5386 -23456
rect 4898 -23496 5386 -23490
rect 2562 -23548 2634 -23544
rect 2562 -23600 2572 -23548
rect 2624 -23600 2634 -23548
rect 2562 -23604 2634 -23600
rect 3076 -23548 3148 -23544
rect 3076 -23600 3086 -23548
rect 3138 -23600 3148 -23548
rect 3076 -23604 3148 -23600
rect 3574 -23548 3646 -23544
rect 3574 -23600 3584 -23548
rect 3636 -23600 3646 -23548
rect 3574 -23604 3646 -23600
rect 4096 -23762 4156 -23496
rect 5118 -23762 5178 -23496
rect 5622 -23544 5682 -23387
rect 6636 -23387 6652 -23353
rect 6686 -23387 6696 -23353
rect 7664 -23353 7710 -23315
rect 7664 -23366 7670 -23353
rect 5916 -23456 6404 -23450
rect 5916 -23490 5963 -23456
rect 5997 -23490 6035 -23456
rect 6069 -23490 6107 -23456
rect 6141 -23490 6179 -23456
rect 6213 -23490 6251 -23456
rect 6285 -23490 6323 -23456
rect 6357 -23490 6404 -23456
rect 5916 -23496 6404 -23490
rect 5616 -23548 5688 -23544
rect 5616 -23600 5626 -23548
rect 5678 -23600 5688 -23548
rect 5616 -23604 5688 -23600
rect 6130 -23656 6190 -23496
rect 6124 -23660 6196 -23656
rect 6124 -23712 6134 -23660
rect 6186 -23712 6196 -23660
rect 6124 -23716 6196 -23712
rect 2104 -23766 2176 -23762
rect 2104 -23818 2114 -23766
rect 2166 -23818 2176 -23766
rect 2104 -23822 2176 -23818
rect 4090 -23766 4162 -23762
rect 4090 -23818 4100 -23766
rect 4152 -23818 4162 -23766
rect 4090 -23822 4162 -23818
rect 5112 -23766 5184 -23762
rect 5112 -23818 5122 -23766
rect 5174 -23818 5184 -23766
rect 5112 -23822 5184 -23818
rect 6636 -23866 6696 -23387
rect 7654 -23387 7670 -23366
rect 7704 -23366 7710 -23353
rect 8674 -22849 8734 -22610
rect 10204 -22644 10264 -22262
rect 11220 -22428 11280 -22262
rect 11724 -22314 11784 -22153
rect 12754 -22153 12760 -22119
rect 12794 -22153 12800 -22119
rect 13772 -21649 13778 -21615
rect 13812 -21649 13818 -21615
rect 14786 -21615 14846 -21332
rect 15282 -21506 15342 -21230
rect 15078 -21512 15566 -21506
rect 15078 -21546 15125 -21512
rect 15159 -21546 15197 -21512
rect 15231 -21546 15269 -21512
rect 15303 -21546 15341 -21512
rect 15375 -21546 15413 -21512
rect 15447 -21546 15485 -21512
rect 15519 -21546 15566 -21512
rect 15078 -21552 15566 -21546
rect 14786 -21644 14796 -21615
rect 13772 -21687 13818 -21649
rect 13772 -21721 13778 -21687
rect 13812 -21721 13818 -21687
rect 13772 -21759 13818 -21721
rect 13772 -21793 13778 -21759
rect 13812 -21793 13818 -21759
rect 13772 -21831 13818 -21793
rect 13772 -21865 13778 -21831
rect 13812 -21865 13818 -21831
rect 13772 -21903 13818 -21865
rect 13772 -21937 13778 -21903
rect 13812 -21937 13818 -21903
rect 13772 -21975 13818 -21937
rect 13772 -22009 13778 -21975
rect 13812 -22009 13818 -21975
rect 13772 -22047 13818 -22009
rect 13772 -22081 13778 -22047
rect 13812 -22081 13818 -22047
rect 13772 -22119 13818 -22081
rect 13772 -22120 13778 -22119
rect 12754 -22184 12800 -22153
rect 13766 -22153 13778 -22120
rect 13812 -22120 13818 -22119
rect 14790 -21649 14796 -21644
rect 14830 -21644 14846 -21615
rect 15800 -21615 15860 -21222
rect 16308 -21506 16368 -21130
rect 16808 -21276 16880 -21272
rect 16808 -21328 16818 -21276
rect 16870 -21328 16880 -21276
rect 16808 -21332 16880 -21328
rect 16096 -21512 16584 -21506
rect 16096 -21546 16143 -21512
rect 16177 -21546 16215 -21512
rect 16249 -21546 16287 -21512
rect 16321 -21546 16359 -21512
rect 16393 -21546 16431 -21512
rect 16465 -21546 16503 -21512
rect 16537 -21546 16584 -21512
rect 16096 -21552 16584 -21546
rect 15800 -21632 15814 -21615
rect 14830 -21649 14836 -21644
rect 14790 -21687 14836 -21649
rect 14790 -21721 14796 -21687
rect 14830 -21721 14836 -21687
rect 14790 -21759 14836 -21721
rect 14790 -21793 14796 -21759
rect 14830 -21793 14836 -21759
rect 14790 -21831 14836 -21793
rect 14790 -21865 14796 -21831
rect 14830 -21865 14836 -21831
rect 14790 -21903 14836 -21865
rect 14790 -21937 14796 -21903
rect 14830 -21937 14836 -21903
rect 14790 -21975 14836 -21937
rect 14790 -22009 14796 -21975
rect 14830 -22009 14836 -21975
rect 14790 -22047 14836 -22009
rect 14790 -22081 14796 -22047
rect 14830 -22081 14836 -22047
rect 14790 -22119 14836 -22081
rect 13812 -22153 13826 -22120
rect 12024 -22222 12512 -22216
rect 12024 -22256 12071 -22222
rect 12105 -22256 12143 -22222
rect 12177 -22256 12215 -22222
rect 12249 -22256 12287 -22222
rect 12321 -22256 12359 -22222
rect 12393 -22256 12431 -22222
rect 12465 -22256 12512 -22222
rect 12024 -22262 12512 -22256
rect 13042 -22222 13530 -22216
rect 13042 -22256 13089 -22222
rect 13123 -22256 13161 -22222
rect 13195 -22256 13233 -22222
rect 13267 -22256 13305 -22222
rect 13339 -22256 13377 -22222
rect 13411 -22256 13449 -22222
rect 13483 -22256 13530 -22222
rect 13042 -22262 13530 -22256
rect 13766 -22314 13826 -22153
rect 14790 -22153 14796 -22119
rect 14830 -22153 14836 -22119
rect 15808 -21649 15814 -21632
rect 15848 -21632 15860 -21615
rect 16814 -21615 16874 -21332
rect 17328 -21506 17388 -21030
rect 17840 -21398 17900 -20921
rect 18852 -20921 18868 -20896
rect 18902 -20896 18908 -20887
rect 19880 -20455 19926 -20422
rect 19880 -20489 19886 -20455
rect 19920 -20489 19926 -20455
rect 19880 -20527 19926 -20489
rect 19880 -20561 19886 -20527
rect 19920 -20561 19926 -20527
rect 19880 -20599 19926 -20561
rect 19880 -20633 19886 -20599
rect 19920 -20633 19926 -20599
rect 19880 -20671 19926 -20633
rect 19880 -20705 19886 -20671
rect 19920 -20705 19926 -20671
rect 19880 -20743 19926 -20705
rect 19880 -20777 19886 -20743
rect 19920 -20777 19926 -20743
rect 19880 -20815 19926 -20777
rect 19880 -20849 19886 -20815
rect 19920 -20849 19926 -20815
rect 19880 -20887 19926 -20849
rect 20898 -20455 20944 -20417
rect 20898 -20489 20904 -20455
rect 20938 -20489 20944 -20455
rect 20898 -20527 20944 -20489
rect 20898 -20561 20904 -20527
rect 20938 -20561 20944 -20527
rect 20898 -20599 20944 -20561
rect 20898 -20633 20904 -20599
rect 20938 -20633 20944 -20599
rect 20898 -20671 20944 -20633
rect 20898 -20705 20904 -20671
rect 20938 -20705 20944 -20671
rect 20898 -20743 20944 -20705
rect 20898 -20777 20904 -20743
rect 20938 -20777 20944 -20743
rect 20898 -20815 20944 -20777
rect 20898 -20849 20904 -20815
rect 20938 -20849 20944 -20815
rect 20898 -20886 20944 -20849
rect 21916 -20417 21922 -20383
rect 21956 -20417 21962 -20383
rect 21916 -20455 21962 -20417
rect 21916 -20489 21922 -20455
rect 21956 -20489 21962 -20455
rect 21916 -20527 21962 -20489
rect 21916 -20561 21922 -20527
rect 21956 -20561 21962 -20527
rect 21916 -20599 21962 -20561
rect 21916 -20633 21922 -20599
rect 21956 -20633 21962 -20599
rect 21916 -20671 21962 -20633
rect 21916 -20705 21922 -20671
rect 21956 -20705 21962 -20671
rect 21916 -20743 21962 -20705
rect 21916 -20777 21922 -20743
rect 21956 -20777 21962 -20743
rect 21916 -20815 21962 -20777
rect 21916 -20849 21922 -20815
rect 21956 -20849 21962 -20815
rect 18902 -20921 18912 -20896
rect 19880 -20900 19886 -20887
rect 18132 -20990 18620 -20984
rect 18132 -21024 18179 -20990
rect 18213 -21024 18251 -20990
rect 18285 -21024 18323 -20990
rect 18357 -21024 18395 -20990
rect 18429 -21024 18467 -20990
rect 18501 -21024 18539 -20990
rect 18573 -21024 18620 -20990
rect 18132 -21030 18620 -21024
rect 17834 -21402 17906 -21398
rect 17834 -21454 17844 -21402
rect 17896 -21454 17906 -21402
rect 17834 -21458 17906 -21454
rect 17114 -21512 17602 -21506
rect 17114 -21546 17161 -21512
rect 17195 -21546 17233 -21512
rect 17267 -21546 17305 -21512
rect 17339 -21546 17377 -21512
rect 17411 -21546 17449 -21512
rect 17483 -21546 17521 -21512
rect 17555 -21546 17602 -21512
rect 17114 -21552 17602 -21546
rect 15848 -21649 15854 -21632
rect 16814 -21644 16832 -21615
rect 15808 -21687 15854 -21649
rect 15808 -21721 15814 -21687
rect 15848 -21721 15854 -21687
rect 15808 -21759 15854 -21721
rect 15808 -21793 15814 -21759
rect 15848 -21793 15854 -21759
rect 15808 -21831 15854 -21793
rect 15808 -21865 15814 -21831
rect 15848 -21865 15854 -21831
rect 15808 -21903 15854 -21865
rect 15808 -21937 15814 -21903
rect 15848 -21937 15854 -21903
rect 15808 -21975 15854 -21937
rect 15808 -22009 15814 -21975
rect 15848 -22009 15854 -21975
rect 15808 -22047 15854 -22009
rect 15808 -22081 15814 -22047
rect 15848 -22081 15854 -22047
rect 15808 -22119 15854 -22081
rect 15808 -22128 15814 -22119
rect 14790 -22184 14836 -22153
rect 15802 -22153 15814 -22128
rect 15848 -22128 15854 -22119
rect 16826 -21649 16832 -21644
rect 16866 -21644 16874 -21615
rect 17840 -21615 17900 -21458
rect 18344 -21506 18404 -21030
rect 18852 -21272 18912 -20921
rect 19870 -20921 19886 -20900
rect 19920 -20900 19926 -20887
rect 20892 -20887 20952 -20886
rect 19920 -20921 19930 -20900
rect 19150 -20990 19638 -20984
rect 19150 -21024 19197 -20990
rect 19231 -21024 19269 -20990
rect 19303 -21024 19341 -20990
rect 19375 -21024 19413 -20990
rect 19447 -21024 19485 -20990
rect 19519 -21024 19557 -20990
rect 19591 -21024 19638 -20990
rect 19150 -21030 19638 -21024
rect 18846 -21276 18918 -21272
rect 18846 -21328 18856 -21276
rect 18908 -21328 18918 -21276
rect 18846 -21332 18918 -21328
rect 19378 -21506 19438 -21030
rect 19870 -21398 19930 -20921
rect 20892 -20921 20904 -20887
rect 20938 -20921 20952 -20887
rect 21916 -20887 21962 -20849
rect 21916 -20894 21922 -20887
rect 20168 -20990 20656 -20984
rect 20168 -21024 20215 -20990
rect 20249 -21024 20287 -20990
rect 20321 -21024 20359 -20990
rect 20393 -21024 20431 -20990
rect 20465 -21024 20503 -20990
rect 20537 -21024 20575 -20990
rect 20609 -21024 20656 -20990
rect 20168 -21030 20656 -21024
rect 19864 -21402 19936 -21398
rect 19864 -21454 19874 -21402
rect 19926 -21454 19936 -21402
rect 19864 -21458 19936 -21454
rect 20396 -21400 20456 -21030
rect 20892 -21272 20952 -20921
rect 21906 -20921 21922 -20894
rect 21956 -20894 21962 -20887
rect 22934 -20383 22980 -20352
rect 22934 -20417 22940 -20383
rect 22974 -20417 22980 -20383
rect 22934 -20455 22980 -20417
rect 22934 -20489 22940 -20455
rect 22974 -20489 22980 -20455
rect 22934 -20527 22980 -20489
rect 22934 -20561 22940 -20527
rect 22974 -20561 22980 -20527
rect 22934 -20599 22980 -20561
rect 22934 -20633 22940 -20599
rect 22974 -20633 22980 -20599
rect 22934 -20671 22980 -20633
rect 22934 -20705 22940 -20671
rect 22974 -20705 22980 -20671
rect 22934 -20743 22980 -20705
rect 22934 -20777 22940 -20743
rect 22974 -20777 22980 -20743
rect 22934 -20815 22980 -20777
rect 22934 -20849 22940 -20815
rect 22974 -20849 22980 -20815
rect 22934 -20887 22980 -20849
rect 21956 -20921 21966 -20894
rect 22934 -20912 22940 -20887
rect 21186 -20990 21674 -20984
rect 21186 -21024 21233 -20990
rect 21267 -21024 21305 -20990
rect 21339 -21024 21377 -20990
rect 21411 -21024 21449 -20990
rect 21483 -21024 21521 -20990
rect 21555 -21024 21593 -20990
rect 21627 -21024 21674 -20990
rect 21186 -21030 21674 -21024
rect 21410 -21268 21470 -21030
rect 21906 -21066 21966 -20921
rect 22926 -20921 22940 -20912
rect 22974 -20912 22980 -20887
rect 22974 -20921 22986 -20912
rect 22204 -20990 22692 -20984
rect 22204 -21024 22251 -20990
rect 22285 -21024 22323 -20990
rect 22357 -21024 22395 -20990
rect 22429 -21024 22467 -20990
rect 22501 -21024 22539 -20990
rect 22573 -21024 22611 -20990
rect 22645 -21024 22692 -20990
rect 22204 -21030 22692 -21024
rect 22412 -21064 22472 -21030
rect 22926 -21064 22986 -20921
rect 22412 -21066 22986 -21064
rect 21906 -21126 22986 -21066
rect 21906 -21162 21966 -21126
rect 21900 -21166 21972 -21162
rect 21900 -21218 21910 -21166
rect 21962 -21218 21972 -21166
rect 21900 -21222 21972 -21218
rect 21404 -21272 21476 -21268
rect 20886 -21276 20958 -21272
rect 20886 -21328 20896 -21276
rect 20948 -21328 20958 -21276
rect 21404 -21324 21414 -21272
rect 21466 -21324 21476 -21272
rect 21404 -21328 21476 -21324
rect 20886 -21332 20958 -21328
rect 20396 -21452 20400 -21400
rect 20452 -21452 20456 -21400
rect 18132 -21512 18620 -21506
rect 18132 -21546 18179 -21512
rect 18213 -21546 18251 -21512
rect 18285 -21546 18323 -21512
rect 18357 -21546 18395 -21512
rect 18429 -21546 18467 -21512
rect 18501 -21546 18539 -21512
rect 18573 -21546 18620 -21512
rect 18132 -21552 18620 -21546
rect 19150 -21512 19638 -21506
rect 19150 -21546 19197 -21512
rect 19231 -21546 19269 -21512
rect 19303 -21546 19341 -21512
rect 19375 -21546 19413 -21512
rect 19447 -21546 19485 -21512
rect 19519 -21546 19557 -21512
rect 19591 -21546 19638 -21512
rect 19150 -21552 19638 -21546
rect 17840 -21642 17850 -21615
rect 16866 -21649 16872 -21644
rect 16826 -21687 16872 -21649
rect 16826 -21721 16832 -21687
rect 16866 -21721 16872 -21687
rect 16826 -21759 16872 -21721
rect 16826 -21793 16832 -21759
rect 16866 -21793 16872 -21759
rect 16826 -21831 16872 -21793
rect 16826 -21865 16832 -21831
rect 16866 -21865 16872 -21831
rect 16826 -21903 16872 -21865
rect 16826 -21937 16832 -21903
rect 16866 -21937 16872 -21903
rect 16826 -21975 16872 -21937
rect 16826 -22009 16832 -21975
rect 16866 -22009 16872 -21975
rect 16826 -22047 16872 -22009
rect 16826 -22081 16832 -22047
rect 16866 -22081 16872 -22047
rect 16826 -22119 16872 -22081
rect 17844 -21649 17850 -21642
rect 17884 -21642 17900 -21615
rect 18862 -21615 18908 -21584
rect 17884 -21649 17890 -21642
rect 17844 -21687 17890 -21649
rect 17844 -21721 17850 -21687
rect 17884 -21721 17890 -21687
rect 17844 -21759 17890 -21721
rect 17844 -21793 17850 -21759
rect 17884 -21793 17890 -21759
rect 17844 -21831 17890 -21793
rect 17844 -21865 17850 -21831
rect 17884 -21865 17890 -21831
rect 17844 -21903 17890 -21865
rect 17844 -21937 17850 -21903
rect 17884 -21937 17890 -21903
rect 17844 -21975 17890 -21937
rect 17844 -22009 17850 -21975
rect 17884 -22009 17890 -21975
rect 17844 -22047 17890 -22009
rect 17844 -22081 17850 -22047
rect 17884 -22081 17890 -22047
rect 17844 -22112 17890 -22081
rect 18862 -21649 18868 -21615
rect 18902 -21649 18908 -21615
rect 19870 -21615 19930 -21458
rect 20396 -21506 20456 -21452
rect 21410 -21506 21470 -21328
rect 21908 -21396 22986 -21338
rect 21902 -21398 22986 -21396
rect 21902 -21400 21974 -21398
rect 21902 -21452 21912 -21400
rect 21964 -21452 21974 -21400
rect 21902 -21456 21974 -21452
rect 20168 -21512 20656 -21506
rect 20168 -21546 20215 -21512
rect 20249 -21546 20287 -21512
rect 20321 -21546 20359 -21512
rect 20393 -21546 20431 -21512
rect 20465 -21546 20503 -21512
rect 20537 -21546 20575 -21512
rect 20609 -21546 20656 -21512
rect 20168 -21552 20656 -21546
rect 21186 -21512 21674 -21506
rect 21186 -21546 21233 -21512
rect 21267 -21546 21305 -21512
rect 21339 -21546 21377 -21512
rect 21411 -21546 21449 -21512
rect 21483 -21546 21521 -21512
rect 21555 -21546 21593 -21512
rect 21627 -21546 21674 -21512
rect 21186 -21552 21674 -21546
rect 19870 -21642 19886 -21615
rect 18862 -21687 18908 -21649
rect 18862 -21721 18868 -21687
rect 18902 -21721 18908 -21687
rect 18862 -21759 18908 -21721
rect 18862 -21793 18868 -21759
rect 18902 -21793 18908 -21759
rect 18862 -21831 18908 -21793
rect 18862 -21865 18868 -21831
rect 18902 -21865 18908 -21831
rect 18862 -21903 18908 -21865
rect 18862 -21937 18868 -21903
rect 18902 -21937 18908 -21903
rect 18862 -21975 18908 -21937
rect 18862 -22009 18868 -21975
rect 18902 -22009 18908 -21975
rect 18862 -22047 18908 -22009
rect 18862 -22081 18868 -22047
rect 18902 -22081 18908 -22047
rect 15848 -22153 15862 -22128
rect 14060 -22222 14548 -22216
rect 14060 -22256 14107 -22222
rect 14141 -22256 14179 -22222
rect 14213 -22256 14251 -22222
rect 14285 -22256 14323 -22222
rect 14357 -22256 14395 -22222
rect 14429 -22256 14467 -22222
rect 14501 -22256 14548 -22222
rect 14060 -22262 14548 -22256
rect 15078 -22222 15566 -22216
rect 15078 -22256 15125 -22222
rect 15159 -22256 15197 -22222
rect 15231 -22256 15269 -22222
rect 15303 -22256 15341 -22222
rect 15375 -22256 15413 -22222
rect 15447 -22256 15485 -22222
rect 15519 -22256 15566 -22222
rect 15078 -22262 15566 -22256
rect 15802 -22314 15862 -22153
rect 16826 -22153 16832 -22119
rect 16866 -22153 16872 -22119
rect 16826 -22184 16872 -22153
rect 17838 -22119 17898 -22112
rect 17838 -22153 17850 -22119
rect 17884 -22153 17898 -22119
rect 18862 -22119 18908 -22081
rect 18862 -22128 18868 -22119
rect 16096 -22222 16584 -22216
rect 16096 -22256 16143 -22222
rect 16177 -22256 16215 -22222
rect 16249 -22256 16287 -22222
rect 16321 -22256 16359 -22222
rect 16393 -22256 16431 -22222
rect 16465 -22256 16503 -22222
rect 16537 -22256 16584 -22222
rect 16096 -22262 16584 -22256
rect 17114 -22222 17602 -22216
rect 17114 -22256 17161 -22222
rect 17195 -22256 17233 -22222
rect 17267 -22256 17305 -22222
rect 17339 -22256 17377 -22222
rect 17411 -22256 17449 -22222
rect 17483 -22256 17521 -22222
rect 17555 -22256 17602 -22222
rect 17114 -22262 17602 -22256
rect 11718 -22318 11790 -22314
rect 11718 -22370 11728 -22318
rect 11780 -22370 11790 -22318
rect 11718 -22374 11790 -22370
rect 13760 -22318 13832 -22314
rect 13760 -22370 13770 -22318
rect 13822 -22370 13832 -22318
rect 13760 -22374 13832 -22370
rect 15796 -22318 15868 -22314
rect 15796 -22370 15806 -22318
rect 15858 -22370 15868 -22318
rect 15796 -22374 15868 -22370
rect 16308 -22424 16368 -22262
rect 16302 -22428 16374 -22424
rect 11214 -22432 11286 -22428
rect 11214 -22484 11224 -22432
rect 11276 -22484 11286 -22432
rect 16302 -22480 16312 -22428
rect 16364 -22480 16374 -22428
rect 16302 -22484 16374 -22480
rect 11214 -22488 11286 -22484
rect 10706 -22554 10778 -22550
rect 10706 -22606 10716 -22554
rect 10768 -22606 10778 -22554
rect 10706 -22610 10778 -22606
rect 12736 -22554 12808 -22550
rect 12736 -22606 12746 -22554
rect 12798 -22606 12808 -22554
rect 12736 -22610 12808 -22606
rect 14774 -22554 14846 -22550
rect 14774 -22606 14784 -22554
rect 14836 -22606 14846 -22554
rect 14774 -22610 14846 -22606
rect 16810 -22554 16882 -22550
rect 16810 -22606 16820 -22554
rect 16872 -22606 16882 -22554
rect 16810 -22610 16882 -22606
rect 10198 -22648 10270 -22644
rect 10198 -22700 10208 -22648
rect 10260 -22700 10270 -22648
rect 10198 -22704 10270 -22700
rect 8970 -22746 9458 -22740
rect 8970 -22780 9017 -22746
rect 9051 -22780 9089 -22746
rect 9123 -22780 9161 -22746
rect 9195 -22780 9233 -22746
rect 9267 -22780 9305 -22746
rect 9339 -22780 9377 -22746
rect 9411 -22780 9458 -22746
rect 8970 -22786 9458 -22780
rect 9988 -22746 10476 -22740
rect 9988 -22780 10035 -22746
rect 10069 -22780 10107 -22746
rect 10141 -22780 10179 -22746
rect 10213 -22780 10251 -22746
rect 10285 -22780 10323 -22746
rect 10357 -22780 10395 -22746
rect 10429 -22780 10476 -22746
rect 9988 -22786 10476 -22780
rect 8674 -22883 8688 -22849
rect 8722 -22883 8734 -22849
rect 8674 -22921 8734 -22883
rect 8674 -22955 8688 -22921
rect 8722 -22955 8734 -22921
rect 8674 -22993 8734 -22955
rect 8674 -23027 8688 -22993
rect 8722 -23027 8734 -22993
rect 8674 -23065 8734 -23027
rect 8674 -23099 8688 -23065
rect 8722 -23099 8734 -23065
rect 8674 -23137 8734 -23099
rect 8674 -23171 8688 -23137
rect 8722 -23171 8734 -23137
rect 8674 -23209 8734 -23171
rect 8674 -23243 8688 -23209
rect 8722 -23243 8734 -23209
rect 8674 -23281 8734 -23243
rect 8674 -23315 8688 -23281
rect 8722 -23315 8734 -23281
rect 8674 -23353 8734 -23315
rect 7704 -23387 7714 -23366
rect 6934 -23456 7422 -23450
rect 6934 -23490 6981 -23456
rect 7015 -23490 7053 -23456
rect 7087 -23490 7125 -23456
rect 7159 -23490 7197 -23456
rect 7231 -23490 7269 -23456
rect 7303 -23490 7341 -23456
rect 7375 -23490 7422 -23456
rect 6934 -23496 7422 -23490
rect 7142 -23656 7202 -23496
rect 7654 -23544 7714 -23387
rect 8674 -23387 8688 -23353
rect 8722 -23387 8734 -23353
rect 9700 -22849 9746 -22818
rect 9700 -22883 9706 -22849
rect 9740 -22883 9746 -22849
rect 9700 -22921 9746 -22883
rect 10712 -22849 10772 -22610
rect 11218 -22686 12288 -22626
rect 11218 -22740 11278 -22686
rect 11006 -22746 11494 -22740
rect 11006 -22780 11053 -22746
rect 11087 -22780 11125 -22746
rect 11159 -22780 11197 -22746
rect 11231 -22780 11269 -22746
rect 11303 -22780 11341 -22746
rect 11375 -22780 11413 -22746
rect 11447 -22780 11494 -22746
rect 11006 -22786 11494 -22780
rect 10712 -22883 10724 -22849
rect 10758 -22883 10772 -22849
rect 11730 -22849 11790 -22686
rect 12228 -22740 12288 -22686
rect 12024 -22746 12512 -22740
rect 12024 -22780 12071 -22746
rect 12105 -22780 12143 -22746
rect 12177 -22780 12215 -22746
rect 12249 -22780 12287 -22746
rect 12321 -22780 12359 -22746
rect 12393 -22780 12431 -22746
rect 12465 -22780 12512 -22746
rect 12024 -22786 12512 -22780
rect 11730 -22866 11742 -22849
rect 10712 -22886 10772 -22883
rect 11736 -22883 11742 -22866
rect 11776 -22866 11790 -22849
rect 12742 -22849 12802 -22610
rect 13242 -22682 14330 -22622
rect 13242 -22740 13302 -22682
rect 13042 -22746 13530 -22740
rect 13042 -22780 13089 -22746
rect 13123 -22780 13161 -22746
rect 13195 -22780 13233 -22746
rect 13267 -22780 13305 -22746
rect 13339 -22780 13377 -22746
rect 13411 -22780 13449 -22746
rect 13483 -22780 13530 -22746
rect 13042 -22786 13530 -22780
rect 11776 -22883 11782 -22866
rect 12742 -22880 12760 -22849
rect 9700 -22955 9706 -22921
rect 9740 -22955 9746 -22921
rect 9700 -22993 9746 -22955
rect 9700 -23027 9706 -22993
rect 9740 -23027 9746 -22993
rect 9700 -23065 9746 -23027
rect 9700 -23099 9706 -23065
rect 9740 -23099 9746 -23065
rect 9700 -23137 9746 -23099
rect 9700 -23171 9706 -23137
rect 9740 -23171 9746 -23137
rect 9700 -23209 9746 -23171
rect 9700 -23243 9706 -23209
rect 9740 -23243 9746 -23209
rect 9700 -23281 9746 -23243
rect 9700 -23315 9706 -23281
rect 9740 -23315 9746 -23281
rect 9700 -23353 9746 -23315
rect 9700 -23366 9706 -23353
rect 7952 -23456 8440 -23450
rect 7952 -23490 7999 -23456
rect 8033 -23490 8071 -23456
rect 8105 -23490 8143 -23456
rect 8177 -23490 8215 -23456
rect 8249 -23490 8287 -23456
rect 8321 -23490 8359 -23456
rect 8393 -23490 8440 -23456
rect 7952 -23496 8440 -23490
rect 7648 -23548 7720 -23544
rect 7648 -23600 7658 -23548
rect 7710 -23600 7720 -23548
rect 7648 -23604 7720 -23600
rect 8156 -23656 8216 -23496
rect 7136 -23660 7208 -23656
rect 7136 -23712 7146 -23660
rect 7198 -23712 7208 -23660
rect 7136 -23716 7208 -23712
rect 8150 -23660 8222 -23656
rect 8150 -23712 8160 -23660
rect 8212 -23712 8222 -23660
rect 8150 -23716 8222 -23712
rect 7650 -23766 7722 -23762
rect 7650 -23818 7660 -23766
rect 7712 -23818 7722 -23766
rect 7650 -23822 7722 -23818
rect 8162 -23766 8234 -23762
rect 8162 -23818 8172 -23766
rect 8224 -23818 8234 -23766
rect 8162 -23822 8234 -23818
rect 1698 -23870 1770 -23866
rect 1698 -23922 1708 -23870
rect 1760 -23922 1770 -23870
rect 1698 -23926 1770 -23922
rect 6126 -23870 6198 -23866
rect 6126 -23922 6136 -23870
rect 6188 -23922 6198 -23870
rect 6126 -23926 6198 -23922
rect 6630 -23870 6702 -23866
rect 6630 -23922 6640 -23870
rect 6692 -23922 6702 -23870
rect 6630 -23926 6702 -23922
rect 7146 -23870 7218 -23866
rect 7146 -23922 7156 -23870
rect 7208 -23922 7218 -23870
rect 7146 -23926 7218 -23922
rect 1070 -24918 1142 -24914
rect 1070 -24970 1080 -24918
rect 1132 -24970 1142 -24918
rect 1070 -24974 1142 -24970
rect -2132 -25944 -2060 -25940
rect -2132 -25996 -2122 -25944
rect -2070 -25996 -2060 -25944
rect -2132 -26000 -2060 -25996
rect -944 -25944 -872 -25940
rect -944 -25996 -934 -25944
rect -882 -25996 -872 -25944
rect -944 -26000 -872 -25996
rect 252 -25944 324 -25940
rect 252 -25996 262 -25944
rect 314 -25996 324 -25944
rect 252 -26000 324 -25996
rect 946 -25944 1018 -25940
rect 946 -25996 956 -25944
rect 1008 -25996 1018 -25944
rect 946 -26000 1018 -25996
rect 1704 -26430 1764 -23926
rect 6132 -23974 6192 -23926
rect 2862 -23980 3350 -23974
rect 2862 -24014 2909 -23980
rect 2943 -24014 2981 -23980
rect 3015 -24014 3053 -23980
rect 3087 -24014 3125 -23980
rect 3159 -24014 3197 -23980
rect 3231 -24014 3269 -23980
rect 3303 -24014 3350 -23980
rect 2862 -24020 3350 -24014
rect 3880 -23980 4368 -23974
rect 3880 -24014 3927 -23980
rect 3961 -24014 3999 -23980
rect 4033 -24014 4071 -23980
rect 4105 -24014 4143 -23980
rect 4177 -24014 4215 -23980
rect 4249 -24014 4287 -23980
rect 4321 -24014 4368 -23980
rect 3880 -24020 4368 -24014
rect 4898 -23980 5386 -23974
rect 4898 -24014 4945 -23980
rect 4979 -24014 5017 -23980
rect 5051 -24014 5089 -23980
rect 5123 -24014 5161 -23980
rect 5195 -24014 5233 -23980
rect 5267 -24014 5305 -23980
rect 5339 -24014 5386 -23980
rect 4898 -24020 5386 -24014
rect 5916 -23980 6404 -23974
rect 5916 -24014 5963 -23980
rect 5997 -24014 6035 -23980
rect 6069 -24014 6107 -23980
rect 6141 -24014 6179 -23980
rect 6213 -24014 6251 -23980
rect 6285 -24014 6323 -23980
rect 6357 -24014 6404 -23980
rect 5916 -24020 6404 -24014
rect 2574 -24083 2620 -24052
rect 2574 -24117 2580 -24083
rect 2614 -24117 2620 -24083
rect 2574 -24155 2620 -24117
rect 2574 -24189 2580 -24155
rect 2614 -24189 2620 -24155
rect 2574 -24227 2620 -24189
rect 2574 -24261 2580 -24227
rect 2614 -24261 2620 -24227
rect 2574 -24299 2620 -24261
rect 2574 -24333 2580 -24299
rect 2614 -24333 2620 -24299
rect 2574 -24371 2620 -24333
rect 2574 -24405 2580 -24371
rect 2614 -24405 2620 -24371
rect 2574 -24443 2620 -24405
rect 2574 -24477 2580 -24443
rect 2614 -24477 2620 -24443
rect 2574 -24515 2620 -24477
rect 2574 -24549 2580 -24515
rect 2614 -24549 2620 -24515
rect 2574 -24587 2620 -24549
rect 2574 -24614 2580 -24587
rect 2568 -24621 2580 -24614
rect 2614 -24614 2620 -24587
rect 3592 -24083 3638 -24052
rect 3592 -24117 3598 -24083
rect 3632 -24117 3638 -24083
rect 3592 -24155 3638 -24117
rect 3592 -24189 3598 -24155
rect 3632 -24189 3638 -24155
rect 3592 -24227 3638 -24189
rect 3592 -24261 3598 -24227
rect 3632 -24261 3638 -24227
rect 3592 -24299 3638 -24261
rect 3592 -24333 3598 -24299
rect 3632 -24333 3638 -24299
rect 3592 -24371 3638 -24333
rect 3592 -24405 3598 -24371
rect 3632 -24405 3638 -24371
rect 3592 -24443 3638 -24405
rect 3592 -24477 3598 -24443
rect 3632 -24477 3638 -24443
rect 3592 -24515 3638 -24477
rect 3592 -24549 3598 -24515
rect 3632 -24549 3638 -24515
rect 3592 -24587 3638 -24549
rect 3592 -24612 3598 -24587
rect 2614 -24621 2628 -24614
rect 2568 -25096 2628 -24621
rect 3580 -24621 3598 -24612
rect 3632 -24612 3638 -24587
rect 4610 -24083 4656 -24052
rect 4610 -24117 4616 -24083
rect 4650 -24117 4656 -24083
rect 4610 -24155 4656 -24117
rect 4610 -24189 4616 -24155
rect 4650 -24189 4656 -24155
rect 4610 -24227 4656 -24189
rect 4610 -24261 4616 -24227
rect 4650 -24261 4656 -24227
rect 4610 -24299 4656 -24261
rect 4610 -24333 4616 -24299
rect 4650 -24333 4656 -24299
rect 4610 -24371 4656 -24333
rect 4610 -24405 4616 -24371
rect 4650 -24405 4656 -24371
rect 4610 -24443 4656 -24405
rect 4610 -24477 4616 -24443
rect 4650 -24477 4656 -24443
rect 4610 -24515 4656 -24477
rect 4610 -24549 4616 -24515
rect 4650 -24549 4656 -24515
rect 4610 -24587 4656 -24549
rect 4610 -24608 4616 -24587
rect 3632 -24621 3640 -24612
rect 2862 -24690 3350 -24684
rect 2862 -24724 2909 -24690
rect 2943 -24724 2981 -24690
rect 3015 -24724 3053 -24690
rect 3087 -24724 3125 -24690
rect 3159 -24724 3197 -24690
rect 3231 -24724 3269 -24690
rect 3303 -24724 3350 -24690
rect 2862 -24730 3350 -24724
rect 2562 -25100 2634 -25096
rect 2562 -25152 2572 -25100
rect 2624 -25152 2634 -25100
rect 2562 -25156 2634 -25152
rect 2568 -25315 2628 -25156
rect 3066 -25206 3126 -24730
rect 3580 -24998 3640 -24621
rect 4598 -24621 4616 -24608
rect 4650 -24608 4656 -24587
rect 5628 -24083 5674 -24052
rect 5628 -24117 5634 -24083
rect 5668 -24117 5674 -24083
rect 6636 -24083 6696 -23926
rect 7152 -23974 7212 -23926
rect 6934 -23980 7422 -23974
rect 6934 -24014 6981 -23980
rect 7015 -24014 7053 -23980
rect 7087 -24014 7125 -23980
rect 7159 -24014 7197 -23980
rect 7231 -24014 7269 -23980
rect 7303 -24014 7341 -23980
rect 7375 -24014 7422 -23980
rect 6934 -24020 7422 -24014
rect 7656 -24064 7716 -23822
rect 8168 -23974 8228 -23822
rect 8674 -23866 8734 -23387
rect 9686 -23387 9706 -23366
rect 9740 -23387 9746 -23353
rect 10718 -22921 10764 -22886
rect 10718 -22955 10724 -22921
rect 10758 -22955 10764 -22921
rect 10718 -22993 10764 -22955
rect 10718 -23027 10724 -22993
rect 10758 -23027 10764 -22993
rect 10718 -23065 10764 -23027
rect 10718 -23099 10724 -23065
rect 10758 -23099 10764 -23065
rect 10718 -23137 10764 -23099
rect 10718 -23171 10724 -23137
rect 10758 -23171 10764 -23137
rect 10718 -23209 10764 -23171
rect 10718 -23243 10724 -23209
rect 10758 -23243 10764 -23209
rect 10718 -23281 10764 -23243
rect 10718 -23315 10724 -23281
rect 10758 -23315 10764 -23281
rect 10718 -23353 10764 -23315
rect 10718 -23354 10724 -23353
rect 8970 -23456 9458 -23450
rect 8970 -23490 9017 -23456
rect 9051 -23490 9089 -23456
rect 9123 -23490 9161 -23456
rect 9195 -23490 9233 -23456
rect 9267 -23490 9305 -23456
rect 9339 -23490 9377 -23456
rect 9411 -23490 9458 -23456
rect 8970 -23496 9458 -23490
rect 9186 -23762 9246 -23496
rect 9686 -23544 9746 -23387
rect 10712 -23387 10724 -23354
rect 10758 -23354 10764 -23353
rect 11736 -22921 11782 -22883
rect 11736 -22955 11742 -22921
rect 11776 -22955 11782 -22921
rect 11736 -22993 11782 -22955
rect 11736 -23027 11742 -22993
rect 11776 -23027 11782 -22993
rect 11736 -23065 11782 -23027
rect 11736 -23099 11742 -23065
rect 11776 -23099 11782 -23065
rect 11736 -23137 11782 -23099
rect 11736 -23171 11742 -23137
rect 11776 -23171 11782 -23137
rect 11736 -23209 11782 -23171
rect 11736 -23243 11742 -23209
rect 11776 -23243 11782 -23209
rect 11736 -23281 11782 -23243
rect 11736 -23315 11742 -23281
rect 11776 -23315 11782 -23281
rect 11736 -23353 11782 -23315
rect 10758 -23387 10772 -23354
rect 11736 -23362 11742 -23353
rect 11728 -23370 11742 -23362
rect 9988 -23456 10476 -23450
rect 9988 -23490 10035 -23456
rect 10069 -23490 10107 -23456
rect 10141 -23490 10179 -23456
rect 10213 -23490 10251 -23456
rect 10285 -23490 10323 -23456
rect 10357 -23490 10395 -23456
rect 10429 -23490 10476 -23456
rect 9988 -23496 10476 -23490
rect 9680 -23548 9752 -23544
rect 9680 -23600 9690 -23548
rect 9742 -23600 9752 -23548
rect 9680 -23604 9752 -23600
rect 10198 -23762 10258 -23496
rect 9180 -23766 9252 -23762
rect 9180 -23818 9190 -23766
rect 9242 -23818 9252 -23766
rect 9180 -23822 9252 -23818
rect 9686 -23766 9758 -23762
rect 9686 -23818 9696 -23766
rect 9748 -23818 9758 -23766
rect 9686 -23822 9758 -23818
rect 10192 -23766 10264 -23762
rect 10192 -23818 10202 -23766
rect 10254 -23818 10264 -23766
rect 10192 -23822 10264 -23818
rect 8668 -23870 8740 -23866
rect 8668 -23922 8678 -23870
rect 8730 -23922 8740 -23870
rect 8668 -23926 8740 -23922
rect 7952 -23980 8440 -23974
rect 7952 -24014 7999 -23980
rect 8033 -24014 8071 -23980
rect 8105 -24014 8143 -23980
rect 8177 -24014 8215 -23980
rect 8249 -24014 8287 -23980
rect 8321 -24014 8359 -23980
rect 8393 -24014 8440 -23980
rect 7952 -24020 8440 -24014
rect 6636 -24116 6652 -24083
rect 5628 -24155 5674 -24117
rect 5628 -24189 5634 -24155
rect 5668 -24189 5674 -24155
rect 5628 -24227 5674 -24189
rect 5628 -24261 5634 -24227
rect 5668 -24261 5674 -24227
rect 5628 -24299 5674 -24261
rect 5628 -24333 5634 -24299
rect 5668 -24333 5674 -24299
rect 5628 -24371 5674 -24333
rect 5628 -24405 5634 -24371
rect 5668 -24405 5674 -24371
rect 5628 -24443 5674 -24405
rect 5628 -24477 5634 -24443
rect 5668 -24477 5674 -24443
rect 5628 -24515 5674 -24477
rect 5628 -24549 5634 -24515
rect 5668 -24549 5674 -24515
rect 5628 -24587 5674 -24549
rect 5628 -24600 5634 -24587
rect 4650 -24621 4658 -24608
rect 3880 -24690 4368 -24684
rect 3880 -24724 3927 -24690
rect 3961 -24724 3999 -24690
rect 4033 -24724 4071 -24690
rect 4105 -24724 4143 -24690
rect 4177 -24724 4215 -24690
rect 4249 -24724 4287 -24690
rect 4321 -24724 4368 -24690
rect 3880 -24730 4368 -24724
rect 3574 -25002 3646 -24998
rect 3574 -25054 3584 -25002
rect 3636 -25054 3646 -25002
rect 3574 -25058 3646 -25054
rect 2862 -25212 3350 -25206
rect 2862 -25246 2909 -25212
rect 2943 -25246 2981 -25212
rect 3015 -25246 3053 -25212
rect 3087 -25246 3125 -25212
rect 3159 -25246 3197 -25212
rect 3231 -25246 3269 -25212
rect 3303 -25246 3350 -25212
rect 2862 -25252 3350 -25246
rect 2568 -25349 2580 -25315
rect 2614 -25349 2628 -25315
rect 3580 -25315 3640 -25058
rect 4088 -25206 4148 -24730
rect 4598 -25096 4658 -24621
rect 5618 -24621 5634 -24600
rect 5668 -24600 5674 -24587
rect 6646 -24117 6652 -24116
rect 6686 -24116 6696 -24083
rect 7654 -24083 7716 -24064
rect 6686 -24117 6692 -24116
rect 6646 -24155 6692 -24117
rect 7654 -24117 7670 -24083
rect 7704 -24116 7716 -24083
rect 8674 -24083 8734 -23926
rect 9186 -23974 9246 -23822
rect 8970 -23980 9458 -23974
rect 8970 -24014 9017 -23980
rect 9051 -24014 9089 -23980
rect 9123 -24014 9161 -23980
rect 9195 -24014 9233 -23980
rect 9267 -24014 9305 -23980
rect 9339 -24014 9377 -23980
rect 9411 -24014 9458 -23980
rect 8970 -24020 9458 -24014
rect 9692 -24064 9752 -23822
rect 10198 -23974 10258 -23822
rect 10712 -23866 10772 -23387
rect 11722 -23387 11742 -23370
rect 11776 -23362 11782 -23353
rect 12754 -22883 12760 -22880
rect 12794 -22880 12802 -22849
rect 13766 -22849 13826 -22682
rect 14270 -22740 14330 -22682
rect 14060 -22746 14548 -22740
rect 14060 -22780 14107 -22746
rect 14141 -22780 14179 -22746
rect 14213 -22780 14251 -22746
rect 14285 -22780 14323 -22746
rect 14357 -22780 14395 -22746
rect 14429 -22780 14467 -22746
rect 14501 -22780 14548 -22746
rect 14060 -22786 14548 -22780
rect 13766 -22862 13778 -22849
rect 12794 -22883 12800 -22880
rect 12754 -22921 12800 -22883
rect 12754 -22955 12760 -22921
rect 12794 -22955 12800 -22921
rect 12754 -22993 12800 -22955
rect 12754 -23027 12760 -22993
rect 12794 -23027 12800 -22993
rect 12754 -23065 12800 -23027
rect 12754 -23099 12760 -23065
rect 12794 -23099 12800 -23065
rect 12754 -23137 12800 -23099
rect 12754 -23171 12760 -23137
rect 12794 -23171 12800 -23137
rect 12754 -23209 12800 -23171
rect 12754 -23243 12760 -23209
rect 12794 -23243 12800 -23209
rect 12754 -23281 12800 -23243
rect 12754 -23315 12760 -23281
rect 12794 -23315 12800 -23281
rect 12754 -23353 12800 -23315
rect 13772 -22883 13778 -22862
rect 13812 -22862 13826 -22849
rect 14780 -22849 14840 -22610
rect 15078 -22746 15566 -22740
rect 15078 -22780 15125 -22746
rect 15159 -22780 15197 -22746
rect 15231 -22780 15269 -22746
rect 15303 -22780 15341 -22746
rect 15375 -22780 15413 -22746
rect 15447 -22780 15485 -22746
rect 15519 -22780 15566 -22746
rect 15078 -22786 15566 -22780
rect 16096 -22746 16584 -22740
rect 16096 -22780 16143 -22746
rect 16177 -22780 16215 -22746
rect 16249 -22780 16287 -22746
rect 16321 -22780 16359 -22746
rect 16393 -22780 16431 -22746
rect 16465 -22780 16503 -22746
rect 16537 -22780 16584 -22746
rect 16096 -22786 16584 -22780
rect 13812 -22883 13818 -22862
rect 14780 -22874 14796 -22849
rect 13772 -22921 13818 -22883
rect 13772 -22955 13778 -22921
rect 13812 -22955 13818 -22921
rect 13772 -22993 13818 -22955
rect 13772 -23027 13778 -22993
rect 13812 -23027 13818 -22993
rect 13772 -23065 13818 -23027
rect 13772 -23099 13778 -23065
rect 13812 -23099 13818 -23065
rect 13772 -23137 13818 -23099
rect 13772 -23171 13778 -23137
rect 13812 -23171 13818 -23137
rect 13772 -23209 13818 -23171
rect 13772 -23243 13778 -23209
rect 13812 -23243 13818 -23209
rect 13772 -23281 13818 -23243
rect 13772 -23315 13778 -23281
rect 13812 -23315 13818 -23281
rect 13772 -23352 13818 -23315
rect 14790 -22883 14796 -22874
rect 14830 -22874 14840 -22849
rect 15808 -22849 15854 -22818
rect 14830 -22883 14836 -22874
rect 14790 -22921 14836 -22883
rect 14790 -22955 14796 -22921
rect 14830 -22955 14836 -22921
rect 14790 -22993 14836 -22955
rect 14790 -23027 14796 -22993
rect 14830 -23027 14836 -22993
rect 14790 -23065 14836 -23027
rect 14790 -23099 14796 -23065
rect 14830 -23099 14836 -23065
rect 14790 -23137 14836 -23099
rect 14790 -23171 14796 -23137
rect 14830 -23171 14836 -23137
rect 14790 -23209 14836 -23171
rect 14790 -23243 14796 -23209
rect 14830 -23243 14836 -23209
rect 14790 -23281 14836 -23243
rect 14790 -23315 14796 -23281
rect 14830 -23315 14836 -23281
rect 12754 -23356 12760 -23353
rect 11776 -23387 11788 -23362
rect 11722 -23406 11788 -23387
rect 11006 -23456 11494 -23450
rect 11006 -23490 11053 -23456
rect 11087 -23490 11125 -23456
rect 11159 -23490 11197 -23456
rect 11231 -23490 11269 -23456
rect 11303 -23490 11341 -23456
rect 11375 -23490 11413 -23456
rect 11447 -23490 11494 -23456
rect 11006 -23496 11494 -23490
rect 11062 -23660 11134 -23656
rect 11062 -23712 11072 -23660
rect 11124 -23712 11134 -23660
rect 11062 -23716 11134 -23712
rect 10706 -23870 10778 -23866
rect 10706 -23922 10716 -23870
rect 10768 -23922 10778 -23870
rect 10706 -23926 10778 -23922
rect 9988 -23980 10476 -23974
rect 9988 -24014 10035 -23980
rect 10069 -24014 10107 -23980
rect 10141 -24014 10179 -23980
rect 10213 -24014 10251 -23980
rect 10285 -24014 10323 -23980
rect 10357 -24014 10395 -23980
rect 10429 -24014 10476 -23980
rect 9988 -24020 10476 -24014
rect 8674 -24114 8688 -24083
rect 7704 -24117 7714 -24116
rect 7654 -24120 7714 -24117
rect 8682 -24117 8688 -24114
rect 8722 -24114 8734 -24083
rect 9686 -24083 9752 -24064
rect 8722 -24117 8728 -24114
rect 6646 -24189 6652 -24155
rect 6686 -24189 6692 -24155
rect 6646 -24227 6692 -24189
rect 6646 -24261 6652 -24227
rect 6686 -24261 6692 -24227
rect 6646 -24299 6692 -24261
rect 6646 -24333 6652 -24299
rect 6686 -24333 6692 -24299
rect 6646 -24371 6692 -24333
rect 6646 -24405 6652 -24371
rect 6686 -24405 6692 -24371
rect 6646 -24443 6692 -24405
rect 6646 -24477 6652 -24443
rect 6686 -24477 6692 -24443
rect 6646 -24515 6692 -24477
rect 6646 -24549 6652 -24515
rect 6686 -24549 6692 -24515
rect 6646 -24587 6692 -24549
rect 5668 -24621 5678 -24600
rect 4898 -24690 5386 -24684
rect 4898 -24724 4945 -24690
rect 4979 -24724 5017 -24690
rect 5051 -24724 5089 -24690
rect 5123 -24724 5161 -24690
rect 5195 -24724 5233 -24690
rect 5267 -24724 5305 -24690
rect 5339 -24724 5386 -24690
rect 4898 -24730 5386 -24724
rect 4592 -25100 4664 -25096
rect 4592 -25152 4602 -25100
rect 4654 -25152 4664 -25100
rect 4592 -25156 4664 -25152
rect 3880 -25212 4368 -25206
rect 3880 -25246 3927 -25212
rect 3961 -25246 3999 -25212
rect 4033 -25246 4071 -25212
rect 4105 -25246 4143 -25212
rect 4177 -25246 4215 -25212
rect 4249 -25246 4287 -25212
rect 4321 -25246 4368 -25212
rect 3880 -25252 4368 -25246
rect 3580 -25334 3598 -25315
rect 2568 -25352 2628 -25349
rect 3592 -25349 3598 -25334
rect 3632 -25334 3640 -25315
rect 4598 -25315 4658 -25156
rect 5114 -25206 5174 -24730
rect 5618 -24998 5678 -24621
rect 6646 -24621 6652 -24587
rect 6686 -24621 6692 -24587
rect 7664 -24155 7710 -24120
rect 7664 -24189 7670 -24155
rect 7704 -24189 7710 -24155
rect 7664 -24227 7710 -24189
rect 7664 -24261 7670 -24227
rect 7704 -24261 7710 -24227
rect 7664 -24299 7710 -24261
rect 7664 -24333 7670 -24299
rect 7704 -24333 7710 -24299
rect 7664 -24371 7710 -24333
rect 7664 -24405 7670 -24371
rect 7704 -24405 7710 -24371
rect 7664 -24443 7710 -24405
rect 7664 -24477 7670 -24443
rect 7704 -24477 7710 -24443
rect 7664 -24515 7710 -24477
rect 7664 -24549 7670 -24515
rect 7704 -24549 7710 -24515
rect 7664 -24587 7710 -24549
rect 7664 -24598 7670 -24587
rect 6646 -24652 6692 -24621
rect 7654 -24621 7670 -24598
rect 7704 -24598 7710 -24587
rect 8682 -24155 8728 -24117
rect 9686 -24117 9706 -24083
rect 9740 -24104 9752 -24083
rect 10712 -24083 10772 -23926
rect 11068 -23974 11128 -23716
rect 11210 -23762 11270 -23496
rect 11590 -23548 11650 -23538
rect 11590 -23600 11594 -23548
rect 11646 -23600 11650 -23548
rect 11204 -23766 11276 -23762
rect 11204 -23818 11214 -23766
rect 11266 -23818 11276 -23766
rect 11204 -23822 11276 -23818
rect 11590 -23774 11650 -23600
rect 11728 -23654 11788 -23406
rect 12748 -23387 12760 -23356
rect 12794 -23356 12800 -23353
rect 13764 -23353 13824 -23352
rect 12794 -23387 12808 -23356
rect 12024 -23456 12512 -23450
rect 12024 -23490 12071 -23456
rect 12105 -23490 12143 -23456
rect 12177 -23490 12215 -23456
rect 12249 -23490 12287 -23456
rect 12321 -23490 12359 -23456
rect 12393 -23490 12431 -23456
rect 12465 -23490 12512 -23456
rect 12024 -23496 12512 -23490
rect 11722 -23658 11794 -23654
rect 11722 -23710 11732 -23658
rect 11784 -23710 11794 -23658
rect 11722 -23714 11794 -23710
rect 12230 -23762 12290 -23496
rect 12350 -23662 12422 -23658
rect 12350 -23714 12360 -23662
rect 12412 -23714 12422 -23662
rect 12350 -23718 12422 -23714
rect 12224 -23766 12296 -23762
rect 11590 -23834 11790 -23774
rect 12224 -23818 12234 -23766
rect 12286 -23818 12296 -23766
rect 12224 -23822 12296 -23818
rect 11006 -23980 11494 -23974
rect 11006 -24014 11053 -23980
rect 11087 -24014 11125 -23980
rect 11159 -24014 11197 -23980
rect 11231 -24014 11269 -23980
rect 11303 -24014 11341 -23980
rect 11375 -24014 11413 -23980
rect 11447 -24014 11494 -23980
rect 11006 -24020 11494 -24014
rect 9740 -24117 9746 -24104
rect 9686 -24130 9746 -24117
rect 10712 -24117 10724 -24083
rect 10758 -24117 10772 -24083
rect 11730 -24083 11790 -23834
rect 12356 -23974 12416 -23718
rect 12748 -23866 12808 -23387
rect 13764 -23387 13778 -23353
rect 13812 -23387 13824 -23353
rect 14790 -23353 14836 -23315
rect 15808 -22883 15814 -22849
rect 15848 -22883 15854 -22849
rect 16816 -22849 16876 -22610
rect 17326 -22644 17386 -22262
rect 17838 -22550 17898 -22153
rect 18856 -22153 18868 -22128
rect 18902 -22128 18908 -22119
rect 19880 -21649 19886 -21642
rect 19920 -21642 19930 -21615
rect 20898 -21615 20944 -21584
rect 19920 -21649 19926 -21642
rect 19880 -21687 19926 -21649
rect 19880 -21721 19886 -21687
rect 19920 -21721 19926 -21687
rect 19880 -21759 19926 -21721
rect 19880 -21793 19886 -21759
rect 19920 -21793 19926 -21759
rect 19880 -21831 19926 -21793
rect 19880 -21865 19886 -21831
rect 19920 -21865 19926 -21831
rect 19880 -21903 19926 -21865
rect 19880 -21937 19886 -21903
rect 19920 -21937 19926 -21903
rect 19880 -21975 19926 -21937
rect 19880 -22009 19886 -21975
rect 19920 -22009 19926 -21975
rect 19880 -22047 19926 -22009
rect 19880 -22081 19886 -22047
rect 19920 -22081 19926 -22047
rect 19880 -22119 19926 -22081
rect 19880 -22124 19886 -22119
rect 18902 -22153 18916 -22128
rect 18132 -22222 18620 -22216
rect 18132 -22256 18179 -22222
rect 18213 -22256 18251 -22222
rect 18285 -22256 18323 -22222
rect 18357 -22256 18395 -22222
rect 18429 -22256 18467 -22222
rect 18501 -22256 18539 -22222
rect 18573 -22256 18620 -22222
rect 18132 -22262 18620 -22256
rect 17832 -22554 17904 -22550
rect 17832 -22606 17842 -22554
rect 17894 -22606 17904 -22554
rect 17832 -22610 17904 -22606
rect 18346 -22644 18406 -22262
rect 18856 -22314 18916 -22153
rect 19872 -22153 19886 -22124
rect 19920 -22124 19926 -22119
rect 20898 -21649 20904 -21615
rect 20938 -21649 20944 -21615
rect 21908 -21615 21968 -21456
rect 22410 -21506 22470 -21398
rect 22204 -21512 22692 -21506
rect 22204 -21546 22251 -21512
rect 22285 -21546 22323 -21512
rect 22357 -21546 22395 -21512
rect 22429 -21546 22467 -21512
rect 22501 -21546 22539 -21512
rect 22573 -21546 22611 -21512
rect 22645 -21546 22692 -21512
rect 22204 -21552 22692 -21546
rect 21908 -21630 21922 -21615
rect 20898 -21687 20944 -21649
rect 20898 -21721 20904 -21687
rect 20938 -21721 20944 -21687
rect 20898 -21759 20944 -21721
rect 20898 -21793 20904 -21759
rect 20938 -21793 20944 -21759
rect 20898 -21831 20944 -21793
rect 20898 -21865 20904 -21831
rect 20938 -21865 20944 -21831
rect 20898 -21903 20944 -21865
rect 20898 -21937 20904 -21903
rect 20938 -21937 20944 -21903
rect 20898 -21975 20944 -21937
rect 20898 -22009 20904 -21975
rect 20938 -22009 20944 -21975
rect 20898 -22047 20944 -22009
rect 20898 -22081 20904 -22047
rect 20938 -22081 20944 -22047
rect 20898 -22119 20944 -22081
rect 19920 -22153 19932 -22124
rect 20898 -22128 20904 -22119
rect 19150 -22222 19638 -22216
rect 19150 -22256 19197 -22222
rect 19231 -22256 19269 -22222
rect 19303 -22256 19341 -22222
rect 19375 -22256 19413 -22222
rect 19447 -22256 19485 -22222
rect 19519 -22256 19557 -22222
rect 19591 -22256 19638 -22222
rect 19150 -22262 19638 -22256
rect 18850 -22318 18922 -22314
rect 18850 -22370 18860 -22318
rect 18912 -22370 18922 -22318
rect 18850 -22374 18922 -22370
rect 18852 -22554 18924 -22550
rect 18852 -22606 18862 -22554
rect 18914 -22606 18924 -22554
rect 18852 -22610 18924 -22606
rect 17320 -22648 17392 -22644
rect 17320 -22700 17330 -22648
rect 17382 -22700 17392 -22648
rect 17320 -22704 17392 -22700
rect 18340 -22648 18412 -22644
rect 18340 -22700 18350 -22648
rect 18402 -22700 18412 -22648
rect 18340 -22704 18412 -22700
rect 17326 -22740 17386 -22704
rect 18346 -22740 18406 -22704
rect 17114 -22746 17602 -22740
rect 17114 -22780 17161 -22746
rect 17195 -22780 17233 -22746
rect 17267 -22780 17305 -22746
rect 17339 -22780 17377 -22746
rect 17411 -22780 17449 -22746
rect 17483 -22780 17521 -22746
rect 17555 -22780 17602 -22746
rect 17114 -22786 17602 -22780
rect 18132 -22746 18620 -22740
rect 18132 -22780 18179 -22746
rect 18213 -22780 18251 -22746
rect 18285 -22780 18323 -22746
rect 18357 -22780 18395 -22746
rect 18429 -22780 18467 -22746
rect 18501 -22780 18539 -22746
rect 18573 -22780 18620 -22746
rect 18132 -22786 18620 -22780
rect 16816 -22874 16832 -22849
rect 15808 -22921 15854 -22883
rect 15808 -22955 15814 -22921
rect 15848 -22955 15854 -22921
rect 15808 -22993 15854 -22955
rect 15808 -23027 15814 -22993
rect 15848 -23027 15854 -22993
rect 15808 -23065 15854 -23027
rect 15808 -23099 15814 -23065
rect 15848 -23099 15854 -23065
rect 15808 -23137 15854 -23099
rect 15808 -23171 15814 -23137
rect 15848 -23171 15854 -23137
rect 15808 -23209 15854 -23171
rect 15808 -23243 15814 -23209
rect 15848 -23243 15854 -23209
rect 15808 -23281 15854 -23243
rect 15808 -23315 15814 -23281
rect 15848 -23315 15854 -23281
rect 15808 -23346 15854 -23315
rect 16826 -22883 16832 -22874
rect 16866 -22874 16876 -22849
rect 17844 -22849 17890 -22818
rect 16866 -22883 16872 -22874
rect 16826 -22921 16872 -22883
rect 16826 -22955 16832 -22921
rect 16866 -22955 16872 -22921
rect 16826 -22993 16872 -22955
rect 16826 -23027 16832 -22993
rect 16866 -23027 16872 -22993
rect 16826 -23065 16872 -23027
rect 16826 -23099 16832 -23065
rect 16866 -23099 16872 -23065
rect 16826 -23137 16872 -23099
rect 16826 -23171 16832 -23137
rect 16866 -23171 16872 -23137
rect 16826 -23209 16872 -23171
rect 16826 -23243 16832 -23209
rect 16866 -23243 16872 -23209
rect 16826 -23281 16872 -23243
rect 16826 -23315 16832 -23281
rect 16866 -23315 16872 -23281
rect 14790 -23368 14796 -23353
rect 13042 -23456 13530 -23450
rect 13042 -23490 13089 -23456
rect 13123 -23490 13161 -23456
rect 13195 -23490 13233 -23456
rect 13267 -23490 13305 -23456
rect 13339 -23490 13377 -23456
rect 13411 -23490 13449 -23456
rect 13483 -23490 13530 -23456
rect 13042 -23496 13530 -23490
rect 13252 -23762 13312 -23496
rect 13396 -23662 13468 -23658
rect 13396 -23714 13406 -23662
rect 13458 -23714 13468 -23662
rect 13396 -23718 13468 -23714
rect 13246 -23766 13318 -23762
rect 13246 -23818 13256 -23766
rect 13308 -23818 13318 -23766
rect 13246 -23822 13318 -23818
rect 12742 -23870 12814 -23866
rect 12742 -23922 12752 -23870
rect 12804 -23922 12814 -23870
rect 12742 -23926 12814 -23922
rect 12024 -23980 12512 -23974
rect 12024 -24014 12071 -23980
rect 12105 -24014 12143 -23980
rect 12177 -24014 12215 -23980
rect 12249 -24014 12287 -23980
rect 12321 -24014 12359 -23980
rect 12393 -24014 12431 -23980
rect 12465 -24014 12512 -23980
rect 12024 -24020 12512 -24014
rect 11730 -24092 11742 -24083
rect 10712 -24124 10772 -24117
rect 11736 -24117 11742 -24092
rect 11776 -24092 11790 -24083
rect 12748 -24083 12808 -23926
rect 13402 -23974 13462 -23718
rect 13764 -23762 13824 -23387
rect 14784 -23387 14796 -23368
rect 14830 -23368 14836 -23353
rect 15800 -23353 15860 -23346
rect 16826 -23352 16872 -23315
rect 17844 -22883 17850 -22849
rect 17884 -22883 17890 -22849
rect 17844 -22921 17890 -22883
rect 18858 -22849 18918 -22610
rect 19360 -22644 19420 -22262
rect 19872 -22550 19932 -22153
rect 20888 -22153 20904 -22128
rect 20938 -22128 20944 -22119
rect 21916 -21649 21922 -21630
rect 21956 -21630 21968 -21615
rect 22926 -21615 22986 -21398
rect 21956 -21649 21962 -21630
rect 22926 -21634 22940 -21615
rect 21916 -21687 21962 -21649
rect 21916 -21721 21922 -21687
rect 21956 -21721 21962 -21687
rect 21916 -21759 21962 -21721
rect 21916 -21793 21922 -21759
rect 21956 -21793 21962 -21759
rect 21916 -21831 21962 -21793
rect 21916 -21865 21922 -21831
rect 21956 -21865 21962 -21831
rect 21916 -21903 21962 -21865
rect 21916 -21937 21922 -21903
rect 21956 -21937 21962 -21903
rect 21916 -21975 21962 -21937
rect 21916 -22009 21922 -21975
rect 21956 -22009 21962 -21975
rect 21916 -22047 21962 -22009
rect 21916 -22081 21922 -22047
rect 21956 -22081 21962 -22047
rect 21916 -22119 21962 -22081
rect 20938 -22153 20948 -22128
rect 20168 -22222 20656 -22216
rect 20168 -22256 20215 -22222
rect 20249 -22256 20287 -22222
rect 20321 -22256 20359 -22222
rect 20393 -22256 20431 -22222
rect 20465 -22256 20503 -22222
rect 20537 -22256 20575 -22222
rect 20609 -22256 20656 -22222
rect 20168 -22262 20656 -22256
rect 19866 -22554 19938 -22550
rect 19866 -22606 19876 -22554
rect 19928 -22606 19938 -22554
rect 19866 -22610 19938 -22606
rect 20396 -22644 20456 -22262
rect 20888 -22314 20948 -22153
rect 21916 -22153 21922 -22119
rect 21956 -22153 21962 -22119
rect 21916 -22184 21962 -22153
rect 22934 -21649 22940 -21634
rect 22974 -21634 22986 -21615
rect 22974 -21649 22980 -21634
rect 22934 -21687 22980 -21649
rect 22934 -21721 22940 -21687
rect 22974 -21721 22980 -21687
rect 22934 -21759 22980 -21721
rect 22934 -21793 22940 -21759
rect 22974 -21793 22980 -21759
rect 22934 -21831 22980 -21793
rect 22934 -21865 22940 -21831
rect 22974 -21865 22980 -21831
rect 22934 -21903 22980 -21865
rect 22934 -21937 22940 -21903
rect 22974 -21937 22980 -21903
rect 22934 -21975 22980 -21937
rect 22934 -22009 22940 -21975
rect 22974 -22009 22980 -21975
rect 22934 -22047 22980 -22009
rect 22934 -22081 22940 -22047
rect 22974 -22081 22980 -22047
rect 22934 -22119 22980 -22081
rect 22934 -22153 22940 -22119
rect 22974 -22153 22980 -22119
rect 22934 -22184 22980 -22153
rect 21186 -22222 21674 -22216
rect 21186 -22256 21233 -22222
rect 21267 -22256 21305 -22222
rect 21339 -22256 21521 -22222
rect 21555 -22256 21593 -22222
rect 21627 -22256 21674 -22222
rect 21186 -22262 21674 -22256
rect 22204 -22222 22692 -22216
rect 22204 -22256 22251 -22222
rect 22285 -22256 22323 -22222
rect 22357 -22256 22395 -22222
rect 22429 -22256 22467 -22222
rect 22501 -22256 22539 -22222
rect 22573 -22256 22611 -22222
rect 22645 -22256 22692 -22222
rect 22204 -22262 22692 -22256
rect 20882 -22318 20954 -22314
rect 20882 -22370 20892 -22318
rect 20944 -22370 20954 -22318
rect 20882 -22374 20954 -22370
rect 21408 -22424 21468 -22262
rect 23034 -22314 23094 -16524
rect 23156 -17382 23228 -17378
rect 23156 -17434 23166 -17382
rect 23218 -17434 23228 -17382
rect 23156 -17438 23228 -17434
rect 23162 -18936 23222 -17438
rect 23278 -17702 23338 -16410
rect 23394 -17604 23466 -17600
rect 23394 -17656 23404 -17604
rect 23456 -17656 23466 -17604
rect 23394 -17660 23466 -17656
rect 23272 -17706 23344 -17702
rect 23272 -17758 23282 -17706
rect 23334 -17758 23344 -17706
rect 23272 -17762 23344 -17758
rect 23156 -18940 23228 -18936
rect 23156 -18992 23166 -18940
rect 23218 -18992 23228 -18940
rect 23156 -18996 23228 -18992
rect 23152 -19842 23224 -19838
rect 23152 -19894 23162 -19842
rect 23214 -19894 23224 -19842
rect 23152 -19898 23224 -19894
rect 23158 -21162 23218 -19898
rect 23278 -21064 23338 -17762
rect 23272 -21068 23344 -21064
rect 23272 -21120 23282 -21068
rect 23334 -21120 23344 -21068
rect 23272 -21124 23344 -21120
rect 23152 -21166 23224 -21162
rect 23152 -21218 23162 -21166
rect 23214 -21218 23224 -21166
rect 23152 -21222 23224 -21218
rect 23400 -21396 23460 -17660
rect 23528 -18828 23588 -16306
rect 23526 -18838 23588 -18828
rect 23526 -18890 23530 -18838
rect 23582 -18890 23588 -18838
rect 23526 -18900 23588 -18890
rect 23528 -21268 23588 -18900
rect 23522 -21272 23594 -21268
rect 23522 -21324 23532 -21272
rect 23584 -21324 23594 -21272
rect 23522 -21328 23594 -21324
rect 23394 -21400 23466 -21396
rect 23394 -21452 23404 -21400
rect 23456 -21452 23466 -21400
rect 23394 -21456 23466 -21452
rect 23028 -22318 23100 -22314
rect 23028 -22370 23038 -22318
rect 23090 -22370 23100 -22318
rect 23028 -22374 23100 -22370
rect 21402 -22428 21474 -22424
rect 21402 -22480 21412 -22428
rect 21464 -22480 21474 -22428
rect 21402 -22484 21474 -22480
rect 21408 -22548 21468 -22484
rect 20888 -22554 20960 -22550
rect 20888 -22606 20898 -22554
rect 20950 -22606 20960 -22554
rect 20888 -22610 20960 -22606
rect 21408 -22608 23154 -22548
rect 19354 -22648 19426 -22644
rect 19354 -22700 19364 -22648
rect 19416 -22700 19426 -22648
rect 19354 -22704 19426 -22700
rect 20390 -22648 20462 -22644
rect 20390 -22700 20400 -22648
rect 20452 -22700 20462 -22648
rect 20390 -22704 20462 -22700
rect 19360 -22740 19420 -22704
rect 19150 -22746 19420 -22740
rect 19428 -22746 19638 -22740
rect 19150 -22780 19197 -22746
rect 19231 -22780 19269 -22746
rect 19303 -22780 19341 -22746
rect 19375 -22780 19413 -22746
rect 19447 -22780 19485 -22746
rect 19519 -22780 19557 -22746
rect 19591 -22780 19638 -22746
rect 19150 -22786 19638 -22780
rect 20168 -22746 20656 -22740
rect 20168 -22780 20215 -22746
rect 20249 -22780 20287 -22746
rect 20321 -22780 20359 -22746
rect 20393 -22780 20431 -22746
rect 20465 -22780 20503 -22746
rect 20537 -22780 20575 -22746
rect 20609 -22780 20656 -22746
rect 20168 -22786 20656 -22780
rect 19368 -22790 19428 -22786
rect 18858 -22883 18868 -22849
rect 18902 -22883 18918 -22849
rect 18858 -22896 18918 -22883
rect 19880 -22849 19926 -22818
rect 19880 -22883 19886 -22849
rect 19920 -22883 19926 -22849
rect 17844 -22955 17850 -22921
rect 17884 -22955 17890 -22921
rect 17844 -22993 17890 -22955
rect 17844 -23027 17850 -22993
rect 17884 -23027 17890 -22993
rect 17844 -23065 17890 -23027
rect 17844 -23099 17850 -23065
rect 17884 -23099 17890 -23065
rect 17844 -23137 17890 -23099
rect 17844 -23171 17850 -23137
rect 17884 -23171 17890 -23137
rect 17844 -23209 17890 -23171
rect 17844 -23243 17850 -23209
rect 17884 -23243 17890 -23209
rect 17844 -23281 17890 -23243
rect 17844 -23315 17850 -23281
rect 17884 -23315 17890 -23281
rect 14830 -23387 14844 -23368
rect 14060 -23456 14548 -23450
rect 14060 -23490 14107 -23456
rect 14141 -23490 14179 -23456
rect 14213 -23490 14251 -23456
rect 14285 -23490 14323 -23456
rect 14357 -23490 14395 -23456
rect 14429 -23490 14467 -23456
rect 14501 -23490 14548 -23456
rect 14060 -23496 14548 -23490
rect 13950 -23546 14010 -23536
rect 13950 -23598 13954 -23546
rect 14006 -23598 14010 -23546
rect 13758 -23766 13830 -23762
rect 13758 -23818 13768 -23766
rect 13820 -23818 13830 -23766
rect 13758 -23822 13830 -23818
rect 13950 -23870 14010 -23598
rect 14270 -23762 14330 -23496
rect 14264 -23766 14336 -23762
rect 14264 -23818 14274 -23766
rect 14326 -23818 14336 -23766
rect 14264 -23822 14336 -23818
rect 13766 -23930 14010 -23870
rect 13042 -23980 13530 -23974
rect 13042 -24014 13089 -23980
rect 13123 -24014 13161 -23980
rect 13195 -24014 13233 -23980
rect 13267 -24014 13305 -23980
rect 13339 -24014 13377 -23980
rect 13411 -24014 13449 -23980
rect 13483 -24014 13530 -23980
rect 13042 -24020 13530 -24014
rect 11776 -24117 11782 -24092
rect 8682 -24189 8688 -24155
rect 8722 -24189 8728 -24155
rect 8682 -24227 8728 -24189
rect 8682 -24261 8688 -24227
rect 8722 -24261 8728 -24227
rect 8682 -24299 8728 -24261
rect 8682 -24333 8688 -24299
rect 8722 -24333 8728 -24299
rect 8682 -24371 8728 -24333
rect 8682 -24405 8688 -24371
rect 8722 -24405 8728 -24371
rect 8682 -24443 8728 -24405
rect 8682 -24477 8688 -24443
rect 8722 -24477 8728 -24443
rect 8682 -24515 8728 -24477
rect 8682 -24549 8688 -24515
rect 8722 -24549 8728 -24515
rect 8682 -24587 8728 -24549
rect 7704 -24621 7714 -24598
rect 5916 -24690 6404 -24684
rect 5916 -24724 5963 -24690
rect 5997 -24724 6035 -24690
rect 6069 -24724 6107 -24690
rect 6141 -24724 6179 -24690
rect 6213 -24724 6251 -24690
rect 6285 -24724 6323 -24690
rect 6357 -24724 6404 -24690
rect 5916 -24730 6404 -24724
rect 6934 -24690 7422 -24684
rect 6934 -24724 6981 -24690
rect 7015 -24724 7053 -24690
rect 7087 -24724 7125 -24690
rect 7159 -24724 7197 -24690
rect 7231 -24724 7269 -24690
rect 7303 -24724 7341 -24690
rect 7375 -24724 7422 -24690
rect 6934 -24730 7422 -24724
rect 7654 -24784 7714 -24621
rect 8682 -24621 8688 -24587
rect 8722 -24621 8728 -24587
rect 9700 -24155 9746 -24130
rect 9700 -24189 9706 -24155
rect 9740 -24189 9746 -24155
rect 9700 -24227 9746 -24189
rect 9700 -24261 9706 -24227
rect 9740 -24261 9746 -24227
rect 9700 -24299 9746 -24261
rect 9700 -24333 9706 -24299
rect 9740 -24333 9746 -24299
rect 9700 -24371 9746 -24333
rect 9700 -24405 9706 -24371
rect 9740 -24405 9746 -24371
rect 9700 -24443 9746 -24405
rect 9700 -24477 9706 -24443
rect 9740 -24477 9746 -24443
rect 9700 -24515 9746 -24477
rect 9700 -24549 9706 -24515
rect 9740 -24549 9746 -24515
rect 9700 -24587 9746 -24549
rect 9700 -24606 9706 -24587
rect 8682 -24652 8728 -24621
rect 9692 -24621 9706 -24606
rect 9740 -24606 9746 -24587
rect 10718 -24155 10764 -24124
rect 10718 -24189 10724 -24155
rect 10758 -24189 10764 -24155
rect 10718 -24227 10764 -24189
rect 10718 -24261 10724 -24227
rect 10758 -24261 10764 -24227
rect 10718 -24299 10764 -24261
rect 10718 -24333 10724 -24299
rect 10758 -24333 10764 -24299
rect 10718 -24371 10764 -24333
rect 10718 -24405 10724 -24371
rect 10758 -24405 10764 -24371
rect 10718 -24443 10764 -24405
rect 10718 -24477 10724 -24443
rect 10758 -24477 10764 -24443
rect 10718 -24515 10764 -24477
rect 10718 -24549 10724 -24515
rect 10758 -24549 10764 -24515
rect 10718 -24587 10764 -24549
rect 9740 -24621 9752 -24606
rect 7952 -24690 8440 -24684
rect 7952 -24724 7999 -24690
rect 8033 -24724 8071 -24690
rect 8105 -24724 8143 -24690
rect 8177 -24724 8215 -24690
rect 8249 -24724 8287 -24690
rect 8321 -24724 8359 -24690
rect 8393 -24724 8440 -24690
rect 7952 -24730 8440 -24724
rect 8970 -24690 9458 -24684
rect 8970 -24724 9017 -24690
rect 9051 -24724 9089 -24690
rect 9123 -24724 9161 -24690
rect 9195 -24724 9233 -24690
rect 9267 -24724 9305 -24690
rect 9339 -24724 9377 -24690
rect 9411 -24724 9458 -24690
rect 8970 -24730 9458 -24724
rect 8158 -24784 8218 -24730
rect 7654 -24844 8218 -24784
rect 9174 -24792 9234 -24730
rect 9692 -24792 9752 -24621
rect 10718 -24621 10724 -24587
rect 10758 -24621 10764 -24587
rect 11736 -24155 11782 -24117
rect 12748 -24117 12760 -24083
rect 12794 -24117 12808 -24083
rect 13766 -24083 13826 -23930
rect 14270 -23974 14330 -23822
rect 14784 -23866 14844 -23387
rect 15800 -23387 15814 -23353
rect 15848 -23387 15860 -23353
rect 15078 -23456 15566 -23450
rect 15078 -23490 15125 -23456
rect 15159 -23490 15197 -23456
rect 15231 -23490 15269 -23456
rect 15303 -23490 15341 -23456
rect 15375 -23490 15413 -23456
rect 15447 -23490 15485 -23456
rect 15519 -23490 15566 -23456
rect 15078 -23496 15566 -23490
rect 15288 -23762 15348 -23496
rect 15800 -23544 15860 -23387
rect 16816 -23353 16876 -23352
rect 16816 -23387 16832 -23353
rect 16866 -23387 16876 -23353
rect 17844 -23353 17890 -23315
rect 17844 -23374 17850 -23353
rect 16096 -23456 16584 -23450
rect 16096 -23490 16143 -23456
rect 16177 -23490 16215 -23456
rect 16249 -23490 16287 -23456
rect 16321 -23490 16359 -23456
rect 16393 -23490 16431 -23456
rect 16465 -23490 16503 -23456
rect 16537 -23490 16584 -23456
rect 16096 -23496 16584 -23490
rect 15794 -23548 15866 -23544
rect 15794 -23600 15804 -23548
rect 15856 -23600 15866 -23548
rect 15794 -23604 15866 -23600
rect 16308 -23762 16368 -23496
rect 15282 -23766 15354 -23762
rect 15282 -23818 15292 -23766
rect 15344 -23818 15354 -23766
rect 15282 -23822 15354 -23818
rect 15794 -23766 15866 -23762
rect 15794 -23818 15804 -23766
rect 15856 -23818 15866 -23766
rect 15794 -23822 15866 -23818
rect 16302 -23766 16374 -23762
rect 16302 -23818 16312 -23766
rect 16364 -23818 16374 -23766
rect 16302 -23822 16374 -23818
rect 14778 -23870 14850 -23866
rect 14778 -23922 14788 -23870
rect 14840 -23922 14850 -23870
rect 14778 -23926 14850 -23922
rect 14060 -23980 14548 -23974
rect 14060 -24014 14107 -23980
rect 14141 -24014 14179 -23980
rect 14213 -24014 14251 -23980
rect 14285 -24014 14323 -23980
rect 14357 -24014 14395 -23980
rect 14429 -24014 14467 -23980
rect 14501 -24014 14548 -23980
rect 14060 -24020 14548 -24014
rect 13766 -24098 13778 -24083
rect 12748 -24130 12808 -24117
rect 13772 -24117 13778 -24098
rect 13812 -24098 13826 -24083
rect 14784 -24083 14844 -23926
rect 15288 -23974 15348 -23822
rect 15078 -23980 15566 -23974
rect 15078 -24014 15125 -23980
rect 15159 -24014 15197 -23980
rect 15231 -24014 15269 -23980
rect 15303 -24014 15341 -23980
rect 15375 -24014 15413 -23980
rect 15447 -24014 15485 -23980
rect 15519 -24014 15566 -23980
rect 15078 -24020 15566 -24014
rect 15800 -24064 15860 -23822
rect 16308 -23974 16368 -23822
rect 16816 -23866 16876 -23387
rect 17834 -23387 17850 -23374
rect 17884 -23374 17890 -23353
rect 18862 -22921 18908 -22896
rect 18862 -22955 18868 -22921
rect 18902 -22955 18908 -22921
rect 18862 -22993 18908 -22955
rect 18862 -23027 18868 -22993
rect 18902 -23027 18908 -22993
rect 18862 -23065 18908 -23027
rect 18862 -23099 18868 -23065
rect 18902 -23099 18908 -23065
rect 18862 -23137 18908 -23099
rect 18862 -23171 18868 -23137
rect 18902 -23171 18908 -23137
rect 18862 -23209 18908 -23171
rect 18862 -23243 18868 -23209
rect 18902 -23243 18908 -23209
rect 18862 -23281 18908 -23243
rect 18862 -23315 18868 -23281
rect 18902 -23315 18908 -23281
rect 18862 -23353 18908 -23315
rect 18862 -23358 18868 -23353
rect 17884 -23387 17894 -23374
rect 17114 -23456 17602 -23450
rect 17114 -23490 17161 -23456
rect 17195 -23490 17233 -23456
rect 17267 -23490 17305 -23456
rect 17339 -23490 17377 -23456
rect 17411 -23490 17449 -23456
rect 17483 -23490 17521 -23456
rect 17555 -23490 17602 -23456
rect 17114 -23496 17602 -23490
rect 17330 -23658 17390 -23496
rect 17834 -23544 17894 -23387
rect 18854 -23387 18868 -23358
rect 18902 -23358 18908 -23353
rect 19880 -22921 19926 -22883
rect 20894 -22849 20954 -22610
rect 21186 -22746 21674 -22740
rect 21186 -22780 21233 -22746
rect 21267 -22780 21305 -22746
rect 21339 -22780 21377 -22746
rect 21411 -22780 21449 -22746
rect 21483 -22780 21521 -22746
rect 21555 -22780 21593 -22746
rect 21627 -22780 21674 -22746
rect 21186 -22786 21674 -22780
rect 22204 -22746 22692 -22740
rect 22204 -22780 22251 -22746
rect 22285 -22780 22323 -22746
rect 22357 -22780 22395 -22746
rect 22429 -22780 22467 -22746
rect 22501 -22780 22539 -22746
rect 22573 -22780 22611 -22746
rect 22645 -22780 22692 -22746
rect 22204 -22786 22692 -22780
rect 20894 -22883 20904 -22849
rect 20938 -22883 20954 -22849
rect 20894 -22890 20954 -22883
rect 21916 -22849 21962 -22818
rect 21916 -22883 21922 -22849
rect 21956 -22883 21962 -22849
rect 19880 -22955 19886 -22921
rect 19920 -22955 19926 -22921
rect 19880 -22993 19926 -22955
rect 19880 -23027 19886 -22993
rect 19920 -23027 19926 -22993
rect 19880 -23065 19926 -23027
rect 19880 -23099 19886 -23065
rect 19920 -23099 19926 -23065
rect 19880 -23137 19926 -23099
rect 19880 -23171 19886 -23137
rect 19920 -23171 19926 -23137
rect 19880 -23209 19926 -23171
rect 19880 -23243 19886 -23209
rect 19920 -23243 19926 -23209
rect 19880 -23281 19926 -23243
rect 19880 -23315 19886 -23281
rect 19920 -23315 19926 -23281
rect 19880 -23353 19926 -23315
rect 19880 -23356 19886 -23353
rect 18902 -23387 18914 -23358
rect 18132 -23456 18620 -23450
rect 18132 -23490 18179 -23456
rect 18213 -23490 18251 -23456
rect 18285 -23490 18323 -23456
rect 18357 -23490 18395 -23456
rect 18429 -23490 18467 -23456
rect 18501 -23490 18539 -23456
rect 18573 -23490 18620 -23456
rect 18132 -23496 18620 -23490
rect 17828 -23548 17900 -23544
rect 17828 -23600 17838 -23548
rect 17890 -23600 17900 -23548
rect 17828 -23604 17900 -23600
rect 18348 -23658 18408 -23496
rect 17324 -23662 17396 -23658
rect 17324 -23714 17334 -23662
rect 17386 -23714 17396 -23662
rect 17324 -23718 17396 -23714
rect 18342 -23662 18414 -23658
rect 18342 -23714 18352 -23662
rect 18404 -23714 18414 -23662
rect 18342 -23718 18414 -23714
rect 18854 -23866 18914 -23387
rect 19868 -23387 19886 -23356
rect 19920 -23356 19926 -23353
rect 20898 -22921 20944 -22890
rect 20898 -22955 20904 -22921
rect 20938 -22955 20944 -22921
rect 20898 -22993 20944 -22955
rect 20898 -23027 20904 -22993
rect 20938 -23027 20944 -22993
rect 20898 -23065 20944 -23027
rect 20898 -23099 20904 -23065
rect 20938 -23099 20944 -23065
rect 20898 -23137 20944 -23099
rect 20898 -23171 20904 -23137
rect 20938 -23171 20944 -23137
rect 20898 -23209 20944 -23171
rect 20898 -23243 20904 -23209
rect 20938 -23243 20944 -23209
rect 20898 -23281 20944 -23243
rect 20898 -23315 20904 -23281
rect 20938 -23315 20944 -23281
rect 20898 -23353 20944 -23315
rect 19920 -23387 19928 -23356
rect 19150 -23456 19638 -23450
rect 19150 -23490 19197 -23456
rect 19231 -23490 19269 -23456
rect 19303 -23490 19341 -23456
rect 19375 -23490 19413 -23456
rect 19447 -23490 19485 -23456
rect 19519 -23490 19557 -23456
rect 19591 -23490 19638 -23456
rect 19150 -23496 19638 -23490
rect 19356 -23652 19416 -23496
rect 19868 -23544 19928 -23387
rect 20898 -23387 20904 -23353
rect 20938 -23387 20944 -23353
rect 21916 -22921 21962 -22883
rect 21916 -22955 21922 -22921
rect 21956 -22955 21962 -22921
rect 21916 -22993 21962 -22955
rect 21916 -23027 21922 -22993
rect 21956 -23027 21962 -22993
rect 21916 -23065 21962 -23027
rect 21916 -23099 21922 -23065
rect 21956 -23099 21962 -23065
rect 21916 -23137 21962 -23099
rect 21916 -23171 21922 -23137
rect 21956 -23171 21962 -23137
rect 21916 -23209 21962 -23171
rect 21916 -23243 21922 -23209
rect 21956 -23243 21962 -23209
rect 21916 -23281 21962 -23243
rect 21916 -23315 21922 -23281
rect 21956 -23315 21962 -23281
rect 21916 -23353 21962 -23315
rect 21916 -23362 21922 -23353
rect 20898 -23418 20944 -23387
rect 21910 -23387 21922 -23362
rect 21956 -23362 21962 -23353
rect 22934 -22849 22980 -22818
rect 22934 -22883 22940 -22849
rect 22974 -22883 22980 -22849
rect 22934 -22921 22980 -22883
rect 22934 -22955 22940 -22921
rect 22974 -22955 22980 -22921
rect 22934 -22993 22980 -22955
rect 22934 -23027 22940 -22993
rect 22974 -23027 22980 -22993
rect 22934 -23065 22980 -23027
rect 22934 -23099 22940 -23065
rect 22974 -23099 22980 -23065
rect 22934 -23137 22980 -23099
rect 22934 -23171 22940 -23137
rect 22974 -23171 22980 -23137
rect 22934 -23209 22980 -23171
rect 22934 -23243 22940 -23209
rect 22974 -23243 22980 -23209
rect 22934 -23281 22980 -23243
rect 22934 -23315 22940 -23281
rect 22974 -23315 22980 -23281
rect 22934 -23353 22980 -23315
rect 21956 -23387 21970 -23362
rect 22934 -23364 22940 -23353
rect 20168 -23456 20656 -23450
rect 20168 -23490 20215 -23456
rect 20249 -23490 20287 -23456
rect 20321 -23490 20359 -23456
rect 20393 -23490 20431 -23456
rect 20465 -23490 20503 -23456
rect 20537 -23490 20575 -23456
rect 20609 -23490 20656 -23456
rect 20168 -23496 20656 -23490
rect 21186 -23456 21674 -23450
rect 21186 -23490 21233 -23456
rect 21267 -23490 21305 -23456
rect 21339 -23490 21377 -23456
rect 21411 -23490 21449 -23456
rect 21483 -23490 21521 -23456
rect 21555 -23490 21593 -23456
rect 21627 -23490 21674 -23456
rect 21186 -23496 21674 -23490
rect 19862 -23548 19934 -23544
rect 19862 -23600 19872 -23548
rect 19924 -23600 19934 -23548
rect 19862 -23604 19934 -23600
rect 19356 -23662 19418 -23652
rect 19356 -23714 19362 -23662
rect 19414 -23714 19418 -23662
rect 19356 -23724 19418 -23714
rect 16810 -23870 16882 -23866
rect 16810 -23922 16820 -23870
rect 16872 -23922 16882 -23870
rect 16810 -23926 16882 -23922
rect 17332 -23870 17404 -23866
rect 17332 -23922 17342 -23870
rect 17394 -23922 17404 -23870
rect 17332 -23926 17404 -23922
rect 17832 -23870 17904 -23866
rect 17832 -23922 17842 -23870
rect 17894 -23922 17904 -23870
rect 17832 -23926 17904 -23922
rect 18340 -23870 18412 -23866
rect 18340 -23922 18350 -23870
rect 18402 -23922 18412 -23870
rect 18340 -23926 18412 -23922
rect 18848 -23870 18920 -23866
rect 18848 -23922 18858 -23870
rect 18910 -23922 18920 -23870
rect 18848 -23926 18920 -23922
rect 19198 -23870 19270 -23866
rect 19198 -23922 19208 -23870
rect 19260 -23922 19270 -23870
rect 19198 -23926 19270 -23922
rect 19356 -23868 19416 -23724
rect 20380 -23762 20440 -23496
rect 21382 -23762 21442 -23496
rect 21910 -23544 21970 -23387
rect 22928 -23387 22940 -23364
rect 22974 -23364 22980 -23353
rect 22974 -23387 22988 -23364
rect 22204 -23456 22692 -23450
rect 22204 -23490 22251 -23456
rect 22285 -23490 22323 -23456
rect 22357 -23490 22395 -23456
rect 22429 -23490 22467 -23456
rect 22501 -23490 22539 -23456
rect 22573 -23490 22611 -23456
rect 22645 -23490 22692 -23456
rect 22204 -23496 22692 -23490
rect 22422 -23544 22482 -23496
rect 22928 -23544 22988 -23387
rect 21904 -23548 21976 -23544
rect 21904 -23600 21914 -23548
rect 21966 -23600 21976 -23548
rect 21904 -23604 21976 -23600
rect 22416 -23548 22488 -23544
rect 22416 -23600 22426 -23548
rect 22478 -23600 22488 -23548
rect 22416 -23604 22488 -23600
rect 22922 -23548 22994 -23544
rect 22922 -23600 22932 -23548
rect 22984 -23600 22994 -23548
rect 22922 -23604 22994 -23600
rect 20374 -23766 20446 -23762
rect 20374 -23818 20384 -23766
rect 20436 -23818 20446 -23766
rect 20374 -23822 20446 -23818
rect 21376 -23766 21448 -23762
rect 21376 -23818 21386 -23766
rect 21438 -23818 21448 -23766
rect 21376 -23822 21448 -23818
rect 16096 -23980 16584 -23974
rect 16096 -24014 16143 -23980
rect 16177 -24014 16215 -23980
rect 16249 -24014 16287 -23980
rect 16321 -24014 16359 -23980
rect 16393 -24014 16431 -23980
rect 16465 -24014 16503 -23980
rect 16537 -24014 16584 -23980
rect 16096 -24020 16584 -24014
rect 13812 -24117 13818 -24098
rect 11736 -24189 11742 -24155
rect 11776 -24189 11782 -24155
rect 11736 -24227 11782 -24189
rect 11736 -24261 11742 -24227
rect 11776 -24261 11782 -24227
rect 11736 -24299 11782 -24261
rect 11736 -24333 11742 -24299
rect 11776 -24333 11782 -24299
rect 11736 -24371 11782 -24333
rect 11736 -24405 11742 -24371
rect 11776 -24405 11782 -24371
rect 11736 -24443 11782 -24405
rect 11736 -24477 11742 -24443
rect 11776 -24477 11782 -24443
rect 11736 -24515 11782 -24477
rect 11736 -24549 11742 -24515
rect 11776 -24549 11782 -24515
rect 11736 -24587 11782 -24549
rect 11736 -24616 11742 -24587
rect 10718 -24652 10764 -24621
rect 11730 -24621 11742 -24616
rect 11776 -24616 11782 -24587
rect 12754 -24155 12800 -24130
rect 12754 -24189 12760 -24155
rect 12794 -24189 12800 -24155
rect 12754 -24227 12800 -24189
rect 12754 -24261 12760 -24227
rect 12794 -24261 12800 -24227
rect 12754 -24299 12800 -24261
rect 12754 -24333 12760 -24299
rect 12794 -24333 12800 -24299
rect 12754 -24371 12800 -24333
rect 12754 -24405 12760 -24371
rect 12794 -24405 12800 -24371
rect 12754 -24443 12800 -24405
rect 12754 -24477 12760 -24443
rect 12794 -24477 12800 -24443
rect 12754 -24515 12800 -24477
rect 12754 -24549 12760 -24515
rect 12794 -24549 12800 -24515
rect 12754 -24587 12800 -24549
rect 13772 -24155 13818 -24117
rect 14784 -24117 14796 -24083
rect 14830 -24117 14844 -24083
rect 15796 -24083 15860 -24064
rect 15796 -24114 15814 -24083
rect 14784 -24140 14844 -24117
rect 15808 -24117 15814 -24114
rect 15848 -24112 15860 -24083
rect 16816 -24083 16876 -23926
rect 17338 -23974 17398 -23926
rect 17114 -23980 17602 -23974
rect 17114 -24014 17161 -23980
rect 17195 -24014 17233 -23980
rect 17267 -24014 17305 -23980
rect 17339 -24014 17377 -23980
rect 17411 -24014 17449 -23980
rect 17483 -24014 17521 -23980
rect 17555 -24014 17602 -23980
rect 17114 -24020 17602 -24014
rect 17338 -24026 17398 -24020
rect 17838 -24064 17898 -23926
rect 18346 -23974 18406 -23926
rect 18132 -23980 18620 -23974
rect 18132 -24014 18179 -23980
rect 18213 -24014 18251 -23980
rect 18285 -24014 18323 -23980
rect 18357 -24014 18395 -23980
rect 18429 -24014 18467 -23980
rect 18501 -24014 18539 -23980
rect 18573 -24014 18620 -23980
rect 18132 -24020 18620 -24014
rect 15848 -24114 15856 -24112
rect 15848 -24117 15854 -24114
rect 13772 -24189 13778 -24155
rect 13812 -24189 13818 -24155
rect 13772 -24227 13818 -24189
rect 13772 -24261 13778 -24227
rect 13812 -24261 13818 -24227
rect 13772 -24299 13818 -24261
rect 13772 -24333 13778 -24299
rect 13812 -24333 13818 -24299
rect 13772 -24371 13818 -24333
rect 13772 -24405 13778 -24371
rect 13812 -24405 13818 -24371
rect 13772 -24443 13818 -24405
rect 13772 -24477 13778 -24443
rect 13812 -24477 13818 -24443
rect 13772 -24515 13818 -24477
rect 13772 -24549 13778 -24515
rect 13812 -24549 13818 -24515
rect 13772 -24574 13818 -24549
rect 14790 -24155 14836 -24140
rect 14790 -24189 14796 -24155
rect 14830 -24189 14836 -24155
rect 14790 -24227 14836 -24189
rect 14790 -24261 14796 -24227
rect 14830 -24261 14836 -24227
rect 14790 -24299 14836 -24261
rect 14790 -24333 14796 -24299
rect 14830 -24333 14836 -24299
rect 14790 -24371 14836 -24333
rect 14790 -24405 14796 -24371
rect 14830 -24405 14836 -24371
rect 14790 -24443 14836 -24405
rect 14790 -24477 14796 -24443
rect 14830 -24477 14836 -24443
rect 14790 -24515 14836 -24477
rect 14790 -24549 14796 -24515
rect 14830 -24549 14836 -24515
rect 11776 -24621 11790 -24616
rect 9988 -24690 10476 -24684
rect 9988 -24724 10035 -24690
rect 10069 -24724 10107 -24690
rect 10141 -24724 10179 -24690
rect 10213 -24724 10251 -24690
rect 10285 -24724 10323 -24690
rect 10357 -24724 10395 -24690
rect 10429 -24724 10476 -24690
rect 9988 -24730 10476 -24724
rect 11006 -24690 11494 -24684
rect 11006 -24724 11053 -24690
rect 11087 -24724 11125 -24690
rect 11159 -24724 11197 -24690
rect 11231 -24724 11269 -24690
rect 11303 -24724 11341 -24690
rect 11375 -24724 11413 -24690
rect 11447 -24724 11494 -24690
rect 11006 -24730 11494 -24724
rect 10200 -24792 10260 -24730
rect 9174 -24852 10260 -24792
rect 11220 -24902 11280 -24730
rect 11730 -24798 11790 -24621
rect 12754 -24621 12760 -24587
rect 12794 -24621 12800 -24587
rect 12754 -24652 12800 -24621
rect 13766 -24587 13826 -24574
rect 13766 -24621 13778 -24587
rect 13812 -24621 13826 -24587
rect 12024 -24690 12512 -24684
rect 12024 -24724 12071 -24690
rect 12105 -24724 12143 -24690
rect 12177 -24724 12215 -24690
rect 12249 -24724 12287 -24690
rect 12321 -24724 12359 -24690
rect 12393 -24724 12431 -24690
rect 12465 -24724 12512 -24690
rect 12024 -24730 12512 -24724
rect 13042 -24690 13530 -24684
rect 13042 -24724 13089 -24690
rect 13123 -24724 13161 -24690
rect 13195 -24724 13233 -24690
rect 13267 -24724 13305 -24690
rect 13339 -24724 13377 -24690
rect 13411 -24724 13449 -24690
rect 13483 -24724 13530 -24690
rect 13042 -24730 13530 -24724
rect 11724 -24802 11796 -24798
rect 11724 -24854 11734 -24802
rect 11786 -24854 11796 -24802
rect 11724 -24858 11796 -24854
rect 12232 -24902 12292 -24730
rect 13258 -24902 13318 -24730
rect 13766 -24798 13826 -24621
rect 14790 -24587 14836 -24549
rect 14790 -24621 14796 -24587
rect 14830 -24621 14836 -24587
rect 15808 -24155 15854 -24117
rect 16816 -24117 16832 -24083
rect 16866 -24117 16876 -24083
rect 16816 -24120 16876 -24117
rect 17832 -24083 17898 -24064
rect 17832 -24117 17850 -24083
rect 17884 -24117 17898 -24083
rect 18854 -24083 18914 -23926
rect 19204 -23974 19264 -23926
rect 19356 -23928 19934 -23868
rect 19150 -23980 19638 -23974
rect 19150 -24014 19197 -23980
rect 19231 -24014 19269 -23980
rect 19303 -24014 19341 -23980
rect 19375 -24014 19413 -23980
rect 19447 -24014 19485 -23980
rect 19519 -24014 19557 -23980
rect 19591 -24014 19638 -23980
rect 19150 -24020 19638 -24014
rect 18854 -24098 18868 -24083
rect 15808 -24189 15814 -24155
rect 15848 -24189 15854 -24155
rect 15808 -24227 15854 -24189
rect 15808 -24261 15814 -24227
rect 15848 -24261 15854 -24227
rect 15808 -24299 15854 -24261
rect 15808 -24333 15814 -24299
rect 15848 -24333 15854 -24299
rect 15808 -24371 15854 -24333
rect 15808 -24405 15814 -24371
rect 15848 -24405 15854 -24371
rect 15808 -24443 15854 -24405
rect 15808 -24477 15814 -24443
rect 15848 -24477 15854 -24443
rect 15808 -24515 15854 -24477
rect 15808 -24549 15814 -24515
rect 15848 -24549 15854 -24515
rect 15808 -24587 15854 -24549
rect 15808 -24608 15814 -24587
rect 14790 -24652 14836 -24621
rect 15798 -24621 15814 -24608
rect 15848 -24608 15854 -24587
rect 16826 -24155 16872 -24120
rect 17832 -24124 17898 -24117
rect 18862 -24117 18868 -24098
rect 18902 -24098 18914 -24083
rect 19874 -24083 19934 -23928
rect 23094 -23930 23154 -22608
rect 20168 -23980 20656 -23974
rect 20168 -24014 20215 -23980
rect 20249 -24014 20287 -23980
rect 20321 -24014 20359 -23980
rect 20393 -24014 20431 -23980
rect 20465 -24014 20503 -23980
rect 20537 -24014 20575 -23980
rect 20609 -24014 20656 -23980
rect 20168 -24020 20656 -24014
rect 21186 -23980 21674 -23974
rect 21186 -24014 21233 -23980
rect 21267 -24014 21305 -23980
rect 21339 -24014 21377 -23980
rect 21411 -24014 21449 -23980
rect 21483 -24014 21521 -23980
rect 21555 -24014 21593 -23980
rect 21627 -24014 21674 -23980
rect 21186 -24020 21674 -24014
rect 22204 -23980 22692 -23974
rect 22204 -24014 22251 -23980
rect 22285 -24014 22323 -23980
rect 22357 -24014 22395 -23980
rect 22429 -24014 22467 -23980
rect 22501 -24014 22539 -23980
rect 22573 -24014 22611 -23980
rect 22645 -24014 22692 -23980
rect 22204 -24020 22692 -24014
rect 22934 -23990 23154 -23930
rect 18902 -24117 18908 -24098
rect 19874 -24102 19886 -24083
rect 16826 -24189 16832 -24155
rect 16866 -24189 16872 -24155
rect 16826 -24227 16872 -24189
rect 16826 -24261 16832 -24227
rect 16866 -24261 16872 -24227
rect 16826 -24299 16872 -24261
rect 16826 -24333 16832 -24299
rect 16866 -24333 16872 -24299
rect 16826 -24371 16872 -24333
rect 16826 -24405 16832 -24371
rect 16866 -24405 16872 -24371
rect 16826 -24443 16872 -24405
rect 16826 -24477 16832 -24443
rect 16866 -24477 16872 -24443
rect 16826 -24515 16872 -24477
rect 16826 -24549 16832 -24515
rect 16866 -24549 16872 -24515
rect 16826 -24587 16872 -24549
rect 15848 -24621 15858 -24608
rect 14060 -24690 14548 -24684
rect 14060 -24724 14107 -24690
rect 14141 -24724 14179 -24690
rect 14213 -24724 14251 -24690
rect 14285 -24724 14323 -24690
rect 14357 -24724 14395 -24690
rect 14429 -24724 14467 -24690
rect 14501 -24724 14548 -24690
rect 14060 -24730 14548 -24724
rect 15078 -24690 15566 -24684
rect 15078 -24724 15125 -24690
rect 15159 -24724 15197 -24690
rect 15231 -24724 15269 -24690
rect 15303 -24724 15341 -24690
rect 15375 -24724 15413 -24690
rect 15447 -24724 15485 -24690
rect 15519 -24724 15566 -24690
rect 15078 -24730 15566 -24724
rect 15286 -24790 15346 -24730
rect 15798 -24790 15858 -24621
rect 16826 -24621 16832 -24587
rect 16866 -24621 16872 -24587
rect 17844 -24155 17890 -24124
rect 17844 -24189 17850 -24155
rect 17884 -24189 17890 -24155
rect 17844 -24227 17890 -24189
rect 17844 -24261 17850 -24227
rect 17884 -24261 17890 -24227
rect 17844 -24299 17890 -24261
rect 17844 -24333 17850 -24299
rect 17884 -24333 17890 -24299
rect 17844 -24371 17890 -24333
rect 17844 -24405 17850 -24371
rect 17884 -24405 17890 -24371
rect 17844 -24443 17890 -24405
rect 17844 -24477 17850 -24443
rect 17884 -24477 17890 -24443
rect 17844 -24515 17890 -24477
rect 17844 -24549 17850 -24515
rect 17884 -24549 17890 -24515
rect 17844 -24587 17890 -24549
rect 17844 -24602 17850 -24587
rect 16826 -24652 16872 -24621
rect 17834 -24621 17850 -24602
rect 17884 -24602 17890 -24587
rect 18862 -24155 18908 -24117
rect 18862 -24189 18868 -24155
rect 18902 -24189 18908 -24155
rect 18862 -24227 18908 -24189
rect 18862 -24261 18868 -24227
rect 18902 -24261 18908 -24227
rect 18862 -24299 18908 -24261
rect 18862 -24333 18868 -24299
rect 18902 -24333 18908 -24299
rect 18862 -24371 18908 -24333
rect 18862 -24405 18868 -24371
rect 18902 -24405 18908 -24371
rect 18862 -24443 18908 -24405
rect 18862 -24477 18868 -24443
rect 18902 -24477 18908 -24443
rect 18862 -24515 18908 -24477
rect 18862 -24549 18868 -24515
rect 18902 -24549 18908 -24515
rect 18862 -24587 18908 -24549
rect 17884 -24621 17894 -24602
rect 17834 -24640 17894 -24621
rect 18862 -24621 18868 -24587
rect 18902 -24621 18908 -24587
rect 18862 -24652 18908 -24621
rect 19880 -24117 19886 -24102
rect 19920 -24102 19934 -24083
rect 20898 -24083 20944 -24052
rect 19920 -24117 19926 -24102
rect 19880 -24155 19926 -24117
rect 19880 -24189 19886 -24155
rect 19920 -24189 19926 -24155
rect 19880 -24227 19926 -24189
rect 19880 -24261 19886 -24227
rect 19920 -24261 19926 -24227
rect 19880 -24299 19926 -24261
rect 19880 -24333 19886 -24299
rect 19920 -24333 19926 -24299
rect 19880 -24371 19926 -24333
rect 19880 -24405 19886 -24371
rect 19920 -24405 19926 -24371
rect 19880 -24443 19926 -24405
rect 19880 -24477 19886 -24443
rect 19920 -24477 19926 -24443
rect 19880 -24515 19926 -24477
rect 19880 -24549 19886 -24515
rect 19920 -24549 19926 -24515
rect 19880 -24587 19926 -24549
rect 19880 -24621 19886 -24587
rect 19920 -24621 19926 -24587
rect 20898 -24117 20904 -24083
rect 20938 -24117 20944 -24083
rect 20898 -24155 20944 -24117
rect 20898 -24189 20904 -24155
rect 20938 -24189 20944 -24155
rect 20898 -24227 20944 -24189
rect 20898 -24261 20904 -24227
rect 20938 -24261 20944 -24227
rect 20898 -24299 20944 -24261
rect 20898 -24333 20904 -24299
rect 20938 -24333 20944 -24299
rect 20898 -24371 20944 -24333
rect 20898 -24405 20904 -24371
rect 20938 -24405 20944 -24371
rect 20898 -24443 20944 -24405
rect 20898 -24477 20904 -24443
rect 20938 -24477 20944 -24443
rect 20898 -24515 20944 -24477
rect 20898 -24549 20904 -24515
rect 20938 -24549 20944 -24515
rect 20898 -24587 20944 -24549
rect 20898 -24608 20904 -24587
rect 19880 -24652 19926 -24621
rect 20888 -24621 20904 -24608
rect 20938 -24608 20944 -24587
rect 21916 -24083 21962 -24052
rect 21916 -24117 21922 -24083
rect 21956 -24117 21962 -24083
rect 21916 -24155 21962 -24117
rect 21916 -24189 21922 -24155
rect 21956 -24189 21962 -24155
rect 21916 -24227 21962 -24189
rect 21916 -24261 21922 -24227
rect 21956 -24261 21962 -24227
rect 21916 -24299 21962 -24261
rect 21916 -24333 21922 -24299
rect 21956 -24333 21962 -24299
rect 21916 -24371 21962 -24333
rect 21916 -24405 21922 -24371
rect 21956 -24405 21962 -24371
rect 21916 -24443 21962 -24405
rect 21916 -24477 21922 -24443
rect 21956 -24477 21962 -24443
rect 21916 -24515 21962 -24477
rect 21916 -24549 21922 -24515
rect 21956 -24549 21962 -24515
rect 21916 -24587 21962 -24549
rect 21916 -24592 21922 -24587
rect 20938 -24621 20948 -24608
rect 16096 -24690 16584 -24684
rect 16096 -24724 16143 -24690
rect 16177 -24724 16215 -24690
rect 16249 -24724 16287 -24690
rect 16321 -24724 16359 -24690
rect 16393 -24724 16431 -24690
rect 16465 -24724 16503 -24690
rect 16537 -24724 16584 -24690
rect 16096 -24730 16584 -24724
rect 17114 -24690 17602 -24684
rect 17114 -24724 17161 -24690
rect 17195 -24724 17233 -24690
rect 17267 -24724 17305 -24690
rect 17339 -24724 17377 -24690
rect 17411 -24724 17449 -24690
rect 17483 -24724 17521 -24690
rect 17555 -24724 17602 -24690
rect 17114 -24730 17330 -24724
rect 17390 -24730 17602 -24724
rect 18132 -24690 18620 -24684
rect 18132 -24724 18179 -24690
rect 18213 -24724 18251 -24690
rect 18285 -24724 18323 -24690
rect 18357 -24724 18395 -24690
rect 18429 -24724 18467 -24690
rect 18501 -24724 18539 -24690
rect 18573 -24724 18620 -24690
rect 18132 -24730 18620 -24724
rect 19150 -24690 19638 -24684
rect 19150 -24724 19197 -24690
rect 19231 -24724 19269 -24690
rect 19303 -24724 19341 -24690
rect 19375 -24724 19413 -24690
rect 19447 -24724 19485 -24690
rect 19519 -24724 19557 -24690
rect 19591 -24724 19638 -24690
rect 19150 -24730 19638 -24724
rect 20168 -24690 20656 -24684
rect 20168 -24724 20215 -24690
rect 20249 -24724 20287 -24690
rect 20321 -24724 20359 -24690
rect 20393 -24724 20431 -24690
rect 20465 -24724 20503 -24690
rect 20537 -24724 20575 -24690
rect 20609 -24724 20656 -24690
rect 20168 -24730 20656 -24724
rect 16304 -24790 16364 -24730
rect 13760 -24802 13832 -24798
rect 13760 -24854 13770 -24802
rect 13822 -24854 13832 -24802
rect 15286 -24850 16364 -24790
rect 13760 -24858 13832 -24854
rect 11220 -24962 13318 -24902
rect 5612 -25002 5684 -24998
rect 5612 -25054 5622 -25002
rect 5674 -25054 5684 -25002
rect 5612 -25058 5684 -25054
rect 7650 -25002 7722 -24998
rect 7650 -25054 7660 -25002
rect 7712 -25054 7722 -25002
rect 7650 -25058 7722 -25054
rect 9682 -25002 9754 -24998
rect 9682 -25054 9692 -25002
rect 9744 -25054 9754 -25002
rect 9682 -25058 9754 -25054
rect 11720 -25002 11792 -24998
rect 11720 -25054 11730 -25002
rect 11782 -25054 11792 -25002
rect 11720 -25058 11792 -25054
rect 13754 -25002 13826 -24998
rect 13754 -25054 13764 -25002
rect 13816 -25054 13826 -25002
rect 13754 -25058 13826 -25054
rect 15794 -25002 15866 -24998
rect 15794 -25054 15804 -25002
rect 15856 -25054 15866 -25002
rect 15794 -25058 15866 -25054
rect 17828 -25002 17900 -24998
rect 17828 -25054 17838 -25002
rect 17890 -25054 17900 -25002
rect 17828 -25058 17900 -25054
rect 19862 -25002 19934 -24998
rect 19862 -25054 19872 -25002
rect 19924 -25054 19934 -25002
rect 19862 -25058 19934 -25054
rect 4898 -25212 5386 -25206
rect 4898 -25246 4945 -25212
rect 4979 -25246 5017 -25212
rect 5051 -25246 5089 -25212
rect 5123 -25246 5161 -25212
rect 5195 -25246 5233 -25212
rect 5267 -25246 5305 -25212
rect 5339 -25246 5386 -25212
rect 4898 -25252 5386 -25246
rect 3632 -25349 3638 -25334
rect 4598 -25344 4616 -25315
rect 2574 -25387 2620 -25352
rect 2574 -25421 2580 -25387
rect 2614 -25421 2620 -25387
rect 2574 -25459 2620 -25421
rect 2574 -25493 2580 -25459
rect 2614 -25493 2620 -25459
rect 2574 -25531 2620 -25493
rect 2574 -25565 2580 -25531
rect 2614 -25565 2620 -25531
rect 2574 -25603 2620 -25565
rect 2574 -25637 2580 -25603
rect 2614 -25637 2620 -25603
rect 2574 -25675 2620 -25637
rect 2574 -25709 2580 -25675
rect 2614 -25709 2620 -25675
rect 2574 -25747 2620 -25709
rect 2574 -25781 2580 -25747
rect 2614 -25781 2620 -25747
rect 2574 -25819 2620 -25781
rect 2574 -25853 2580 -25819
rect 2614 -25853 2620 -25819
rect 3592 -25387 3638 -25349
rect 3592 -25421 3598 -25387
rect 3632 -25421 3638 -25387
rect 3592 -25459 3638 -25421
rect 3592 -25493 3598 -25459
rect 3632 -25493 3638 -25459
rect 3592 -25531 3638 -25493
rect 3592 -25565 3598 -25531
rect 3632 -25565 3638 -25531
rect 3592 -25603 3638 -25565
rect 3592 -25637 3598 -25603
rect 3632 -25637 3638 -25603
rect 3592 -25675 3638 -25637
rect 3592 -25709 3598 -25675
rect 3632 -25709 3638 -25675
rect 3592 -25747 3638 -25709
rect 3592 -25781 3598 -25747
rect 3632 -25781 3638 -25747
rect 3592 -25819 3638 -25781
rect 3592 -25822 3598 -25819
rect 2574 -25884 2620 -25853
rect 3582 -25853 3598 -25822
rect 3632 -25822 3638 -25819
rect 4610 -25349 4616 -25344
rect 4650 -25344 4658 -25315
rect 5618 -25315 5678 -25058
rect 6630 -25100 6702 -25096
rect 6630 -25152 6640 -25100
rect 6692 -25152 6702 -25100
rect 6630 -25156 6702 -25152
rect 5916 -25212 6404 -25206
rect 5916 -25246 5963 -25212
rect 5997 -25246 6035 -25212
rect 6069 -25246 6107 -25212
rect 6141 -25246 6179 -25212
rect 6213 -25246 6251 -25212
rect 6285 -25246 6323 -25212
rect 6357 -25246 6404 -25212
rect 5916 -25252 6404 -25246
rect 5618 -25328 5634 -25315
rect 4650 -25349 4656 -25344
rect 4610 -25387 4656 -25349
rect 4610 -25421 4616 -25387
rect 4650 -25421 4656 -25387
rect 4610 -25459 4656 -25421
rect 4610 -25493 4616 -25459
rect 4650 -25493 4656 -25459
rect 4610 -25531 4656 -25493
rect 4610 -25565 4616 -25531
rect 4650 -25565 4656 -25531
rect 4610 -25603 4656 -25565
rect 4610 -25637 4616 -25603
rect 4650 -25637 4656 -25603
rect 4610 -25675 4656 -25637
rect 4610 -25709 4616 -25675
rect 4650 -25709 4656 -25675
rect 4610 -25747 4656 -25709
rect 4610 -25781 4616 -25747
rect 4650 -25781 4656 -25747
rect 4610 -25819 4656 -25781
rect 5628 -25349 5634 -25328
rect 5668 -25328 5678 -25315
rect 6636 -25315 6696 -25156
rect 6934 -25212 7422 -25206
rect 6934 -25246 6981 -25212
rect 7015 -25246 7053 -25212
rect 7087 -25246 7125 -25212
rect 7159 -25246 7197 -25212
rect 7231 -25246 7269 -25212
rect 7303 -25246 7341 -25212
rect 7375 -25246 7422 -25212
rect 6934 -25252 7422 -25246
rect 5668 -25349 5674 -25328
rect 5628 -25387 5674 -25349
rect 6636 -25349 6652 -25315
rect 6686 -25349 6696 -25315
rect 7656 -25315 7716 -25058
rect 8666 -25100 8738 -25096
rect 8666 -25152 8676 -25100
rect 8728 -25152 8738 -25100
rect 8666 -25156 8738 -25152
rect 7952 -25212 8440 -25206
rect 7952 -25246 7999 -25212
rect 8033 -25246 8071 -25212
rect 8105 -25246 8143 -25212
rect 8177 -25246 8215 -25212
rect 8249 -25246 8287 -25212
rect 8321 -25246 8359 -25212
rect 8393 -25246 8440 -25212
rect 7952 -25252 8440 -25246
rect 7656 -25342 7670 -25315
rect 6636 -25352 6696 -25349
rect 7664 -25349 7670 -25342
rect 7704 -25342 7716 -25315
rect 8672 -25315 8732 -25156
rect 8970 -25212 9458 -25206
rect 8970 -25246 9017 -25212
rect 9051 -25246 9089 -25212
rect 9123 -25246 9161 -25212
rect 9195 -25246 9233 -25212
rect 9267 -25246 9305 -25212
rect 9339 -25246 9377 -25212
rect 9411 -25246 9458 -25212
rect 8970 -25252 9458 -25246
rect 7704 -25349 7710 -25342
rect 8672 -25346 8688 -25315
rect 5628 -25421 5634 -25387
rect 5668 -25421 5674 -25387
rect 5628 -25459 5674 -25421
rect 5628 -25493 5634 -25459
rect 5668 -25493 5674 -25459
rect 5628 -25531 5674 -25493
rect 5628 -25565 5634 -25531
rect 5668 -25565 5674 -25531
rect 5628 -25603 5674 -25565
rect 5628 -25637 5634 -25603
rect 5668 -25637 5674 -25603
rect 5628 -25675 5674 -25637
rect 5628 -25709 5634 -25675
rect 5668 -25709 5674 -25675
rect 5628 -25747 5674 -25709
rect 5628 -25781 5634 -25747
rect 5668 -25781 5674 -25747
rect 5628 -25782 5674 -25781
rect 6646 -25387 6692 -25352
rect 6646 -25421 6652 -25387
rect 6686 -25421 6692 -25387
rect 6646 -25459 6692 -25421
rect 6646 -25493 6652 -25459
rect 6686 -25493 6692 -25459
rect 6646 -25531 6692 -25493
rect 6646 -25565 6652 -25531
rect 6686 -25565 6692 -25531
rect 6646 -25603 6692 -25565
rect 6646 -25637 6652 -25603
rect 6686 -25637 6692 -25603
rect 6646 -25675 6692 -25637
rect 6646 -25709 6652 -25675
rect 6686 -25709 6692 -25675
rect 6646 -25747 6692 -25709
rect 6646 -25781 6652 -25747
rect 6686 -25781 6692 -25747
rect 3632 -25853 3642 -25822
rect 2862 -25922 3350 -25916
rect 2862 -25956 2909 -25922
rect 2943 -25956 2981 -25922
rect 3015 -25956 3053 -25922
rect 3087 -25956 3125 -25922
rect 3159 -25956 3197 -25922
rect 3231 -25956 3269 -25922
rect 3303 -25956 3350 -25922
rect 2862 -25962 3350 -25956
rect 3066 -26028 3126 -25962
rect 3582 -26028 3642 -25853
rect 4610 -25853 4616 -25819
rect 4650 -25853 4656 -25819
rect 5634 -25819 5668 -25782
rect 4610 -25884 4656 -25853
rect 5620 -25853 5634 -25844
rect 6646 -25819 6692 -25781
rect 5668 -25853 5680 -25844
rect 3880 -25922 4368 -25916
rect 3880 -25956 3927 -25922
rect 3961 -25956 3999 -25922
rect 4033 -25956 4071 -25922
rect 4105 -25956 4143 -25922
rect 4177 -25956 4215 -25922
rect 4249 -25956 4287 -25922
rect 4321 -25956 4368 -25922
rect 3880 -25962 4368 -25956
rect 4898 -25922 5386 -25916
rect 4898 -25956 4945 -25922
rect 4979 -25956 5017 -25922
rect 5051 -25956 5089 -25922
rect 5123 -25956 5161 -25922
rect 5195 -25956 5233 -25922
rect 5267 -25956 5305 -25922
rect 5339 -25956 5386 -25922
rect 4898 -25962 5386 -25956
rect 4114 -26028 4174 -25962
rect 5104 -26028 5164 -25962
rect 5620 -26028 5680 -25853
rect 6646 -25853 6652 -25819
rect 6686 -25853 6692 -25819
rect 7664 -25387 7710 -25349
rect 7664 -25421 7670 -25387
rect 7704 -25421 7710 -25387
rect 7664 -25459 7710 -25421
rect 7664 -25493 7670 -25459
rect 7704 -25493 7710 -25459
rect 7664 -25531 7710 -25493
rect 7664 -25565 7670 -25531
rect 7704 -25565 7710 -25531
rect 7664 -25603 7710 -25565
rect 7664 -25637 7670 -25603
rect 7704 -25637 7710 -25603
rect 7664 -25675 7710 -25637
rect 7664 -25709 7670 -25675
rect 7704 -25709 7710 -25675
rect 7664 -25747 7710 -25709
rect 7664 -25781 7670 -25747
rect 7704 -25781 7710 -25747
rect 7664 -25819 7710 -25781
rect 7664 -25844 7670 -25819
rect 6646 -25884 6692 -25853
rect 7656 -25853 7670 -25844
rect 7704 -25844 7710 -25819
rect 8682 -25349 8688 -25346
rect 8722 -25346 8732 -25315
rect 9688 -25315 9748 -25058
rect 10702 -25100 10774 -25096
rect 10702 -25152 10712 -25100
rect 10764 -25152 10774 -25100
rect 10702 -25156 10774 -25152
rect 9988 -25212 10476 -25206
rect 9988 -25246 10035 -25212
rect 10069 -25246 10107 -25212
rect 10141 -25246 10179 -25212
rect 10213 -25246 10251 -25212
rect 10285 -25246 10323 -25212
rect 10357 -25246 10395 -25212
rect 10429 -25246 10476 -25212
rect 9988 -25252 10476 -25246
rect 8722 -25349 8728 -25346
rect 8682 -25387 8728 -25349
rect 9688 -25349 9706 -25315
rect 9740 -25349 9748 -25315
rect 10708 -25315 10768 -25156
rect 11006 -25212 11494 -25206
rect 11006 -25246 11053 -25212
rect 11087 -25246 11125 -25212
rect 11159 -25246 11197 -25212
rect 11231 -25246 11269 -25212
rect 11303 -25246 11341 -25212
rect 11375 -25246 11413 -25212
rect 11447 -25246 11494 -25212
rect 11006 -25252 11494 -25246
rect 10708 -25344 10724 -25315
rect 9688 -25352 9748 -25349
rect 10718 -25349 10724 -25344
rect 10758 -25344 10768 -25315
rect 11726 -25315 11786 -25058
rect 12738 -25100 12810 -25096
rect 12738 -25152 12748 -25100
rect 12800 -25152 12810 -25100
rect 12738 -25156 12810 -25152
rect 12024 -25212 12512 -25206
rect 12024 -25246 12071 -25212
rect 12105 -25246 12143 -25212
rect 12177 -25246 12215 -25212
rect 12249 -25246 12287 -25212
rect 12321 -25246 12359 -25212
rect 12393 -25246 12431 -25212
rect 12465 -25246 12512 -25212
rect 12024 -25252 12512 -25246
rect 11726 -25340 11742 -25315
rect 10758 -25349 10764 -25344
rect 8682 -25421 8688 -25387
rect 8722 -25421 8728 -25387
rect 8682 -25459 8728 -25421
rect 8682 -25493 8688 -25459
rect 8722 -25493 8728 -25459
rect 8682 -25531 8728 -25493
rect 8682 -25565 8688 -25531
rect 8722 -25565 8728 -25531
rect 8682 -25603 8728 -25565
rect 8682 -25637 8688 -25603
rect 8722 -25637 8728 -25603
rect 8682 -25675 8728 -25637
rect 8682 -25709 8688 -25675
rect 8722 -25709 8728 -25675
rect 8682 -25747 8728 -25709
rect 8682 -25781 8688 -25747
rect 8722 -25781 8728 -25747
rect 8682 -25819 8728 -25781
rect 7704 -25853 7716 -25844
rect 5916 -25922 6404 -25916
rect 5916 -25956 5963 -25922
rect 5997 -25956 6035 -25922
rect 6069 -25956 6107 -25922
rect 6141 -25956 6179 -25922
rect 6213 -25956 6251 -25922
rect 6285 -25956 6323 -25922
rect 6357 -25956 6404 -25922
rect 5916 -25962 6404 -25956
rect 6934 -25922 7422 -25916
rect 6934 -25956 6981 -25922
rect 7015 -25956 7053 -25922
rect 7087 -25956 7125 -25922
rect 7159 -25956 7197 -25922
rect 7231 -25956 7269 -25922
rect 7303 -25956 7341 -25922
rect 7375 -25956 7422 -25922
rect 6934 -25962 7422 -25956
rect 6126 -26028 6186 -25962
rect 7148 -26028 7208 -25962
rect 7656 -26028 7716 -25853
rect 8682 -25853 8688 -25819
rect 8722 -25853 8728 -25819
rect 9700 -25387 9746 -25352
rect 9700 -25421 9706 -25387
rect 9740 -25421 9746 -25387
rect 9700 -25459 9746 -25421
rect 9700 -25493 9706 -25459
rect 9740 -25493 9746 -25459
rect 9700 -25531 9746 -25493
rect 9700 -25565 9706 -25531
rect 9740 -25565 9746 -25531
rect 9700 -25603 9746 -25565
rect 9700 -25637 9706 -25603
rect 9740 -25637 9746 -25603
rect 9700 -25675 9746 -25637
rect 9700 -25709 9706 -25675
rect 9740 -25709 9746 -25675
rect 9700 -25747 9746 -25709
rect 9700 -25781 9706 -25747
rect 9740 -25781 9746 -25747
rect 9700 -25819 9746 -25781
rect 9700 -25838 9706 -25819
rect 8682 -25884 8728 -25853
rect 9690 -25853 9706 -25838
rect 9740 -25838 9746 -25819
rect 10718 -25387 10764 -25349
rect 10718 -25421 10724 -25387
rect 10758 -25421 10764 -25387
rect 10718 -25459 10764 -25421
rect 10718 -25493 10724 -25459
rect 10758 -25493 10764 -25459
rect 10718 -25531 10764 -25493
rect 10718 -25565 10724 -25531
rect 10758 -25565 10764 -25531
rect 10718 -25603 10764 -25565
rect 10718 -25637 10724 -25603
rect 10758 -25637 10764 -25603
rect 10718 -25675 10764 -25637
rect 10718 -25709 10724 -25675
rect 10758 -25709 10764 -25675
rect 10718 -25747 10764 -25709
rect 10718 -25781 10724 -25747
rect 10758 -25781 10764 -25747
rect 10718 -25819 10764 -25781
rect 11736 -25349 11742 -25340
rect 11776 -25340 11786 -25315
rect 12744 -25315 12804 -25156
rect 13042 -25212 13530 -25206
rect 13042 -25246 13089 -25212
rect 13123 -25246 13161 -25212
rect 13195 -25246 13233 -25212
rect 13267 -25246 13305 -25212
rect 13339 -25246 13377 -25212
rect 13411 -25246 13449 -25212
rect 13483 -25246 13530 -25212
rect 13042 -25252 13530 -25246
rect 12744 -25338 12760 -25315
rect 11776 -25349 11782 -25340
rect 11736 -25387 11782 -25349
rect 11736 -25421 11742 -25387
rect 11776 -25421 11782 -25387
rect 11736 -25459 11782 -25421
rect 11736 -25493 11742 -25459
rect 11776 -25493 11782 -25459
rect 11736 -25531 11782 -25493
rect 11736 -25565 11742 -25531
rect 11776 -25565 11782 -25531
rect 11736 -25603 11782 -25565
rect 11736 -25637 11742 -25603
rect 11776 -25637 11782 -25603
rect 11736 -25675 11782 -25637
rect 11736 -25709 11742 -25675
rect 11776 -25709 11782 -25675
rect 11736 -25747 11782 -25709
rect 11736 -25781 11742 -25747
rect 11776 -25781 11782 -25747
rect 11736 -25814 11782 -25781
rect 12754 -25349 12760 -25338
rect 12794 -25338 12804 -25315
rect 13760 -25315 13820 -25058
rect 14772 -25100 14844 -25096
rect 14772 -25152 14782 -25100
rect 14834 -25152 14844 -25100
rect 14772 -25156 14844 -25152
rect 14060 -25212 14548 -25206
rect 14060 -25246 14107 -25212
rect 14141 -25246 14179 -25212
rect 14213 -25246 14251 -25212
rect 14285 -25246 14323 -25212
rect 14357 -25246 14395 -25212
rect 14429 -25246 14467 -25212
rect 14501 -25246 14548 -25212
rect 14060 -25252 14548 -25246
rect 12794 -25349 12800 -25338
rect 12754 -25387 12800 -25349
rect 13760 -25349 13778 -25315
rect 13812 -25349 13820 -25315
rect 14778 -25315 14838 -25156
rect 15078 -25212 15566 -25206
rect 15078 -25246 15125 -25212
rect 15159 -25246 15197 -25212
rect 15231 -25246 15269 -25212
rect 15303 -25246 15341 -25212
rect 15375 -25246 15413 -25212
rect 15447 -25246 15485 -25212
rect 15519 -25246 15566 -25212
rect 15078 -25252 15566 -25246
rect 14778 -25338 14796 -25315
rect 13760 -25352 13820 -25349
rect 14790 -25349 14796 -25338
rect 14830 -25338 14838 -25315
rect 15800 -25315 15860 -25058
rect 16808 -25100 16880 -25096
rect 16808 -25152 16818 -25100
rect 16870 -25152 16880 -25100
rect 16808 -25156 16880 -25152
rect 16096 -25212 16584 -25206
rect 16096 -25246 16143 -25212
rect 16177 -25246 16215 -25212
rect 16249 -25246 16287 -25212
rect 16321 -25246 16359 -25212
rect 16393 -25246 16431 -25212
rect 16465 -25246 16503 -25212
rect 16537 -25246 16584 -25212
rect 16096 -25252 16584 -25246
rect 14830 -25349 14836 -25338
rect 15800 -25342 15814 -25315
rect 12754 -25421 12760 -25387
rect 12794 -25421 12800 -25387
rect 12754 -25459 12800 -25421
rect 12754 -25493 12760 -25459
rect 12794 -25493 12800 -25459
rect 12754 -25531 12800 -25493
rect 12754 -25565 12760 -25531
rect 12794 -25565 12800 -25531
rect 12754 -25603 12800 -25565
rect 12754 -25637 12760 -25603
rect 12794 -25637 12800 -25603
rect 12754 -25675 12800 -25637
rect 12754 -25709 12760 -25675
rect 12794 -25709 12800 -25675
rect 12754 -25747 12800 -25709
rect 12754 -25781 12760 -25747
rect 12794 -25781 12800 -25747
rect 9740 -25853 9750 -25838
rect 7952 -25922 8440 -25916
rect 7952 -25956 7999 -25922
rect 8033 -25956 8071 -25922
rect 8105 -25956 8143 -25922
rect 8177 -25956 8215 -25922
rect 8249 -25956 8287 -25922
rect 8321 -25956 8359 -25922
rect 8393 -25956 8440 -25922
rect 7952 -25962 8440 -25956
rect 8970 -25922 9458 -25916
rect 8970 -25956 9017 -25922
rect 9051 -25956 9089 -25922
rect 9123 -25956 9161 -25922
rect 9195 -25956 9233 -25922
rect 9267 -25956 9305 -25922
rect 9339 -25956 9377 -25922
rect 9411 -25956 9458 -25922
rect 8970 -25962 9458 -25956
rect 8170 -26028 8230 -25962
rect 9180 -26028 9240 -25962
rect 9690 -26028 9750 -25853
rect 10718 -25853 10724 -25819
rect 10758 -25853 10764 -25819
rect 10718 -25884 10764 -25853
rect 11730 -25819 11790 -25814
rect 11730 -25853 11742 -25819
rect 11776 -25853 11790 -25819
rect 9988 -25922 10476 -25916
rect 9988 -25956 10035 -25922
rect 10069 -25956 10107 -25922
rect 10141 -25956 10179 -25922
rect 10213 -25956 10251 -25922
rect 10285 -25956 10323 -25922
rect 10357 -25956 10395 -25922
rect 10429 -25956 10476 -25922
rect 9988 -25962 10476 -25956
rect 11006 -25922 11494 -25916
rect 11006 -25956 11053 -25922
rect 11087 -25956 11125 -25922
rect 11159 -25956 11197 -25922
rect 11231 -25956 11269 -25922
rect 11303 -25956 11341 -25922
rect 11375 -25956 11413 -25922
rect 11447 -25956 11494 -25922
rect 11006 -25962 11494 -25956
rect 10208 -26028 10268 -25962
rect 11226 -26028 11286 -25962
rect 11730 -26028 11790 -25853
rect 12754 -25819 12800 -25781
rect 12754 -25853 12760 -25819
rect 12794 -25853 12800 -25819
rect 13772 -25387 13818 -25352
rect 13772 -25421 13778 -25387
rect 13812 -25421 13818 -25387
rect 13772 -25459 13818 -25421
rect 13772 -25493 13778 -25459
rect 13812 -25493 13818 -25459
rect 13772 -25531 13818 -25493
rect 13772 -25565 13778 -25531
rect 13812 -25565 13818 -25531
rect 13772 -25603 13818 -25565
rect 13772 -25637 13778 -25603
rect 13812 -25637 13818 -25603
rect 13772 -25675 13818 -25637
rect 13772 -25709 13778 -25675
rect 13812 -25709 13818 -25675
rect 13772 -25747 13818 -25709
rect 13772 -25781 13778 -25747
rect 13812 -25781 13818 -25747
rect 13772 -25819 13818 -25781
rect 13772 -25842 13778 -25819
rect 12754 -25884 12800 -25853
rect 13768 -25853 13778 -25842
rect 13812 -25842 13818 -25819
rect 14790 -25387 14836 -25349
rect 14790 -25421 14796 -25387
rect 14830 -25421 14836 -25387
rect 14790 -25459 14836 -25421
rect 14790 -25493 14796 -25459
rect 14830 -25493 14836 -25459
rect 14790 -25531 14836 -25493
rect 14790 -25565 14796 -25531
rect 14830 -25565 14836 -25531
rect 14790 -25603 14836 -25565
rect 14790 -25637 14796 -25603
rect 14830 -25637 14836 -25603
rect 14790 -25675 14836 -25637
rect 14790 -25709 14796 -25675
rect 14830 -25709 14836 -25675
rect 14790 -25747 14836 -25709
rect 14790 -25781 14796 -25747
rect 14830 -25781 14836 -25747
rect 14790 -25819 14836 -25781
rect 13812 -25853 13828 -25842
rect 12024 -25922 12512 -25916
rect 12024 -25956 12071 -25922
rect 12105 -25956 12143 -25922
rect 12177 -25956 12215 -25922
rect 12249 -25956 12287 -25922
rect 12321 -25956 12359 -25922
rect 12393 -25956 12431 -25922
rect 12465 -25956 12512 -25922
rect 12024 -25962 12512 -25956
rect 13042 -25922 13530 -25916
rect 13042 -25956 13089 -25922
rect 13123 -25956 13161 -25922
rect 13195 -25956 13233 -25922
rect 13267 -25956 13305 -25922
rect 13339 -25956 13377 -25922
rect 13411 -25956 13449 -25922
rect 13483 -25956 13530 -25922
rect 13042 -25962 13530 -25956
rect 12242 -26028 12302 -25962
rect 13264 -26028 13324 -25962
rect 13768 -26028 13828 -25853
rect 14790 -25853 14796 -25819
rect 14830 -25853 14836 -25819
rect 15808 -25349 15814 -25342
rect 15848 -25342 15860 -25315
rect 16814 -25315 16874 -25156
rect 17114 -25212 17602 -25206
rect 17114 -25246 17161 -25212
rect 17195 -25246 17233 -25212
rect 17267 -25246 17305 -25212
rect 17339 -25246 17377 -25212
rect 17411 -25246 17449 -25212
rect 17483 -25246 17521 -25212
rect 17555 -25246 17602 -25212
rect 17114 -25252 17602 -25246
rect 16814 -25342 16832 -25315
rect 15848 -25349 15854 -25342
rect 15808 -25387 15854 -25349
rect 15808 -25421 15814 -25387
rect 15848 -25421 15854 -25387
rect 15808 -25459 15854 -25421
rect 15808 -25493 15814 -25459
rect 15848 -25493 15854 -25459
rect 15808 -25531 15854 -25493
rect 15808 -25565 15814 -25531
rect 15848 -25565 15854 -25531
rect 15808 -25603 15854 -25565
rect 15808 -25637 15814 -25603
rect 15848 -25637 15854 -25603
rect 15808 -25675 15854 -25637
rect 15808 -25709 15814 -25675
rect 15848 -25709 15854 -25675
rect 15808 -25747 15854 -25709
rect 15808 -25781 15814 -25747
rect 15848 -25781 15854 -25747
rect 15808 -25819 15854 -25781
rect 15808 -25828 15814 -25819
rect 14790 -25884 14836 -25853
rect 15802 -25853 15814 -25828
rect 15848 -25828 15854 -25819
rect 16826 -25349 16832 -25342
rect 16866 -25342 16874 -25315
rect 17834 -25315 17894 -25058
rect 18848 -25100 18920 -25096
rect 18848 -25152 18858 -25100
rect 18910 -25152 18920 -25100
rect 18848 -25156 18920 -25152
rect 18132 -25212 18620 -25206
rect 18132 -25246 18179 -25212
rect 18213 -25246 18251 -25212
rect 18285 -25246 18323 -25212
rect 18357 -25246 18395 -25212
rect 18429 -25246 18467 -25212
rect 18501 -25246 18539 -25212
rect 18573 -25246 18620 -25212
rect 18132 -25252 18620 -25246
rect 16866 -25349 16872 -25342
rect 16826 -25387 16872 -25349
rect 17834 -25349 17850 -25315
rect 17884 -25349 17894 -25315
rect 18854 -25315 18914 -25156
rect 19150 -25212 19638 -25206
rect 19150 -25246 19197 -25212
rect 19231 -25246 19269 -25212
rect 19303 -25246 19341 -25212
rect 19375 -25246 19413 -25212
rect 19447 -25246 19485 -25212
rect 19519 -25246 19557 -25212
rect 19591 -25246 19638 -25212
rect 19150 -25252 19638 -25246
rect 18854 -25328 18868 -25315
rect 17834 -25354 17894 -25349
rect 18862 -25349 18868 -25328
rect 18902 -25328 18914 -25315
rect 19868 -25315 19928 -25058
rect 20366 -25206 20426 -24730
rect 20888 -25096 20948 -24621
rect 21906 -24621 21922 -24592
rect 21956 -24592 21962 -24587
rect 22934 -24083 22994 -23990
rect 22934 -24117 22940 -24083
rect 22974 -24117 22994 -24083
rect 22934 -24140 22994 -24117
rect 22934 -24155 22980 -24140
rect 22934 -24189 22940 -24155
rect 22974 -24189 22980 -24155
rect 22934 -24227 22980 -24189
rect 22934 -24261 22940 -24227
rect 22974 -24261 22980 -24227
rect 22934 -24299 22980 -24261
rect 22934 -24333 22940 -24299
rect 22974 -24333 22980 -24299
rect 22934 -24371 22980 -24333
rect 22934 -24405 22940 -24371
rect 22974 -24405 22980 -24371
rect 22934 -24443 22980 -24405
rect 22934 -24477 22940 -24443
rect 22974 -24477 22980 -24443
rect 22934 -24515 22980 -24477
rect 22934 -24549 22940 -24515
rect 22974 -24549 22980 -24515
rect 22934 -24587 22980 -24549
rect 21956 -24621 21966 -24592
rect 22934 -24606 22940 -24587
rect 21186 -24690 21674 -24684
rect 21186 -24724 21233 -24690
rect 21267 -24724 21305 -24690
rect 21339 -24724 21377 -24690
rect 21411 -24724 21449 -24690
rect 21483 -24724 21521 -24690
rect 21555 -24724 21593 -24690
rect 21627 -24724 21674 -24690
rect 21186 -24730 21674 -24724
rect 20882 -25100 20954 -25096
rect 20882 -25152 20892 -25100
rect 20944 -25152 20954 -25100
rect 20882 -25156 20954 -25152
rect 20168 -25212 20656 -25206
rect 20168 -25246 20215 -25212
rect 20249 -25246 20287 -25212
rect 20321 -25246 20359 -25212
rect 20393 -25246 20431 -25212
rect 20465 -25246 20503 -25212
rect 20537 -25246 20575 -25212
rect 20609 -25246 20656 -25212
rect 20168 -25252 20656 -25246
rect 18902 -25349 18908 -25328
rect 19868 -25338 19886 -25315
rect 16826 -25421 16832 -25387
rect 16866 -25421 16872 -25387
rect 16826 -25459 16872 -25421
rect 16826 -25493 16832 -25459
rect 16866 -25493 16872 -25459
rect 16826 -25531 16872 -25493
rect 16826 -25565 16832 -25531
rect 16866 -25565 16872 -25531
rect 16826 -25603 16872 -25565
rect 16826 -25637 16832 -25603
rect 16866 -25637 16872 -25603
rect 16826 -25675 16872 -25637
rect 16826 -25709 16832 -25675
rect 16866 -25709 16872 -25675
rect 16826 -25747 16872 -25709
rect 16826 -25781 16832 -25747
rect 16866 -25781 16872 -25747
rect 16826 -25819 16872 -25781
rect 15848 -25853 15862 -25828
rect 14060 -25922 14548 -25916
rect 14060 -25956 14107 -25922
rect 14141 -25956 14179 -25922
rect 14213 -25956 14251 -25922
rect 14285 -25956 14323 -25922
rect 14357 -25956 14395 -25922
rect 14429 -25956 14467 -25922
rect 14501 -25956 14548 -25922
rect 14060 -25962 14548 -25956
rect 15078 -25922 15566 -25916
rect 15078 -25956 15125 -25922
rect 15159 -25956 15197 -25922
rect 15231 -25956 15269 -25922
rect 15303 -25956 15341 -25922
rect 15375 -25956 15413 -25922
rect 15447 -25956 15485 -25922
rect 15519 -25956 15566 -25922
rect 15078 -25962 15566 -25956
rect 14286 -26028 14346 -25962
rect 15294 -26028 15354 -25962
rect 15802 -26028 15862 -25853
rect 16826 -25853 16832 -25819
rect 16866 -25853 16872 -25819
rect 17844 -25387 17890 -25354
rect 17844 -25421 17850 -25387
rect 17884 -25421 17890 -25387
rect 17844 -25459 17890 -25421
rect 17844 -25493 17850 -25459
rect 17884 -25493 17890 -25459
rect 17844 -25531 17890 -25493
rect 17844 -25565 17850 -25531
rect 17884 -25565 17890 -25531
rect 17844 -25603 17890 -25565
rect 17844 -25637 17850 -25603
rect 17884 -25637 17890 -25603
rect 17844 -25675 17890 -25637
rect 17844 -25709 17850 -25675
rect 17884 -25709 17890 -25675
rect 17844 -25747 17890 -25709
rect 17844 -25781 17850 -25747
rect 17884 -25781 17890 -25747
rect 17844 -25819 17890 -25781
rect 17844 -25832 17850 -25819
rect 16826 -25884 16872 -25853
rect 17838 -25853 17850 -25832
rect 17884 -25832 17890 -25819
rect 18862 -25387 18908 -25349
rect 18862 -25421 18868 -25387
rect 18902 -25421 18908 -25387
rect 18862 -25459 18908 -25421
rect 18862 -25493 18868 -25459
rect 18902 -25493 18908 -25459
rect 18862 -25531 18908 -25493
rect 18862 -25565 18868 -25531
rect 18902 -25565 18908 -25531
rect 18862 -25603 18908 -25565
rect 18862 -25637 18868 -25603
rect 18902 -25637 18908 -25603
rect 18862 -25675 18908 -25637
rect 18862 -25709 18868 -25675
rect 18902 -25709 18908 -25675
rect 18862 -25747 18908 -25709
rect 18862 -25781 18868 -25747
rect 18902 -25781 18908 -25747
rect 18862 -25819 18908 -25781
rect 17884 -25853 17898 -25832
rect 16298 -25916 16358 -25914
rect 16096 -25922 16584 -25916
rect 16096 -25956 16143 -25922
rect 16177 -25956 16215 -25922
rect 16249 -25956 16287 -25922
rect 16321 -25956 16359 -25922
rect 16393 -25956 16431 -25922
rect 16465 -25956 16503 -25922
rect 16537 -25956 16584 -25922
rect 16096 -25962 16584 -25956
rect 17114 -25922 17602 -25916
rect 17114 -25956 17161 -25922
rect 17195 -25956 17233 -25922
rect 17267 -25956 17305 -25922
rect 17339 -25956 17377 -25922
rect 17411 -25956 17449 -25922
rect 17483 -25956 17521 -25922
rect 17555 -25956 17602 -25922
rect 17114 -25962 17602 -25956
rect 16298 -26028 16358 -25962
rect 17344 -26028 17404 -25962
rect 17838 -26028 17898 -25853
rect 18862 -25853 18868 -25819
rect 18902 -25853 18908 -25819
rect 19880 -25349 19886 -25338
rect 19920 -25338 19928 -25315
rect 20888 -25315 20948 -25156
rect 21394 -25206 21454 -24730
rect 21906 -24998 21966 -24621
rect 22924 -24621 22940 -24606
rect 22974 -24606 22980 -24587
rect 22974 -24621 22984 -24606
rect 22204 -24690 22692 -24684
rect 22204 -24724 22251 -24690
rect 22285 -24724 22323 -24690
rect 22357 -24724 22395 -24690
rect 22429 -24724 22467 -24690
rect 22501 -24724 22539 -24690
rect 22573 -24724 22611 -24690
rect 22645 -24724 22692 -24690
rect 22204 -24730 22692 -24724
rect 21900 -25002 21972 -24998
rect 21900 -25054 21910 -25002
rect 21962 -25054 21972 -25002
rect 21900 -25058 21972 -25054
rect 21186 -25212 21674 -25206
rect 21186 -25246 21233 -25212
rect 21267 -25246 21305 -25212
rect 21339 -25246 21377 -25212
rect 21411 -25246 21449 -25212
rect 21483 -25246 21521 -25212
rect 21555 -25246 21593 -25212
rect 21627 -25246 21674 -25212
rect 21186 -25252 21674 -25246
rect 20888 -25336 20904 -25315
rect 19920 -25349 19926 -25338
rect 19880 -25387 19926 -25349
rect 19880 -25421 19886 -25387
rect 19920 -25421 19926 -25387
rect 19880 -25459 19926 -25421
rect 19880 -25493 19886 -25459
rect 19920 -25493 19926 -25459
rect 19880 -25531 19926 -25493
rect 19880 -25565 19886 -25531
rect 19920 -25565 19926 -25531
rect 19880 -25603 19926 -25565
rect 19880 -25637 19886 -25603
rect 19920 -25637 19926 -25603
rect 19880 -25675 19926 -25637
rect 19880 -25709 19886 -25675
rect 19920 -25709 19926 -25675
rect 19880 -25747 19926 -25709
rect 19880 -25781 19886 -25747
rect 19920 -25781 19926 -25747
rect 19880 -25819 19926 -25781
rect 19880 -25838 19886 -25819
rect 18862 -25884 18908 -25853
rect 19876 -25853 19886 -25838
rect 19920 -25838 19926 -25819
rect 20898 -25349 20904 -25336
rect 20938 -25336 20948 -25315
rect 21906 -25315 21966 -25058
rect 22386 -25206 22446 -24730
rect 22924 -25096 22984 -24621
rect 23648 -24998 23708 -12606
rect 24816 -12629 24855 -12595
rect 24889 -12629 24928 -12595
rect 24816 -12667 24928 -12629
rect 24816 -12701 24855 -12667
rect 24889 -12701 24928 -12667
rect 24816 -12739 24928 -12701
rect 24816 -12773 24855 -12739
rect 24889 -12773 24928 -12739
rect 24816 -12811 24928 -12773
rect 24816 -12845 24855 -12811
rect 24889 -12845 24928 -12811
rect 24816 -12883 24928 -12845
rect 24816 -12917 24855 -12883
rect 24889 -12917 24928 -12883
rect 24816 -12955 24928 -12917
rect 24816 -12989 24855 -12955
rect 24889 -12989 24928 -12955
rect 24816 -13027 24928 -12989
rect 24816 -13061 24855 -13027
rect 24889 -13061 24928 -13027
rect 24816 -13099 24928 -13061
rect 24816 -13133 24855 -13099
rect 24889 -13133 24928 -13099
rect 24816 -13171 24928 -13133
rect 24816 -13205 24855 -13171
rect 24889 -13205 24928 -13171
rect 24816 -13243 24928 -13205
rect 24816 -13277 24855 -13243
rect 24889 -13277 24928 -13243
rect 24816 -13315 24928 -13277
rect 24816 -13349 24855 -13315
rect 24889 -13349 24928 -13315
rect 24816 -13387 24928 -13349
rect 24816 -13421 24855 -13387
rect 24889 -13421 24928 -13387
rect 24816 -13459 24928 -13421
rect 24816 -13493 24855 -13459
rect 24889 -13493 24928 -13459
rect 24816 -13531 24928 -13493
rect 24816 -13565 24855 -13531
rect 24889 -13565 24928 -13531
rect 24816 -13603 24928 -13565
rect 24816 -13637 24855 -13603
rect 24889 -13637 24928 -13603
rect 24816 -13675 24928 -13637
rect 24816 -13709 24855 -13675
rect 24889 -13709 24928 -13675
rect 24816 -13747 24928 -13709
rect 24816 -13781 24855 -13747
rect 24889 -13781 24928 -13747
rect 24816 -13819 24928 -13781
rect 24816 -13853 24855 -13819
rect 24889 -13853 24928 -13819
rect 24816 -13891 24928 -13853
rect 24816 -13925 24855 -13891
rect 24889 -13925 24928 -13891
rect 24816 -13963 24928 -13925
rect 24816 -13997 24855 -13963
rect 24889 -13997 24928 -13963
rect 24816 -14035 24928 -13997
rect 24816 -14069 24855 -14035
rect 24889 -14069 24928 -14035
rect 24816 -14107 24928 -14069
rect 24816 -14141 24855 -14107
rect 24889 -14141 24928 -14107
rect 24816 -14179 24928 -14141
rect 24816 -14213 24855 -14179
rect 24889 -14213 24928 -14179
rect 24816 -14251 24928 -14213
rect 24816 -14285 24855 -14251
rect 24889 -14285 24928 -14251
rect 24816 -14323 24928 -14285
rect 24816 -14357 24855 -14323
rect 24889 -14357 24928 -14323
rect 24816 -14395 24928 -14357
rect 24816 -14429 24855 -14395
rect 24889 -14429 24928 -14395
rect 24816 -14467 24928 -14429
rect 24816 -14501 24855 -14467
rect 24889 -14501 24928 -14467
rect 24816 -14539 24928 -14501
rect 24816 -14573 24855 -14539
rect 24889 -14573 24928 -14539
rect 24816 -14611 24928 -14573
rect 24816 -14645 24855 -14611
rect 24889 -14645 24928 -14611
rect 24816 -14683 24928 -14645
rect 24816 -14717 24855 -14683
rect 24889 -14717 24928 -14683
rect 24816 -14755 24928 -14717
rect 24816 -14789 24855 -14755
rect 24889 -14789 24928 -14755
rect 24816 -14827 24928 -14789
rect 24816 -14861 24855 -14827
rect 24889 -14861 24928 -14827
rect 24816 -14899 24928 -14861
rect 24816 -14933 24855 -14899
rect 24889 -14933 24928 -14899
rect 24816 -14971 24928 -14933
rect 24816 -15005 24855 -14971
rect 24889 -15005 24928 -14971
rect 24816 -15043 24928 -15005
rect 24816 -15077 24855 -15043
rect 24889 -15077 24928 -15043
rect 24816 -15115 24928 -15077
rect 24816 -15149 24855 -15115
rect 24889 -15149 24928 -15115
rect 24816 -15187 24928 -15149
rect 24816 -15221 24855 -15187
rect 24889 -15221 24928 -15187
rect 24816 -15259 24928 -15221
rect 24816 -15293 24855 -15259
rect 24889 -15293 24928 -15259
rect 24816 -15331 24928 -15293
rect 24816 -15365 24855 -15331
rect 24889 -15365 24928 -15331
rect 24816 -15403 24928 -15365
rect 24816 -15437 24855 -15403
rect 24889 -15437 24928 -15403
rect 24816 -15475 24928 -15437
rect 24816 -15509 24855 -15475
rect 24889 -15509 24928 -15475
rect 24816 -15547 24928 -15509
rect 24816 -15581 24855 -15547
rect 24889 -15581 24928 -15547
rect 24816 -15619 24928 -15581
rect 24816 -15653 24855 -15619
rect 24889 -15653 24928 -15619
rect 24816 -15691 24928 -15653
rect 24816 -15725 24855 -15691
rect 24889 -15725 24928 -15691
rect 24816 -15763 24928 -15725
rect 24816 -15797 24855 -15763
rect 24889 -15797 24928 -15763
rect 24816 -15835 24928 -15797
rect 24816 -15869 24855 -15835
rect 24889 -15869 24928 -15835
rect 24816 -15907 24928 -15869
rect 24816 -15941 24855 -15907
rect 24889 -15941 24928 -15907
rect 24816 -15979 24928 -15941
rect 24816 -16013 24855 -15979
rect 24889 -16013 24928 -15979
rect 24816 -16051 24928 -16013
rect 24816 -16085 24855 -16051
rect 24889 -16085 24928 -16051
rect 24816 -16123 24928 -16085
rect 24816 -16157 24855 -16123
rect 24889 -16157 24928 -16123
rect 24816 -16195 24928 -16157
rect 24816 -16229 24855 -16195
rect 24889 -16229 24928 -16195
rect 24816 -16267 24928 -16229
rect 24816 -16301 24855 -16267
rect 24889 -16301 24928 -16267
rect 24816 -16339 24928 -16301
rect 24816 -16373 24855 -16339
rect 24889 -16373 24928 -16339
rect 24816 -16411 24928 -16373
rect 24816 -16445 24855 -16411
rect 24889 -16445 24928 -16411
rect 24816 -16483 24928 -16445
rect 24816 -16517 24855 -16483
rect 24889 -16517 24928 -16483
rect 24816 -16555 24928 -16517
rect 24816 -16589 24855 -16555
rect 24889 -16589 24928 -16555
rect 24816 -16627 24928 -16589
rect 24816 -16661 24855 -16627
rect 24889 -16661 24928 -16627
rect 24816 -16699 24928 -16661
rect 24816 -16733 24855 -16699
rect 24889 -16733 24928 -16699
rect 24816 -16771 24928 -16733
rect 24816 -16805 24855 -16771
rect 24889 -16805 24928 -16771
rect 24816 -16843 24928 -16805
rect 24816 -16877 24855 -16843
rect 24889 -16877 24928 -16843
rect 24816 -16915 24928 -16877
rect 24816 -16949 24855 -16915
rect 24889 -16949 24928 -16915
rect 24816 -16987 24928 -16949
rect 24816 -17021 24855 -16987
rect 24889 -17021 24928 -16987
rect 24816 -17059 24928 -17021
rect 24816 -17093 24855 -17059
rect 24889 -17093 24928 -17059
rect 24816 -17131 24928 -17093
rect 24816 -17165 24855 -17131
rect 24889 -17165 24928 -17131
rect 24816 -17203 24928 -17165
rect 24816 -17237 24855 -17203
rect 24889 -17237 24928 -17203
rect 24816 -17275 24928 -17237
rect 24816 -17309 24855 -17275
rect 24889 -17309 24928 -17275
rect 24816 -17347 24928 -17309
rect 24816 -17381 24855 -17347
rect 24889 -17381 24928 -17347
rect 24816 -17419 24928 -17381
rect 24816 -17453 24855 -17419
rect 24889 -17453 24928 -17419
rect 24816 -17491 24928 -17453
rect 24816 -17525 24855 -17491
rect 24889 -17525 24928 -17491
rect 24816 -17563 24928 -17525
rect 24816 -17597 24855 -17563
rect 24889 -17597 24928 -17563
rect 24816 -17635 24928 -17597
rect 24816 -17669 24855 -17635
rect 24889 -17669 24928 -17635
rect 24816 -17707 24928 -17669
rect 24816 -17741 24855 -17707
rect 24889 -17741 24928 -17707
rect 24816 -17779 24928 -17741
rect 24816 -17813 24855 -17779
rect 24889 -17813 24928 -17779
rect 24816 -17851 24928 -17813
rect 24816 -17885 24855 -17851
rect 24889 -17885 24928 -17851
rect 24816 -17923 24928 -17885
rect 24816 -17957 24855 -17923
rect 24889 -17957 24928 -17923
rect 24816 -17995 24928 -17957
rect 24816 -18029 24855 -17995
rect 24889 -18029 24928 -17995
rect 24816 -18067 24928 -18029
rect 24816 -18101 24855 -18067
rect 24889 -18101 24928 -18067
rect 24816 -18139 24928 -18101
rect 24816 -18173 24855 -18139
rect 24889 -18173 24928 -18139
rect 24816 -18211 24928 -18173
rect 24816 -18245 24855 -18211
rect 24889 -18245 24928 -18211
rect 24816 -18283 24928 -18245
rect 24816 -18317 24855 -18283
rect 24889 -18317 24928 -18283
rect 24816 -18355 24928 -18317
rect 24816 -18389 24855 -18355
rect 24889 -18389 24928 -18355
rect 24816 -18427 24928 -18389
rect 24816 -18461 24855 -18427
rect 24889 -18461 24928 -18427
rect 24816 -18499 24928 -18461
rect 24816 -18533 24855 -18499
rect 24889 -18533 24928 -18499
rect 24816 -18571 24928 -18533
rect 24816 -18605 24855 -18571
rect 24889 -18605 24928 -18571
rect 24816 -18643 24928 -18605
rect 24816 -18677 24855 -18643
rect 24889 -18677 24928 -18643
rect 24816 -18715 24928 -18677
rect 24816 -18749 24855 -18715
rect 24889 -18749 24928 -18715
rect 24816 -18787 24928 -18749
rect 24816 -18821 24855 -18787
rect 24889 -18821 24928 -18787
rect 24816 -18859 24928 -18821
rect 24816 -18893 24855 -18859
rect 24889 -18893 24928 -18859
rect 24816 -18931 24928 -18893
rect 24816 -18965 24855 -18931
rect 24889 -18965 24928 -18931
rect 24816 -19003 24928 -18965
rect 24816 -19037 24855 -19003
rect 24889 -19037 24928 -19003
rect 24816 -19075 24928 -19037
rect 24816 -19109 24855 -19075
rect 24889 -19109 24928 -19075
rect 24816 -19147 24928 -19109
rect 24816 -19181 24855 -19147
rect 24889 -19181 24928 -19147
rect 24816 -19219 24928 -19181
rect 24816 -19253 24855 -19219
rect 24889 -19253 24928 -19219
rect 24816 -19291 24928 -19253
rect 24816 -19325 24855 -19291
rect 24889 -19325 24928 -19291
rect 24816 -19363 24928 -19325
rect 24816 -19397 24855 -19363
rect 24889 -19397 24928 -19363
rect 24816 -19435 24928 -19397
rect 24816 -19469 24855 -19435
rect 24889 -19469 24928 -19435
rect 24816 -19507 24928 -19469
rect 24816 -19541 24855 -19507
rect 24889 -19541 24928 -19507
rect 24816 -19579 24928 -19541
rect 24816 -19613 24855 -19579
rect 24889 -19613 24928 -19579
rect 24816 -19651 24928 -19613
rect 24816 -19685 24855 -19651
rect 24889 -19685 24928 -19651
rect 24816 -19723 24928 -19685
rect 24816 -19757 24855 -19723
rect 24889 -19757 24928 -19723
rect 24816 -19795 24928 -19757
rect 24816 -19829 24855 -19795
rect 24889 -19829 24928 -19795
rect 24816 -19867 24928 -19829
rect 24816 -19901 24855 -19867
rect 24889 -19901 24928 -19867
rect 24816 -19939 24928 -19901
rect 24816 -19973 24855 -19939
rect 24889 -19973 24928 -19939
rect 24816 -20011 24928 -19973
rect 24816 -20045 24855 -20011
rect 24889 -20045 24928 -20011
rect 24816 -20083 24928 -20045
rect 24816 -20117 24855 -20083
rect 24889 -20117 24928 -20083
rect 24816 -20155 24928 -20117
rect 24816 -20189 24855 -20155
rect 24889 -20189 24928 -20155
rect 24816 -20227 24928 -20189
rect 24816 -20261 24855 -20227
rect 24889 -20261 24928 -20227
rect 24816 -20299 24928 -20261
rect 24816 -20333 24855 -20299
rect 24889 -20333 24928 -20299
rect 24816 -20371 24928 -20333
rect 24816 -20405 24855 -20371
rect 24889 -20405 24928 -20371
rect 24816 -20443 24928 -20405
rect 24816 -20477 24855 -20443
rect 24889 -20477 24928 -20443
rect 24816 -20515 24928 -20477
rect 24816 -20549 24855 -20515
rect 24889 -20549 24928 -20515
rect 24816 -20587 24928 -20549
rect 24816 -20621 24855 -20587
rect 24889 -20621 24928 -20587
rect 24816 -20659 24928 -20621
rect 24816 -20693 24855 -20659
rect 24889 -20693 24928 -20659
rect 24816 -20731 24928 -20693
rect 24816 -20765 24855 -20731
rect 24889 -20765 24928 -20731
rect 24816 -20803 24928 -20765
rect 24816 -20837 24855 -20803
rect 24889 -20837 24928 -20803
rect 24816 -20875 24928 -20837
rect 24816 -20909 24855 -20875
rect 24889 -20909 24928 -20875
rect 24816 -20947 24928 -20909
rect 24816 -20981 24855 -20947
rect 24889 -20981 24928 -20947
rect 24816 -21019 24928 -20981
rect 24816 -21053 24855 -21019
rect 24889 -21053 24928 -21019
rect 24816 -21091 24928 -21053
rect 24816 -21125 24855 -21091
rect 24889 -21125 24928 -21091
rect 24816 -21163 24928 -21125
rect 24816 -21197 24855 -21163
rect 24889 -21197 24928 -21163
rect 24816 -21235 24928 -21197
rect 24816 -21269 24855 -21235
rect 24889 -21269 24928 -21235
rect 24816 -21307 24928 -21269
rect 24816 -21341 24855 -21307
rect 24889 -21341 24928 -21307
rect 24816 -21379 24928 -21341
rect 24816 -21413 24855 -21379
rect 24889 -21413 24928 -21379
rect 24816 -21451 24928 -21413
rect 24816 -21485 24855 -21451
rect 24889 -21485 24928 -21451
rect 24816 -21523 24928 -21485
rect 24816 -21557 24855 -21523
rect 24889 -21557 24928 -21523
rect 24816 -21595 24928 -21557
rect 24816 -21629 24855 -21595
rect 24889 -21629 24928 -21595
rect 24816 -21667 24928 -21629
rect 24816 -21701 24855 -21667
rect 24889 -21701 24928 -21667
rect 24816 -21739 24928 -21701
rect 24816 -21773 24855 -21739
rect 24889 -21773 24928 -21739
rect 24816 -21811 24928 -21773
rect 24816 -21845 24855 -21811
rect 24889 -21845 24928 -21811
rect 24816 -21883 24928 -21845
rect 24816 -21917 24855 -21883
rect 24889 -21917 24928 -21883
rect 24816 -21955 24928 -21917
rect 24816 -21989 24855 -21955
rect 24889 -21989 24928 -21955
rect 24816 -22027 24928 -21989
rect 24816 -22061 24855 -22027
rect 24889 -22061 24928 -22027
rect 24816 -22099 24928 -22061
rect 24816 -22133 24855 -22099
rect 24889 -22133 24928 -22099
rect 24816 -22171 24928 -22133
rect 24816 -22205 24855 -22171
rect 24889 -22205 24928 -22171
rect 24816 -22243 24928 -22205
rect 24816 -22277 24855 -22243
rect 24889 -22277 24928 -22243
rect 24816 -22315 24928 -22277
rect 24816 -22349 24855 -22315
rect 24889 -22349 24928 -22315
rect 24816 -22387 24928 -22349
rect 24816 -22421 24855 -22387
rect 24889 -22421 24928 -22387
rect 24816 -22459 24928 -22421
rect 24816 -22493 24855 -22459
rect 24889 -22493 24928 -22459
rect 24816 -22531 24928 -22493
rect 24816 -22565 24855 -22531
rect 24889 -22565 24928 -22531
rect 24816 -22603 24928 -22565
rect 24816 -22637 24855 -22603
rect 24889 -22637 24928 -22603
rect 24816 -22675 24928 -22637
rect 24816 -22709 24855 -22675
rect 24889 -22709 24928 -22675
rect 24816 -22747 24928 -22709
rect 24816 -22781 24855 -22747
rect 24889 -22781 24928 -22747
rect 24816 -22819 24928 -22781
rect 24816 -22853 24855 -22819
rect 24889 -22853 24928 -22819
rect 24816 -22891 24928 -22853
rect 24816 -22925 24855 -22891
rect 24889 -22925 24928 -22891
rect 24816 -22963 24928 -22925
rect 24816 -22997 24855 -22963
rect 24889 -22997 24928 -22963
rect 24816 -23035 24928 -22997
rect 24816 -23069 24855 -23035
rect 24889 -23069 24928 -23035
rect 24816 -23107 24928 -23069
rect 24816 -23141 24855 -23107
rect 24889 -23141 24928 -23107
rect 24816 -23179 24928 -23141
rect 24816 -23213 24855 -23179
rect 24889 -23213 24928 -23179
rect 24816 -23251 24928 -23213
rect 24816 -23285 24855 -23251
rect 24889 -23285 24928 -23251
rect 24816 -23323 24928 -23285
rect 24816 -23357 24855 -23323
rect 24889 -23357 24928 -23323
rect 24816 -23395 24928 -23357
rect 24816 -23429 24855 -23395
rect 24889 -23429 24928 -23395
rect 24816 -23467 24928 -23429
rect 24816 -23501 24855 -23467
rect 24889 -23501 24928 -23467
rect 24816 -23539 24928 -23501
rect 24816 -23573 24855 -23539
rect 24889 -23573 24928 -23539
rect 24816 -23611 24928 -23573
rect 24816 -23645 24855 -23611
rect 24889 -23645 24928 -23611
rect 24816 -23683 24928 -23645
rect 24816 -23717 24855 -23683
rect 24889 -23717 24928 -23683
rect 24816 -23755 24928 -23717
rect 24816 -23789 24855 -23755
rect 24889 -23789 24928 -23755
rect 24816 -23827 24928 -23789
rect 24816 -23861 24855 -23827
rect 24889 -23861 24928 -23827
rect 23800 -23870 23872 -23866
rect 23800 -23922 23810 -23870
rect 23862 -23922 23872 -23870
rect 23800 -23926 23872 -23922
rect 24816 -23899 24928 -23861
rect 23642 -25002 23714 -24998
rect 23642 -25054 23652 -25002
rect 23704 -25054 23714 -25002
rect 23642 -25058 23714 -25054
rect 22918 -25100 22990 -25096
rect 22918 -25152 22928 -25100
rect 22980 -25152 22990 -25100
rect 22918 -25156 22990 -25152
rect 22204 -25212 22692 -25206
rect 22204 -25246 22251 -25212
rect 22285 -25246 22323 -25212
rect 22357 -25246 22395 -25212
rect 22429 -25246 22467 -25212
rect 22501 -25246 22539 -25212
rect 22573 -25246 22611 -25212
rect 22645 -25246 22692 -25212
rect 22204 -25252 22692 -25246
rect 22386 -25254 22446 -25252
rect 21906 -25326 21922 -25315
rect 20938 -25349 20944 -25336
rect 20898 -25387 20944 -25349
rect 20898 -25421 20904 -25387
rect 20938 -25421 20944 -25387
rect 20898 -25459 20944 -25421
rect 20898 -25493 20904 -25459
rect 20938 -25493 20944 -25459
rect 20898 -25531 20944 -25493
rect 20898 -25565 20904 -25531
rect 20938 -25565 20944 -25531
rect 20898 -25603 20944 -25565
rect 20898 -25637 20904 -25603
rect 20938 -25637 20944 -25603
rect 20898 -25675 20944 -25637
rect 20898 -25709 20904 -25675
rect 20938 -25709 20944 -25675
rect 20898 -25747 20944 -25709
rect 20898 -25781 20904 -25747
rect 20938 -25781 20944 -25747
rect 20898 -25819 20944 -25781
rect 19920 -25853 19936 -25838
rect 18132 -25922 18620 -25916
rect 18132 -25956 18179 -25922
rect 18213 -25956 18251 -25922
rect 18285 -25956 18323 -25922
rect 18357 -25956 18395 -25922
rect 18429 -25956 18467 -25922
rect 18501 -25956 18539 -25922
rect 18573 -25956 18620 -25922
rect 18132 -25962 18620 -25956
rect 19150 -25922 19638 -25916
rect 19150 -25956 19197 -25922
rect 19231 -25956 19269 -25922
rect 19303 -25956 19341 -25922
rect 19375 -25956 19413 -25922
rect 19447 -25956 19485 -25922
rect 19519 -25956 19557 -25922
rect 19591 -25956 19638 -25922
rect 19150 -25962 19638 -25956
rect 18342 -26028 18402 -25962
rect 19354 -26028 19414 -25962
rect 19876 -26028 19936 -25853
rect 20898 -25853 20904 -25819
rect 20938 -25853 20944 -25819
rect 21916 -25349 21922 -25326
rect 21956 -25326 21966 -25315
rect 22924 -25315 22984 -25156
rect 21956 -25349 21962 -25326
rect 22924 -25332 22940 -25315
rect 21916 -25387 21962 -25349
rect 21916 -25421 21922 -25387
rect 21956 -25421 21962 -25387
rect 21916 -25459 21962 -25421
rect 21916 -25493 21922 -25459
rect 21956 -25493 21962 -25459
rect 21916 -25531 21962 -25493
rect 21916 -25565 21922 -25531
rect 21956 -25565 21962 -25531
rect 21916 -25603 21962 -25565
rect 21916 -25637 21922 -25603
rect 21956 -25637 21962 -25603
rect 21916 -25675 21962 -25637
rect 21916 -25709 21922 -25675
rect 21956 -25709 21962 -25675
rect 21916 -25747 21962 -25709
rect 21916 -25781 21922 -25747
rect 21956 -25781 21962 -25747
rect 21916 -25819 21962 -25781
rect 21916 -25844 21922 -25819
rect 20898 -25884 20944 -25853
rect 21904 -25853 21922 -25844
rect 21956 -25844 21962 -25819
rect 22934 -25349 22940 -25332
rect 22974 -25332 22984 -25315
rect 22974 -25349 22980 -25332
rect 22934 -25387 22980 -25349
rect 22934 -25421 22940 -25387
rect 22974 -25421 22980 -25387
rect 22934 -25459 22980 -25421
rect 22934 -25493 22940 -25459
rect 22974 -25493 22980 -25459
rect 22934 -25531 22980 -25493
rect 22934 -25565 22940 -25531
rect 22974 -25565 22980 -25531
rect 22934 -25603 22980 -25565
rect 22934 -25637 22940 -25603
rect 22974 -25637 22980 -25603
rect 22934 -25675 22980 -25637
rect 22934 -25709 22940 -25675
rect 22974 -25709 22980 -25675
rect 22934 -25747 22980 -25709
rect 22934 -25781 22940 -25747
rect 22974 -25781 22980 -25747
rect 22934 -25819 22980 -25781
rect 21956 -25853 21964 -25844
rect 20168 -25922 20656 -25916
rect 20168 -25956 20215 -25922
rect 20249 -25956 20287 -25922
rect 20321 -25956 20359 -25922
rect 20393 -25956 20431 -25922
rect 20465 -25956 20503 -25922
rect 20537 -25956 20575 -25922
rect 20609 -25956 20656 -25922
rect 20168 -25962 20656 -25956
rect 21186 -25922 21674 -25916
rect 21186 -25956 21233 -25922
rect 21267 -25956 21305 -25922
rect 21339 -25956 21377 -25922
rect 21411 -25956 21449 -25922
rect 21483 -25956 21521 -25922
rect 21555 -25956 21593 -25922
rect 21627 -25956 21674 -25922
rect 21186 -25962 21674 -25956
rect 20376 -26028 20436 -25962
rect 21442 -26028 21502 -25962
rect 21904 -26028 21964 -25853
rect 22934 -25853 22940 -25819
rect 22974 -25853 22980 -25819
rect 22934 -25884 22980 -25853
rect 22204 -25922 22692 -25916
rect 22204 -25956 22251 -25922
rect 22285 -25956 22323 -25922
rect 22357 -25956 22395 -25922
rect 22429 -25956 22467 -25922
rect 22501 -25956 22539 -25922
rect 22573 -25956 22611 -25922
rect 22645 -25956 22692 -25922
rect 22204 -25962 22692 -25956
rect 22404 -26028 22464 -25962
rect 3066 -26088 22464 -26028
rect 23806 -26430 23866 -23926
rect 24816 -23933 24855 -23899
rect 24889 -23933 24928 -23899
rect 24816 -23971 24928 -23933
rect 24816 -24005 24855 -23971
rect 24889 -24005 24928 -23971
rect 24816 -24043 24928 -24005
rect 24816 -24077 24855 -24043
rect 24889 -24077 24928 -24043
rect 24816 -24115 24928 -24077
rect 24816 -24149 24855 -24115
rect 24889 -24149 24928 -24115
rect 24816 -24187 24928 -24149
rect 24816 -24221 24855 -24187
rect 24889 -24221 24928 -24187
rect 24816 -24259 24928 -24221
rect 24816 -24293 24855 -24259
rect 24889 -24293 24928 -24259
rect 24816 -24331 24928 -24293
rect 24816 -24365 24855 -24331
rect 24889 -24365 24928 -24331
rect 24816 -24403 24928 -24365
rect 24816 -24437 24855 -24403
rect 24889 -24437 24928 -24403
rect 24816 -24475 24928 -24437
rect 24816 -24509 24855 -24475
rect 24889 -24509 24928 -24475
rect 24816 -24547 24928 -24509
rect 24816 -24581 24855 -24547
rect 24889 -24581 24928 -24547
rect 24816 -24619 24928 -24581
rect 24816 -24653 24855 -24619
rect 24889 -24653 24928 -24619
rect 24816 -24691 24928 -24653
rect 24816 -24725 24855 -24691
rect 24889 -24725 24928 -24691
rect 24816 -24763 24928 -24725
rect 24816 -24797 24855 -24763
rect 24889 -24797 24928 -24763
rect 24816 -24835 24928 -24797
rect 24816 -24869 24855 -24835
rect 24889 -24869 24928 -24835
rect 24816 -24907 24928 -24869
rect 24816 -24941 24855 -24907
rect 24889 -24941 24928 -24907
rect 24816 -24979 24928 -24941
rect 24816 -25013 24855 -24979
rect 24889 -25013 24928 -24979
rect 24816 -25051 24928 -25013
rect 24816 -25085 24855 -25051
rect 24889 -25085 24928 -25051
rect 24816 -25123 24928 -25085
rect 24816 -25157 24855 -25123
rect 24889 -25157 24928 -25123
rect 24816 -25195 24928 -25157
rect 24816 -25229 24855 -25195
rect 24889 -25229 24928 -25195
rect 24816 -25267 24928 -25229
rect 24816 -25301 24855 -25267
rect 24889 -25301 24928 -25267
rect 24816 -25339 24928 -25301
rect 24816 -25373 24855 -25339
rect 24889 -25373 24928 -25339
rect 24816 -25411 24928 -25373
rect 24816 -25445 24855 -25411
rect 24889 -25445 24928 -25411
rect 24816 -25483 24928 -25445
rect 24816 -25517 24855 -25483
rect 24889 -25517 24928 -25483
rect 24816 -25555 24928 -25517
rect 24816 -25589 24855 -25555
rect 24889 -25589 24928 -25555
rect 24816 -25627 24928 -25589
rect 24816 -25661 24855 -25627
rect 24889 -25661 24928 -25627
rect 24816 -25699 24928 -25661
rect 24816 -25733 24855 -25699
rect 24889 -25733 24928 -25699
rect 24816 -25771 24928 -25733
rect 24816 -25805 24855 -25771
rect 24889 -25805 24928 -25771
rect 24816 -25843 24928 -25805
rect 24816 -25877 24855 -25843
rect 24889 -25877 24928 -25843
rect 24816 -25915 24928 -25877
rect 24816 -25949 24855 -25915
rect 24889 -25949 24928 -25915
rect 24816 -25987 24928 -25949
rect 24816 -26021 24855 -25987
rect 24889 -26021 24928 -25987
rect 24816 -26059 24928 -26021
rect 24816 -26093 24855 -26059
rect 24889 -26093 24928 -26059
rect 24816 -26131 24928 -26093
rect 24816 -26165 24855 -26131
rect 24889 -26165 24928 -26131
rect 24816 -26203 24928 -26165
rect 24816 -26237 24855 -26203
rect 24889 -26237 24928 -26203
rect 24816 -26275 24928 -26237
rect 24816 -26309 24855 -26275
rect 24889 -26309 24928 -26275
rect -7518 -26495 23968 -26430
rect -7518 -26611 -7446 -26495
rect 23902 -26611 23968 -26495
rect -7518 -26676 23968 -26611
rect 24816 -26816 24928 -26309
rect -12328 -26844 -11606 -26816
rect -12328 -27088 -12198 -26844
rect -11634 -27088 -11606 -26844
rect -12328 -27116 -11606 -27088
rect 24206 -26844 24928 -26816
rect 24206 -27088 24234 -26844
rect 24798 -27088 24928 -26844
rect 24206 -27116 24928 -27088
rect -12328 -27155 24928 -27116
rect -12328 -27189 -12221 -27155
rect -12187 -27189 -12149 -27155
rect -12115 -27189 -12077 -27155
rect -12043 -27189 -12005 -27155
rect -11971 -27189 -11933 -27155
rect -11899 -27189 -11861 -27155
rect -11827 -27189 -11789 -27155
rect -11755 -27189 -11717 -27155
rect -11683 -27189 -11645 -27155
rect -11611 -27189 -11573 -27155
rect -11539 -27189 -11501 -27155
rect -11467 -27189 -11429 -27155
rect -11395 -27189 -11357 -27155
rect -11323 -27189 -11285 -27155
rect -11251 -27189 -11213 -27155
rect -11179 -27189 -11141 -27155
rect -11107 -27189 -11069 -27155
rect -11035 -27189 -10997 -27155
rect -10963 -27189 -10925 -27155
rect -10891 -27189 -10853 -27155
rect -10819 -27189 -10781 -27155
rect -10747 -27189 -10709 -27155
rect -10675 -27189 -10637 -27155
rect -10603 -27189 -10565 -27155
rect -10531 -27189 -10493 -27155
rect -10459 -27189 -10421 -27155
rect -10387 -27189 -10349 -27155
rect -10315 -27189 -10277 -27155
rect -10243 -27189 -10205 -27155
rect -10171 -27189 -10133 -27155
rect -10099 -27189 -10061 -27155
rect -10027 -27189 -9989 -27155
rect -9955 -27189 -9917 -27155
rect -9883 -27189 -9845 -27155
rect -9811 -27189 -9773 -27155
rect -9739 -27189 -9701 -27155
rect -9667 -27189 -9629 -27155
rect -9595 -27189 -9557 -27155
rect -9523 -27189 -9485 -27155
rect -9451 -27189 -9413 -27155
rect -9379 -27189 -9341 -27155
rect -9307 -27189 -9269 -27155
rect -9235 -27189 -9197 -27155
rect -9163 -27189 -9125 -27155
rect -9091 -27189 -9053 -27155
rect -9019 -27189 -8981 -27155
rect -8947 -27189 -8909 -27155
rect -8875 -27189 -8837 -27155
rect -8803 -27189 -8765 -27155
rect -8731 -27189 -8693 -27155
rect -8659 -27189 -8621 -27155
rect -8587 -27189 -8549 -27155
rect -8515 -27189 -8477 -27155
rect -8443 -27189 -8405 -27155
rect -8371 -27189 -8333 -27155
rect -8299 -27189 -8261 -27155
rect -8227 -27189 -8189 -27155
rect -8155 -27189 -8117 -27155
rect -8083 -27189 -8045 -27155
rect -8011 -27189 -7973 -27155
rect -7939 -27189 -7901 -27155
rect -7867 -27189 -7829 -27155
rect -7795 -27189 -7757 -27155
rect -7723 -27189 -7685 -27155
rect -7651 -27189 -7613 -27155
rect -7579 -27189 -7541 -27155
rect -7507 -27189 -7469 -27155
rect -7435 -27189 -7397 -27155
rect -7363 -27189 -7325 -27155
rect -7291 -27189 -7253 -27155
rect -7219 -27189 -7181 -27155
rect -7147 -27189 -7109 -27155
rect -7075 -27189 -7037 -27155
rect -7003 -27189 -6965 -27155
rect -6931 -27189 -6893 -27155
rect -6859 -27189 -6821 -27155
rect -6787 -27189 -6749 -27155
rect -6715 -27189 -6677 -27155
rect -6643 -27189 -6605 -27155
rect -6571 -27189 -6533 -27155
rect -6499 -27189 -6461 -27155
rect -6427 -27189 -6389 -27155
rect -6355 -27189 -6317 -27155
rect -6283 -27189 -6245 -27155
rect -6211 -27189 -6173 -27155
rect -6139 -27189 -6101 -27155
rect -6067 -27189 -6029 -27155
rect -5995 -27189 -5957 -27155
rect -5923 -27189 -5885 -27155
rect -5851 -27189 -5813 -27155
rect -5779 -27189 -5741 -27155
rect -5707 -27189 -5669 -27155
rect -5635 -27189 -5597 -27155
rect -5563 -27189 -5525 -27155
rect -5491 -27189 -5453 -27155
rect -5419 -27189 -5381 -27155
rect -5347 -27189 -5309 -27155
rect -5275 -27189 -5237 -27155
rect -5203 -27189 -5165 -27155
rect -5131 -27189 -5093 -27155
rect -5059 -27189 -5021 -27155
rect -4987 -27189 -4949 -27155
rect -4915 -27189 -4877 -27155
rect -4843 -27189 -4805 -27155
rect -4771 -27189 -4733 -27155
rect -4699 -27189 -4661 -27155
rect -4627 -27189 -4589 -27155
rect -4555 -27189 -4517 -27155
rect -4483 -27189 -4445 -27155
rect -4411 -27189 -4373 -27155
rect -4339 -27189 -4301 -27155
rect -4267 -27189 -4229 -27155
rect -4195 -27189 -4157 -27155
rect -4123 -27189 -4085 -27155
rect -4051 -27189 -4013 -27155
rect -3979 -27189 -3941 -27155
rect -3907 -27189 -3869 -27155
rect -3835 -27189 -3797 -27155
rect -3763 -27189 -3725 -27155
rect -3691 -27189 -3653 -27155
rect -3619 -27189 -3581 -27155
rect -3547 -27189 -3509 -27155
rect -3475 -27189 -3437 -27155
rect -3403 -27189 -3365 -27155
rect -3331 -27189 -3293 -27155
rect -3259 -27189 -3221 -27155
rect -3187 -27189 -3149 -27155
rect -3115 -27189 -3077 -27155
rect -3043 -27189 -3005 -27155
rect -2971 -27189 -2933 -27155
rect -2899 -27189 -2861 -27155
rect -2827 -27189 -2789 -27155
rect -2755 -27189 -2717 -27155
rect -2683 -27189 -2645 -27155
rect -2611 -27189 -2573 -27155
rect -2539 -27189 -2501 -27155
rect -2467 -27189 -2429 -27155
rect -2395 -27189 -2357 -27155
rect -2323 -27189 -2285 -27155
rect -2251 -27189 -2213 -27155
rect -2179 -27189 -2141 -27155
rect -2107 -27189 -2069 -27155
rect -2035 -27189 -1997 -27155
rect -1963 -27189 -1925 -27155
rect -1891 -27189 -1853 -27155
rect -1819 -27189 -1781 -27155
rect -1747 -27189 -1709 -27155
rect -1675 -27189 -1637 -27155
rect -1603 -27189 -1565 -27155
rect -1531 -27189 -1493 -27155
rect -1459 -27189 -1421 -27155
rect -1387 -27189 -1349 -27155
rect -1315 -27189 -1277 -27155
rect -1243 -27189 -1205 -27155
rect -1171 -27189 -1133 -27155
rect -1099 -27189 -1061 -27155
rect -1027 -27189 -989 -27155
rect -955 -27189 -917 -27155
rect -883 -27189 -845 -27155
rect -811 -27189 -773 -27155
rect -739 -27189 -701 -27155
rect -667 -27189 -629 -27155
rect -595 -27189 -557 -27155
rect -523 -27189 -485 -27155
rect -451 -27189 -413 -27155
rect -379 -27189 -341 -27155
rect -307 -27189 -269 -27155
rect -235 -27189 -197 -27155
rect -163 -27189 -125 -27155
rect -91 -27189 -53 -27155
rect -19 -27189 19 -27155
rect 53 -27189 91 -27155
rect 125 -27189 163 -27155
rect 197 -27189 235 -27155
rect 269 -27189 307 -27155
rect 341 -27189 379 -27155
rect 413 -27189 451 -27155
rect 485 -27189 523 -27155
rect 557 -27189 595 -27155
rect 629 -27189 667 -27155
rect 701 -27189 739 -27155
rect 773 -27189 811 -27155
rect 845 -27189 883 -27155
rect 917 -27189 955 -27155
rect 989 -27189 1027 -27155
rect 1061 -27189 1099 -27155
rect 1133 -27189 1171 -27155
rect 1205 -27189 1243 -27155
rect 1277 -27189 1315 -27155
rect 1349 -27189 1387 -27155
rect 1421 -27189 1459 -27155
rect 1493 -27189 1531 -27155
rect 1565 -27189 1603 -27155
rect 1637 -27189 1675 -27155
rect 1709 -27189 1747 -27155
rect 1781 -27189 1819 -27155
rect 1853 -27189 1891 -27155
rect 1925 -27189 1963 -27155
rect 1997 -27189 2035 -27155
rect 2069 -27189 2107 -27155
rect 2141 -27189 2179 -27155
rect 2213 -27189 2251 -27155
rect 2285 -27189 2323 -27155
rect 2357 -27189 2395 -27155
rect 2429 -27189 2467 -27155
rect 2501 -27189 2539 -27155
rect 2573 -27189 2611 -27155
rect 2645 -27189 2683 -27155
rect 2717 -27189 2755 -27155
rect 2789 -27189 2827 -27155
rect 2861 -27189 2899 -27155
rect 2933 -27189 2971 -27155
rect 3005 -27189 3043 -27155
rect 3077 -27189 3115 -27155
rect 3149 -27189 3187 -27155
rect 3221 -27189 3259 -27155
rect 3293 -27189 3331 -27155
rect 3365 -27189 3403 -27155
rect 3437 -27189 3475 -27155
rect 3509 -27189 3547 -27155
rect 3581 -27189 3619 -27155
rect 3653 -27189 3691 -27155
rect 3725 -27189 3763 -27155
rect 3797 -27189 3835 -27155
rect 3869 -27189 3907 -27155
rect 3941 -27189 3979 -27155
rect 4013 -27189 4051 -27155
rect 4085 -27189 4123 -27155
rect 4157 -27189 4195 -27155
rect 4229 -27189 4267 -27155
rect 4301 -27189 4339 -27155
rect 4373 -27189 4411 -27155
rect 4445 -27189 4483 -27155
rect 4517 -27189 4555 -27155
rect 4589 -27189 4627 -27155
rect 4661 -27189 4699 -27155
rect 4733 -27189 4771 -27155
rect 4805 -27189 4843 -27155
rect 4877 -27189 4915 -27155
rect 4949 -27189 4987 -27155
rect 5021 -27189 5059 -27155
rect 5093 -27189 5131 -27155
rect 5165 -27189 5203 -27155
rect 5237 -27189 5275 -27155
rect 5309 -27189 5347 -27155
rect 5381 -27189 5419 -27155
rect 5453 -27189 5491 -27155
rect 5525 -27189 5563 -27155
rect 5597 -27189 5635 -27155
rect 5669 -27189 5707 -27155
rect 5741 -27189 5779 -27155
rect 5813 -27189 5851 -27155
rect 5885 -27189 5923 -27155
rect 5957 -27189 5995 -27155
rect 6029 -27189 6067 -27155
rect 6101 -27189 6139 -27155
rect 6173 -27189 6211 -27155
rect 6245 -27189 6283 -27155
rect 6317 -27189 6355 -27155
rect 6389 -27189 6427 -27155
rect 6461 -27189 6499 -27155
rect 6533 -27189 6571 -27155
rect 6605 -27189 6643 -27155
rect 6677 -27189 6715 -27155
rect 6749 -27189 6787 -27155
rect 6821 -27189 6859 -27155
rect 6893 -27189 6931 -27155
rect 6965 -27189 7003 -27155
rect 7037 -27189 7075 -27155
rect 7109 -27189 7147 -27155
rect 7181 -27189 7219 -27155
rect 7253 -27189 7291 -27155
rect 7325 -27189 7363 -27155
rect 7397 -27189 7435 -27155
rect 7469 -27189 7507 -27155
rect 7541 -27189 7579 -27155
rect 7613 -27189 7651 -27155
rect 7685 -27189 7723 -27155
rect 7757 -27189 7795 -27155
rect 7829 -27189 7867 -27155
rect 7901 -27189 7939 -27155
rect 7973 -27189 8011 -27155
rect 8045 -27189 8083 -27155
rect 8117 -27189 8155 -27155
rect 8189 -27189 8227 -27155
rect 8261 -27189 8299 -27155
rect 8333 -27189 8371 -27155
rect 8405 -27189 8443 -27155
rect 8477 -27189 8515 -27155
rect 8549 -27189 8587 -27155
rect 8621 -27189 8659 -27155
rect 8693 -27189 8731 -27155
rect 8765 -27189 8803 -27155
rect 8837 -27189 8875 -27155
rect 8909 -27189 8947 -27155
rect 8981 -27189 9019 -27155
rect 9053 -27189 9091 -27155
rect 9125 -27189 9163 -27155
rect 9197 -27189 9235 -27155
rect 9269 -27189 9307 -27155
rect 9341 -27189 9379 -27155
rect 9413 -27189 9451 -27155
rect 9485 -27189 9523 -27155
rect 9557 -27189 9595 -27155
rect 9629 -27189 9667 -27155
rect 9701 -27189 9739 -27155
rect 9773 -27189 9811 -27155
rect 9845 -27189 9883 -27155
rect 9917 -27189 9955 -27155
rect 9989 -27189 10027 -27155
rect 10061 -27189 10099 -27155
rect 10133 -27189 10171 -27155
rect 10205 -27189 10243 -27155
rect 10277 -27189 10315 -27155
rect 10349 -27189 10387 -27155
rect 10421 -27189 10459 -27155
rect 10493 -27189 10531 -27155
rect 10565 -27189 10603 -27155
rect 10637 -27189 10675 -27155
rect 10709 -27189 10747 -27155
rect 10781 -27189 10819 -27155
rect 10853 -27189 10891 -27155
rect 10925 -27189 10963 -27155
rect 10997 -27189 11035 -27155
rect 11069 -27189 11107 -27155
rect 11141 -27189 11179 -27155
rect 11213 -27189 11251 -27155
rect 11285 -27189 11323 -27155
rect 11357 -27189 11395 -27155
rect 11429 -27189 11467 -27155
rect 11501 -27189 11539 -27155
rect 11573 -27189 11611 -27155
rect 11645 -27189 11683 -27155
rect 11717 -27189 11755 -27155
rect 11789 -27189 11827 -27155
rect 11861 -27189 11899 -27155
rect 11933 -27189 11971 -27155
rect 12005 -27189 12043 -27155
rect 12077 -27189 12115 -27155
rect 12149 -27189 12187 -27155
rect 12221 -27189 12259 -27155
rect 12293 -27189 12331 -27155
rect 12365 -27189 12403 -27155
rect 12437 -27189 12475 -27155
rect 12509 -27189 12547 -27155
rect 12581 -27189 12619 -27155
rect 12653 -27189 12691 -27155
rect 12725 -27189 12763 -27155
rect 12797 -27189 12835 -27155
rect 12869 -27189 12907 -27155
rect 12941 -27189 12979 -27155
rect 13013 -27189 13051 -27155
rect 13085 -27189 13123 -27155
rect 13157 -27189 13195 -27155
rect 13229 -27189 13267 -27155
rect 13301 -27189 13339 -27155
rect 13373 -27189 13411 -27155
rect 13445 -27189 13483 -27155
rect 13517 -27189 13555 -27155
rect 13589 -27189 13627 -27155
rect 13661 -27189 13699 -27155
rect 13733 -27189 13771 -27155
rect 13805 -27189 13843 -27155
rect 13877 -27189 13915 -27155
rect 13949 -27189 13987 -27155
rect 14021 -27189 14059 -27155
rect 14093 -27189 14131 -27155
rect 14165 -27189 14203 -27155
rect 14237 -27189 14275 -27155
rect 14309 -27189 14347 -27155
rect 14381 -27189 14419 -27155
rect 14453 -27189 14491 -27155
rect 14525 -27189 14563 -27155
rect 14597 -27189 14635 -27155
rect 14669 -27189 14707 -27155
rect 14741 -27189 14779 -27155
rect 14813 -27189 14851 -27155
rect 14885 -27189 14923 -27155
rect 14957 -27189 14995 -27155
rect 15029 -27189 15067 -27155
rect 15101 -27189 15139 -27155
rect 15173 -27189 15211 -27155
rect 15245 -27189 15283 -27155
rect 15317 -27189 15355 -27155
rect 15389 -27189 15427 -27155
rect 15461 -27189 15499 -27155
rect 15533 -27189 15571 -27155
rect 15605 -27189 15643 -27155
rect 15677 -27189 15715 -27155
rect 15749 -27189 15787 -27155
rect 15821 -27189 15859 -27155
rect 15893 -27189 15931 -27155
rect 15965 -27189 16003 -27155
rect 16037 -27189 16075 -27155
rect 16109 -27189 16147 -27155
rect 16181 -27189 16219 -27155
rect 16253 -27189 16291 -27155
rect 16325 -27189 16363 -27155
rect 16397 -27189 16435 -27155
rect 16469 -27189 16507 -27155
rect 16541 -27189 16579 -27155
rect 16613 -27189 16651 -27155
rect 16685 -27189 16723 -27155
rect 16757 -27189 16795 -27155
rect 16829 -27189 16867 -27155
rect 16901 -27189 16939 -27155
rect 16973 -27189 17011 -27155
rect 17045 -27189 17083 -27155
rect 17117 -27189 17155 -27155
rect 17189 -27189 17227 -27155
rect 17261 -27189 17299 -27155
rect 17333 -27189 17371 -27155
rect 17405 -27189 17443 -27155
rect 17477 -27189 17515 -27155
rect 17549 -27189 17587 -27155
rect 17621 -27189 17659 -27155
rect 17693 -27189 17731 -27155
rect 17765 -27189 17803 -27155
rect 17837 -27189 17875 -27155
rect 17909 -27189 17947 -27155
rect 17981 -27189 18019 -27155
rect 18053 -27189 18091 -27155
rect 18125 -27189 18163 -27155
rect 18197 -27189 18235 -27155
rect 18269 -27189 18307 -27155
rect 18341 -27189 18379 -27155
rect 18413 -27189 18451 -27155
rect 18485 -27189 18523 -27155
rect 18557 -27189 18595 -27155
rect 18629 -27189 18667 -27155
rect 18701 -27189 18739 -27155
rect 18773 -27189 18811 -27155
rect 18845 -27189 18883 -27155
rect 18917 -27189 18955 -27155
rect 18989 -27189 19027 -27155
rect 19061 -27189 19099 -27155
rect 19133 -27189 19171 -27155
rect 19205 -27189 19243 -27155
rect 19277 -27189 19315 -27155
rect 19349 -27189 19387 -27155
rect 19421 -27189 19459 -27155
rect 19493 -27189 19531 -27155
rect 19565 -27189 19603 -27155
rect 19637 -27189 19675 -27155
rect 19709 -27189 19747 -27155
rect 19781 -27189 19819 -27155
rect 19853 -27189 19891 -27155
rect 19925 -27189 19963 -27155
rect 19997 -27189 20035 -27155
rect 20069 -27189 20107 -27155
rect 20141 -27189 20179 -27155
rect 20213 -27189 20251 -27155
rect 20285 -27189 20323 -27155
rect 20357 -27189 20395 -27155
rect 20429 -27189 20467 -27155
rect 20501 -27189 20539 -27155
rect 20573 -27189 20611 -27155
rect 20645 -27189 20683 -27155
rect 20717 -27189 20755 -27155
rect 20789 -27189 20827 -27155
rect 20861 -27189 20899 -27155
rect 20933 -27189 20971 -27155
rect 21005 -27189 21043 -27155
rect 21077 -27189 21115 -27155
rect 21149 -27189 21187 -27155
rect 21221 -27189 21259 -27155
rect 21293 -27189 21331 -27155
rect 21365 -27189 21403 -27155
rect 21437 -27189 21475 -27155
rect 21509 -27189 21547 -27155
rect 21581 -27189 21619 -27155
rect 21653 -27189 21691 -27155
rect 21725 -27189 21763 -27155
rect 21797 -27189 21835 -27155
rect 21869 -27189 21907 -27155
rect 21941 -27189 21979 -27155
rect 22013 -27189 22051 -27155
rect 22085 -27189 22123 -27155
rect 22157 -27189 22195 -27155
rect 22229 -27189 22267 -27155
rect 22301 -27189 22339 -27155
rect 22373 -27189 22411 -27155
rect 22445 -27189 22483 -27155
rect 22517 -27189 22555 -27155
rect 22589 -27189 22627 -27155
rect 22661 -27189 22699 -27155
rect 22733 -27189 22771 -27155
rect 22805 -27189 22843 -27155
rect 22877 -27189 22915 -27155
rect 22949 -27189 22987 -27155
rect 23021 -27189 23059 -27155
rect 23093 -27189 23131 -27155
rect 23165 -27189 23203 -27155
rect 23237 -27189 23275 -27155
rect 23309 -27189 23347 -27155
rect 23381 -27189 23419 -27155
rect 23453 -27189 23491 -27155
rect 23525 -27189 23563 -27155
rect 23597 -27189 23635 -27155
rect 23669 -27189 23707 -27155
rect 23741 -27189 23779 -27155
rect 23813 -27189 23851 -27155
rect 23885 -27189 23923 -27155
rect 23957 -27189 23995 -27155
rect 24029 -27189 24067 -27155
rect 24101 -27189 24139 -27155
rect 24173 -27189 24211 -27155
rect 24245 -27189 24283 -27155
rect 24317 -27189 24355 -27155
rect 24389 -27189 24427 -27155
rect 24461 -27189 24499 -27155
rect 24533 -27189 24571 -27155
rect 24605 -27189 24643 -27155
rect 24677 -27189 24715 -27155
rect 24749 -27189 24787 -27155
rect 24821 -27189 24928 -27155
rect -12328 -27228 24928 -27189
<< via1 >>
rect 502 1344 1066 1588
rect 24134 1344 24698 1588
rect 4075 1037 20831 1217
rect 4160 -4558 4212 -4506
rect 4272 -4558 4324 -4506
rect 4382 -4558 4434 -4506
rect 3496 -5270 3548 -5218
rect 3836 -5270 3888 -5218
rect 3946 -5270 3998 -5218
rect 2114 -6216 2166 -6164
rect 5032 -4558 5084 -4506
rect 5142 -4558 5194 -4506
rect 5250 -4558 5302 -4506
rect 4596 -5270 4648 -5218
rect 4708 -5270 4760 -5218
rect 4816 -5270 4868 -5218
rect 7990 828 8042 880
rect 9072 828 9124 880
rect 10030 828 10082 880
rect 8516 582 8568 634
rect 11066 828 11118 880
rect 12072 828 12124 880
rect 10552 582 10604 634
rect 11570 694 11622 746
rect 13094 828 13146 880
rect 14112 828 14164 880
rect 12590 584 12642 636
rect 15136 828 15188 880
rect 16148 828 16200 880
rect 14620 584 14672 636
rect 17166 828 17218 880
rect 18178 828 18230 880
rect 16662 586 16714 638
rect 17674 694 17726 746
rect 19206 828 19258 880
rect 20218 828 20270 880
rect 18694 586 18746 638
rect 21236 828 21288 880
rect 20730 586 20782 638
rect 6334 -350 6386 -298
rect 7498 -350 7550 -298
rect 6204 -554 6256 -502
rect 7498 -554 7550 -502
rect 9534 -454 9586 -402
rect 11570 -454 11622 -402
rect 13608 -350 13660 -298
rect 13604 -554 13656 -502
rect 15642 -350 15694 -298
rect 15640 -554 15692 -502
rect 17676 -454 17728 -402
rect 17818 -558 17870 -506
rect 19710 -454 19762 -402
rect 19712 -558 19764 -506
rect 21750 -350 21802 -298
rect 22888 -350 22940 -298
rect 8514 -1488 8566 -1436
rect 10550 -1488 10602 -1436
rect 9532 -1584 9584 -1532
rect 10238 -1588 10290 -1536
rect 11410 -1588 11462 -1536
rect 11570 -1694 11622 -1642
rect 12584 -1488 12636 -1436
rect 14622 -1490 14674 -1438
rect 15642 -1588 15694 -1536
rect 16658 -1490 16710 -1438
rect 17676 -1694 17728 -1642
rect 18694 -1490 18746 -1438
rect 19712 -1694 19764 -1642
rect 20728 -1492 20780 -1440
rect 21750 -1588 21802 -1536
rect 8514 -2626 8566 -2574
rect 9532 -2738 9584 -2686
rect 7494 -2876 7546 -2824
rect 6334 -3024 6386 -2972
rect 7316 -3024 7368 -2972
rect 6920 -3360 6972 -3308
rect 6052 -4558 6104 -4506
rect 5468 -5270 5520 -5218
rect 5578 -5270 5630 -5218
rect 4052 -5376 4104 -5324
rect 4488 -5376 4540 -5324
rect 4926 -5376 4978 -5324
rect 5360 -5376 5412 -5324
rect 4272 -5492 4324 -5440
rect 3836 -6216 3888 -6164
rect 5142 -5492 5194 -5440
rect 4052 -6320 4104 -6268
rect 3946 -6418 3998 -6366
rect 4270 -6216 4322 -6164
rect 4160 -6418 4212 -6366
rect 4488 -6320 4540 -6268
rect 4380 -6418 4432 -6366
rect 3496 -7054 3548 -7002
rect 4706 -6216 4758 -6164
rect 5936 -5492 5988 -5440
rect 4926 -6320 4978 -6268
rect 4598 -6418 4650 -6366
rect 4708 -6418 4760 -6366
rect 4814 -6418 4866 -6366
rect 3836 -7154 3888 -7102
rect 5142 -6216 5194 -6164
rect 5032 -6418 5084 -6366
rect 5360 -6320 5412 -6268
rect 5250 -6418 5302 -6366
rect 5580 -6216 5632 -6164
rect 5466 -6418 5518 -6366
rect 4706 -7154 4758 -7102
rect 5580 -7154 5632 -7102
rect 5936 -7154 5988 -7102
rect 4052 -7252 4104 -7200
rect 4488 -7252 4540 -7200
rect 4926 -7252 4978 -7200
rect 5360 -7252 5412 -7200
rect 3496 -7370 3548 -7318
rect 4162 -7370 4214 -7318
rect 4270 -7370 4322 -7318
rect 4378 -7370 4430 -7318
rect 5024 -7370 5076 -7318
rect 5142 -7370 5194 -7318
rect 5250 -7371 5302 -7319
rect 6806 -5664 6858 -5612
rect 10550 -2626 10602 -2574
rect 9532 -3172 9584 -3120
rect 7316 -3460 7368 -3408
rect 8482 -3460 8534 -3408
rect 7048 -4506 7100 -4454
rect 6920 -5768 6972 -5716
rect 3836 -8090 3888 -8038
rect 3946 -8090 3998 -8038
rect 4600 -8090 4652 -8038
rect 4706 -8090 4758 -8038
rect 4816 -8090 4868 -8038
rect 5468 -8090 5520 -8038
rect 5580 -8090 5632 -8038
rect 6052 -8090 6104 -8038
rect 7184 -4604 7236 -4552
rect 7048 -8178 7100 -8126
rect 12044 -2630 12096 -2578
rect 11568 -3360 11620 -3308
rect 10518 -3460 10570 -3408
rect 12568 -2627 12620 -2575
rect 13044 -2626 13096 -2574
rect 8486 -4714 8538 -4662
rect 9500 -4408 9552 -4356
rect 9500 -4604 9552 -4552
rect 10520 -4602 10572 -4550
rect 10520 -4714 10572 -4662
rect 14088 -2624 14140 -2572
rect 13604 -2876 13656 -2824
rect 13604 -3160 13656 -3108
rect 14606 -2626 14658 -2574
rect 15104 -2624 15156 -2572
rect 16132 -2624 16184 -2572
rect 15640 -2876 15692 -2824
rect 16642 -2629 16694 -2577
rect 17154 -2634 17206 -2582
rect 17642 -2630 17694 -2578
rect 18154 -2634 18206 -2582
rect 18694 -2630 18746 -2578
rect 20728 -2630 20780 -2578
rect 19712 -2738 19764 -2686
rect 21748 -2876 21800 -2824
rect 21718 -3154 21770 -3102
rect 22888 -3160 22940 -3108
rect 18664 -3460 18716 -3408
rect 20698 -3460 20750 -3408
rect 23142 -3460 23194 -3408
rect 11536 -4408 11588 -4356
rect 13576 -4716 13628 -4664
rect 15610 -4716 15662 -4664
rect 18666 -4716 18718 -4664
rect 19680 -4408 19732 -4356
rect 20700 -4716 20752 -4664
rect 21716 -4408 21768 -4356
rect 22982 -4602 23034 -4550
rect 9502 -5768 9554 -5716
rect 9502 -5972 9554 -5920
rect 13572 -5664 13624 -5612
rect 11538 -5768 11590 -5716
rect 11536 -5870 11588 -5818
rect 11536 -5972 11588 -5920
rect 14592 -5664 14644 -5612
rect 14592 -5970 14644 -5918
rect 15610 -5970 15662 -5918
rect 16628 -5664 16680 -5612
rect 16626 -5970 16678 -5918
rect 18662 -5768 18714 -5716
rect 19530 -5650 19582 -5598
rect 19678 -5760 19730 -5708
rect 19530 -5970 19582 -5918
rect 19682 -5968 19734 -5916
rect 20698 -5870 20750 -5818
rect 21718 -5760 21770 -5708
rect 22850 -5760 22902 -5708
rect 21716 -5968 21768 -5916
rect 8484 -6920 8536 -6868
rect 7316 -7128 7368 -7076
rect 9498 -7230 9550 -7178
rect 10520 -6920 10572 -6868
rect 10520 -7028 10572 -6976
rect 11532 -7230 11584 -7178
rect 11736 -7224 11788 -7172
rect 13574 -6918 13626 -6866
rect 15610 -6918 15662 -6866
rect 18664 -6916 18716 -6864
rect 13570 -7224 13622 -7172
rect 14590 -7228 14642 -7176
rect 16624 -7228 16676 -7176
rect 16838 -7232 16890 -7180
rect 19174 -7232 19226 -7180
rect 19686 -7230 19738 -7178
rect 20700 -6916 20752 -6864
rect 22982 -5968 23034 -5916
rect 22850 -7028 22902 -6976
rect 21720 -7230 21772 -7178
rect 8480 -8178 8532 -8126
rect 10516 -8178 10568 -8126
rect 7184 -8308 7236 -8256
rect 2114 -8448 2166 -8396
rect 1958 -8554 2010 -8502
rect 18668 -8178 18720 -8126
rect 20704 -8178 20756 -8126
rect 11538 -8448 11590 -8396
rect 23142 -8448 23194 -8396
rect 1188 -8672 1240 -8620
rect -12008 -11211 -11956 -11202
rect -10214 -11211 -10162 -11202
rect -7614 -11211 -7562 -11202
rect -5014 -11211 -4962 -11200
rect -2414 -11211 -2362 -11200
rect -610 -11211 -558 -11200
rect -12008 -11245 -12005 -11211
rect -12005 -11245 -11971 -11211
rect -11971 -11245 -11956 -11211
rect -10214 -11245 -10205 -11211
rect -10205 -11245 -10171 -11211
rect -10171 -11245 -10162 -11211
rect -7614 -11245 -7613 -11211
rect -7613 -11245 -7579 -11211
rect -7579 -11245 -7562 -11211
rect -5014 -11245 -4987 -11211
rect -4987 -11245 -4962 -11211
rect -2414 -11245 -2395 -11211
rect -2395 -11245 -2362 -11211
rect -610 -11245 -595 -11211
rect -595 -11245 -558 -11211
rect -12008 -11254 -11956 -11245
rect -10214 -11254 -10162 -11245
rect -7614 -11254 -7562 -11245
rect -5014 -11252 -4962 -11245
rect -2414 -11252 -2362 -11245
rect -610 -11252 -558 -11245
rect 1958 -11404 2010 -11352
rect 2114 -11404 2166 -11352
rect 1188 -12390 1240 -12338
rect 1854 -12504 1906 -12452
rect 2340 -11412 2392 -11360
rect 2116 -13844 2168 -13792
rect 1980 -14056 2032 -14004
rect 1854 -14958 1906 -14906
rect 694 -18944 746 -18892
rect -2972 -20216 -2920 -20164
rect -7382 -21656 -7330 -21604
rect -5342 -21656 -5290 -21604
rect -9534 -22560 -9482 -22508
rect -8396 -22560 -8344 -22508
rect -7382 -22656 -7330 -22604
rect -6360 -22772 -6308 -22720
rect -5342 -22656 -5290 -22604
rect -4322 -22560 -4270 -22508
rect -810 -19180 -758 -19128
rect 102 -19180 154 -19128
rect -1680 -19290 -1628 -19238
rect -2594 -19398 -2542 -19346
rect -2464 -19506 -2412 -19454
rect -916 -19398 -864 -19346
rect -1134 -19506 -1082 -19454
rect -2006 -20006 -1954 -19954
rect -18 -19290 34 -19238
rect -698 -19398 -646 -19346
rect -480 -19506 -428 -19454
rect -1898 -20106 -1846 -20054
rect -1896 -20216 -1844 -20164
rect -1350 -20006 -1298 -19954
rect -1460 -20106 -1408 -20054
rect -1462 -20216 -1410 -20164
rect -1788 -20326 -1736 -20274
rect -1568 -20326 -1516 -20274
rect -2464 -20830 -2412 -20778
rect -2594 -20952 -2542 -20900
rect -2006 -20830 -1954 -20778
rect -1788 -20952 -1736 -20900
rect -2114 -21076 -2062 -21024
rect -480 -20006 -428 -19954
rect -1134 -20216 -1082 -20164
rect -1024 -20216 -972 -20164
rect -588 -20216 -536 -20164
rect -914 -20326 -862 -20274
rect -698 -20326 -646 -20274
rect -1350 -20830 -1298 -20778
rect -1570 -20952 -1518 -20900
rect -1676 -21202 -1624 -21150
rect -18 -19780 34 -19728
rect -370 -20126 -318 -20074
rect -806 -20830 -754 -20778
rect -1134 -20950 -1082 -20898
rect -478 -20950 -426 -20898
rect -18 -20830 34 -20778
rect -1244 -21076 -1192 -21024
rect -372 -21076 -320 -21024
rect 224 -20006 276 -19954
rect 224 -20252 276 -20200
rect 102 -21202 154 -21150
rect -1346 -21312 -1294 -21260
rect 956 -18914 1008 -18862
rect -2666 -21636 -2614 -21584
rect -8250 -23672 -8198 -23620
rect -8398 -23780 -8346 -23728
rect -3198 -22772 -3146 -22720
rect -7380 -23892 -7328 -23840
rect -6364 -23672 -6312 -23620
rect -6362 -23780 -6310 -23728
rect -5342 -23892 -5290 -23840
rect -4494 -23672 -4442 -23620
rect -4326 -23780 -4274 -23728
rect -8396 -24876 -8344 -24824
rect -9534 -24982 -9482 -24930
rect -7378 -24774 -7326 -24722
rect -6362 -24982 -6310 -24930
rect -5348 -24774 -5296 -24722
rect -7892 -25926 -7840 -25874
rect -2118 -21536 -2066 -21484
rect -928 -21536 -876 -21484
rect 266 -21536 318 -21484
rect 956 -21536 1008 -21484
rect -1674 -21636 -1622 -21584
rect -1376 -21636 -1324 -21584
rect -480 -21636 -428 -21584
rect -184 -21636 -132 -21584
rect -2538 -22670 -2486 -22618
rect -2122 -22670 -2070 -22618
rect -1826 -22538 -1774 -22486
rect -1970 -22778 -1918 -22726
rect -1222 -22538 -1170 -22486
rect -1528 -22670 -1476 -22618
rect -1672 -22778 -1620 -22726
rect -1372 -22778 -1320 -22726
rect -930 -22670 -878 -22618
rect -1078 -22778 -1026 -22726
rect -631 -22538 -579 -22486
rect -782 -22778 -730 -22726
rect -34 -22538 18 -22486
rect -336 -22670 -284 -22618
rect -482 -22778 -430 -22726
rect -180 -22778 -128 -22726
rect -2666 -23676 -2614 -23624
rect -4328 -24876 -4276 -24824
rect -3198 -24876 -3146 -24824
rect -6866 -25926 -6814 -25874
rect -5842 -25926 -5790 -25874
rect -1972 -23676 -1920 -23624
rect 262 -22670 314 -22618
rect 110 -22778 162 -22726
rect 562 -22538 614 -22486
rect 414 -22778 466 -22726
rect -1526 -23784 -1474 -23732
rect -1076 -23676 -1024 -23624
rect -782 -23676 -730 -23624
rect -332 -23784 -280 -23732
rect -1824 -24768 -1772 -24716
rect -2422 -24862 -2370 -24810
rect -1974 -24970 -1922 -24918
rect -1530 -24862 -1478 -24810
rect -1676 -24970 -1624 -24918
rect 112 -23676 164 -23624
rect 414 -23676 466 -23624
rect -1230 -24768 -1178 -24716
rect -1380 -24970 -1328 -24918
rect -630 -24768 -578 -24716
rect -932 -24862 -880 -24810
rect -1076 -24970 -1024 -24918
rect -780 -24970 -728 -24918
rect -334 -24862 -282 -24810
rect -482 -24970 -430 -24918
rect 956 -23784 1008 -23732
rect -36 -24768 16 -24716
rect -186 -24970 -134 -24918
rect 558 -24768 610 -24716
rect 266 -24862 318 -24810
rect 110 -24970 162 -24918
rect 414 -24970 466 -24918
rect -4942 -25926 -4890 -25874
rect -2666 -25896 -2614 -25844
rect -1676 -25896 -1624 -25844
rect -1378 -25896 -1326 -25844
rect -482 -25896 -430 -25844
rect -180 -25896 -128 -25844
rect 1080 -22778 1132 -22726
rect 1980 -23600 2032 -23548
rect 2572 -12504 2624 -12452
rect 3590 -12602 3642 -12550
rect 4608 -12504 4660 -12452
rect 6642 -12504 6694 -12452
rect 8682 -12504 8734 -12452
rect 10718 -12504 10770 -12452
rect 12752 -12504 12804 -12452
rect 14788 -12504 14840 -12452
rect 16824 -12504 16876 -12452
rect 18860 -12504 18912 -12452
rect 5628 -12602 5680 -12550
rect 7662 -12602 7714 -12550
rect 9696 -12602 9748 -12550
rect 11736 -12602 11788 -12550
rect 13770 -12602 13822 -12550
rect 15808 -12602 15860 -12550
rect 17840 -12602 17892 -12550
rect 19878 -12602 19930 -12550
rect 11736 -12814 11788 -12762
rect 13768 -12814 13820 -12762
rect 6276 -13734 6328 -13682
rect 6646 -13734 6698 -13682
rect 7148 -13734 7200 -13682
rect 7660 -13734 7712 -13682
rect 8188 -13734 8240 -13682
rect 8680 -13734 8732 -13682
rect 4100 -13844 4152 -13792
rect 5122 -13844 5174 -13792
rect 2576 -14056 2628 -14004
rect 3074 -14056 3126 -14004
rect 3586 -14056 3638 -14004
rect 6142 -13948 6194 -13896
rect 5628 -14056 5680 -14004
rect 4090 -14958 4142 -14906
rect 2340 -15172 2392 -15120
rect 7142 -13948 7194 -13896
rect 8162 -13948 8214 -13896
rect 7662 -14056 7714 -14004
rect 10712 -13734 10764 -13682
rect 9194 -13844 9246 -13792
rect 9698 -13844 9750 -13792
rect 10214 -13844 10266 -13792
rect 9696 -14056 9748 -14004
rect 5106 -14946 5158 -14894
rect 6126 -14946 6178 -14894
rect 4602 -15050 4654 -14998
rect 4608 -15284 4660 -15232
rect 5626 -15050 5678 -14998
rect 11234 -13844 11286 -13792
rect 11736 -13844 11788 -13792
rect 12236 -13844 12288 -13792
rect 11852 -14056 11904 -14004
rect 12748 -13734 12800 -13682
rect 12376 -13948 12428 -13896
rect 13262 -13844 13314 -13792
rect 13384 -13948 13436 -13896
rect 13772 -13844 13824 -13792
rect 14280 -13844 14332 -13792
rect 13576 -14058 13628 -14006
rect 20898 -12504 20950 -12452
rect 14784 -13734 14836 -13682
rect 14426 -13948 14478 -13896
rect 7138 -14946 7190 -14894
rect 8164 -14946 8216 -14894
rect 6638 -15050 6690 -14998
rect 6644 -15284 6696 -15232
rect 7658 -15050 7710 -14998
rect 16822 -13734 16874 -13682
rect 15288 -13844 15340 -13792
rect 15810 -13844 15862 -13792
rect 16300 -13844 16352 -13792
rect 15810 -14056 15862 -14004
rect 21916 -12602 21968 -12550
rect 22928 -12504 22980 -12452
rect 23652 -12602 23704 -12550
rect 18346 -13734 18398 -13682
rect 18860 -13734 18912 -13682
rect 19368 -13734 19420 -13682
rect 17332 -13844 17384 -13792
rect 17844 -13844 17896 -13792
rect 17318 -13948 17370 -13896
rect 18356 -13948 18408 -13896
rect 17842 -14056 17894 -14004
rect 8680 -15050 8732 -14998
rect 10716 -15050 10768 -14998
rect 12754 -15050 12806 -14998
rect 14784 -15050 14836 -14998
rect 9700 -15172 9752 -15120
rect 11734 -15172 11786 -15120
rect 13764 -15172 13816 -15120
rect 2452 -16214 2504 -16162
rect 3590 -16214 3642 -16162
rect 2340 -16414 2392 -16362
rect 2234 -16516 2286 -16464
rect 2340 -17650 2392 -17598
rect 2234 -20006 2286 -19954
rect 3588 -16414 3640 -16362
rect 4606 -16294 4658 -16242
rect 5624 -16190 5676 -16138
rect 5120 -16408 5172 -16356
rect 6646 -16294 6698 -16242
rect 6124 -16408 6176 -16356
rect 7660 -16190 7712 -16138
rect 7136 -16408 7188 -16356
rect 3588 -17446 3640 -17394
rect 4094 -17548 4146 -17496
rect 8678 -16294 8730 -16242
rect 15804 -15050 15856 -14998
rect 8156 -16408 8208 -16356
rect 8678 -16406 8730 -16354
rect 10712 -16294 10764 -16242
rect 9696 -16516 9748 -16464
rect 10714 -16406 10766 -16354
rect 11730 -16516 11782 -16464
rect 5626 -17446 5678 -17394
rect 5624 -17650 5676 -17598
rect 20388 -13844 20440 -13792
rect 21408 -13844 21460 -13792
rect 19356 -13948 19408 -13896
rect 19874 -14056 19926 -14004
rect 21916 -14056 21968 -14004
rect 22420 -14056 22472 -14004
rect 22930 -14056 22982 -14004
rect 17320 -14946 17372 -14894
rect 18356 -14946 18408 -14894
rect 16822 -15050 16874 -14998
rect 17842 -15050 17894 -14998
rect 12752 -16294 12804 -16242
rect 19372 -14946 19424 -14894
rect 18858 -15050 18910 -14998
rect 20894 -15050 20946 -14998
rect 12750 -16406 12802 -16354
rect 14786 -16294 14838 -16242
rect 14982 -16298 15034 -16246
rect 13770 -16516 13822 -16464
rect 14786 -16406 14838 -16354
rect 15804 -16190 15856 -16138
rect 14982 -16516 15034 -16464
rect 15276 -16514 15328 -16462
rect 16820 -16406 16872 -16354
rect 16304 -16514 16356 -16462
rect 16822 -16520 16874 -16468
rect 7662 -17446 7714 -17394
rect 4608 -17750 4660 -17698
rect 6132 -17656 6184 -17604
rect 7154 -17656 7206 -17604
rect 6642 -17750 6694 -17698
rect 9694 -17446 9746 -17394
rect 9186 -17548 9238 -17496
rect 8168 -17656 8220 -17604
rect 9186 -17656 9238 -17604
rect 8678 -17750 8730 -17698
rect 4090 -18674 4142 -18622
rect 5000 -18674 5052 -18622
rect 4090 -18890 4142 -18838
rect 2454 -18994 2506 -18942
rect 2340 -20252 2392 -20200
rect 2242 -21312 2294 -21260
rect 6002 -18674 6054 -18622
rect 5128 -18890 5180 -18838
rect 7154 -18674 7206 -18622
rect 6642 -18776 6694 -18724
rect 6142 -18890 6194 -18838
rect 10206 -17656 10258 -17604
rect 17840 -16190 17892 -16138
rect 18858 -16406 18910 -16354
rect 23038 -15284 23090 -15232
rect 19874 -16298 19926 -16246
rect 20378 -16302 20430 -16250
rect 20898 -16406 20950 -16354
rect 18858 -16520 18910 -16468
rect 20896 -16520 20948 -16468
rect 14276 -17434 14328 -17382
rect 13770 -17562 13822 -17510
rect 15806 -17760 15858 -17708
rect 8164 -18674 8216 -18622
rect 9170 -18674 9222 -18622
rect 10214 -18674 10266 -18622
rect 10714 -18668 10766 -18616
rect 9168 -18890 9220 -18838
rect 10208 -18890 10260 -18838
rect 9692 -18994 9744 -18942
rect 4088 -19902 4140 -19850
rect 3590 -20006 3642 -19954
rect 3586 -20216 3638 -20164
rect 5096 -19902 5148 -19850
rect 4606 -20118 4658 -20066
rect 6110 -19902 6162 -19850
rect 11222 -18890 11274 -18838
rect 12750 -18668 12802 -18616
rect 12230 -18890 12282 -18838
rect 13274 -18890 13326 -18838
rect 11734 -18994 11786 -18942
rect 21914 -16190 21966 -16138
rect 22932 -16172 22984 -16120
rect 23532 -16302 23584 -16250
rect 23282 -16406 23334 -16354
rect 17318 -17656 17370 -17604
rect 19370 -17434 19422 -17382
rect 19508 -17430 19560 -17378
rect 23038 -16520 23090 -16468
rect 20390 -17430 20442 -17378
rect 21396 -17430 21448 -17378
rect 21914 -17434 21966 -17382
rect 18348 -17656 18400 -17604
rect 19508 -17656 19560 -17604
rect 19876 -17656 19928 -17604
rect 19876 -17760 19928 -17708
rect 21914 -17562 21966 -17510
rect 20892 -17758 20944 -17706
rect 14786 -18668 14838 -18616
rect 14264 -18890 14316 -18838
rect 15282 -18890 15334 -18838
rect 13772 -18994 13824 -18942
rect 7148 -19902 7200 -19850
rect 6644 -20118 6696 -20066
rect 5624 -20216 5676 -20164
rect 8166 -19902 8218 -19850
rect 8682 -19896 8734 -19844
rect 16824 -18668 16876 -18616
rect 16816 -18776 16868 -18724
rect 16316 -18890 16368 -18838
rect 15806 -18994 15858 -18942
rect 16318 -18998 16370 -18946
rect 17340 -18998 17392 -18946
rect 17840 -18992 17892 -18940
rect 18860 -18668 18912 -18616
rect 18856 -18776 18908 -18724
rect 19348 -18890 19400 -18838
rect 20898 -18668 20950 -18616
rect 20894 -18776 20946 -18724
rect 20386 -18890 20438 -18838
rect 19874 -18992 19926 -18940
rect 21412 -18890 21464 -18838
rect 21916 -18992 21968 -18940
rect 10718 -19896 10770 -19844
rect 7664 -20216 7716 -20164
rect 2452 -21238 2504 -21186
rect 3592 -21454 3644 -21402
rect 12750 -19896 12802 -19844
rect 14784 -19896 14836 -19844
rect 11734 -20006 11786 -19954
rect 13770 -20006 13822 -19954
rect 10716 -20118 10768 -20066
rect 9700 -20216 9752 -20164
rect 4606 -21140 4658 -21088
rect 4610 -21334 4662 -21282
rect 5624 -21238 5676 -21186
rect 6642 -21140 6694 -21088
rect 7148 -21238 7200 -21186
rect 6646 -21334 6698 -21282
rect 8680 -21140 8732 -21088
rect 8170 -21238 8222 -21186
rect 7660 -21454 7712 -21402
rect 9192 -21238 9244 -21186
rect 8674 -21334 8726 -21282
rect 15806 -19894 15858 -19842
rect 16160 -19894 16212 -19842
rect 15802 -20006 15854 -19954
rect 15312 -20104 15364 -20052
rect 10542 -21120 10594 -21068
rect 10196 -21238 10248 -21186
rect 9694 -21454 9746 -21402
rect 10712 -21120 10764 -21068
rect 10542 -21334 10594 -21282
rect 10718 -21328 10770 -21276
rect 16350 -20104 16402 -20052
rect 17326 -20104 17378 -20052
rect 19878 -19894 19930 -19842
rect 18342 -20104 18394 -20052
rect 20368 -20104 20420 -20052
rect 16160 -20212 16212 -20160
rect 17840 -20216 17892 -20164
rect 19876 -20216 19928 -20164
rect 12754 -21120 12806 -21068
rect 14786 -21120 14838 -21068
rect 21398 -20104 21450 -20052
rect 21912 -20216 21964 -20164
rect 16826 -21120 16878 -21068
rect 15804 -21218 15856 -21166
rect 12746 -21328 12798 -21276
rect 2340 -22370 2392 -22318
rect 2234 -22496 2286 -22444
rect 5624 -22496 5676 -22444
rect 6144 -22484 6196 -22432
rect 4606 -22606 4658 -22554
rect 6642 -22606 6694 -22554
rect 6260 -22700 6312 -22648
rect 7662 -22606 7714 -22554
rect 14790 -21328 14842 -21276
rect 8678 -22606 8730 -22554
rect 9698 -22606 9750 -22554
rect 7144 -22700 7196 -22648
rect 8166 -22700 8218 -22648
rect 2572 -23600 2624 -23548
rect 3086 -23600 3138 -23548
rect 3584 -23600 3636 -23548
rect 5626 -23600 5678 -23548
rect 6134 -23712 6186 -23660
rect 2114 -23818 2166 -23766
rect 4100 -23818 4152 -23766
rect 5122 -23818 5174 -23766
rect 16818 -21328 16870 -21276
rect 17844 -21454 17896 -21402
rect 18856 -21328 18908 -21276
rect 19874 -21454 19926 -21402
rect 21910 -21218 21962 -21166
rect 20896 -21328 20948 -21276
rect 21414 -21324 21466 -21272
rect 20400 -21452 20452 -21400
rect 21912 -21452 21964 -21400
rect 11728 -22370 11780 -22318
rect 13770 -22370 13822 -22318
rect 15806 -22370 15858 -22318
rect 11224 -22484 11276 -22432
rect 16312 -22480 16364 -22428
rect 10716 -22606 10768 -22554
rect 12746 -22606 12798 -22554
rect 14784 -22606 14836 -22554
rect 16820 -22606 16872 -22554
rect 10208 -22700 10260 -22648
rect 7658 -23600 7710 -23548
rect 7146 -23712 7198 -23660
rect 8160 -23712 8212 -23660
rect 7660 -23818 7712 -23766
rect 8172 -23818 8224 -23766
rect 1708 -23922 1760 -23870
rect 6136 -23922 6188 -23870
rect 6640 -23922 6692 -23870
rect 7156 -23922 7208 -23870
rect 1080 -24970 1132 -24918
rect -2122 -25996 -2070 -25944
rect -934 -25996 -882 -25944
rect 262 -25996 314 -25944
rect 956 -25996 1008 -25944
rect 2572 -25152 2624 -25100
rect 9690 -23600 9742 -23548
rect 9190 -23818 9242 -23766
rect 9696 -23818 9748 -23766
rect 10202 -23818 10254 -23766
rect 8678 -23922 8730 -23870
rect 3584 -25054 3636 -25002
rect 11072 -23712 11124 -23660
rect 10716 -23922 10768 -23870
rect 4602 -25152 4654 -25100
rect 11594 -23600 11646 -23548
rect 11214 -23818 11266 -23766
rect 11732 -23710 11784 -23658
rect 12360 -23714 12412 -23662
rect 12234 -23818 12286 -23766
rect 17842 -22606 17894 -22554
rect 18860 -22370 18912 -22318
rect 18862 -22606 18914 -22554
rect 17330 -22700 17382 -22648
rect 18350 -22700 18402 -22648
rect 13406 -23714 13458 -23662
rect 13256 -23818 13308 -23766
rect 12752 -23922 12804 -23870
rect 19876 -22606 19928 -22554
rect 20892 -22370 20944 -22318
rect 23166 -17434 23218 -17382
rect 23404 -17656 23456 -17604
rect 23282 -17758 23334 -17706
rect 23166 -18992 23218 -18940
rect 23162 -19894 23214 -19842
rect 23282 -21120 23334 -21068
rect 23162 -21218 23214 -21166
rect 23530 -18890 23582 -18838
rect 23532 -21324 23584 -21272
rect 23404 -21452 23456 -21400
rect 23038 -22370 23090 -22318
rect 21412 -22480 21464 -22428
rect 20898 -22606 20950 -22554
rect 19364 -22700 19416 -22648
rect 20400 -22700 20452 -22648
rect 13954 -23598 14006 -23546
rect 13768 -23818 13820 -23766
rect 14274 -23818 14326 -23766
rect 15804 -23600 15856 -23548
rect 15292 -23818 15344 -23766
rect 15804 -23818 15856 -23766
rect 16312 -23818 16364 -23766
rect 14788 -23922 14840 -23870
rect 17838 -23600 17890 -23548
rect 17334 -23714 17386 -23662
rect 18352 -23714 18404 -23662
rect 19872 -23600 19924 -23548
rect 19362 -23714 19414 -23662
rect 16820 -23922 16872 -23870
rect 17342 -23922 17394 -23870
rect 17842 -23922 17894 -23870
rect 18350 -23922 18402 -23870
rect 18858 -23922 18910 -23870
rect 19208 -23922 19260 -23870
rect 21914 -23600 21966 -23548
rect 22426 -23600 22478 -23548
rect 22932 -23600 22984 -23548
rect 20384 -23818 20436 -23766
rect 21386 -23818 21438 -23766
rect 11734 -24854 11786 -24802
rect 13770 -24854 13822 -24802
rect 5622 -25054 5674 -25002
rect 7660 -25054 7712 -25002
rect 9692 -25054 9744 -25002
rect 11730 -25054 11782 -25002
rect 13764 -25054 13816 -25002
rect 15804 -25054 15856 -25002
rect 17838 -25054 17890 -25002
rect 19872 -25054 19924 -25002
rect 6640 -25152 6692 -25100
rect 8676 -25152 8728 -25100
rect 10712 -25152 10764 -25100
rect 12748 -25152 12800 -25100
rect 14782 -25152 14834 -25100
rect 16818 -25152 16870 -25100
rect 18858 -25152 18910 -25100
rect 20892 -25152 20944 -25100
rect 21910 -25054 21962 -25002
rect 23810 -23922 23862 -23870
rect 23652 -25054 23704 -25002
rect 22928 -25152 22980 -25100
rect -7446 -26611 23902 -26495
rect -12198 -27088 -11634 -26844
rect 24234 -27088 24798 -26844
<< metal2 >>
rect 484 1614 1084 1626
rect 484 1588 516 1614
rect 1052 1588 1084 1614
rect 484 1344 502 1588
rect 1066 1344 1084 1588
rect 484 1318 516 1344
rect 1052 1318 1084 1344
rect 484 1306 1084 1318
rect 24116 1614 24716 1626
rect 24116 1588 24148 1614
rect 24684 1588 24716 1614
rect 24116 1344 24134 1588
rect 24698 1344 24716 1588
rect 24116 1318 24148 1344
rect 24684 1318 24716 1344
rect 24116 1306 24716 1318
rect 3998 1217 20878 1266
rect 3998 1195 4075 1217
rect 20831 1195 20878 1217
rect 3998 1059 4065 1195
rect 20841 1059 20878 1195
rect 3998 1037 4075 1059
rect 20831 1037 20878 1059
rect 3998 1000 20878 1037
rect 3998 998 8352 1000
rect 7986 884 8046 890
rect 9068 884 9128 890
rect 10026 884 10086 890
rect 11062 884 11122 890
rect 12068 884 12128 890
rect 13090 884 13150 890
rect 14108 884 14168 890
rect 15132 884 15192 890
rect 16144 884 16204 890
rect 17162 884 17222 890
rect 18174 884 18234 890
rect 19202 884 19262 890
rect 20214 884 20274 890
rect 21232 884 21292 890
rect 7986 880 21292 884
rect 7986 828 7990 880
rect 8042 828 9072 880
rect 9124 828 10030 880
rect 10082 828 11066 880
rect 11118 828 12072 880
rect 12124 828 13094 880
rect 13146 828 14112 880
rect 14164 828 15136 880
rect 15188 828 16148 880
rect 16200 828 17166 880
rect 17218 828 18178 880
rect 18230 828 19206 880
rect 19258 828 20218 880
rect 20270 828 21236 880
rect 21288 828 21292 880
rect 7986 824 21292 828
rect 7986 818 8046 824
rect 9068 818 9128 824
rect 10026 818 10086 824
rect 11062 818 11122 824
rect 12068 818 12128 824
rect 13090 818 13150 824
rect 14108 818 14168 824
rect 15132 818 15192 824
rect 16144 818 16204 824
rect 17162 818 17222 824
rect 18174 818 18234 824
rect 19202 818 19262 824
rect 20214 818 20274 824
rect 21232 818 21292 824
rect 11566 750 11626 756
rect 17670 750 17730 756
rect 11566 746 17730 750
rect 11566 694 11570 746
rect 11622 694 17674 746
rect 17726 694 17730 746
rect 11566 690 17730 694
rect 11566 684 11626 690
rect 17670 684 17730 690
rect 8512 638 8572 644
rect 10548 638 10608 644
rect 12586 640 12646 646
rect 14616 640 14676 646
rect 16658 642 16718 648
rect 18690 642 18750 648
rect 20726 642 20786 648
rect 16658 640 20786 642
rect 12586 638 20786 640
rect 8512 636 16662 638
rect 8512 634 12590 636
rect 8512 582 8516 634
rect 8568 582 10552 634
rect 10604 584 12590 634
rect 12642 584 14620 636
rect 14672 586 16662 636
rect 16714 586 18694 638
rect 18746 586 20730 638
rect 20782 586 20786 638
rect 14672 584 20786 586
rect 10604 582 20786 584
rect 8512 580 16856 582
rect 8512 578 12768 580
rect 8512 572 8572 578
rect 10548 572 10608 578
rect 12586 574 12646 578
rect 14616 574 14676 580
rect 16658 576 16718 580
rect 18690 576 18750 582
rect 20726 576 20786 582
rect 6330 -294 6390 -288
rect 7494 -294 7554 -288
rect 13604 -294 13664 -288
rect 6330 -298 13664 -294
rect 6330 -350 6334 -298
rect 6386 -350 7498 -298
rect 7550 -350 13608 -298
rect 13660 -350 13664 -298
rect 6330 -354 13664 -350
rect 6330 -360 6390 -354
rect 7494 -360 7554 -354
rect 13604 -360 13664 -354
rect 15638 -294 15698 -288
rect 21746 -294 21806 -288
rect 22884 -294 22944 -288
rect 15638 -298 22944 -294
rect 15638 -350 15642 -298
rect 15694 -350 21750 -298
rect 21802 -350 22888 -298
rect 22940 -350 22944 -298
rect 15638 -354 22944 -350
rect 15638 -360 15698 -354
rect 21746 -360 21806 -354
rect 22884 -360 22944 -354
rect 9530 -398 9590 -392
rect 11566 -398 11626 -392
rect 17672 -398 17732 -392
rect 19706 -398 19766 -392
rect 9530 -402 12044 -398
rect 9530 -454 9534 -402
rect 9586 -454 11570 -402
rect 11622 -406 12044 -402
rect 12260 -402 19766 -398
rect 12260 -406 17676 -402
rect 11622 -452 17676 -406
rect 11622 -454 14060 -452
rect 9530 -456 14060 -454
rect 9530 -458 13034 -456
rect 13272 -458 14060 -456
rect 14276 -454 17676 -452
rect 17728 -454 19710 -402
rect 19762 -454 19766 -402
rect 14276 -458 19766 -454
rect 9530 -464 9590 -458
rect 11566 -464 11626 -458
rect 17672 -464 17732 -458
rect 19706 -464 19766 -458
rect 6200 -498 6260 -492
rect 7494 -498 7554 -492
rect 13600 -498 13660 -492
rect 15636 -498 15696 -492
rect 6200 -502 15696 -498
rect 6200 -554 6204 -502
rect 6256 -554 7498 -502
rect 7550 -554 13604 -502
rect 13656 -554 15640 -502
rect 15692 -554 15696 -502
rect 6200 -558 15696 -554
rect 6200 -564 6260 -558
rect 7494 -564 7554 -558
rect 13600 -564 13660 -558
rect 15636 -564 15696 -558
rect 17814 -502 17874 -496
rect 19708 -502 19768 -496
rect 17814 -506 19768 -502
rect 17814 -558 17818 -506
rect 17870 -558 19712 -506
rect 19764 -558 19768 -506
rect 17814 -562 19768 -558
rect 17814 -568 17874 -562
rect 19708 -568 19768 -562
rect 8510 -1432 8570 -1426
rect 10546 -1432 10606 -1426
rect 12580 -1432 12640 -1426
rect 14618 -1432 14678 -1428
rect 8510 -1434 14822 -1432
rect 16654 -1434 16714 -1428
rect 18690 -1434 18750 -1428
rect 8510 -1436 19560 -1434
rect 20724 -1436 20784 -1430
rect 8510 -1488 8514 -1436
rect 8566 -1488 10550 -1436
rect 10602 -1488 12584 -1436
rect 12636 -1438 20784 -1436
rect 12636 -1488 14622 -1438
rect 8510 -1490 14622 -1488
rect 14674 -1490 16658 -1438
rect 16710 -1490 18694 -1438
rect 18746 -1440 20784 -1438
rect 18746 -1490 20728 -1440
rect 8510 -1492 20728 -1490
rect 20780 -1492 20784 -1440
rect 8510 -1498 8570 -1492
rect 10546 -1498 10606 -1492
rect 12580 -1498 12640 -1492
rect 14618 -1494 20784 -1492
rect 14618 -1500 14678 -1494
rect 16654 -1500 16714 -1494
rect 18589 -1496 19104 -1494
rect 19354 -1496 20784 -1494
rect 18690 -1500 18750 -1496
rect 20724 -1502 20784 -1496
rect 9528 -1528 9588 -1522
rect 9528 -1532 10100 -1528
rect 9528 -1584 9532 -1532
rect 9584 -1584 10100 -1532
rect 9528 -1588 10100 -1584
rect 9528 -1594 9588 -1588
rect 10040 -1638 10100 -1588
rect 10232 -1530 10296 -1524
rect 11404 -1530 11468 -1524
rect 10232 -1536 11468 -1530
rect 10232 -1588 10238 -1536
rect 10290 -1588 11410 -1536
rect 11462 -1588 11468 -1536
rect 10232 -1594 11468 -1588
rect 10232 -1600 10296 -1594
rect 11404 -1600 11468 -1594
rect 15638 -1532 15698 -1526
rect 21746 -1532 21806 -1526
rect 15638 -1536 21806 -1532
rect 15638 -1588 15642 -1536
rect 15694 -1588 21750 -1536
rect 21802 -1588 21806 -1536
rect 15638 -1592 21806 -1588
rect 15638 -1598 15698 -1592
rect 21746 -1598 21806 -1592
rect 11566 -1638 11626 -1632
rect 17672 -1638 17732 -1632
rect 19708 -1638 19768 -1632
rect 10040 -1642 19768 -1638
rect 10040 -1694 11570 -1642
rect 11622 -1694 17676 -1642
rect 17728 -1694 19712 -1642
rect 19764 -1694 19768 -1642
rect 10040 -1698 19768 -1694
rect 11566 -1704 11626 -1698
rect 17672 -1704 17732 -1698
rect 19708 -1704 19768 -1698
rect 8510 -2570 8570 -2564
rect 10546 -2570 10606 -2564
rect 12580 -2570 12640 -2564
rect 13040 -2570 13100 -2564
rect 14618 -2568 14678 -2566
rect 14078 -2570 14150 -2568
rect 14580 -2570 14678 -2568
rect 15094 -2570 15166 -2568
rect 16122 -2570 16194 -2568
rect 8510 -2572 16500 -2570
rect 16654 -2572 16714 -2566
rect 18690 -2572 18750 -2568
rect 8510 -2574 14088 -2572
rect 8510 -2626 8514 -2574
rect 8566 -2626 10550 -2574
rect 10602 -2575 13044 -2574
rect 10602 -2578 12568 -2575
rect 10602 -2626 12044 -2578
rect 8510 -2630 12044 -2626
rect 12096 -2627 12568 -2578
rect 12620 -2626 13044 -2575
rect 13096 -2624 14088 -2574
rect 14140 -2574 15104 -2572
rect 14140 -2624 14606 -2574
rect 13096 -2626 14606 -2624
rect 14658 -2624 15104 -2574
rect 15156 -2624 16132 -2572
rect 16184 -2574 18878 -2572
rect 20724 -2574 20784 -2568
rect 16184 -2577 20784 -2574
rect 16184 -2624 16642 -2577
rect 14658 -2626 16642 -2624
rect 12620 -2627 16642 -2626
rect 12096 -2629 16642 -2627
rect 16694 -2578 20784 -2577
rect 16694 -2582 17642 -2578
rect 16694 -2629 17154 -2582
rect 12096 -2630 17154 -2629
rect 8510 -2636 8570 -2630
rect 10546 -2636 10606 -2630
rect 12034 -2634 12106 -2630
rect 12542 -2632 12640 -2630
rect 12580 -2636 12640 -2632
rect 13040 -2636 13100 -2630
rect 14618 -2632 15066 -2630
rect 15272 -2632 16086 -2630
rect 16292 -2632 17154 -2630
rect 14618 -2638 14678 -2632
rect 16616 -2634 16714 -2632
rect 16654 -2638 16714 -2634
rect 17144 -2634 17154 -2632
rect 17206 -2630 17642 -2582
rect 17694 -2582 18694 -2578
rect 17694 -2630 18154 -2582
rect 17206 -2632 18154 -2630
rect 17206 -2634 17216 -2632
rect 17632 -2634 17704 -2632
rect 18144 -2634 18154 -2632
rect 18206 -2630 18694 -2582
rect 18746 -2630 20728 -2578
rect 20780 -2630 20784 -2578
rect 18206 -2632 20784 -2630
rect 18206 -2634 18216 -2632
rect 17144 -2638 17216 -2634
rect 18144 -2638 18216 -2634
rect 18690 -2634 20784 -2632
rect 18690 -2640 18750 -2634
rect 20724 -2640 20784 -2634
rect 9526 -2680 9590 -2674
rect 19706 -2680 19770 -2674
rect 9526 -2686 23354 -2680
rect 9526 -2738 9532 -2686
rect 9584 -2738 19712 -2686
rect 19764 -2738 23354 -2686
rect 9526 -2744 23354 -2738
rect 9526 -2750 9590 -2744
rect 19706 -2750 19770 -2744
rect 7488 -2818 7552 -2812
rect 13598 -2818 13662 -2812
rect 7488 -2824 13662 -2818
rect 7488 -2876 7494 -2824
rect 7546 -2876 13604 -2824
rect 13656 -2876 13662 -2824
rect 7488 -2882 13662 -2876
rect 7488 -2888 7552 -2882
rect 13598 -2888 13662 -2882
rect 15634 -2818 15698 -2812
rect 21742 -2818 21806 -2812
rect 15634 -2824 18074 -2818
rect 15634 -2876 15640 -2824
rect 15692 -2826 18074 -2824
rect 18456 -2824 21806 -2818
rect 18456 -2826 21748 -2824
rect 15692 -2876 21748 -2826
rect 21800 -2876 21806 -2824
rect 15634 -2882 21806 -2876
rect 15634 -2888 15698 -2882
rect 6330 -2968 6390 -2962
rect 15838 -2968 15898 -2882
rect 21742 -2888 21806 -2882
rect 6330 -2972 15898 -2968
rect 6330 -3024 6334 -2972
rect 6386 -3024 7316 -2972
rect 7368 -3024 15898 -2972
rect 6330 -3028 15898 -3024
rect 6330 -3034 6390 -3028
rect 21708 -3100 21780 -3098
rect 13598 -3102 22944 -3100
rect 13592 -3108 21718 -3102
rect 9526 -3114 9590 -3108
rect 690 -3120 9590 -3114
rect 690 -3172 9532 -3120
rect 9584 -3172 9590 -3120
rect 13592 -3160 13604 -3108
rect 13656 -3154 21718 -3108
rect 21770 -3104 22944 -3102
rect 21770 -3108 22950 -3104
rect 21770 -3154 22888 -3108
rect 13656 -3160 22888 -3154
rect 22940 -3160 22950 -3108
rect 13592 -3164 22950 -3160
rect 13592 -3166 13668 -3164
rect 690 -3178 9590 -3172
rect -12032 -11183 -11932 -11172
rect -10238 -11183 -10138 -11172
rect -7638 -11183 -7538 -11172
rect -5038 -11181 -4938 -11170
rect -2438 -11181 -2338 -11170
rect -634 -11181 -534 -11170
rect -12036 -11200 -11928 -11183
rect -12036 -11256 -12010 -11200
rect -11954 -11256 -11928 -11200
rect -12036 -11273 -11928 -11256
rect -10242 -11200 -10134 -11183
rect -10242 -11256 -10216 -11200
rect -10160 -11256 -10134 -11200
rect -10242 -11273 -10134 -11256
rect -7642 -11200 -7534 -11183
rect -7642 -11256 -7616 -11200
rect -7560 -11256 -7534 -11200
rect -7642 -11273 -7534 -11256
rect -5042 -11198 -4934 -11181
rect -5042 -11254 -5016 -11198
rect -4960 -11254 -4934 -11198
rect -5042 -11271 -4934 -11254
rect -2442 -11198 -2334 -11181
rect -2442 -11254 -2416 -11198
rect -2360 -11254 -2334 -11198
rect -2442 -11271 -2334 -11254
rect -638 -11198 -530 -11181
rect -638 -11254 -612 -11198
rect -556 -11254 -530 -11198
rect -638 -11271 -530 -11254
rect -12032 -11284 -11932 -11273
rect -10238 -11284 -10138 -11273
rect -7638 -11284 -7538 -11273
rect -5038 -11282 -4938 -11271
rect -2438 -11282 -2338 -11271
rect -634 -11282 -534 -11271
rect 690 -18888 750 -3178
rect 9526 -3184 9590 -3178
rect 11564 -3304 11624 -3298
rect 952 -3308 11624 -3304
rect 952 -3360 6920 -3308
rect 6972 -3360 11568 -3308
rect 11620 -3360 11624 -3308
rect 952 -3364 11624 -3360
rect 952 -18858 1012 -3364
rect 11564 -3370 11624 -3364
rect 7312 -3404 7372 -3398
rect 8478 -3404 8538 -3398
rect 10514 -3404 10574 -3398
rect 7312 -3408 10574 -3404
rect 7312 -3460 7316 -3408
rect 7368 -3460 8482 -3408
rect 8534 -3460 10518 -3408
rect 10570 -3460 10574 -3408
rect 7312 -3464 10574 -3460
rect 7312 -3470 7372 -3464
rect 8478 -3470 8538 -3464
rect 10514 -3470 10574 -3464
rect 18660 -3404 18720 -3398
rect 20694 -3404 20754 -3398
rect 23138 -3404 23198 -3398
rect 18660 -3408 23198 -3404
rect 18660 -3460 18664 -3408
rect 18716 -3460 20698 -3408
rect 20750 -3460 23142 -3408
rect 23194 -3460 23198 -3408
rect 18660 -3464 23198 -3460
rect 18660 -3470 18720 -3464
rect 20694 -3470 20754 -3464
rect 23138 -3470 23198 -3464
rect 9496 -4352 9556 -4346
rect 11532 -4352 11592 -4346
rect 9496 -4356 11592 -4352
rect 9496 -4408 9500 -4356
rect 9552 -4408 11536 -4356
rect 11588 -4408 11592 -4356
rect 9496 -4412 11592 -4408
rect 9496 -4418 9556 -4412
rect 11532 -4418 11592 -4412
rect 19676 -4352 19736 -4346
rect 21712 -4352 21772 -4346
rect 19676 -4356 21772 -4352
rect 19676 -4408 19680 -4356
rect 19732 -4408 21716 -4356
rect 21768 -4408 21772 -4356
rect 19676 -4412 21772 -4408
rect 19676 -4418 19736 -4412
rect 7044 -4450 7104 -4444
rect 19784 -4450 19844 -4412
rect 21712 -4418 21772 -4412
rect 7044 -4454 19844 -4450
rect 4156 -4502 4216 -4496
rect 4268 -4502 4328 -4496
rect 4378 -4502 4438 -4496
rect 5028 -4502 5088 -4496
rect 5138 -4502 5198 -4496
rect 5246 -4502 5306 -4496
rect 6048 -4502 6108 -4496
rect 1330 -4506 6108 -4502
rect 1330 -4558 4160 -4506
rect 4212 -4558 4272 -4506
rect 4324 -4558 4382 -4506
rect 4434 -4558 5032 -4506
rect 5084 -4558 5142 -4506
rect 5194 -4558 5250 -4506
rect 5302 -4558 6052 -4506
rect 6104 -4558 6108 -4506
rect 7044 -4506 7048 -4454
rect 7100 -4506 19844 -4454
rect 7044 -4510 19844 -4506
rect 7044 -4516 7104 -4510
rect 1330 -4562 6108 -4558
rect 1178 -8620 1250 -8616
rect 1178 -8672 1188 -8620
rect 1240 -8672 1250 -8620
rect 1178 -8676 1250 -8672
rect 1184 -12334 1244 -8676
rect 1178 -12338 1250 -12334
rect 1178 -12390 1188 -12338
rect 1240 -12390 1250 -12338
rect 1178 -12394 1250 -12390
rect 946 -18862 1018 -18858
rect 684 -18892 756 -18888
rect 684 -18944 694 -18892
rect 746 -18944 756 -18892
rect 946 -18914 956 -18862
rect 1008 -18914 1018 -18862
rect 946 -18918 1018 -18914
rect 684 -18948 756 -18944
rect -814 -19124 -754 -19118
rect 98 -19124 158 -19118
rect 1330 -19124 1390 -4562
rect 4156 -4568 4216 -4562
rect 4268 -4568 4328 -4562
rect 4378 -4568 4438 -4562
rect 5028 -4568 5088 -4562
rect 5138 -4568 5198 -4562
rect 5246 -4568 5306 -4562
rect 6048 -4568 6108 -4562
rect 7180 -4548 7240 -4542
rect 9496 -4548 9556 -4542
rect 7180 -4552 9556 -4548
rect 7180 -4604 7184 -4552
rect 7236 -4604 9500 -4552
rect 9552 -4604 9556 -4552
rect 7180 -4608 9556 -4604
rect 7180 -4614 7240 -4608
rect 9496 -4614 9556 -4608
rect 10516 -4546 10576 -4540
rect 22978 -4546 23038 -4540
rect 10516 -4550 23038 -4546
rect 10516 -4602 10520 -4550
rect 10572 -4602 22982 -4550
rect 23034 -4602 23038 -4550
rect 10516 -4606 23038 -4602
rect 10516 -4612 10576 -4606
rect 22978 -4612 23038 -4606
rect 8482 -4658 8542 -4652
rect 10516 -4658 10576 -4652
rect 8482 -4662 10576 -4658
rect 8482 -4714 8486 -4662
rect 8538 -4714 10520 -4662
rect 10572 -4714 10576 -4662
rect 8482 -4718 10576 -4714
rect 8482 -4724 8542 -4718
rect 10516 -4724 10576 -4718
rect 13572 -4660 13632 -4654
rect 15606 -4660 15666 -4654
rect 13572 -4664 15666 -4660
rect 13572 -4716 13576 -4664
rect 13628 -4716 15610 -4664
rect 15662 -4716 15666 -4664
rect 13572 -4720 15666 -4716
rect 13572 -4726 13632 -4720
rect 15606 -4726 15666 -4720
rect 18662 -4660 18722 -4654
rect 20696 -4658 20756 -4654
rect 23290 -4658 23354 -2744
rect 20628 -4660 23354 -4658
rect 18662 -4664 23354 -4660
rect 18662 -4716 18666 -4664
rect 18718 -4716 20700 -4664
rect 20752 -4716 23354 -4664
rect 18662 -4720 23354 -4716
rect 18662 -4726 18722 -4720
rect 20628 -4722 23354 -4720
rect 20696 -4726 20756 -4722
rect 3492 -5214 3552 -5208
rect 3832 -5214 3892 -5208
rect 3942 -5214 4002 -5208
rect 4592 -5214 4652 -5208
rect 4704 -5214 4764 -5208
rect 4812 -5214 4872 -5208
rect 5464 -5214 5524 -5208
rect 5574 -5214 5634 -5208
rect 3492 -5218 5634 -5214
rect 3492 -5270 3496 -5218
rect 3548 -5270 3836 -5218
rect 3888 -5270 3946 -5218
rect 3998 -5270 4596 -5218
rect 4648 -5270 4708 -5218
rect 4760 -5270 4816 -5218
rect 4868 -5270 5468 -5218
rect 5520 -5270 5578 -5218
rect 5630 -5270 5634 -5218
rect 3492 -5274 5634 -5270
rect 3492 -5280 3552 -5274
rect 3832 -5280 3892 -5274
rect 3942 -5280 4002 -5274
rect 4592 -5280 4652 -5274
rect 4704 -5280 4764 -5274
rect 4812 -5280 4872 -5274
rect 5464 -5280 5524 -5274
rect 5574 -5280 5634 -5274
rect 4048 -5320 4108 -5314
rect 4484 -5320 4544 -5314
rect 4922 -5320 4982 -5314
rect 5356 -5320 5416 -5314
rect 4048 -5324 5416 -5320
rect 4048 -5376 4052 -5324
rect 4104 -5376 4488 -5324
rect 4540 -5376 4926 -5324
rect 4978 -5376 5360 -5324
rect 5412 -5376 5416 -5324
rect 4048 -5380 5416 -5376
rect 4048 -5386 4108 -5380
rect 4484 -5386 4544 -5380
rect 4922 -5386 4982 -5380
rect 5356 -5386 5416 -5380
rect 4268 -5436 4328 -5430
rect 5138 -5436 5198 -5430
rect 5932 -5436 5992 -5430
rect 4268 -5440 5992 -5436
rect 4268 -5492 4272 -5440
rect 4324 -5492 5142 -5440
rect 5194 -5492 5936 -5440
rect 5988 -5492 5992 -5440
rect 4268 -5496 5992 -5492
rect 4268 -5502 4328 -5496
rect 5138 -5502 5198 -5496
rect 5932 -5502 5992 -5496
rect 19526 -5594 19586 -5588
rect 19526 -5598 23948 -5594
rect 6802 -5608 6862 -5602
rect 13568 -5608 13628 -5602
rect 14588 -5608 14648 -5602
rect 16624 -5608 16684 -5602
rect 6802 -5612 16684 -5608
rect 6802 -5664 6806 -5612
rect 6858 -5664 13572 -5612
rect 13624 -5664 14592 -5612
rect 14644 -5664 16628 -5612
rect 16680 -5664 16684 -5612
rect 19526 -5650 19530 -5598
rect 19582 -5650 23948 -5598
rect 19526 -5654 23948 -5650
rect 19526 -5660 19586 -5654
rect 6802 -5668 16684 -5664
rect 6802 -5674 6862 -5668
rect 13568 -5674 13628 -5668
rect 14588 -5674 14648 -5668
rect 16624 -5674 16684 -5668
rect 19674 -5704 19734 -5698
rect 21714 -5704 21774 -5698
rect 22846 -5704 22906 -5698
rect 6916 -5712 6976 -5706
rect 11534 -5712 11594 -5706
rect 18658 -5712 18718 -5706
rect 6916 -5716 18718 -5712
rect 6916 -5768 6920 -5716
rect 6972 -5768 9502 -5716
rect 9554 -5768 11538 -5716
rect 11590 -5768 18662 -5716
rect 18714 -5768 18718 -5716
rect 6916 -5772 18718 -5768
rect 19674 -5708 22906 -5704
rect 19674 -5760 19678 -5708
rect 19730 -5760 21718 -5708
rect 21770 -5760 22850 -5708
rect 22902 -5760 22906 -5708
rect 19674 -5764 22906 -5760
rect 19674 -5770 19734 -5764
rect 21714 -5770 21774 -5764
rect 22846 -5770 22906 -5764
rect 6916 -5778 6976 -5772
rect 11534 -5778 11594 -5772
rect 18658 -5778 18718 -5772
rect 11532 -5814 11592 -5808
rect 20694 -5814 20754 -5808
rect 11532 -5818 20754 -5814
rect 11532 -5870 11536 -5818
rect 11588 -5870 20698 -5818
rect 20750 -5870 20754 -5818
rect 11532 -5874 20754 -5870
rect 11532 -5880 11592 -5874
rect 20694 -5880 20754 -5874
rect 9498 -5916 9558 -5910
rect 11532 -5916 11592 -5910
rect 9498 -5920 11592 -5916
rect 9498 -5972 9502 -5920
rect 9554 -5972 11536 -5920
rect 11588 -5972 11592 -5920
rect 9498 -5976 11592 -5972
rect 9498 -5982 9558 -5976
rect 11532 -5982 11592 -5976
rect 14588 -5914 14648 -5908
rect 15606 -5914 15666 -5908
rect 16622 -5914 16682 -5908
rect 19526 -5914 19586 -5908
rect 14588 -5918 19586 -5914
rect 14588 -5970 14592 -5918
rect 14644 -5970 15610 -5918
rect 15662 -5970 16626 -5918
rect 16678 -5970 19530 -5918
rect 19582 -5970 19586 -5918
rect 14588 -5974 19586 -5970
rect 14588 -5980 14648 -5974
rect 15606 -5980 15666 -5974
rect 16622 -5980 16682 -5974
rect 19526 -5980 19586 -5974
rect 19678 -5912 19738 -5906
rect 21712 -5912 21772 -5906
rect 22978 -5912 23038 -5906
rect 19678 -5916 23820 -5912
rect 19678 -5968 19682 -5916
rect 19734 -5968 21716 -5916
rect 21768 -5968 22982 -5916
rect 23034 -5968 23820 -5916
rect 19678 -5972 23820 -5968
rect 19678 -5978 19738 -5972
rect 21712 -5978 21772 -5972
rect 22978 -5978 23038 -5972
rect 2110 -6160 2170 -6154
rect 3832 -6160 3892 -6154
rect 4266 -6160 4326 -6154
rect 4702 -6160 4762 -6154
rect 5138 -6160 5198 -6154
rect 5576 -6160 5636 -6154
rect 2110 -6164 5636 -6160
rect 2110 -6216 2114 -6164
rect 2166 -6216 3836 -6164
rect 3888 -6216 4270 -6164
rect 4322 -6216 4706 -6164
rect 4758 -6216 5142 -6164
rect 5194 -6216 5580 -6164
rect 5632 -6216 5636 -6164
rect 2110 -6220 5636 -6216
rect 2110 -6226 2170 -6220
rect 3832 -6226 3892 -6220
rect 4266 -6226 4326 -6220
rect 4702 -6226 4762 -6220
rect 5138 -6226 5198 -6220
rect 5576 -6226 5636 -6220
rect 4048 -6264 4108 -6258
rect 4484 -6264 4544 -6258
rect 4922 -6264 4982 -6258
rect 5356 -6264 5416 -6258
rect 4048 -6268 5416 -6264
rect 4048 -6320 4052 -6268
rect 4104 -6320 4488 -6268
rect 4540 -6320 4926 -6268
rect 4978 -6320 5360 -6268
rect 5412 -6320 5416 -6268
rect 4048 -6324 5416 -6320
rect 4048 -6330 4108 -6324
rect 4484 -6330 4544 -6324
rect 4922 -6330 4982 -6324
rect 5356 -6330 5416 -6324
rect 3942 -6362 4002 -6356
rect 4156 -6362 4216 -6356
rect 4376 -6362 4436 -6356
rect 4594 -6362 4654 -6356
rect 4704 -6362 4764 -6356
rect 4810 -6362 4870 -6356
rect 5028 -6362 5088 -6356
rect 5246 -6362 5306 -6356
rect 5462 -6362 5522 -6356
rect 3942 -6366 5522 -6362
rect 3942 -6418 3946 -6366
rect 3998 -6418 4160 -6366
rect 4212 -6418 4380 -6366
rect 4432 -6418 4598 -6366
rect 4650 -6418 4708 -6366
rect 4760 -6418 4814 -6366
rect 4866 -6418 5032 -6366
rect 5084 -6418 5250 -6366
rect 5302 -6418 5466 -6366
rect 5518 -6418 5522 -6366
rect 3942 -6422 5522 -6418
rect 3942 -6428 4002 -6422
rect 4156 -6428 4216 -6422
rect 4376 -6428 4436 -6422
rect 4594 -6428 4654 -6422
rect 4704 -6428 4764 -6422
rect 4810 -6428 4870 -6422
rect 5028 -6428 5088 -6422
rect 5246 -6428 5306 -6422
rect 5462 -6428 5522 -6422
rect 8480 -6864 8540 -6858
rect 10516 -6864 10576 -6858
rect 6914 -6868 10576 -6864
rect 6914 -6920 8484 -6868
rect 8536 -6920 10520 -6868
rect 10572 -6920 10576 -6868
rect 6914 -6924 10576 -6920
rect -814 -19128 1390 -19124
rect -814 -19180 -810 -19128
rect -758 -19180 102 -19128
rect 154 -19180 1390 -19128
rect -814 -19184 1390 -19180
rect 1468 -7002 3558 -6998
rect 1468 -7054 3496 -7002
rect 3548 -7054 3558 -7002
rect 1468 -7058 3558 -7054
rect -814 -19190 -754 -19184
rect 98 -19190 158 -19184
rect -1684 -19234 -1624 -19228
rect -22 -19234 38 -19228
rect -1684 -19238 38 -19234
rect -1684 -19290 -1680 -19238
rect -1628 -19290 -18 -19238
rect 34 -19290 38 -19238
rect -1684 -19294 38 -19290
rect -1684 -19300 -1624 -19294
rect -22 -19300 38 -19294
rect -2598 -19342 -2538 -19336
rect -920 -19342 -860 -19336
rect -702 -19342 -642 -19336
rect -2598 -19346 -642 -19342
rect -2598 -19398 -2594 -19346
rect -2542 -19398 -916 -19346
rect -864 -19398 -698 -19346
rect -646 -19398 -642 -19346
rect -2598 -19402 -642 -19398
rect -2598 -19408 -2538 -19402
rect -920 -19408 -860 -19402
rect -702 -19408 -642 -19402
rect -2468 -19450 -2408 -19444
rect -1138 -19450 -1078 -19444
rect -484 -19450 -424 -19444
rect -2468 -19454 -424 -19450
rect -2468 -19506 -2464 -19454
rect -2412 -19506 -1134 -19454
rect -1082 -19506 -480 -19454
rect -428 -19506 -424 -19454
rect -2468 -19510 -424 -19506
rect -2468 -19516 -2408 -19510
rect -1138 -19516 -1078 -19510
rect -484 -19516 -424 -19510
rect 1468 -19724 1528 -7058
rect 3832 -7098 3892 -7092
rect 4702 -7098 4762 -7092
rect 5576 -7098 5636 -7092
rect 5932 -7098 5992 -7092
rect -28 -19728 1528 -19724
rect -28 -19780 -18 -19728
rect 34 -19780 1528 -19728
rect -28 -19784 1528 -19780
rect 1586 -7102 5992 -7098
rect 1586 -7154 3836 -7102
rect 3888 -7154 4706 -7102
rect 4758 -7154 5580 -7102
rect 5632 -7154 5936 -7102
rect 5988 -7154 5992 -7102
rect 1586 -7158 5992 -7154
rect -2010 -19950 -1950 -19944
rect -1354 -19950 -1294 -19944
rect -484 -19950 -424 -19944
rect 220 -19950 280 -19944
rect -2010 -19954 280 -19950
rect -2010 -20006 -2006 -19954
rect -1954 -20006 -1350 -19954
rect -1298 -20006 -480 -19954
rect -428 -20006 224 -19954
rect 276 -20006 280 -19954
rect -2010 -20010 280 -20006
rect -2010 -20016 -1950 -20010
rect -1354 -20016 -1294 -20010
rect -484 -20016 -424 -20010
rect 220 -20016 280 -20010
rect -1902 -20050 -1842 -20044
rect -1464 -20050 -1404 -20044
rect -3096 -20054 -968 -20050
rect -3096 -20106 -1898 -20054
rect -1846 -20106 -1460 -20054
rect -1408 -20106 -968 -20054
rect -3096 -20110 -968 -20106
rect -7386 -21600 -7326 -21594
rect -5346 -21600 -5286 -21594
rect -7386 -21604 -5286 -21600
rect -7386 -21656 -7382 -21604
rect -7330 -21656 -5342 -21604
rect -5290 -21656 -5286 -21604
rect -7386 -21660 -5286 -21656
rect -7386 -21666 -7326 -21660
rect -5346 -21666 -5286 -21660
rect -9538 -22504 -9478 -22498
rect -8400 -22504 -8340 -22498
rect -4326 -22504 -4266 -22498
rect -9538 -22508 -4266 -22504
rect -9538 -22560 -9534 -22508
rect -9482 -22560 -8396 -22508
rect -8344 -22560 -4322 -22508
rect -4270 -22560 -4266 -22508
rect -9538 -22564 -4266 -22560
rect -9538 -22570 -9478 -22564
rect -8400 -22570 -8340 -22564
rect -4326 -22570 -4266 -22564
rect -7386 -22600 -7326 -22594
rect -5346 -22600 -5286 -22594
rect -7386 -22604 -5286 -22600
rect -7386 -22656 -7382 -22604
rect -7330 -22656 -5342 -22604
rect -5290 -22656 -5286 -22604
rect -7386 -22660 -5286 -22656
rect -7386 -22666 -7326 -22660
rect -5346 -22666 -5286 -22660
rect -6364 -22716 -6304 -22710
rect -3202 -22716 -3142 -22710
rect -6364 -22720 -3142 -22716
rect -6364 -22772 -6360 -22720
rect -6308 -22772 -3198 -22720
rect -3146 -22772 -3142 -22720
rect -6364 -22776 -3142 -22772
rect -6364 -22782 -6304 -22776
rect -3202 -22782 -3142 -22776
rect -8254 -23616 -8194 -23610
rect -6368 -23616 -6308 -23610
rect -4498 -23616 -4438 -23610
rect -3096 -23616 -3036 -20110
rect -1902 -20116 -1842 -20110
rect -1464 -20116 -1404 -20110
rect -2976 -20160 -2916 -20154
rect -1900 -20160 -1840 -20154
rect -1466 -20160 -1406 -20154
rect -1138 -20160 -1078 -20154
rect -2976 -20164 -1078 -20160
rect -2976 -20216 -2972 -20164
rect -2920 -20216 -1896 -20164
rect -1844 -20216 -1462 -20164
rect -1410 -20216 -1134 -20164
rect -1082 -20216 -1078 -20164
rect -2976 -20220 -1078 -20216
rect -2976 -20226 -2916 -20220
rect -1900 -20226 -1840 -20220
rect -1466 -20226 -1406 -20220
rect -1138 -20226 -1078 -20220
rect -1028 -20160 -968 -20110
rect -374 -20070 -314 -20064
rect 1586 -20070 1646 -7158
rect 3832 -7164 3892 -7158
rect 4702 -7164 4762 -7158
rect 5576 -7164 5636 -7158
rect 5932 -7164 5992 -7158
rect 4048 -7196 4108 -7190
rect 4484 -7196 4544 -7190
rect 4922 -7196 4982 -7190
rect 5356 -7196 5416 -7190
rect 4048 -7200 5416 -7196
rect 4048 -7252 4052 -7200
rect 4104 -7252 4488 -7200
rect 4540 -7252 4926 -7200
rect 4978 -7252 5360 -7200
rect 5412 -7252 5416 -7200
rect 4048 -7256 5416 -7252
rect 4048 -7262 4108 -7256
rect 4484 -7262 4544 -7256
rect 4922 -7262 4982 -7256
rect 5356 -7262 5416 -7256
rect 3492 -7314 3552 -7308
rect 4158 -7314 4218 -7308
rect 4266 -7314 4326 -7308
rect 4374 -7314 4434 -7308
rect 5020 -7314 5080 -7308
rect 5138 -7314 5198 -7308
rect 3492 -7316 5198 -7314
rect 5247 -7316 5305 -7310
rect 3492 -7318 5305 -7316
rect 3492 -7370 3496 -7318
rect 3548 -7370 4162 -7318
rect 4214 -7370 4270 -7318
rect 4322 -7370 4378 -7318
rect 4430 -7370 5024 -7318
rect 5076 -7370 5142 -7318
rect 5194 -7319 5305 -7318
rect 5194 -7370 5250 -7319
rect 3492 -7371 5250 -7370
rect 5302 -7371 5305 -7319
rect 3492 -7374 5305 -7371
rect 3492 -7380 3552 -7374
rect 4158 -7380 4218 -7374
rect 4266 -7380 4326 -7374
rect 4374 -7380 4434 -7374
rect 5020 -7380 5080 -7374
rect 5138 -7380 5198 -7374
rect 5247 -7380 5305 -7374
rect 2318 -7644 2426 -7627
rect 2318 -7700 2344 -7644
rect 2400 -7700 2426 -7644
rect 2318 -7717 2426 -7700
rect 2110 -8396 2170 -8386
rect 2110 -8448 2114 -8396
rect 2166 -8448 2170 -8396
rect 1948 -8502 2020 -8498
rect 1948 -8554 1958 -8502
rect 2010 -8554 2020 -8502
rect 1948 -8558 2020 -8554
rect 1696 -10140 1804 -10123
rect 1696 -10196 1722 -10140
rect 1778 -10196 1804 -10140
rect 1696 -10213 1804 -10196
rect 1720 -11476 1780 -10213
rect 1954 -11352 2014 -8558
rect 1954 -11404 1958 -11352
rect 2010 -11404 2014 -11352
rect 1954 -11414 2014 -11404
rect 2110 -11352 2170 -8448
rect 2110 -11404 2114 -11352
rect 2166 -11404 2170 -11352
rect 2336 -11356 2396 -7717
rect 3832 -8034 3892 -8028
rect 3942 -8034 4002 -8028
rect 4596 -8034 4656 -8028
rect 4702 -8034 4762 -8028
rect 4812 -8034 4872 -8028
rect 5464 -8034 5524 -8028
rect 5576 -8034 5636 -8028
rect 6048 -8034 6108 -8028
rect 3832 -8038 6108 -8034
rect 3832 -8090 3836 -8038
rect 3888 -8090 3946 -8038
rect 3998 -8090 4600 -8038
rect 4652 -8090 4706 -8038
rect 4758 -8090 4816 -8038
rect 4868 -8090 5468 -8038
rect 5520 -8090 5580 -8038
rect 5632 -8090 6052 -8038
rect 6104 -8090 6108 -8038
rect 3832 -8094 6108 -8090
rect 3832 -8100 3892 -8094
rect 3942 -8100 4002 -8094
rect 4596 -8100 4656 -8094
rect 4702 -8100 4762 -8094
rect 4812 -8100 4872 -8094
rect 5464 -8100 5524 -8094
rect 5576 -8100 5636 -8094
rect 6048 -8100 6108 -8094
rect 2110 -11414 2170 -11404
rect 2330 -11360 2402 -11356
rect 2330 -11412 2340 -11360
rect 2392 -11412 2402 -11360
rect 2330 -11416 2402 -11412
rect 6914 -11476 6974 -6924
rect 8480 -6930 8540 -6924
rect 10516 -6930 10576 -6924
rect 13570 -6862 13630 -6856
rect 15606 -6862 15666 -6856
rect 13570 -6866 15666 -6862
rect 13570 -6918 13574 -6866
rect 13626 -6918 15610 -6866
rect 15662 -6918 15666 -6866
rect 13570 -6922 15666 -6918
rect 13570 -6928 13630 -6922
rect 15606 -6928 15666 -6922
rect 18660 -6860 18720 -6854
rect 20696 -6860 20756 -6854
rect 18660 -6864 20756 -6860
rect 18660 -6916 18664 -6864
rect 18716 -6916 20700 -6864
rect 20752 -6916 20756 -6864
rect 18660 -6920 20756 -6916
rect 18660 -6926 18720 -6920
rect 20696 -6926 20756 -6920
rect 10516 -6972 10576 -6966
rect 22846 -6972 22906 -6966
rect 10516 -6976 22906 -6972
rect 10516 -7028 10520 -6976
rect 10572 -7028 22850 -6976
rect 22902 -7028 22906 -6976
rect 10516 -7032 22906 -7028
rect 10516 -7038 10576 -7032
rect 22846 -7038 22906 -7032
rect 7312 -7072 7372 -7066
rect 7312 -7076 19896 -7072
rect 7312 -7128 7316 -7076
rect 7368 -7128 19896 -7076
rect 7312 -7132 19896 -7128
rect 7312 -7138 7372 -7132
rect 11732 -7168 11792 -7162
rect 9494 -7174 9554 -7168
rect 11528 -7174 11588 -7168
rect 9494 -7178 11588 -7174
rect 9494 -7230 9498 -7178
rect 9550 -7230 11532 -7178
rect 11584 -7230 11588 -7178
rect 9494 -7234 11588 -7230
rect 11732 -7172 13632 -7168
rect 11732 -7224 11736 -7172
rect 11788 -7224 13570 -7172
rect 13622 -7224 13632 -7172
rect 11732 -7228 13632 -7224
rect 14586 -7172 14646 -7166
rect 16620 -7172 16680 -7166
rect 14586 -7176 16680 -7172
rect 14586 -7228 14590 -7176
rect 14642 -7228 16624 -7176
rect 16676 -7228 16680 -7176
rect 11732 -7234 11792 -7228
rect 14586 -7232 16680 -7228
rect 9494 -7240 9554 -7234
rect 11528 -7240 11588 -7234
rect 14586 -7238 14646 -7232
rect 16620 -7238 16680 -7232
rect 16834 -7176 16894 -7170
rect 19682 -7174 19742 -7168
rect 19836 -7174 19896 -7132
rect 21716 -7174 21776 -7168
rect 16834 -7180 19236 -7176
rect 16834 -7232 16838 -7180
rect 16890 -7232 19174 -7180
rect 19226 -7232 19236 -7180
rect 16834 -7236 19236 -7232
rect 19682 -7178 21776 -7174
rect 19682 -7230 19686 -7178
rect 19738 -7230 21720 -7178
rect 21772 -7230 21776 -7178
rect 19682 -7234 21776 -7230
rect 16834 -7242 16894 -7236
rect 19682 -7240 19742 -7234
rect 21716 -7240 21776 -7234
rect 7044 -8122 7104 -8116
rect 8476 -8122 8536 -8116
rect 10512 -8122 10572 -8116
rect 7044 -8126 10572 -8122
rect 7044 -8178 7048 -8126
rect 7100 -8178 8480 -8126
rect 8532 -8178 10516 -8126
rect 10568 -8178 10572 -8126
rect 7044 -8182 10572 -8178
rect 7044 -8188 7104 -8182
rect 8476 -8188 8536 -8182
rect 10512 -8188 10572 -8182
rect 18664 -8122 18724 -8116
rect 20700 -8122 20760 -8116
rect 18664 -8126 20760 -8122
rect 18664 -8178 18668 -8126
rect 18720 -8178 20704 -8126
rect 20756 -8178 20760 -8126
rect 18664 -8182 20760 -8178
rect 18664 -8188 18724 -8182
rect 7180 -8252 7240 -8246
rect 18794 -8252 18854 -8182
rect 20700 -8188 20760 -8182
rect 7180 -8256 18854 -8252
rect 7180 -8308 7184 -8256
rect 7236 -8308 18854 -8256
rect 7180 -8312 18854 -8308
rect 7180 -8318 7240 -8312
rect 11534 -8392 11594 -8386
rect 23138 -8392 23198 -8386
rect 11534 -8396 23198 -8392
rect 11534 -8448 11538 -8396
rect 11590 -8448 23142 -8396
rect 23194 -8448 23198 -8396
rect 11534 -8452 23198 -8448
rect 11534 -8458 11594 -8452
rect 1720 -11536 6974 -11476
rect 1720 -16460 1780 -11536
rect 1850 -12448 1910 -12442
rect 2568 -12448 2628 -12442
rect 4604 -12448 4664 -12442
rect 6638 -12448 6698 -12442
rect 8678 -12448 8738 -12442
rect 10714 -12448 10774 -12442
rect 12748 -12448 12808 -12442
rect 14784 -12448 14844 -12442
rect 16820 -12448 16880 -12442
rect 18856 -12448 18916 -12442
rect 20894 -12448 20954 -12442
rect 22924 -12448 22984 -12442
rect 1850 -12452 22984 -12448
rect 1850 -12504 1854 -12452
rect 1906 -12504 2572 -12452
rect 2624 -12504 4608 -12452
rect 4660 -12504 6642 -12452
rect 6694 -12504 8682 -12452
rect 8734 -12504 10718 -12452
rect 10770 -12504 12752 -12452
rect 12804 -12504 14788 -12452
rect 14840 -12504 16824 -12452
rect 16876 -12504 18860 -12452
rect 18912 -12504 20898 -12452
rect 20950 -12504 22928 -12452
rect 22980 -12504 22984 -12452
rect 1850 -12508 22984 -12504
rect 1850 -12514 1910 -12508
rect 2568 -12514 2628 -12508
rect 4604 -12514 4664 -12508
rect 6638 -12514 6698 -12508
rect 8678 -12514 8738 -12508
rect 10714 -12514 10774 -12508
rect 12748 -12514 12808 -12508
rect 14784 -12514 14844 -12508
rect 16820 -12514 16880 -12508
rect 18856 -12514 18916 -12508
rect 20894 -12514 20954 -12508
rect 22924 -12514 22984 -12508
rect 3586 -12546 3646 -12540
rect 5624 -12546 5684 -12540
rect 7658 -12546 7718 -12540
rect 9692 -12546 9752 -12540
rect 11732 -12546 11792 -12540
rect 13766 -12546 13826 -12540
rect 15804 -12546 15864 -12540
rect 17836 -12546 17896 -12540
rect 19874 -12546 19934 -12540
rect 21912 -12546 21972 -12540
rect 23046 -12546 23106 -8452
rect 23138 -8458 23198 -8452
rect 23648 -12546 23708 -12540
rect 3586 -12550 23708 -12546
rect 3586 -12602 3590 -12550
rect 3642 -12602 5628 -12550
rect 5680 -12602 7662 -12550
rect 7714 -12602 9696 -12550
rect 9748 -12602 11736 -12550
rect 11788 -12602 13770 -12550
rect 13822 -12602 15808 -12550
rect 15860 -12602 17840 -12550
rect 17892 -12602 19878 -12550
rect 19930 -12602 21916 -12550
rect 21968 -12602 23652 -12550
rect 23704 -12602 23708 -12550
rect 3586 -12606 23708 -12602
rect 3586 -12612 3646 -12606
rect 5624 -12612 5684 -12606
rect 7658 -12612 7718 -12606
rect 9692 -12612 9752 -12606
rect 11732 -12612 11792 -12606
rect 13766 -12612 13826 -12606
rect 15804 -12612 15864 -12606
rect 17836 -12612 17896 -12606
rect 19874 -12612 19934 -12606
rect 21912 -12612 21972 -12606
rect 23648 -12612 23708 -12606
rect 11732 -12758 11792 -12752
rect 13764 -12758 13824 -12752
rect 11732 -12762 13824 -12758
rect 11732 -12814 11736 -12762
rect 11788 -12814 13768 -12762
rect 13820 -12814 13824 -12762
rect 11732 -12818 13824 -12814
rect 11732 -12824 11792 -12818
rect 13764 -12824 13824 -12818
rect 6272 -13678 6332 -13672
rect 6642 -13678 6702 -13672
rect 7144 -13678 7204 -13672
rect 7656 -13678 7716 -13672
rect 8184 -13678 8244 -13672
rect 8676 -13678 8736 -13672
rect 10708 -13678 10768 -13672
rect 12744 -13678 12804 -13672
rect 14780 -13678 14840 -13672
rect 16818 -13678 16878 -13672
rect 18856 -13678 18916 -13672
rect 19364 -13678 19424 -13672
rect 6272 -13682 19424 -13678
rect 6272 -13734 6276 -13682
rect 6328 -13734 6646 -13682
rect 6698 -13734 7148 -13682
rect 7200 -13734 7660 -13682
rect 7712 -13734 8188 -13682
rect 8240 -13734 8680 -13682
rect 8732 -13734 10712 -13682
rect 10764 -13734 12748 -13682
rect 12800 -13734 14784 -13682
rect 14836 -13734 16822 -13682
rect 16874 -13734 18346 -13682
rect 18398 -13734 18860 -13682
rect 18912 -13734 19368 -13682
rect 19420 -13734 19424 -13682
rect 6272 -13738 19424 -13734
rect 6272 -13744 6332 -13738
rect 6642 -13744 6702 -13738
rect 7144 -13744 7204 -13738
rect 7656 -13744 7716 -13738
rect 8184 -13744 8244 -13738
rect 8676 -13744 8736 -13738
rect 10708 -13744 10768 -13738
rect 12744 -13744 12804 -13738
rect 14780 -13744 14840 -13738
rect 16818 -13744 16878 -13738
rect 18856 -13744 18916 -13738
rect 19364 -13744 19424 -13738
rect 4096 -13788 4156 -13782
rect 5118 -13788 5178 -13782
rect 9190 -13788 9250 -13782
rect 9694 -13788 9754 -13782
rect 10210 -13788 10270 -13782
rect 11230 -13788 11290 -13782
rect 11732 -13788 11792 -13782
rect 12232 -13788 12292 -13782
rect 13258 -13788 13318 -13782
rect 13768 -13788 13828 -13782
rect 14276 -13788 14336 -13782
rect 15284 -13788 15344 -13782
rect 15806 -13788 15866 -13782
rect 16296 -13788 16356 -13782
rect 17328 -13788 17388 -13782
rect 17840 -13788 17900 -13782
rect 20384 -13788 20444 -13782
rect 21404 -13788 21464 -13782
rect 2106 -13792 21464 -13788
rect 2106 -13844 2116 -13792
rect 2168 -13844 4100 -13792
rect 4152 -13844 5122 -13792
rect 5174 -13844 9194 -13792
rect 9246 -13844 9698 -13792
rect 9750 -13844 10214 -13792
rect 10266 -13844 11234 -13792
rect 11286 -13844 11736 -13792
rect 11788 -13844 12236 -13792
rect 12288 -13844 13262 -13792
rect 13314 -13844 13772 -13792
rect 13824 -13844 14280 -13792
rect 14332 -13844 15288 -13792
rect 15340 -13844 15810 -13792
rect 15862 -13844 16300 -13792
rect 16352 -13844 17332 -13792
rect 17384 -13844 17844 -13792
rect 17896 -13844 20388 -13792
rect 20440 -13844 21408 -13792
rect 21460 -13844 21464 -13792
rect 2106 -13848 21464 -13844
rect 4096 -13854 4156 -13848
rect 5118 -13854 5178 -13848
rect 9190 -13854 9250 -13848
rect 9694 -13854 9754 -13848
rect 10210 -13854 10270 -13848
rect 11230 -13854 11290 -13848
rect 11732 -13854 11792 -13848
rect 12232 -13854 12292 -13848
rect 13258 -13854 13318 -13848
rect 13768 -13854 13828 -13848
rect 14276 -13854 14336 -13848
rect 15284 -13854 15344 -13848
rect 15806 -13854 15866 -13848
rect 16296 -13854 16356 -13848
rect 17328 -13854 17388 -13848
rect 17840 -13854 17900 -13848
rect 20384 -13854 20444 -13848
rect 21404 -13854 21464 -13848
rect 7138 -13892 7198 -13886
rect 8158 -13892 8218 -13886
rect 12372 -13892 12432 -13886
rect 13380 -13892 13440 -13886
rect 14422 -13892 14482 -13886
rect 17314 -13892 17374 -13886
rect 18352 -13892 18412 -13886
rect 19352 -13892 19412 -13886
rect 6132 -13896 19412 -13892
rect 6132 -13948 6142 -13896
rect 6194 -13948 7142 -13896
rect 7194 -13948 8162 -13896
rect 8214 -13948 12376 -13896
rect 12428 -13948 13384 -13896
rect 13436 -13948 14426 -13896
rect 14478 -13948 17318 -13896
rect 17370 -13948 18356 -13896
rect 18408 -13948 19356 -13896
rect 19408 -13948 19412 -13896
rect 6132 -13952 19412 -13948
rect 7138 -13958 7198 -13952
rect 8158 -13958 8218 -13952
rect 12372 -13958 12432 -13952
rect 13380 -13958 13440 -13952
rect 14422 -13958 14482 -13952
rect 17314 -13958 17374 -13952
rect 18352 -13958 18412 -13952
rect 19352 -13958 19412 -13952
rect 1976 -14000 2036 -13994
rect 2572 -14000 2632 -13994
rect 3070 -14000 3130 -13994
rect 3582 -14000 3642 -13994
rect 5624 -14000 5684 -13994
rect 7658 -14000 7718 -13994
rect 9692 -14000 9752 -13994
rect 15806 -14000 15866 -13994
rect 17838 -14000 17898 -13994
rect 19870 -14000 19930 -13994
rect 21912 -14000 21972 -13994
rect 22416 -14000 22476 -13994
rect 22926 -14000 22986 -13994
rect 1976 -14004 22986 -14000
rect 1976 -14056 1980 -14004
rect 2032 -14056 2576 -14004
rect 2628 -14056 3074 -14004
rect 3126 -14056 3586 -14004
rect 3638 -14056 5628 -14004
rect 5680 -14056 7662 -14004
rect 7714 -14056 9696 -14004
rect 9748 -14056 11852 -14004
rect 11904 -14006 15810 -14004
rect 11904 -14056 13576 -14006
rect 1976 -14058 13576 -14056
rect 13628 -14056 15810 -14006
rect 15862 -14056 17842 -14004
rect 17894 -14056 19874 -14004
rect 19926 -14056 21916 -14004
rect 21968 -14056 22420 -14004
rect 22472 -14056 22930 -14004
rect 22982 -14056 22986 -14004
rect 13628 -14058 22986 -14056
rect 1976 -14060 22986 -14058
rect 1976 -14066 2036 -14060
rect 2572 -14066 2632 -14060
rect 3070 -14066 3130 -14060
rect 3582 -14066 3642 -14060
rect 5624 -14066 5684 -14060
rect 7658 -14066 7718 -14060
rect 9692 -14066 9752 -14060
rect 13566 -14062 13638 -14060
rect 15806 -14066 15866 -14060
rect 17838 -14066 17898 -14060
rect 19870 -14066 19930 -14060
rect 21912 -14066 21972 -14060
rect 22416 -14066 22476 -14060
rect 22926 -14066 22986 -14060
rect 5102 -14890 5162 -14884
rect 6122 -14890 6182 -14884
rect 7134 -14890 7194 -14884
rect 8160 -14890 8220 -14884
rect 17316 -14890 17376 -14884
rect 18352 -14890 18412 -14884
rect 19368 -14890 19428 -14884
rect 5102 -14894 19428 -14890
rect 1850 -14902 1910 -14896
rect 4086 -14902 4146 -14896
rect 1850 -14906 4146 -14902
rect 1850 -14958 1854 -14906
rect 1906 -14958 4090 -14906
rect 4142 -14958 4146 -14906
rect 5102 -14946 5106 -14894
rect 5158 -14946 6126 -14894
rect 6178 -14946 7138 -14894
rect 7190 -14946 8164 -14894
rect 8216 -14946 17320 -14894
rect 17372 -14946 18356 -14894
rect 18408 -14946 19372 -14894
rect 19424 -14946 19428 -14894
rect 5102 -14950 19428 -14946
rect 5102 -14956 5162 -14950
rect 6122 -14956 6182 -14950
rect 7134 -14956 7194 -14950
rect 8160 -14956 8220 -14950
rect 17316 -14956 17376 -14950
rect 18352 -14956 18412 -14950
rect 19368 -14956 19428 -14950
rect 1850 -14962 4146 -14958
rect 1850 -14968 1910 -14962
rect 4086 -14968 4146 -14962
rect 4598 -14994 4658 -14988
rect 5622 -14994 5682 -14988
rect 6634 -14994 6694 -14988
rect 7654 -14994 7714 -14988
rect 8676 -14994 8736 -14988
rect 10712 -14994 10772 -14988
rect 12750 -14994 12810 -14988
rect 14780 -14994 14840 -14988
rect 15800 -14994 15860 -14988
rect 16818 -14994 16878 -14988
rect 17838 -14994 17898 -14988
rect 18854 -14994 18914 -14988
rect 20890 -14994 20950 -14988
rect 4598 -14998 20950 -14994
rect 4598 -15050 4602 -14998
rect 4654 -15050 5626 -14998
rect 5678 -15050 6638 -14998
rect 6690 -15050 7658 -14998
rect 7710 -15050 8680 -14998
rect 8732 -15050 10716 -14998
rect 10768 -15050 12754 -14998
rect 12806 -15050 14784 -14998
rect 14836 -15050 15804 -14998
rect 15856 -15050 16822 -14998
rect 16874 -15050 17842 -14998
rect 17894 -15050 18858 -14998
rect 18910 -15050 20894 -14998
rect 20946 -15050 20950 -14998
rect 4598 -15054 20950 -15050
rect 4598 -15060 4658 -15054
rect 5622 -15060 5682 -15054
rect 6634 -15060 6694 -15054
rect 7654 -15060 7714 -15054
rect 8676 -15060 8736 -15054
rect 10712 -15060 10772 -15054
rect 12750 -15060 12810 -15054
rect 14780 -15060 14840 -15054
rect 15800 -15060 15860 -15054
rect 16818 -15060 16878 -15054
rect 17838 -15060 17898 -15054
rect 18854 -15060 18914 -15054
rect 20890 -15060 20950 -15054
rect 2336 -15116 2396 -15110
rect 9696 -15116 9756 -15110
rect 11730 -15116 11790 -15110
rect 13760 -15116 13820 -15110
rect 23760 -15116 23820 -5972
rect 2336 -15120 23820 -15116
rect 2336 -15172 2340 -15120
rect 2392 -15172 9700 -15120
rect 9752 -15172 11734 -15120
rect 11786 -15172 13764 -15120
rect 13816 -15172 23820 -15120
rect 2336 -15176 23820 -15172
rect 2336 -15182 2396 -15176
rect 9696 -15182 9756 -15176
rect 11730 -15182 11790 -15176
rect 13760 -15182 13820 -15176
rect 4604 -15228 4664 -15222
rect 6640 -15228 6700 -15222
rect 23034 -15228 23094 -15222
rect 4604 -15232 23094 -15228
rect 4604 -15284 4608 -15232
rect 4660 -15284 6644 -15232
rect 6696 -15284 23038 -15232
rect 23090 -15284 23094 -15232
rect 4604 -15288 23094 -15284
rect 4604 -15294 4664 -15288
rect 6640 -15294 6700 -15288
rect 23034 -15294 23094 -15288
rect 22928 -16116 22988 -16110
rect 23888 -16116 23948 -5654
rect 22928 -16120 23948 -16116
rect 5620 -16134 5680 -16128
rect 7656 -16134 7716 -16128
rect 15800 -16134 15860 -16128
rect 17836 -16134 17896 -16128
rect 21910 -16134 21970 -16128
rect 5620 -16138 21970 -16134
rect 2448 -16158 2508 -16152
rect 3586 -16158 3646 -16152
rect 2448 -16162 4468 -16158
rect 2448 -16214 2452 -16162
rect 2504 -16214 3590 -16162
rect 3642 -16214 4468 -16162
rect 5620 -16190 5624 -16138
rect 5676 -16190 7660 -16138
rect 7712 -16190 15804 -16138
rect 15856 -16190 17840 -16138
rect 17892 -16190 21914 -16138
rect 21966 -16190 21970 -16138
rect 22928 -16172 22932 -16120
rect 22984 -16172 23948 -16120
rect 22928 -16176 23948 -16172
rect 22928 -16182 22988 -16176
rect 5620 -16194 21970 -16190
rect 5620 -16200 5680 -16194
rect 7656 -16200 7716 -16194
rect 15800 -16200 15860 -16194
rect 17836 -16200 17896 -16194
rect 21910 -16200 21970 -16194
rect 2448 -16218 4468 -16214
rect 2448 -16224 2508 -16218
rect 3586 -16224 3646 -16218
rect 2336 -16358 2396 -16352
rect 3584 -16358 3644 -16352
rect 2336 -16362 3644 -16358
rect 2336 -16414 2340 -16362
rect 2392 -16414 3588 -16362
rect 3640 -16414 3644 -16362
rect 4408 -16354 4468 -16218
rect 4602 -16238 4662 -16232
rect 6642 -16238 6702 -16232
rect 8674 -16238 8734 -16232
rect 10708 -16238 10768 -16232
rect 12748 -16238 12808 -16232
rect 14782 -16238 14842 -16232
rect 4602 -16242 14842 -16238
rect 4602 -16294 4606 -16242
rect 4658 -16294 6646 -16242
rect 6698 -16294 8678 -16242
rect 8730 -16294 10712 -16242
rect 10764 -16294 12752 -16242
rect 12804 -16294 14786 -16242
rect 14838 -16294 14842 -16242
rect 4602 -16298 14842 -16294
rect 4602 -16304 4662 -16298
rect 6642 -16304 6702 -16298
rect 8674 -16304 8734 -16298
rect 10708 -16304 10768 -16298
rect 12748 -16304 12808 -16298
rect 14782 -16304 14842 -16298
rect 14978 -16242 15038 -16236
rect 19870 -16242 19930 -16236
rect 14978 -16246 19930 -16242
rect 23528 -16246 23588 -16240
rect 14978 -16298 14982 -16246
rect 15034 -16298 19874 -16246
rect 19926 -16298 19930 -16246
rect 14978 -16302 19930 -16298
rect 14978 -16308 15038 -16302
rect 19870 -16308 19930 -16302
rect 20368 -16250 23588 -16246
rect 20368 -16302 20378 -16250
rect 20430 -16302 23532 -16250
rect 23584 -16302 23588 -16250
rect 20368 -16306 23588 -16302
rect 23528 -16312 23588 -16306
rect 5116 -16352 5176 -16346
rect 8674 -16350 8734 -16344
rect 10710 -16350 10770 -16344
rect 12746 -16350 12806 -16344
rect 14782 -16350 14842 -16344
rect 16816 -16350 16876 -16344
rect 18854 -16350 18914 -16344
rect 20894 -16350 20954 -16344
rect 23278 -16350 23338 -16344
rect 5116 -16354 8218 -16352
rect 4408 -16356 8218 -16354
rect 4408 -16408 5120 -16356
rect 5172 -16408 6124 -16356
rect 6176 -16408 7136 -16356
rect 7188 -16408 8156 -16356
rect 8208 -16408 8218 -16356
rect 4408 -16412 8218 -16408
rect 8674 -16354 23338 -16350
rect 8674 -16406 8678 -16354
rect 8730 -16406 10714 -16354
rect 10766 -16406 12750 -16354
rect 12802 -16406 14786 -16354
rect 14838 -16406 16820 -16354
rect 16872 -16406 18858 -16354
rect 18910 -16406 20898 -16354
rect 20950 -16406 23282 -16354
rect 23334 -16406 23338 -16354
rect 8674 -16410 23338 -16406
rect 4408 -16414 5458 -16412
rect 2336 -16418 3644 -16414
rect 5116 -16418 5176 -16414
rect 8674 -16416 8734 -16410
rect 10710 -16416 10770 -16410
rect 12746 -16416 12806 -16410
rect 14782 -16416 14842 -16410
rect 16816 -16416 16876 -16410
rect 18854 -16416 18914 -16410
rect 20894 -16416 20954 -16410
rect 23278 -16416 23338 -16410
rect 2336 -16424 2396 -16418
rect 3584 -16424 3644 -16418
rect 2230 -16460 2290 -16454
rect 9692 -16460 9752 -16454
rect 11726 -16460 11786 -16454
rect 13766 -16460 13826 -16454
rect 14978 -16460 15038 -16454
rect 1720 -16464 15038 -16460
rect 1720 -16516 2234 -16464
rect 2286 -16516 9696 -16464
rect 9748 -16516 11730 -16464
rect 11782 -16516 13770 -16464
rect 13822 -16516 14982 -16464
rect 15034 -16516 15038 -16464
rect 1720 -16520 15038 -16516
rect 2230 -16526 2290 -16520
rect 9692 -16526 9752 -16520
rect 11726 -16526 11786 -16520
rect 13766 -16526 13826 -16520
rect 14978 -16526 15038 -16520
rect 15272 -16458 15332 -16452
rect 15272 -16462 16366 -16458
rect 15272 -16514 15276 -16462
rect 15328 -16514 16304 -16462
rect 16356 -16514 16366 -16462
rect 15272 -16518 16366 -16514
rect 16818 -16464 16878 -16458
rect 18854 -16464 18914 -16458
rect 20892 -16464 20952 -16458
rect 23034 -16464 23094 -16458
rect 16818 -16468 23094 -16464
rect 15272 -16524 15332 -16518
rect 16818 -16520 16822 -16468
rect 16874 -16520 18858 -16468
rect 18910 -16520 20896 -16468
rect 20948 -16520 23038 -16468
rect 23090 -16520 23094 -16468
rect 16818 -16524 23094 -16520
rect 16818 -16530 16878 -16524
rect 18854 -16530 18914 -16524
rect 20892 -16530 20952 -16524
rect 23034 -16530 23094 -16524
rect 19366 -17378 19426 -17372
rect 14266 -17382 19426 -17378
rect 3584 -17390 3644 -17384
rect 5622 -17390 5682 -17384
rect 7658 -17390 7718 -17384
rect 9690 -17390 9750 -17384
rect 3584 -17394 9750 -17390
rect 3584 -17446 3588 -17394
rect 3640 -17446 5626 -17394
rect 5678 -17446 7662 -17394
rect 7714 -17446 9694 -17394
rect 9746 -17446 9750 -17394
rect 14266 -17434 14276 -17382
rect 14328 -17434 19370 -17382
rect 19422 -17434 19426 -17382
rect 14266 -17438 19426 -17434
rect 19366 -17444 19426 -17438
rect 19504 -17374 19564 -17368
rect 20386 -17374 20446 -17368
rect 21392 -17374 21452 -17368
rect 19504 -17378 21452 -17374
rect 19504 -17430 19508 -17378
rect 19560 -17430 20390 -17378
rect 20442 -17430 21396 -17378
rect 21448 -17430 21452 -17378
rect 19504 -17434 21452 -17430
rect 19504 -17440 19564 -17434
rect 20386 -17440 20446 -17434
rect 21392 -17440 21452 -17434
rect 21910 -17378 21970 -17372
rect 23162 -17378 23222 -17372
rect 21910 -17382 23222 -17378
rect 21910 -17434 21914 -17382
rect 21966 -17434 23166 -17382
rect 23218 -17434 23222 -17382
rect 21910 -17438 23222 -17434
rect 21910 -17444 21970 -17438
rect 23162 -17444 23222 -17438
rect 3584 -17450 9750 -17446
rect 3584 -17456 3644 -17450
rect 5622 -17456 5682 -17450
rect 7658 -17456 7718 -17450
rect 9690 -17456 9750 -17450
rect 4090 -17492 4150 -17486
rect 9182 -17492 9242 -17486
rect 4090 -17496 9242 -17492
rect 4090 -17548 4094 -17496
rect 4146 -17548 9186 -17496
rect 9238 -17548 9242 -17496
rect 4090 -17552 9242 -17548
rect 4090 -17558 4150 -17552
rect 9182 -17558 9242 -17552
rect 13766 -17506 13826 -17500
rect 21910 -17506 21970 -17500
rect 13766 -17510 21970 -17506
rect 13766 -17562 13770 -17510
rect 13822 -17562 21914 -17510
rect 21966 -17562 21970 -17510
rect 13766 -17566 21970 -17562
rect 13766 -17572 13826 -17566
rect 21910 -17572 21970 -17566
rect 2336 -17594 2396 -17588
rect 5620 -17594 5680 -17588
rect 2336 -17598 5680 -17594
rect 2336 -17650 2340 -17598
rect 2392 -17650 5624 -17598
rect 5676 -17650 5680 -17598
rect 2336 -17654 5680 -17650
rect 2336 -17660 2396 -17654
rect 5620 -17660 5680 -17654
rect 6128 -17600 6188 -17594
rect 7150 -17600 7210 -17594
rect 8164 -17600 8224 -17594
rect 9182 -17600 9242 -17594
rect 10202 -17600 10262 -17594
rect 17314 -17600 17374 -17594
rect 18344 -17600 18404 -17594
rect 19504 -17600 19564 -17594
rect 6128 -17604 19564 -17600
rect 6128 -17656 6132 -17604
rect 6184 -17656 7154 -17604
rect 7206 -17656 8168 -17604
rect 8220 -17656 9186 -17604
rect 9238 -17656 10206 -17604
rect 10258 -17656 17318 -17604
rect 17370 -17656 18348 -17604
rect 18400 -17656 19508 -17604
rect 19560 -17656 19564 -17604
rect 6128 -17660 19564 -17656
rect 6128 -17666 6188 -17660
rect 7150 -17666 7210 -17660
rect 8164 -17666 8224 -17660
rect 9182 -17666 9242 -17660
rect 10202 -17666 10262 -17660
rect 17314 -17666 17374 -17660
rect 18344 -17666 18404 -17660
rect 19504 -17666 19564 -17660
rect 19872 -17600 19932 -17594
rect 23400 -17600 23460 -17594
rect 19872 -17604 23460 -17600
rect 19872 -17656 19876 -17604
rect 19928 -17656 23404 -17604
rect 23456 -17656 23460 -17604
rect 19872 -17660 23460 -17656
rect 19872 -17666 19932 -17660
rect 23400 -17666 23460 -17660
rect 4604 -17694 4664 -17688
rect 6638 -17694 6698 -17688
rect 8674 -17694 8734 -17688
rect 4604 -17698 8734 -17694
rect 4604 -17750 4608 -17698
rect 4660 -17750 6642 -17698
rect 6694 -17750 8678 -17698
rect 8730 -17750 8734 -17698
rect 4604 -17754 8734 -17750
rect 4604 -17760 4664 -17754
rect 6638 -17760 6698 -17754
rect 8674 -17760 8734 -17754
rect 15802 -17704 15862 -17698
rect 19872 -17704 19932 -17698
rect 15802 -17708 19932 -17704
rect 15802 -17760 15806 -17708
rect 15858 -17760 19876 -17708
rect 19928 -17760 19932 -17708
rect 15802 -17764 19932 -17760
rect 15802 -17770 15862 -17764
rect 19872 -17770 19932 -17764
rect 20888 -17702 20948 -17696
rect 23278 -17702 23338 -17696
rect 20888 -17706 23338 -17702
rect 20888 -17758 20892 -17706
rect 20944 -17758 23282 -17706
rect 23334 -17758 23338 -17706
rect 20888 -17762 23338 -17758
rect 20888 -17768 20948 -17762
rect 23278 -17768 23338 -17762
rect 10710 -18612 10770 -18606
rect 12746 -18612 12806 -18606
rect 14782 -18612 14842 -18606
rect 16820 -18612 16880 -18606
rect 4086 -18618 4146 -18612
rect 4996 -18618 5056 -18612
rect 5998 -18618 6058 -18612
rect 7150 -18618 7210 -18612
rect 8160 -18618 8220 -18612
rect 9166 -18618 9226 -18612
rect 10210 -18618 10270 -18612
rect 4086 -18622 10270 -18618
rect 4086 -18674 4090 -18622
rect 4142 -18674 5000 -18622
rect 5052 -18674 6002 -18622
rect 6054 -18674 7154 -18622
rect 7206 -18674 8164 -18622
rect 8216 -18674 9170 -18622
rect 9222 -18674 10214 -18622
rect 10266 -18674 10270 -18622
rect 4086 -18678 10270 -18674
rect 10710 -18616 16880 -18612
rect 10710 -18668 10714 -18616
rect 10766 -18668 12750 -18616
rect 12802 -18668 14786 -18616
rect 14838 -18668 16824 -18616
rect 16876 -18668 16880 -18616
rect 10710 -18672 16880 -18668
rect 10710 -18678 10770 -18672
rect 12746 -18678 12806 -18672
rect 14782 -18678 14842 -18672
rect 16820 -18678 16880 -18672
rect 18856 -18612 18916 -18606
rect 20894 -18612 20954 -18606
rect 18856 -18616 20954 -18612
rect 18856 -18668 18860 -18616
rect 18912 -18668 20898 -18616
rect 20950 -18668 20954 -18616
rect 18856 -18672 20954 -18668
rect 18856 -18678 18916 -18672
rect 20894 -18678 20954 -18672
rect 4086 -18684 4146 -18678
rect 4996 -18684 5056 -18678
rect 5998 -18684 6058 -18678
rect 7150 -18684 7210 -18678
rect 8160 -18684 8220 -18678
rect 9166 -18684 9226 -18678
rect 10210 -18684 10270 -18678
rect 6638 -18720 6698 -18714
rect 16812 -18720 16872 -18714
rect 18852 -18720 18912 -18714
rect 20890 -18720 20950 -18714
rect 6638 -18724 20950 -18720
rect 6638 -18776 6642 -18724
rect 6694 -18776 16816 -18724
rect 16868 -18776 18856 -18724
rect 18908 -18776 20894 -18724
rect 20946 -18776 20950 -18724
rect 6638 -18780 20950 -18776
rect 6638 -18786 6698 -18780
rect 16812 -18786 16872 -18780
rect 18852 -18786 18912 -18780
rect 20890 -18786 20950 -18780
rect 4086 -18834 4146 -18828
rect 6138 -18834 6198 -18828
rect 9164 -18834 9224 -18828
rect 10204 -18834 10264 -18828
rect 11218 -18834 11278 -18828
rect 12226 -18834 12286 -18828
rect 13270 -18834 13330 -18828
rect 14260 -18834 14320 -18828
rect 15278 -18834 15338 -18828
rect 16312 -18834 16372 -18828
rect 19344 -18834 19404 -18828
rect 20382 -18834 20442 -18828
rect 21408 -18834 21468 -18828
rect 4086 -18838 23592 -18834
rect 4086 -18890 4090 -18838
rect 4142 -18890 5128 -18838
rect 5180 -18890 6142 -18838
rect 6194 -18890 9168 -18838
rect 9220 -18890 10208 -18838
rect 10260 -18890 11222 -18838
rect 11274 -18890 12230 -18838
rect 12282 -18890 13274 -18838
rect 13326 -18890 14264 -18838
rect 14316 -18890 15282 -18838
rect 15334 -18890 16316 -18838
rect 16368 -18890 19348 -18838
rect 19400 -18890 20386 -18838
rect 20438 -18890 21412 -18838
rect 21464 -18890 23530 -18838
rect 23582 -18890 23592 -18838
rect 4086 -18894 23592 -18890
rect 4086 -18900 4146 -18894
rect 6138 -18900 6198 -18894
rect 9164 -18900 9224 -18894
rect 10204 -18900 10264 -18894
rect 11218 -18900 11278 -18894
rect 12226 -18900 12286 -18894
rect 13270 -18900 13330 -18894
rect 14260 -18900 14320 -18894
rect 15278 -18900 15338 -18894
rect 16312 -18900 16372 -18894
rect 19344 -18900 19404 -18894
rect 20382 -18900 20442 -18894
rect 21408 -18900 21468 -18894
rect 9688 -18938 9748 -18932
rect 11730 -18938 11790 -18932
rect 13768 -18938 13828 -18932
rect 15802 -18938 15862 -18932
rect 17836 -18936 17896 -18930
rect 19870 -18936 19930 -18930
rect 21912 -18936 21972 -18930
rect 23162 -18936 23222 -18930
rect 2444 -18942 15862 -18938
rect 2444 -18994 2454 -18942
rect 2506 -18994 9692 -18942
rect 9744 -18994 11734 -18942
rect 11786 -18994 13772 -18942
rect 13824 -18994 15806 -18942
rect 15858 -18994 15862 -18942
rect 2444 -18998 15862 -18994
rect 9688 -19004 9748 -18998
rect 11730 -19004 11790 -18998
rect 13768 -19004 13828 -18998
rect 15802 -19004 15862 -18998
rect 16314 -18942 16374 -18936
rect 17336 -18942 17396 -18936
rect 16314 -18946 17396 -18942
rect 16314 -18998 16318 -18946
rect 16370 -18998 17340 -18946
rect 17392 -18998 17396 -18946
rect 16314 -19002 17396 -18998
rect 17836 -18940 23222 -18936
rect 17836 -18992 17840 -18940
rect 17892 -18992 19874 -18940
rect 19926 -18992 21916 -18940
rect 21968 -18992 23166 -18940
rect 23218 -18992 23222 -18940
rect 17836 -18996 23222 -18992
rect 17836 -19002 17896 -18996
rect 19870 -19002 19930 -18996
rect 21912 -19002 21972 -18996
rect 23162 -19002 23222 -18996
rect 16314 -19008 16374 -19002
rect 17336 -19008 17396 -19002
rect 8678 -19840 8738 -19834
rect 12746 -19840 12806 -19834
rect 14780 -19840 14840 -19834
rect 4084 -19846 4144 -19840
rect 5092 -19846 5152 -19840
rect 6106 -19846 6166 -19840
rect 7144 -19846 7204 -19840
rect 8162 -19846 8222 -19840
rect 4084 -19850 8222 -19846
rect 4084 -19902 4088 -19850
rect 4140 -19902 5096 -19850
rect 5148 -19902 6110 -19850
rect 6162 -19902 7148 -19850
rect 7200 -19902 8166 -19850
rect 8218 -19902 8222 -19850
rect 4084 -19906 8222 -19902
rect 8678 -19844 14840 -19840
rect 8678 -19896 8682 -19844
rect 8734 -19896 10718 -19844
rect 10770 -19896 12750 -19844
rect 12802 -19896 14784 -19844
rect 14836 -19896 14840 -19844
rect 8678 -19900 14840 -19896
rect 8678 -19906 8738 -19900
rect 12746 -19906 12806 -19900
rect 14780 -19906 14840 -19900
rect 15802 -19838 15862 -19832
rect 16156 -19838 16216 -19832
rect 15802 -19842 16216 -19838
rect 15802 -19894 15806 -19842
rect 15858 -19894 16160 -19842
rect 16212 -19894 16216 -19842
rect 15802 -19898 16216 -19894
rect 15802 -19904 15862 -19898
rect 16156 -19904 16216 -19898
rect 19874 -19838 19934 -19832
rect 23158 -19838 23218 -19832
rect 19874 -19842 23218 -19838
rect 19874 -19894 19878 -19842
rect 19930 -19894 23162 -19842
rect 23214 -19894 23218 -19842
rect 19874 -19898 23218 -19894
rect 19874 -19904 19934 -19898
rect 23158 -19904 23218 -19898
rect 4084 -19912 4144 -19906
rect 5092 -19912 5152 -19906
rect 6106 -19912 6166 -19906
rect 7144 -19912 7204 -19906
rect 8162 -19912 8222 -19906
rect 2230 -19950 2290 -19944
rect 3586 -19950 3646 -19944
rect 11730 -19950 11790 -19944
rect 13766 -19950 13826 -19944
rect 15798 -19950 15858 -19944
rect 2230 -19954 15858 -19950
rect 2230 -20006 2234 -19954
rect 2286 -20006 3590 -19954
rect 3642 -20006 11734 -19954
rect 11786 -20006 13770 -19954
rect 13822 -20006 15802 -19954
rect 15854 -20006 15858 -19954
rect 2230 -20010 15858 -20006
rect 2230 -20016 2290 -20010
rect 3586 -20016 3646 -20010
rect 11730 -20016 11790 -20010
rect 13766 -20016 13826 -20010
rect 15798 -20016 15858 -20010
rect 15308 -20048 15368 -20042
rect 16346 -20048 16406 -20042
rect 17322 -20048 17382 -20042
rect 18338 -20048 18398 -20042
rect 20364 -20048 20424 -20042
rect 21394 -20048 21454 -20042
rect 15308 -20052 21454 -20048
rect -374 -20074 1646 -20070
rect -374 -20126 -370 -20074
rect -318 -20126 1646 -20074
rect -374 -20130 1646 -20126
rect 4602 -20062 4662 -20056
rect 6640 -20062 6700 -20056
rect 10712 -20062 10772 -20056
rect 4602 -20066 10772 -20062
rect 4602 -20118 4606 -20066
rect 4658 -20118 6644 -20066
rect 6696 -20118 10716 -20066
rect 10768 -20118 10772 -20066
rect 15308 -20104 15312 -20052
rect 15364 -20104 16350 -20052
rect 16402 -20104 17326 -20052
rect 17378 -20104 18342 -20052
rect 18394 -20104 20368 -20052
rect 20420 -20104 21398 -20052
rect 21450 -20104 21454 -20052
rect 15308 -20108 21454 -20104
rect 15308 -20114 15368 -20108
rect 16346 -20114 16406 -20108
rect 17322 -20114 17382 -20108
rect 18338 -20114 18398 -20108
rect 20364 -20114 20424 -20108
rect 21394 -20114 21454 -20108
rect 4602 -20122 10772 -20118
rect 4602 -20128 4662 -20122
rect 6640 -20128 6700 -20122
rect 10712 -20128 10772 -20122
rect -374 -20136 -314 -20130
rect -592 -20160 -532 -20154
rect -1028 -20164 -532 -20160
rect -1028 -20216 -1024 -20164
rect -972 -20216 -588 -20164
rect -536 -20216 -532 -20164
rect 3582 -20160 3642 -20154
rect 5620 -20160 5680 -20154
rect 7660 -20160 7720 -20154
rect 9696 -20160 9756 -20154
rect 15800 -20160 15860 -20154
rect 16150 -20160 16222 -20156
rect 17836 -20160 17896 -20154
rect 19872 -20160 19932 -20154
rect 21908 -20160 21968 -20154
rect 3582 -20164 16160 -20160
rect 2336 -20196 2396 -20190
rect -1028 -20220 -532 -20216
rect -1028 -20226 -968 -20220
rect -592 -20226 -532 -20220
rect 214 -20200 2396 -20196
rect 214 -20252 224 -20200
rect 276 -20252 2340 -20200
rect 2392 -20252 2396 -20200
rect 3582 -20216 3586 -20164
rect 3638 -20216 5624 -20164
rect 5676 -20216 7664 -20164
rect 7716 -20216 9700 -20164
rect 9752 -20212 16160 -20164
rect 16212 -20164 21968 -20160
rect 16212 -20212 17840 -20164
rect 9752 -20216 17840 -20212
rect 17892 -20216 19876 -20164
rect 19928 -20216 21912 -20164
rect 21964 -20216 21968 -20164
rect 3582 -20220 21968 -20216
rect 3582 -20226 3642 -20220
rect 5620 -20226 5680 -20220
rect 7660 -20226 7720 -20220
rect 9696 -20226 9756 -20220
rect 15800 -20226 15860 -20220
rect 17836 -20226 17896 -20220
rect 19872 -20226 19932 -20220
rect 21908 -20226 21968 -20220
rect 214 -20256 2396 -20252
rect 2336 -20262 2396 -20256
rect -1792 -20270 -1732 -20264
rect -1572 -20270 -1512 -20264
rect -918 -20270 -858 -20264
rect -702 -20270 -642 -20264
rect -1792 -20274 -642 -20270
rect -1792 -20326 -1788 -20274
rect -1736 -20326 -1568 -20274
rect -1516 -20326 -914 -20274
rect -862 -20326 -698 -20274
rect -646 -20326 -642 -20274
rect -1792 -20330 -642 -20326
rect -1792 -20336 -1732 -20330
rect -1572 -20336 -1512 -20330
rect -918 -20336 -858 -20330
rect -702 -20336 -642 -20330
rect -2468 -20774 -2408 -20768
rect -2010 -20774 -1950 -20768
rect -1354 -20774 -1294 -20768
rect -2468 -20778 -1294 -20774
rect -2468 -20830 -2464 -20778
rect -2412 -20830 -2006 -20778
rect -1954 -20830 -1350 -20778
rect -1298 -20830 -1294 -20778
rect -2468 -20834 -1294 -20830
rect -2468 -20840 -2408 -20834
rect -2010 -20840 -1950 -20834
rect -1354 -20840 -1294 -20834
rect -810 -20774 -750 -20768
rect -22 -20774 38 -20768
rect -810 -20778 38 -20774
rect -810 -20830 -806 -20778
rect -754 -20830 -18 -20778
rect 34 -20830 38 -20778
rect -810 -20834 38 -20830
rect -810 -20840 -750 -20834
rect -22 -20840 38 -20834
rect -2598 -20896 -2538 -20890
rect -1792 -20896 -1732 -20890
rect -1574 -20896 -1514 -20890
rect -2598 -20900 -1514 -20896
rect -2598 -20952 -2594 -20900
rect -2542 -20952 -1788 -20900
rect -1736 -20952 -1570 -20900
rect -1518 -20952 -1514 -20900
rect -2598 -20956 -1514 -20952
rect -2598 -20962 -2538 -20956
rect -1792 -20962 -1732 -20956
rect -1574 -20962 -1514 -20956
rect -1138 -20894 -1078 -20888
rect -482 -20894 -422 -20888
rect -1138 -20898 -422 -20894
rect -1138 -20950 -1134 -20898
rect -1082 -20950 -478 -20898
rect -426 -20950 -422 -20898
rect -1138 -20954 -422 -20950
rect -1138 -20960 -1078 -20954
rect -482 -20960 -422 -20954
rect -2118 -21020 -2058 -21014
rect -1248 -21020 -1188 -21014
rect -376 -21020 -316 -21014
rect -2118 -21024 -316 -21020
rect -2118 -21076 -2114 -21024
rect -2062 -21076 -1244 -21024
rect -1192 -21076 -372 -21024
rect -320 -21076 -316 -21024
rect 10708 -21064 10768 -21058
rect 12750 -21064 12810 -21058
rect 14782 -21064 14842 -21058
rect 16822 -21064 16882 -21058
rect 23278 -21064 23338 -21058
rect -2118 -21080 -316 -21076
rect 10532 -21068 23338 -21064
rect -2118 -21086 -2058 -21080
rect -1248 -21086 -1188 -21080
rect -376 -21086 -316 -21080
rect 4602 -21084 4662 -21078
rect 6638 -21084 6698 -21078
rect 8676 -21084 8736 -21078
rect 4602 -21088 8736 -21084
rect 4602 -21140 4606 -21088
rect 4658 -21140 6642 -21088
rect 6694 -21140 8680 -21088
rect 8732 -21140 8736 -21088
rect 10532 -21120 10542 -21068
rect 10594 -21120 10712 -21068
rect 10764 -21120 12754 -21068
rect 12806 -21120 14786 -21068
rect 14838 -21120 16826 -21068
rect 16878 -21120 23282 -21068
rect 23334 -21120 23338 -21068
rect 10532 -21124 23338 -21120
rect 10708 -21130 10768 -21124
rect 12750 -21130 12810 -21124
rect 14782 -21130 14842 -21124
rect 16822 -21130 16882 -21124
rect 23278 -21130 23338 -21124
rect -1680 -21146 -1620 -21140
rect 98 -21146 158 -21140
rect -1680 -21150 158 -21146
rect 4602 -21144 8736 -21140
rect 4602 -21150 4662 -21144
rect 6638 -21150 6698 -21144
rect 8676 -21150 8736 -21144
rect -1680 -21202 -1676 -21150
rect -1624 -21202 102 -21150
rect 154 -21202 158 -21150
rect 15800 -21162 15860 -21156
rect 21906 -21162 21966 -21156
rect 23158 -21162 23218 -21156
rect 15800 -21166 23218 -21162
rect -1680 -21206 158 -21202
rect -1680 -21212 -1620 -21206
rect 98 -21212 158 -21206
rect 2448 -21182 2508 -21176
rect 5620 -21182 5680 -21176
rect 2448 -21186 5680 -21182
rect 2448 -21238 2452 -21186
rect 2504 -21238 5624 -21186
rect 5676 -21238 5680 -21186
rect 2448 -21242 5680 -21238
rect 2448 -21248 2508 -21242
rect 5620 -21248 5680 -21242
rect 7144 -21182 7204 -21176
rect 10192 -21182 10252 -21176
rect 7144 -21186 10252 -21182
rect 7144 -21238 7148 -21186
rect 7200 -21238 8170 -21186
rect 8222 -21238 9192 -21186
rect 9244 -21238 10196 -21186
rect 10248 -21238 10252 -21186
rect 15800 -21218 15804 -21166
rect 15856 -21218 21910 -21166
rect 21962 -21218 23162 -21166
rect 23214 -21218 23218 -21166
rect 15800 -21222 23218 -21218
rect 15800 -21228 15860 -21222
rect 21906 -21228 21966 -21222
rect 23158 -21228 23218 -21222
rect 7144 -21242 10252 -21238
rect 7144 -21248 7204 -21242
rect 10192 -21248 10252 -21242
rect -1346 -21260 -1294 -21254
rect 2236 -21262 2242 -21260
rect -1294 -21310 2242 -21262
rect 2236 -21312 2242 -21310
rect 2294 -21312 2300 -21260
rect 10714 -21272 10774 -21266
rect 12742 -21272 12802 -21266
rect 14786 -21272 14846 -21266
rect 16814 -21272 16874 -21266
rect 18852 -21272 18912 -21266
rect 20892 -21272 20952 -21266
rect 4606 -21278 4666 -21272
rect 6642 -21278 6702 -21272
rect 8670 -21278 8730 -21272
rect 10538 -21278 10598 -21272
rect 4606 -21282 10598 -21278
rect -1346 -21318 -1294 -21312
rect 4606 -21334 4610 -21282
rect 4662 -21334 6646 -21282
rect 6698 -21334 8674 -21282
rect 8726 -21334 10542 -21282
rect 10594 -21334 10598 -21282
rect 4606 -21338 10598 -21334
rect 10714 -21276 20952 -21272
rect 10714 -21328 10718 -21276
rect 10770 -21328 12746 -21276
rect 12798 -21328 14790 -21276
rect 14842 -21328 16818 -21276
rect 16870 -21328 18856 -21276
rect 18908 -21328 20896 -21276
rect 20948 -21328 20952 -21276
rect 10714 -21332 20952 -21328
rect 10714 -21338 10774 -21332
rect 12742 -21338 12802 -21332
rect 14786 -21338 14846 -21332
rect 16814 -21338 16874 -21332
rect 18852 -21338 18912 -21332
rect 20892 -21338 20952 -21332
rect 21410 -21268 21470 -21262
rect 23528 -21268 23588 -21262
rect 21410 -21272 23588 -21268
rect 21410 -21324 21414 -21272
rect 21466 -21324 23532 -21272
rect 23584 -21324 23588 -21272
rect 21410 -21328 23588 -21324
rect 21410 -21334 21470 -21328
rect 23528 -21334 23588 -21328
rect 4606 -21344 4666 -21338
rect 6642 -21344 6702 -21338
rect 8670 -21344 8730 -21338
rect 10538 -21344 10598 -21338
rect 3588 -21398 3648 -21392
rect 7656 -21398 7716 -21392
rect 9690 -21398 9750 -21392
rect 17840 -21398 17900 -21392
rect 19870 -21398 19930 -21392
rect 21908 -21396 21968 -21390
rect 23400 -21396 23460 -21390
rect 3588 -21402 19930 -21398
rect 3588 -21454 3592 -21402
rect 3644 -21454 7660 -21402
rect 7712 -21454 9694 -21402
rect 9746 -21454 17844 -21402
rect 17896 -21454 19874 -21402
rect 19926 -21454 19930 -21402
rect 3588 -21458 19930 -21454
rect 20390 -21400 23460 -21396
rect 20390 -21452 20400 -21400
rect 20452 -21452 21912 -21400
rect 21964 -21452 23404 -21400
rect 23456 -21452 23460 -21400
rect 20390 -21456 23460 -21452
rect 3588 -21464 3648 -21458
rect 7656 -21464 7716 -21458
rect 9690 -21464 9750 -21458
rect 17840 -21464 17900 -21458
rect 19870 -21464 19930 -21458
rect 21908 -21462 21968 -21456
rect 23400 -21462 23460 -21456
rect -932 -21480 -872 -21474
rect 262 -21480 322 -21474
rect 952 -21480 1012 -21474
rect -2128 -21484 1012 -21480
rect -2128 -21536 -2118 -21484
rect -2066 -21536 -928 -21484
rect -876 -21536 266 -21484
rect 318 -21536 956 -21484
rect 1008 -21536 1012 -21484
rect -2128 -21540 1012 -21536
rect -932 -21546 -872 -21540
rect 262 -21546 322 -21540
rect 952 -21546 1012 -21540
rect -2670 -21580 -2610 -21574
rect -1678 -21580 -1618 -21574
rect -1380 -21580 -1320 -21574
rect -484 -21580 -424 -21574
rect -188 -21580 -128 -21574
rect -2670 -21584 -128 -21580
rect -2670 -21636 -2666 -21584
rect -2614 -21636 -1674 -21584
rect -1622 -21636 -1376 -21584
rect -1324 -21636 -480 -21584
rect -428 -21636 -184 -21584
rect -132 -21636 -128 -21584
rect -2670 -21640 -128 -21636
rect -2670 -21646 -2610 -21640
rect -1678 -21646 -1618 -21640
rect -1380 -21646 -1320 -21640
rect -484 -21646 -424 -21640
rect -188 -21646 -128 -21640
rect 2336 -22314 2396 -22308
rect 11724 -22314 11784 -22308
rect 13766 -22314 13826 -22308
rect 15802 -22314 15862 -22308
rect 2336 -22318 15862 -22314
rect 2336 -22370 2340 -22318
rect 2392 -22370 11728 -22318
rect 11780 -22370 13770 -22318
rect 13822 -22370 15806 -22318
rect 15858 -22370 15862 -22318
rect 2336 -22374 15862 -22370
rect 2336 -22380 2396 -22374
rect 11724 -22380 11784 -22374
rect 13766 -22380 13826 -22374
rect 15802 -22380 15862 -22374
rect 18856 -22314 18916 -22308
rect 20888 -22314 20948 -22308
rect 23034 -22314 23094 -22308
rect 18856 -22318 23094 -22314
rect 18856 -22370 18860 -22318
rect 18912 -22370 20892 -22318
rect 20944 -22370 23038 -22318
rect 23090 -22370 23094 -22318
rect 18856 -22374 23094 -22370
rect 18856 -22380 18916 -22374
rect 20888 -22380 20948 -22374
rect 23034 -22380 23094 -22374
rect 6140 -22428 6200 -22422
rect 11220 -22428 11280 -22422
rect 6140 -22432 11280 -22428
rect 2230 -22440 2290 -22434
rect 5620 -22440 5680 -22434
rect 2230 -22444 5680 -22440
rect -1829 -22483 -1771 -22477
rect -1225 -22483 -1167 -22477
rect -634 -22483 -576 -22477
rect -1829 -22486 623 -22483
rect -1829 -22538 -1826 -22486
rect -1774 -22538 -1222 -22486
rect -1170 -22538 -631 -22486
rect -579 -22538 -34 -22486
rect 18 -22538 562 -22486
rect 614 -22538 623 -22486
rect 2230 -22496 2234 -22444
rect 2286 -22496 5624 -22444
rect 5676 -22496 5680 -22444
rect 6140 -22484 6144 -22432
rect 6196 -22484 11224 -22432
rect 11276 -22484 11280 -22432
rect 6140 -22488 11280 -22484
rect 6140 -22494 6200 -22488
rect 11220 -22494 11280 -22488
rect 16308 -22424 16368 -22418
rect 21408 -22424 21468 -22418
rect 16308 -22428 21468 -22424
rect 16308 -22480 16312 -22428
rect 16364 -22480 21412 -22428
rect 21464 -22480 21468 -22428
rect 16308 -22484 21468 -22480
rect 16308 -22490 16368 -22484
rect 21408 -22490 21468 -22484
rect 2230 -22500 5680 -22496
rect 2230 -22506 2290 -22500
rect 5620 -22506 5680 -22500
rect -1829 -22541 623 -22538
rect -1829 -22547 -1771 -22541
rect -1225 -22547 -1167 -22541
rect -634 -22547 -576 -22541
rect 4602 -22550 4662 -22544
rect 6638 -22550 6698 -22544
rect 7658 -22550 7718 -22544
rect 8674 -22550 8734 -22544
rect 9694 -22550 9754 -22544
rect 10712 -22550 10772 -22544
rect 12742 -22550 12802 -22544
rect 14780 -22550 14840 -22544
rect 16816 -22550 16876 -22544
rect 17838 -22550 17898 -22544
rect 18858 -22550 18918 -22544
rect 19872 -22550 19932 -22544
rect 20894 -22550 20954 -22544
rect 4602 -22554 20954 -22550
rect 4602 -22606 4606 -22554
rect 4658 -22606 6642 -22554
rect 6694 -22606 7662 -22554
rect 7714 -22606 8678 -22554
rect 8730 -22606 9698 -22554
rect 9750 -22606 10716 -22554
rect 10768 -22606 12746 -22554
rect 12798 -22606 14784 -22554
rect 14836 -22606 16820 -22554
rect 16872 -22606 17842 -22554
rect 17894 -22606 18862 -22554
rect 18914 -22606 19876 -22554
rect 19928 -22606 20898 -22554
rect 20950 -22606 20954 -22554
rect -2542 -22614 -2482 -22608
rect -1532 -22614 -1472 -22608
rect -934 -22614 -874 -22608
rect -340 -22614 -280 -22608
rect 258 -22614 318 -22608
rect -2542 -22618 318 -22614
rect 4602 -22610 20954 -22606
rect 4602 -22616 4662 -22610
rect 6638 -22616 6698 -22610
rect 7658 -22616 7718 -22610
rect 8674 -22616 8734 -22610
rect 9694 -22616 9754 -22610
rect 10712 -22616 10772 -22610
rect 12742 -22616 12802 -22610
rect 14780 -22616 14840 -22610
rect 16816 -22616 16876 -22610
rect 17838 -22616 17898 -22610
rect 18858 -22616 18918 -22610
rect 19872 -22616 19932 -22610
rect 20894 -22616 20954 -22610
rect -2542 -22670 -2538 -22618
rect -2486 -22670 -2122 -22618
rect -2070 -22670 -1528 -22618
rect -1476 -22670 -930 -22618
rect -878 -22670 -336 -22618
rect -284 -22670 262 -22618
rect 314 -22670 318 -22618
rect -2542 -22674 318 -22670
rect -2542 -22680 -2482 -22674
rect -1532 -22680 -1472 -22674
rect -934 -22680 -874 -22674
rect -340 -22680 -280 -22674
rect 258 -22680 318 -22674
rect 6256 -22644 6316 -22638
rect 7140 -22644 7200 -22638
rect 8162 -22644 8222 -22638
rect 10204 -22644 10264 -22638
rect 6256 -22648 10264 -22644
rect 6256 -22700 6260 -22648
rect 6312 -22700 7144 -22648
rect 7196 -22700 8166 -22648
rect 8218 -22700 10208 -22648
rect 10260 -22700 10264 -22648
rect 6256 -22704 10264 -22700
rect 6256 -22710 6316 -22704
rect 7140 -22710 7200 -22704
rect 8162 -22710 8222 -22704
rect 10204 -22710 10264 -22704
rect 17326 -22644 17386 -22638
rect 18346 -22644 18406 -22638
rect 19360 -22644 19420 -22638
rect 20396 -22644 20456 -22638
rect 17326 -22648 20456 -22644
rect 17326 -22700 17330 -22648
rect 17382 -22700 18350 -22648
rect 18402 -22700 19364 -22648
rect 19416 -22700 20400 -22648
rect 20452 -22700 20456 -22648
rect 17326 -22704 20456 -22700
rect 17326 -22710 17386 -22704
rect 18346 -22710 18406 -22704
rect 19360 -22710 19420 -22704
rect 20396 -22710 20456 -22704
rect -1974 -22722 -1914 -22716
rect -1676 -22722 -1616 -22716
rect -1376 -22722 -1316 -22716
rect -1082 -22722 -1022 -22716
rect -786 -22722 -726 -22716
rect -486 -22722 -426 -22716
rect -184 -22722 -124 -22716
rect 106 -22722 166 -22716
rect 410 -22722 470 -22716
rect -1974 -22726 1142 -22722
rect -1974 -22778 -1970 -22726
rect -1918 -22778 -1672 -22726
rect -1620 -22778 -1372 -22726
rect -1320 -22778 -1078 -22726
rect -1026 -22778 -782 -22726
rect -730 -22778 -482 -22726
rect -430 -22778 -180 -22726
rect -128 -22778 110 -22726
rect 162 -22778 414 -22726
rect 466 -22778 1080 -22726
rect 1132 -22778 1142 -22726
rect -1974 -22782 1142 -22778
rect -1974 -22788 -1914 -22782
rect -1676 -22788 -1616 -22782
rect -1376 -22788 -1316 -22782
rect -1082 -22788 -1022 -22782
rect -786 -22788 -726 -22782
rect -486 -22788 -426 -22782
rect -184 -22788 -124 -22782
rect 106 -22788 166 -22782
rect 410 -22788 470 -22782
rect 1976 -23544 2036 -23538
rect 2568 -23544 2628 -23538
rect 3082 -23544 3142 -23538
rect 3580 -23544 3640 -23538
rect 5622 -23544 5682 -23538
rect 7654 -23544 7714 -23538
rect 9686 -23544 9746 -23538
rect 13944 -23544 14016 -23542
rect 15800 -23544 15860 -23538
rect 17834 -23544 17894 -23538
rect 19868 -23544 19928 -23538
rect 21910 -23544 21970 -23538
rect 22422 -23544 22482 -23538
rect 22928 -23544 22988 -23538
rect 1544 -23546 22988 -23544
rect 1400 -23548 13954 -23546
rect 1400 -23600 1980 -23548
rect 2032 -23600 2572 -23548
rect 2624 -23600 3086 -23548
rect 3138 -23600 3584 -23548
rect 3636 -23600 5626 -23548
rect 5678 -23600 7658 -23548
rect 7710 -23600 9690 -23548
rect 9742 -23600 11594 -23548
rect 11646 -23598 13954 -23548
rect 14006 -23548 22988 -23546
rect 14006 -23598 15804 -23548
rect 11646 -23600 15804 -23598
rect 15856 -23600 17838 -23548
rect 17890 -23600 19872 -23548
rect 19924 -23600 21914 -23548
rect 21966 -23600 22426 -23548
rect 22478 -23600 22932 -23548
rect 22984 -23600 22988 -23548
rect 1400 -23604 22988 -23600
rect 1400 -23606 1636 -23604
rect -8254 -23620 -3036 -23616
rect -8254 -23672 -8250 -23620
rect -8198 -23672 -6364 -23620
rect -6312 -23672 -4494 -23620
rect -4442 -23672 -3036 -23620
rect -8254 -23676 -3036 -23672
rect -2670 -23620 -2610 -23614
rect -1976 -23620 -1916 -23614
rect -1080 -23620 -1020 -23614
rect -786 -23620 -726 -23614
rect 108 -23620 168 -23614
rect 410 -23620 470 -23614
rect -2670 -23624 470 -23620
rect -2670 -23676 -2666 -23624
rect -2614 -23676 -1972 -23624
rect -1920 -23676 -1076 -23624
rect -1024 -23676 -782 -23624
rect -730 -23676 112 -23624
rect 164 -23676 414 -23624
rect 466 -23676 470 -23624
rect -8254 -23682 -8194 -23676
rect -6368 -23682 -6308 -23676
rect -4498 -23682 -4438 -23676
rect -2670 -23680 470 -23676
rect -2670 -23686 -2610 -23680
rect -1976 -23686 -1916 -23680
rect -1080 -23686 -1020 -23680
rect -786 -23686 -726 -23680
rect 108 -23686 168 -23680
rect 410 -23686 470 -23680
rect -8402 -23724 -8342 -23718
rect -6366 -23724 -6306 -23718
rect -4330 -23724 -4270 -23718
rect -8402 -23728 -4270 -23724
rect -8402 -23780 -8398 -23728
rect -8346 -23780 -6362 -23728
rect -6310 -23780 -4326 -23728
rect -4274 -23780 -4270 -23728
rect -8402 -23784 -4270 -23780
rect -8402 -23790 -8342 -23784
rect -6366 -23790 -6306 -23784
rect -4330 -23790 -4270 -23784
rect -1530 -23728 -1470 -23722
rect -336 -23728 -276 -23722
rect -1530 -23732 1018 -23728
rect -1530 -23784 -1526 -23732
rect -1474 -23784 -332 -23732
rect -280 -23784 956 -23732
rect 1008 -23784 1018 -23732
rect -1530 -23788 1018 -23784
rect -1530 -23794 -1470 -23788
rect -336 -23794 -276 -23788
rect -7384 -23836 -7324 -23830
rect -7384 -23840 -5280 -23836
rect -7384 -23892 -7380 -23840
rect -7328 -23892 -5342 -23840
rect -5290 -23892 -5280 -23840
rect -7384 -23896 -5280 -23892
rect -7384 -23902 -7324 -23896
rect -1828 -24712 -1768 -24706
rect -1234 -24712 -1174 -24706
rect -634 -24712 -574 -24706
rect -40 -24712 20 -24706
rect 554 -24712 614 -24706
rect 1400 -24712 1460 -23606
rect 1976 -23610 2036 -23604
rect 2568 -23610 2628 -23604
rect 3082 -23610 3142 -23604
rect 3580 -23610 3640 -23604
rect 5622 -23610 5682 -23604
rect 7654 -23610 7714 -23604
rect 9686 -23610 9746 -23604
rect 15800 -23610 15860 -23604
rect 17834 -23610 17894 -23604
rect 19868 -23610 19928 -23604
rect 21910 -23610 21970 -23604
rect 22422 -23610 22482 -23604
rect 22928 -23610 22988 -23604
rect 6130 -23656 6190 -23650
rect 7142 -23656 7202 -23650
rect 8156 -23656 8216 -23650
rect 11068 -23656 11128 -23650
rect 6130 -23660 11128 -23656
rect 6130 -23712 6134 -23660
rect 6186 -23712 7146 -23660
rect 7198 -23712 8160 -23660
rect 8212 -23712 11072 -23660
rect 11124 -23712 11128 -23660
rect 6130 -23716 11128 -23712
rect 6130 -23722 6190 -23716
rect 7142 -23722 7202 -23716
rect 8156 -23722 8216 -23716
rect 11068 -23722 11128 -23716
rect 11728 -23658 11788 -23648
rect 11728 -23710 11732 -23658
rect 11784 -23710 11788 -23658
rect 2110 -23762 2170 -23756
rect 4096 -23762 4156 -23756
rect 5118 -23762 5178 -23756
rect 7656 -23762 7716 -23756
rect 8168 -23762 8228 -23756
rect 9186 -23762 9246 -23756
rect 9692 -23762 9752 -23756
rect 10198 -23762 10258 -23756
rect 11210 -23762 11270 -23756
rect 11728 -23762 11788 -23710
rect 12356 -23658 12416 -23652
rect 13402 -23658 13462 -23652
rect 17330 -23658 17390 -23652
rect 18348 -23658 18408 -23652
rect 12356 -23662 19424 -23658
rect 12356 -23714 12360 -23662
rect 12412 -23714 13406 -23662
rect 13458 -23714 17334 -23662
rect 17386 -23714 18352 -23662
rect 18404 -23714 19362 -23662
rect 19414 -23714 19424 -23662
rect 12356 -23718 19424 -23714
rect 12356 -23724 12416 -23718
rect 13402 -23724 13462 -23718
rect 17330 -23724 17390 -23718
rect 18348 -23724 18408 -23718
rect 12230 -23762 12290 -23756
rect 13252 -23762 13312 -23756
rect 13764 -23762 13824 -23756
rect 14270 -23762 14330 -23756
rect 15288 -23762 15348 -23756
rect 15800 -23762 15860 -23756
rect 16308 -23762 16368 -23756
rect 20380 -23762 20440 -23756
rect 21382 -23762 21442 -23756
rect 2110 -23766 21442 -23762
rect 2110 -23818 2114 -23766
rect 2166 -23818 4100 -23766
rect 4152 -23818 5122 -23766
rect 5174 -23818 7660 -23766
rect 7712 -23818 8172 -23766
rect 8224 -23818 9190 -23766
rect 9242 -23818 9696 -23766
rect 9748 -23818 10202 -23766
rect 10254 -23818 11214 -23766
rect 11266 -23818 12234 -23766
rect 12286 -23818 13256 -23766
rect 13308 -23818 13768 -23766
rect 13820 -23818 14274 -23766
rect 14326 -23818 15292 -23766
rect 15344 -23818 15804 -23766
rect 15856 -23818 16312 -23766
rect 16364 -23818 20384 -23766
rect 20436 -23818 21386 -23766
rect 21438 -23818 21442 -23766
rect 2110 -23822 21442 -23818
rect 2110 -23828 2170 -23822
rect 4096 -23828 4156 -23822
rect 5118 -23828 5178 -23822
rect 7656 -23828 7716 -23822
rect 8168 -23828 8228 -23822
rect 9186 -23828 9246 -23822
rect 9692 -23828 9752 -23822
rect 10198 -23828 10258 -23822
rect 11210 -23828 11270 -23822
rect 12230 -23828 12290 -23822
rect 13252 -23828 13312 -23822
rect 13764 -23828 13824 -23822
rect 14270 -23828 14330 -23822
rect 15288 -23828 15348 -23822
rect 15800 -23828 15860 -23822
rect 16308 -23828 16368 -23822
rect 20380 -23828 20440 -23822
rect 21382 -23828 21442 -23822
rect 1704 -23866 1764 -23860
rect 6132 -23866 6192 -23860
rect 6636 -23866 6696 -23860
rect 7152 -23866 7212 -23860
rect 8674 -23866 8734 -23860
rect 10712 -23866 10772 -23860
rect 12748 -23866 12808 -23860
rect 14784 -23866 14844 -23860
rect 16816 -23866 16876 -23860
rect 17338 -23866 17398 -23860
rect 17838 -23866 17898 -23860
rect 18346 -23866 18406 -23860
rect 18854 -23866 18914 -23860
rect 19204 -23866 19264 -23860
rect 23806 -23866 23866 -23860
rect 1704 -23870 23866 -23866
rect 1704 -23922 1708 -23870
rect 1760 -23922 6136 -23870
rect 6188 -23922 6640 -23870
rect 6692 -23922 7156 -23870
rect 7208 -23922 8678 -23870
rect 8730 -23922 10716 -23870
rect 10768 -23922 12752 -23870
rect 12804 -23922 14788 -23870
rect 14840 -23922 16820 -23870
rect 16872 -23922 17342 -23870
rect 17394 -23922 17842 -23870
rect 17894 -23922 18350 -23870
rect 18402 -23922 18858 -23870
rect 18910 -23922 19208 -23870
rect 19260 -23922 23810 -23870
rect 23862 -23922 23866 -23870
rect 1704 -23926 23866 -23922
rect 1704 -23932 1764 -23926
rect 6132 -23932 6192 -23926
rect 6636 -23932 6696 -23926
rect 7152 -23932 7212 -23926
rect 8674 -23932 8734 -23926
rect 10712 -23932 10772 -23926
rect 12748 -23932 12808 -23926
rect 14784 -23932 14844 -23926
rect 16816 -23932 16876 -23926
rect 17338 -23932 17398 -23926
rect 17838 -23932 17898 -23926
rect 18346 -23932 18406 -23926
rect 18854 -23932 18914 -23926
rect 19204 -23932 19264 -23926
rect 23806 -23932 23866 -23926
rect -7382 -24718 -7322 -24712
rect -1828 -24716 1460 -24712
rect -7382 -24722 -5286 -24718
rect -7382 -24774 -7378 -24722
rect -7326 -24774 -5348 -24722
rect -5296 -24774 -5286 -24722
rect -7382 -24778 -5286 -24774
rect -1828 -24768 -1824 -24716
rect -1772 -24768 -1230 -24716
rect -1178 -24768 -630 -24716
rect -578 -24768 -36 -24716
rect 16 -24768 558 -24716
rect 610 -24768 1460 -24716
rect -1828 -24772 1460 -24768
rect -1828 -24778 -1768 -24772
rect -1234 -24778 -1174 -24772
rect -634 -24778 -574 -24772
rect -40 -24778 20 -24772
rect 554 -24778 614 -24772
rect -7382 -24784 -7322 -24778
rect 11730 -24798 11790 -24792
rect 13766 -24798 13826 -24792
rect -1534 -24806 -1474 -24800
rect -936 -24806 -876 -24800
rect -338 -24806 -278 -24800
rect 262 -24806 322 -24800
rect -2432 -24810 322 -24806
rect -8400 -24820 -8340 -24814
rect -4332 -24820 -4272 -24814
rect -3202 -24820 -3142 -24814
rect -8400 -24824 -3142 -24820
rect -8400 -24876 -8396 -24824
rect -8344 -24876 -4328 -24824
rect -4276 -24876 -3198 -24824
rect -3146 -24876 -3142 -24824
rect -2432 -24862 -2422 -24810
rect -2370 -24862 -1530 -24810
rect -1478 -24862 -932 -24810
rect -880 -24862 -334 -24810
rect -282 -24862 266 -24810
rect 318 -24862 322 -24810
rect -2432 -24866 322 -24862
rect 11730 -24802 13826 -24798
rect 11730 -24854 11734 -24802
rect 11786 -24854 13770 -24802
rect 13822 -24854 13826 -24802
rect 11730 -24858 13826 -24854
rect 11730 -24864 11790 -24858
rect 13766 -24864 13826 -24858
rect -1534 -24872 -1474 -24866
rect -936 -24872 -876 -24866
rect -338 -24872 -278 -24866
rect 262 -24872 322 -24866
rect -8400 -24880 -3142 -24876
rect -8400 -24886 -8340 -24880
rect -4332 -24886 -4272 -24880
rect -3202 -24886 -3142 -24880
rect -1978 -24914 -1918 -24908
rect -1680 -24914 -1620 -24908
rect -1384 -24914 -1324 -24908
rect -1080 -24914 -1020 -24908
rect -784 -24914 -724 -24908
rect -486 -24914 -426 -24908
rect -190 -24914 -130 -24908
rect 106 -24914 166 -24908
rect 410 -24914 470 -24908
rect 1076 -24914 1136 -24908
rect -1978 -24918 1136 -24914
rect -9538 -24926 -9478 -24920
rect -6366 -24926 -6306 -24920
rect -9538 -24930 -6306 -24926
rect -9538 -24982 -9534 -24930
rect -9482 -24982 -6362 -24930
rect -6310 -24982 -6306 -24930
rect -1978 -24970 -1974 -24918
rect -1922 -24970 -1676 -24918
rect -1624 -24970 -1380 -24918
rect -1328 -24970 -1076 -24918
rect -1024 -24970 -780 -24918
rect -728 -24970 -482 -24918
rect -430 -24970 -186 -24918
rect -134 -24970 110 -24918
rect 162 -24970 414 -24918
rect 466 -24970 1080 -24918
rect 1132 -24970 1136 -24918
rect -1978 -24974 1136 -24970
rect -1978 -24980 -1918 -24974
rect -1680 -24980 -1620 -24974
rect -1384 -24980 -1324 -24974
rect -1080 -24980 -1020 -24974
rect -784 -24980 -724 -24974
rect -486 -24980 -426 -24974
rect -190 -24980 -130 -24974
rect 106 -24980 166 -24974
rect 410 -24980 470 -24974
rect 1076 -24980 1136 -24974
rect -9538 -24986 -6306 -24982
rect -9538 -24992 -9478 -24986
rect -6366 -24992 -6306 -24986
rect 3580 -24998 3640 -24992
rect 5618 -24998 5678 -24992
rect 7656 -24998 7716 -24992
rect 9688 -24998 9748 -24992
rect 11726 -24998 11786 -24992
rect 13760 -24998 13820 -24992
rect 15800 -24998 15860 -24992
rect 17834 -24998 17894 -24992
rect 19868 -24998 19928 -24992
rect 21906 -24998 21966 -24992
rect 23648 -24998 23708 -24992
rect 3580 -25002 23708 -24998
rect 3580 -25054 3584 -25002
rect 3636 -25054 5622 -25002
rect 5674 -25054 7660 -25002
rect 7712 -25054 9692 -25002
rect 9744 -25054 11730 -25002
rect 11782 -25054 13764 -25002
rect 13816 -25054 15804 -25002
rect 15856 -25054 17838 -25002
rect 17890 -25054 19872 -25002
rect 19924 -25054 21910 -25002
rect 21962 -25054 23652 -25002
rect 23704 -25054 23708 -25002
rect 3580 -25058 23708 -25054
rect 3580 -25064 3640 -25058
rect 5618 -25064 5678 -25058
rect 7656 -25064 7716 -25058
rect 9688 -25064 9748 -25058
rect 11726 -25064 11786 -25058
rect 13760 -25064 13820 -25058
rect 15800 -25064 15860 -25058
rect 17834 -25064 17894 -25058
rect 19868 -25064 19928 -25058
rect 21906 -25064 21966 -25058
rect 23648 -25064 23708 -25058
rect 2568 -25096 2628 -25090
rect 4598 -25096 4658 -25090
rect 6636 -25096 6696 -25090
rect 8672 -25096 8732 -25090
rect 10708 -25096 10768 -25090
rect 12744 -25096 12804 -25090
rect 14778 -25096 14838 -25090
rect 16814 -25096 16874 -25090
rect 18854 -25096 18914 -25090
rect 20888 -25096 20948 -25090
rect 22924 -25096 22984 -25090
rect 2568 -25100 22984 -25096
rect 2568 -25152 2572 -25100
rect 2624 -25152 4602 -25100
rect 4654 -25152 6640 -25100
rect 6692 -25152 8676 -25100
rect 8728 -25152 10712 -25100
rect 10764 -25152 12748 -25100
rect 12800 -25152 14782 -25100
rect 14834 -25152 16818 -25100
rect 16870 -25152 18858 -25100
rect 18910 -25152 20892 -25100
rect 20944 -25152 22928 -25100
rect 22980 -25152 22984 -25100
rect 2568 -25156 22984 -25152
rect 2568 -25162 2628 -25156
rect 4598 -25162 4658 -25156
rect 6636 -25162 6696 -25156
rect 8672 -25162 8732 -25156
rect 10708 -25162 10768 -25156
rect 12744 -25162 12804 -25156
rect 14778 -25162 14838 -25156
rect 16814 -25162 16874 -25156
rect 18854 -25162 18914 -25156
rect 20888 -25162 20948 -25156
rect 22924 -25162 22984 -25156
rect -2670 -25840 -2610 -25834
rect -1680 -25840 -1620 -25834
rect -1382 -25840 -1322 -25834
rect -486 -25840 -426 -25834
rect -184 -25840 -124 -25834
rect -2670 -25844 -124 -25840
rect -7896 -25870 -7836 -25864
rect -6870 -25870 -6810 -25864
rect -5846 -25870 -5786 -25864
rect -7896 -25874 -4880 -25870
rect -7896 -25926 -7892 -25874
rect -7840 -25926 -6866 -25874
rect -6814 -25926 -5842 -25874
rect -5790 -25926 -4942 -25874
rect -4890 -25926 -4880 -25874
rect -2670 -25896 -2666 -25844
rect -2614 -25896 -1676 -25844
rect -1624 -25896 -1378 -25844
rect -1326 -25896 -482 -25844
rect -430 -25896 -180 -25844
rect -128 -25896 -124 -25844
rect -2670 -25900 -124 -25896
rect -2670 -25906 -2610 -25900
rect -1680 -25906 -1620 -25900
rect -1382 -25906 -1322 -25900
rect -486 -25906 -426 -25900
rect -184 -25906 -124 -25900
rect -7896 -25930 -4880 -25926
rect -7896 -25936 -7836 -25930
rect -6870 -25936 -6810 -25930
rect -5846 -25936 -5786 -25930
rect -2126 -25940 -2066 -25934
rect -938 -25940 -878 -25934
rect 258 -25940 318 -25934
rect 952 -25940 1012 -25934
rect -2126 -25944 1012 -25940
rect -2126 -25996 -2122 -25944
rect -2070 -25996 -934 -25944
rect -882 -25996 262 -25944
rect 314 -25996 956 -25944
rect 1008 -25996 1012 -25944
rect -2126 -26000 1012 -25996
rect -2126 -26006 -2066 -26000
rect -938 -26006 -878 -26000
rect 258 -26006 318 -26000
rect 952 -26006 1012 -26000
rect -7518 -26485 23968 -26430
rect -7518 -26495 -7440 -26485
rect 23896 -26495 23968 -26485
rect -7518 -26611 -7446 -26495
rect 23902 -26611 23968 -26495
rect -7518 -26621 -7440 -26611
rect 23896 -26621 23968 -26611
rect -7518 -26676 23968 -26621
rect -12216 -26818 -11616 -26806
rect -12216 -26844 -12184 -26818
rect -11648 -26844 -11616 -26818
rect -12216 -27088 -12198 -26844
rect -11634 -27088 -11616 -26844
rect -12216 -27114 -12184 -27088
rect -11648 -27114 -11616 -27088
rect -12216 -27126 -11616 -27114
rect 24216 -26818 24816 -26806
rect 24216 -26844 24248 -26818
rect 24784 -26844 24816 -26818
rect 24216 -27088 24234 -26844
rect 24798 -27088 24816 -26844
rect 24216 -27114 24248 -27088
rect 24784 -27114 24816 -27088
rect 24216 -27126 24816 -27114
<< via2 >>
rect 516 1588 1052 1614
rect 516 1344 1052 1588
rect 516 1318 1052 1344
rect 24148 1588 24684 1614
rect 24148 1344 24684 1588
rect 24148 1318 24684 1344
rect 4065 1059 4075 1195
rect 4075 1059 20831 1195
rect 20831 1059 20841 1195
rect -12010 -11202 -11954 -11200
rect -12010 -11254 -12008 -11202
rect -12008 -11254 -11956 -11202
rect -11956 -11254 -11954 -11202
rect -12010 -11256 -11954 -11254
rect -10216 -11202 -10160 -11200
rect -10216 -11254 -10214 -11202
rect -10214 -11254 -10162 -11202
rect -10162 -11254 -10160 -11202
rect -10216 -11256 -10160 -11254
rect -7616 -11202 -7560 -11200
rect -7616 -11254 -7614 -11202
rect -7614 -11254 -7562 -11202
rect -7562 -11254 -7560 -11202
rect -7616 -11256 -7560 -11254
rect -5016 -11200 -4960 -11198
rect -5016 -11252 -5014 -11200
rect -5014 -11252 -4962 -11200
rect -4962 -11252 -4960 -11200
rect -5016 -11254 -4960 -11252
rect -2416 -11200 -2360 -11198
rect -2416 -11252 -2414 -11200
rect -2414 -11252 -2362 -11200
rect -2362 -11252 -2360 -11200
rect -2416 -11254 -2360 -11252
rect -612 -11200 -556 -11198
rect -612 -11252 -610 -11200
rect -610 -11252 -558 -11200
rect -558 -11252 -556 -11200
rect -612 -11254 -556 -11252
rect 2344 -7700 2400 -7644
rect 1722 -10196 1778 -10140
rect -7440 -26495 23896 -26485
rect -7440 -26611 23896 -26495
rect -7440 -26621 23896 -26611
rect -12184 -26844 -11648 -26818
rect -12184 -27088 -11648 -26844
rect -12184 -27114 -11648 -27088
rect 24248 -26844 24784 -26818
rect 24248 -27088 24784 -26844
rect 24248 -27114 24784 -27088
<< metal3 >>
rect 474 1614 1094 1621
rect 474 1578 516 1614
rect 1052 1578 1094 1614
rect 474 1354 512 1578
rect 1056 1354 1094 1578
rect 474 1318 516 1354
rect 1052 1318 1094 1354
rect 474 1311 1094 1318
rect 24106 1614 24726 1621
rect 24106 1578 24148 1614
rect 24684 1578 24726 1614
rect 24106 1354 24144 1578
rect 24688 1354 24726 1578
rect 24106 1318 24148 1354
rect 24684 1318 24726 1354
rect 24106 1311 24726 1318
rect 3998 1199 20878 1266
rect 3998 1055 4061 1199
rect 20845 1055 20878 1199
rect 3998 1000 20878 1055
rect 3998 998 8352 1000
rect -10238 -1378 -10138 32
rect -11658 -1478 -8642 -1378
rect -10238 -2894 -10138 -1478
rect -7638 -2894 -7538 48
rect -6524 -1478 -6042 -1378
rect -5038 -2894 -4938 26
rect -2438 -1378 -2338 22
rect -3924 -1478 -818 -1378
rect -2438 -2894 -2338 -1478
rect -11678 -3978 -8642 -3878
rect -6524 -3978 -6042 -3878
rect -3924 -3978 -812 -3878
rect -10238 -5394 -10138 -4982
rect -7638 -5394 -7538 -4982
rect -5038 -5394 -4938 -4982
rect -2438 -5394 -2338 -4982
rect -11678 -6478 -8642 -6378
rect -6524 -6478 -6042 -6378
rect -3924 -6478 -850 -6378
rect -10238 -8878 -10138 -7482
rect -11674 -8978 -8642 -8878
rect -12032 -11200 -11932 -10854
rect -12032 -11256 -12010 -11200
rect -11954 -11256 -11932 -11200
rect -12032 -11278 -11932 -11256
rect -10238 -11200 -10138 -8978
rect -10238 -11256 -10216 -11200
rect -10160 -11256 -10138 -11200
rect -10238 -11278 -10138 -11256
rect -7638 -11200 -7538 -7482
rect -6524 -8978 -6042 -8878
rect -7638 -11256 -7616 -11200
rect -7560 -11256 -7538 -11200
rect -7638 -11278 -7538 -11256
rect -5038 -11198 -4938 -7482
rect -2438 -8878 -2338 -7482
rect -1749 -7622 -1651 -7617
rect -1750 -7640 2422 -7622
rect -1750 -7704 -1732 -7640
rect -1668 -7644 2422 -7640
rect -1668 -7700 2344 -7644
rect 2400 -7700 2422 -7644
rect -1668 -7704 2422 -7700
rect -1750 -7722 2422 -7704
rect -1749 -7727 -1651 -7722
rect -3924 -8978 -844 -8878
rect -5038 -11254 -5016 -11198
rect -4960 -11254 -4938 -11198
rect -5038 -11276 -4938 -11254
rect -2438 -11198 -2338 -8978
rect -1089 -10118 -991 -10113
rect -1090 -10136 1800 -10118
rect -1090 -10200 -1072 -10136
rect -1008 -10140 1800 -10136
rect -1008 -10196 1722 -10140
rect 1778 -10196 1800 -10140
rect -1008 -10200 1800 -10196
rect -1090 -10218 1800 -10200
rect -1089 -10223 -991 -10218
rect -2438 -11254 -2416 -11198
rect -2360 -11254 -2338 -11198
rect -2438 -11276 -2338 -11254
rect -634 -11198 -534 -10856
rect -634 -11254 -612 -11198
rect -556 -11254 -534 -11198
rect -634 -11276 -534 -11254
rect -7518 -26481 23968 -26430
rect -7518 -26625 -7444 -26481
rect 23900 -26625 23968 -26481
rect -7518 -26676 23968 -26625
rect -12226 -26818 -11606 -26811
rect -12226 -26854 -12184 -26818
rect -11648 -26854 -11606 -26818
rect -12226 -27078 -12188 -26854
rect -11644 -27078 -11606 -26854
rect -12226 -27114 -12184 -27078
rect -11648 -27114 -11606 -27078
rect -12226 -27121 -11606 -27114
rect 24206 -26818 24826 -26811
rect 24206 -26854 24248 -26818
rect 24784 -26854 24826 -26818
rect 24206 -27078 24244 -26854
rect 24788 -27078 24826 -26854
rect 24206 -27114 24248 -27078
rect 24784 -27114 24826 -27078
rect 24206 -27121 24826 -27114
<< via3 >>
rect 512 1354 516 1578
rect 516 1354 1052 1578
rect 1052 1354 1056 1578
rect 24144 1354 24148 1578
rect 24148 1354 24684 1578
rect 24684 1354 24688 1578
rect 4061 1195 20845 1199
rect 4061 1059 4065 1195
rect 4065 1059 20841 1195
rect 20841 1059 20845 1195
rect 4061 1055 20845 1059
rect -1732 -7704 -1668 -7640
rect -1072 -10200 -1008 -10136
rect -7444 -26485 23900 -26481
rect -7444 -26621 -7440 -26485
rect -7440 -26621 23896 -26485
rect 23896 -26621 23900 -26485
rect -7444 -26625 23900 -26621
rect -12188 -27078 -12184 -26854
rect -12184 -27078 -11648 -26854
rect -11648 -27078 -11644 -26854
rect 24244 -27078 24248 -26854
rect 24248 -27078 24784 -26854
rect 24784 -27078 24788 -26854
<< metal4 >>
rect -12400 1578 25000 1800
rect -12400 1354 512 1578
rect 1056 1354 24144 1578
rect 24688 1354 25000 1578
rect -12400 1199 25000 1354
rect -12400 1055 4061 1199
rect 20845 1055 25000 1199
rect -12400 1000 25000 1055
rect -12032 226 -186 326
rect -12032 -10566 -11932 226
rect -11680 -10566 -11580 226
rect -10230 -220 -992 -120
rect -10230 -542 -10130 -220
rect -5000 -566 -4900 -220
rect -7608 -2622 -7508 -2200
rect -2424 -2622 -2324 -2240
rect -11478 -2722 -2324 -2622
rect -11478 -7622 -11378 -2722
rect -10238 -3078 -10138 -2722
rect -5000 -3078 -4900 -2722
rect -7622 -5122 -7522 -4754
rect -2432 -5122 -2332 -4746
rect -1092 -5122 -992 -220
rect -10246 -5222 -992 -5122
rect -10246 -5600 -10146 -5222
rect -5008 -5592 -4908 -5222
rect -7630 -7622 -7530 -7266
rect -2440 -7622 -2340 -7242
rect -11478 -7640 -1650 -7622
rect -11478 -7704 -1732 -7640
rect -1668 -7704 -1650 -7640
rect -11478 -7722 -1650 -7704
rect -10254 -8080 -10154 -7722
rect -5008 -8096 -4908 -7722
rect -7646 -10118 -7546 -9780
rect -2440 -10118 -2340 -9786
rect -1092 -10118 -992 -5222
rect -7646 -10136 -990 -10118
rect -7646 -10200 -1072 -10136
rect -1008 -10200 -990 -10136
rect -7646 -10218 -990 -10200
rect -636 -10566 -536 226
rect -286 -10566 -186 226
rect -12032 -10666 -186 -10566
rect -12032 -10668 -11932 -10666
rect -11680 -10668 -11580 -10666
rect -636 -10668 -536 -10666
rect -286 -10668 -186 -10666
rect -12400 -26481 25000 -26400
rect -12400 -26625 -7444 -26481
rect 23900 -26625 25000 -26481
rect -12400 -26854 25000 -26625
rect -12400 -27078 -12188 -26854
rect -11644 -27078 24244 -26854
rect 24788 -27078 25000 -26854
rect -12400 -27200 25000 -27078
use sky130_fd_pr__pfet_01v8_LEMKJU  sky130_fd_pr__pfet_01v8_LEMKJU_3
timestamp 1626065694
transform 1 0 4733 0 1 -7704
box -1155 -300 1155 300
use sky130_fd_pr__pfet_01v8_LEMKJU  sky130_fd_pr__pfet_01v8_LEMKJU_2
timestamp 1626065694
transform 1 0 4733 0 1 -6766
box -1155 -300 1155 300
use sky130_fd_pr__pfet_01v8_LEMKJU  sky130_fd_pr__pfet_01v8_LEMKJU_1
timestamp 1626065694
transform 1 0 4733 0 1 -5828
box -1155 -300 1155 300
use sky130_fd_pr__pfet_01v8_LEMKJU  sky130_fd_pr__pfet_01v8_LEMKJU_0
timestamp 1626065694
transform 1 0 4733 0 1 -4890
box -1155 -300 1155 300
use sky130_fd_pr__cap_mim_m3_1_KB5CJD  sky130_fd_pr__cap_mim_m3_1_KB5CJD_15
timestamp 1626065694
transform 1 0 -10133 0 1 -8921
box -1150 -1100 1149 1100
use sky130_fd_pr__cap_mim_m3_1_KB5CJD  sky130_fd_pr__cap_mim_m3_1_KB5CJD_14
timestamp 1626065694
transform 1 0 -7533 0 1 -8921
box -1150 -1100 1149 1100
use sky130_fd_pr__cap_mim_m3_1_KB5CJD  sky130_fd_pr__cap_mim_m3_1_KB5CJD_13
timestamp 1626065694
transform 1 0 -4933 0 1 -8921
box -1150 -1100 1149 1100
use sky130_fd_pr__cap_mim_m3_1_KB5CJD  sky130_fd_pr__cap_mim_m3_1_KB5CJD_12
timestamp 1626065694
transform 1 0 -2333 0 1 -8921
box -1150 -1100 1149 1100
use sky130_fd_pr__cap_mim_m3_1_KB5CJD  sky130_fd_pr__cap_mim_m3_1_KB5CJD_11
timestamp 1626065694
transform 1 0 -10133 0 1 -6421
box -1150 -1100 1149 1100
use sky130_fd_pr__cap_mim_m3_1_KB5CJD  sky130_fd_pr__cap_mim_m3_1_KB5CJD_10
timestamp 1626065694
transform 1 0 -2333 0 1 -6421
box -1150 -1100 1149 1100
use sky130_fd_pr__cap_mim_m3_1_KB5CJD  sky130_fd_pr__cap_mim_m3_1_KB5CJD_9
timestamp 1626065694
transform 1 0 -4933 0 1 -6421
box -1150 -1100 1149 1100
use sky130_fd_pr__cap_mim_m3_1_KB5CJD  sky130_fd_pr__cap_mim_m3_1_KB5CJD_8
timestamp 1626065694
transform 1 0 -7533 0 1 -6421
box -1150 -1100 1149 1100
use sky130_fd_pr__cap_mim_m3_1_KB5CJD  sky130_fd_pr__cap_mim_m3_1_KB5CJD_7
timestamp 1626065694
transform 1 0 -10133 0 1 -3921
box -1150 -1100 1149 1100
use sky130_fd_pr__cap_mim_m3_1_KB5CJD  sky130_fd_pr__cap_mim_m3_1_KB5CJD_6
timestamp 1626065694
transform 1 0 -2333 0 1 -3921
box -1150 -1100 1149 1100
use sky130_fd_pr__cap_mim_m3_1_KB5CJD  sky130_fd_pr__cap_mim_m3_1_KB5CJD_5
timestamp 1626065694
transform 1 0 -4933 0 1 -3921
box -1150 -1100 1149 1100
use sky130_fd_pr__cap_mim_m3_1_KB5CJD  sky130_fd_pr__cap_mim_m3_1_KB5CJD_4
timestamp 1626065694
transform 1 0 -7533 0 1 -3921
box -1150 -1100 1149 1100
use sky130_fd_pr__cap_mim_m3_1_KB5CJD  sky130_fd_pr__cap_mim_m3_1_KB5CJD_3
timestamp 1626065694
transform 1 0 -10133 0 1 -1420
box -1150 -1100 1149 1100
use sky130_fd_pr__cap_mim_m3_1_KB5CJD  sky130_fd_pr__cap_mim_m3_1_KB5CJD_2
timestamp 1626065694
transform 1 0 -2333 0 1 -1420
box -1150 -1100 1149 1100
use sky130_fd_pr__cap_mim_m3_1_KB5CJD  sky130_fd_pr__cap_mim_m3_1_KB5CJD_1
timestamp 1626065694
transform 1 0 -4933 0 1 -1420
box -1150 -1100 1149 1100
use sky130_fd_pr__cap_mim_m3_1_KB5CJD  sky130_fd_pr__cap_mim_m3_1_KB5CJD_0
timestamp 1626065694
transform 1 0 -7533 0 1 -1420
box -1150 -1100 1149 1100
use sky130_fd_pr__cap_mim_m3_1_P3BUE2  sky130_fd_pr__cap_mim_m3_1_P3BUE2_7
timestamp 1626065694
transform 1 0 -10134 0 1 -10619
box -1150 -300 1149 300
use sky130_fd_pr__cap_mim_m3_1_P3BUE2  sky130_fd_pr__cap_mim_m3_1_P3BUE2_6
timestamp 1626065694
transform 1 0 -7534 0 1 -10619
box -1150 -300 1149 300
use sky130_fd_pr__cap_mim_m3_1_P3BUE2  sky130_fd_pr__cap_mim_m3_1_P3BUE2_5
timestamp 1626065694
transform 1 0 -4934 0 1 -10619
box -1150 -300 1149 300
use sky130_fd_pr__cap_mim_m3_1_P3BUE2  sky130_fd_pr__cap_mim_m3_1_P3BUE2_4
timestamp 1626065694
transform 1 0 -2334 0 1 -10619
box -1150 -300 1149 300
use sky130_fd_pr__cap_mim_m3_1_P3BUE2  sky130_fd_pr__cap_mim_m3_1_P3BUE2_3
timestamp 1626065694
transform 1 0 -10134 0 1 281
box -1150 -300 1149 300
use sky130_fd_pr__cap_mim_m3_1_P3BUE2  sky130_fd_pr__cap_mim_m3_1_P3BUE2_2
timestamp 1626065694
transform 1 0 -4934 0 1 281
box -1150 -300 1149 300
use sky130_fd_pr__cap_mim_m3_1_P3BUE2  sky130_fd_pr__cap_mim_m3_1_P3BUE2_1
timestamp 1626065694
transform 1 0 -7534 0 1 281
box -1150 -300 1149 300
use sky130_fd_pr__cap_mim_m3_1_P3BUE2  sky130_fd_pr__cap_mim_m3_1_P3BUE2_0
timestamp 1626065694
transform 1 0 -2334 0 1 281
box -1150 -300 1149 300
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_3
timestamp 1626065694
transform 1 0 -11932 0 1 -10618
box -350 -300 349 300
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_2
timestamp 1626065694
transform 1 0 -534 0 1 -10618
box -350 -300 349 300
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_1
timestamp 1626065694
transform 1 0 -11928 0 1 280
box -350 -300 349 300
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_0
timestamp 1626065694
transform 1 0 -534 0 1 280
box -350 -300 349 300
use sky130_fd_pr__nfet_01v8_lvt_LYGCX9  sky130_fd_pr__nfet_01v8_lvt_LYGCX9_1
timestamp 1626065694
transform 1 0 -1217 0 1 -20554
box -1145 -188 1145 188
use sky130_fd_pr__nfet_01v8_lvt_LYGCX9  sky130_fd_pr__nfet_01v8_lvt_LYGCX9_0
timestamp 1626065694
transform 1 0 -1217 0 1 -19722
box -1145 -188 1145 188
use sky130_fd_pr__nfet_01v8_lvt_DHUKXE  sky130_fd_pr__nfet_01v8_lvt_DHUKXE_3
timestamp 1626065694
transform 1 0 -756 0 1 -25414
box -1694 -388 1694 388
use sky130_fd_pr__nfet_01v8_lvt_DHUKXE  sky130_fd_pr__nfet_01v8_lvt_DHUKXE_2
timestamp 1626065694
transform 1 0 -756 0 1 -24304
box -1694 -388 1694 388
use sky130_fd_pr__nfet_01v8_lvt_DHUKXE  sky130_fd_pr__nfet_01v8_lvt_DHUKXE_1
timestamp 1626065694
transform 1 0 -754 0 1 -23192
box -1694 -388 1694 388
use sky130_fd_pr__nfet_01v8_lvt_DHUKXE  sky130_fd_pr__nfet_01v8_lvt_DHUKXE_0
timestamp 1626065694
transform 1 0 -754 0 1 -22080
box -1694 -388 1694 388
use sky130_fd_pr__nfet_01v8_Y4K3TH  sky130_fd_pr__nfet_01v8_Y4K3TH_3
timestamp 1626065694
transform 1 0 -6335 0 1 -25418
box -3109 -388 3109 388
use sky130_fd_pr__nfet_01v8_Y4K3TH  sky130_fd_pr__nfet_01v8_Y4K3TH_2
timestamp 1626065694
transform 1 0 -6334 0 1 -24305
box -3109 -388 3109 388
use sky130_fd_pr__nfet_01v8_Y4K3TH  sky130_fd_pr__nfet_01v8_Y4K3TH_1
timestamp 1626065694
transform 1 0 -6335 0 1 -23194
box -3109 -388 3109 388
use sky130_fd_pr__nfet_01v8_Y4K3TH  sky130_fd_pr__nfet_01v8_Y4K3TH_0
timestamp 1626065694
transform 1 0 -6334 0 1 -22081
box -3109 -388 3109 388
use sky130_fd_pr__pfet_01v8_lvt_V2JKJ2  sky130_fd_pr__pfet_01v8_lvt_V2JKJ2_2
timestamp 1626065694
transform 1 0 14649 0 1 -2132
box -8209 -400 8209 400
use sky130_fd_pr__pfet_01v8_lvt_V2JKJ2  sky130_fd_pr__pfet_01v8_lvt_V2JKJ2_1
timestamp 1626065694
transform 1 0 14649 0 1 -996
box -8209 -400 8209 400
use sky130_fd_pr__pfet_01v8_lvt_V2JKJ2  sky130_fd_pr__pfet_01v8_lvt_V2JKJ2_0
timestamp 1626065694
transform 1 0 14649 0 1 140
box -8209 -400 8209 400
use sky130_fd_pr__pfet_01v8_MSJKJ2  sky130_fd_pr__pfet_01v8_MSJKJ2_3
timestamp 1626065694
transform 1 0 15126 0 1 -7674
box -7700 -400 7700 400
use sky130_fd_pr__pfet_01v8_MSJKJ2  sky130_fd_pr__pfet_01v8_MSJKJ2_2
timestamp 1626065694
transform 1 0 15126 0 1 -6418
box -7700 -400 7700 400
use sky130_fd_pr__pfet_01v8_MSJKJ2  sky130_fd_pr__pfet_01v8_MSJKJ2_1
timestamp 1626065694
transform 1 0 15126 0 1 -5162
box -7700 -400 7700 400
use sky130_fd_pr__pfet_01v8_MSJKJ2  sky130_fd_pr__pfet_01v8_MSJKJ2_0
timestamp 1626065694
transform 1 0 15126 0 1 -3906
box -7700 -400 7700 400
use sky130_fd_pr__nfet_01v8_lvt_XH9Q8F  sky130_fd_pr__nfet_01v8_lvt_XH9Q8F_1
timestamp 1626065694
transform 1 0 -4586 0 1 -17311
box -4636 -1615 4636 1615
use sky130_fd_pr__nfet_01v8_lvt_XH9Q8F  sky130_fd_pr__nfet_01v8_lvt_XH9Q8F_0
timestamp 1626065694
transform 1 0 -4586 0 1 -14039
box -4636 -1615 4636 1615
use sky130_fd_pr__nfet_01v8_MCKC3T  sky130_fd_pr__nfet_01v8_MCKC3T_11
timestamp 1626065694
transform 1 0 12777 0 1 -25584
box -10235 -388 10235 388
use sky130_fd_pr__nfet_01v8_MCKC3T  sky130_fd_pr__nfet_01v8_MCKC3T_10
timestamp 1626065694
transform 1 0 12777 0 1 -24352
box -10235 -388 10235 388
use sky130_fd_pr__nfet_01v8_MCKC3T  sky130_fd_pr__nfet_01v8_MCKC3T_9
timestamp 1626065694
transform 1 0 12777 0 1 -23118
box -10235 -388 10235 388
use sky130_fd_pr__nfet_01v8_MCKC3T  sky130_fd_pr__nfet_01v8_MCKC3T_8
timestamp 1626065694
transform 1 0 12777 0 1 -21884
box -10235 -388 10235 388
use sky130_fd_pr__nfet_01v8_MCKC3T  sky130_fd_pr__nfet_01v8_MCKC3T_7
timestamp 1626065694
transform 1 0 12777 0 1 -20652
box -10235 -388 10235 388
use sky130_fd_pr__nfet_01v8_MCKC3T  sky130_fd_pr__nfet_01v8_MCKC3T_6
timestamp 1626065694
transform 1 0 12777 0 1 -19418
box -10235 -388 10235 388
use sky130_fd_pr__nfet_01v8_MCKC3T  sky130_fd_pr__nfet_01v8_MCKC3T_5
timestamp 1626065694
transform 1 0 12777 0 1 -18184
box -10235 -388 10235 388
use sky130_fd_pr__nfet_01v8_MCKC3T  sky130_fd_pr__nfet_01v8_MCKC3T_4
timestamp 1626065694
transform 1 0 12777 0 1 -16952
box -10235 -388 10235 388
use sky130_fd_pr__nfet_01v8_MCKC3T  sky130_fd_pr__nfet_01v8_MCKC3T_3
timestamp 1626065694
transform 1 0 12777 0 1 -15718
box -10235 -388 10235 388
use sky130_fd_pr__nfet_01v8_MCKC3T  sky130_fd_pr__nfet_01v8_MCKC3T_2
timestamp 1626065694
transform 1 0 12779 0 1 -14484
box -10235 -388 10235 388
use sky130_fd_pr__nfet_01v8_MCKC3T  sky130_fd_pr__nfet_01v8_MCKC3T_1
timestamp 1626065694
transform 1 0 12779 0 1 -13252
box -10235 -388 10235 388
use sky130_fd_pr__nfet_01v8_MCKC3T  sky130_fd_pr__nfet_01v8_MCKC3T_0
timestamp 1626065694
transform 1 0 12779 0 1 -12018
box -10235 -388 10235 388
use ptap  ptap_361
timestamp 1626065694
transform 1 0 -6976 0 1 -26218
box 62 116 196 250
use ptap  ptap_360
timestamp 1626065694
transform 1 0 -9012 0 1 -26218
box 62 116 196 250
use ptap  ptap_359
timestamp 1626065694
transform 1 0 -7994 0 1 -26218
box 62 116 196 250
use ptap  ptap_358
timestamp 1626065694
transform 1 0 -384 0 1 -26272
box 62 116 196 250
use ptap  ptap_357
timestamp 1626065694
transform 1 0 -2420 0 1 -26272
box 62 116 196 250
use ptap  ptap_356
timestamp 1626065694
transform 1 0 -1402 0 1 -26272
box 62 116 196 250
use ptap  ptap_355
timestamp 1626065694
transform 1 0 -4940 0 1 -26218
box 62 116 196 250
use ptap  ptap_354
timestamp 1626065694
transform 1 0 -3922 0 1 -26218
box 62 116 196 250
use ptap  ptap_353
timestamp 1626065694
transform 1 0 -5958 0 1 -26218
box 62 116 196 250
use ptap  ptap_352
timestamp 1626065694
transform 1 0 634 0 1 -26272
box 62 116 196 250
use ptap  ptap_351
timestamp 1626065694
transform 1 0 -8986 0 1 -25024
box 62 116 196 250
use ptap  ptap_350
timestamp 1626065694
transform 1 0 -7968 0 1 -25024
box 62 116 196 250
use ptap  ptap_349
timestamp 1626065694
transform 1 0 -6950 0 1 -25024
box 62 116 196 250
use ptap  ptap_348
timestamp 1626065694
transform 1 0 -3896 0 1 -25024
box 62 116 196 250
use ptap  ptap_347
timestamp 1626065694
transform 1 0 -2394 0 1 -25038
box 62 116 196 250
use ptap  ptap_346
timestamp 1626065694
transform 1 0 -1376 0 1 -25038
box 62 116 196 250
use ptap  ptap_345
timestamp 1626065694
transform 1 0 -358 0 1 -25038
box 62 116 196 250
use ptap  ptap_344
timestamp 1626065694
transform 1 0 -5932 0 1 -25024
box 62 116 196 250
use ptap  ptap_343
timestamp 1626065694
transform 1 0 -4914 0 1 -25024
box 62 116 196 250
use ptap  ptap_342
timestamp 1626065694
transform 1 0 5014 0 1 -25132
box 62 116 196 250
use ptap  ptap_341
timestamp 1626065694
transform 1 0 3996 0 1 -25132
box 62 116 196 250
use ptap  ptap_340
timestamp 1626065694
transform 1 0 2978 0 1 -25132
box 62 116 196 250
use ptap  ptap_339
timestamp 1626065694
transform 1 0 660 0 1 -25038
box 62 116 196 250
use ptap  ptap_338
timestamp 1626065694
transform 1 0 6032 0 1 -25132
box 62 116 196 250
use ptap  ptap_337
timestamp 1626065694
transform 1 0 7050 0 1 -25132
box 62 116 196 250
use ptap  ptap_336
timestamp 1626065694
transform 1 0 8068 0 1 -25132
box 62 116 196 250
use ptap  ptap_335
timestamp 1626065694
transform 1 0 9086 0 1 -25132
box 62 116 196 250
use ptap  ptap_334
timestamp 1626065694
transform 1 0 10104 0 1 -25132
box 62 116 196 250
use ptap  ptap_333
timestamp 1626065694
transform 1 0 11122 0 1 -25132
box 62 116 196 250
use ptap  ptap_332
timestamp 1626065694
transform 1 0 12140 0 1 -25132
box 62 116 196 250
use ptap  ptap_331
timestamp 1626065694
transform 1 0 13158 0 1 -25132
box 62 116 196 250
use ptap  ptap_330
timestamp 1626065694
transform 1 0 14176 0 1 -25132
box 62 116 196 250
use ptap  ptap_329
timestamp 1626065694
transform 1 0 15194 0 1 -25132
box 62 116 196 250
use ptap  ptap_328
timestamp 1626065694
transform 1 0 16212 0 1 -25132
box 62 116 196 250
use ptap  ptap_327
timestamp 1626065694
transform 1 0 17230 0 1 -25132
box 62 116 196 250
use ptap  ptap_326
timestamp 1626065694
transform 1 0 18248 0 1 -25132
box 62 116 196 250
use ptap  ptap_325
timestamp 1626065694
transform 1 0 19266 0 1 -25132
box 62 116 196 250
use ptap  ptap_324
timestamp 1626065694
transform 1 0 20284 0 1 -25132
box 62 116 196 250
use ptap  ptap_323
timestamp 1626065694
transform 1 0 21302 0 1 -25132
box 62 116 196 250
use ptap  ptap_322
timestamp 1626065694
transform 1 0 22320 0 1 -25132
box 62 116 196 250
use ptap  ptap_321
timestamp 1626065694
transform 1 0 -9012 0 1 -23926
box 62 116 196 250
use ptap  ptap_320
timestamp 1626065694
transform 1 0 -7994 0 1 -23926
box 62 116 196 250
use ptap  ptap_319
timestamp 1626065694
transform 1 0 -6976 0 1 -23926
box 62 116 196 250
use ptap  ptap_318
timestamp 1626065694
transform 1 0 -3922 0 1 -23926
box 62 116 196 250
use ptap  ptap_317
timestamp 1626065694
transform 1 0 -2448 0 1 -23926
box 62 116 196 250
use ptap  ptap_316
timestamp 1626065694
transform 1 0 -1430 0 1 -23926
box 62 116 196 250
use ptap  ptap_315
timestamp 1626065694
transform 1 0 -412 0 1 -23926
box 62 116 196 250
use ptap  ptap_314
timestamp 1626065694
transform 1 0 -5958 0 1 -23926
box 62 116 196 250
use ptap  ptap_313
timestamp 1626065694
transform 1 0 -4940 0 1 -23926
box 62 116 196 250
use ptap  ptap_312
timestamp 1626065694
transform 1 0 3996 0 1 -23912
box 62 116 196 250
use ptap  ptap_311
timestamp 1626065694
transform 1 0 5014 0 1 -23912
box 62 116 196 250
use ptap  ptap_310
timestamp 1626065694
transform 1 0 2978 0 1 -23912
box 62 116 196 250
use ptap  ptap_309
timestamp 1626065694
transform 1 0 606 0 1 -23926
box 62 116 196 250
use ptap  ptap_308
timestamp 1626065694
transform 1 0 6032 0 1 -23912
box 62 116 196 250
use ptap  ptap_307
timestamp 1626065694
transform 1 0 7050 0 1 -23912
box 62 116 196 250
use ptap  ptap_306
timestamp 1626065694
transform 1 0 8068 0 1 -23912
box 62 116 196 250
use ptap  ptap_305
timestamp 1626065694
transform 1 0 9086 0 1 -23912
box 62 116 196 250
use ptap  ptap_304
timestamp 1626065694
transform 1 0 10104 0 1 -23912
box 62 116 196 250
use ptap  ptap_303
timestamp 1626065694
transform 1 0 11122 0 1 -23912
box 62 116 196 250
use ptap  ptap_302
timestamp 1626065694
transform 1 0 12140 0 1 -23912
box 62 116 196 250
use ptap  ptap_301
timestamp 1626065694
transform 1 0 13158 0 1 -23912
box 62 116 196 250
use ptap  ptap_300
timestamp 1626065694
transform 1 0 14176 0 1 -23912
box 62 116 196 250
use ptap  ptap_299
timestamp 1626065694
transform 1 0 15194 0 1 -23912
box 62 116 196 250
use ptap  ptap_298
timestamp 1626065694
transform 1 0 16212 0 1 -23912
box 62 116 196 250
use ptap  ptap_297
timestamp 1626065694
transform 1 0 17230 0 1 -23912
box 62 116 196 250
use ptap  ptap_296
timestamp 1626065694
transform 1 0 18248 0 1 -23912
box 62 116 196 250
use ptap  ptap_295
timestamp 1626065694
transform 1 0 19266 0 1 -23912
box 62 116 196 250
use ptap  ptap_294
timestamp 1626065694
transform 1 0 20284 0 1 -23912
box 62 116 196 250
use ptap  ptap_293
timestamp 1626065694
transform 1 0 21302 0 1 -23912
box 62 116 196 250
use ptap  ptap_292
timestamp 1626065694
transform 1 0 22320 0 1 -23912
box 62 116 196 250
use ptap  ptap_291
timestamp 1626065694
transform 1 0 -6950 0 1 -22800
box 62 116 196 250
use ptap  ptap_290
timestamp 1626065694
transform 1 0 -7968 0 1 -22800
box 62 116 196 250
use ptap  ptap_289
timestamp 1626065694
transform 1 0 -8986 0 1 -22800
box 62 116 196 250
use ptap  ptap_288
timestamp 1626065694
transform 1 0 -412 0 1 -22812
box 62 116 196 250
use ptap  ptap_287
timestamp 1626065694
transform 1 0 -1430 0 1 -22812
box 62 116 196 250
use ptap  ptap_286
timestamp 1626065694
transform 1 0 -2448 0 1 -22812
box 62 116 196 250
use ptap  ptap_285
timestamp 1626065694
transform 1 0 -3896 0 1 -22800
box 62 116 196 250
use ptap  ptap_284
timestamp 1626065694
transform 1 0 -4914 0 1 -22800
box 62 116 196 250
use ptap  ptap_283
timestamp 1626065694
transform 1 0 -5932 0 1 -22800
box 62 116 196 250
use ptap  ptap_282
timestamp 1626065694
transform 1 0 5028 0 1 -22690
box 62 116 196 250
use ptap  ptap_281
timestamp 1626065694
transform 1 0 4010 0 1 -22690
box 62 116 196 250
use ptap  ptap_280
timestamp 1626065694
transform 1 0 2992 0 1 -22690
box 62 116 196 250
use ptap  ptap_279
timestamp 1626065694
transform 1 0 606 0 1 -22812
box 62 116 196 250
use ptap  ptap_278
timestamp 1626065694
transform 1 0 6046 0 1 -22690
box 62 116 196 250
use ptap  ptap_277
timestamp 1626065694
transform 1 0 7064 0 1 -22690
box 62 116 196 250
use ptap  ptap_276
timestamp 1626065694
transform 1 0 8082 0 1 -22690
box 62 116 196 250
use ptap  ptap_275
timestamp 1626065694
transform 1 0 9100 0 1 -22690
box 62 116 196 250
use ptap  ptap_274
timestamp 1626065694
transform 1 0 10118 0 1 -22690
box 62 116 196 250
use ptap  ptap_273
timestamp 1626065694
transform 1 0 11136 0 1 -22690
box 62 116 196 250
use ptap  ptap_272
timestamp 1626065694
transform 1 0 12154 0 1 -22690
box 62 116 196 250
use ptap  ptap_271
timestamp 1626065694
transform 1 0 13172 0 1 -22690
box 62 116 196 250
use ptap  ptap_270
timestamp 1626065694
transform 1 0 14190 0 1 -22690
box 62 116 196 250
use ptap  ptap_269
timestamp 1626065694
transform 1 0 15208 0 1 -22690
box 62 116 196 250
use ptap  ptap_268
timestamp 1626065694
transform 1 0 16226 0 1 -22690
box 62 116 196 250
use ptap  ptap_267
timestamp 1626065694
transform 1 0 17244 0 1 -22690
box 62 116 196 250
use ptap  ptap_266
timestamp 1626065694
transform 1 0 18262 0 1 -22690
box 62 116 196 250
use ptap  ptap_265
timestamp 1626065694
transform 1 0 19280 0 1 -22690
box 62 116 196 250
use ptap  ptap_264
timestamp 1626065694
transform 1 0 20298 0 1 -22690
box 62 116 196 250
use ptap  ptap_263
timestamp 1626065694
transform 1 0 21316 0 1 -22690
box 62 116 196 250
use ptap  ptap_262
timestamp 1626065694
transform 1 0 22334 0 1 -22690
box 62 116 196 250
use ptap  ptap_261
timestamp 1626065694
transform 1 0 -9000 0 1 -21674
box 62 116 196 250
use ptap  ptap_260
timestamp 1626065694
transform 1 0 -6964 0 1 -21674
box 62 116 196 250
use ptap  ptap_259
timestamp 1626065694
transform 1 0 -5946 0 1 -21674
box 62 116 196 250
use ptap  ptap_258
timestamp 1626065694
transform 1 0 -7982 0 1 -21674
box 62 116 196 250
use ptap  ptap_257
timestamp 1626065694
transform 1 0 -2408 0 1 -21618
box 62 116 196 250
use ptap  ptap_256
timestamp 1626065694
transform 1 0 -4928 0 1 -21674
box 62 116 196 250
use ptap  ptap_255
timestamp 1626065694
transform 1 0 -3910 0 1 -21674
box 62 116 196 250
use ptap  ptap_254
timestamp 1626065694
transform 1 0 646 0 1 -21618
box 62 116 196 250
use ptap  ptap_253
timestamp 1626065694
transform 1 0 -1390 0 1 -21618
box 62 116 196 250
use ptap  ptap_252
timestamp 1626065694
transform 1 0 -372 0 1 -21618
box 62 116 196 250
use ptap  ptap_251
timestamp 1626065694
transform 1 0 2992 0 1 -21442
box 62 116 196 250
use ptap  ptap_250
timestamp 1626065694
transform 1 0 5028 0 1 -21442
box 62 116 196 250
use ptap  ptap_249
timestamp 1626065694
transform 1 0 4010 0 1 -21442
box 62 116 196 250
use ptap  ptap_248
timestamp 1626065694
transform 1 0 6046 0 1 -21442
box 62 116 196 250
use ptap  ptap_247
timestamp 1626065694
transform 1 0 8082 0 1 -21442
box 62 116 196 250
use ptap  ptap_246
timestamp 1626065694
transform 1 0 7064 0 1 -21442
box 62 116 196 250
use ptap  ptap_245
timestamp 1626065694
transform 1 0 10118 0 1 -21442
box 62 116 196 250
use ptap  ptap_244
timestamp 1626065694
transform 1 0 9100 0 1 -21442
box 62 116 196 250
use ptap  ptap_243
timestamp 1626065694
transform 1 0 12154 0 1 -21442
box 62 116 196 250
use ptap  ptap_242
timestamp 1626065694
transform 1 0 11136 0 1 -21442
box 62 116 196 250
use ptap  ptap_241
timestamp 1626065694
transform 1 0 13172 0 1 -21442
box 62 116 196 250
use ptap  ptap_240
timestamp 1626065694
transform 1 0 15208 0 1 -21442
box 62 116 196 250
use ptap  ptap_239
timestamp 1626065694
transform 1 0 14190 0 1 -21442
box 62 116 196 250
use ptap  ptap_238
timestamp 1626065694
transform 1 0 17244 0 1 -21442
box 62 116 196 250
use ptap  ptap_237
timestamp 1626065694
transform 1 0 16226 0 1 -21442
box 62 116 196 250
use ptap  ptap_236
timestamp 1626065694
transform 1 0 19280 0 1 -21442
box 62 116 196 250
use ptap  ptap_235
timestamp 1626065694
transform 1 0 18262 0 1 -21442
box 62 116 196 250
use ptap  ptap_234
timestamp 1626065694
transform 1 0 20298 0 1 -21442
box 62 116 196 250
use ptap  ptap_233
timestamp 1626065694
transform 1 0 22334 0 1 -21442
box 62 116 196 250
use ptap  ptap_232
timestamp 1626065694
transform 1 0 21316 0 1 -21442
box 62 116 196 250
use ptap  ptap_231
timestamp 1626065694
transform 1 0 -1688 0 1 -20330
box 62 116 196 250
use ptap  ptap_230
timestamp 1626065694
transform 1 0 -2706 0 1 -20330
box 62 116 196 250
use ptap  ptap_229
timestamp 1626065694
transform 1 0 348 0 1 -20330
box 62 116 196 250
use ptap  ptap_228
timestamp 1626065694
transform 1 0 -670 0 1 -20330
box 62 116 196 250
use ptap  ptap_227
timestamp 1626065694
transform 1 0 2978 0 1 -20222
box 62 116 196 250
use ptap  ptap_226
timestamp 1626065694
transform 1 0 5014 0 1 -20222
box 62 116 196 250
use ptap  ptap_225
timestamp 1626065694
transform 1 0 3996 0 1 -20222
box 62 116 196 250
use ptap  ptap_224
timestamp 1626065694
transform 1 0 7050 0 1 -20222
box 62 116 196 250
use ptap  ptap_223
timestamp 1626065694
transform 1 0 6032 0 1 -20222
box 62 116 196 250
use ptap  ptap_222
timestamp 1626065694
transform 1 0 9086 0 1 -20222
box 62 116 196 250
use ptap  ptap_221
timestamp 1626065694
transform 1 0 8068 0 1 -20222
box 62 116 196 250
use ptap  ptap_220
timestamp 1626065694
transform 1 0 12140 0 1 -20222
box 62 116 196 250
use ptap  ptap_219
timestamp 1626065694
transform 1 0 11122 0 1 -20222
box 62 116 196 250
use ptap  ptap_218
timestamp 1626065694
transform 1 0 10104 0 1 -20222
box 62 116 196 250
use ptap  ptap_217
timestamp 1626065694
transform 1 0 14176 0 1 -20222
box 62 116 196 250
use ptap  ptap_216
timestamp 1626065694
transform 1 0 13158 0 1 -20222
box 62 116 196 250
use ptap  ptap_215
timestamp 1626065694
transform 1 0 16212 0 1 -20222
box 62 116 196 250
use ptap  ptap_214
timestamp 1626065694
transform 1 0 15194 0 1 -20222
box 62 116 196 250
use ptap  ptap_213
timestamp 1626065694
transform 1 0 18248 0 1 -20222
box 62 116 196 250
use ptap  ptap_212
timestamp 1626065694
transform 1 0 17230 0 1 -20222
box 62 116 196 250
use ptap  ptap_211
timestamp 1626065694
transform 1 0 20284 0 1 -20222
box 62 116 196 250
use ptap  ptap_210
timestamp 1626065694
transform 1 0 19266 0 1 -20222
box 62 116 196 250
use ptap  ptap_209
timestamp 1626065694
transform 1 0 22320 0 1 -20222
box 62 116 196 250
use ptap  ptap_208
timestamp 1626065694
transform 1 0 21302 0 1 -20222
box 62 116 196 250
use ptap  ptap_207
timestamp 1626065694
transform 1 0 -8784 0 1 -19354
box 62 116 196 250
use ptap  ptap_206
timestamp 1626065694
transform 1 0 -7766 0 1 -19354
box 62 116 196 250
use ptap  ptap_205
timestamp 1626065694
transform 1 0 -6748 0 1 -19354
box 62 116 196 250
use ptap  ptap_204
timestamp 1626065694
transform 1 0 -5730 0 1 -19354
box 62 116 196 250
use ptap  ptap_203
timestamp 1626065694
transform 1 0 -4712 0 1 -19354
box 62 116 196 250
use ptap  ptap_202
timestamp 1626065694
transform 1 0 -3694 0 1 -19354
box 62 116 196 250
use ptap  ptap_201
timestamp 1626065694
transform 1 0 -2676 0 1 -19354
box 62 116 196 250
use ptap  ptap_200
timestamp 1626065694
transform 1 0 -1658 0 1 -19354
box 62 116 196 250
use ptap  ptap_199
timestamp 1626065694
transform 1 0 -640 0 1 -19354
box 62 116 196 250
use ptap  ptap_198
timestamp 1626065694
transform 1 0 2978 0 1 -18974
box 62 116 196 250
use ptap  ptap_197
timestamp 1626065694
transform 1 0 3996 0 1 -18974
box 62 116 196 250
use ptap  ptap_196
timestamp 1626065694
transform 1 0 5014 0 1 -18974
box 62 116 196 250
use ptap  ptap_195
timestamp 1626065694
transform 1 0 6032 0 1 -18974
box 62 116 196 250
use ptap  ptap_194
timestamp 1626065694
transform 1 0 7050 0 1 -18974
box 62 116 196 250
use ptap  ptap_193
timestamp 1626065694
transform 1 0 8068 0 1 -18974
box 62 116 196 250
use ptap  ptap_192
timestamp 1626065694
transform 1 0 9086 0 1 -18974
box 62 116 196 250
use ptap  ptap_191
timestamp 1626065694
transform 1 0 10104 0 1 -18974
box 62 116 196 250
use ptap  ptap_190
timestamp 1626065694
transform 1 0 11122 0 1 -18974
box 62 116 196 250
use ptap  ptap_189
timestamp 1626065694
transform 1 0 12140 0 1 -18974
box 62 116 196 250
use ptap  ptap_188
timestamp 1626065694
transform 1 0 13158 0 1 -18974
box 62 116 196 250
use ptap  ptap_187
timestamp 1626065694
transform 1 0 15194 0 1 -18974
box 62 116 196 250
use ptap  ptap_186
timestamp 1626065694
transform 1 0 14176 0 1 -18974
box 62 116 196 250
use ptap  ptap_185
timestamp 1626065694
transform 1 0 17230 0 1 -18974
box 62 116 196 250
use ptap  ptap_184
timestamp 1626065694
transform 1 0 16212 0 1 -18974
box 62 116 196 250
use ptap  ptap_183
timestamp 1626065694
transform 1 0 19266 0 1 -18974
box 62 116 196 250
use ptap  ptap_182
timestamp 1626065694
transform 1 0 18248 0 1 -18974
box 62 116 196 250
use ptap  ptap_181
timestamp 1626065694
transform 1 0 20284 0 1 -18974
box 62 116 196 250
use ptap  ptap_180
timestamp 1626065694
transform 1 0 22320 0 1 -18974
box 62 116 196 250
use ptap  ptap_179
timestamp 1626065694
transform 1 0 21302 0 1 -18974
box 62 116 196 250
use ptap  ptap_178
timestamp 1626065694
transform 1 0 -9294 0 1 -18312
box 62 116 196 250
use ptap  ptap_177
timestamp 1626065694
transform 1 0 -6240 0 1 -18312
box 62 116 196 250
use ptap  ptap_176
timestamp 1626065694
transform 1 0 -7258 0 1 -18312
box 62 116 196 250
use ptap  ptap_175
timestamp 1626065694
transform 1 0 -8276 0 1 -18312
box 62 116 196 250
use ptap  ptap_174
timestamp 1626065694
transform 1 0 -2168 0 1 -18312
box 62 116 196 250
use ptap  ptap_173
timestamp 1626065694
transform 1 0 -3186 0 1 -18312
box 62 116 196 250
use ptap  ptap_172
timestamp 1626065694
transform 1 0 -4204 0 1 -18312
box 62 116 196 250
use ptap  ptap_171
timestamp 1626065694
transform 1 0 -5222 0 1 -18312
box 62 116 196 250
use ptap  ptap_170
timestamp 1626065694
transform 1 0 -132 0 1 -18312
box 62 116 196 250
use ptap  ptap_169
timestamp 1626065694
transform 1 0 -1150 0 1 -18312
box 62 116 196 250
use ptap  ptap_168
timestamp 1626065694
transform 1 0 -9294 0 1 -17494
box 62 116 196 250
use ptap  ptap_167
timestamp 1626065694
transform 1 0 -8276 0 1 -17494
box 62 116 196 250
use ptap  ptap_166
timestamp 1626065694
transform 1 0 -7258 0 1 -17494
box 62 116 196 250
use ptap  ptap_165
timestamp 1626065694
transform 1 0 -6240 0 1 -17494
box 62 116 196 250
use ptap  ptap_164
timestamp 1626065694
transform 1 0 -4204 0 1 -17494
box 62 116 196 250
use ptap  ptap_163
timestamp 1626065694
transform 1 0 -5222 0 1 -17494
box 62 116 196 250
use ptap  ptap_162
timestamp 1626065694
transform 1 0 -3186 0 1 -17494
box 62 116 196 250
use ptap  ptap_161
timestamp 1626065694
transform 1 0 -2168 0 1 -17494
box 62 116 196 250
use ptap  ptap_160
timestamp 1626065694
transform 1 0 -1150 0 1 -17494
box 62 116 196 250
use ptap  ptap_159
timestamp 1626065694
transform 1 0 -132 0 1 -17494
box 62 116 196 250
use ptap  ptap_158
timestamp 1626065694
transform 1 0 4010 0 1 -17752
box 62 116 196 250
use ptap  ptap_157
timestamp 1626065694
transform 1 0 2992 0 1 -17752
box 62 116 196 250
use ptap  ptap_156
timestamp 1626065694
transform 1 0 5028 0 1 -17752
box 62 116 196 250
use ptap  ptap_155
timestamp 1626065694
transform 1 0 6046 0 1 -17752
box 62 116 196 250
use ptap  ptap_154
timestamp 1626065694
transform 1 0 7064 0 1 -17752
box 62 116 196 250
use ptap  ptap_153
timestamp 1626065694
transform 1 0 8082 0 1 -17752
box 62 116 196 250
use ptap  ptap_152
timestamp 1626065694
transform 1 0 9100 0 1 -17752
box 62 116 196 250
use ptap  ptap_151
timestamp 1626065694
transform 1 0 11136 0 1 -17752
box 62 116 196 250
use ptap  ptap_150
timestamp 1626065694
transform 1 0 10118 0 1 -17752
box 62 116 196 250
use ptap  ptap_149
timestamp 1626065694
transform 1 0 12154 0 1 -17752
box 62 116 196 250
use ptap  ptap_148
timestamp 1626065694
transform 1 0 13172 0 1 -17752
box 62 116 196 250
use ptap  ptap_147
timestamp 1626065694
transform 1 0 14190 0 1 -17752
box 62 116 196 250
use ptap  ptap_146
timestamp 1626065694
transform 1 0 15208 0 1 -17752
box 62 116 196 250
use ptap  ptap_145
timestamp 1626065694
transform 1 0 16226 0 1 -17752
box 62 116 196 250
use ptap  ptap_144
timestamp 1626065694
transform 1 0 17244 0 1 -17752
box 62 116 196 250
use ptap  ptap_143
timestamp 1626065694
transform 1 0 19280 0 1 -17752
box 62 116 196 250
use ptap  ptap_142
timestamp 1626065694
transform 1 0 18262 0 1 -17752
box 62 116 196 250
use ptap  ptap_141
timestamp 1626065694
transform 1 0 20298 0 1 -17752
box 62 116 196 250
use ptap  ptap_140
timestamp 1626065694
transform 1 0 21316 0 1 -17752
box 62 116 196 250
use ptap  ptap_139
timestamp 1626065694
transform 1 0 22334 0 1 -17752
box 62 116 196 250
use ptap  ptap_138
timestamp 1626065694
transform 1 0 -9294 0 1 -16676
box 62 116 196 250
use ptap  ptap_137
timestamp 1626065694
transform 1 0 -6240 0 1 -16676
box 62 116 196 250
use ptap  ptap_136
timestamp 1626065694
transform 1 0 -7258 0 1 -16676
box 62 116 196 250
use ptap  ptap_135
timestamp 1626065694
transform 1 0 -8276 0 1 -16676
box 62 116 196 250
use ptap  ptap_134
timestamp 1626065694
transform 1 0 -2168 0 1 -16676
box 62 116 196 250
use ptap  ptap_133
timestamp 1626065694
transform 1 0 -3186 0 1 -16676
box 62 116 196 250
use ptap  ptap_132
timestamp 1626065694
transform 1 0 -4204 0 1 -16676
box 62 116 196 250
use ptap  ptap_131
timestamp 1626065694
transform 1 0 -5222 0 1 -16676
box 62 116 196 250
use ptap  ptap_130
timestamp 1626065694
transform 1 0 -132 0 1 -16676
box 62 116 196 250
use ptap  ptap_129
timestamp 1626065694
transform 1 0 -1150 0 1 -16676
box 62 116 196 250
use ptap  ptap_128
timestamp 1626065694
transform 1 0 2978 0 1 -16504
box 62 116 196 250
use ptap  ptap_127
timestamp 1626065694
transform 1 0 5014 0 1 -16504
box 62 116 196 250
use ptap  ptap_126
timestamp 1626065694
transform 1 0 3996 0 1 -16504
box 62 116 196 250
use ptap  ptap_125
timestamp 1626065694
transform 1 0 6032 0 1 -16504
box 62 116 196 250
use ptap  ptap_124
timestamp 1626065694
transform 1 0 8068 0 1 -16504
box 62 116 196 250
use ptap  ptap_123
timestamp 1626065694
transform 1 0 7050 0 1 -16504
box 62 116 196 250
use ptap  ptap_122
timestamp 1626065694
transform 1 0 10104 0 1 -16504
box 62 116 196 250
use ptap  ptap_121
timestamp 1626065694
transform 1 0 9086 0 1 -16504
box 62 116 196 250
use ptap  ptap_120
timestamp 1626065694
transform 1 0 12140 0 1 -16504
box 62 116 196 250
use ptap  ptap_119
timestamp 1626065694
transform 1 0 11122 0 1 -16504
box 62 116 196 250
use ptap  ptap_118
timestamp 1626065694
transform 1 0 13158 0 1 -16504
box 62 116 196 250
use ptap  ptap_117
timestamp 1626065694
transform 1 0 15194 0 1 -16504
box 62 116 196 250
use ptap  ptap_116
timestamp 1626065694
transform 1 0 14176 0 1 -16504
box 62 116 196 250
use ptap  ptap_115
timestamp 1626065694
transform 1 0 17230 0 1 -16504
box 62 116 196 250
use ptap  ptap_114
timestamp 1626065694
transform 1 0 16212 0 1 -16504
box 62 116 196 250
use ptap  ptap_113
timestamp 1626065694
transform 1 0 19266 0 1 -16504
box 62 116 196 250
use ptap  ptap_112
timestamp 1626065694
transform 1 0 18248 0 1 -16504
box 62 116 196 250
use ptap  ptap_111
timestamp 1626065694
transform 1 0 20284 0 1 -16504
box 62 116 196 250
use ptap  ptap_110
timestamp 1626065694
transform 1 0 22320 0 1 -16504
box 62 116 196 250
use ptap  ptap_109
timestamp 1626065694
transform 1 0 21302 0 1 -16504
box 62 116 196 250
use ptap  ptap_108
timestamp 1626065694
transform 1 0 -9294 0 1 -15858
box 62 116 196 250
use ptap  ptap_107
timestamp 1626065694
transform 1 0 -6240 0 1 -15858
box 62 116 196 250
use ptap  ptap_106
timestamp 1626065694
transform 1 0 -7258 0 1 -15858
box 62 116 196 250
use ptap  ptap_105
timestamp 1626065694
transform 1 0 -8276 0 1 -15858
box 62 116 196 250
use ptap  ptap_104
timestamp 1626065694
transform 1 0 -2168 0 1 -15858
box 62 116 196 250
use ptap  ptap_103
timestamp 1626065694
transform 1 0 -3186 0 1 -15858
box 62 116 196 250
use ptap  ptap_102
timestamp 1626065694
transform 1 0 -4204 0 1 -15858
box 62 116 196 250
use ptap  ptap_101
timestamp 1626065694
transform 1 0 -5222 0 1 -15858
box 62 116 196 250
use ptap  ptap_100
timestamp 1626065694
transform 1 0 -132 0 1 -15858
box 62 116 196 250
use ptap  ptap_99
timestamp 1626065694
transform 1 0 -1150 0 1 -15858
box 62 116 196 250
use ptap  ptap_98
timestamp 1626065694
transform 1 0 -9294 0 1 -15040
box 62 116 196 250
use ptap  ptap_97
timestamp 1626065694
transform 1 0 -8276 0 1 -15040
box 62 116 196 250
use ptap  ptap_96
timestamp 1626065694
transform 1 0 -7258 0 1 -15040
box 62 116 196 250
use ptap  ptap_95
timestamp 1626065694
transform 1 0 -6240 0 1 -15040
box 62 116 196 250
use ptap  ptap_94
timestamp 1626065694
transform 1 0 -4204 0 1 -15040
box 62 116 196 250
use ptap  ptap_93
timestamp 1626065694
transform 1 0 -5222 0 1 -15040
box 62 116 196 250
use ptap  ptap_92
timestamp 1626065694
transform 1 0 -3186 0 1 -15040
box 62 116 196 250
use ptap  ptap_91
timestamp 1626065694
transform 1 0 -2168 0 1 -15040
box 62 116 196 250
use ptap  ptap_90
timestamp 1626065694
transform 1 0 -1150 0 1 -15040
box 62 116 196 250
use ptap  ptap_89
timestamp 1626065694
transform 1 0 -132 0 1 -15040
box 62 116 196 250
use ptap  ptap_88
timestamp 1626065694
transform 1 0 3996 0 1 -15284
box 62 116 196 250
use ptap  ptap_87
timestamp 1626065694
transform 1 0 2978 0 1 -15284
box 62 116 196 250
use ptap  ptap_86
timestamp 1626065694
transform 1 0 5014 0 1 -15284
box 62 116 196 250
use ptap  ptap_85
timestamp 1626065694
transform 1 0 6032 0 1 -15284
box 62 116 196 250
use ptap  ptap_84
timestamp 1626065694
transform 1 0 7050 0 1 -15284
box 62 116 196 250
use ptap  ptap_83
timestamp 1626065694
transform 1 0 8068 0 1 -15284
box 62 116 196 250
use ptap  ptap_82
timestamp 1626065694
transform 1 0 9086 0 1 -15284
box 62 116 196 250
use ptap  ptap_81
timestamp 1626065694
transform 1 0 11122 0 1 -15284
box 62 116 196 250
use ptap  ptap_80
timestamp 1626065694
transform 1 0 10104 0 1 -15284
box 62 116 196 250
use ptap  ptap_79
timestamp 1626065694
transform 1 0 12140 0 1 -15284
box 62 116 196 250
use ptap  ptap_78
timestamp 1626065694
transform 1 0 13158 0 1 -15284
box 62 116 196 250
use ptap  ptap_77
timestamp 1626065694
transform 1 0 14176 0 1 -15284
box 62 116 196 250
use ptap  ptap_76
timestamp 1626065694
transform 1 0 15194 0 1 -15284
box 62 116 196 250
use ptap  ptap_75
timestamp 1626065694
transform 1 0 16212 0 1 -15284
box 62 116 196 250
use ptap  ptap_74
timestamp 1626065694
transform 1 0 17230 0 1 -15284
box 62 116 196 250
use ptap  ptap_73
timestamp 1626065694
transform 1 0 19266 0 1 -15284
box 62 116 196 250
use ptap  ptap_72
timestamp 1626065694
transform 1 0 18248 0 1 -15284
box 62 116 196 250
use ptap  ptap_71
timestamp 1626065694
transform 1 0 20284 0 1 -15284
box 62 116 196 250
use ptap  ptap_70
timestamp 1626065694
transform 1 0 21302 0 1 -15284
box 62 116 196 250
use ptap  ptap_69
timestamp 1626065694
transform 1 0 22320 0 1 -15284
box 62 116 196 250
use ptap  ptap_68
timestamp 1626065694
transform 1 0 -9294 0 1 -14222
box 62 116 196 250
use ptap  ptap_67
timestamp 1626065694
transform 1 0 -6240 0 1 -14222
box 62 116 196 250
use ptap  ptap_66
timestamp 1626065694
transform 1 0 -7258 0 1 -14222
box 62 116 196 250
use ptap  ptap_65
timestamp 1626065694
transform 1 0 -8276 0 1 -14222
box 62 116 196 250
use ptap  ptap_64
timestamp 1626065694
transform 1 0 -2168 0 1 -14222
box 62 116 196 250
use ptap  ptap_63
timestamp 1626065694
transform 1 0 -3186 0 1 -14222
box 62 116 196 250
use ptap  ptap_62
timestamp 1626065694
transform 1 0 -4204 0 1 -14222
box 62 116 196 250
use ptap  ptap_61
timestamp 1626065694
transform 1 0 -5222 0 1 -14222
box 62 116 196 250
use ptap  ptap_60
timestamp 1626065694
transform 1 0 -132 0 1 -14222
box 62 116 196 250
use ptap  ptap_59
timestamp 1626065694
transform 1 0 -1150 0 1 -14222
box 62 116 196 250
use ptap  ptap_58
timestamp 1626065694
transform 1 0 2966 0 1 -14050
box 62 116 196 250
use ptap  ptap_57
timestamp 1626065694
transform 1 0 5002 0 1 -14050
box 62 116 196 250
use ptap  ptap_56
timestamp 1626065694
transform 1 0 3984 0 1 -14050
box 62 116 196 250
use ptap  ptap_55
timestamp 1626065694
transform 1 0 7038 0 1 -14050
box 62 116 196 250
use ptap  ptap_54
timestamp 1626065694
transform 1 0 6020 0 1 -14050
box 62 116 196 250
use ptap  ptap_53
timestamp 1626065694
transform 1 0 8056 0 1 -14050
box 62 116 196 250
use ptap  ptap_52
timestamp 1626065694
transform 1 0 10092 0 1 -14050
box 62 116 196 250
use ptap  ptap_51
timestamp 1626065694
transform 1 0 9074 0 1 -14050
box 62 116 196 250
use ptap  ptap_50
timestamp 1626065694
transform 1 0 12128 0 1 -14050
box 62 116 196 250
use ptap  ptap_49
timestamp 1626065694
transform 1 0 11110 0 1 -14050
box 62 116 196 250
use ptap  ptap_48
timestamp 1626065694
transform 1 0 13146 0 1 -14050
box 62 116 196 250
use ptap  ptap_47
timestamp 1626065694
transform 1 0 15182 0 1 -14050
box 62 116 196 250
use ptap  ptap_46
timestamp 1626065694
transform 1 0 14164 0 1 -14050
box 62 116 196 250
use ptap  ptap_45
timestamp 1626065694
transform 1 0 17218 0 1 -14050
box 62 116 196 250
use ptap  ptap_44
timestamp 1626065694
transform 1 0 16200 0 1 -14050
box 62 116 196 250
use ptap  ptap_43
timestamp 1626065694
transform 1 0 19254 0 1 -14050
box 62 116 196 250
use ptap  ptap_42
timestamp 1626065694
transform 1 0 18236 0 1 -14050
box 62 116 196 250
use ptap  ptap_41
timestamp 1626065694
transform 1 0 20272 0 1 -14050
box 62 116 196 250
use ptap  ptap_40
timestamp 1626065694
transform 1 0 22308 0 1 -14050
box 62 116 196 250
use ptap  ptap_39
timestamp 1626065694
transform 1 0 21290 0 1 -14050
box 62 116 196 250
use ptap  ptap_38
timestamp 1626065694
transform 1 0 -9294 0 1 -13404
box 62 116 196 250
use ptap  ptap_37
timestamp 1626065694
transform 1 0 -7258 0 1 -13404
box 62 116 196 250
use ptap  ptap_36
timestamp 1626065694
transform 1 0 -6240 0 1 -13404
box 62 116 196 250
use ptap  ptap_35
timestamp 1626065694
transform 1 0 -8276 0 1 -13404
box 62 116 196 250
use ptap  ptap_34
timestamp 1626065694
transform 1 0 -3186 0 1 -13404
box 62 116 196 250
use ptap  ptap_33
timestamp 1626065694
transform 1 0 -2168 0 1 -13404
box 62 116 196 250
use ptap  ptap_32
timestamp 1626065694
transform 1 0 -5222 0 1 -13404
box 62 116 196 250
use ptap  ptap_31
timestamp 1626065694
transform 1 0 -4204 0 1 -13404
box 62 116 196 250
use ptap  ptap_30
timestamp 1626065694
transform 1 0 -1150 0 1 -13404
box 62 116 196 250
use ptap  ptap_29
timestamp 1626065694
transform 1 0 -132 0 1 -13404
box 62 116 196 250
use ptap  ptap_28
timestamp 1626065694
transform 1 0 -8756 0 1 -12422
box 62 116 196 250
use ptap  ptap_27
timestamp 1626065694
transform 1 0 -7738 0 1 -12422
box 62 116 196 250
use ptap  ptap_26
timestamp 1626065694
transform 1 0 -6720 0 1 -12422
box 62 116 196 250
use ptap  ptap_25
timestamp 1626065694
transform 1 0 -5702 0 1 -12422
box 62 116 196 250
use ptap  ptap_24
timestamp 1626065694
transform 1 0 -4684 0 1 -12422
box 62 116 196 250
use ptap  ptap_23
timestamp 1626065694
transform 1 0 -3666 0 1 -12422
box 62 116 196 250
use ptap  ptap_22
timestamp 1626065694
transform 1 0 -2648 0 1 -12422
box 62 116 196 250
use ptap  ptap_21
timestamp 1626065694
transform 1 0 -1630 0 1 -12422
box 62 116 196 250
use ptap  ptap_20
timestamp 1626065694
transform 1 0 -612 0 1 -12422
box 62 116 196 250
use ptap  ptap_19
timestamp 1626065694
transform 1 0 2978 0 1 -12814
box 62 116 196 250
use ptap  ptap_18
timestamp 1626065694
transform 1 0 3996 0 1 -12814
box 62 116 196 250
use ptap  ptap_17
timestamp 1626065694
transform 1 0 5014 0 1 -12814
box 62 116 196 250
use ptap  ptap_16
timestamp 1626065694
transform 1 0 6032 0 1 -12814
box 62 116 196 250
use ptap  ptap_15
timestamp 1626065694
transform 1 0 7050 0 1 -12814
box 62 116 196 250
use ptap  ptap_14
timestamp 1626065694
transform 1 0 8068 0 1 -12814
box 62 116 196 250
use ptap  ptap_13
timestamp 1626065694
transform 1 0 9086 0 1 -12814
box 62 116 196 250
use ptap  ptap_12
timestamp 1626065694
transform 1 0 10104 0 1 -12814
box 62 116 196 250
use ptap  ptap_11
timestamp 1626065694
transform 1 0 11122 0 1 -12814
box 62 116 196 250
use ptap  ptap_10
timestamp 1626065694
transform 1 0 12140 0 1 -12814
box 62 116 196 250
use ptap  ptap_9
timestamp 1626065694
transform 1 0 13158 0 1 -12814
box 62 116 196 250
use ptap  ptap_8
timestamp 1626065694
transform 1 0 14176 0 1 -12814
box 62 116 196 250
use ptap  ptap_7
timestamp 1626065694
transform 1 0 15194 0 1 -12814
box 62 116 196 250
use ptap  ptap_6
timestamp 1626065694
transform 1 0 16212 0 1 -12814
box 62 116 196 250
use ptap  ptap_5
timestamp 1626065694
transform 1 0 17230 0 1 -12814
box 62 116 196 250
use ptap  ptap_4
timestamp 1626065694
transform 1 0 18248 0 1 -12814
box 62 116 196 250
use ptap  ptap_3
timestamp 1626065694
transform 1 0 19266 0 1 -12814
box 62 116 196 250
use ptap  ptap_2
timestamp 1626065694
transform 1 0 20284 0 1 -12814
box 62 116 196 250
use ptap  ptap_1
timestamp 1626065694
transform 1 0 21302 0 1 -12814
box 62 116 196 250
use ptap  ptap_0
timestamp 1626065694
transform 1 0 22320 0 1 -12814
box 62 116 196 250
use ntap  ntap_102
timestamp 1626065694
transform 1 0 3326 0 1 -7550
box 250 218 480 436
use ntap  ntap_101
timestamp 1626065694
transform 1 0 4344 0 1 -7550
box 250 218 480 436
use ntap  ntap_100
timestamp 1626065694
transform 1 0 5362 0 1 -7550
box 250 218 480 436
use ntap  ntap_99
timestamp 1626065694
transform 1 0 7628 0 1 -7356
box 250 218 480 436
use ntap  ntap_98
timestamp 1626065694
transform 1 0 8646 0 1 -7356
box 250 218 480 436
use ntap  ntap_97
timestamp 1626065694
transform 1 0 9664 0 1 -7356
box 250 218 480 436
use ntap  ntap_96
timestamp 1626065694
transform 1 0 11700 0 1 -7356
box 250 218 480 436
use ntap  ntap_95
timestamp 1626065694
transform 1 0 10682 0 1 -7356
box 250 218 480 436
use ntap  ntap_94
timestamp 1626065694
transform 1 0 12718 0 1 -7356
box 250 218 480 436
use ntap  ntap_93
timestamp 1626065694
transform 1 0 13736 0 1 -7356
box 250 218 480 436
use ntap  ntap_92
timestamp 1626065694
transform 1 0 15772 0 1 -7356
box 250 218 480 436
use ntap  ntap_91
timestamp 1626065694
transform 1 0 14754 0 1 -7356
box 250 218 480 436
use ntap  ntap_90
timestamp 1626065694
transform 1 0 16790 0 1 -7356
box 250 218 480 436
use ntap  ntap_89
timestamp 1626065694
transform 1 0 17808 0 1 -7356
box 250 218 480 436
use ntap  ntap_88
timestamp 1626065694
transform 1 0 19844 0 1 -7356
box 250 218 480 436
use ntap  ntap_87
timestamp 1626065694
transform 1 0 18826 0 1 -7356
box 250 218 480 436
use ntap  ntap_86
timestamp 1626065694
transform 1 0 20862 0 1 -7356
box 250 218 480 436
use ntap  ntap_85
timestamp 1626065694
transform 1 0 21880 0 1 -7356
box 250 218 480 436
use ntap  ntap_84
timestamp 1626065694
transform 1 0 4344 0 1 -6636
box 250 218 480 436
use ntap  ntap_83
timestamp 1626065694
transform 1 0 3326 0 1 -6636
box 250 218 480 436
use ntap  ntap_82
timestamp 1626065694
transform 1 0 5362 0 1 -6636
box 250 218 480 436
use ntap  ntap_81
timestamp 1626065694
transform 1 0 9664 0 1 -6118
box 250 218 480 436
use ntap  ntap_80
timestamp 1626065694
transform 1 0 8646 0 1 -6118
box 250 218 480 436
use ntap  ntap_79
timestamp 1626065694
transform 1 0 7628 0 1 -6118
box 250 218 480 436
use ntap  ntap_78
timestamp 1626065694
transform 1 0 3354 0 1 -5694
box 250 218 480 436
use ntap  ntap_77
timestamp 1626065694
transform 1 0 4372 0 1 -5694
box 250 218 480 436
use ntap  ntap_76
timestamp 1626065694
transform 1 0 5390 0 1 -5694
box 250 218 480 436
use ntap  ntap_75
timestamp 1626065694
transform 1 0 10682 0 1 -6118
box 250 218 480 436
use ntap  ntap_74
timestamp 1626065694
transform 1 0 11700 0 1 -6118
box 250 218 480 436
use ntap  ntap_73
timestamp 1626065694
transform 1 0 12718 0 1 -6118
box 250 218 480 436
use ntap  ntap_72
timestamp 1626065694
transform 1 0 13736 0 1 -6118
box 250 218 480 436
use ntap  ntap_71
timestamp 1626065694
transform 1 0 14754 0 1 -6118
box 250 218 480 436
use ntap  ntap_70
timestamp 1626065694
transform 1 0 15772 0 1 -6118
box 250 218 480 436
use ntap  ntap_69
timestamp 1626065694
transform 1 0 16790 0 1 -6118
box 250 218 480 436
use ntap  ntap_68
timestamp 1626065694
transform 1 0 17808 0 1 -6118
box 250 218 480 436
use ntap  ntap_67
timestamp 1626065694
transform 1 0 3396 0 1 -4610
box 250 218 480 436
use ntap  ntap_66
timestamp 1626065694
transform 1 0 4414 0 1 -4610
box 250 218 480 436
use ntap  ntap_65
timestamp 1626065694
transform 1 0 5432 0 1 -4610
box 250 218 480 436
use ntap  ntap_64
timestamp 1626065694
transform 1 0 7670 0 1 -4850
box 250 218 480 436
use ntap  ntap_63
timestamp 1626065694
transform 1 0 8688 0 1 -4850
box 250 218 480 436
use ntap  ntap_62
timestamp 1626065694
transform 1 0 9706 0 1 -4850
box 250 218 480 436
use ntap  ntap_61
timestamp 1626065694
transform 1 0 10724 0 1 -4850
box 250 218 480 436
use ntap  ntap_60
timestamp 1626065694
transform 1 0 11742 0 1 -4850
box 250 218 480 436
use ntap  ntap_59
timestamp 1626065694
transform 1 0 12760 0 1 -4850
box 250 218 480 436
use ntap  ntap_58
timestamp 1626065694
transform 1 0 13778 0 1 -4850
box 250 218 480 436
use ntap  ntap_57
timestamp 1626065694
transform 1 0 14796 0 1 -4850
box 250 218 480 436
use ntap  ntap_56
timestamp 1626065694
transform 1 0 15814 0 1 -4850
box 250 218 480 436
use ntap  ntap_55
timestamp 1626065694
transform 1 0 16832 0 1 -4850
box 250 218 480 436
use ntap  ntap_54
timestamp 1626065694
transform 1 0 17850 0 1 -4850
box 250 218 480 436
use ntap  ntap_53
timestamp 1626065694
transform 1 0 19844 0 1 -6118
box 250 218 480 436
use ntap  ntap_52
timestamp 1626065694
transform 1 0 18826 0 1 -6118
box 250 218 480 436
use ntap  ntap_51
timestamp 1626065694
transform 1 0 20862 0 1 -6118
box 250 218 480 436
use ntap  ntap_50
timestamp 1626065694
transform 1 0 21880 0 1 -6118
box 250 218 480 436
use ntap  ntap_49
timestamp 1626065694
transform 1 0 19886 0 1 -4850
box 250 218 480 436
use ntap  ntap_48
timestamp 1626065694
transform 1 0 18868 0 1 -4850
box 250 218 480 436
use ntap  ntap_47
timestamp 1626065694
transform 1 0 20904 0 1 -4850
box 250 218 480 436
use ntap  ntap_46
timestamp 1626065694
transform 1 0 21922 0 1 -4850
box 250 218 480 436
use ntap  ntap_45
timestamp 1626065694
transform 1 0 7670 0 1 -3338
box 250 218 480 436
use ntap  ntap_44
timestamp 1626065694
transform 1 0 8688 0 1 -3338
box 250 218 480 436
use ntap  ntap_43
timestamp 1626065694
transform 1 0 9706 0 1 -3338
box 250 218 480 436
use ntap  ntap_42
timestamp 1626065694
transform 1 0 10724 0 1 -3338
box 250 218 480 436
use ntap  ntap_41
timestamp 1626065694
transform 1 0 11742 0 1 -3338
box 250 218 480 436
use ntap  ntap_40
timestamp 1626065694
transform 1 0 12760 0 1 -3338
box 250 218 480 436
use ntap  ntap_39
timestamp 1626065694
transform 1 0 13778 0 1 -3338
box 250 218 480 436
use ntap  ntap_38
timestamp 1626065694
transform 1 0 14796 0 1 -3338
box 250 218 480 436
use ntap  ntap_37
timestamp 1626065694
transform 1 0 15814 0 1 -3338
box 250 218 480 436
use ntap  ntap_36
timestamp 1626065694
transform 1 0 16832 0 1 -3338
box 250 218 480 436
use ntap  ntap_35
timestamp 1626065694
transform 1 0 17850 0 1 -3338
box 250 218 480 436
use ntap  ntap_34
timestamp 1626065694
transform 1 0 18868 0 1 -3338
box 250 218 480 436
use ntap  ntap_33
timestamp 1626065694
transform 1 0 19886 0 1 -3338
box 250 218 480 436
use ntap  ntap_32
timestamp 1626065694
transform 1 0 6652 0 1 -1894
box 250 218 480 436
use ntap  ntap_31
timestamp 1626065694
transform 1 0 7670 0 1 -1894
box 250 218 480 436
use ntap  ntap_30
timestamp 1626065694
transform 1 0 9706 0 1 -1894
box 250 218 480 436
use ntap  ntap_29
timestamp 1626065694
transform 1 0 8688 0 1 -1894
box 250 218 480 436
use ntap  ntap_28
timestamp 1626065694
transform 1 0 10724 0 1 -1894
box 250 218 480 436
use ntap  ntap_27
timestamp 1626065694
transform 1 0 11742 0 1 -1894
box 250 218 480 436
use ntap  ntap_26
timestamp 1626065694
transform 1 0 12760 0 1 -1894
box 250 218 480 436
use ntap  ntap_25
timestamp 1626065694
transform 1 0 13778 0 1 -1894
box 250 218 480 436
use ntap  ntap_24
timestamp 1626065694
transform 1 0 14796 0 1 -1894
box 250 218 480 436
use ntap  ntap_23
timestamp 1626065694
transform 1 0 15814 0 1 -1894
box 250 218 480 436
use ntap  ntap_22
timestamp 1626065694
transform 1 0 16832 0 1 -1894
box 250 218 480 436
use ntap  ntap_21
timestamp 1626065694
transform 1 0 17850 0 1 -1894
box 250 218 480 436
use ntap  ntap_20
timestamp 1626065694
transform 1 0 18868 0 1 -1894
box 250 218 480 436
use ntap  ntap_19
timestamp 1626065694
transform 1 0 19886 0 1 -1894
box 250 218 480 436
use ntap  ntap_18
timestamp 1626065694
transform 1 0 7670 0 1 -742
box 250 218 480 436
use ntap  ntap_17
timestamp 1626065694
transform 1 0 8688 0 1 -742
box 250 218 480 436
use ntap  ntap_16
timestamp 1626065694
transform 1 0 9706 0 1 -742
box 250 218 480 436
use ntap  ntap_15
timestamp 1626065694
transform 1 0 10724 0 1 -742
box 250 218 480 436
use ntap  ntap_14
timestamp 1626065694
transform 1 0 11742 0 1 -742
box 250 218 480 436
use ntap  ntap_13
timestamp 1626065694
transform 1 0 12760 0 1 -742
box 250 218 480 436
use ntap  ntap_12
timestamp 1626065694
transform 1 0 13778 0 1 -742
box 250 218 480 436
use ntap  ntap_11
timestamp 1626065694
transform 1 0 14796 0 1 -742
box 250 218 480 436
use ntap  ntap_10
timestamp 1626065694
transform 1 0 15814 0 1 -742
box 250 218 480 436
use ntap  ntap_9
timestamp 1626065694
transform 1 0 16832 0 1 -742
box 250 218 480 436
use ntap  ntap_8
timestamp 1626065694
transform 1 0 17850 0 1 -742
box 250 218 480 436
use ntap  ntap_7
timestamp 1626065694
transform 1 0 18868 0 1 -742
box 250 218 480 436
use ntap  ntap_6
timestamp 1626065694
transform 1 0 19886 0 1 -742
box 250 218 480 436
use ntap  ntap_5
timestamp 1626065694
transform 1 0 20904 0 1 -3338
box 250 218 480 436
use ntap  ntap_4
timestamp 1626065694
transform 1 0 20904 0 1 -1894
box 250 218 480 436
use ntap  ntap_3
timestamp 1626065694
transform 1 0 21922 0 1 -3338
box 250 218 480 436
use ntap  ntap_2
timestamp 1626065694
transform 1 0 21922 0 1 -1894
box 250 218 480 436
use ntap  ntap_1
timestamp 1626065694
transform 1 0 21922 0 1 -742
box 250 218 480 436
use ntap  ntap_0
timestamp 1626065694
transform 1 0 20904 0 1 -742
box 250 218 480 436
use sky130_fd_pr__cap_mim_m3_1_VQCCU2  sky130_fd_pr__cap_mim_m3_1_VQCCU2_0
timestamp 1626065694
transform 1 0 -536 0 1 -1420
box -350 -1100 349 1100
use sky130_fd_pr__cap_mim_m3_1_VQCCU2  sky130_fd_pr__cap_mim_m3_1_VQCCU2_1
timestamp 1626065694
transform 1 0 -11930 0 1 -1420
box -350 -1100 349 1100
use sky130_fd_pr__cap_mim_m3_1_VQCCU2  sky130_fd_pr__cap_mim_m3_1_VQCCU2_2
timestamp 1626065694
transform 1 0 -536 0 1 -3920
box -350 -1100 349 1100
use sky130_fd_pr__cap_mim_m3_1_VQCCU2  sky130_fd_pr__cap_mim_m3_1_VQCCU2_3
timestamp 1626065694
transform 1 0 -11930 0 1 -3920
box -350 -1100 349 1100
use sky130_fd_pr__cap_mim_m3_1_VQCCU2  sky130_fd_pr__cap_mim_m3_1_VQCCU2_4
timestamp 1626065694
transform 1 0 -536 0 1 -6420
box -350 -1100 349 1100
use sky130_fd_pr__cap_mim_m3_1_VQCCU2  sky130_fd_pr__cap_mim_m3_1_VQCCU2_5
timestamp 1626065694
transform 1 0 -11930 0 1 -6420
box -350 -1100 349 1100
use sky130_fd_pr__cap_mim_m3_1_VQCCU2  sky130_fd_pr__cap_mim_m3_1_VQCCU2_6
timestamp 1626065694
transform 1 0 -536 0 1 -8920
box -350 -1100 349 1100
use sky130_fd_pr__cap_mim_m3_1_VQCCU2  sky130_fd_pr__cap_mim_m3_1_VQCCU2_7
timestamp 1626065694
transform 1 0 -11930 0 1 -8920
box -350 -1100 349 1100
<< labels >>
flabel metal2 s 9924 -2710 9924 -2710 1 FreeSans 600 0 0 0 vfoldm
flabel metal1 s 6356 -500 6356 -500 1 FreeSans 600 0 0 0 M1d
flabel metal1 s 7520 -2684 7520 -2684 1 FreeSans 600 0 0 0 M2d
flabel metal2 s 7798 -524 7798 -524 1 FreeSans 600 0 0 0 M6d
flabel metal1 s 7340 -3616 7340 -3616 1 FreeSans 600 0 0 0 M1d
flabel metal2 s 7618 -4582 7618 -4582 1 FreeSans 600 0 0 0 vbias1
flabel metal2 s 7514 -8154 7514 -8154 1 FreeSans 600 0 0 0 M2d
flabel metal2 s 16472 -5648 16472 -5648 1 FreeSans 600 0 0 0 M6d
flabel metal1 s 16668 -6000 16668 -6000 1 FreeSans 600 0 0 0 M13d
flabel metal2 s 11872 -8432 11872 -8432 1 FreeSans 600 0 0 0 M3d
flabel metal1 s 20726 -5618 20726 -5618 1 FreeSans 600 0 0 0 vfoldm
flabel metal2 s 20598 -6894 20598 -6894 1 FreeSans 600 0 0 0 vfoldp
flabel metal2 s 11830 716 11830 716 1 FreeSans 600 0 0 0 vfoldp
flabel metal2 s 3964 -6186 3964 -6186 1 FreeSans 600 0 0 0 vcmc_casc
flabel metal2 s 5800 -7134 5800 -7134 1 FreeSans 600 0 0 0 vcmcn_casc
flabel metal1 s 6080 -7670 6080 -7670 1 FreeSans 600 0 0 0 vcmcn2_casc
flabel metal1 s 3524 -7256 3524 -7256 1 FreeSans 600 0 0 0 vcmcn1_casc
flabel metal2 s 8324 850 8324 850 1 FreeSans 600 0 0 0 vbias1
flabel metal2 s 9302 588 9332 616 1 FreeSans 600 0 0 0 VDD
flabel metal1 s 2248 -17074 2270 -17046 1 FreeSans 600 0 0 0 vom
flabel metal2 s 12404 -15160 12436 -15142 1 FreeSans 600 0 0 0 vop
flabel metal1 s 23180 -18038 23204 -18008 1 FreeSans 600 0 0 0 VSS
flabel metal1 s 23556 -17190 23556 -17190 1 FreeSans 600 0 0 0 vbias3
flabel metal1 s 2144 -12732 2144 -12732 1 FreeSans 600 0 0 0 vcmc_casc
flabel metal1 s -2940 -20628 -2940 -20628 1 FreeSans 600 0 0 0 vcmn_casc_tail2
flabel metal2 s -3068 -20216 -3068 -20216 1 FreeSans 600 0 0 0 vcmn_casc_tail1
flabel metal1 s 132 -19622 132 -19622 1 FreeSans 600 0 0 0 vcmcn2_casc
flabel metal1 s -338 -20144 -338 -20144 1 FreeSans 600 0 0 0 vcmcn_casc
flabel metal1 s 18 -19488 18 -19488 1 FreeSans 600 0 0 0 vcmcn1_casc
flabel metal2 s -1114 -21516 -1114 -21516 1 FreeSans 600 0 0 0 vfoldp
flabel metal1 s 4648 -16436 4648 -16436 1 FreeSans 600 0 0 0 vcascnp
flabel metal1 s 23300 -16984 23300 -16984 1 FreeSans 600 0 0 0 vcascnm
flabel metal1 s 23436 -21216 23436 -21216 1 FreeSans 600 0 0 0 vbias4
flabel metal1 s 2006 -14484 2006 -14484 1 FreeSans 600 0 0 0 vtail_casc
flabel metal1 s 23678 -12816 23678 -12816 1 FreeSans 600 0 0 0 M3d
flabel metal1 s 22954 -15336 22954 -15336 1 FreeSans 600 0 0 0 M13d
flabel metal1 s 592 -22748 592 -22748 1 FreeSans 600 0 0 0 vtail_casc
flabel metal1 s -2092 -23816 -2092 -23816 1 FreeSans 600 0 0 0 vfoldm
flabel metal1 s -9506 -22906 -9506 -22906 1 FreeSans 600 0 0 0 vcmn_casc_tail2
flabel metal1 s -8364 -23636 -8364 -23636 1 FreeSans 600 0 0 0 vbias2
flabel metal1 s -4292 -23864 -4292 -23864 1 FreeSans 600 0 0 0 vcmn_casc_tail1
flabel metal1 s -8078 -12352 -8078 -12352 1 FreeSans 600 0 0 0 vbias1
flabel metal1 s -6206 -19026 -6206 -19026 1 FreeSans 600 0 0 0 vbias2
flabel metal4 s -1342 -5198 -1266 -5156 1 FreeSans 600 0 0 0 vom
flabel metal4 s -10820 -2704 -10756 -2664 1 FreeSans 600 0 0 0 vop
flabel metal1 s -2450 -19926 -2422 -19890 1 FreeSans 600 0 0 0 vom
flabel metal2 s -768 -19990 -736 -19968 1 FreeSans 600 0 0 0 vop
flabel metal1 s 17510 -4394 17546 -4366 1 FreeSans 600 0 0 0 VDD
flabel metal4 s -12400 -26800 -12400 -26800 3 FreeSans 4000 0 0 0 VSS
flabel metal1 s 1096 -23294 1122 -23264 1 FreeSans 600 0 0 0 vim
port 1 nsew
flabel metal1 s -2656 -23502 -2622 -23470 1 FreeSans 600 0 0 0 vip
port 2 nsew
flabel metal1 s -5330 -24996 -5294 -24960 1 FreeSans 600 0 0 0 VSS
port 3 nsew
flabel metal1 s -6348 -21586 -6316 -21566 1 FreeSans 600 0 0 0 ibiasn
port 4 nsew
flabel metal2 s -2498 -19392 -2424 -19358 1 FreeSans 600 0 0 0 vocm
port 5 nsew
flabel metal2 s 22386 -5742 22418 -5726 1 FreeSans 600 0 0 0 vom
port 6 nsew
flabel metal1 s 22574 -6900 22616 -6878 1 FreeSans 600 0 0 0 vop
port 7 nsew
flabel metal4 s -12400 1400 -12400 1400 3 FreeSans 4000 0 0 0 VDD
port 8 nsew
<< properties >>
string FIXED_BBOX -10872 -26372 24872 -10428
<< end >>
