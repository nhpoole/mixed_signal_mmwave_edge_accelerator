magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect -88575 -57856 91452 29600
<< nwell >>
rect -12082 15478 -10232 16318
rect -8617 15502 -7946 15800
rect -8617 15479 -8084 15502
rect -7962 15479 -7946 15502
<< locali >>
rect -8052 15471 -8004 15478
rect -8052 15437 -8045 15471
rect -8011 15437 -8004 15471
rect -8052 15430 -8004 15437
rect -7950 15475 -7902 15482
rect -7950 15441 -7943 15475
rect -7909 15441 -7902 15475
rect -7950 15434 -7902 15441
<< viali >>
rect -8045 15437 -8011 15471
rect -7943 15441 -7909 15475
<< metal1 >>
rect 47792 27680 48000 27710
rect -1414 27638 -1354 27648
rect -1414 27586 -1410 27638
rect -1358 27586 -1354 27638
rect -11462 16348 -10092 16408
rect -8742 16404 -8682 16414
rect -1414 16408 -1354 27586
rect 47792 27564 47854 27680
rect 47970 27564 48000 27680
rect 47022 25478 47376 25538
rect 47792 25514 48000 27564
rect 48306 27680 48488 27710
rect 48306 27564 48326 27680
rect 48442 27564 48488 27680
rect 48306 25497 48488 27564
rect 47022 23538 47082 25478
rect 47244 23930 47316 23934
rect 47244 23878 47254 23930
rect 47306 23878 47316 23930
rect 47244 23874 47316 23878
rect 47022 23478 47802 23538
rect 48682 23478 50478 23538
rect 46972 21916 47310 21920
rect 46972 21864 46982 21916
rect 47034 21864 47310 21916
rect 46972 21860 47310 21864
rect -8742 16352 -8738 16404
rect -8686 16352 -8682 16404
rect -8742 16342 -8682 16352
rect -1420 16404 -1348 16408
rect -1420 16352 -1410 16404
rect -1358 16352 -1348 16404
rect -1420 16348 -1348 16352
rect -8340 15714 -8100 15810
rect -8299 15471 -7992 15484
rect -8299 15437 -8045 15471
rect -8011 15437 -7992 15471
rect -8299 15424 -7992 15437
rect -7962 15475 -7734 15488
rect -7962 15441 -7943 15475
rect -7909 15441 -7734 15475
rect -7962 15428 -7734 15441
rect -8340 15170 -8100 15266
rect -12478 14956 -12418 15054
rect -12484 14952 -12412 14956
rect -9878 14952 -9818 15078
rect -12484 14900 -12474 14952
rect -12422 14900 -12412 14952
rect -12484 14896 -12412 14900
rect -9884 14948 -9812 14952
rect -9884 14896 -9874 14948
rect -9822 14896 -9812 14948
rect -9884 14892 -9812 14896
rect -10006 14833 -9946 14843
rect -10006 14781 -10002 14833
rect -9950 14781 -9946 14833
rect -10006 14771 -9946 14781
rect -10508 14712 -10502 14730
rect -11460 14652 -9402 14712
rect -8750 14708 -8690 14718
rect -8750 14656 -8746 14708
rect -8694 14656 -8690 14708
rect -8750 14646 -8690 14656
rect -1792 14712 -1732 14718
rect -1792 14708 -1294 14712
rect -1792 14656 -1788 14708
rect -1736 14656 -1294 14708
rect -1792 14652 -1294 14656
rect -1792 14646 -1732 14652
rect 48494 8574 48554 8578
rect 48494 8514 49142 8574
rect 50076 8546 50476 23478
rect 50938 9104 51010 9108
rect 50938 9052 50948 9104
rect 51000 9052 51010 9104
rect 50938 9048 51010 9052
rect 48358 7547 48430 7551
rect 48358 7495 48368 7547
rect 48420 7495 48430 7547
rect 48358 7491 48430 7495
rect 48364 6176 48424 7491
rect 48494 6610 48554 8514
rect 50944 7650 51004 9048
rect 50812 7590 51004 7650
rect 49766 6818 52704 6878
rect 48494 6550 48854 6610
rect 48358 6172 48430 6176
rect 48358 6120 48368 6172
rect 48420 6120 48430 6172
rect 48358 6116 48430 6120
rect 8274 5200 8346 5204
rect 8274 5148 8284 5200
rect 8336 5148 8346 5200
rect 8274 5144 8346 5148
rect 3944 4926 4244 4986
rect 8280 4788 8340 5144
rect 48494 4610 48554 6550
rect 50810 5626 51006 5686
rect 57932 4926 58226 4986
rect 49930 4854 52710 4914
rect 48494 4550 48994 4610
rect 48494 2520 48554 4550
rect 49960 2854 52704 2914
rect 48494 2462 49148 2520
rect 48498 2460 49148 2462
rect 50008 764 52706 824
<< via1 >>
rect -1410 27586 -1358 27638
rect 47854 27564 47970 27680
rect 48326 27564 48442 27680
rect 47254 23878 47306 23930
rect 46982 21864 47034 21916
rect -8738 16352 -8686 16404
rect -1410 16352 -1358 16404
rect -12474 14900 -12422 14952
rect -9874 14896 -9822 14948
rect -10002 14781 -9950 14833
rect -8746 14656 -8694 14708
rect -1788 14656 -1736 14708
rect 50948 9052 51000 9104
rect 48368 7495 48420 7547
rect 48368 6120 48420 6172
rect 8284 5148 8336 5200
<< metal2 >>
rect 47796 27680 48490 27702
rect -1414 27642 -1354 27651
rect 47796 27650 47854 27680
rect 47970 27650 48326 27680
rect 48442 27650 48490 27680
rect -1420 27640 -1348 27642
rect -1420 27584 -1412 27640
rect -1356 27584 -1348 27640
rect -1420 27582 -1348 27584
rect 47796 27594 47835 27650
rect 47971 27594 47995 27650
rect 48051 27594 48075 27650
rect 48131 27594 48155 27650
rect 48211 27594 48235 27650
rect 48291 27594 48315 27650
rect 48451 27594 48490 27650
rect -1414 27573 -1354 27582
rect 47796 27564 47854 27594
rect 47970 27564 48326 27594
rect 48442 27564 48490 27594
rect 47796 27536 48490 27564
rect 48230 24662 48467 24664
rect 48230 24606 48400 24662
rect 48456 24606 48467 24662
rect 48230 24604 48467 24606
rect 47615 24513 47782 24515
rect 47615 24457 47626 24513
rect 47682 24457 47782 24513
rect 47615 24455 47782 24457
rect 47250 23934 47310 23940
rect 42781 23932 47310 23934
rect 42781 23876 42792 23932
rect 42848 23930 47310 23932
rect 42848 23878 47254 23930
rect 47306 23878 47310 23930
rect 42848 23876 47310 23878
rect 42781 23874 47310 23876
rect 47250 23868 47310 23874
rect 38874 23861 38964 23866
rect 38870 23849 38968 23861
rect 38870 23793 38891 23849
rect 38947 23793 38968 23849
rect 38870 23781 38968 23793
rect 38874 23705 38964 23781
rect 38874 23615 41091 23705
rect 41001 23510 41091 23615
rect 41001 23454 41018 23510
rect 41074 23454 41091 23510
rect 41001 23428 41091 23454
rect 47867 22662 48046 22664
rect 47867 22606 47878 22662
rect 47934 22606 48046 22662
rect 47867 22604 48046 22606
rect 48514 22513 48725 22515
rect 48514 22457 48658 22513
rect 48714 22457 48725 22513
rect 48514 22455 48725 22457
rect 49519 22328 49579 24074
rect 46978 21920 47038 21926
rect 42791 21918 47038 21920
rect 42791 21862 42802 21918
rect 42858 21916 47038 21918
rect 42858 21864 46982 21916
rect 47034 21864 47038 21916
rect 42858 21862 47038 21864
rect 42791 21860 47038 21862
rect 46978 21854 47038 21860
rect 40228 21414 40328 21423
rect 36254 21392 40328 21414
rect 36254 21336 40250 21392
rect 40306 21336 40328 21392
rect 36254 21314 40328 21336
rect 11206 18913 11306 18918
rect 11202 18896 11310 18913
rect 11202 18840 11228 18896
rect 11284 18840 11310 18896
rect 11202 18823 11310 18840
rect -1414 16408 -1354 16414
rect -8748 16404 -1354 16408
rect -8748 16352 -8738 16404
rect -8686 16352 -1410 16404
rect -1358 16352 -1354 16404
rect -8748 16348 -1354 16352
rect -1414 16342 -1354 16348
rect 10953 16396 11071 16418
rect 10953 16340 10984 16396
rect 11040 16340 11071 16396
rect 10953 16318 11071 16340
rect -13295 15383 -12580 15385
rect -13295 15327 -13284 15383
rect -13228 15327 -12580 15383
rect -13295 15325 -12580 15327
rect -10629 15383 -10006 15385
rect -10629 15327 -10618 15383
rect -10562 15327 -10006 15383
rect -10629 15325 -10006 15327
rect -1933 15150 -1855 15152
rect -1933 15094 -1922 15150
rect -1866 15094 -1855 15150
rect -1933 15092 -1855 15094
rect -12478 14952 -12418 14962
rect -12478 14900 -12474 14952
rect -12422 14900 -12418 14952
rect -13467 14610 -13377 14614
rect -12478 14610 -12418 14900
rect -9878 14948 -9818 14958
rect -9878 14896 -9874 14948
rect -9822 14896 -9818 14948
rect -10838 14833 -9940 14837
rect -10838 14781 -10002 14833
rect -9950 14781 -9940 14833
rect -10838 14777 -9940 14781
rect -13472 14588 -12418 14610
rect -13472 14532 -13450 14588
rect -13394 14532 -12418 14588
rect -13472 14510 -12418 14532
rect -13467 14506 -13377 14510
rect -9878 14306 -9818 14896
rect -1924 14838 -1864 15092
rect 10962 14983 11062 16318
rect 11206 15882 11306 18823
rect 36254 16193 36354 21314
rect 40228 21305 40328 21314
rect 65088 18913 65188 18918
rect 65084 18896 65192 18913
rect 65084 18840 65110 18896
rect 65166 18840 65192 18896
rect 65084 18823 65192 18840
rect 43134 17841 43262 17846
rect 38968 17829 39076 17834
rect 38964 17808 39080 17829
rect 38964 17752 38994 17808
rect 39050 17752 39080 17808
rect 38964 17731 39080 17752
rect 43130 17810 43266 17841
rect 47326 17831 47436 17836
rect 43130 17754 43170 17810
rect 43226 17754 43266 17810
rect 38968 17668 39076 17731
rect 43130 17723 43266 17754
rect 47322 17809 47440 17831
rect 47322 17753 47353 17809
rect 47409 17753 47440 17809
rect 47322 17731 47440 17753
rect 43134 17694 43262 17723
rect 38968 17560 41102 17668
rect 43134 17566 45316 17694
rect 40994 17490 41102 17560
rect 40994 17434 41020 17490
rect 41076 17434 41102 17490
rect 40994 17399 41102 17434
rect 45188 17490 45316 17566
rect 47326 17669 47436 17731
rect 47326 17559 49393 17669
rect 45188 17434 45224 17490
rect 45280 17434 45316 17490
rect 45188 17389 45316 17434
rect 49283 17480 49393 17559
rect 49283 17424 49310 17480
rect 49366 17424 49393 17480
rect 49283 17388 49393 17424
rect 36250 16176 36358 16193
rect 36250 16120 36276 16176
rect 36332 16120 36358 16176
rect 36250 16103 36358 16120
rect 36254 16098 36354 16103
rect 11197 15860 11315 15882
rect 11197 15804 11228 15860
rect 11284 15804 11315 15860
rect 11197 15782 11315 15804
rect 10958 14966 11066 14983
rect 10958 14910 10984 14966
rect 11040 14910 11066 14966
rect 10958 14893 11066 14910
rect 10962 14888 11062 14893
rect -8360 14778 -1864 14838
rect 11206 14812 11306 15782
rect 11197 14790 11315 14812
rect 11197 14734 11228 14790
rect 11284 14734 11315 14790
rect 65088 14738 65188 18823
rect 11197 14712 11315 14734
rect 65079 14716 65197 14738
rect -8756 14708 -1726 14712
rect -8756 14656 -8746 14708
rect -8694 14656 -1788 14708
rect -1736 14656 -1726 14708
rect -8756 14652 -1726 14656
rect 65079 14660 65110 14716
rect 65166 14660 65197 14716
rect 65079 14638 65197 14660
rect -9878 14246 -9628 14306
rect -9688 13120 -9628 14246
rect 36456 13814 36556 13823
rect 39253 13814 39343 13818
rect 36456 13792 39348 13814
rect 36456 13736 36478 13792
rect 36534 13736 39270 13792
rect 39326 13736 39348 13792
rect 36456 13714 39348 13736
rect 36456 13705 36556 13714
rect 39253 13710 39343 13714
rect -9688 13064 -9686 13120
rect -9630 13064 -9628 13120
rect -9688 13053 -9628 13064
rect 42994 11727 43130 11732
rect 38844 11711 38950 11716
rect 38840 11691 38954 11711
rect 38840 11635 38869 11691
rect 38925 11635 38954 11691
rect 38840 11615 38954 11635
rect 42990 11690 43134 11727
rect 42990 11634 43034 11690
rect 43090 11634 43134 11690
rect 38844 11553 38950 11615
rect 42990 11597 43134 11634
rect 42994 11590 43134 11597
rect 38844 11447 40991 11553
rect 42994 11454 45158 11590
rect 40885 11356 40991 11447
rect 40885 11300 40910 11356
rect 40966 11300 40991 11356
rect 40885 11266 40991 11300
rect 45050 11366 45158 11454
rect 45050 11310 45076 11366
rect 45132 11310 45158 11366
rect 45050 11275 45158 11310
rect -9960 11043 -9846 11048
rect -9964 11019 -9842 11043
rect -5826 11027 -5720 11032
rect -9964 10963 -9931 11019
rect -9875 10963 -9842 11019
rect -9964 10939 -9842 10963
rect -5830 11007 -5716 11027
rect -5830 10951 -5801 11007
rect -5745 10951 -5716 11007
rect -9960 10871 -9846 10939
rect -5830 10931 -5716 10951
rect -5826 10891 -5720 10931
rect -9960 10757 -8667 10871
rect -5826 10785 -4683 10891
rect -8781 10696 -8667 10757
rect -8781 10640 -8752 10696
rect -8696 10640 -8667 10696
rect -8781 10602 -8667 10640
rect -4789 10690 -4683 10785
rect -4789 10634 -4764 10690
rect -4708 10634 -4683 10690
rect -4789 10600 -4683 10634
rect 36060 9306 36160 9315
rect 39009 9306 39099 9310
rect 36056 9284 39104 9306
rect 36056 9228 36082 9284
rect 36138 9228 39026 9284
rect 39082 9228 39104 9284
rect 36056 9206 39104 9228
rect 36060 9197 36160 9206
rect 39009 9202 39099 9206
rect 35833 9132 35935 9136
rect 35828 9104 51026 9132
rect 35828 9048 35856 9104
rect 35912 9052 50948 9104
rect 51000 9052 51026 9104
rect 35912 9048 51026 9052
rect 35828 9020 51026 9048
rect 35833 9016 35935 9020
rect 49704 7698 49891 7700
rect 49704 7642 49824 7698
rect 49880 7642 49891 7698
rect 49704 7640 49891 7642
rect 48364 7551 48424 7557
rect 48364 7547 49184 7551
rect 48364 7495 48368 7547
rect 48420 7495 49184 7547
rect 48364 7491 49184 7495
rect 48364 7485 48424 7491
rect 11382 7198 11442 7207
rect 9888 7196 11442 7198
rect 9888 7140 11384 7196
rect 11440 7140 11442 7196
rect 9888 7138 11442 7140
rect 62341 7196 62660 7198
rect 62341 7140 62352 7196
rect 62408 7140 62660 7196
rect 62341 7138 62660 7140
rect 11382 7129 11442 7138
rect 50834 6944 51160 7004
rect 45907 6176 48434 6198
rect 45907 6120 45938 6176
rect 45994 6172 48434 6176
rect 45994 6120 48368 6172
rect 48420 6120 48434 6172
rect 45907 6098 48434 6120
rect 49297 5734 49510 5736
rect 49297 5678 49308 5734
rect 49364 5678 49510 5734
rect 49297 5676 49510 5678
rect 49931 5585 50009 5587
rect 49931 5529 49942 5585
rect 49998 5529 50009 5585
rect 49931 5527 50009 5529
rect 8280 5204 8340 5210
rect 8271 5202 8349 5204
rect 8271 5146 8282 5202
rect 8338 5146 8349 5202
rect 8271 5144 8349 5146
rect 8280 5138 8340 5144
rect 38910 4099 39020 4104
rect 38906 4077 39024 4099
rect 43082 4097 43192 4102
rect 38906 4021 38937 4077
rect 38993 4021 39024 4077
rect 38906 3999 39024 4021
rect 43078 4075 43196 4097
rect 43078 4019 43109 4075
rect 43165 4019 43196 4075
rect 38910 3971 39020 3999
rect 43078 3997 43196 4019
rect 38910 3861 40895 3971
rect -10820 3835 -10716 3840
rect -10824 3816 -10712 3835
rect -6742 3827 -6642 3832
rect -10824 3760 -10796 3816
rect -10740 3760 -10712 3816
rect -10824 3741 -10712 3760
rect -6746 3810 -6638 3827
rect -6746 3754 -6720 3810
rect -6664 3754 -6638 3810
rect -10820 3688 -10716 3741
rect -6746 3737 -6638 3754
rect 40785 3772 40895 3861
rect 43082 3957 43192 3997
rect 43082 3847 45171 3957
rect -10820 3584 -8906 3688
rect -6742 3686 -6642 3737
rect 40785 3716 40812 3772
rect 40868 3716 40895 3772
rect -6742 3586 -4536 3686
rect 40785 3680 40895 3716
rect 45061 3760 45171 3847
rect 45061 3704 45088 3760
rect 45144 3704 45171 3760
rect 45061 3668 45171 3704
rect 49293 3734 49472 3736
rect 49293 3678 49304 3734
rect 49360 3678 49472 3734
rect 49293 3676 49472 3678
rect -9010 3490 -8906 3584
rect -9010 3434 -8986 3490
rect -8930 3434 -8906 3490
rect -9010 3401 -8906 3434
rect -4636 3488 -4536 3586
rect 49940 3585 50151 3587
rect 49940 3529 50084 3585
rect 50140 3529 50151 3585
rect 49940 3527 50151 3529
rect -4636 3432 -4614 3488
rect -4558 3432 -4536 3488
rect -4636 3401 -4536 3432
rect 50945 3400 51005 5146
rect 46079 1668 46157 1670
rect 8042 1566 9100 1626
rect 46079 1612 46090 1668
rect 46146 1612 46157 1668
rect 46079 1610 46157 1612
rect 49734 1644 49897 1646
rect 8042 582 8102 1566
rect 46088 1497 46148 1610
rect 49734 1588 49830 1644
rect 49886 1588 49897 1644
rect 51100 1596 51160 6944
rect 66017 4934 66095 4936
rect 66017 4878 66028 4934
rect 66084 4878 66095 4934
rect 66017 4876 66095 4878
rect 66026 3818 66086 4876
rect 65964 3758 66086 3818
rect 62153 2920 62243 2942
rect 62153 2916 62414 2920
rect 62153 2860 62170 2916
rect 62226 2860 62414 2916
rect 62153 2834 62243 2860
rect 49734 1586 49897 1588
rect 50940 1536 51160 1596
rect 46088 1437 49196 1497
rect 8033 580 8111 582
rect 8033 524 8044 580
rect 8100 524 8111 580
rect 8033 522 8111 524
<< via2 >>
rect -1412 27638 -1356 27640
rect -1412 27586 -1410 27638
rect -1410 27586 -1358 27638
rect -1358 27586 -1356 27638
rect -1412 27584 -1356 27586
rect 47835 27594 47854 27650
rect 47854 27594 47891 27650
rect 47915 27594 47970 27650
rect 47970 27594 47971 27650
rect 47995 27594 48051 27650
rect 48075 27594 48131 27650
rect 48155 27594 48211 27650
rect 48235 27594 48291 27650
rect 48315 27594 48326 27650
rect 48326 27594 48371 27650
rect 48395 27594 48442 27650
rect 48442 27594 48451 27650
rect 48400 24606 48456 24662
rect 47626 24457 47682 24513
rect 42792 23876 42848 23932
rect 38891 23793 38947 23849
rect 41018 23454 41074 23510
rect 47878 22606 47934 22662
rect 48658 22457 48714 22513
rect 42802 21862 42858 21918
rect 40250 21336 40306 21392
rect 11228 18840 11284 18896
rect 10984 16340 11040 16396
rect -13284 15327 -13228 15383
rect -10618 15327 -10562 15383
rect -1922 15094 -1866 15150
rect -13450 14532 -13394 14588
rect 65110 18840 65166 18896
rect 38994 17752 39050 17808
rect 43170 17754 43226 17810
rect 47353 17753 47409 17809
rect 41020 17434 41076 17490
rect 45224 17434 45280 17490
rect 49310 17424 49366 17480
rect 36276 16120 36332 16176
rect 11228 15804 11284 15860
rect 10984 14910 11040 14966
rect 11228 14734 11284 14790
rect 65110 14660 65166 14716
rect 36478 13736 36534 13792
rect 39270 13736 39326 13792
rect -9686 13064 -9630 13120
rect 38869 11635 38925 11691
rect 43034 11634 43090 11690
rect 40910 11300 40966 11356
rect 45076 11310 45132 11366
rect -9931 10963 -9875 11019
rect -5801 10951 -5745 11007
rect -8752 10640 -8696 10696
rect -4764 10634 -4708 10690
rect 36082 9228 36138 9284
rect 39026 9228 39082 9284
rect 35856 9048 35912 9104
rect 49824 7642 49880 7698
rect 11384 7140 11440 7196
rect 62352 7140 62408 7196
rect 45938 6120 45994 6176
rect 49308 5678 49364 5734
rect 49942 5529 49998 5585
rect 8282 5200 8338 5202
rect 8282 5148 8284 5200
rect 8284 5148 8336 5200
rect 8336 5148 8338 5200
rect 8282 5146 8338 5148
rect 38937 4021 38993 4077
rect 43109 4019 43165 4075
rect -10796 3760 -10740 3816
rect -6720 3754 -6664 3810
rect 40812 3716 40868 3772
rect 45088 3704 45144 3760
rect 49304 3678 49360 3734
rect -8986 3434 -8930 3490
rect 50084 3529 50140 3585
rect -4614 3432 -4558 3488
rect 46090 1612 46146 1668
rect 49830 1588 49886 1644
rect 66028 4878 66084 4934
rect 62170 2860 62226 2916
rect 8044 524 8100 580
<< metal3 >>
rect -1436 27647 -1330 27668
rect -1436 27583 -1416 27647
rect -1352 27583 -1330 27647
rect -1436 27562 -1330 27583
rect 47796 27654 48490 27702
rect 47796 27590 47831 27654
rect 47895 27590 47911 27654
rect 47975 27590 47991 27654
rect 48055 27590 48071 27654
rect 48135 27590 48151 27654
rect 48215 27590 48231 27654
rect 48295 27590 48311 27654
rect 48375 27590 48391 27654
rect 48455 27590 48490 27654
rect 47796 27536 48490 27590
rect 38430 26566 38578 26574
rect 38430 26494 38432 26566
rect 37160 26422 38432 26494
rect 38576 26494 38578 26566
rect 41348 26561 41506 26574
rect 41348 26494 41355 26561
rect 38576 26422 41355 26494
rect 37160 26417 41355 26422
rect 41499 26494 41506 26561
rect 41499 26417 42865 26494
rect 37160 25893 42865 26417
rect 37160 24776 37761 25893
rect 41522 25880 42865 25893
rect 37044 24742 37761 24776
rect 37044 24678 37084 24742
rect 37148 24678 37761 24742
rect 37044 24644 37761 24678
rect 36462 23552 36574 23570
rect 36462 23488 36486 23552
rect 36550 23488 36574 23552
rect 36462 23470 36574 23488
rect 36468 20168 36568 23470
rect 37160 22676 37761 24644
rect 42251 24768 42865 25880
rect 42251 24732 43054 24768
rect 42251 24668 42948 24732
rect 43012 24668 43054 24732
rect 42251 24632 43054 24668
rect 48378 24662 51894 24688
rect 38874 23849 38964 23912
rect 40401 23870 40503 24099
rect 42251 23932 42865 24632
rect 48378 24606 48400 24662
rect 48456 24606 51894 24662
rect 48378 24588 51894 24606
rect 46576 24534 46676 24540
rect 46576 24516 47704 24534
rect 46576 24452 46594 24516
rect 46658 24513 47704 24516
rect 46658 24457 47626 24513
rect 47682 24457 47704 24513
rect 46658 24452 47704 24457
rect 46576 24434 47704 24452
rect 46576 24428 46676 24434
rect 42251 23876 42792 23932
rect 42848 23876 42865 23932
rect 38874 23793 38891 23849
rect 38947 23793 38964 23849
rect 38874 23776 38964 23793
rect 40396 23852 40508 23870
rect 40396 23788 40420 23852
rect 40484 23788 40508 23852
rect 40396 23770 40508 23788
rect 40401 23769 40503 23770
rect 41563 23712 41661 23717
rect 42030 23712 42130 23718
rect 41562 23694 42130 23712
rect 41562 23630 41580 23694
rect 41644 23630 42048 23694
rect 42112 23630 42130 23694
rect 41562 23612 42130 23630
rect 41563 23607 41661 23612
rect 42030 23606 42130 23612
rect 39492 23567 39592 23568
rect 39487 23550 39597 23567
rect 39487 23486 39510 23550
rect 39574 23486 39597 23550
rect 39487 23469 39597 23486
rect 40996 23510 41096 23532
rect 39492 23348 39592 23469
rect 40996 23454 41018 23510
rect 41074 23454 41096 23510
rect 40996 23432 41096 23454
rect 41001 23229 41091 23432
rect 37070 22648 37761 22676
rect 37070 22584 37104 22648
rect 37168 22584 37761 22648
rect 37070 22556 37761 22584
rect 37160 21038 37761 22556
rect 42251 22658 42865 23876
rect 46404 22662 47952 22684
rect 42251 22620 43010 22658
rect 42251 22556 42902 22620
rect 42966 22556 43010 22620
rect 42251 22518 43010 22556
rect 46404 22606 47878 22662
rect 47934 22606 47952 22662
rect 46404 22584 47952 22606
rect 40228 21419 40328 22002
rect 42251 21918 42865 22518
rect 42251 21862 42802 21918
rect 42858 21862 42865 21918
rect 40223 21392 40333 21419
rect 40223 21336 40250 21392
rect 40306 21336 40333 21392
rect 40223 21309 40333 21336
rect 42251 21038 42865 21862
rect 46404 21381 46504 22584
rect 48640 22513 49860 22532
rect 48640 22457 48658 22513
rect 48714 22457 49860 22513
rect 48640 22432 49860 22457
rect 49760 21682 49860 22432
rect 49760 21618 49778 21682
rect 49842 21618 49860 21682
rect 49760 21594 49860 21618
rect 46399 21364 46509 21381
rect 46399 21300 46422 21364
rect 46486 21300 46509 21364
rect 46399 21283 46509 21300
rect 46404 21282 46504 21283
rect 51794 21066 51894 24588
rect 52138 23696 52250 23714
rect 52138 23632 52162 23696
rect 52226 23632 52250 23696
rect 52138 23614 52250 23632
rect 51788 21048 51900 21066
rect 37160 20828 51393 21038
rect 51788 20984 51812 21048
rect 51876 20984 51900 21048
rect 51788 20966 51900 20984
rect 37160 20473 40646 20828
rect 37160 20437 38511 20473
rect 37279 20420 38511 20437
rect 36468 19925 36572 20168
rect 36467 19908 36577 19925
rect 36467 19844 36490 19908
rect 36554 19844 36577 19908
rect 36467 19827 36577 19844
rect 11036 18896 11638 18918
rect 11036 18840 11228 18896
rect 11284 18840 11638 18896
rect 11036 18818 11638 18840
rect 36468 17152 36572 19827
rect 37279 19649 37879 20420
rect 38494 20329 38511 20420
rect 38655 20456 40646 20473
rect 40846 20473 51393 20828
rect 40846 20456 40911 20473
rect 38655 20420 40911 20456
rect 38655 20329 38672 20420
rect 38494 20306 38672 20329
rect 40894 20329 40911 20420
rect 41055 20420 43311 20473
rect 41055 20329 41072 20420
rect 40894 20306 41072 20329
rect 43294 20329 43311 20420
rect 43455 20420 45437 20473
rect 43455 20329 43472 20420
rect 43294 20306 43472 20329
rect 45420 20329 45437 20420
rect 45581 20420 47611 20473
rect 45581 20329 45598 20420
rect 45420 20306 45598 20329
rect 47594 20329 47611 20420
rect 47755 20420 50011 20473
rect 47755 20329 47772 20420
rect 47594 20306 47772 20329
rect 49994 20329 50011 20420
rect 50155 20420 51393 20473
rect 50155 20329 50172 20420
rect 49994 20306 50172 20329
rect 39072 19908 46764 19926
rect 39072 19844 39096 19908
rect 39160 19844 46764 19908
rect 39072 19826 46764 19844
rect 37279 18790 37881 19649
rect 39682 19460 39782 19826
rect 42460 19512 42560 19826
rect 46664 19432 46764 19826
rect 37144 18758 37881 18790
rect 37144 18614 37182 18758
rect 37326 18614 37881 18758
rect 37144 18582 37881 18614
rect 36468 17048 36852 17152
rect 10957 16396 11067 16423
rect 10957 16340 10984 16396
rect 11040 16340 11067 16396
rect 10957 16313 11067 16340
rect 11464 16322 36558 16422
rect 36254 16176 36354 16198
rect 36254 16120 36276 16176
rect 36332 16120 36354 16176
rect 11201 15882 11311 15887
rect 11201 15860 36158 15882
rect 11201 15804 11228 15860
rect 11284 15804 36158 15860
rect 11201 15782 36158 15804
rect 11201 15777 11311 15782
rect -13304 15383 -13204 15396
rect -13304 15327 -13284 15383
rect -13228 15327 -13204 15383
rect -13304 14732 -13204 15327
rect -10642 15383 -10542 15410
rect -10642 15327 -10618 15383
rect -10562 15327 -10542 15383
rect -10642 14732 -10542 15327
rect -1950 15150 35940 15182
rect -1950 15094 -1922 15150
rect -1866 15094 35940 15150
rect -1950 15070 35940 15094
rect -13304 14632 -10542 14732
rect -2396 14966 11062 14988
rect -2396 14910 10984 14966
rect 11040 14910 11062 14966
rect -2396 14888 11062 14910
rect -13472 14588 -13372 14610
rect -13472 14532 -13450 14588
rect -13394 14532 -13372 14588
rect -13472 10731 -13372 14532
rect -13477 10714 -13367 10731
rect -13477 10650 -13454 10714
rect -13390 10650 -13367 10714
rect -13477 10633 -13367 10650
rect -13472 10632 -13372 10633
rect -13304 3537 -13204 14632
rect -11154 14167 -11008 14174
rect -11154 14023 -11153 14167
rect -11009 14023 -11008 14167
rect -11154 14002 -11008 14023
rect -8836 14151 -8646 14180
rect -3940 14161 -3782 14174
rect -8836 14007 -8813 14151
rect -8669 14007 -8646 14151
rect -8836 14002 -8646 14007
rect -6346 14134 -6170 14156
rect -6346 14002 -6330 14134
rect -12476 13990 -6330 14002
rect -6186 14002 -6170 14134
rect -3940 14017 -3933 14161
rect -3789 14017 -3782 14161
rect -3940 14002 -3782 14017
rect -6186 13990 -2606 14002
rect -12476 13400 -2606 13990
rect -12476 13398 -7666 13400
rect -13108 13137 -13008 13138
rect -13113 13120 -13003 13137
rect -13113 13056 -13090 13120
rect -13026 13056 -13003 13120
rect -13113 13039 -13003 13056
rect -13108 12772 -13006 13039
rect -13106 9154 -13006 12772
rect -12476 11974 -11875 13398
rect -10580 13120 -7214 13138
rect -10580 13056 -10556 13120
rect -10492 13064 -9686 13120
rect -9630 13064 -7214 13120
rect -10492 13056 -7214 13064
rect -10580 13038 -7214 13056
rect -9994 12784 -9894 13038
rect -12630 11959 -11875 11974
rect -12630 11895 -12609 11959
rect -12545 11895 -11875 11959
rect -12630 11880 -11875 11895
rect -12476 10010 -11875 11880
rect -9960 11192 -9894 12784
rect -7314 12716 -7214 13038
rect -3207 12166 -2606 13400
rect -2396 12904 -2296 14888
rect 11201 14812 11311 14817
rect 10974 14810 11311 14812
rect -1756 14790 11311 14810
rect -1756 14734 11228 14790
rect 11284 14734 11311 14790
rect -1756 14710 11311 14734
rect -2402 12886 -2290 12904
rect -2402 12822 -2378 12886
rect -2314 12822 -2290 12886
rect -2402 12804 -2290 12822
rect -3207 11856 -2604 12166
rect -3207 11842 -2426 11856
rect -3207 11778 -2510 11842
rect -2446 11778 -2426 11842
rect -3207 11764 -2426 11778
rect -3207 11566 -2604 11764
rect -9960 11019 -9846 11128
rect -9226 11029 -9126 11252
rect -9960 10963 -9931 11019
rect -9875 10963 -9846 11019
rect -9960 10934 -9846 10963
rect -9231 11012 -9121 11029
rect -9231 10948 -9208 11012
rect -9144 10948 -9121 11012
rect -9231 10931 -9121 10948
rect -5826 11007 -5720 11164
rect -5270 11029 -5170 11234
rect -5826 10951 -5801 11007
rect -5745 10951 -5720 11007
rect -9226 10930 -9126 10931
rect -5826 10926 -5720 10951
rect -5275 11012 -5165 11029
rect -5275 10948 -5252 11012
rect -5188 10948 -5165 11012
rect -5275 10931 -5165 10948
rect -5270 10930 -5170 10931
rect -8101 10882 -8003 10887
rect -7570 10882 -7470 10888
rect -8102 10864 -7470 10882
rect -3901 10880 -3803 10885
rect -3392 10880 -3292 10886
rect -8102 10800 -8084 10864
rect -8020 10800 -7552 10864
rect -7488 10800 -7470 10864
rect -8102 10782 -7470 10800
rect -8101 10777 -8003 10782
rect -7570 10776 -7470 10782
rect -3902 10862 -3288 10880
rect -3902 10798 -3884 10862
rect -3820 10798 -3374 10862
rect -3310 10798 -3288 10862
rect -3902 10780 -3288 10798
rect -3901 10775 -3803 10780
rect -3392 10774 -3292 10780
rect -6556 10733 -6456 10734
rect -10356 10731 -10256 10732
rect -10361 10714 -10251 10731
rect -10361 10650 -10338 10714
rect -10274 10650 -10251 10714
rect -10361 10633 -10251 10650
rect -8786 10696 -8662 10730
rect -8786 10640 -8752 10696
rect -8696 10640 -8662 10696
rect -6561 10716 -6451 10733
rect -10356 10588 -10256 10633
rect -8786 10606 -8662 10640
rect -10356 10476 -10202 10588
rect -10302 10450 -10202 10476
rect -12640 10002 -11875 10010
rect -12640 9938 -12626 10002
rect -12562 9938 -11875 10002
rect -12640 9930 -11875 9938
rect -13106 9054 -12632 9154
rect -13100 8619 -13000 8620
rect -13105 8602 -12995 8619
rect -13105 8538 -13082 8602
rect -13018 8538 -12995 8602
rect -13105 8521 -12995 8538
rect -13309 3520 -13199 3537
rect -13309 3456 -13286 3520
rect -13222 3456 -13199 3520
rect -13309 3439 -13199 3456
rect -13304 3438 -13204 3439
rect -13100 1627 -13000 8521
rect -12732 5665 -12632 9054
rect -12476 8260 -11875 9930
rect -10132 8620 -10032 10450
rect -8781 10315 -8667 10606
rect -7192 10492 -7190 10684
rect -6561 10652 -6538 10716
rect -6474 10652 -6451 10716
rect -6561 10635 -6451 10652
rect -4794 10690 -4678 10720
rect -6556 10476 -6456 10635
rect -4794 10634 -4764 10690
rect -4708 10634 -4678 10690
rect -4794 10604 -4678 10634
rect -4789 10433 -4683 10604
rect -3207 9848 -2606 11566
rect -1756 11018 -1656 14710
rect 11201 14707 11311 14710
rect -3207 9827 -2406 9848
rect -3207 9763 -2497 9827
rect -2433 9763 -2406 9827
rect -3207 9742 -2406 9763
rect -7192 8620 -7092 9154
rect -10540 8602 -7092 8620
rect -10540 8538 -10516 8602
rect -10452 8538 -7092 8602
rect -10540 8520 -7092 8538
rect -6953 8262 -6351 8264
rect -5974 8262 -4547 8264
rect -4183 8262 -3581 8264
rect -3207 8262 -2606 9742
rect -1758 8863 -1656 11018
rect 35828 9104 35940 15070
rect 36058 9716 36158 15782
rect 36254 15375 36354 16120
rect 36249 15358 36359 15375
rect 36249 15294 36272 15358
rect 36336 15294 36359 15358
rect 36249 15277 36359 15294
rect 35828 9048 35856 9104
rect 35912 9048 35940 9104
rect 35828 9020 35940 9048
rect 36054 9311 36158 9716
rect 36254 9541 36354 15277
rect 36458 13819 36558 16322
rect 36451 13792 36561 13819
rect 36451 13736 36478 13792
rect 36534 13736 36561 13792
rect 36451 13709 36561 13736
rect 36249 9524 36359 9541
rect 36249 9460 36272 9524
rect 36336 9460 36359 9524
rect 36249 9443 36359 9460
rect 36254 9442 36354 9443
rect 36054 9284 36165 9311
rect 36054 9228 36082 9284
rect 36138 9228 36165 9284
rect 36054 9201 36165 9228
rect -1761 8846 -1651 8863
rect -1761 8782 -1738 8846
rect -1674 8782 -1651 8846
rect -1761 8765 -1651 8782
rect -11351 8260 -2606 8262
rect -12476 7662 -2606 8260
rect 35229 7738 35327 7743
rect 11362 7720 35328 7738
rect -12476 7660 -6020 7662
rect -4183 7660 -3581 7662
rect -11204 7638 -10950 7660
rect -11204 7414 -11189 7638
rect -10965 7556 -10950 7638
rect -8792 7638 -8538 7660
rect -10965 7414 -10951 7556
rect -11204 7406 -10951 7414
rect -8792 7414 -8777 7638
rect -8553 7556 -8538 7638
rect -6380 7638 -6126 7660
rect -8553 7414 -8539 7556
rect -8792 7406 -8539 7414
rect -6380 7414 -6365 7638
rect -6141 7556 -6126 7638
rect -3968 7638 -3714 7660
rect -6141 7414 -6127 7556
rect -6380 7406 -6127 7414
rect -3968 7414 -3953 7638
rect -3729 7556 -3714 7638
rect 11362 7656 35246 7720
rect 35310 7656 35328 7720
rect 11362 7638 35328 7656
rect -3729 7414 -3715 7556
rect -3968 7406 -3715 7414
rect -11204 7047 -10954 7406
rect -11204 6823 -11189 7047
rect -10965 6823 -10954 7047
rect -11204 6812 -10954 6823
rect -8792 7047 -8542 7406
rect -8792 6823 -8777 7047
rect -8553 6823 -8542 7047
rect -8792 6812 -8542 6823
rect -6380 7047 -6130 7406
rect -6380 6823 -6365 7047
rect -6141 6823 -6130 7047
rect -6380 6812 -6130 6823
rect -3968 7047 -3718 7406
rect 11362 7196 11462 7638
rect 35229 7633 35327 7638
rect 11362 7140 11384 7196
rect 11440 7140 11462 7196
rect 11362 7102 11462 7140
rect -3968 6823 -3953 7047
rect -3729 6823 -3718 7047
rect -3968 6812 -3718 6823
rect -12474 6798 -2604 6812
rect -12475 6712 -2604 6798
rect -12475 6198 -2607 6712
rect -12737 5648 -12627 5665
rect -12737 5584 -12714 5648
rect -12650 5584 -12627 5648
rect -12737 5567 -12627 5584
rect -12732 5566 -12632 5567
rect -12475 4766 -11875 6198
rect -12592 4763 -11875 4766
rect -12592 4619 -12583 4763
rect -12439 4619 -11875 4763
rect -12592 4616 -11875 4619
rect -12475 2650 -11875 4616
rect -9948 5852 -7198 5952
rect -9948 4138 -9848 5852
rect -7298 5478 -7198 5852
rect -3207 4716 -2607 6198
rect -2426 5665 -2322 5666
rect -2427 5648 -2317 5665
rect -2427 5584 -2404 5648
rect -2340 5584 -2317 5648
rect -2427 5567 -2317 5584
rect -2426 5228 -2322 5567
rect -2426 5226 8314 5228
rect -2426 5202 8366 5226
rect -2426 5146 8282 5202
rect 8338 5146 8366 5202
rect -2426 5126 8366 5146
rect -2426 5124 8314 5126
rect -3207 4711 -2500 4716
rect -3207 4567 -2655 4711
rect -2511 4567 -2500 4711
rect -3207 4562 -2500 4567
rect -10820 3816 -10716 3856
rect -9366 3827 -9266 4098
rect -10820 3760 -10796 3816
rect -10740 3760 -10716 3816
rect -10820 3736 -10716 3760
rect -9371 3810 -9261 3827
rect -9371 3746 -9348 3810
rect -9284 3746 -9261 3810
rect -9371 3729 -9261 3746
rect -6742 3810 -6642 3888
rect -5144 3839 -5028 4060
rect -6742 3754 -6720 3810
rect -6664 3754 -6642 3810
rect -6742 3732 -6642 3754
rect -5149 3814 -5023 3839
rect -5149 3750 -5118 3814
rect -5054 3750 -5023 3814
rect -9366 3728 -9266 3729
rect -5149 3725 -5023 3750
rect -5144 3724 -5028 3725
rect -8085 3682 -7987 3687
rect -7554 3682 -7454 3688
rect -3885 3684 -3787 3689
rect -3382 3684 -3282 3690
rect -8086 3664 -7454 3682
rect -8086 3600 -8068 3664
rect -8004 3600 -7536 3664
rect -7472 3600 -7454 3664
rect -8086 3582 -7454 3600
rect -3886 3666 -3282 3684
rect -3886 3602 -3868 3666
rect -3804 3602 -3364 3666
rect -3300 3602 -3282 3666
rect -3886 3584 -3282 3602
rect -8085 3577 -7987 3582
rect -7554 3576 -7454 3582
rect -3885 3579 -3787 3584
rect -3382 3578 -3282 3584
rect -10168 3537 -10068 3538
rect -10173 3520 -10063 3537
rect -10173 3456 -10150 3520
rect -10086 3456 -10063 3520
rect -10173 3439 -10063 3456
rect -9015 3490 -8901 3519
rect -10168 3194 -10068 3439
rect -9015 3434 -8986 3490
rect -8930 3434 -8901 3490
rect -5914 3516 -5786 3542
rect -5914 3452 -5882 3516
rect -5818 3452 -5786 3516
rect -9015 3405 -8901 3434
rect -9010 3238 -8906 3405
rect -7176 3254 -7174 3446
rect -5914 3426 -5786 3452
rect -4641 3488 -4531 3515
rect -4641 3432 -4614 3488
rect -4558 3432 -4531 3488
rect -5908 3332 -5792 3426
rect -4641 3405 -4531 3432
rect -4636 3174 -4536 3405
rect -12586 2619 -11875 2650
rect -12586 2555 -12549 2619
rect -12485 2555 -11875 2619
rect -12586 2524 -11875 2555
rect -13103 1610 -12993 1627
rect -13103 1546 -13080 1610
rect -13016 1546 -12993 1610
rect -13103 1529 -12993 1546
rect -13100 1528 -13000 1529
rect -12475 1062 -11875 2524
rect -10086 1422 -9986 3082
rect -3207 3060 -2607 4562
rect -3207 2664 -2608 3060
rect -3207 2656 -2500 2664
rect -3207 2512 -2658 2656
rect -2514 2512 -2500 2656
rect -3207 2504 -2500 2512
rect -3207 2202 -2608 2504
rect 36054 2238 36158 9201
rect 36458 6197 36558 13709
rect 36748 13581 36852 17048
rect 37279 16650 37881 18582
rect 50792 18732 51393 20420
rect 50792 18723 51506 18732
rect 50792 18579 51347 18723
rect 51491 18579 51506 18723
rect 50792 18570 51506 18579
rect 38968 17808 39076 17892
rect 40416 17829 40516 18064
rect 38968 17752 38994 17808
rect 39050 17752 39076 17808
rect 38968 17726 39076 17752
rect 40411 17812 40521 17829
rect 40411 17748 40434 17812
rect 40498 17748 40521 17812
rect 40411 17731 40521 17748
rect 43134 17810 43262 17960
rect 44642 17817 44742 18054
rect 43134 17754 43170 17810
rect 43226 17754 43262 17810
rect 40416 17730 40516 17731
rect 43134 17718 43262 17754
rect 44637 17800 44747 17817
rect 44637 17736 44660 17800
rect 44724 17736 44747 17800
rect 44637 17719 44747 17736
rect 47326 17809 47436 17902
rect 48764 17827 48864 18046
rect 47326 17753 47353 17809
rect 47409 17753 47436 17809
rect 47326 17726 47436 17753
rect 48759 17810 48869 17827
rect 48759 17746 48782 17810
rect 48846 17746 48869 17810
rect 48759 17729 48869 17746
rect 48764 17728 48864 17729
rect 44642 17718 44742 17719
rect 41673 17678 41771 17683
rect 42204 17678 42304 17684
rect 45873 17678 45971 17683
rect 46404 17678 46504 17684
rect 50073 17678 50171 17683
rect 50604 17678 50704 17684
rect 41672 17660 42304 17678
rect 41672 17596 41690 17660
rect 41754 17596 42222 17660
rect 42286 17596 42304 17660
rect 41672 17578 42304 17596
rect 45872 17660 46504 17678
rect 45872 17596 45890 17660
rect 45954 17596 46422 17660
rect 46486 17596 46504 17660
rect 45872 17578 46504 17596
rect 50072 17660 50704 17678
rect 50072 17596 50090 17660
rect 50154 17596 50622 17660
rect 50686 17596 50704 17660
rect 50072 17578 50704 17596
rect 41673 17573 41771 17578
rect 42204 17572 42304 17578
rect 45873 17573 45971 17578
rect 46404 17572 46504 17578
rect 50073 17573 50171 17578
rect 50604 17572 50704 17578
rect 39618 17523 39718 17524
rect 43818 17523 43918 17524
rect 39613 17506 39723 17523
rect 39613 17442 39636 17506
rect 39700 17442 39723 17506
rect 39613 17425 39723 17442
rect 40989 17490 41107 17521
rect 40989 17434 41020 17490
rect 41076 17434 41107 17490
rect 39618 17384 39718 17425
rect 40989 17403 41107 17434
rect 43813 17506 43923 17523
rect 43813 17442 43836 17506
rect 43900 17442 43923 17506
rect 43813 17425 43923 17442
rect 45183 17490 45321 17531
rect 48018 17521 48118 17522
rect 45183 17434 45224 17490
rect 45280 17434 45321 17490
rect 39618 17272 39772 17384
rect 37073 16629 37881 16650
rect 37073 16485 37100 16629
rect 37244 16485 37881 16629
rect 37073 16464 37881 16485
rect 37279 14870 37881 16464
rect 39672 15376 39772 17272
rect 40994 17156 41102 17403
rect 43818 17272 43918 17425
rect 45183 17393 45321 17434
rect 48013 17504 48123 17521
rect 48013 17440 48036 17504
rect 48100 17440 48123 17504
rect 48013 17423 48123 17440
rect 49278 17480 49398 17512
rect 49278 17424 49310 17480
rect 49366 17424 49398 17480
rect 45188 17194 45316 17393
rect 48018 17272 48118 17423
rect 49278 17392 49398 17424
rect 49283 17165 49393 17392
rect 50792 16638 51393 18570
rect 50792 16626 51538 16638
rect 50792 16482 51376 16626
rect 51520 16482 51538 16626
rect 50792 16470 51538 16482
rect 42582 15376 42682 15950
rect 46660 15376 46760 15844
rect 39292 15358 46760 15376
rect 39292 15294 39316 15358
rect 39380 15294 46760 15358
rect 39292 15276 46760 15294
rect 50792 14870 51393 16470
rect 37131 14309 51393 14870
rect 52144 14738 52244 23614
rect 65088 18896 65188 18918
rect 65088 18840 65110 18896
rect 65166 18840 65188 18896
rect 65088 18818 65188 18840
rect 52380 15100 52480 15106
rect 64976 15100 65076 16422
rect 52380 15082 65076 15100
rect 52380 15018 52398 15082
rect 52462 15018 65076 15082
rect 52380 15000 65076 15018
rect 52380 14994 52480 15000
rect 65083 14738 65193 14743
rect 52144 14716 65193 14738
rect 52144 14660 65110 14716
rect 65166 14660 65193 14716
rect 52144 14638 65193 14660
rect 65083 14633 65193 14638
rect 37131 14260 38485 14309
rect 36743 13564 36853 13581
rect 36743 13500 36766 13564
rect 36830 13500 36853 13564
rect 36743 13483 36853 13500
rect 37131 13527 37731 14260
rect 38478 14165 38485 14260
rect 38629 14260 40897 14309
rect 38629 14165 38636 14260
rect 38478 14152 38636 14165
rect 40890 14165 40897 14260
rect 41041 14260 43297 14309
rect 41041 14165 41048 14260
rect 40890 14152 41048 14165
rect 43290 14165 43297 14260
rect 43441 14260 45697 14309
rect 43441 14165 43448 14260
rect 43290 14152 43448 14165
rect 45690 14165 45697 14260
rect 45841 14268 47697 14309
rect 45841 14260 46992 14268
rect 45841 14165 45848 14260
rect 45690 14152 45848 14165
rect 39248 13792 42430 13814
rect 39248 13736 39270 13792
rect 39326 13736 42430 13792
rect 39248 13714 42430 13736
rect 36748 13480 36852 13483
rect 37131 12668 37733 13527
rect 39568 13134 39668 13714
rect 42330 13394 42430 13714
rect 36996 12636 37733 12668
rect 36996 12492 37034 12636
rect 37178 12492 37733 12636
rect 36996 12460 37733 12492
rect 37131 10528 37733 12460
rect 46399 12734 46992 14260
rect 47690 14165 47697 14268
rect 47841 14268 50097 14309
rect 47841 14165 47848 14268
rect 47690 14152 47848 14165
rect 50090 14165 50097 14268
rect 50241 14268 51393 14309
rect 50241 14165 50248 14268
rect 50792 14264 51393 14268
rect 50090 14152 50248 14165
rect 46399 12610 46999 12734
rect 46399 12601 47198 12610
rect 46399 12457 47039 12601
rect 47183 12457 47198 12601
rect 46399 12448 47198 12457
rect 46399 12380 46999 12448
rect 38844 11691 38950 11868
rect 40292 11709 40392 11914
rect 38844 11635 38869 11691
rect 38925 11635 38950 11691
rect 38844 11610 38950 11635
rect 40287 11692 40397 11709
rect 40287 11628 40310 11692
rect 40374 11628 40397 11692
rect 40287 11611 40397 11628
rect 42994 11690 43130 11854
rect 44512 11709 44612 11890
rect 42994 11634 43034 11690
rect 43090 11634 43130 11690
rect 40292 11610 40392 11611
rect 42994 11592 43130 11634
rect 44507 11692 44617 11709
rect 44507 11628 44530 11692
rect 44594 11628 44617 11692
rect 44507 11611 44617 11628
rect 44512 11610 44612 11611
rect 41543 11560 41641 11565
rect 42074 11560 42174 11566
rect 45743 11560 45841 11565
rect 46218 11560 46318 11566
rect 41542 11542 42174 11560
rect 41542 11478 41560 11542
rect 41624 11478 42092 11542
rect 42156 11478 42174 11542
rect 41542 11460 42174 11478
rect 45742 11542 46318 11560
rect 45742 11478 45760 11542
rect 45824 11478 46236 11542
rect 46300 11478 46318 11542
rect 45742 11460 46318 11478
rect 41543 11455 41641 11460
rect 42074 11454 42174 11460
rect 45743 11455 45841 11460
rect 46218 11454 46318 11460
rect 39488 11411 39588 11412
rect 39483 11394 39593 11411
rect 39483 11330 39506 11394
rect 39570 11330 39593 11394
rect 43688 11393 43788 11394
rect 39483 11313 39593 11330
rect 40880 11356 40996 11386
rect 39488 11266 39588 11313
rect 40880 11300 40910 11356
rect 40966 11300 40996 11356
rect 40880 11270 40996 11300
rect 43683 11376 43793 11393
rect 43683 11312 43706 11376
rect 43770 11312 43793 11376
rect 43683 11295 43793 11312
rect 45045 11366 45163 11397
rect 45045 11310 45076 11366
rect 45132 11310 45163 11366
rect 39488 11154 39642 11266
rect 36925 10507 37733 10528
rect 36925 10363 36952 10507
rect 37096 10363 37733 10507
rect 36925 10342 37733 10363
rect 37131 8932 37733 10342
rect 39542 9306 39642 11154
rect 40885 10991 40991 11270
rect 43688 11154 43788 11295
rect 45045 11279 45163 11310
rect 45050 11168 45158 11279
rect 45008 11090 45158 11168
rect 45050 11088 45158 11090
rect 45010 11078 45158 11088
rect 45010 10952 45146 11078
rect 46399 10634 46992 12380
rect 46399 10510 46999 10634
rect 46399 10498 47166 10510
rect 46399 10354 47004 10498
rect 47148 10354 47166 10498
rect 46399 10342 47166 10354
rect 46399 9958 46999 10342
rect 42452 9306 42552 9832
rect 39004 9284 42552 9306
rect 39004 9228 39026 9284
rect 39082 9228 42552 9284
rect 39004 9206 42552 9228
rect 46399 9218 47037 9958
rect 46399 8932 46999 9218
rect 37131 8398 46999 8932
rect 37131 8330 38478 8398
rect 37131 8328 37731 8330
rect 38476 8174 38478 8330
rect 38702 8396 46999 8398
rect 38702 8328 40890 8396
rect 38702 8174 38704 8328
rect 40886 8312 40890 8328
rect 38476 8166 38704 8174
rect 40888 8172 40890 8312
rect 41114 8328 43234 8396
rect 41114 8172 41116 8328
rect 43230 8312 43234 8328
rect 40888 8164 41116 8172
rect 43232 8172 43234 8312
rect 43458 8330 45622 8396
rect 43458 8328 44542 8330
rect 43458 8172 43460 8328
rect 43232 8164 43460 8172
rect 45620 8172 45622 8330
rect 45846 8348 46999 8396
rect 45846 8330 46992 8348
rect 45846 8310 45850 8330
rect 45846 8172 45848 8310
rect 45620 8164 45848 8172
rect 36990 7720 47596 7738
rect 53050 7722 53150 7728
rect 36990 7656 37014 7720
rect 37078 7656 47596 7720
rect 36990 7638 47596 7656
rect 47496 7222 47596 7638
rect 49800 7704 53150 7722
rect 49800 7698 53068 7704
rect 49800 7642 49824 7698
rect 49880 7642 53068 7698
rect 49800 7640 53068 7642
rect 53132 7640 53150 7704
rect 49800 7622 53150 7640
rect 53050 7616 53150 7622
rect 47494 7196 62432 7222
rect 38428 7155 38610 7180
rect 38428 7078 38447 7155
rect 37150 7064 38447 7078
rect 37149 7011 38447 7064
rect 38591 7078 38610 7155
rect 40828 7155 41010 7180
rect 40828 7078 40847 7155
rect 38591 7011 40847 7078
rect 40991 7078 41010 7155
rect 43240 7155 43422 7180
rect 43240 7078 43259 7155
rect 40991 7011 43259 7078
rect 43403 7078 43422 7155
rect 45640 7155 45822 7180
rect 45640 7078 45659 7155
rect 43403 7011 45659 7078
rect 45803 7078 45822 7155
rect 47494 7140 62352 7196
rect 62408 7140 62432 7196
rect 47494 7122 62432 7140
rect 45803 7011 47017 7078
rect 37149 6464 47017 7011
rect 36453 6180 36563 6197
rect 36453 6116 36476 6180
rect 36540 6116 36563 6180
rect 36453 6099 36563 6116
rect 36458 6098 36558 6099
rect 37149 5066 37749 6464
rect 45911 6198 46021 6203
rect 39048 6180 46021 6198
rect 39048 6116 39072 6180
rect 39136 6176 46021 6180
rect 39136 6120 45938 6176
rect 45994 6120 46021 6176
rect 39136 6116 46021 6120
rect 39048 6098 46021 6116
rect 39368 5682 39468 6098
rect 42330 5794 42430 6098
rect 45911 6093 46021 6098
rect 37014 5034 37749 5066
rect 37014 4890 37052 5034
rect 37196 4890 37749 5034
rect 37014 4858 37749 4890
rect 37149 2926 37749 4858
rect 46417 5008 47017 6464
rect 48476 5981 48576 5982
rect 48471 5964 48581 5981
rect 48471 5900 48494 5964
rect 48558 5900 48581 5964
rect 48471 5883 48581 5900
rect 48476 5758 48576 5883
rect 48476 5734 49388 5758
rect 48476 5678 49308 5734
rect 49364 5678 49388 5734
rect 48476 5658 49388 5678
rect 53048 5604 53148 5610
rect 49924 5586 53148 5604
rect 49924 5585 53066 5586
rect 49924 5529 49942 5585
rect 49998 5529 53066 5585
rect 49924 5522 53066 5529
rect 53130 5522 53148 5586
rect 49924 5504 53148 5522
rect 53048 5498 53148 5504
rect 46417 4999 47216 5008
rect 46417 4855 47057 4999
rect 47201 4855 47216 4999
rect 46417 4846 47216 4855
rect 52183 4956 52281 4961
rect 52183 4938 66110 4956
rect 52183 4874 52200 4938
rect 52264 4934 66110 4938
rect 52264 4878 66028 4934
rect 66084 4878 66110 4934
rect 52264 4874 66110 4878
rect 52183 4856 66110 4874
rect 52183 4851 52281 4856
rect 38910 4077 39020 4204
rect 40278 4105 40378 4356
rect 38910 4021 38937 4077
rect 38993 4021 39020 4077
rect 38910 3994 39020 4021
rect 40273 4088 40383 4105
rect 40273 4024 40296 4088
rect 40360 4024 40383 4088
rect 40273 4007 40383 4024
rect 43082 4075 43192 4226
rect 44490 4089 44590 4350
rect 43082 4019 43109 4075
rect 43165 4019 43192 4075
rect 40278 4006 40378 4007
rect 43082 3992 43192 4019
rect 44485 4072 44595 4089
rect 44485 4008 44508 4072
rect 44572 4008 44595 4072
rect 44485 3991 44595 4008
rect 44490 3990 44590 3991
rect 41543 3960 41641 3965
rect 42074 3960 42174 3966
rect 45743 3960 45841 3965
rect 46238 3960 46338 3966
rect 41542 3942 42174 3960
rect 41542 3878 41560 3942
rect 41624 3878 42092 3942
rect 42156 3878 42174 3942
rect 41542 3860 42174 3878
rect 45742 3942 46338 3960
rect 45742 3878 45760 3942
rect 45824 3878 46256 3942
rect 46320 3878 46338 3942
rect 45742 3860 46338 3878
rect 41543 3855 41641 3860
rect 42074 3854 42174 3860
rect 45743 3855 45841 3860
rect 46238 3854 46338 3860
rect 39488 3797 39588 3798
rect 39483 3780 39593 3797
rect 39483 3716 39506 3780
rect 39570 3716 39593 3780
rect 39483 3699 39593 3716
rect 40780 3772 40900 3804
rect 43688 3799 43788 3800
rect 40780 3716 40812 3772
rect 40868 3716 40900 3772
rect 39488 3666 39588 3699
rect 40780 3684 40900 3716
rect 43683 3782 43793 3799
rect 43683 3718 43706 3782
rect 43770 3718 43793 3782
rect 43683 3701 43793 3718
rect 45056 3760 45176 3792
rect 45056 3704 45088 3760
rect 45144 3704 45176 3760
rect 39488 3554 39642 3666
rect 36943 2905 37749 2926
rect 36943 2761 36970 2905
rect 37114 2761 37749 2905
rect 36943 2740 37749 2761
rect -7176 1422 -7076 1916
rect -10086 1322 -7076 1422
rect -3207 1064 -2607 2202
rect 36054 1691 36154 2238
rect 36049 1674 36159 1691
rect -2334 1625 -2234 1626
rect -2339 1608 -2229 1625
rect -2339 1544 -2316 1608
rect -2252 1544 -2229 1608
rect 36049 1610 36072 1674
rect 36136 1610 36159 1674
rect 36049 1593 36159 1610
rect 36054 1592 36154 1593
rect -2339 1527 -2229 1544
rect -7140 1062 -2607 1064
rect -12475 505 -2607 1062
rect -12475 460 -11149 505
rect -11156 281 -11149 460
rect -10925 460 -8737 505
rect -10925 281 -10918 460
rect -11156 268 -10918 281
rect -8744 281 -8737 460
rect -8513 460 -6325 505
rect -8513 281 -8506 460
rect -8744 268 -8506 281
rect -6332 281 -6325 460
rect -6101 462 -3913 505
rect -6101 460 -5990 462
rect -3978 460 -3913 462
rect -6101 281 -6094 460
rect -6332 268 -6094 281
rect -3920 281 -3913 460
rect -3689 462 -2607 505
rect -2334 602 -2230 1527
rect 37149 1330 37749 2740
rect 39542 1692 39642 3554
rect 40785 3463 40895 3684
rect 43688 3554 43788 3701
rect 45056 3672 45176 3704
rect 45061 3381 45171 3672
rect 46417 2908 47017 4846
rect 48482 3756 48582 3762
rect 48482 3738 49378 3756
rect 48482 3674 48500 3738
rect 48564 3734 49378 3738
rect 48564 3678 49304 3734
rect 49360 3678 49378 3734
rect 48564 3674 49378 3678
rect 48482 3656 49378 3674
rect 48482 3650 48582 3656
rect 52181 3604 52283 3611
rect 50066 3586 52283 3604
rect 50066 3585 52200 3586
rect 50066 3529 50084 3585
rect 50140 3529 52200 3585
rect 50066 3522 52200 3529
rect 52264 3522 52283 3586
rect 50066 3504 52283 3522
rect 52181 3497 52283 3504
rect 61918 2916 62248 2938
rect 46417 2896 47184 2908
rect 46417 2752 47022 2896
rect 47166 2752 47184 2896
rect 61918 2860 62170 2916
rect 62226 2860 62248 2916
rect 46417 2740 47184 2752
rect 53051 2834 53149 2839
rect 61918 2838 62248 2860
rect 61918 2834 62018 2838
rect 53051 2816 62018 2834
rect 53051 2752 53068 2816
rect 53132 2752 62018 2816
rect 42452 1692 42552 2232
rect 39160 1674 46162 1692
rect 39160 1610 39184 1674
rect 39248 1668 46162 1674
rect 39248 1612 46090 1668
rect 46146 1612 46162 1668
rect 39248 1610 46162 1612
rect 39160 1592 46162 1610
rect 46417 1330 47017 2740
rect 53051 2734 62018 2752
rect 53051 2729 53149 2734
rect 52177 1672 52287 1678
rect 49806 1649 52287 1672
rect 49806 1644 52200 1649
rect 49806 1588 49830 1644
rect 49886 1588 52200 1644
rect 49806 1585 52200 1588
rect 52264 1585 52287 1649
rect 49806 1562 52287 1585
rect 52177 1556 52287 1562
rect 37149 796 47017 1330
rect 37149 728 38496 796
rect 37149 726 37749 728
rect -2334 580 8126 602
rect -2334 524 8044 580
rect 8100 524 8126 580
rect 38494 572 38496 728
rect 38720 794 47017 796
rect 38720 726 40908 794
rect 38720 572 38722 726
rect 40904 710 40908 726
rect 38494 564 38722 572
rect 40906 570 40908 710
rect 41132 726 43252 794
rect 41132 570 41134 726
rect 43248 710 43252 726
rect 40906 562 41134 570
rect 43250 570 43252 710
rect 43476 728 45640 794
rect 43476 726 44560 728
rect 43476 570 43478 726
rect 43250 562 43478 570
rect 45638 570 45640 728
rect 45864 746 47017 794
rect 45864 728 47016 746
rect 45864 708 45868 728
rect 45864 570 45866 708
rect 45638 562 45866 570
rect -2334 502 8126 524
rect -2334 500 -2234 502
rect -3689 460 -3578 462
rect -3689 281 -3682 460
rect -3920 268 -3682 281
<< via3 >>
rect -1416 27640 -1352 27647
rect -1416 27584 -1412 27640
rect -1412 27584 -1356 27640
rect -1356 27584 -1352 27640
rect -1416 27583 -1352 27584
rect 47831 27650 47895 27654
rect 47831 27594 47835 27650
rect 47835 27594 47891 27650
rect 47891 27594 47895 27650
rect 47831 27590 47895 27594
rect 47911 27650 47975 27654
rect 47911 27594 47915 27650
rect 47915 27594 47971 27650
rect 47971 27594 47975 27650
rect 47911 27590 47975 27594
rect 47991 27650 48055 27654
rect 47991 27594 47995 27650
rect 47995 27594 48051 27650
rect 48051 27594 48055 27650
rect 47991 27590 48055 27594
rect 48071 27650 48135 27654
rect 48071 27594 48075 27650
rect 48075 27594 48131 27650
rect 48131 27594 48135 27650
rect 48071 27590 48135 27594
rect 48151 27650 48215 27654
rect 48151 27594 48155 27650
rect 48155 27594 48211 27650
rect 48211 27594 48215 27650
rect 48151 27590 48215 27594
rect 48231 27650 48295 27654
rect 48231 27594 48235 27650
rect 48235 27594 48291 27650
rect 48291 27594 48295 27650
rect 48231 27590 48295 27594
rect 48311 27650 48375 27654
rect 48311 27594 48315 27650
rect 48315 27594 48371 27650
rect 48371 27594 48375 27650
rect 48311 27590 48375 27594
rect 48391 27650 48455 27654
rect 48391 27594 48395 27650
rect 48395 27594 48451 27650
rect 48451 27594 48455 27650
rect 48391 27590 48455 27594
rect 38432 26422 38576 26566
rect 41355 26417 41499 26561
rect 37084 24678 37148 24742
rect 36486 23488 36550 23552
rect 42948 24668 43012 24732
rect 46594 24452 46658 24516
rect 40420 23788 40484 23852
rect 41580 23630 41644 23694
rect 42048 23630 42112 23694
rect 39510 23486 39574 23550
rect 37104 22584 37168 22648
rect 42902 22556 42966 22620
rect 49778 21618 49842 21682
rect 46422 21300 46486 21364
rect 52162 23632 52226 23696
rect 51812 20984 51876 21048
rect 36490 19844 36554 19908
rect 38511 20329 38655 20473
rect 40911 20329 41055 20473
rect 43311 20329 43455 20473
rect 45437 20329 45581 20473
rect 47611 20329 47755 20473
rect 50011 20329 50155 20473
rect 39096 19844 39160 19908
rect 37182 18614 37326 18758
rect -13454 10650 -13390 10714
rect -11153 14023 -11009 14167
rect -8813 14007 -8669 14151
rect -6330 13990 -6186 14134
rect -3933 14017 -3789 14161
rect -13090 13056 -13026 13120
rect -10556 13056 -10492 13120
rect -12609 11895 -12545 11959
rect -2378 12822 -2314 12886
rect -2510 11778 -2446 11842
rect -9208 10948 -9144 11012
rect -5252 10948 -5188 11012
rect -8084 10800 -8020 10864
rect -7552 10800 -7488 10864
rect -3884 10798 -3820 10862
rect -3374 10798 -3310 10862
rect -10338 10650 -10274 10714
rect -12626 9938 -12562 10002
rect -13082 8538 -13018 8602
rect -13286 3456 -13222 3520
rect -6538 10652 -6474 10716
rect -2497 9763 -2433 9827
rect -10516 8538 -10452 8602
rect 36272 15294 36336 15358
rect 36272 9460 36336 9524
rect -1738 8782 -1674 8846
rect -11189 7414 -10965 7638
rect -8777 7414 -8553 7638
rect -6365 7414 -6141 7638
rect -3953 7414 -3729 7638
rect 35246 7656 35310 7720
rect -11189 6823 -10965 7047
rect -8777 6823 -8553 7047
rect -6365 6823 -6141 7047
rect -3953 6823 -3729 7047
rect -12714 5584 -12650 5648
rect -12583 4619 -12439 4763
rect -2404 5584 -2340 5648
rect -2655 4567 -2511 4711
rect -9348 3746 -9284 3810
rect -5118 3750 -5054 3814
rect -8068 3600 -8004 3664
rect -7536 3600 -7472 3664
rect -3868 3602 -3804 3666
rect -3364 3602 -3300 3666
rect -10150 3456 -10086 3520
rect -5882 3452 -5818 3516
rect -12549 2555 -12485 2619
rect -13080 1546 -13016 1610
rect -2658 2512 -2514 2656
rect 51347 18579 51491 18723
rect 40434 17748 40498 17812
rect 44660 17736 44724 17800
rect 48782 17746 48846 17810
rect 41690 17596 41754 17660
rect 42222 17596 42286 17660
rect 45890 17596 45954 17660
rect 46422 17596 46486 17660
rect 50090 17596 50154 17660
rect 50622 17596 50686 17660
rect 39636 17442 39700 17506
rect 43836 17442 43900 17506
rect 37100 16485 37244 16629
rect 48036 17440 48100 17504
rect 51376 16482 51520 16626
rect 39316 15294 39380 15358
rect 52398 15018 52462 15082
rect 36766 13500 36830 13564
rect 38485 14165 38629 14309
rect 40897 14165 41041 14309
rect 43297 14165 43441 14309
rect 45697 14165 45841 14309
rect 37034 12492 37178 12636
rect 47697 14165 47841 14309
rect 50097 14165 50241 14309
rect 47039 12457 47183 12601
rect 40310 11628 40374 11692
rect 44530 11628 44594 11692
rect 41560 11478 41624 11542
rect 42092 11478 42156 11542
rect 45760 11478 45824 11542
rect 46236 11478 46300 11542
rect 39506 11330 39570 11394
rect 43706 11312 43770 11376
rect 36952 10363 37096 10507
rect 47004 10354 47148 10498
rect 38478 8174 38702 8398
rect 40890 8172 41114 8396
rect 43234 8172 43458 8396
rect 45622 8172 45846 8396
rect 37014 7656 37078 7720
rect 53068 7640 53132 7704
rect 38447 7011 38591 7155
rect 40847 7011 40991 7155
rect 43259 7011 43403 7155
rect 45659 7011 45803 7155
rect 36476 6116 36540 6180
rect 39072 6116 39136 6180
rect 37052 4890 37196 5034
rect 48494 5900 48558 5964
rect 53066 5522 53130 5586
rect 47057 4855 47201 4999
rect 52200 4874 52264 4938
rect 40296 4024 40360 4088
rect 44508 4008 44572 4072
rect 41560 3878 41624 3942
rect 42092 3878 42156 3942
rect 45760 3878 45824 3942
rect 46256 3878 46320 3942
rect 39506 3716 39570 3780
rect 43706 3718 43770 3782
rect 36970 2761 37114 2905
rect -2316 1544 -2252 1608
rect 36072 1610 36136 1674
rect -11149 281 -10925 505
rect -8737 281 -8513 505
rect -6325 281 -6101 505
rect -3913 281 -3689 505
rect 48500 3674 48564 3738
rect 52200 3522 52264 3586
rect 47022 2752 47166 2896
rect 53068 2752 53132 2816
rect 39184 1610 39248 1674
rect 52200 1585 52264 1649
rect 38496 572 38720 796
rect 40908 570 41132 794
rect 43252 570 43476 794
rect 45640 570 45864 794
<< metal4 >>
rect 33530 27654 55572 28340
rect -1420 27647 -1348 27648
rect -1420 27583 -1416 27647
rect -1352 27583 -1348 27647
rect -1420 27582 -1348 27583
rect 33530 27590 47831 27654
rect 47895 27590 47911 27654
rect 47975 27590 47991 27654
rect 48055 27590 48071 27654
rect 48135 27590 48151 27654
rect 48215 27590 48231 27654
rect 48295 27590 48311 27654
rect 48375 27590 48391 27654
rect 48455 27590 55572 27654
rect 33530 27540 55572 27590
rect 38429 26566 38579 26569
rect 38429 26422 38432 26566
rect 38576 26422 38579 26566
rect 38429 26419 38579 26422
rect 41347 26561 41507 26569
rect 38430 26166 38578 26419
rect 41347 26417 41355 26561
rect 41499 26417 41507 26561
rect 41347 26409 41507 26417
rect 41348 26105 41506 26409
rect 39530 25634 46676 25734
rect 39530 25280 39630 25634
rect 37049 24776 37183 24777
rect 37049 24742 37586 24776
rect 37049 24678 37084 24742
rect 37148 24678 37586 24742
rect 37049 24644 37586 24678
rect 37049 24643 37183 24644
rect 41418 24614 41928 24714
rect 40401 23852 40503 23871
rect 40401 23788 40420 23852
rect 40484 23788 40503 23852
rect 36467 23568 36569 23571
rect 40401 23568 40503 23788
rect 36462 23552 40503 23568
rect 36462 23488 36486 23552
rect 36550 23550 40503 23552
rect 36550 23488 39510 23550
rect 36462 23486 39510 23488
rect 39574 23486 40503 23550
rect 36462 23468 40503 23486
rect 40401 23467 40503 23468
rect 41562 23694 41662 23712
rect 41562 23630 41580 23694
rect 41644 23630 41662 23694
rect 41562 23212 41662 23630
rect 37075 22676 37197 22677
rect 37075 22648 37492 22676
rect 37075 22584 37104 22648
rect 37168 22584 37492 22648
rect 37075 22556 37492 22584
rect 37075 22555 37197 22556
rect 39512 21694 39612 22074
rect 41828 21694 41928 24614
rect 42030 23714 42130 25634
rect 42911 24768 43049 24769
rect 42584 24732 43049 24768
rect 42584 24668 42948 24732
rect 43012 24668 43049 24732
rect 42584 24632 43049 24668
rect 42911 24631 43049 24632
rect 46576 24535 46676 25634
rect 46575 24516 46677 24535
rect 46575 24452 46594 24516
rect 46658 24452 46677 24516
rect 46575 24433 46677 24452
rect 52143 23714 52245 23715
rect 42030 23713 52245 23714
rect 42029 23696 52245 23713
rect 42029 23694 52162 23696
rect 42029 23630 42048 23694
rect 42112 23632 52162 23694
rect 52226 23632 52245 23696
rect 42112 23630 52245 23632
rect 42029 23614 52245 23630
rect 42029 23611 42131 23614
rect 52143 23613 52245 23614
rect 42863 22658 43005 22659
rect 42582 22620 43005 22658
rect 42582 22556 42902 22620
rect 42966 22556 43005 22620
rect 42582 22518 43005 22556
rect 42863 22517 43005 22518
rect 49759 21694 49861 21701
rect 52380 21694 52480 21696
rect 39512 21682 52480 21694
rect 39512 21618 49778 21682
rect 49842 21618 52480 21682
rect 39512 21594 52480 21618
rect 46404 21364 46504 21382
rect 46404 21300 46422 21364
rect 46486 21300 46504 21364
rect 38494 20491 38672 20787
rect 40894 20491 41072 20787
rect 43294 20491 43472 20787
rect 45420 20491 45598 20787
rect 38493 20473 38673 20491
rect 38493 20329 38511 20473
rect 38655 20329 38673 20473
rect 38493 20311 38673 20329
rect 40893 20473 41073 20491
rect 40893 20329 40911 20473
rect 41055 20329 41073 20473
rect 40893 20311 41073 20329
rect 43293 20473 43473 20491
rect 43293 20329 43311 20473
rect 43455 20329 43473 20473
rect 43293 20311 43473 20329
rect 45419 20473 45599 20491
rect 45419 20329 45437 20473
rect 45581 20329 45599 20473
rect 45419 20311 45599 20329
rect 39077 19926 39179 19927
rect 36472 19908 39179 19926
rect 36472 19844 36490 19908
rect 36554 19844 39096 19908
rect 39160 19844 39179 19908
rect 36472 19826 39179 19844
rect 39077 19825 39179 19826
rect 46404 19700 46504 21300
rect 51793 21066 51895 21067
rect 51793 21048 52248 21066
rect 51793 20984 51812 21048
rect 51876 20984 52248 21048
rect 51793 20966 52248 20984
rect 51793 20965 51895 20966
rect 47594 20491 47772 20787
rect 49994 20491 50172 20787
rect 47593 20473 47773 20491
rect 47593 20329 47611 20473
rect 47755 20329 47773 20473
rect 47593 20311 47773 20329
rect 49993 20473 50173 20491
rect 49993 20329 50011 20473
rect 50155 20329 50173 20473
rect 49993 20311 50173 20329
rect 39640 19600 50704 19700
rect 39640 19246 39740 19600
rect 37149 18790 37359 18791
rect 37149 18758 37676 18790
rect 37149 18614 37182 18758
rect 37326 18614 37676 18758
rect 37149 18582 37676 18614
rect 37149 18581 37359 18582
rect 41528 18580 42068 18680
rect 40416 17812 40516 17830
rect 40416 17748 40434 17812
rect 40498 17748 40516 17812
rect 40416 17524 40516 17748
rect 39618 17506 40516 17524
rect 39618 17442 39636 17506
rect 39700 17442 40516 17506
rect 39618 17424 40516 17442
rect 41672 17660 41772 17678
rect 41672 17596 41690 17660
rect 41754 17596 41772 17660
rect 41672 17178 41772 17596
rect 37078 16650 37266 16651
rect 37078 16629 37629 16650
rect 37078 16485 37100 16629
rect 37244 16485 37629 16629
rect 37078 16464 37629 16485
rect 37078 16463 37266 16464
rect 39622 15660 39722 16040
rect 41968 15660 42068 18580
rect 42204 17679 42304 19600
rect 43840 19246 43940 19600
rect 45728 18580 46268 18680
rect 44642 17800 44742 17818
rect 44642 17736 44660 17800
rect 44724 17736 44742 17800
rect 42203 17660 42305 17679
rect 42203 17596 42222 17660
rect 42286 17596 42305 17660
rect 42203 17577 42305 17596
rect 44642 17524 44742 17736
rect 43818 17506 44742 17524
rect 43818 17442 43836 17506
rect 43900 17442 44742 17506
rect 43818 17424 44742 17442
rect 45872 17660 45972 17678
rect 45872 17596 45890 17660
rect 45954 17596 45972 17660
rect 45872 17178 45972 17596
rect 43822 15660 43922 16040
rect 46168 15660 46268 18580
rect 46404 17679 46504 19600
rect 48040 19246 48140 19600
rect 49928 18580 50468 18680
rect 48764 17810 48864 17828
rect 48764 17746 48782 17810
rect 48846 17746 48864 17810
rect 46403 17660 46505 17679
rect 46403 17596 46422 17660
rect 46486 17596 46505 17660
rect 46403 17577 46505 17596
rect 48764 17522 48864 17746
rect 48018 17504 48864 17522
rect 48018 17440 48036 17504
rect 48100 17440 48864 17504
rect 48018 17422 48864 17440
rect 50072 17660 50172 17678
rect 50072 17596 50090 17660
rect 50154 17596 50172 17660
rect 50072 17178 50172 17596
rect 48022 15660 48122 16040
rect 50368 15660 50468 18580
rect 50604 17679 50704 19600
rect 51337 18732 51501 18733
rect 51037 18723 51501 18732
rect 51037 18579 51347 18723
rect 51491 18579 51501 18723
rect 51037 18570 51501 18579
rect 51337 18569 51501 18570
rect 50603 17660 50705 17679
rect 50603 17596 50622 17660
rect 50686 17596 50705 17660
rect 50603 17577 50705 17596
rect 51363 16638 51533 16639
rect 51014 16626 51533 16638
rect 51014 16482 51376 16626
rect 51520 16482 51533 16626
rect 51014 16470 51533 16482
rect 51363 16469 51533 16470
rect 52148 15660 52248 20966
rect 39622 15560 52248 15660
rect 39297 15376 39399 15377
rect 36254 15358 39399 15376
rect 36254 15294 36272 15358
rect 36336 15294 39316 15358
rect 39380 15294 39399 15358
rect 36254 15276 39399 15294
rect 39297 15275 39399 15276
rect 52380 15101 52480 21594
rect 52379 15082 52481 15101
rect 52379 15018 52398 15082
rect 52462 15018 52481 15082
rect 52379 14999 52481 15018
rect 38478 14317 38636 14613
rect 40890 14317 41048 14613
rect 43290 14317 43448 14613
rect 45690 14317 45848 14613
rect 47690 14317 47848 14613
rect 50090 14317 50248 14613
rect 38477 14309 38637 14317
rect -11155 14167 -11007 14169
rect -11155 14023 -11153 14167
rect -11009 14023 -11007 14167
rect -11155 14021 -11007 14023
rect -8837 14151 -8645 14175
rect -3941 14161 -3781 14169
rect -11154 13679 -11008 14021
rect -8837 14007 -8813 14151
rect -8669 14007 -8645 14151
rect -8837 13983 -8645 14007
rect -6347 14134 -6169 14151
rect -6347 13990 -6330 14134
rect -6186 13990 -6169 14134
rect -3941 14017 -3933 14161
rect -3789 14017 -3781 14161
rect 38477 14165 38485 14309
rect 38629 14165 38637 14309
rect 38477 14157 38637 14165
rect 40889 14309 41049 14317
rect 40889 14165 40897 14309
rect 41041 14165 41049 14309
rect 40889 14157 41049 14165
rect 43289 14309 43449 14317
rect 43289 14165 43297 14309
rect 43441 14165 43449 14309
rect 43289 14157 43449 14165
rect 45689 14309 45849 14317
rect 45689 14165 45697 14309
rect 45841 14165 45849 14309
rect 45689 14157 45849 14165
rect 47689 14309 47849 14317
rect 47689 14165 47697 14309
rect 47841 14165 47849 14309
rect 47689 14157 47849 14165
rect 50089 14309 50249 14317
rect 50089 14165 50097 14309
rect 50241 14165 50249 14309
rect 50089 14157 50249 14165
rect -3941 14009 -3781 14017
rect -8836 13619 -8646 13983
rect -6347 13973 -6169 13990
rect -6346 13602 -6170 13973
rect -3940 13667 -3782 14009
rect 36748 13564 46318 13582
rect 36748 13500 36766 13564
rect 36830 13500 46318 13564
rect 36748 13482 46318 13500
rect -10575 13138 -10473 13139
rect -13108 13120 -10473 13138
rect 39510 13128 39610 13482
rect -13108 13056 -13090 13120
rect -13026 13056 -10556 13120
rect -10492 13056 -10473 13120
rect -13108 13038 -10473 13056
rect -10575 13037 -10473 13038
rect -2397 12904 -2295 12905
rect -10164 12886 -2295 12904
rect -10164 12822 -2378 12886
rect -2314 12822 -2295 12886
rect -10164 12804 -2295 12822
rect -10164 12450 -10064 12804
rect -12625 11974 -12529 11975
rect -12625 11959 -12207 11974
rect -12625 11895 -12609 11959
rect -12545 11895 -12207 11959
rect -12625 11880 -12207 11895
rect -12625 11879 -12529 11880
rect -8246 11784 -7706 11884
rect -9226 11012 -9126 11030
rect -9226 10948 -9208 11012
rect -9144 10948 -9126 11012
rect -9226 10732 -9126 10948
rect -13472 10714 -9126 10732
rect -13472 10650 -13454 10714
rect -13390 10650 -10338 10714
rect -10274 10650 -9126 10714
rect -13472 10632 -9126 10650
rect -8102 10864 -8002 10882
rect -8102 10800 -8084 10864
rect -8020 10800 -8002 10864
rect -8102 10382 -8002 10800
rect -12635 10010 -12553 10011
rect -12635 10002 -12204 10010
rect -12635 9938 -12626 10002
rect -12562 9938 -12204 10002
rect -12635 9930 -12204 9938
rect -12635 9929 -12553 9930
rect -10182 8864 -10082 9244
rect -7806 8864 -7706 11784
rect -7570 10883 -7470 12804
rect -5934 12450 -5834 12804
rect -4046 11784 -3506 11884
rect -5270 11012 -5170 11030
rect -5270 10948 -5252 11012
rect -5188 10948 -5170 11012
rect -7571 10864 -7469 10883
rect -7571 10800 -7552 10864
rect -7488 10800 -7469 10864
rect -7571 10781 -7469 10800
rect -5270 10734 -5170 10948
rect -6556 10716 -5170 10734
rect -6556 10652 -6538 10716
rect -6474 10652 -5170 10716
rect -6556 10634 -5170 10652
rect -3902 10862 -3802 10880
rect -3902 10798 -3884 10862
rect -3820 10798 -3802 10862
rect -3902 10382 -3802 10798
rect -5952 8864 -5852 9244
rect -3606 8864 -3506 11784
rect -3392 10881 -3292 12804
rect -2397 12803 -2295 12804
rect 37001 12668 37211 12669
rect 37001 12636 37528 12668
rect 37001 12492 37034 12636
rect 37178 12492 37528 12636
rect 37001 12460 37528 12492
rect 41398 12462 41938 12562
rect 37001 12459 37211 12460
rect -2525 11856 -2431 11857
rect -2892 11842 -2431 11856
rect -2892 11778 -2510 11842
rect -2446 11778 -2431 11842
rect -2892 11764 -2431 11778
rect -2525 11763 -2431 11764
rect 40292 11692 40392 11710
rect 40292 11628 40310 11692
rect 40374 11628 40392 11692
rect 40292 11412 40392 11628
rect 39488 11394 40392 11412
rect 39488 11330 39506 11394
rect 39570 11330 40392 11394
rect 39488 11312 40392 11330
rect 41542 11542 41642 11560
rect 41542 11478 41560 11542
rect 41624 11478 41642 11542
rect 41542 11060 41642 11478
rect -3393 10862 -3291 10881
rect -3393 10798 -3374 10862
rect -3310 10798 -3291 10862
rect -3393 10779 -3291 10798
rect -3392 10776 -3292 10779
rect 36930 10528 37118 10529
rect 36930 10507 37481 10528
rect 36930 10363 36952 10507
rect 37096 10363 37481 10507
rect 36930 10342 37481 10363
rect 36930 10341 37118 10342
rect -2519 9848 -2411 9849
rect -2891 9827 -2411 9848
rect -2891 9763 -2497 9827
rect -2433 9763 -2411 9827
rect -2891 9742 -2411 9763
rect -2519 9741 -2411 9742
rect 39492 9542 39592 9922
rect 41838 9542 41938 12462
rect 42074 11561 42174 13482
rect 43710 13128 43810 13482
rect 45598 12462 46138 12562
rect 44512 11692 44612 11710
rect 44512 11628 44530 11692
rect 44594 11628 44612 11692
rect 42073 11542 42175 11561
rect 42073 11478 42092 11542
rect 42156 11478 42175 11542
rect 42073 11459 42175 11478
rect 44512 11394 44612 11628
rect 43688 11376 44612 11394
rect 43688 11312 43706 11376
rect 43770 11312 44612 11376
rect 43688 11294 44612 11312
rect 45742 11542 45842 11560
rect 45742 11478 45760 11542
rect 45824 11478 45842 11542
rect 45742 11060 45842 11478
rect 43692 9542 43792 9922
rect 46038 9542 46138 12462
rect 46218 11561 46318 13482
rect 47029 12610 47193 12611
rect 46679 12601 47193 12610
rect 46679 12457 47039 12601
rect 47183 12457 47193 12601
rect 46679 12448 47193 12457
rect 47029 12447 47193 12448
rect 46217 11556 46319 11561
rect 46217 11542 53150 11556
rect 46217 11478 46236 11542
rect 46300 11478 53150 11542
rect 46217 11459 53150 11478
rect 46218 11456 53150 11459
rect 46991 10510 47161 10511
rect 46658 10498 47161 10510
rect 46658 10354 47004 10498
rect 47148 10354 47161 10498
rect 46658 10342 47161 10354
rect 46991 10341 47161 10342
rect 36254 9524 52282 9542
rect 36254 9460 36272 9524
rect 36336 9460 52282 9524
rect 36254 9442 52282 9460
rect -10182 8846 -1656 8864
rect -10182 8782 -1738 8846
rect -1674 8782 -1656 8846
rect -10182 8764 -1656 8782
rect 38476 8638 38704 8726
rect -10535 8620 -10433 8621
rect -13100 8602 -10433 8620
rect -13100 8538 -13082 8602
rect -13018 8538 -10516 8602
rect -10452 8538 -10433 8602
rect -13100 8520 -10433 8538
rect -10535 8519 -10433 8520
rect 38394 8398 38748 8638
rect 40888 8600 41116 8726
rect 38394 8174 38478 8398
rect 38702 8174 38748 8398
rect -11198 7638 -10956 8059
rect -11198 7414 -11189 7638
rect -10965 7414 -10956 7638
rect -11198 7057 -10956 7414
rect -8786 7638 -8544 8059
rect -8786 7414 -8777 7638
rect -8553 7414 -8544 7638
rect -8786 7057 -8544 7414
rect -6374 7638 -6132 8059
rect -6374 7414 -6365 7638
rect -6141 7414 -6132 7638
rect -6374 7057 -6132 7414
rect -3962 7638 -3720 8059
rect 36995 7738 37097 7739
rect 35228 7720 37097 7738
rect 35228 7656 35246 7720
rect 35310 7656 37014 7720
rect 37078 7656 37097 7720
rect 35228 7638 37097 7656
rect -3962 7414 -3953 7638
rect -3729 7414 -3720 7638
rect 36995 7637 37097 7638
rect -3962 7057 -3720 7414
rect 38394 7155 38748 8174
rect -11199 7047 -10955 7057
rect -11199 6823 -11189 7047
rect -10965 6823 -10955 7047
rect -11199 6813 -10955 6823
rect -8787 7047 -8543 7057
rect -8787 6823 -8777 7047
rect -8553 6823 -8543 7047
rect -8787 6813 -8543 6823
rect -6375 7047 -6131 7057
rect -6375 6823 -6365 7047
rect -6141 6823 -6131 7047
rect -6375 6813 -6131 6823
rect -3963 7047 -3719 7057
rect -3963 6823 -3953 7047
rect -3729 6823 -3719 7047
rect -3963 6813 -3719 6823
rect 38394 7011 38447 7155
rect 38591 7011 38748 7155
rect -11198 6413 -10956 6813
rect -9421 6658 -9070 6659
rect -9421 6338 -9420 6658
rect -8786 6413 -8544 6813
rect -6374 6413 -6132 6813
rect -3962 6413 -3720 6813
rect 38394 6640 38748 7011
rect 40796 8396 41150 8600
rect 40796 8172 40890 8396
rect 41114 8172 41150 8396
rect 40796 7155 41150 8172
rect 40796 7011 40847 7155
rect 40991 7011 41150 7155
rect 38428 6635 38610 6640
rect 40796 6630 41150 7011
rect 43168 8396 43504 8730
rect 43168 8172 43234 8396
rect 43458 8172 43504 8396
rect 43168 7155 43504 8172
rect 43168 7011 43259 7155
rect 43403 7011 43504 7155
rect 43168 6620 43504 7011
rect 45576 8396 45872 8746
rect 45576 8172 45622 8396
rect 45846 8172 45872 8396
rect 45576 7155 45872 8172
rect 45576 7011 45659 7155
rect 45803 7011 45872 7155
rect 45576 6630 45872 7011
rect -9421 6337 -9070 6338
rect 39053 6198 39155 6199
rect 36458 6180 39155 6198
rect 36458 6116 36476 6180
rect 36540 6116 39072 6180
rect 39136 6116 39155 6180
rect 36458 6098 39155 6116
rect 39053 6097 39155 6098
rect 39510 5964 48576 5982
rect 39510 5900 48494 5964
rect 48558 5900 48576 5964
rect 39510 5882 48576 5900
rect -12732 5648 -2322 5666
rect -12732 5584 -12714 5648
rect -12650 5584 -2404 5648
rect -2340 5584 -2322 5648
rect -12732 5566 -2322 5584
rect -10118 5212 -10018 5566
rect -12587 4766 -12435 4767
rect -12587 4763 -12157 4766
rect -12587 4619 -12583 4763
rect -12439 4619 -12157 4763
rect -12587 4616 -12157 4619
rect -12587 4615 -12435 4616
rect -8230 4546 -7690 4646
rect -9366 3810 -9266 3828
rect -9366 3746 -9348 3810
rect -9284 3746 -9266 3810
rect -9366 3538 -9266 3746
rect -13304 3520 -9266 3538
rect -13304 3456 -13286 3520
rect -13222 3456 -10150 3520
rect -10086 3456 -9266 3520
rect -13304 3438 -9266 3456
rect -8086 3664 -7986 3682
rect -8086 3600 -8068 3664
rect -8004 3600 -7986 3664
rect -8086 3144 -7986 3600
rect -12581 2650 -12453 2651
rect -12581 2619 -12079 2650
rect -12581 2555 -12549 2619
rect -12485 2555 -12079 2619
rect -12581 2524 -12079 2555
rect -12581 2523 -12453 2524
rect -10136 1628 -10036 2006
rect -13098 1626 -9512 1628
rect -7790 1626 -7690 4546
rect -7554 3683 -7454 5566
rect -5918 5212 -5818 5566
rect -4030 4546 -3490 4646
rect -5144 3814 -5028 3840
rect -5144 3750 -5118 3814
rect -5054 3750 -5028 3814
rect -7555 3664 -7453 3683
rect -7555 3600 -7536 3664
rect -7472 3600 -7453 3664
rect -7555 3581 -7453 3600
rect -5909 3542 -5791 3543
rect -5144 3542 -5028 3750
rect -5909 3516 -5028 3542
rect -5909 3452 -5882 3516
rect -5818 3452 -5028 3516
rect -5909 3426 -5028 3452
rect -3886 3666 -3786 3684
rect -3886 3602 -3868 3666
rect -3804 3602 -3786 3666
rect -5909 3425 -5791 3426
rect -3886 3144 -3786 3602
rect -5936 1626 -5836 2006
rect -3590 1626 -3490 4546
rect -3382 3685 -3282 5566
rect 39510 5528 39610 5882
rect 37019 5066 37229 5067
rect 37019 5034 37546 5066
rect 37019 4890 37052 5034
rect 37196 4890 37546 5034
rect 37019 4858 37546 4890
rect 41398 4862 41938 4962
rect 37019 4857 37229 4858
rect -2661 4716 -2505 4717
rect -2943 4711 -2505 4716
rect -2943 4567 -2655 4711
rect -2511 4567 -2505 4711
rect -2943 4562 -2505 4567
rect -2661 4561 -2505 4562
rect 40278 4088 40378 4106
rect 40278 4024 40296 4088
rect 40360 4024 40378 4088
rect 40278 3798 40378 4024
rect 39488 3780 40378 3798
rect 39488 3716 39506 3780
rect 39570 3716 40378 3780
rect 39488 3698 40378 3716
rect 41542 3942 41642 3960
rect 41542 3878 41560 3942
rect 41624 3878 41642 3942
rect -3383 3666 -3281 3685
rect -3383 3602 -3364 3666
rect -3300 3602 -3281 3666
rect -3383 3583 -3281 3602
rect 41542 3460 41642 3878
rect 36948 2926 37136 2927
rect 36948 2905 37499 2926
rect 36948 2761 36970 2905
rect 37114 2761 37499 2905
rect 36948 2740 37499 2761
rect 36948 2739 37136 2740
rect -2667 2664 -2505 2665
rect -2926 2656 -2505 2664
rect -2926 2512 -2658 2656
rect -2514 2512 -2505 2656
rect -2926 2504 -2505 2512
rect -2667 2503 -2505 2504
rect 39492 1942 39592 2322
rect 41838 1942 41938 4862
rect 42074 3961 42174 5882
rect 43710 5528 43810 5882
rect 45598 4862 46138 4962
rect 44490 4072 44590 4090
rect 44490 4008 44508 4072
rect 44572 4008 44590 4072
rect 42073 3942 42175 3961
rect 42073 3878 42092 3942
rect 42156 3878 42175 3942
rect 42073 3859 42175 3878
rect 44490 3800 44590 4008
rect 43688 3782 44590 3800
rect 43688 3718 43706 3782
rect 43770 3718 44590 3782
rect 43688 3700 44590 3718
rect 45742 3942 45842 3960
rect 45742 3878 45760 3942
rect 45824 3878 45842 3942
rect 45742 3460 45842 3878
rect 43692 1942 43792 2322
rect 46038 1942 46138 4862
rect 46238 3961 46338 5882
rect 47047 5008 47211 5009
rect 46697 4999 47211 5008
rect 46697 4855 47057 4999
rect 47201 4855 47211 4999
rect 46697 4846 47211 4855
rect 47047 4845 47211 4846
rect 52182 4938 52282 9442
rect 53050 7723 53150 11456
rect 53049 7704 53151 7723
rect 53049 7640 53068 7704
rect 53132 7640 53151 7704
rect 53049 7621 53151 7640
rect 53050 5605 53150 7621
rect 53047 5586 53150 5605
rect 53047 5522 53066 5586
rect 53130 5522 53150 5586
rect 53047 5503 53150 5522
rect 52182 4874 52200 4938
rect 52264 4874 52282 4938
rect 52182 4087 52282 4874
rect 46237 3942 46339 3961
rect 46237 3878 46256 3942
rect 46320 3878 46339 3942
rect 46237 3859 46339 3878
rect 48481 3738 48583 3757
rect 48481 3674 48500 3738
rect 48564 3674 48583 3738
rect 48481 3655 48583 3674
rect 47009 2908 47179 2909
rect 46676 2896 47179 2908
rect 46676 2752 47022 2896
rect 47166 2752 47179 2896
rect 46676 2740 47179 2752
rect 47009 2739 47179 2740
rect 48482 1942 48582 3655
rect 52181 3606 52283 4087
rect 52180 3586 52284 3606
rect 52180 3522 52200 3586
rect 52264 3522 52284 3586
rect 52180 3502 52284 3522
rect 39492 1842 48582 1942
rect 52181 1897 52283 3502
rect 53050 2816 53150 5503
rect 53050 2752 53068 2816
rect 53132 2752 53150 2816
rect 53050 2734 53150 2752
rect 39165 1692 39267 1693
rect 36054 1674 39267 1692
rect -13098 1610 -2234 1626
rect -13098 1546 -13080 1610
rect -13016 1608 -2234 1610
rect -13016 1546 -2316 1608
rect -13098 1544 -2316 1546
rect -2252 1544 -2234 1608
rect 36054 1610 36072 1674
rect 36136 1610 39184 1674
rect 39248 1610 39267 1674
rect 52177 1673 52287 1897
rect 36054 1592 39267 1610
rect 39165 1591 39267 1592
rect 52176 1649 52288 1673
rect 52176 1585 52200 1649
rect 52264 1585 52288 1649
rect 52176 1561 52288 1585
rect -13098 1528 -2234 1544
rect -10136 1526 -2234 1528
rect -11156 513 -10918 859
rect -8744 513 -8506 859
rect -6332 513 -6094 859
rect -3920 513 -3682 859
rect 38494 799 38722 1124
rect 38493 796 38723 799
rect 40906 797 41134 1124
rect 43250 797 43478 1124
rect 45638 797 45866 1124
rect 38493 572 38496 796
rect 38720 572 38723 796
rect 38493 569 38723 572
rect 40905 794 41135 797
rect 40905 570 40908 794
rect 41132 570 41135 794
rect -11157 505 -10917 513
rect -11157 281 -11149 505
rect -10925 281 -10917 505
rect -11157 273 -10917 281
rect -8745 505 -8505 513
rect -8745 281 -8737 505
rect -8513 281 -8505 505
rect -8745 273 -8505 281
rect -6333 505 -6093 513
rect -6333 281 -6325 505
rect -6101 281 -6093 505
rect -6333 273 -6093 281
rect -3921 505 -3681 513
rect -3921 281 -3913 505
rect -3689 281 -3681 505
rect -3921 273 -3681 281
rect -11156 140 -10918 273
rect -8744 140 -8506 273
rect -6332 140 -6094 273
rect -3920 140 -3682 273
rect 38494 140 38722 569
rect 40905 567 41135 570
rect 43249 794 43479 797
rect 43249 570 43252 794
rect 43476 570 43479 794
rect 43249 567 43479 570
rect 45637 794 45867 797
rect 45637 570 45640 794
rect 45864 570 45867 794
rect 45637 567 45867 570
rect 40906 140 41134 567
rect 43250 140 43478 567
rect 45638 140 45866 567
rect -13292 -660 378 140
rect 34882 -660 90192 140
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_21
timestamp 1626486988
transform 1 0 -8610 0 1 762
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_46
timestamp 1626486988
transform 1 0 -10678 0 1 2584
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_47
timestamp 1626486988
transform 1 0 -8648 0 1 2584
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_23
timestamp 1626486988
transform 1 0 -12124 0 1 2580
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_19
timestamp 1626486988
transform -1 0 -11093 0 1 762
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_20
timestamp 1626486988
transform -1 0 -6322 0 1 764
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_45
timestamp 1626486988
transform 1 0 -6488 0 1 2584
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_44
timestamp 1626486988
transform 1 0 -4448 0 1 2584
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_22
timestamp 1626486988
transform -1 0 -2958 0 1 2582
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_18
timestamp 1626486988
transform 1 0 -3839 0 1 764
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_19
timestamp 1626486988
transform 1 0 -8610 0 1 6498
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_42
timestamp 1626486988
transform 1 0 -10678 0 1 4684
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_43
timestamp 1626486988
transform 1 0 -8648 0 1 4684
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_21
timestamp 1626486988
transform 1 0 -12124 0 1 4684
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_17
timestamp 1626486988
transform -1 0 -11093 0 1 6498
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_18
timestamp 1626486988
transform -1 0 -6322 0 1 6500
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_41
timestamp 1626486988
transform 1 0 -6488 0 1 4684
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_40
timestamp 1626486988
transform 1 0 -4448 0 1 4684
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_20
timestamp 1626486988
transform -1 0 -2958 0 1 4686
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_16
timestamp 1626486988
transform 1 0 -3839 0 1 6500
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_17
timestamp 1626486988
transform 1 0 -8610 0 1 7962
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_38
timestamp 1626486988
transform 1 0 -8648 0 1 9784
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_39
timestamp 1626486988
transform 1 0 -10678 0 1 9784
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_19
timestamp 1626486988
transform 1 0 -12124 0 1 9780
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_15
timestamp 1626486988
transform -1 0 -11093 0 1 7962
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_16
timestamp 1626486988
transform -1 0 -6322 0 1 7964
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_37
timestamp 1626486988
transform 1 0 -6488 0 1 9784
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_36
timestamp 1626486988
transform 1 0 -4448 0 1 9784
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_18
timestamp 1626486988
transform -1 0 -2958 0 1 9782
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_14
timestamp 1626486988
transform 1 0 -3839 0 1 7964
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_15
timestamp 1626486988
transform 1 0 -8610 0 1 13698
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_34
timestamp 1626486988
transform 1 0 -8648 0 1 11884
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_35
timestamp 1626486988
transform 1 0 -10678 0 1 11884
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_17
timestamp 1626486988
transform 1 0 -12124 0 1 11884
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_13
timestamp 1626486988
transform -1 0 -11093 0 1 13698
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_14
timestamp 1626486988
transform -1 0 -6322 0 1 13700
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_33
timestamp 1626486988
transform 1 0 -6488 0 1 11884
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_32
timestamp 1626486988
transform 1 0 -4448 0 1 11884
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_16
timestamp 1626486988
transform -1 0 -2958 0 1 11886
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_12
timestamp 1626486988
transform 1 0 -3839 0 1 13700
box -1350 -300 1232 300
use txgate  txgate_7
timestamp 1626486988
transform 1 0 -84715 0 1 -42708
box 74185 57360 76542 59116
use txgate  txgate_6
timestamp 1626486988
transform 1 0 -87315 0 1 -42708
box 74185 57360 76542 59116
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0
timestamp 1626486988
transform -1 0 -7834 0 1 15218
box -38 -48 314 592
use diff_fold_casc_ota  diff_fold_casc_ota_1
timestamp 1626486988
transform 1 0 10950 0 1 26540
box -12400 -27248 25000 1800
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_31
timestamp 1626486988
transform 1 0 38946 0 1 2850
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_15
timestamp 1626486988
transform 1 0 37500 0 1 2846
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_11
timestamp 1626486988
transform -1 0 38531 0 1 1028
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_12
timestamp 1626486988
transform -1 0 43302 0 1 1030
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_13
timestamp 1626486988
transform 1 0 41014 0 1 1028
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_29
timestamp 1626486988
transform 1 0 40976 0 1 2850
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_30
timestamp 1626486988
transform 1 0 43136 0 1 2850
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_28
timestamp 1626486988
transform 1 0 45176 0 1 2850
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_10
timestamp 1626486988
transform 1 0 45785 0 1 1030
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_14
timestamp 1626486988
transform -1 0 46666 0 1 2848
box -350 -900 244 900
use txgate  txgate_4
timestamp 1626486988
transform 1 0 -25531 0 1 -54506
box 74185 57360 76542 59116
use txgate  txgate_5
timestamp 1626486988
transform 1 0 -25531 0 1 -56596
box 74185 57360 76542 59116
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_27
timestamp 1626486988
transform 1 0 38946 0 1 4950
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_13
timestamp 1626486988
transform 1 0 37500 0 1 4950
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_9
timestamp 1626486988
transform -1 0 38531 0 1 6764
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_10
timestamp 1626486988
transform -1 0 43302 0 1 6766
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_11
timestamp 1626486988
transform 1 0 41014 0 1 6764
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_25
timestamp 1626486988
transform 1 0 40976 0 1 4950
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_26
timestamp 1626486988
transform 1 0 43136 0 1 4950
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_24
timestamp 1626486988
transform 1 0 45176 0 1 4950
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_8
timestamp 1626486988
transform 1 0 45785 0 1 6766
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_12
timestamp 1626486988
transform -1 0 46666 0 1 4952
box -350 -900 244 900
use txgate  txgate_3
timestamp 1626486988
transform 1 0 -25531 0 1 -52506
box 74185 57360 76542 59116
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_23
timestamp 1626486988
transform 1 0 38928 0 1 10452
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_11
timestamp 1626486988
transform 1 0 37482 0 1 10448
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_7
timestamp 1626486988
transform -1 0 38513 0 1 8630
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_8
timestamp 1626486988
transform 1 0 40996 0 1 8630
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_9
timestamp 1626486988
transform -1 0 43284 0 1 8632
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_21
timestamp 1626486988
transform 1 0 43118 0 1 10452
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_22
timestamp 1626486988
transform 1 0 40958 0 1 10452
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_20
timestamp 1626486988
transform 1 0 45158 0 1 10452
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_6
timestamp 1626486988
transform 1 0 45767 0 1 8632
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_10
timestamp 1626486988
transform -1 0 46648 0 1 10450
box -350 -900 244 900
use txgate  txgate_2
timestamp 1626486988
transform 1 0 -25531 0 1 -50542
box 74185 57360 76542 59116
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_19
timestamp 1626486988
transform 1 0 38928 0 1 12552
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_9
timestamp 1626486988
transform 1 0 37482 0 1 12552
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_17
timestamp 1626486988
transform 1 0 43118 0 1 12552
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_18
timestamp 1626486988
transform 1 0 40958 0 1 12552
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_16
timestamp 1626486988
transform 1 0 45158 0 1 12552
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_8
timestamp 1626486988
transform -1 0 46648 0 1 12554
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_15
timestamp 1626486988
transform 1 0 39076 0 1 16574
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_7
timestamp 1626486988
transform 1 0 37630 0 1 16570
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_5
timestamp 1626486988
transform -1 0 38513 0 1 14566
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_6
timestamp 1626486988
transform -1 0 43284 0 1 14568
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_7
timestamp 1626486988
transform 1 0 40996 0 1 14566
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_13
timestamp 1626486988
transform 1 0 43266 0 1 16574
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_14
timestamp 1626486988
transform 1 0 41106 0 1 16574
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_5
timestamp 1626486988
transform -1 0 45566 0 1 14568
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_12
timestamp 1626486988
transform 1 0 45306 0 1 16574
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_4
timestamp 1626486988
transform -1 0 47678 0 1 14568
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_10
timestamp 1626486988
transform 1 0 49502 0 1 16574
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_11
timestamp 1626486988
transform 1 0 47462 0 1 16574
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_4
timestamp 1626486988
transform 1 0 50161 0 1 14568
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_6
timestamp 1626486988
transform -1 0 51042 0 1 16570
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_9
timestamp 1626486988
transform 1 0 39076 0 1 18674
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_5
timestamp 1626486988
transform 1 0 37630 0 1 18674
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_3
timestamp 1626486988
transform -1 0 38513 0 1 20726
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_2
timestamp 1626486988
transform -1 0 43284 0 1 20728
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_3
timestamp 1626486988
transform 1 0 40996 0 1 20726
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_7
timestamp 1626486988
transform 1 0 43266 0 1 18674
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_8
timestamp 1626486988
transform 1 0 41106 0 1 18674
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_1
timestamp 1626486988
transform -1 0 45392 0 1 20728
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_6
timestamp 1626486988
transform 1 0 45306 0 1 18674
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_0
timestamp 1626486988
transform -1 0 47678 0 1 20728
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_4
timestamp 1626486988
transform 1 0 49502 0 1 18674
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_5
timestamp 1626486988
transform 1 0 47462 0 1 18674
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_2
timestamp 1626486988
transform 1 0 50161 0 1 20728
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_4
timestamp 1626486988
transform -1 0 51042 0 1 18674
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_2
timestamp 1626486988
transform 1 0 38968 0 1 22612
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_3
timestamp 1626486988
transform 1 0 38968 0 1 24712
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_2
timestamp 1626486988
transform 1 0 37516 0 1 24716
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_3
timestamp 1626486988
transform 1 0 37516 0 1 22612
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_0
timestamp 1626486988
transform 1 0 40998 0 1 22612
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_1
timestamp 1626486988
transform 1 0 40998 0 1 24712
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_0
timestamp 1626486988
transform 1 0 42616 0 1 24716
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_1
timestamp 1626486988
transform 1 0 42616 0 1 22612
box -350 -900 244 900
use txgate  txgate_0
timestamp 1626486988
transform 1 0 -26957 0 1 -33578
box 74185 57360 76542 59116
use txgate  txgate_1
timestamp 1626486988
transform 1 0 -26957 0 1 -35578
box 74185 57360 76542 59116
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_1
timestamp 1626486988
transform -1 0 38400 0 1 26180
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_0
timestamp 1626486988
transform -1 0 41400 0 1 26180
box -1350 -300 1232 300
use diff_fold_casc_ota  diff_fold_casc_ota_0
timestamp 1626486988
transform 1 0 64950 0 1 26540
box -12400 -27248 25000 1800
<< labels >>
flabel metal4 s -9700 5602 -9690 5614 1 FreeSans 600 0 0 0 vip1
flabel metal4 s -9752 1570 -9732 1586 1 FreeSans 600 0 0 0 vim1
flabel metal4 s -5616 -342 -5562 -296 1 FreeSans 600 0 0 0 VSS
flabel metal4 s 39914 1890 39924 1898 1 FreeSans 600 0 0 0 venp1
flabel metal4 s 39912 5932 39922 5950 1 FreeSans 600 0 0 0 venm1
flabel metal4 s 39872 9472 39892 9486 1 FreeSans 600 0 0 0 vim2
flabel metal4 s 39942 13524 39962 13540 1 FreeSans 600 0 0 0 vip2
flabel metal4 s 40082 15590 40102 15606 1 FreeSans 600 0 0 0 venp2
flabel metal4 s 40024 19636 40048 19656 1 FreeSans 600 0 0 0 venm2
flabel metal4 s 40068 25698 40084 25712 1 FreeSans 600 0 0 0 vop
flabel metal4 s 49508 27900 49618 28008 1 FreeSans 600 0 0 0 VDD
flabel metal2 s 50956 4528 50982 4554 1 FreeSans 600 0 0 0 gain_ctrl_0
flabel metal2 s 49538 23440 49558 23458 1 FreeSans 600 0 0 0 gain_ctrl_1
flabel metal4 s 36296 7672 36328 7702 1 FreeSans 600 0 0 0 vocm
flabel metal1 s 3968 4954 3982 4962 1 FreeSans 600 0 0 0 ibiasn1
flabel metal1 s 57962 4966 57978 4972 1 FreeSans 600 0 0 0 ibiasn2
flabel metal1 s -7768 15456 -7762 15460 1 FreeSans 600 0 0 0 rst_n
flabel metal1 s -8136 15450 -8128 15458 1 FreeSans 600 0 0 0 rst
flabel metal4 s -9728 8802 -9684 8828 1 FreeSans 600 0 0 0 vop1
flabel metal4 s -9734 12846 -9714 12872 1 FreeSans 600 0 0 0 vom1
flabel metal3 s -9770 8556 -9744 8576 1 FreeSans 600 0 0 0 vim1
flabel metal3 s -9338 5886 -9298 5918 1 FreeSans 600 0 0 0 vhpf
flabel metal3 s -9718 1372 -9700 1386 1 FreeSans 600 0 0 0 vincm
flabel metal3 s 39912 1630 39926 1644 1 FreeSans 600 0 0 0 vop1
flabel metal3 s 39900 6144 39910 6156 1 FreeSans 600 0 0 0 vom1
flabel metal3 s 39848 9234 39866 9256 1 FreeSans 600 0 0 0 vop1
flabel metal3 s 39924 13774 39940 13786 1 FreeSans 600 0 0 0 vom1
flabel metal3 s 40106 19872 40122 19884 1 FreeSans 600 0 0 0 vip2
flabel metal3 s 40076 15316 40096 15328 1 FreeSans 600 0 0 0 vim2
flabel metal2 s 40896 23642 40916 23660 1 FreeSans 600 0 0 0 vim2
flabel metal4 s 39646 23514 39664 23536 1 FreeSans 600 0 0 0 vip2
flabel metal4 s 41878 23258 41900 23278 1 FreeSans 600 0 0 0 vom
flabel metal3 s -10202 13080 -10184 13090 1 FreeSans 600 0 0 0 vip1
<< end >>
