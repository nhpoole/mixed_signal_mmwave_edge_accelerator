magic
tech sky130A
magscale 1 2
timestamp 1620620197
<< error_p >>
rect -560 172 -502 178
rect -442 172 -384 178
rect -324 172 -266 178
rect -206 172 -148 178
rect -88 172 -30 178
rect 30 172 88 178
rect 148 172 206 178
rect 266 172 324 178
rect 384 172 442 178
rect 502 172 560 178
rect -560 138 -548 172
rect -442 138 -430 172
rect -324 138 -312 172
rect -206 138 -194 172
rect -88 138 -76 172
rect 30 138 42 172
rect 148 138 160 172
rect 266 138 278 172
rect 384 138 396 172
rect 502 138 514 172
rect -560 132 -502 138
rect -442 132 -384 138
rect -324 132 -266 138
rect -206 132 -148 138
rect -88 132 -30 138
rect 30 132 88 138
rect 148 132 206 138
rect 266 132 324 138
rect 384 132 442 138
rect 502 132 560 138
rect -560 -138 -502 -132
rect -442 -138 -384 -132
rect -324 -138 -266 -132
rect -206 -138 -148 -132
rect -88 -138 -30 -132
rect 30 -138 88 -132
rect 148 -138 206 -132
rect 266 -138 324 -132
rect 384 -138 442 -132
rect 502 -138 560 -132
rect -560 -172 -548 -138
rect -442 -172 -430 -138
rect -324 -172 -312 -138
rect -206 -172 -194 -138
rect -88 -172 -76 -138
rect 30 -172 42 -138
rect 148 -172 160 -138
rect 266 -172 278 -138
rect 384 -172 396 -138
rect 502 -172 514 -138
rect -560 -178 -502 -172
rect -442 -178 -384 -172
rect -324 -178 -266 -172
rect -206 -178 -148 -172
rect -88 -178 -30 -172
rect 30 -178 88 -172
rect 148 -178 206 -172
rect 266 -178 324 -172
rect 384 -178 442 -172
rect 502 -178 560 -172
<< nmoslvt >>
rect -561 -100 -501 100
rect -443 -100 -383 100
rect -325 -100 -265 100
rect -207 -100 -147 100
rect -89 -100 -29 100
rect 29 -100 89 100
rect 147 -100 207 100
rect 265 -100 325 100
rect 383 -100 443 100
rect 501 -100 561 100
<< ndiff >>
rect -619 88 -561 100
rect -619 -88 -607 88
rect -573 -88 -561 88
rect -619 -100 -561 -88
rect -501 88 -443 100
rect -501 -88 -489 88
rect -455 -88 -443 88
rect -501 -100 -443 -88
rect -383 88 -325 100
rect -383 -88 -371 88
rect -337 -88 -325 88
rect -383 -100 -325 -88
rect -265 88 -207 100
rect -265 -88 -253 88
rect -219 -88 -207 88
rect -265 -100 -207 -88
rect -147 88 -89 100
rect -147 -88 -135 88
rect -101 -88 -89 88
rect -147 -100 -89 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 89 88 147 100
rect 89 -88 101 88
rect 135 -88 147 88
rect 89 -100 147 -88
rect 207 88 265 100
rect 207 -88 219 88
rect 253 -88 265 88
rect 207 -100 265 -88
rect 325 88 383 100
rect 325 -88 337 88
rect 371 -88 383 88
rect 325 -100 383 -88
rect 443 88 501 100
rect 443 -88 455 88
rect 489 -88 501 88
rect 443 -100 501 -88
rect 561 88 619 100
rect 561 -88 573 88
rect 607 -88 619 88
rect 561 -100 619 -88
<< ndiffc >>
rect -607 -88 -573 88
rect -489 -88 -455 88
rect -371 -88 -337 88
rect -253 -88 -219 88
rect -135 -88 -101 88
rect -17 -88 17 88
rect 101 -88 135 88
rect 219 -88 253 88
rect 337 -88 371 88
rect 455 -88 489 88
rect 573 -88 607 88
<< poly >>
rect -564 172 -498 188
rect -564 138 -548 172
rect -514 138 -498 172
rect -564 122 -498 138
rect -446 172 -380 188
rect -446 138 -430 172
rect -396 138 -380 172
rect -446 122 -380 138
rect -328 172 -262 188
rect -328 138 -312 172
rect -278 138 -262 172
rect -328 122 -262 138
rect -210 172 -144 188
rect -210 138 -194 172
rect -160 138 -144 172
rect -210 122 -144 138
rect -92 172 -26 188
rect -92 138 -76 172
rect -42 138 -26 172
rect -92 122 -26 138
rect 26 172 92 188
rect 26 138 42 172
rect 76 138 92 172
rect 26 122 92 138
rect 144 172 210 188
rect 144 138 160 172
rect 194 138 210 172
rect 144 122 210 138
rect 262 172 328 188
rect 262 138 278 172
rect 312 138 328 172
rect 262 122 328 138
rect 380 172 446 188
rect 380 138 396 172
rect 430 138 446 172
rect 380 122 446 138
rect 498 172 564 188
rect 498 138 514 172
rect 548 138 564 172
rect 498 122 564 138
rect -561 100 -501 122
rect -443 100 -383 122
rect -325 100 -265 122
rect -207 100 -147 122
rect -89 100 -29 122
rect 29 100 89 122
rect 147 100 207 122
rect 265 100 325 122
rect 383 100 443 122
rect 501 100 561 122
rect -561 -122 -501 -100
rect -443 -122 -383 -100
rect -325 -122 -265 -100
rect -207 -122 -147 -100
rect -89 -122 -29 -100
rect 29 -122 89 -100
rect 147 -122 207 -100
rect 265 -122 325 -100
rect 383 -122 443 -100
rect 501 -122 561 -100
rect -564 -138 -498 -122
rect -564 -172 -548 -138
rect -514 -172 -498 -138
rect -564 -188 -498 -172
rect -446 -138 -380 -122
rect -446 -172 -430 -138
rect -396 -172 -380 -138
rect -446 -188 -380 -172
rect -328 -138 -262 -122
rect -328 -172 -312 -138
rect -278 -172 -262 -138
rect -328 -188 -262 -172
rect -210 -138 -144 -122
rect -210 -172 -194 -138
rect -160 -172 -144 -138
rect -210 -188 -144 -172
rect -92 -138 -26 -122
rect -92 -172 -76 -138
rect -42 -172 -26 -138
rect -92 -188 -26 -172
rect 26 -138 92 -122
rect 26 -172 42 -138
rect 76 -172 92 -138
rect 26 -188 92 -172
rect 144 -138 210 -122
rect 144 -172 160 -138
rect 194 -172 210 -138
rect 144 -188 210 -172
rect 262 -138 328 -122
rect 262 -172 278 -138
rect 312 -172 328 -138
rect 262 -188 328 -172
rect 380 -138 446 -122
rect 380 -172 396 -138
rect 430 -172 446 -138
rect 380 -188 446 -172
rect 498 -138 564 -122
rect 498 -172 514 -138
rect 548 -172 564 -138
rect 498 -188 564 -172
<< polycont >>
rect -548 138 -514 172
rect -430 138 -396 172
rect -312 138 -278 172
rect -194 138 -160 172
rect -76 138 -42 172
rect 42 138 76 172
rect 160 138 194 172
rect 278 138 312 172
rect 396 138 430 172
rect 514 138 548 172
rect -548 -172 -514 -138
rect -430 -172 -396 -138
rect -312 -172 -278 -138
rect -194 -172 -160 -138
rect -76 -172 -42 -138
rect 42 -172 76 -138
rect 160 -172 194 -138
rect 278 -172 312 -138
rect 396 -172 430 -138
rect 514 -172 548 -138
<< locali >>
rect -564 138 -548 172
rect -514 138 -498 172
rect -446 138 -430 172
rect -396 138 -380 172
rect -328 138 -312 172
rect -278 138 -262 172
rect -210 138 -194 172
rect -160 138 -144 172
rect -92 138 -76 172
rect -42 138 -26 172
rect 26 138 42 172
rect 76 138 92 172
rect 144 138 160 172
rect 194 138 210 172
rect 262 138 278 172
rect 312 138 328 172
rect 380 138 396 172
rect 430 138 446 172
rect 498 138 514 172
rect 548 138 564 172
rect -607 88 -573 104
rect -607 -104 -573 -88
rect -489 88 -455 104
rect -489 -104 -455 -88
rect -371 88 -337 104
rect -371 -104 -337 -88
rect -253 88 -219 104
rect -253 -104 -219 -88
rect -135 88 -101 104
rect -135 -104 -101 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 101 88 135 104
rect 101 -104 135 -88
rect 219 88 253 104
rect 219 -104 253 -88
rect 337 88 371 104
rect 337 -104 371 -88
rect 455 88 489 104
rect 455 -104 489 -88
rect 573 88 607 104
rect 573 -104 607 -88
rect -564 -172 -548 -138
rect -514 -172 -498 -138
rect -446 -172 -430 -138
rect -396 -172 -380 -138
rect -328 -172 -312 -138
rect -278 -172 -262 -138
rect -210 -172 -194 -138
rect -160 -172 -144 -138
rect -92 -172 -76 -138
rect -42 -172 -26 -138
rect 26 -172 42 -138
rect 76 -172 92 -138
rect 144 -172 160 -138
rect 194 -172 210 -138
rect 262 -172 278 -138
rect 312 -172 328 -138
rect 380 -172 396 -138
rect 430 -172 446 -138
rect 498 -172 514 -138
rect 548 -172 564 -138
<< viali >>
rect -548 138 -514 172
rect -430 138 -396 172
rect -312 138 -278 172
rect -194 138 -160 172
rect -76 138 -42 172
rect 42 138 76 172
rect 160 138 194 172
rect 278 138 312 172
rect 396 138 430 172
rect 514 138 548 172
rect -607 -88 -573 88
rect -489 -88 -455 88
rect -371 -88 -337 88
rect -253 -88 -219 88
rect -135 -88 -101 88
rect -17 -88 17 88
rect 101 -88 135 88
rect 219 -88 253 88
rect 337 -88 371 88
rect 455 -88 489 88
rect 573 -88 607 88
rect -548 -172 -514 -138
rect -430 -172 -396 -138
rect -312 -172 -278 -138
rect -194 -172 -160 -138
rect -76 -172 -42 -138
rect 42 -172 76 -138
rect 160 -172 194 -138
rect 278 -172 312 -138
rect 396 -172 430 -138
rect 514 -172 548 -138
<< metal1 >>
rect -560 172 -502 178
rect -560 138 -548 172
rect -514 138 -502 172
rect -560 132 -502 138
rect -442 172 -384 178
rect -442 138 -430 172
rect -396 138 -384 172
rect -442 132 -384 138
rect -324 172 -266 178
rect -324 138 -312 172
rect -278 138 -266 172
rect -324 132 -266 138
rect -206 172 -148 178
rect -206 138 -194 172
rect -160 138 -148 172
rect -206 132 -148 138
rect -88 172 -30 178
rect -88 138 -76 172
rect -42 138 -30 172
rect -88 132 -30 138
rect 30 172 88 178
rect 30 138 42 172
rect 76 138 88 172
rect 30 132 88 138
rect 148 172 206 178
rect 148 138 160 172
rect 194 138 206 172
rect 148 132 206 138
rect 266 172 324 178
rect 266 138 278 172
rect 312 138 324 172
rect 266 132 324 138
rect 384 172 442 178
rect 384 138 396 172
rect 430 138 442 172
rect 384 132 442 138
rect 502 172 560 178
rect 502 138 514 172
rect 548 138 560 172
rect 502 132 560 138
rect -613 88 -567 100
rect -613 -88 -607 88
rect -573 -88 -567 88
rect -613 -100 -567 -88
rect -495 88 -449 100
rect -495 -88 -489 88
rect -455 -88 -449 88
rect -495 -100 -449 -88
rect -377 88 -331 100
rect -377 -88 -371 88
rect -337 -88 -331 88
rect -377 -100 -331 -88
rect -259 88 -213 100
rect -259 -88 -253 88
rect -219 -88 -213 88
rect -259 -100 -213 -88
rect -141 88 -95 100
rect -141 -88 -135 88
rect -101 -88 -95 88
rect -141 -100 -95 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 95 88 141 100
rect 95 -88 101 88
rect 135 -88 141 88
rect 95 -100 141 -88
rect 213 88 259 100
rect 213 -88 219 88
rect 253 -88 259 88
rect 213 -100 259 -88
rect 331 88 377 100
rect 331 -88 337 88
rect 371 -88 377 88
rect 331 -100 377 -88
rect 449 88 495 100
rect 449 -88 455 88
rect 489 -88 495 88
rect 449 -100 495 -88
rect 567 88 613 100
rect 567 -88 573 88
rect 607 -88 613 88
rect 567 -100 613 -88
rect -560 -138 -502 -132
rect -560 -172 -548 -138
rect -514 -172 -502 -138
rect -560 -178 -502 -172
rect -442 -138 -384 -132
rect -442 -172 -430 -138
rect -396 -172 -384 -138
rect -442 -178 -384 -172
rect -324 -138 -266 -132
rect -324 -172 -312 -138
rect -278 -172 -266 -138
rect -324 -178 -266 -172
rect -206 -138 -148 -132
rect -206 -172 -194 -138
rect -160 -172 -148 -138
rect -206 -178 -148 -172
rect -88 -138 -30 -132
rect -88 -172 -76 -138
rect -42 -172 -30 -138
rect -88 -178 -30 -172
rect 30 -138 88 -132
rect 30 -172 42 -138
rect 76 -172 88 -138
rect 30 -178 88 -172
rect 148 -138 206 -132
rect 148 -172 160 -138
rect 194 -172 206 -138
rect 148 -178 206 -172
rect 266 -138 324 -132
rect 266 -172 278 -138
rect 312 -172 324 -138
rect 266 -178 324 -172
rect 384 -138 442 -132
rect 384 -172 396 -138
rect 430 -172 442 -138
rect 384 -178 442 -172
rect 502 -138 560 -132
rect 502 -172 514 -138
rect 548 -172 560 -138
rect 502 -178 560 -172
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string parameters w 1 l 0.3 m 1 nf 10 diffcov 100 polycov 60 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
