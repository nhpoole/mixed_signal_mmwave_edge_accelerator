* Stimulus file.

.param Ibias_comp=10u vincm_comp=0.9 vsig=0 vdd=1.8 Wp_comp=4 Wn_comp=2

vdd VDD GND 'vdd'
vip vip GND pwl(0 'vincm_comp' 10n 'vincm_comp' 10.1n 'vincm_comp+5m' 50n 'vincm_comp+5m' 50.1n 'vincm_comp-5m' 90n 'vincm_comp-5m' 90.1n 'vincm_comp+5m' 130n 'vincm_comp+5m')
vim vim GND pwl(0 'vincm_comp' 10n 'vincm_comp' 10.1n 'vincm_comp-5m' 50n 'vincm_comp-5m' 50.1n 'vincm_comp+5m' 90n 'vincm_comp+5m' 90.1n 'vincm_comp-5m' 130n 'vincm_comp-5m')
*vip vip GND dc 'vincm_comp+vsig' ac 0.5 0
*vim vim GND dc 'vincm_comp-vsig' ac 0.5 180

.control
options savecurrents
save all
+ @m.xm1.msky130_fd_pr__nfet_01v8_lvt[id]
+ @m.xm1.msky130_fd_pr__nfet_01v8_lvt[vth]
+ @m.xm2.msky130_fd_pr__nfet_01v8[gm]
+ @m.xm2.msky130_fd_pr__nfet_01v8[id]
+ @m.xm2.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm3.msky130_fd_pr__pfet_01v8[id]
+ @m.xm3.msky130_fd_pr__pfet_01v8[vth]
+ @m.xm4.msky130_fd_pr__nfet_01v8_lvt[id]
+ @m.xm4.msky130_fd_pr__nfet_01v8_lvt[vth]
+ @m.xm5.msky130_fd_pr__pfet_01v8[id]
+ @m.xm5.msky130_fd_pr__pfet_01v8[vth]
+ @m.xm6.msky130_fd_pr__pfet_01v8[id]
+ @m.xm6.msky130_fd_pr__pfet_01v8[vth]
+ @m.xm7.msky130_fd_pr__pfet_01v8[id]
+ @m.xm7.msky130_fd_pr__pfet_01v8[vth]
+ @m.xm8.msky130_fd_pr__pfet_01v8[id]
+ @m.xm8.msky130_fd_pr__pfet_01v8[vth]
+ @m.xm9.msky130_fd_pr__nfet_01v8[id]
+ @m.xm9.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm10.msky130_fd_pr__pfet_01v8[id]
+ @m.xm10.msky130_fd_pr__pfet_01v8[vth]
+ @m.xm11.msky130_fd_pr__nfet_01v8[id]
+ @m.xm11.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm12.msky130_fd_pr__nfet_01v8[id]
+ @m.xm12.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm13.msky130_fd_pr__nfet_01v8[id]
+ @m.xm13.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm14.msky130_fd_pr__nfet_01v8[id]
+ @m.xm14.msky130_fd_pr__nfet_01v8[vth]
+ @m.xm15.msky130_fd_pr__pfet_01v8_hvt[id]
+ @m.xm15.msky130_fd_pr__pfet_01v8_hvt[vth]

op
run
print all
*write comparator_op.raw

tran 0.1n 130n
run
write comparator_tran.raw

*dc vip 0.8999 0.9001 1e-7
*run
*write comparator_dc.raw

*ac dec 100 0.1 1g
*run
*write comparator_ac.raw
quit
.endc
