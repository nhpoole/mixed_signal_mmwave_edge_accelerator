magic
tech sky130A
magscale 1 2
timestamp 1626065694
<< checkpaint >>
rect -1610 -2360 1609 2360
<< metal3 >>
rect -350 1072 349 1100
rect -350 1008 265 1072
rect 329 1008 349 1072
rect -350 992 349 1008
rect -350 928 265 992
rect 329 928 349 992
rect -350 912 349 928
rect -350 848 265 912
rect 329 848 349 912
rect -350 832 349 848
rect -350 768 265 832
rect 329 768 349 832
rect -350 752 349 768
rect -350 688 265 752
rect 329 688 349 752
rect -350 672 349 688
rect -350 608 265 672
rect 329 608 349 672
rect -350 592 349 608
rect -350 528 265 592
rect 329 528 349 592
rect -350 512 349 528
rect -350 448 265 512
rect 329 448 349 512
rect -350 432 349 448
rect -350 368 265 432
rect 329 368 349 432
rect -350 352 349 368
rect -350 288 265 352
rect 329 288 349 352
rect -350 272 349 288
rect -350 208 265 272
rect 329 208 349 272
rect -350 192 349 208
rect -350 128 265 192
rect 329 128 349 192
rect -350 112 349 128
rect -350 48 265 112
rect 329 48 349 112
rect -350 32 349 48
rect -350 -32 265 32
rect 329 -32 349 32
rect -350 -48 349 -32
rect -350 -112 265 -48
rect 329 -112 349 -48
rect -350 -128 349 -112
rect -350 -192 265 -128
rect 329 -192 349 -128
rect -350 -208 349 -192
rect -350 -272 265 -208
rect 329 -272 349 -208
rect -350 -288 349 -272
rect -350 -352 265 -288
rect 329 -352 349 -288
rect -350 -368 349 -352
rect -350 -432 265 -368
rect 329 -432 349 -368
rect -350 -448 349 -432
rect -350 -512 265 -448
rect 329 -512 349 -448
rect -350 -528 349 -512
rect -350 -592 265 -528
rect 329 -592 349 -528
rect -350 -608 349 -592
rect -350 -672 265 -608
rect 329 -672 349 -608
rect -350 -688 349 -672
rect -350 -752 265 -688
rect 329 -752 349 -688
rect -350 -768 349 -752
rect -350 -832 265 -768
rect 329 -832 349 -768
rect -350 -848 349 -832
rect -350 -912 265 -848
rect 329 -912 349 -848
rect -350 -928 349 -912
rect -350 -992 265 -928
rect 329 -992 349 -928
rect -350 -1008 349 -992
rect -350 -1072 265 -1008
rect 329 -1072 349 -1008
rect -350 -1100 349 -1072
<< via3 >>
rect 265 1008 329 1072
rect 265 928 329 992
rect 265 848 329 912
rect 265 768 329 832
rect 265 688 329 752
rect 265 608 329 672
rect 265 528 329 592
rect 265 448 329 512
rect 265 368 329 432
rect 265 288 329 352
rect 265 208 329 272
rect 265 128 329 192
rect 265 48 329 112
rect 265 -32 329 32
rect 265 -112 329 -48
rect 265 -192 329 -128
rect 265 -272 329 -208
rect 265 -352 329 -288
rect 265 -432 329 -368
rect 265 -512 329 -448
rect 265 -592 329 -528
rect 265 -672 329 -608
rect 265 -752 329 -688
rect 265 -832 329 -768
rect 265 -912 329 -848
rect 265 -992 329 -928
rect 265 -1072 329 -1008
<< mimcap >>
rect -250 952 150 1000
rect -250 -952 -202 952
rect 102 -952 150 952
rect -250 -1000 150 -952
<< mimcapcontact >>
rect -202 -952 102 952
<< metal4 >>
rect 249 1072 345 1088
rect 249 1008 265 1072
rect 329 1008 345 1072
rect 249 992 345 1008
rect -211 952 111 961
rect -211 -952 -202 952
rect 102 -952 111 952
rect -211 -961 111 -952
rect 249 928 265 992
rect 329 928 345 992
rect 249 912 345 928
rect 249 848 265 912
rect 329 848 345 912
rect 249 832 345 848
rect 249 768 265 832
rect 329 768 345 832
rect 249 752 345 768
rect 249 688 265 752
rect 329 688 345 752
rect 249 672 345 688
rect 249 608 265 672
rect 329 608 345 672
rect 249 592 345 608
rect 249 528 265 592
rect 329 528 345 592
rect 249 512 345 528
rect 249 448 265 512
rect 329 448 345 512
rect 249 432 345 448
rect 249 368 265 432
rect 329 368 345 432
rect 249 352 345 368
rect 249 288 265 352
rect 329 288 345 352
rect 249 272 345 288
rect 249 208 265 272
rect 329 208 345 272
rect 249 192 345 208
rect 249 128 265 192
rect 329 128 345 192
rect 249 112 345 128
rect 249 48 265 112
rect 329 48 345 112
rect 249 32 345 48
rect 249 -32 265 32
rect 329 -32 345 32
rect 249 -48 345 -32
rect 249 -112 265 -48
rect 329 -112 345 -48
rect 249 -128 345 -112
rect 249 -192 265 -128
rect 329 -192 345 -128
rect 249 -208 345 -192
rect 249 -272 265 -208
rect 329 -272 345 -208
rect 249 -288 345 -272
rect 249 -352 265 -288
rect 329 -352 345 -288
rect 249 -368 345 -352
rect 249 -432 265 -368
rect 329 -432 345 -368
rect 249 -448 345 -432
rect 249 -512 265 -448
rect 329 -512 345 -448
rect 249 -528 345 -512
rect 249 -592 265 -528
rect 329 -592 345 -528
rect 249 -608 345 -592
rect 249 -672 265 -608
rect 329 -672 345 -608
rect 249 -688 345 -672
rect 249 -752 265 -688
rect 329 -752 345 -688
rect 249 -768 345 -752
rect 249 -832 265 -768
rect 329 -832 345 -768
rect 249 -848 345 -832
rect 249 -912 265 -848
rect 329 -912 345 -848
rect 249 -928 345 -912
rect 249 -992 265 -928
rect 329 -992 345 -928
rect 249 -1008 345 -992
rect 249 -1072 265 -1008
rect 329 -1072 345 -1008
rect 249 -1088 345 -1072
<< properties >>
string FIXED_BBOX -350 -1100 250 1100
<< end >>
