magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect -1216 -1260 4524 1750
<< nwell >>
rect 1756 0 3264 490
<< poly >>
rect 77 155 136 185
rect 1588 155 1784 185
<< locali >>
rect 60 137 94 203
rect 829 103 3246 137
<< metal1 >>
rect 848 0 876 395
rect 2496 0 2524 395
use sky130_sram_2kbyte_1rw1r_32x512_8_nmos_m1_w7_000_sli_dli_da_p  sky130_sram_2kbyte_1rw1r_32x512_8_nmos_m1_w7_000_sli_dli_da_p_0
timestamp 1626486988
transform 0 1 162 -1 0 245
box -26 -26 176 1426
use sky130_sram_2kbyte_1rw1r_32x512_8_pmos_m1_w7_000_sli_dli_da_p  sky130_sram_2kbyte_1rw1r_32x512_8_pmos_m1_w7_000_sli_dli_da_p_0
timestamp 1626486988
transform 0 1 1810 -1 0 245
box -59 -54 209 1454
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_15  sky130_sram_2kbyte_1rw1r_32x512_8_contact_15_0
timestamp 1626486988
transform 1 0 837 0 1 354
box -26 -26 76 108
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_0
timestamp 1626486988
transform 1 0 2481 0 1 187
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1
timestamp 1626486988
transform 1 0 833 0 1 187
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_16  sky130_sram_2kbyte_1rw1r_32x512_8_contact_16_0
timestamp 1626486988
transform 1 0 44 0 1 137
box 0 0 66 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_2
timestamp 1626486988
transform 1 0 833 0 1 362
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_3
timestamp 1626486988
transform 1 0 2481 0 1 362
box 0 0 58 66
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_13  sky130_sram_2kbyte_1rw1r_32x512_8_contact_13_0
timestamp 1626486988
transform 1 0 2485 0 1 354
box -59 -43 109 125
<< labels >>
rlabel metal1 s 848 0 876 395 4 gnd
rlabel metal1 s 2496 0 2524 395 4 vdd
rlabel locali s 77 170 77 170 4 A
rlabel locali s 2037 120 2037 120 4 Z
<< properties >>
string FIXED_BBOX 0 0 3246 395
<< end >>
