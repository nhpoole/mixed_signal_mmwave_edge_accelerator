magic
tech sky130A
timestamp 1626065694
<< checkpaint >>
rect -677 -654 677 654
<< metal1 >>
rect -47 13 47 24
rect -47 -13 -45 13
rect -19 -13 -13 13
rect 13 -13 19 13
rect 45 -13 47 13
rect -47 -24 47 -13
<< via1 >>
rect -45 -13 -19 13
rect -13 -13 13 13
rect 19 -13 45 13
<< metal2 >>
rect -47 13 47 24
rect -47 -13 -45 13
rect -19 -13 -13 13
rect 13 -13 19 13
rect 45 -13 47 13
rect -47 -24 47 -13
<< end >>
