magic
tech sky130A
magscale 1 2
timestamp 1621053618
<< error_p >>
rect -3549 3500 -3489 5700
rect -3469 3500 -3409 5700
rect -1230 3500 -1170 5700
rect -1150 3500 -1090 5700
rect 1089 3500 1149 5700
rect 1169 3500 1229 5700
rect 3408 3500 3468 5700
rect 3488 3500 3548 5700
rect -3549 1200 -3489 3400
rect -3469 1200 -3409 3400
rect -1230 1200 -1170 3400
rect -1150 1200 -1090 3400
rect 1089 1200 1149 3400
rect 1169 1200 1229 3400
rect 3408 1200 3468 3400
rect 3488 1200 3548 3400
rect -3549 -1100 -3489 1100
rect -3469 -1100 -3409 1100
rect -1230 -1100 -1170 1100
rect -1150 -1100 -1090 1100
rect 1089 -1100 1149 1100
rect 1169 -1100 1229 1100
rect 3408 -1100 3468 1100
rect 3488 -1100 3548 1100
rect -3549 -3400 -3489 -1200
rect -3469 -3400 -3409 -1200
rect -1230 -3400 -1170 -1200
rect -1150 -3400 -1090 -1200
rect 1089 -3400 1149 -1200
rect 1169 -3400 1229 -1200
rect 3408 -3400 3468 -1200
rect 3488 -3400 3548 -1200
rect -3549 -5700 -3489 -3500
rect -3469 -5700 -3409 -3500
rect -1230 -5700 -1170 -3500
rect -1150 -5700 -1090 -3500
rect 1089 -5700 1149 -3500
rect 1169 -5700 1229 -3500
rect 3408 -5700 3468 -3500
rect 3488 -5700 3548 -3500
<< metal3 >>
rect -5788 5672 -3489 5700
rect -5788 3528 -3573 5672
rect -3509 3528 -3489 5672
rect -5788 3500 -3489 3528
rect -3469 5672 -1170 5700
rect -3469 3528 -1254 5672
rect -1190 3528 -1170 5672
rect -3469 3500 -1170 3528
rect -1150 5672 1149 5700
rect -1150 3528 1065 5672
rect 1129 3528 1149 5672
rect -1150 3500 1149 3528
rect 1169 5672 3468 5700
rect 1169 3528 3384 5672
rect 3448 3528 3468 5672
rect 1169 3500 3468 3528
rect 3488 5672 5787 5700
rect 3488 3528 5703 5672
rect 5767 3528 5787 5672
rect 3488 3500 5787 3528
rect -5788 3372 -3489 3400
rect -5788 1228 -3573 3372
rect -3509 1228 -3489 3372
rect -5788 1200 -3489 1228
rect -3469 3372 -1170 3400
rect -3469 1228 -1254 3372
rect -1190 1228 -1170 3372
rect -3469 1200 -1170 1228
rect -1150 3372 1149 3400
rect -1150 1228 1065 3372
rect 1129 1228 1149 3372
rect -1150 1200 1149 1228
rect 1169 3372 3468 3400
rect 1169 1228 3384 3372
rect 3448 1228 3468 3372
rect 1169 1200 3468 1228
rect 3488 3372 5787 3400
rect 3488 1228 5703 3372
rect 5767 1228 5787 3372
rect 3488 1200 5787 1228
rect -5788 1072 -3489 1100
rect -5788 -1072 -3573 1072
rect -3509 -1072 -3489 1072
rect -5788 -1100 -3489 -1072
rect -3469 1072 -1170 1100
rect -3469 -1072 -1254 1072
rect -1190 -1072 -1170 1072
rect -3469 -1100 -1170 -1072
rect -1150 1072 1149 1100
rect -1150 -1072 1065 1072
rect 1129 -1072 1149 1072
rect -1150 -1100 1149 -1072
rect 1169 1072 3468 1100
rect 1169 -1072 3384 1072
rect 3448 -1072 3468 1072
rect 1169 -1100 3468 -1072
rect 3488 1072 5787 1100
rect 3488 -1072 5703 1072
rect 5767 -1072 5787 1072
rect 3488 -1100 5787 -1072
rect -5788 -1228 -3489 -1200
rect -5788 -3372 -3573 -1228
rect -3509 -3372 -3489 -1228
rect -5788 -3400 -3489 -3372
rect -3469 -1228 -1170 -1200
rect -3469 -3372 -1254 -1228
rect -1190 -3372 -1170 -1228
rect -3469 -3400 -1170 -3372
rect -1150 -1228 1149 -1200
rect -1150 -3372 1065 -1228
rect 1129 -3372 1149 -1228
rect -1150 -3400 1149 -3372
rect 1169 -1228 3468 -1200
rect 1169 -3372 3384 -1228
rect 3448 -3372 3468 -1228
rect 1169 -3400 3468 -3372
rect 3488 -1228 5787 -1200
rect 3488 -3372 5703 -1228
rect 5767 -3372 5787 -1228
rect 3488 -3400 5787 -3372
rect -5788 -3528 -3489 -3500
rect -5788 -5672 -3573 -3528
rect -3509 -5672 -3489 -3528
rect -5788 -5700 -3489 -5672
rect -3469 -3528 -1170 -3500
rect -3469 -5672 -1254 -3528
rect -1190 -5672 -1170 -3528
rect -3469 -5700 -1170 -5672
rect -1150 -3528 1149 -3500
rect -1150 -5672 1065 -3528
rect 1129 -5672 1149 -3528
rect -1150 -5700 1149 -5672
rect 1169 -3528 3468 -3500
rect 1169 -5672 3384 -3528
rect 3448 -5672 3468 -3528
rect 1169 -5700 3468 -5672
rect 3488 -3528 5787 -3500
rect 3488 -5672 5703 -3528
rect 5767 -5672 5787 -3528
rect 3488 -5700 5787 -5672
<< via3 >>
rect -3573 3528 -3509 5672
rect -1254 3528 -1190 5672
rect 1065 3528 1129 5672
rect 3384 3528 3448 5672
rect 5703 3528 5767 5672
rect -3573 1228 -3509 3372
rect -1254 1228 -1190 3372
rect 1065 1228 1129 3372
rect 3384 1228 3448 3372
rect 5703 1228 5767 3372
rect -3573 -1072 -3509 1072
rect -1254 -1072 -1190 1072
rect 1065 -1072 1129 1072
rect 3384 -1072 3448 1072
rect 5703 -1072 5767 1072
rect -3573 -3372 -3509 -1228
rect -1254 -3372 -1190 -1228
rect 1065 -3372 1129 -1228
rect 3384 -3372 3448 -1228
rect 5703 -3372 5767 -1228
rect -3573 -5672 -3509 -3528
rect -1254 -5672 -1190 -3528
rect 1065 -5672 1129 -3528
rect 3384 -5672 3448 -3528
rect 5703 -5672 5767 -3528
<< mimcap >>
rect -5688 5560 -3688 5600
rect -5688 3640 -5648 5560
rect -3728 3640 -3688 5560
rect -5688 3600 -3688 3640
rect -3369 5560 -1369 5600
rect -3369 3640 -3329 5560
rect -1409 3640 -1369 5560
rect -3369 3600 -1369 3640
rect -1050 5560 950 5600
rect -1050 3640 -1010 5560
rect 910 3640 950 5560
rect -1050 3600 950 3640
rect 1269 5560 3269 5600
rect 1269 3640 1309 5560
rect 3229 3640 3269 5560
rect 1269 3600 3269 3640
rect 3588 5560 5588 5600
rect 3588 3640 3628 5560
rect 5548 3640 5588 5560
rect 3588 3600 5588 3640
rect -5688 3260 -3688 3300
rect -5688 1340 -5648 3260
rect -3728 1340 -3688 3260
rect -5688 1300 -3688 1340
rect -3369 3260 -1369 3300
rect -3369 1340 -3329 3260
rect -1409 1340 -1369 3260
rect -3369 1300 -1369 1340
rect -1050 3260 950 3300
rect -1050 1340 -1010 3260
rect 910 1340 950 3260
rect -1050 1300 950 1340
rect 1269 3260 3269 3300
rect 1269 1340 1309 3260
rect 3229 1340 3269 3260
rect 1269 1300 3269 1340
rect 3588 3260 5588 3300
rect 3588 1340 3628 3260
rect 5548 1340 5588 3260
rect 3588 1300 5588 1340
rect -5688 960 -3688 1000
rect -5688 -960 -5648 960
rect -3728 -960 -3688 960
rect -5688 -1000 -3688 -960
rect -3369 960 -1369 1000
rect -3369 -960 -3329 960
rect -1409 -960 -1369 960
rect -3369 -1000 -1369 -960
rect -1050 960 950 1000
rect -1050 -960 -1010 960
rect 910 -960 950 960
rect -1050 -1000 950 -960
rect 1269 960 3269 1000
rect 1269 -960 1309 960
rect 3229 -960 3269 960
rect 1269 -1000 3269 -960
rect 3588 960 5588 1000
rect 3588 -960 3628 960
rect 5548 -960 5588 960
rect 3588 -1000 5588 -960
rect -5688 -1340 -3688 -1300
rect -5688 -3260 -5648 -1340
rect -3728 -3260 -3688 -1340
rect -5688 -3300 -3688 -3260
rect -3369 -1340 -1369 -1300
rect -3369 -3260 -3329 -1340
rect -1409 -3260 -1369 -1340
rect -3369 -3300 -1369 -3260
rect -1050 -1340 950 -1300
rect -1050 -3260 -1010 -1340
rect 910 -3260 950 -1340
rect -1050 -3300 950 -3260
rect 1269 -1340 3269 -1300
rect 1269 -3260 1309 -1340
rect 3229 -3260 3269 -1340
rect 1269 -3300 3269 -3260
rect 3588 -1340 5588 -1300
rect 3588 -3260 3628 -1340
rect 5548 -3260 5588 -1340
rect 3588 -3300 5588 -3260
rect -5688 -3640 -3688 -3600
rect -5688 -5560 -5648 -3640
rect -3728 -5560 -3688 -3640
rect -5688 -5600 -3688 -5560
rect -3369 -3640 -1369 -3600
rect -3369 -5560 -3329 -3640
rect -1409 -5560 -1369 -3640
rect -3369 -5600 -1369 -5560
rect -1050 -3640 950 -3600
rect -1050 -5560 -1010 -3640
rect 910 -5560 950 -3640
rect -1050 -5600 950 -5560
rect 1269 -3640 3269 -3600
rect 1269 -5560 1309 -3640
rect 3229 -5560 3269 -3640
rect 1269 -5600 3269 -5560
rect 3588 -3640 5588 -3600
rect 3588 -5560 3628 -3640
rect 5548 -5560 5588 -3640
rect 3588 -5600 5588 -5560
<< mimcapcontact >>
rect -5648 3640 -3728 5560
rect -3329 3640 -1409 5560
rect -1010 3640 910 5560
rect 1309 3640 3229 5560
rect 3628 3640 5548 5560
rect -5648 1340 -3728 3260
rect -3329 1340 -1409 3260
rect -1010 1340 910 3260
rect 1309 1340 3229 3260
rect 3628 1340 5548 3260
rect -5648 -960 -3728 960
rect -3329 -960 -1409 960
rect -1010 -960 910 960
rect 1309 -960 3229 960
rect 3628 -960 5548 960
rect -5648 -3260 -3728 -1340
rect -3329 -3260 -1409 -1340
rect -1010 -3260 910 -1340
rect 1309 -3260 3229 -1340
rect 3628 -3260 5548 -1340
rect -5648 -5560 -3728 -3640
rect -3329 -5560 -1409 -3640
rect -1010 -5560 910 -3640
rect 1309 -5560 3229 -3640
rect 3628 -5560 5548 -3640
<< metal4 >>
rect -3589 5672 -3493 5688
rect -5649 5560 -3727 5561
rect -5649 3640 -5648 5560
rect -3728 3640 -3727 5560
rect -5649 3639 -3727 3640
rect -3589 3528 -3573 5672
rect -3509 3528 -3493 5672
rect -1270 5672 -1174 5688
rect -3330 5560 -1408 5561
rect -3330 3640 -3329 5560
rect -1409 3640 -1408 5560
rect -3330 3639 -1408 3640
rect -3589 3512 -3493 3528
rect -1270 3528 -1254 5672
rect -1190 3528 -1174 5672
rect 1049 5672 1145 5688
rect -1011 5560 911 5561
rect -1011 3640 -1010 5560
rect 910 3640 911 5560
rect -1011 3639 911 3640
rect -1270 3512 -1174 3528
rect 1049 3528 1065 5672
rect 1129 3528 1145 5672
rect 3368 5672 3464 5688
rect 1308 5560 3230 5561
rect 1308 3640 1309 5560
rect 3229 3640 3230 5560
rect 1308 3639 3230 3640
rect 1049 3512 1145 3528
rect 3368 3528 3384 5672
rect 3448 3528 3464 5672
rect 5687 5672 5783 5688
rect 3627 5560 5549 5561
rect 3627 3640 3628 5560
rect 5548 3640 5549 5560
rect 3627 3639 5549 3640
rect 3368 3512 3464 3528
rect 5687 3528 5703 5672
rect 5767 3528 5783 5672
rect 5687 3512 5783 3528
rect -3589 3372 -3493 3388
rect -5649 3260 -3727 3261
rect -5649 1340 -5648 3260
rect -3728 1340 -3727 3260
rect -5649 1339 -3727 1340
rect -3589 1228 -3573 3372
rect -3509 1228 -3493 3372
rect -1270 3372 -1174 3388
rect -3330 3260 -1408 3261
rect -3330 1340 -3329 3260
rect -1409 1340 -1408 3260
rect -3330 1339 -1408 1340
rect -3589 1212 -3493 1228
rect -1270 1228 -1254 3372
rect -1190 1228 -1174 3372
rect 1049 3372 1145 3388
rect -1011 3260 911 3261
rect -1011 1340 -1010 3260
rect 910 1340 911 3260
rect -1011 1339 911 1340
rect -1270 1212 -1174 1228
rect 1049 1228 1065 3372
rect 1129 1228 1145 3372
rect 3368 3372 3464 3388
rect 1308 3260 3230 3261
rect 1308 1340 1309 3260
rect 3229 1340 3230 3260
rect 1308 1339 3230 1340
rect 1049 1212 1145 1228
rect 3368 1228 3384 3372
rect 3448 1228 3464 3372
rect 5687 3372 5783 3388
rect 3627 3260 5549 3261
rect 3627 1340 3628 3260
rect 5548 1340 5549 3260
rect 3627 1339 5549 1340
rect 3368 1212 3464 1228
rect 5687 1228 5703 3372
rect 5767 1228 5783 3372
rect 5687 1212 5783 1228
rect -3589 1072 -3493 1088
rect -5649 960 -3727 961
rect -5649 -960 -5648 960
rect -3728 -960 -3727 960
rect -5649 -961 -3727 -960
rect -3589 -1072 -3573 1072
rect -3509 -1072 -3493 1072
rect -1270 1072 -1174 1088
rect -3330 960 -1408 961
rect -3330 -960 -3329 960
rect -1409 -960 -1408 960
rect -3330 -961 -1408 -960
rect -3589 -1088 -3493 -1072
rect -1270 -1072 -1254 1072
rect -1190 -1072 -1174 1072
rect 1049 1072 1145 1088
rect -1011 960 911 961
rect -1011 -960 -1010 960
rect 910 -960 911 960
rect -1011 -961 911 -960
rect -1270 -1088 -1174 -1072
rect 1049 -1072 1065 1072
rect 1129 -1072 1145 1072
rect 3368 1072 3464 1088
rect 1308 960 3230 961
rect 1308 -960 1309 960
rect 3229 -960 3230 960
rect 1308 -961 3230 -960
rect 1049 -1088 1145 -1072
rect 3368 -1072 3384 1072
rect 3448 -1072 3464 1072
rect 5687 1072 5783 1088
rect 3627 960 5549 961
rect 3627 -960 3628 960
rect 5548 -960 5549 960
rect 3627 -961 5549 -960
rect 3368 -1088 3464 -1072
rect 5687 -1072 5703 1072
rect 5767 -1072 5783 1072
rect 5687 -1088 5783 -1072
rect -3589 -1228 -3493 -1212
rect -5649 -1340 -3727 -1339
rect -5649 -3260 -5648 -1340
rect -3728 -3260 -3727 -1340
rect -5649 -3261 -3727 -3260
rect -3589 -3372 -3573 -1228
rect -3509 -3372 -3493 -1228
rect -1270 -1228 -1174 -1212
rect -3330 -1340 -1408 -1339
rect -3330 -3260 -3329 -1340
rect -1409 -3260 -1408 -1340
rect -3330 -3261 -1408 -3260
rect -3589 -3388 -3493 -3372
rect -1270 -3372 -1254 -1228
rect -1190 -3372 -1174 -1228
rect 1049 -1228 1145 -1212
rect -1011 -1340 911 -1339
rect -1011 -3260 -1010 -1340
rect 910 -3260 911 -1340
rect -1011 -3261 911 -3260
rect -1270 -3388 -1174 -3372
rect 1049 -3372 1065 -1228
rect 1129 -3372 1145 -1228
rect 3368 -1228 3464 -1212
rect 1308 -1340 3230 -1339
rect 1308 -3260 1309 -1340
rect 3229 -3260 3230 -1340
rect 1308 -3261 3230 -3260
rect 1049 -3388 1145 -3372
rect 3368 -3372 3384 -1228
rect 3448 -3372 3464 -1228
rect 5687 -1228 5783 -1212
rect 3627 -1340 5549 -1339
rect 3627 -3260 3628 -1340
rect 5548 -3260 5549 -1340
rect 3627 -3261 5549 -3260
rect 3368 -3388 3464 -3372
rect 5687 -3372 5703 -1228
rect 5767 -3372 5783 -1228
rect 5687 -3388 5783 -3372
rect -3589 -3528 -3493 -3512
rect -5649 -3640 -3727 -3639
rect -5649 -5560 -5648 -3640
rect -3728 -5560 -3727 -3640
rect -5649 -5561 -3727 -5560
rect -3589 -5672 -3573 -3528
rect -3509 -5672 -3493 -3528
rect -1270 -3528 -1174 -3512
rect -3330 -3640 -1408 -3639
rect -3330 -5560 -3329 -3640
rect -1409 -5560 -1408 -3640
rect -3330 -5561 -1408 -5560
rect -3589 -5688 -3493 -5672
rect -1270 -5672 -1254 -3528
rect -1190 -5672 -1174 -3528
rect 1049 -3528 1145 -3512
rect -1011 -3640 911 -3639
rect -1011 -5560 -1010 -3640
rect 910 -5560 911 -3640
rect -1011 -5561 911 -5560
rect -1270 -5688 -1174 -5672
rect 1049 -5672 1065 -3528
rect 1129 -5672 1145 -3528
rect 3368 -3528 3464 -3512
rect 1308 -3640 3230 -3639
rect 1308 -5560 1309 -3640
rect 3229 -5560 3230 -3640
rect 1308 -5561 3230 -5560
rect 1049 -5688 1145 -5672
rect 3368 -5672 3384 -3528
rect 3448 -5672 3464 -3528
rect 5687 -3528 5783 -3512
rect 3627 -3640 5549 -3639
rect 3627 -5560 3628 -3640
rect 5548 -5560 5549 -3640
rect 3627 -5561 5549 -5560
rect 3368 -5688 3464 -5672
rect 5687 -5672 5703 -3528
rect 5767 -5672 5783 -3528
rect 5687 -5688 5783 -5672
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_1
string FIXED_BBOX 3488 3500 5688 5700
string parameters w 10.00 l 10.00 val 207.6 carea 2.00 cperi 0.19 nx 5 ny 5 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 0 tconnect 0 ccov 100
string library sky130
<< end >>
