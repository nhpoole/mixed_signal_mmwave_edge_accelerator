magic
tech sky130A
magscale 1 2
timestamp 1626065694
<< checkpaint >>
rect 100505 65776 105279 71992
<< metal1 >>
rect 101921 69445 103987 69473
rect 101797 69343 102819 69371
<< metal2 >>
rect 101783 67068 101811 69357
rect 101907 68558 101935 69459
rect 102805 69357 102833 70732
rect 103973 69459 104001 70732
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_0
timestamp 1626065694
transform 1 0 103955 0 1 69427
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_1
timestamp 1626065694
transform 1 0 101889 0 1 68526
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_2
timestamp 1626065694
transform 1 0 101889 0 1 69427
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_3
timestamp 1626065694
transform 1 0 102787 0 1 69325
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_4
timestamp 1626065694
transform 1 0 101765 0 1 67036
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_5
timestamp 1626065694
transform 1 0 101765 0 1 69325
box 0 0 64 64
<< properties >>
string FIXED_BBOX 101765 67036 104019 70732
<< end >>
