magic
tech sky130A
magscale 1 2
timestamp 1624494425
<< nwell >>
rect 428 0 760 490
<< poly >>
rect 77 155 136 185
rect 260 155 456 185
<< locali >>
rect 60 137 94 203
rect 165 103 742 137
<< metal1 >>
rect 184 0 212 395
rect 580 0 608 395
use contact_7  contact_7_0
timestamp 1624494425
transform 1 0 565 0 1 187
box 0 0 58 66
use contact_7  contact_7_1
timestamp 1624494425
transform 1 0 169 0 1 187
box 0 0 58 66
use contact_15  contact_15_0
timestamp 1624494425
transform 1 0 44 0 1 137
box 0 0 66 66
use contact_7  contact_7_2
timestamp 1624494425
transform 1 0 169 0 1 362
box 0 0 58 66
use contact_14  contact_14_0
timestamp 1624494425
transform 1 0 173 0 1 354
box -26 -26 76 108
use contact_7  contact_7_3
timestamp 1624494425
transform 1 0 565 0 1 362
box 0 0 58 66
use contact_13  contact_13_0
timestamp 1624494425
transform 1 0 569 0 1 354
box -59 -43 109 125
use nmos_m1_w0_360_sli_dli_da_p  nmos_m1_w0_360_sli_dli_da_p_0
timestamp 1624494425
transform 0 1 162 -1 0 245
box -26 -26 176 98
use pmos_m1_w1_120_sli_dli_da_p  pmos_m1_w1_120_sli_dli_da_p_0
timestamp 1624494425
transform 0 1 482 -1 0 245
box -59 -54 209 278
<< labels >>
rlabel locali s 77 170 77 170 4 A
rlabel locali s 453 120 453 120 4 Z
rlabel metal1 s 184 0 212 395 4 gnd
rlabel metal1 s 580 0 608 395 4 vdd
<< properties >>
string FIXED_BBOX 0 0 742 395
<< end >>
