magic
tech sky130A
magscale 1 2
timestamp 1626065694
<< checkpaint >>
rect -1787 -1386 1787 1386
<< pwell >>
rect -527 -126 527 126
<< nmos >>
rect -443 -100 -383 100
rect -325 -100 -265 100
rect -207 -100 -147 100
rect -89 -100 -29 100
rect 29 -100 89 100
rect 147 -100 207 100
rect 265 -100 325 100
rect 383 -100 443 100
<< ndiff >>
rect -501 85 -443 100
rect -501 51 -489 85
rect -455 51 -443 85
rect -501 17 -443 51
rect -501 -17 -489 17
rect -455 -17 -443 17
rect -501 -51 -443 -17
rect -501 -85 -489 -51
rect -455 -85 -443 -51
rect -501 -100 -443 -85
rect -383 85 -325 100
rect -383 51 -371 85
rect -337 51 -325 85
rect -383 17 -325 51
rect -383 -17 -371 17
rect -337 -17 -325 17
rect -383 -51 -325 -17
rect -383 -85 -371 -51
rect -337 -85 -325 -51
rect -383 -100 -325 -85
rect -265 85 -207 100
rect -265 51 -253 85
rect -219 51 -207 85
rect -265 17 -207 51
rect -265 -17 -253 17
rect -219 -17 -207 17
rect -265 -51 -207 -17
rect -265 -85 -253 -51
rect -219 -85 -207 -51
rect -265 -100 -207 -85
rect -147 85 -89 100
rect -147 51 -135 85
rect -101 51 -89 85
rect -147 17 -89 51
rect -147 -17 -135 17
rect -101 -17 -89 17
rect -147 -51 -89 -17
rect -147 -85 -135 -51
rect -101 -85 -89 -51
rect -147 -100 -89 -85
rect -29 85 29 100
rect -29 51 -17 85
rect 17 51 29 85
rect -29 17 29 51
rect -29 -17 -17 17
rect 17 -17 29 17
rect -29 -51 29 -17
rect -29 -85 -17 -51
rect 17 -85 29 -51
rect -29 -100 29 -85
rect 89 85 147 100
rect 89 51 101 85
rect 135 51 147 85
rect 89 17 147 51
rect 89 -17 101 17
rect 135 -17 147 17
rect 89 -51 147 -17
rect 89 -85 101 -51
rect 135 -85 147 -51
rect 89 -100 147 -85
rect 207 85 265 100
rect 207 51 219 85
rect 253 51 265 85
rect 207 17 265 51
rect 207 -17 219 17
rect 253 -17 265 17
rect 207 -51 265 -17
rect 207 -85 219 -51
rect 253 -85 265 -51
rect 207 -100 265 -85
rect 325 85 383 100
rect 325 51 337 85
rect 371 51 383 85
rect 325 17 383 51
rect 325 -17 337 17
rect 371 -17 383 17
rect 325 -51 383 -17
rect 325 -85 337 -51
rect 371 -85 383 -51
rect 325 -100 383 -85
rect 443 85 501 100
rect 443 51 455 85
rect 489 51 501 85
rect 443 17 501 51
rect 443 -17 455 17
rect 489 -17 501 17
rect 443 -51 501 -17
rect 443 -85 455 -51
rect 489 -85 501 -51
rect 443 -100 501 -85
<< ndiffc >>
rect -489 51 -455 85
rect -489 -17 -455 17
rect -489 -85 -455 -51
rect -371 51 -337 85
rect -371 -17 -337 17
rect -371 -85 -337 -51
rect -253 51 -219 85
rect -253 -17 -219 17
rect -253 -85 -219 -51
rect -135 51 -101 85
rect -135 -17 -101 17
rect -135 -85 -101 -51
rect -17 51 17 85
rect -17 -17 17 17
rect -17 -85 17 -51
rect 101 51 135 85
rect 101 -17 135 17
rect 101 -85 135 -51
rect 219 51 253 85
rect 219 -17 253 17
rect 219 -85 253 -51
rect 337 51 371 85
rect 337 -17 371 17
rect 337 -85 371 -51
rect 455 51 489 85
rect 455 -17 489 17
rect 455 -85 489 -51
<< poly >>
rect -443 100 -383 126
rect -325 100 -265 126
rect -207 100 -147 126
rect -89 100 -29 126
rect 29 100 89 126
rect 147 100 207 126
rect 265 100 325 126
rect 383 100 443 126
rect -443 -126 -383 -100
rect -325 -126 -265 -100
rect -207 -126 -147 -100
rect -89 -126 -29 -100
rect 29 -126 89 -100
rect 147 -126 207 -100
rect 265 -126 325 -100
rect 383 -126 443 -100
<< locali >>
rect -489 85 -455 104
rect -489 17 -455 19
rect -489 -19 -455 -17
rect -489 -104 -455 -85
rect -371 85 -337 104
rect -371 17 -337 19
rect -371 -19 -337 -17
rect -371 -104 -337 -85
rect -253 85 -219 104
rect -253 17 -219 19
rect -253 -19 -219 -17
rect -253 -104 -219 -85
rect -135 85 -101 104
rect -135 17 -101 19
rect -135 -19 -101 -17
rect -135 -104 -101 -85
rect -17 85 17 104
rect -17 17 17 19
rect -17 -19 17 -17
rect -17 -104 17 -85
rect 101 85 135 104
rect 101 17 135 19
rect 101 -19 135 -17
rect 101 -104 135 -85
rect 219 85 253 104
rect 219 17 253 19
rect 219 -19 253 -17
rect 219 -104 253 -85
rect 337 85 371 104
rect 337 17 371 19
rect 337 -19 371 -17
rect 337 -104 371 -85
rect 455 85 489 104
rect 455 17 489 19
rect 455 -19 489 -17
rect 455 -104 489 -85
<< viali >>
rect -489 51 -455 53
rect -489 19 -455 51
rect -489 -51 -455 -19
rect -489 -53 -455 -51
rect -371 51 -337 53
rect -371 19 -337 51
rect -371 -51 -337 -19
rect -371 -53 -337 -51
rect -253 51 -219 53
rect -253 19 -219 51
rect -253 -51 -219 -19
rect -253 -53 -219 -51
rect -135 51 -101 53
rect -135 19 -101 51
rect -135 -51 -101 -19
rect -135 -53 -101 -51
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect 101 51 135 53
rect 101 19 135 51
rect 101 -51 135 -19
rect 101 -53 135 -51
rect 219 51 253 53
rect 219 19 253 51
rect 219 -51 253 -19
rect 219 -53 253 -51
rect 337 51 371 53
rect 337 19 371 51
rect 337 -51 371 -19
rect 337 -53 371 -51
rect 455 51 489 53
rect 455 19 489 51
rect 455 -51 489 -19
rect 455 -53 489 -51
<< metal1 >>
rect -495 53 -449 100
rect -495 19 -489 53
rect -455 19 -449 53
rect -495 -19 -449 19
rect -495 -53 -489 -19
rect -455 -53 -449 -19
rect -495 -100 -449 -53
rect -377 53 -331 100
rect -377 19 -371 53
rect -337 19 -331 53
rect -377 -19 -331 19
rect -377 -53 -371 -19
rect -337 -53 -331 -19
rect -377 -100 -331 -53
rect -259 53 -213 100
rect -259 19 -253 53
rect -219 19 -213 53
rect -259 -19 -213 19
rect -259 -53 -253 -19
rect -219 -53 -213 -19
rect -259 -100 -213 -53
rect -141 53 -95 100
rect -141 19 -135 53
rect -101 19 -95 53
rect -141 -19 -95 19
rect -141 -53 -135 -19
rect -101 -53 -95 -19
rect -141 -100 -95 -53
rect -23 53 23 100
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -100 23 -53
rect 95 53 141 100
rect 95 19 101 53
rect 135 19 141 53
rect 95 -19 141 19
rect 95 -53 101 -19
rect 135 -53 141 -19
rect 95 -100 141 -53
rect 213 53 259 100
rect 213 19 219 53
rect 253 19 259 53
rect 213 -19 259 19
rect 213 -53 219 -19
rect 253 -53 259 -19
rect 213 -100 259 -53
rect 331 53 377 100
rect 331 19 337 53
rect 371 19 377 53
rect 331 -19 377 19
rect 331 -53 337 -19
rect 371 -53 377 -19
rect 331 -100 377 -53
rect 449 53 495 100
rect 449 19 455 53
rect 489 19 495 53
rect 449 -19 495 19
rect 449 -53 455 -19
rect 489 -53 495 -19
rect 449 -100 495 -53
<< end >>
