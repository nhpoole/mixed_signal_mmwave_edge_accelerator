magic
tech sky130A
magscale 1 2
timestamp 1626065694
<< checkpaint >>
rect -2954 -1648 2954 1648
<< pwell >>
rect -1694 -326 1694 326
<< nmoslvt >>
rect -1610 -300 -1370 300
rect -1312 -300 -1072 300
rect -1014 -300 -774 300
rect -716 -300 -476 300
rect -418 -300 -178 300
rect -120 -300 120 300
rect 178 -300 418 300
rect 476 -300 716 300
rect 774 -300 1014 300
rect 1072 -300 1312 300
rect 1370 -300 1610 300
<< ndiff >>
rect -1668 255 -1610 300
rect -1668 221 -1656 255
rect -1622 221 -1610 255
rect -1668 187 -1610 221
rect -1668 153 -1656 187
rect -1622 153 -1610 187
rect -1668 119 -1610 153
rect -1668 85 -1656 119
rect -1622 85 -1610 119
rect -1668 51 -1610 85
rect -1668 17 -1656 51
rect -1622 17 -1610 51
rect -1668 -17 -1610 17
rect -1668 -51 -1656 -17
rect -1622 -51 -1610 -17
rect -1668 -85 -1610 -51
rect -1668 -119 -1656 -85
rect -1622 -119 -1610 -85
rect -1668 -153 -1610 -119
rect -1668 -187 -1656 -153
rect -1622 -187 -1610 -153
rect -1668 -221 -1610 -187
rect -1668 -255 -1656 -221
rect -1622 -255 -1610 -221
rect -1668 -300 -1610 -255
rect -1370 255 -1312 300
rect -1370 221 -1358 255
rect -1324 221 -1312 255
rect -1370 187 -1312 221
rect -1370 153 -1358 187
rect -1324 153 -1312 187
rect -1370 119 -1312 153
rect -1370 85 -1358 119
rect -1324 85 -1312 119
rect -1370 51 -1312 85
rect -1370 17 -1358 51
rect -1324 17 -1312 51
rect -1370 -17 -1312 17
rect -1370 -51 -1358 -17
rect -1324 -51 -1312 -17
rect -1370 -85 -1312 -51
rect -1370 -119 -1358 -85
rect -1324 -119 -1312 -85
rect -1370 -153 -1312 -119
rect -1370 -187 -1358 -153
rect -1324 -187 -1312 -153
rect -1370 -221 -1312 -187
rect -1370 -255 -1358 -221
rect -1324 -255 -1312 -221
rect -1370 -300 -1312 -255
rect -1072 255 -1014 300
rect -1072 221 -1060 255
rect -1026 221 -1014 255
rect -1072 187 -1014 221
rect -1072 153 -1060 187
rect -1026 153 -1014 187
rect -1072 119 -1014 153
rect -1072 85 -1060 119
rect -1026 85 -1014 119
rect -1072 51 -1014 85
rect -1072 17 -1060 51
rect -1026 17 -1014 51
rect -1072 -17 -1014 17
rect -1072 -51 -1060 -17
rect -1026 -51 -1014 -17
rect -1072 -85 -1014 -51
rect -1072 -119 -1060 -85
rect -1026 -119 -1014 -85
rect -1072 -153 -1014 -119
rect -1072 -187 -1060 -153
rect -1026 -187 -1014 -153
rect -1072 -221 -1014 -187
rect -1072 -255 -1060 -221
rect -1026 -255 -1014 -221
rect -1072 -300 -1014 -255
rect -774 255 -716 300
rect -774 221 -762 255
rect -728 221 -716 255
rect -774 187 -716 221
rect -774 153 -762 187
rect -728 153 -716 187
rect -774 119 -716 153
rect -774 85 -762 119
rect -728 85 -716 119
rect -774 51 -716 85
rect -774 17 -762 51
rect -728 17 -716 51
rect -774 -17 -716 17
rect -774 -51 -762 -17
rect -728 -51 -716 -17
rect -774 -85 -716 -51
rect -774 -119 -762 -85
rect -728 -119 -716 -85
rect -774 -153 -716 -119
rect -774 -187 -762 -153
rect -728 -187 -716 -153
rect -774 -221 -716 -187
rect -774 -255 -762 -221
rect -728 -255 -716 -221
rect -774 -300 -716 -255
rect -476 255 -418 300
rect -476 221 -464 255
rect -430 221 -418 255
rect -476 187 -418 221
rect -476 153 -464 187
rect -430 153 -418 187
rect -476 119 -418 153
rect -476 85 -464 119
rect -430 85 -418 119
rect -476 51 -418 85
rect -476 17 -464 51
rect -430 17 -418 51
rect -476 -17 -418 17
rect -476 -51 -464 -17
rect -430 -51 -418 -17
rect -476 -85 -418 -51
rect -476 -119 -464 -85
rect -430 -119 -418 -85
rect -476 -153 -418 -119
rect -476 -187 -464 -153
rect -430 -187 -418 -153
rect -476 -221 -418 -187
rect -476 -255 -464 -221
rect -430 -255 -418 -221
rect -476 -300 -418 -255
rect -178 255 -120 300
rect -178 221 -166 255
rect -132 221 -120 255
rect -178 187 -120 221
rect -178 153 -166 187
rect -132 153 -120 187
rect -178 119 -120 153
rect -178 85 -166 119
rect -132 85 -120 119
rect -178 51 -120 85
rect -178 17 -166 51
rect -132 17 -120 51
rect -178 -17 -120 17
rect -178 -51 -166 -17
rect -132 -51 -120 -17
rect -178 -85 -120 -51
rect -178 -119 -166 -85
rect -132 -119 -120 -85
rect -178 -153 -120 -119
rect -178 -187 -166 -153
rect -132 -187 -120 -153
rect -178 -221 -120 -187
rect -178 -255 -166 -221
rect -132 -255 -120 -221
rect -178 -300 -120 -255
rect 120 255 178 300
rect 120 221 132 255
rect 166 221 178 255
rect 120 187 178 221
rect 120 153 132 187
rect 166 153 178 187
rect 120 119 178 153
rect 120 85 132 119
rect 166 85 178 119
rect 120 51 178 85
rect 120 17 132 51
rect 166 17 178 51
rect 120 -17 178 17
rect 120 -51 132 -17
rect 166 -51 178 -17
rect 120 -85 178 -51
rect 120 -119 132 -85
rect 166 -119 178 -85
rect 120 -153 178 -119
rect 120 -187 132 -153
rect 166 -187 178 -153
rect 120 -221 178 -187
rect 120 -255 132 -221
rect 166 -255 178 -221
rect 120 -300 178 -255
rect 418 255 476 300
rect 418 221 430 255
rect 464 221 476 255
rect 418 187 476 221
rect 418 153 430 187
rect 464 153 476 187
rect 418 119 476 153
rect 418 85 430 119
rect 464 85 476 119
rect 418 51 476 85
rect 418 17 430 51
rect 464 17 476 51
rect 418 -17 476 17
rect 418 -51 430 -17
rect 464 -51 476 -17
rect 418 -85 476 -51
rect 418 -119 430 -85
rect 464 -119 476 -85
rect 418 -153 476 -119
rect 418 -187 430 -153
rect 464 -187 476 -153
rect 418 -221 476 -187
rect 418 -255 430 -221
rect 464 -255 476 -221
rect 418 -300 476 -255
rect 716 255 774 300
rect 716 221 728 255
rect 762 221 774 255
rect 716 187 774 221
rect 716 153 728 187
rect 762 153 774 187
rect 716 119 774 153
rect 716 85 728 119
rect 762 85 774 119
rect 716 51 774 85
rect 716 17 728 51
rect 762 17 774 51
rect 716 -17 774 17
rect 716 -51 728 -17
rect 762 -51 774 -17
rect 716 -85 774 -51
rect 716 -119 728 -85
rect 762 -119 774 -85
rect 716 -153 774 -119
rect 716 -187 728 -153
rect 762 -187 774 -153
rect 716 -221 774 -187
rect 716 -255 728 -221
rect 762 -255 774 -221
rect 716 -300 774 -255
rect 1014 255 1072 300
rect 1014 221 1026 255
rect 1060 221 1072 255
rect 1014 187 1072 221
rect 1014 153 1026 187
rect 1060 153 1072 187
rect 1014 119 1072 153
rect 1014 85 1026 119
rect 1060 85 1072 119
rect 1014 51 1072 85
rect 1014 17 1026 51
rect 1060 17 1072 51
rect 1014 -17 1072 17
rect 1014 -51 1026 -17
rect 1060 -51 1072 -17
rect 1014 -85 1072 -51
rect 1014 -119 1026 -85
rect 1060 -119 1072 -85
rect 1014 -153 1072 -119
rect 1014 -187 1026 -153
rect 1060 -187 1072 -153
rect 1014 -221 1072 -187
rect 1014 -255 1026 -221
rect 1060 -255 1072 -221
rect 1014 -300 1072 -255
rect 1312 255 1370 300
rect 1312 221 1324 255
rect 1358 221 1370 255
rect 1312 187 1370 221
rect 1312 153 1324 187
rect 1358 153 1370 187
rect 1312 119 1370 153
rect 1312 85 1324 119
rect 1358 85 1370 119
rect 1312 51 1370 85
rect 1312 17 1324 51
rect 1358 17 1370 51
rect 1312 -17 1370 17
rect 1312 -51 1324 -17
rect 1358 -51 1370 -17
rect 1312 -85 1370 -51
rect 1312 -119 1324 -85
rect 1358 -119 1370 -85
rect 1312 -153 1370 -119
rect 1312 -187 1324 -153
rect 1358 -187 1370 -153
rect 1312 -221 1370 -187
rect 1312 -255 1324 -221
rect 1358 -255 1370 -221
rect 1312 -300 1370 -255
rect 1610 255 1668 300
rect 1610 221 1622 255
rect 1656 221 1668 255
rect 1610 187 1668 221
rect 1610 153 1622 187
rect 1656 153 1668 187
rect 1610 119 1668 153
rect 1610 85 1622 119
rect 1656 85 1668 119
rect 1610 51 1668 85
rect 1610 17 1622 51
rect 1656 17 1668 51
rect 1610 -17 1668 17
rect 1610 -51 1622 -17
rect 1656 -51 1668 -17
rect 1610 -85 1668 -51
rect 1610 -119 1622 -85
rect 1656 -119 1668 -85
rect 1610 -153 1668 -119
rect 1610 -187 1622 -153
rect 1656 -187 1668 -153
rect 1610 -221 1668 -187
rect 1610 -255 1622 -221
rect 1656 -255 1668 -221
rect 1610 -300 1668 -255
<< ndiffc >>
rect -1656 221 -1622 255
rect -1656 153 -1622 187
rect -1656 85 -1622 119
rect -1656 17 -1622 51
rect -1656 -51 -1622 -17
rect -1656 -119 -1622 -85
rect -1656 -187 -1622 -153
rect -1656 -255 -1622 -221
rect -1358 221 -1324 255
rect -1358 153 -1324 187
rect -1358 85 -1324 119
rect -1358 17 -1324 51
rect -1358 -51 -1324 -17
rect -1358 -119 -1324 -85
rect -1358 -187 -1324 -153
rect -1358 -255 -1324 -221
rect -1060 221 -1026 255
rect -1060 153 -1026 187
rect -1060 85 -1026 119
rect -1060 17 -1026 51
rect -1060 -51 -1026 -17
rect -1060 -119 -1026 -85
rect -1060 -187 -1026 -153
rect -1060 -255 -1026 -221
rect -762 221 -728 255
rect -762 153 -728 187
rect -762 85 -728 119
rect -762 17 -728 51
rect -762 -51 -728 -17
rect -762 -119 -728 -85
rect -762 -187 -728 -153
rect -762 -255 -728 -221
rect -464 221 -430 255
rect -464 153 -430 187
rect -464 85 -430 119
rect -464 17 -430 51
rect -464 -51 -430 -17
rect -464 -119 -430 -85
rect -464 -187 -430 -153
rect -464 -255 -430 -221
rect -166 221 -132 255
rect -166 153 -132 187
rect -166 85 -132 119
rect -166 17 -132 51
rect -166 -51 -132 -17
rect -166 -119 -132 -85
rect -166 -187 -132 -153
rect -166 -255 -132 -221
rect 132 221 166 255
rect 132 153 166 187
rect 132 85 166 119
rect 132 17 166 51
rect 132 -51 166 -17
rect 132 -119 166 -85
rect 132 -187 166 -153
rect 132 -255 166 -221
rect 430 221 464 255
rect 430 153 464 187
rect 430 85 464 119
rect 430 17 464 51
rect 430 -51 464 -17
rect 430 -119 464 -85
rect 430 -187 464 -153
rect 430 -255 464 -221
rect 728 221 762 255
rect 728 153 762 187
rect 728 85 762 119
rect 728 17 762 51
rect 728 -51 762 -17
rect 728 -119 762 -85
rect 728 -187 762 -153
rect 728 -255 762 -221
rect 1026 221 1060 255
rect 1026 153 1060 187
rect 1026 85 1060 119
rect 1026 17 1060 51
rect 1026 -51 1060 -17
rect 1026 -119 1060 -85
rect 1026 -187 1060 -153
rect 1026 -255 1060 -221
rect 1324 221 1358 255
rect 1324 153 1358 187
rect 1324 85 1358 119
rect 1324 17 1358 51
rect 1324 -51 1358 -17
rect 1324 -119 1358 -85
rect 1324 -187 1358 -153
rect 1324 -255 1358 -221
rect 1622 221 1656 255
rect 1622 153 1656 187
rect 1622 85 1656 119
rect 1622 17 1656 51
rect 1622 -51 1656 -17
rect 1622 -119 1656 -85
rect 1622 -187 1656 -153
rect 1622 -255 1656 -221
<< poly >>
rect -1568 372 -1412 388
rect -1568 355 -1541 372
rect -1610 338 -1541 355
rect -1507 338 -1473 372
rect -1439 355 -1412 372
rect -1270 372 -1114 388
rect -1270 355 -1243 372
rect -1439 338 -1370 355
rect -1610 300 -1370 338
rect -1312 338 -1243 355
rect -1209 338 -1175 372
rect -1141 355 -1114 372
rect -972 372 -816 388
rect -972 355 -945 372
rect -1141 338 -1072 355
rect -1312 300 -1072 338
rect -1014 338 -945 355
rect -911 338 -877 372
rect -843 355 -816 372
rect -674 372 -518 388
rect -674 355 -647 372
rect -843 338 -774 355
rect -1014 300 -774 338
rect -716 338 -647 355
rect -613 338 -579 372
rect -545 355 -518 372
rect -376 372 -220 388
rect -376 355 -349 372
rect -545 338 -476 355
rect -716 300 -476 338
rect -418 338 -349 355
rect -315 338 -281 372
rect -247 355 -220 372
rect -78 372 78 388
rect -78 355 -51 372
rect -247 338 -178 355
rect -418 300 -178 338
rect -120 338 -51 355
rect -17 338 17 372
rect 51 355 78 372
rect 220 372 376 388
rect 220 355 247 372
rect 51 338 120 355
rect -120 300 120 338
rect 178 338 247 355
rect 281 338 315 372
rect 349 355 376 372
rect 518 372 674 388
rect 518 355 545 372
rect 349 338 418 355
rect 178 300 418 338
rect 476 338 545 355
rect 579 338 613 372
rect 647 355 674 372
rect 816 372 972 388
rect 816 355 843 372
rect 647 338 716 355
rect 476 300 716 338
rect 774 338 843 355
rect 877 338 911 372
rect 945 355 972 372
rect 1114 372 1270 388
rect 1114 355 1141 372
rect 945 338 1014 355
rect 774 300 1014 338
rect 1072 338 1141 355
rect 1175 338 1209 372
rect 1243 355 1270 372
rect 1412 372 1568 388
rect 1412 355 1439 372
rect 1243 338 1312 355
rect 1072 300 1312 338
rect 1370 338 1439 355
rect 1473 338 1507 372
rect 1541 355 1568 372
rect 1541 338 1610 355
rect 1370 300 1610 338
rect -1610 -338 -1370 -300
rect -1610 -355 -1541 -338
rect -1568 -372 -1541 -355
rect -1507 -372 -1473 -338
rect -1439 -355 -1370 -338
rect -1312 -338 -1072 -300
rect -1312 -355 -1243 -338
rect -1439 -372 -1412 -355
rect -1568 -388 -1412 -372
rect -1270 -372 -1243 -355
rect -1209 -372 -1175 -338
rect -1141 -355 -1072 -338
rect -1014 -338 -774 -300
rect -1014 -355 -945 -338
rect -1141 -372 -1114 -355
rect -1270 -388 -1114 -372
rect -972 -372 -945 -355
rect -911 -372 -877 -338
rect -843 -355 -774 -338
rect -716 -338 -476 -300
rect -716 -355 -647 -338
rect -843 -372 -816 -355
rect -972 -388 -816 -372
rect -674 -372 -647 -355
rect -613 -372 -579 -338
rect -545 -355 -476 -338
rect -418 -338 -178 -300
rect -418 -355 -349 -338
rect -545 -372 -518 -355
rect -674 -388 -518 -372
rect -376 -372 -349 -355
rect -315 -372 -281 -338
rect -247 -355 -178 -338
rect -120 -338 120 -300
rect -120 -355 -51 -338
rect -247 -372 -220 -355
rect -376 -388 -220 -372
rect -78 -372 -51 -355
rect -17 -372 17 -338
rect 51 -355 120 -338
rect 178 -338 418 -300
rect 178 -355 247 -338
rect 51 -372 78 -355
rect -78 -388 78 -372
rect 220 -372 247 -355
rect 281 -372 315 -338
rect 349 -355 418 -338
rect 476 -338 716 -300
rect 476 -355 545 -338
rect 349 -372 376 -355
rect 220 -388 376 -372
rect 518 -372 545 -355
rect 579 -372 613 -338
rect 647 -355 716 -338
rect 774 -338 1014 -300
rect 774 -355 843 -338
rect 647 -372 674 -355
rect 518 -388 674 -372
rect 816 -372 843 -355
rect 877 -372 911 -338
rect 945 -355 1014 -338
rect 1072 -338 1312 -300
rect 1072 -355 1141 -338
rect 945 -372 972 -355
rect 816 -388 972 -372
rect 1114 -372 1141 -355
rect 1175 -372 1209 -338
rect 1243 -355 1312 -338
rect 1370 -338 1610 -300
rect 1370 -355 1439 -338
rect 1243 -372 1270 -355
rect 1114 -388 1270 -372
rect 1412 -372 1439 -355
rect 1473 -372 1507 -338
rect 1541 -355 1610 -338
rect 1541 -372 1568 -355
rect 1412 -388 1568 -372
<< polycont >>
rect -1541 338 -1507 372
rect -1473 338 -1439 372
rect -1243 338 -1209 372
rect -1175 338 -1141 372
rect -945 338 -911 372
rect -877 338 -843 372
rect -647 338 -613 372
rect -579 338 -545 372
rect -349 338 -315 372
rect -281 338 -247 372
rect -51 338 -17 372
rect 17 338 51 372
rect 247 338 281 372
rect 315 338 349 372
rect 545 338 579 372
rect 613 338 647 372
rect 843 338 877 372
rect 911 338 945 372
rect 1141 338 1175 372
rect 1209 338 1243 372
rect 1439 338 1473 372
rect 1507 338 1541 372
rect -1541 -372 -1507 -338
rect -1473 -372 -1439 -338
rect -1243 -372 -1209 -338
rect -1175 -372 -1141 -338
rect -945 -372 -911 -338
rect -877 -372 -843 -338
rect -647 -372 -613 -338
rect -579 -372 -545 -338
rect -349 -372 -315 -338
rect -281 -372 -247 -338
rect -51 -372 -17 -338
rect 17 -372 51 -338
rect 247 -372 281 -338
rect 315 -372 349 -338
rect 545 -372 579 -338
rect 613 -372 647 -338
rect 843 -372 877 -338
rect 911 -372 945 -338
rect 1141 -372 1175 -338
rect 1209 -372 1243 -338
rect 1439 -372 1473 -338
rect 1507 -372 1541 -338
<< locali >>
rect -1568 338 -1541 372
rect -1439 338 -1412 372
rect -1270 338 -1243 372
rect -1141 338 -1114 372
rect -972 338 -945 372
rect -843 338 -816 372
rect -674 338 -647 372
rect -545 338 -518 372
rect -376 338 -349 372
rect -247 338 -220 372
rect -78 338 -51 372
rect 51 338 78 372
rect 220 338 247 372
rect 349 338 376 372
rect 518 338 545 372
rect 647 338 674 372
rect 816 338 843 372
rect 945 338 972 372
rect 1114 338 1141 372
rect 1243 338 1270 372
rect 1412 338 1439 372
rect 1541 338 1568 372
rect -1656 269 -1622 304
rect -1656 197 -1622 221
rect -1656 125 -1622 153
rect -1656 53 -1622 85
rect -1656 -17 -1622 17
rect -1656 -85 -1622 -53
rect -1656 -153 -1622 -125
rect -1656 -221 -1622 -197
rect -1656 -304 -1622 -269
rect -1358 269 -1324 304
rect -1358 197 -1324 221
rect -1358 125 -1324 153
rect -1358 53 -1324 85
rect -1358 -17 -1324 17
rect -1358 -85 -1324 -53
rect -1358 -153 -1324 -125
rect -1358 -221 -1324 -197
rect -1358 -304 -1324 -269
rect -1060 269 -1026 304
rect -1060 197 -1026 221
rect -1060 125 -1026 153
rect -1060 53 -1026 85
rect -1060 -17 -1026 17
rect -1060 -85 -1026 -53
rect -1060 -153 -1026 -125
rect -1060 -221 -1026 -197
rect -1060 -304 -1026 -269
rect -762 269 -728 304
rect -762 197 -728 221
rect -762 125 -728 153
rect -762 53 -728 85
rect -762 -17 -728 17
rect -762 -85 -728 -53
rect -762 -153 -728 -125
rect -762 -221 -728 -197
rect -762 -304 -728 -269
rect -464 269 -430 304
rect -464 197 -430 221
rect -464 125 -430 153
rect -464 53 -430 85
rect -464 -17 -430 17
rect -464 -85 -430 -53
rect -464 -153 -430 -125
rect -464 -221 -430 -197
rect -464 -304 -430 -269
rect -166 269 -132 304
rect -166 197 -132 221
rect -166 125 -132 153
rect -166 53 -132 85
rect -166 -17 -132 17
rect -166 -85 -132 -53
rect -166 -153 -132 -125
rect -166 -221 -132 -197
rect -166 -304 -132 -269
rect 132 269 166 304
rect 132 197 166 221
rect 132 125 166 153
rect 132 53 166 85
rect 132 -17 166 17
rect 132 -85 166 -53
rect 132 -153 166 -125
rect 132 -221 166 -197
rect 132 -304 166 -269
rect 430 269 464 304
rect 430 197 464 221
rect 430 125 464 153
rect 430 53 464 85
rect 430 -17 464 17
rect 430 -85 464 -53
rect 430 -153 464 -125
rect 430 -221 464 -197
rect 430 -304 464 -269
rect 728 269 762 304
rect 728 197 762 221
rect 728 125 762 153
rect 728 53 762 85
rect 728 -17 762 17
rect 728 -85 762 -53
rect 728 -153 762 -125
rect 728 -221 762 -197
rect 728 -304 762 -269
rect 1026 269 1060 304
rect 1026 197 1060 221
rect 1026 125 1060 153
rect 1026 53 1060 85
rect 1026 -17 1060 17
rect 1026 -85 1060 -53
rect 1026 -153 1060 -125
rect 1026 -221 1060 -197
rect 1026 -304 1060 -269
rect 1324 269 1358 304
rect 1324 197 1358 221
rect 1324 125 1358 153
rect 1324 53 1358 85
rect 1324 -17 1358 17
rect 1324 -85 1358 -53
rect 1324 -153 1358 -125
rect 1324 -221 1358 -197
rect 1324 -304 1358 -269
rect 1622 269 1656 304
rect 1622 197 1656 221
rect 1622 125 1656 153
rect 1622 53 1656 85
rect 1622 -17 1656 17
rect 1622 -85 1656 -53
rect 1622 -153 1656 -125
rect 1622 -221 1656 -197
rect 1622 -304 1656 -269
rect -1568 -372 -1541 -338
rect -1439 -372 -1412 -338
rect -1270 -372 -1243 -338
rect -1141 -372 -1114 -338
rect -972 -372 -945 -338
rect -843 -372 -816 -338
rect -674 -372 -647 -338
rect -545 -372 -518 -338
rect -376 -372 -349 -338
rect -247 -372 -220 -338
rect -78 -372 -51 -338
rect 51 -372 78 -338
rect 220 -372 247 -338
rect 349 -372 376 -338
rect 518 -372 545 -338
rect 647 -372 674 -338
rect 816 -372 843 -338
rect 945 -372 972 -338
rect 1114 -372 1141 -338
rect 1243 -372 1270 -338
rect 1412 -372 1439 -338
rect 1541 -372 1568 -338
<< viali >>
rect -1507 338 -1473 372
rect -1209 338 -1175 372
rect -911 338 -877 372
rect -613 338 -579 372
rect -315 338 -281 372
rect -17 338 17 372
rect 281 338 315 372
rect 579 338 613 372
rect 877 338 911 372
rect 1175 338 1209 372
rect 1473 338 1507 372
rect -1656 255 -1622 269
rect -1656 235 -1622 255
rect -1656 187 -1622 197
rect -1656 163 -1622 187
rect -1656 119 -1622 125
rect -1656 91 -1622 119
rect -1656 51 -1622 53
rect -1656 19 -1622 51
rect -1656 -51 -1622 -19
rect -1656 -53 -1622 -51
rect -1656 -119 -1622 -91
rect -1656 -125 -1622 -119
rect -1656 -187 -1622 -163
rect -1656 -197 -1622 -187
rect -1656 -255 -1622 -235
rect -1656 -269 -1622 -255
rect -1358 255 -1324 269
rect -1358 235 -1324 255
rect -1358 187 -1324 197
rect -1358 163 -1324 187
rect -1358 119 -1324 125
rect -1358 91 -1324 119
rect -1358 51 -1324 53
rect -1358 19 -1324 51
rect -1358 -51 -1324 -19
rect -1358 -53 -1324 -51
rect -1358 -119 -1324 -91
rect -1358 -125 -1324 -119
rect -1358 -187 -1324 -163
rect -1358 -197 -1324 -187
rect -1358 -255 -1324 -235
rect -1358 -269 -1324 -255
rect -1060 255 -1026 269
rect -1060 235 -1026 255
rect -1060 187 -1026 197
rect -1060 163 -1026 187
rect -1060 119 -1026 125
rect -1060 91 -1026 119
rect -1060 51 -1026 53
rect -1060 19 -1026 51
rect -1060 -51 -1026 -19
rect -1060 -53 -1026 -51
rect -1060 -119 -1026 -91
rect -1060 -125 -1026 -119
rect -1060 -187 -1026 -163
rect -1060 -197 -1026 -187
rect -1060 -255 -1026 -235
rect -1060 -269 -1026 -255
rect -762 255 -728 269
rect -762 235 -728 255
rect -762 187 -728 197
rect -762 163 -728 187
rect -762 119 -728 125
rect -762 91 -728 119
rect -762 51 -728 53
rect -762 19 -728 51
rect -762 -51 -728 -19
rect -762 -53 -728 -51
rect -762 -119 -728 -91
rect -762 -125 -728 -119
rect -762 -187 -728 -163
rect -762 -197 -728 -187
rect -762 -255 -728 -235
rect -762 -269 -728 -255
rect -464 255 -430 269
rect -464 235 -430 255
rect -464 187 -430 197
rect -464 163 -430 187
rect -464 119 -430 125
rect -464 91 -430 119
rect -464 51 -430 53
rect -464 19 -430 51
rect -464 -51 -430 -19
rect -464 -53 -430 -51
rect -464 -119 -430 -91
rect -464 -125 -430 -119
rect -464 -187 -430 -163
rect -464 -197 -430 -187
rect -464 -255 -430 -235
rect -464 -269 -430 -255
rect -166 255 -132 269
rect -166 235 -132 255
rect -166 187 -132 197
rect -166 163 -132 187
rect -166 119 -132 125
rect -166 91 -132 119
rect -166 51 -132 53
rect -166 19 -132 51
rect -166 -51 -132 -19
rect -166 -53 -132 -51
rect -166 -119 -132 -91
rect -166 -125 -132 -119
rect -166 -187 -132 -163
rect -166 -197 -132 -187
rect -166 -255 -132 -235
rect -166 -269 -132 -255
rect 132 255 166 269
rect 132 235 166 255
rect 132 187 166 197
rect 132 163 166 187
rect 132 119 166 125
rect 132 91 166 119
rect 132 51 166 53
rect 132 19 166 51
rect 132 -51 166 -19
rect 132 -53 166 -51
rect 132 -119 166 -91
rect 132 -125 166 -119
rect 132 -187 166 -163
rect 132 -197 166 -187
rect 132 -255 166 -235
rect 132 -269 166 -255
rect 430 255 464 269
rect 430 235 464 255
rect 430 187 464 197
rect 430 163 464 187
rect 430 119 464 125
rect 430 91 464 119
rect 430 51 464 53
rect 430 19 464 51
rect 430 -51 464 -19
rect 430 -53 464 -51
rect 430 -119 464 -91
rect 430 -125 464 -119
rect 430 -187 464 -163
rect 430 -197 464 -187
rect 430 -255 464 -235
rect 430 -269 464 -255
rect 728 255 762 269
rect 728 235 762 255
rect 728 187 762 197
rect 728 163 762 187
rect 728 119 762 125
rect 728 91 762 119
rect 728 51 762 53
rect 728 19 762 51
rect 728 -51 762 -19
rect 728 -53 762 -51
rect 728 -119 762 -91
rect 728 -125 762 -119
rect 728 -187 762 -163
rect 728 -197 762 -187
rect 728 -255 762 -235
rect 728 -269 762 -255
rect 1026 255 1060 269
rect 1026 235 1060 255
rect 1026 187 1060 197
rect 1026 163 1060 187
rect 1026 119 1060 125
rect 1026 91 1060 119
rect 1026 51 1060 53
rect 1026 19 1060 51
rect 1026 -51 1060 -19
rect 1026 -53 1060 -51
rect 1026 -119 1060 -91
rect 1026 -125 1060 -119
rect 1026 -187 1060 -163
rect 1026 -197 1060 -187
rect 1026 -255 1060 -235
rect 1026 -269 1060 -255
rect 1324 255 1358 269
rect 1324 235 1358 255
rect 1324 187 1358 197
rect 1324 163 1358 187
rect 1324 119 1358 125
rect 1324 91 1358 119
rect 1324 51 1358 53
rect 1324 19 1358 51
rect 1324 -51 1358 -19
rect 1324 -53 1358 -51
rect 1324 -119 1358 -91
rect 1324 -125 1358 -119
rect 1324 -187 1358 -163
rect 1324 -197 1358 -187
rect 1324 -255 1358 -235
rect 1324 -269 1358 -255
rect 1622 255 1656 269
rect 1622 235 1656 255
rect 1622 187 1656 197
rect 1622 163 1656 187
rect 1622 119 1656 125
rect 1622 91 1656 119
rect 1622 51 1656 53
rect 1622 19 1656 51
rect 1622 -51 1656 -19
rect 1622 -53 1656 -51
rect 1622 -119 1656 -91
rect 1622 -125 1656 -119
rect 1622 -187 1656 -163
rect 1622 -197 1656 -187
rect 1622 -255 1656 -235
rect 1622 -269 1656 -255
rect -1507 -372 -1473 -338
rect -1209 -372 -1175 -338
rect -911 -372 -877 -338
rect -613 -372 -579 -338
rect -315 -372 -281 -338
rect -17 -372 17 -338
rect 281 -372 315 -338
rect 579 -372 613 -338
rect 877 -372 911 -338
rect 1175 -372 1209 -338
rect 1473 -372 1507 -338
<< metal1 >>
rect -1554 372 -1426 378
rect -1554 338 -1507 372
rect -1473 338 -1426 372
rect -1554 332 -1426 338
rect -1256 372 -1128 378
rect -1256 338 -1209 372
rect -1175 338 -1128 372
rect -1256 332 -1128 338
rect -958 372 -830 378
rect -958 338 -911 372
rect -877 338 -830 372
rect -958 332 -830 338
rect -660 372 -532 378
rect -660 338 -613 372
rect -579 338 -532 372
rect -660 332 -532 338
rect -362 372 -234 378
rect -362 338 -315 372
rect -281 338 -234 372
rect -362 332 -234 338
rect -64 372 64 378
rect -64 338 -17 372
rect 17 338 64 372
rect -64 332 64 338
rect 234 372 362 378
rect 234 338 281 372
rect 315 338 362 372
rect 234 332 362 338
rect 532 372 660 378
rect 532 338 579 372
rect 613 338 660 372
rect 532 332 660 338
rect 830 372 958 378
rect 830 338 877 372
rect 911 338 958 372
rect 830 332 958 338
rect 1128 372 1256 378
rect 1128 338 1175 372
rect 1209 338 1256 372
rect 1128 332 1256 338
rect 1426 372 1554 378
rect 1426 338 1473 372
rect 1507 338 1554 372
rect 1426 332 1554 338
rect -1662 269 -1616 300
rect -1662 235 -1656 269
rect -1622 235 -1616 269
rect -1662 197 -1616 235
rect -1662 163 -1656 197
rect -1622 163 -1616 197
rect -1662 125 -1616 163
rect -1662 91 -1656 125
rect -1622 91 -1616 125
rect -1662 53 -1616 91
rect -1662 19 -1656 53
rect -1622 19 -1616 53
rect -1662 -19 -1616 19
rect -1662 -53 -1656 -19
rect -1622 -53 -1616 -19
rect -1662 -91 -1616 -53
rect -1662 -125 -1656 -91
rect -1622 -125 -1616 -91
rect -1662 -163 -1616 -125
rect -1662 -197 -1656 -163
rect -1622 -197 -1616 -163
rect -1662 -235 -1616 -197
rect -1662 -269 -1656 -235
rect -1622 -269 -1616 -235
rect -1662 -300 -1616 -269
rect -1364 269 -1318 300
rect -1364 235 -1358 269
rect -1324 235 -1318 269
rect -1364 197 -1318 235
rect -1364 163 -1358 197
rect -1324 163 -1318 197
rect -1364 125 -1318 163
rect -1364 91 -1358 125
rect -1324 91 -1318 125
rect -1364 53 -1318 91
rect -1364 19 -1358 53
rect -1324 19 -1318 53
rect -1364 -19 -1318 19
rect -1364 -53 -1358 -19
rect -1324 -53 -1318 -19
rect -1364 -91 -1318 -53
rect -1364 -125 -1358 -91
rect -1324 -125 -1318 -91
rect -1364 -163 -1318 -125
rect -1364 -197 -1358 -163
rect -1324 -197 -1318 -163
rect -1364 -235 -1318 -197
rect -1364 -269 -1358 -235
rect -1324 -269 -1318 -235
rect -1364 -300 -1318 -269
rect -1066 269 -1020 300
rect -1066 235 -1060 269
rect -1026 235 -1020 269
rect -1066 197 -1020 235
rect -1066 163 -1060 197
rect -1026 163 -1020 197
rect -1066 125 -1020 163
rect -1066 91 -1060 125
rect -1026 91 -1020 125
rect -1066 53 -1020 91
rect -1066 19 -1060 53
rect -1026 19 -1020 53
rect -1066 -19 -1020 19
rect -1066 -53 -1060 -19
rect -1026 -53 -1020 -19
rect -1066 -91 -1020 -53
rect -1066 -125 -1060 -91
rect -1026 -125 -1020 -91
rect -1066 -163 -1020 -125
rect -1066 -197 -1060 -163
rect -1026 -197 -1020 -163
rect -1066 -235 -1020 -197
rect -1066 -269 -1060 -235
rect -1026 -269 -1020 -235
rect -1066 -300 -1020 -269
rect -768 269 -722 300
rect -768 235 -762 269
rect -728 235 -722 269
rect -768 197 -722 235
rect -768 163 -762 197
rect -728 163 -722 197
rect -768 125 -722 163
rect -768 91 -762 125
rect -728 91 -722 125
rect -768 53 -722 91
rect -768 19 -762 53
rect -728 19 -722 53
rect -768 -19 -722 19
rect -768 -53 -762 -19
rect -728 -53 -722 -19
rect -768 -91 -722 -53
rect -768 -125 -762 -91
rect -728 -125 -722 -91
rect -768 -163 -722 -125
rect -768 -197 -762 -163
rect -728 -197 -722 -163
rect -768 -235 -722 -197
rect -768 -269 -762 -235
rect -728 -269 -722 -235
rect -768 -300 -722 -269
rect -470 269 -424 300
rect -470 235 -464 269
rect -430 235 -424 269
rect -470 197 -424 235
rect -470 163 -464 197
rect -430 163 -424 197
rect -470 125 -424 163
rect -470 91 -464 125
rect -430 91 -424 125
rect -470 53 -424 91
rect -470 19 -464 53
rect -430 19 -424 53
rect -470 -19 -424 19
rect -470 -53 -464 -19
rect -430 -53 -424 -19
rect -470 -91 -424 -53
rect -470 -125 -464 -91
rect -430 -125 -424 -91
rect -470 -163 -424 -125
rect -470 -197 -464 -163
rect -430 -197 -424 -163
rect -470 -235 -424 -197
rect -470 -269 -464 -235
rect -430 -269 -424 -235
rect -470 -300 -424 -269
rect -172 269 -126 300
rect -172 235 -166 269
rect -132 235 -126 269
rect -172 197 -126 235
rect -172 163 -166 197
rect -132 163 -126 197
rect -172 125 -126 163
rect -172 91 -166 125
rect -132 91 -126 125
rect -172 53 -126 91
rect -172 19 -166 53
rect -132 19 -126 53
rect -172 -19 -126 19
rect -172 -53 -166 -19
rect -132 -53 -126 -19
rect -172 -91 -126 -53
rect -172 -125 -166 -91
rect -132 -125 -126 -91
rect -172 -163 -126 -125
rect -172 -197 -166 -163
rect -132 -197 -126 -163
rect -172 -235 -126 -197
rect -172 -269 -166 -235
rect -132 -269 -126 -235
rect -172 -300 -126 -269
rect 126 269 172 300
rect 126 235 132 269
rect 166 235 172 269
rect 126 197 172 235
rect 126 163 132 197
rect 166 163 172 197
rect 126 125 172 163
rect 126 91 132 125
rect 166 91 172 125
rect 126 53 172 91
rect 126 19 132 53
rect 166 19 172 53
rect 126 -19 172 19
rect 126 -53 132 -19
rect 166 -53 172 -19
rect 126 -91 172 -53
rect 126 -125 132 -91
rect 166 -125 172 -91
rect 126 -163 172 -125
rect 126 -197 132 -163
rect 166 -197 172 -163
rect 126 -235 172 -197
rect 126 -269 132 -235
rect 166 -269 172 -235
rect 126 -300 172 -269
rect 424 269 470 300
rect 424 235 430 269
rect 464 235 470 269
rect 424 197 470 235
rect 424 163 430 197
rect 464 163 470 197
rect 424 125 470 163
rect 424 91 430 125
rect 464 91 470 125
rect 424 53 470 91
rect 424 19 430 53
rect 464 19 470 53
rect 424 -19 470 19
rect 424 -53 430 -19
rect 464 -53 470 -19
rect 424 -91 470 -53
rect 424 -125 430 -91
rect 464 -125 470 -91
rect 424 -163 470 -125
rect 424 -197 430 -163
rect 464 -197 470 -163
rect 424 -235 470 -197
rect 424 -269 430 -235
rect 464 -269 470 -235
rect 424 -300 470 -269
rect 722 269 768 300
rect 722 235 728 269
rect 762 235 768 269
rect 722 197 768 235
rect 722 163 728 197
rect 762 163 768 197
rect 722 125 768 163
rect 722 91 728 125
rect 762 91 768 125
rect 722 53 768 91
rect 722 19 728 53
rect 762 19 768 53
rect 722 -19 768 19
rect 722 -53 728 -19
rect 762 -53 768 -19
rect 722 -91 768 -53
rect 722 -125 728 -91
rect 762 -125 768 -91
rect 722 -163 768 -125
rect 722 -197 728 -163
rect 762 -197 768 -163
rect 722 -235 768 -197
rect 722 -269 728 -235
rect 762 -269 768 -235
rect 722 -300 768 -269
rect 1020 269 1066 300
rect 1020 235 1026 269
rect 1060 235 1066 269
rect 1020 197 1066 235
rect 1020 163 1026 197
rect 1060 163 1066 197
rect 1020 125 1066 163
rect 1020 91 1026 125
rect 1060 91 1066 125
rect 1020 53 1066 91
rect 1020 19 1026 53
rect 1060 19 1066 53
rect 1020 -19 1066 19
rect 1020 -53 1026 -19
rect 1060 -53 1066 -19
rect 1020 -91 1066 -53
rect 1020 -125 1026 -91
rect 1060 -125 1066 -91
rect 1020 -163 1066 -125
rect 1020 -197 1026 -163
rect 1060 -197 1066 -163
rect 1020 -235 1066 -197
rect 1020 -269 1026 -235
rect 1060 -269 1066 -235
rect 1020 -300 1066 -269
rect 1318 269 1364 300
rect 1318 235 1324 269
rect 1358 235 1364 269
rect 1318 197 1364 235
rect 1318 163 1324 197
rect 1358 163 1364 197
rect 1318 125 1364 163
rect 1318 91 1324 125
rect 1358 91 1364 125
rect 1318 53 1364 91
rect 1318 19 1324 53
rect 1358 19 1364 53
rect 1318 -19 1364 19
rect 1318 -53 1324 -19
rect 1358 -53 1364 -19
rect 1318 -91 1364 -53
rect 1318 -125 1324 -91
rect 1358 -125 1364 -91
rect 1318 -163 1364 -125
rect 1318 -197 1324 -163
rect 1358 -197 1364 -163
rect 1318 -235 1364 -197
rect 1318 -269 1324 -235
rect 1358 -269 1364 -235
rect 1318 -300 1364 -269
rect 1616 269 1662 300
rect 1616 235 1622 269
rect 1656 235 1662 269
rect 1616 197 1662 235
rect 1616 163 1622 197
rect 1656 163 1662 197
rect 1616 125 1662 163
rect 1616 91 1622 125
rect 1656 91 1662 125
rect 1616 53 1662 91
rect 1616 19 1622 53
rect 1656 19 1662 53
rect 1616 -19 1662 19
rect 1616 -53 1622 -19
rect 1656 -53 1662 -19
rect 1616 -91 1662 -53
rect 1616 -125 1622 -91
rect 1656 -125 1662 -91
rect 1616 -163 1662 -125
rect 1616 -197 1622 -163
rect 1656 -197 1662 -163
rect 1616 -235 1662 -197
rect 1616 -269 1622 -235
rect 1656 -269 1662 -235
rect 1616 -300 1662 -269
rect -1554 -338 -1426 -332
rect -1554 -372 -1507 -338
rect -1473 -372 -1426 -338
rect -1554 -378 -1426 -372
rect -1256 -338 -1128 -332
rect -1256 -372 -1209 -338
rect -1175 -372 -1128 -338
rect -1256 -378 -1128 -372
rect -958 -338 -830 -332
rect -958 -372 -911 -338
rect -877 -372 -830 -338
rect -958 -378 -830 -372
rect -660 -338 -532 -332
rect -660 -372 -613 -338
rect -579 -372 -532 -338
rect -660 -378 -532 -372
rect -362 -338 -234 -332
rect -362 -372 -315 -338
rect -281 -372 -234 -338
rect -362 -378 -234 -372
rect -64 -338 64 -332
rect -64 -372 -17 -338
rect 17 -372 64 -338
rect -64 -378 64 -372
rect 234 -338 362 -332
rect 234 -372 281 -338
rect 315 -372 362 -338
rect 234 -378 362 -372
rect 532 -338 660 -332
rect 532 -372 579 -338
rect 613 -372 660 -338
rect 532 -378 660 -372
rect 830 -338 958 -332
rect 830 -372 877 -338
rect 911 -372 958 -338
rect 830 -378 958 -372
rect 1128 -338 1256 -332
rect 1128 -372 1175 -338
rect 1209 -372 1256 -338
rect 1128 -378 1256 -372
rect 1426 -338 1554 -332
rect 1426 -372 1473 -338
rect 1507 -372 1554 -338
rect 1426 -378 1554 -372
<< end >>
