magic
tech sky130A
magscale 1 2
timestamp 1620626447
<< nwell >>
rect -1257 -1373 1257 1373
<< pmos >>
rect -1061 754 -901 1154
rect -843 754 -683 1154
rect -625 754 -465 1154
rect -407 754 -247 1154
rect -189 754 -29 1154
rect 29 754 189 1154
rect 247 754 407 1154
rect 465 754 625 1154
rect 683 754 843 1154
rect 901 754 1061 1154
rect -1061 118 -901 518
rect -843 118 -683 518
rect -625 118 -465 518
rect -407 118 -247 518
rect -189 118 -29 518
rect 29 118 189 518
rect 247 118 407 518
rect 465 118 625 518
rect 683 118 843 518
rect 901 118 1061 518
rect -1061 -518 -901 -118
rect -843 -518 -683 -118
rect -625 -518 -465 -118
rect -407 -518 -247 -118
rect -189 -518 -29 -118
rect 29 -518 189 -118
rect 247 -518 407 -118
rect 465 -518 625 -118
rect 683 -518 843 -118
rect 901 -518 1061 -118
rect -1061 -1154 -901 -754
rect -843 -1154 -683 -754
rect -625 -1154 -465 -754
rect -407 -1154 -247 -754
rect -189 -1154 -29 -754
rect 29 -1154 189 -754
rect 247 -1154 407 -754
rect 465 -1154 625 -754
rect 683 -1154 843 -754
rect 901 -1154 1061 -754
<< pdiff >>
rect -1119 1142 -1061 1154
rect -1119 766 -1107 1142
rect -1073 766 -1061 1142
rect -1119 754 -1061 766
rect -901 1142 -843 1154
rect -901 766 -889 1142
rect -855 766 -843 1142
rect -901 754 -843 766
rect -683 1142 -625 1154
rect -683 766 -671 1142
rect -637 766 -625 1142
rect -683 754 -625 766
rect -465 1142 -407 1154
rect -465 766 -453 1142
rect -419 766 -407 1142
rect -465 754 -407 766
rect -247 1142 -189 1154
rect -247 766 -235 1142
rect -201 766 -189 1142
rect -247 754 -189 766
rect -29 1142 29 1154
rect -29 766 -17 1142
rect 17 766 29 1142
rect -29 754 29 766
rect 189 1142 247 1154
rect 189 766 201 1142
rect 235 766 247 1142
rect 189 754 247 766
rect 407 1142 465 1154
rect 407 766 419 1142
rect 453 766 465 1142
rect 407 754 465 766
rect 625 1142 683 1154
rect 625 766 637 1142
rect 671 766 683 1142
rect 625 754 683 766
rect 843 1142 901 1154
rect 843 766 855 1142
rect 889 766 901 1142
rect 843 754 901 766
rect 1061 1142 1119 1154
rect 1061 766 1073 1142
rect 1107 766 1119 1142
rect 1061 754 1119 766
rect -1119 506 -1061 518
rect -1119 130 -1107 506
rect -1073 130 -1061 506
rect -1119 118 -1061 130
rect -901 506 -843 518
rect -901 130 -889 506
rect -855 130 -843 506
rect -901 118 -843 130
rect -683 506 -625 518
rect -683 130 -671 506
rect -637 130 -625 506
rect -683 118 -625 130
rect -465 506 -407 518
rect -465 130 -453 506
rect -419 130 -407 506
rect -465 118 -407 130
rect -247 506 -189 518
rect -247 130 -235 506
rect -201 130 -189 506
rect -247 118 -189 130
rect -29 506 29 518
rect -29 130 -17 506
rect 17 130 29 506
rect -29 118 29 130
rect 189 506 247 518
rect 189 130 201 506
rect 235 130 247 506
rect 189 118 247 130
rect 407 506 465 518
rect 407 130 419 506
rect 453 130 465 506
rect 407 118 465 130
rect 625 506 683 518
rect 625 130 637 506
rect 671 130 683 506
rect 625 118 683 130
rect 843 506 901 518
rect 843 130 855 506
rect 889 130 901 506
rect 843 118 901 130
rect 1061 506 1119 518
rect 1061 130 1073 506
rect 1107 130 1119 506
rect 1061 118 1119 130
rect -1119 -130 -1061 -118
rect -1119 -506 -1107 -130
rect -1073 -506 -1061 -130
rect -1119 -518 -1061 -506
rect -901 -130 -843 -118
rect -901 -506 -889 -130
rect -855 -506 -843 -130
rect -901 -518 -843 -506
rect -683 -130 -625 -118
rect -683 -506 -671 -130
rect -637 -506 -625 -130
rect -683 -518 -625 -506
rect -465 -130 -407 -118
rect -465 -506 -453 -130
rect -419 -506 -407 -130
rect -465 -518 -407 -506
rect -247 -130 -189 -118
rect -247 -506 -235 -130
rect -201 -506 -189 -130
rect -247 -518 -189 -506
rect -29 -130 29 -118
rect -29 -506 -17 -130
rect 17 -506 29 -130
rect -29 -518 29 -506
rect 189 -130 247 -118
rect 189 -506 201 -130
rect 235 -506 247 -130
rect 189 -518 247 -506
rect 407 -130 465 -118
rect 407 -506 419 -130
rect 453 -506 465 -130
rect 407 -518 465 -506
rect 625 -130 683 -118
rect 625 -506 637 -130
rect 671 -506 683 -130
rect 625 -518 683 -506
rect 843 -130 901 -118
rect 843 -506 855 -130
rect 889 -506 901 -130
rect 843 -518 901 -506
rect 1061 -130 1119 -118
rect 1061 -506 1073 -130
rect 1107 -506 1119 -130
rect 1061 -518 1119 -506
rect -1119 -766 -1061 -754
rect -1119 -1142 -1107 -766
rect -1073 -1142 -1061 -766
rect -1119 -1154 -1061 -1142
rect -901 -766 -843 -754
rect -901 -1142 -889 -766
rect -855 -1142 -843 -766
rect -901 -1154 -843 -1142
rect -683 -766 -625 -754
rect -683 -1142 -671 -766
rect -637 -1142 -625 -766
rect -683 -1154 -625 -1142
rect -465 -766 -407 -754
rect -465 -1142 -453 -766
rect -419 -1142 -407 -766
rect -465 -1154 -407 -1142
rect -247 -766 -189 -754
rect -247 -1142 -235 -766
rect -201 -1142 -189 -766
rect -247 -1154 -189 -1142
rect -29 -766 29 -754
rect -29 -1142 -17 -766
rect 17 -1142 29 -766
rect -29 -1154 29 -1142
rect 189 -766 247 -754
rect 189 -1142 201 -766
rect 235 -1142 247 -766
rect 189 -1154 247 -1142
rect 407 -766 465 -754
rect 407 -1142 419 -766
rect 453 -1142 465 -766
rect 407 -1154 465 -1142
rect 625 -766 683 -754
rect 625 -1142 637 -766
rect 671 -1142 683 -766
rect 625 -1154 683 -1142
rect 843 -766 901 -754
rect 843 -1142 855 -766
rect 889 -1142 901 -766
rect 843 -1154 901 -1142
rect 1061 -766 1119 -754
rect 1061 -1142 1073 -766
rect 1107 -1142 1119 -766
rect 1061 -1154 1119 -1142
<< pdiffc >>
rect -1107 766 -1073 1142
rect -889 766 -855 1142
rect -671 766 -637 1142
rect -453 766 -419 1142
rect -235 766 -201 1142
rect -17 766 17 1142
rect 201 766 235 1142
rect 419 766 453 1142
rect 637 766 671 1142
rect 855 766 889 1142
rect 1073 766 1107 1142
rect -1107 130 -1073 506
rect -889 130 -855 506
rect -671 130 -637 506
rect -453 130 -419 506
rect -235 130 -201 506
rect -17 130 17 506
rect 201 130 235 506
rect 419 130 453 506
rect 637 130 671 506
rect 855 130 889 506
rect 1073 130 1107 506
rect -1107 -506 -1073 -130
rect -889 -506 -855 -130
rect -671 -506 -637 -130
rect -453 -506 -419 -130
rect -235 -506 -201 -130
rect -17 -506 17 -130
rect 201 -506 235 -130
rect 419 -506 453 -130
rect 637 -506 671 -130
rect 855 -506 889 -130
rect 1073 -506 1107 -130
rect -1107 -1142 -1073 -766
rect -889 -1142 -855 -766
rect -671 -1142 -637 -766
rect -453 -1142 -419 -766
rect -235 -1142 -201 -766
rect -17 -1142 17 -766
rect 201 -1142 235 -766
rect 419 -1142 453 -766
rect 637 -1142 671 -766
rect 855 -1142 889 -766
rect 1073 -1142 1107 -766
<< nsubdiff >>
rect -1221 1303 -1125 1337
rect 1125 1303 1221 1337
rect -1221 1241 -1187 1303
rect 1187 1241 1221 1303
rect -1221 -1303 -1187 -1241
rect 1187 -1303 1221 -1241
rect -1221 -1337 -1125 -1303
rect 1125 -1337 1221 -1303
<< nsubdiffcont >>
rect -1125 1303 1125 1337
rect -1221 -1241 -1187 1241
rect 1187 -1241 1221 1241
rect -1125 -1337 1125 -1303
<< poly >>
rect -1035 1235 -927 1251
rect -1035 1218 -1019 1235
rect -1061 1201 -1019 1218
rect -943 1218 -927 1235
rect -817 1235 -709 1251
rect -817 1218 -801 1235
rect -943 1201 -901 1218
rect -1061 1154 -901 1201
rect -843 1201 -801 1218
rect -725 1218 -709 1235
rect -599 1235 -491 1251
rect -599 1218 -583 1235
rect -725 1201 -683 1218
rect -843 1154 -683 1201
rect -625 1201 -583 1218
rect -507 1218 -491 1235
rect -381 1235 -273 1251
rect -381 1218 -365 1235
rect -507 1201 -465 1218
rect -625 1154 -465 1201
rect -407 1201 -365 1218
rect -289 1218 -273 1235
rect -163 1235 -55 1251
rect -163 1218 -147 1235
rect -289 1201 -247 1218
rect -407 1154 -247 1201
rect -189 1201 -147 1218
rect -71 1218 -55 1235
rect 55 1235 163 1251
rect 55 1218 71 1235
rect -71 1201 -29 1218
rect -189 1154 -29 1201
rect 29 1201 71 1218
rect 147 1218 163 1235
rect 273 1235 381 1251
rect 273 1218 289 1235
rect 147 1201 189 1218
rect 29 1154 189 1201
rect 247 1201 289 1218
rect 365 1218 381 1235
rect 491 1235 599 1251
rect 491 1218 507 1235
rect 365 1201 407 1218
rect 247 1154 407 1201
rect 465 1201 507 1218
rect 583 1218 599 1235
rect 709 1235 817 1251
rect 709 1218 725 1235
rect 583 1201 625 1218
rect 465 1154 625 1201
rect 683 1201 725 1218
rect 801 1218 817 1235
rect 927 1235 1035 1251
rect 927 1218 943 1235
rect 801 1201 843 1218
rect 683 1154 843 1201
rect 901 1201 943 1218
rect 1019 1218 1035 1235
rect 1019 1201 1061 1218
rect 901 1154 1061 1201
rect -1061 707 -901 754
rect -1061 690 -1019 707
rect -1035 673 -1019 690
rect -943 690 -901 707
rect -843 707 -683 754
rect -843 690 -801 707
rect -943 673 -927 690
rect -1035 657 -927 673
rect -817 673 -801 690
rect -725 690 -683 707
rect -625 707 -465 754
rect -625 690 -583 707
rect -725 673 -709 690
rect -817 657 -709 673
rect -599 673 -583 690
rect -507 690 -465 707
rect -407 707 -247 754
rect -407 690 -365 707
rect -507 673 -491 690
rect -599 657 -491 673
rect -381 673 -365 690
rect -289 690 -247 707
rect -189 707 -29 754
rect -189 690 -147 707
rect -289 673 -273 690
rect -381 657 -273 673
rect -163 673 -147 690
rect -71 690 -29 707
rect 29 707 189 754
rect 29 690 71 707
rect -71 673 -55 690
rect -163 657 -55 673
rect 55 673 71 690
rect 147 690 189 707
rect 247 707 407 754
rect 247 690 289 707
rect 147 673 163 690
rect 55 657 163 673
rect 273 673 289 690
rect 365 690 407 707
rect 465 707 625 754
rect 465 690 507 707
rect 365 673 381 690
rect 273 657 381 673
rect 491 673 507 690
rect 583 690 625 707
rect 683 707 843 754
rect 683 690 725 707
rect 583 673 599 690
rect 491 657 599 673
rect 709 673 725 690
rect 801 690 843 707
rect 901 707 1061 754
rect 901 690 943 707
rect 801 673 817 690
rect 709 657 817 673
rect 927 673 943 690
rect 1019 690 1061 707
rect 1019 673 1035 690
rect 927 657 1035 673
rect -1035 599 -927 615
rect -1035 582 -1019 599
rect -1061 565 -1019 582
rect -943 582 -927 599
rect -817 599 -709 615
rect -817 582 -801 599
rect -943 565 -901 582
rect -1061 518 -901 565
rect -843 565 -801 582
rect -725 582 -709 599
rect -599 599 -491 615
rect -599 582 -583 599
rect -725 565 -683 582
rect -843 518 -683 565
rect -625 565 -583 582
rect -507 582 -491 599
rect -381 599 -273 615
rect -381 582 -365 599
rect -507 565 -465 582
rect -625 518 -465 565
rect -407 565 -365 582
rect -289 582 -273 599
rect -163 599 -55 615
rect -163 582 -147 599
rect -289 565 -247 582
rect -407 518 -247 565
rect -189 565 -147 582
rect -71 582 -55 599
rect 55 599 163 615
rect 55 582 71 599
rect -71 565 -29 582
rect -189 518 -29 565
rect 29 565 71 582
rect 147 582 163 599
rect 273 599 381 615
rect 273 582 289 599
rect 147 565 189 582
rect 29 518 189 565
rect 247 565 289 582
rect 365 582 381 599
rect 491 599 599 615
rect 491 582 507 599
rect 365 565 407 582
rect 247 518 407 565
rect 465 565 507 582
rect 583 582 599 599
rect 709 599 817 615
rect 709 582 725 599
rect 583 565 625 582
rect 465 518 625 565
rect 683 565 725 582
rect 801 582 817 599
rect 927 599 1035 615
rect 927 582 943 599
rect 801 565 843 582
rect 683 518 843 565
rect 901 565 943 582
rect 1019 582 1035 599
rect 1019 565 1061 582
rect 901 518 1061 565
rect -1061 71 -901 118
rect -1061 54 -1019 71
rect -1035 37 -1019 54
rect -943 54 -901 71
rect -843 71 -683 118
rect -843 54 -801 71
rect -943 37 -927 54
rect -1035 21 -927 37
rect -817 37 -801 54
rect -725 54 -683 71
rect -625 71 -465 118
rect -625 54 -583 71
rect -725 37 -709 54
rect -817 21 -709 37
rect -599 37 -583 54
rect -507 54 -465 71
rect -407 71 -247 118
rect -407 54 -365 71
rect -507 37 -491 54
rect -599 21 -491 37
rect -381 37 -365 54
rect -289 54 -247 71
rect -189 71 -29 118
rect -189 54 -147 71
rect -289 37 -273 54
rect -381 21 -273 37
rect -163 37 -147 54
rect -71 54 -29 71
rect 29 71 189 118
rect 29 54 71 71
rect -71 37 -55 54
rect -163 21 -55 37
rect 55 37 71 54
rect 147 54 189 71
rect 247 71 407 118
rect 247 54 289 71
rect 147 37 163 54
rect 55 21 163 37
rect 273 37 289 54
rect 365 54 407 71
rect 465 71 625 118
rect 465 54 507 71
rect 365 37 381 54
rect 273 21 381 37
rect 491 37 507 54
rect 583 54 625 71
rect 683 71 843 118
rect 683 54 725 71
rect 583 37 599 54
rect 491 21 599 37
rect 709 37 725 54
rect 801 54 843 71
rect 901 71 1061 118
rect 901 54 943 71
rect 801 37 817 54
rect 709 21 817 37
rect 927 37 943 54
rect 1019 54 1061 71
rect 1019 37 1035 54
rect 927 21 1035 37
rect -1035 -37 -927 -21
rect -1035 -54 -1019 -37
rect -1061 -71 -1019 -54
rect -943 -54 -927 -37
rect -817 -37 -709 -21
rect -817 -54 -801 -37
rect -943 -71 -901 -54
rect -1061 -118 -901 -71
rect -843 -71 -801 -54
rect -725 -54 -709 -37
rect -599 -37 -491 -21
rect -599 -54 -583 -37
rect -725 -71 -683 -54
rect -843 -118 -683 -71
rect -625 -71 -583 -54
rect -507 -54 -491 -37
rect -381 -37 -273 -21
rect -381 -54 -365 -37
rect -507 -71 -465 -54
rect -625 -118 -465 -71
rect -407 -71 -365 -54
rect -289 -54 -273 -37
rect -163 -37 -55 -21
rect -163 -54 -147 -37
rect -289 -71 -247 -54
rect -407 -118 -247 -71
rect -189 -71 -147 -54
rect -71 -54 -55 -37
rect 55 -37 163 -21
rect 55 -54 71 -37
rect -71 -71 -29 -54
rect -189 -118 -29 -71
rect 29 -71 71 -54
rect 147 -54 163 -37
rect 273 -37 381 -21
rect 273 -54 289 -37
rect 147 -71 189 -54
rect 29 -118 189 -71
rect 247 -71 289 -54
rect 365 -54 381 -37
rect 491 -37 599 -21
rect 491 -54 507 -37
rect 365 -71 407 -54
rect 247 -118 407 -71
rect 465 -71 507 -54
rect 583 -54 599 -37
rect 709 -37 817 -21
rect 709 -54 725 -37
rect 583 -71 625 -54
rect 465 -118 625 -71
rect 683 -71 725 -54
rect 801 -54 817 -37
rect 927 -37 1035 -21
rect 927 -54 943 -37
rect 801 -71 843 -54
rect 683 -118 843 -71
rect 901 -71 943 -54
rect 1019 -54 1035 -37
rect 1019 -71 1061 -54
rect 901 -118 1061 -71
rect -1061 -565 -901 -518
rect -1061 -582 -1019 -565
rect -1035 -599 -1019 -582
rect -943 -582 -901 -565
rect -843 -565 -683 -518
rect -843 -582 -801 -565
rect -943 -599 -927 -582
rect -1035 -615 -927 -599
rect -817 -599 -801 -582
rect -725 -582 -683 -565
rect -625 -565 -465 -518
rect -625 -582 -583 -565
rect -725 -599 -709 -582
rect -817 -615 -709 -599
rect -599 -599 -583 -582
rect -507 -582 -465 -565
rect -407 -565 -247 -518
rect -407 -582 -365 -565
rect -507 -599 -491 -582
rect -599 -615 -491 -599
rect -381 -599 -365 -582
rect -289 -582 -247 -565
rect -189 -565 -29 -518
rect -189 -582 -147 -565
rect -289 -599 -273 -582
rect -381 -615 -273 -599
rect -163 -599 -147 -582
rect -71 -582 -29 -565
rect 29 -565 189 -518
rect 29 -582 71 -565
rect -71 -599 -55 -582
rect -163 -615 -55 -599
rect 55 -599 71 -582
rect 147 -582 189 -565
rect 247 -565 407 -518
rect 247 -582 289 -565
rect 147 -599 163 -582
rect 55 -615 163 -599
rect 273 -599 289 -582
rect 365 -582 407 -565
rect 465 -565 625 -518
rect 465 -582 507 -565
rect 365 -599 381 -582
rect 273 -615 381 -599
rect 491 -599 507 -582
rect 583 -582 625 -565
rect 683 -565 843 -518
rect 683 -582 725 -565
rect 583 -599 599 -582
rect 491 -615 599 -599
rect 709 -599 725 -582
rect 801 -582 843 -565
rect 901 -565 1061 -518
rect 901 -582 943 -565
rect 801 -599 817 -582
rect 709 -615 817 -599
rect 927 -599 943 -582
rect 1019 -582 1061 -565
rect 1019 -599 1035 -582
rect 927 -615 1035 -599
rect -1035 -673 -927 -657
rect -1035 -690 -1019 -673
rect -1061 -707 -1019 -690
rect -943 -690 -927 -673
rect -817 -673 -709 -657
rect -817 -690 -801 -673
rect -943 -707 -901 -690
rect -1061 -754 -901 -707
rect -843 -707 -801 -690
rect -725 -690 -709 -673
rect -599 -673 -491 -657
rect -599 -690 -583 -673
rect -725 -707 -683 -690
rect -843 -754 -683 -707
rect -625 -707 -583 -690
rect -507 -690 -491 -673
rect -381 -673 -273 -657
rect -381 -690 -365 -673
rect -507 -707 -465 -690
rect -625 -754 -465 -707
rect -407 -707 -365 -690
rect -289 -690 -273 -673
rect -163 -673 -55 -657
rect -163 -690 -147 -673
rect -289 -707 -247 -690
rect -407 -754 -247 -707
rect -189 -707 -147 -690
rect -71 -690 -55 -673
rect 55 -673 163 -657
rect 55 -690 71 -673
rect -71 -707 -29 -690
rect -189 -754 -29 -707
rect 29 -707 71 -690
rect 147 -690 163 -673
rect 273 -673 381 -657
rect 273 -690 289 -673
rect 147 -707 189 -690
rect 29 -754 189 -707
rect 247 -707 289 -690
rect 365 -690 381 -673
rect 491 -673 599 -657
rect 491 -690 507 -673
rect 365 -707 407 -690
rect 247 -754 407 -707
rect 465 -707 507 -690
rect 583 -690 599 -673
rect 709 -673 817 -657
rect 709 -690 725 -673
rect 583 -707 625 -690
rect 465 -754 625 -707
rect 683 -707 725 -690
rect 801 -690 817 -673
rect 927 -673 1035 -657
rect 927 -690 943 -673
rect 801 -707 843 -690
rect 683 -754 843 -707
rect 901 -707 943 -690
rect 1019 -690 1035 -673
rect 1019 -707 1061 -690
rect 901 -754 1061 -707
rect -1061 -1201 -901 -1154
rect -1061 -1218 -1019 -1201
rect -1035 -1235 -1019 -1218
rect -943 -1218 -901 -1201
rect -843 -1201 -683 -1154
rect -843 -1218 -801 -1201
rect -943 -1235 -927 -1218
rect -1035 -1251 -927 -1235
rect -817 -1235 -801 -1218
rect -725 -1218 -683 -1201
rect -625 -1201 -465 -1154
rect -625 -1218 -583 -1201
rect -725 -1235 -709 -1218
rect -817 -1251 -709 -1235
rect -599 -1235 -583 -1218
rect -507 -1218 -465 -1201
rect -407 -1201 -247 -1154
rect -407 -1218 -365 -1201
rect -507 -1235 -491 -1218
rect -599 -1251 -491 -1235
rect -381 -1235 -365 -1218
rect -289 -1218 -247 -1201
rect -189 -1201 -29 -1154
rect -189 -1218 -147 -1201
rect -289 -1235 -273 -1218
rect -381 -1251 -273 -1235
rect -163 -1235 -147 -1218
rect -71 -1218 -29 -1201
rect 29 -1201 189 -1154
rect 29 -1218 71 -1201
rect -71 -1235 -55 -1218
rect -163 -1251 -55 -1235
rect 55 -1235 71 -1218
rect 147 -1218 189 -1201
rect 247 -1201 407 -1154
rect 247 -1218 289 -1201
rect 147 -1235 163 -1218
rect 55 -1251 163 -1235
rect 273 -1235 289 -1218
rect 365 -1218 407 -1201
rect 465 -1201 625 -1154
rect 465 -1218 507 -1201
rect 365 -1235 381 -1218
rect 273 -1251 381 -1235
rect 491 -1235 507 -1218
rect 583 -1218 625 -1201
rect 683 -1201 843 -1154
rect 683 -1218 725 -1201
rect 583 -1235 599 -1218
rect 491 -1251 599 -1235
rect 709 -1235 725 -1218
rect 801 -1218 843 -1201
rect 901 -1201 1061 -1154
rect 901 -1218 943 -1201
rect 801 -1235 817 -1218
rect 709 -1251 817 -1235
rect 927 -1235 943 -1218
rect 1019 -1218 1061 -1201
rect 1019 -1235 1035 -1218
rect 927 -1251 1035 -1235
<< polycont >>
rect -1019 1201 -943 1235
rect -801 1201 -725 1235
rect -583 1201 -507 1235
rect -365 1201 -289 1235
rect -147 1201 -71 1235
rect 71 1201 147 1235
rect 289 1201 365 1235
rect 507 1201 583 1235
rect 725 1201 801 1235
rect 943 1201 1019 1235
rect -1019 673 -943 707
rect -801 673 -725 707
rect -583 673 -507 707
rect -365 673 -289 707
rect -147 673 -71 707
rect 71 673 147 707
rect 289 673 365 707
rect 507 673 583 707
rect 725 673 801 707
rect 943 673 1019 707
rect -1019 565 -943 599
rect -801 565 -725 599
rect -583 565 -507 599
rect -365 565 -289 599
rect -147 565 -71 599
rect 71 565 147 599
rect 289 565 365 599
rect 507 565 583 599
rect 725 565 801 599
rect 943 565 1019 599
rect -1019 37 -943 71
rect -801 37 -725 71
rect -583 37 -507 71
rect -365 37 -289 71
rect -147 37 -71 71
rect 71 37 147 71
rect 289 37 365 71
rect 507 37 583 71
rect 725 37 801 71
rect 943 37 1019 71
rect -1019 -71 -943 -37
rect -801 -71 -725 -37
rect -583 -71 -507 -37
rect -365 -71 -289 -37
rect -147 -71 -71 -37
rect 71 -71 147 -37
rect 289 -71 365 -37
rect 507 -71 583 -37
rect 725 -71 801 -37
rect 943 -71 1019 -37
rect -1019 -599 -943 -565
rect -801 -599 -725 -565
rect -583 -599 -507 -565
rect -365 -599 -289 -565
rect -147 -599 -71 -565
rect 71 -599 147 -565
rect 289 -599 365 -565
rect 507 -599 583 -565
rect 725 -599 801 -565
rect 943 -599 1019 -565
rect -1019 -707 -943 -673
rect -801 -707 -725 -673
rect -583 -707 -507 -673
rect -365 -707 -289 -673
rect -147 -707 -71 -673
rect 71 -707 147 -673
rect 289 -707 365 -673
rect 507 -707 583 -673
rect 725 -707 801 -673
rect 943 -707 1019 -673
rect -1019 -1235 -943 -1201
rect -801 -1235 -725 -1201
rect -583 -1235 -507 -1201
rect -365 -1235 -289 -1201
rect -147 -1235 -71 -1201
rect 71 -1235 147 -1201
rect 289 -1235 365 -1201
rect 507 -1235 583 -1201
rect 725 -1235 801 -1201
rect 943 -1235 1019 -1201
<< locali >>
rect -1221 1303 -1125 1337
rect 1125 1303 1221 1337
rect -1221 1241 -1187 1303
rect 1187 1241 1221 1303
rect -1035 1201 -1019 1235
rect -943 1201 -927 1235
rect -817 1201 -801 1235
rect -725 1201 -709 1235
rect -599 1201 -583 1235
rect -507 1201 -491 1235
rect -381 1201 -365 1235
rect -289 1201 -273 1235
rect -163 1201 -147 1235
rect -71 1201 -55 1235
rect 55 1201 71 1235
rect 147 1201 163 1235
rect 273 1201 289 1235
rect 365 1201 381 1235
rect 491 1201 507 1235
rect 583 1201 599 1235
rect 709 1201 725 1235
rect 801 1201 817 1235
rect 927 1201 943 1235
rect 1019 1201 1035 1235
rect -1107 1142 -1073 1158
rect -1107 750 -1073 766
rect -889 1142 -855 1158
rect -889 750 -855 766
rect -671 1142 -637 1158
rect -671 750 -637 766
rect -453 1142 -419 1158
rect -453 750 -419 766
rect -235 1142 -201 1158
rect -235 750 -201 766
rect -17 1142 17 1158
rect -17 750 17 766
rect 201 1142 235 1158
rect 201 750 235 766
rect 419 1142 453 1158
rect 419 750 453 766
rect 637 1142 671 1158
rect 637 750 671 766
rect 855 1142 889 1158
rect 855 750 889 766
rect 1073 1142 1107 1158
rect 1073 750 1107 766
rect -1035 673 -1019 707
rect -943 673 -927 707
rect -817 673 -801 707
rect -725 673 -709 707
rect -599 673 -583 707
rect -507 673 -491 707
rect -381 673 -365 707
rect -289 673 -273 707
rect -163 673 -147 707
rect -71 673 -55 707
rect 55 673 71 707
rect 147 673 163 707
rect 273 673 289 707
rect 365 673 381 707
rect 491 673 507 707
rect 583 673 599 707
rect 709 673 725 707
rect 801 673 817 707
rect 927 673 943 707
rect 1019 673 1035 707
rect -1035 565 -1019 599
rect -943 565 -927 599
rect -817 565 -801 599
rect -725 565 -709 599
rect -599 565 -583 599
rect -507 565 -491 599
rect -381 565 -365 599
rect -289 565 -273 599
rect -163 565 -147 599
rect -71 565 -55 599
rect 55 565 71 599
rect 147 565 163 599
rect 273 565 289 599
rect 365 565 381 599
rect 491 565 507 599
rect 583 565 599 599
rect 709 565 725 599
rect 801 565 817 599
rect 927 565 943 599
rect 1019 565 1035 599
rect -1107 506 -1073 522
rect -1107 114 -1073 130
rect -889 506 -855 522
rect -889 114 -855 130
rect -671 506 -637 522
rect -671 114 -637 130
rect -453 506 -419 522
rect -453 114 -419 130
rect -235 506 -201 522
rect -235 114 -201 130
rect -17 506 17 522
rect -17 114 17 130
rect 201 506 235 522
rect 201 114 235 130
rect 419 506 453 522
rect 419 114 453 130
rect 637 506 671 522
rect 637 114 671 130
rect 855 506 889 522
rect 855 114 889 130
rect 1073 506 1107 522
rect 1073 114 1107 130
rect -1035 37 -1019 71
rect -943 37 -927 71
rect -817 37 -801 71
rect -725 37 -709 71
rect -599 37 -583 71
rect -507 37 -491 71
rect -381 37 -365 71
rect -289 37 -273 71
rect -163 37 -147 71
rect -71 37 -55 71
rect 55 37 71 71
rect 147 37 163 71
rect 273 37 289 71
rect 365 37 381 71
rect 491 37 507 71
rect 583 37 599 71
rect 709 37 725 71
rect 801 37 817 71
rect 927 37 943 71
rect 1019 37 1035 71
rect -1035 -71 -1019 -37
rect -943 -71 -927 -37
rect -817 -71 -801 -37
rect -725 -71 -709 -37
rect -599 -71 -583 -37
rect -507 -71 -491 -37
rect -381 -71 -365 -37
rect -289 -71 -273 -37
rect -163 -71 -147 -37
rect -71 -71 -55 -37
rect 55 -71 71 -37
rect 147 -71 163 -37
rect 273 -71 289 -37
rect 365 -71 381 -37
rect 491 -71 507 -37
rect 583 -71 599 -37
rect 709 -71 725 -37
rect 801 -71 817 -37
rect 927 -71 943 -37
rect 1019 -71 1035 -37
rect -1107 -130 -1073 -114
rect -1107 -522 -1073 -506
rect -889 -130 -855 -114
rect -889 -522 -855 -506
rect -671 -130 -637 -114
rect -671 -522 -637 -506
rect -453 -130 -419 -114
rect -453 -522 -419 -506
rect -235 -130 -201 -114
rect -235 -522 -201 -506
rect -17 -130 17 -114
rect -17 -522 17 -506
rect 201 -130 235 -114
rect 201 -522 235 -506
rect 419 -130 453 -114
rect 419 -522 453 -506
rect 637 -130 671 -114
rect 637 -522 671 -506
rect 855 -130 889 -114
rect 855 -522 889 -506
rect 1073 -130 1107 -114
rect 1073 -522 1107 -506
rect -1035 -599 -1019 -565
rect -943 -599 -927 -565
rect -817 -599 -801 -565
rect -725 -599 -709 -565
rect -599 -599 -583 -565
rect -507 -599 -491 -565
rect -381 -599 -365 -565
rect -289 -599 -273 -565
rect -163 -599 -147 -565
rect -71 -599 -55 -565
rect 55 -599 71 -565
rect 147 -599 163 -565
rect 273 -599 289 -565
rect 365 -599 381 -565
rect 491 -599 507 -565
rect 583 -599 599 -565
rect 709 -599 725 -565
rect 801 -599 817 -565
rect 927 -599 943 -565
rect 1019 -599 1035 -565
rect -1035 -707 -1019 -673
rect -943 -707 -927 -673
rect -817 -707 -801 -673
rect -725 -707 -709 -673
rect -599 -707 -583 -673
rect -507 -707 -491 -673
rect -381 -707 -365 -673
rect -289 -707 -273 -673
rect -163 -707 -147 -673
rect -71 -707 -55 -673
rect 55 -707 71 -673
rect 147 -707 163 -673
rect 273 -707 289 -673
rect 365 -707 381 -673
rect 491 -707 507 -673
rect 583 -707 599 -673
rect 709 -707 725 -673
rect 801 -707 817 -673
rect 927 -707 943 -673
rect 1019 -707 1035 -673
rect -1107 -766 -1073 -750
rect -1107 -1158 -1073 -1142
rect -889 -766 -855 -750
rect -889 -1158 -855 -1142
rect -671 -766 -637 -750
rect -671 -1158 -637 -1142
rect -453 -766 -419 -750
rect -453 -1158 -419 -1142
rect -235 -766 -201 -750
rect -235 -1158 -201 -1142
rect -17 -766 17 -750
rect -17 -1158 17 -1142
rect 201 -766 235 -750
rect 201 -1158 235 -1142
rect 419 -766 453 -750
rect 419 -1158 453 -1142
rect 637 -766 671 -750
rect 637 -1158 671 -1142
rect 855 -766 889 -750
rect 855 -1158 889 -1142
rect 1073 -766 1107 -750
rect 1073 -1158 1107 -1142
rect -1035 -1235 -1019 -1201
rect -943 -1235 -927 -1201
rect -817 -1235 -801 -1201
rect -725 -1235 -709 -1201
rect -599 -1235 -583 -1201
rect -507 -1235 -491 -1201
rect -381 -1235 -365 -1201
rect -289 -1235 -273 -1201
rect -163 -1235 -147 -1201
rect -71 -1235 -55 -1201
rect 55 -1235 71 -1201
rect 147 -1235 163 -1201
rect 273 -1235 289 -1201
rect 365 -1235 381 -1201
rect 491 -1235 507 -1201
rect 583 -1235 599 -1201
rect 709 -1235 725 -1201
rect 801 -1235 817 -1201
rect 927 -1235 943 -1201
rect 1019 -1235 1035 -1201
rect -1221 -1303 -1187 -1241
rect 1187 -1303 1221 -1241
rect -1221 -1337 -1125 -1303
rect 1125 -1337 1221 -1303
<< viali >>
rect -1013 1201 -949 1235
rect -795 1201 -731 1235
rect -577 1201 -513 1235
rect -359 1201 -295 1235
rect -141 1201 -77 1235
rect 77 1201 141 1235
rect 295 1201 359 1235
rect 513 1201 577 1235
rect 731 1201 795 1235
rect 949 1201 1013 1235
rect -1107 766 -1073 1142
rect -889 766 -855 1142
rect -671 766 -637 1142
rect -453 766 -419 1142
rect -235 766 -201 1142
rect -17 766 17 1142
rect 201 766 235 1142
rect 419 766 453 1142
rect 637 766 671 1142
rect 855 766 889 1142
rect 1073 766 1107 1142
rect -1013 673 -949 707
rect -795 673 -731 707
rect -577 673 -513 707
rect -359 673 -295 707
rect -141 673 -77 707
rect 77 673 141 707
rect 295 673 359 707
rect 513 673 577 707
rect 731 673 795 707
rect 949 673 1013 707
rect -1013 565 -949 599
rect -795 565 -731 599
rect -577 565 -513 599
rect -359 565 -295 599
rect -141 565 -77 599
rect 77 565 141 599
rect 295 565 359 599
rect 513 565 577 599
rect 731 565 795 599
rect 949 565 1013 599
rect -1107 130 -1073 506
rect -889 130 -855 506
rect -671 130 -637 506
rect -453 130 -419 506
rect -235 130 -201 506
rect -17 130 17 506
rect 201 130 235 506
rect 419 130 453 506
rect 637 130 671 506
rect 855 130 889 506
rect 1073 130 1107 506
rect -1013 37 -949 71
rect -795 37 -731 71
rect -577 37 -513 71
rect -359 37 -295 71
rect -141 37 -77 71
rect 77 37 141 71
rect 295 37 359 71
rect 513 37 577 71
rect 731 37 795 71
rect 949 37 1013 71
rect -1013 -71 -949 -37
rect -795 -71 -731 -37
rect -577 -71 -513 -37
rect -359 -71 -295 -37
rect -141 -71 -77 -37
rect 77 -71 141 -37
rect 295 -71 359 -37
rect 513 -71 577 -37
rect 731 -71 795 -37
rect 949 -71 1013 -37
rect -1107 -506 -1073 -130
rect -889 -506 -855 -130
rect -671 -506 -637 -130
rect -453 -506 -419 -130
rect -235 -506 -201 -130
rect -17 -506 17 -130
rect 201 -506 235 -130
rect 419 -506 453 -130
rect 637 -506 671 -130
rect 855 -506 889 -130
rect 1073 -506 1107 -130
rect -1013 -599 -949 -565
rect -795 -599 -731 -565
rect -577 -599 -513 -565
rect -359 -599 -295 -565
rect -141 -599 -77 -565
rect 77 -599 141 -565
rect 295 -599 359 -565
rect 513 -599 577 -565
rect 731 -599 795 -565
rect 949 -599 1013 -565
rect -1013 -707 -949 -673
rect -795 -707 -731 -673
rect -577 -707 -513 -673
rect -359 -707 -295 -673
rect -141 -707 -77 -673
rect 77 -707 141 -673
rect 295 -707 359 -673
rect 513 -707 577 -673
rect 731 -707 795 -673
rect 949 -707 1013 -673
rect -1107 -1142 -1073 -766
rect -889 -1142 -855 -766
rect -671 -1142 -637 -766
rect -453 -1142 -419 -766
rect -235 -1142 -201 -766
rect -17 -1142 17 -766
rect 201 -1142 235 -766
rect 419 -1142 453 -766
rect 637 -1142 671 -766
rect 855 -1142 889 -766
rect 1073 -1142 1107 -766
rect -1013 -1235 -949 -1201
rect -795 -1235 -731 -1201
rect -577 -1235 -513 -1201
rect -359 -1235 -295 -1201
rect -141 -1235 -77 -1201
rect 77 -1235 141 -1201
rect 295 -1235 359 -1201
rect 513 -1235 577 -1201
rect 731 -1235 795 -1201
rect 949 -1235 1013 -1201
<< metal1 >>
rect -1025 1235 -937 1241
rect -1025 1201 -1013 1235
rect -949 1201 -937 1235
rect -1025 1195 -937 1201
rect -807 1235 -719 1241
rect -807 1201 -795 1235
rect -731 1201 -719 1235
rect -807 1195 -719 1201
rect -589 1235 -501 1241
rect -589 1201 -577 1235
rect -513 1201 -501 1235
rect -589 1195 -501 1201
rect -371 1235 -283 1241
rect -371 1201 -359 1235
rect -295 1201 -283 1235
rect -371 1195 -283 1201
rect -153 1235 -65 1241
rect -153 1201 -141 1235
rect -77 1201 -65 1235
rect -153 1195 -65 1201
rect 65 1235 153 1241
rect 65 1201 77 1235
rect 141 1201 153 1235
rect 65 1195 153 1201
rect 283 1235 371 1241
rect 283 1201 295 1235
rect 359 1201 371 1235
rect 283 1195 371 1201
rect 501 1235 589 1241
rect 501 1201 513 1235
rect 577 1201 589 1235
rect 501 1195 589 1201
rect 719 1235 807 1241
rect 719 1201 731 1235
rect 795 1201 807 1235
rect 719 1195 807 1201
rect 937 1235 1025 1241
rect 937 1201 949 1235
rect 1013 1201 1025 1235
rect 937 1195 1025 1201
rect -1113 1142 -1067 1154
rect -1113 766 -1107 1142
rect -1073 766 -1067 1142
rect -1113 754 -1067 766
rect -895 1142 -849 1154
rect -895 766 -889 1142
rect -855 766 -849 1142
rect -895 754 -849 766
rect -677 1142 -631 1154
rect -677 766 -671 1142
rect -637 766 -631 1142
rect -677 754 -631 766
rect -459 1142 -413 1154
rect -459 766 -453 1142
rect -419 766 -413 1142
rect -459 754 -413 766
rect -241 1142 -195 1154
rect -241 766 -235 1142
rect -201 766 -195 1142
rect -241 754 -195 766
rect -23 1142 23 1154
rect -23 766 -17 1142
rect 17 766 23 1142
rect -23 754 23 766
rect 195 1142 241 1154
rect 195 766 201 1142
rect 235 766 241 1142
rect 195 754 241 766
rect 413 1142 459 1154
rect 413 766 419 1142
rect 453 766 459 1142
rect 413 754 459 766
rect 631 1142 677 1154
rect 631 766 637 1142
rect 671 766 677 1142
rect 631 754 677 766
rect 849 1142 895 1154
rect 849 766 855 1142
rect 889 766 895 1142
rect 849 754 895 766
rect 1067 1142 1113 1154
rect 1067 766 1073 1142
rect 1107 766 1113 1142
rect 1067 754 1113 766
rect -1025 707 -937 713
rect -1025 673 -1013 707
rect -949 673 -937 707
rect -1025 667 -937 673
rect -807 707 -719 713
rect -807 673 -795 707
rect -731 673 -719 707
rect -807 667 -719 673
rect -589 707 -501 713
rect -589 673 -577 707
rect -513 673 -501 707
rect -589 667 -501 673
rect -371 707 -283 713
rect -371 673 -359 707
rect -295 673 -283 707
rect -371 667 -283 673
rect -153 707 -65 713
rect -153 673 -141 707
rect -77 673 -65 707
rect -153 667 -65 673
rect 65 707 153 713
rect 65 673 77 707
rect 141 673 153 707
rect 65 667 153 673
rect 283 707 371 713
rect 283 673 295 707
rect 359 673 371 707
rect 283 667 371 673
rect 501 707 589 713
rect 501 673 513 707
rect 577 673 589 707
rect 501 667 589 673
rect 719 707 807 713
rect 719 673 731 707
rect 795 673 807 707
rect 719 667 807 673
rect 937 707 1025 713
rect 937 673 949 707
rect 1013 673 1025 707
rect 937 667 1025 673
rect -1025 599 -937 605
rect -1025 565 -1013 599
rect -949 565 -937 599
rect -1025 559 -937 565
rect -807 599 -719 605
rect -807 565 -795 599
rect -731 565 -719 599
rect -807 559 -719 565
rect -589 599 -501 605
rect -589 565 -577 599
rect -513 565 -501 599
rect -589 559 -501 565
rect -371 599 -283 605
rect -371 565 -359 599
rect -295 565 -283 599
rect -371 559 -283 565
rect -153 599 -65 605
rect -153 565 -141 599
rect -77 565 -65 599
rect -153 559 -65 565
rect 65 599 153 605
rect 65 565 77 599
rect 141 565 153 599
rect 65 559 153 565
rect 283 599 371 605
rect 283 565 295 599
rect 359 565 371 599
rect 283 559 371 565
rect 501 599 589 605
rect 501 565 513 599
rect 577 565 589 599
rect 501 559 589 565
rect 719 599 807 605
rect 719 565 731 599
rect 795 565 807 599
rect 719 559 807 565
rect 937 599 1025 605
rect 937 565 949 599
rect 1013 565 1025 599
rect 937 559 1025 565
rect -1113 506 -1067 518
rect -1113 130 -1107 506
rect -1073 130 -1067 506
rect -1113 118 -1067 130
rect -895 506 -849 518
rect -895 130 -889 506
rect -855 130 -849 506
rect -895 118 -849 130
rect -677 506 -631 518
rect -677 130 -671 506
rect -637 130 -631 506
rect -677 118 -631 130
rect -459 506 -413 518
rect -459 130 -453 506
rect -419 130 -413 506
rect -459 118 -413 130
rect -241 506 -195 518
rect -241 130 -235 506
rect -201 130 -195 506
rect -241 118 -195 130
rect -23 506 23 518
rect -23 130 -17 506
rect 17 130 23 506
rect -23 118 23 130
rect 195 506 241 518
rect 195 130 201 506
rect 235 130 241 506
rect 195 118 241 130
rect 413 506 459 518
rect 413 130 419 506
rect 453 130 459 506
rect 413 118 459 130
rect 631 506 677 518
rect 631 130 637 506
rect 671 130 677 506
rect 631 118 677 130
rect 849 506 895 518
rect 849 130 855 506
rect 889 130 895 506
rect 849 118 895 130
rect 1067 506 1113 518
rect 1067 130 1073 506
rect 1107 130 1113 506
rect 1067 118 1113 130
rect -1025 71 -937 77
rect -1025 37 -1013 71
rect -949 37 -937 71
rect -1025 31 -937 37
rect -807 71 -719 77
rect -807 37 -795 71
rect -731 37 -719 71
rect -807 31 -719 37
rect -589 71 -501 77
rect -589 37 -577 71
rect -513 37 -501 71
rect -589 31 -501 37
rect -371 71 -283 77
rect -371 37 -359 71
rect -295 37 -283 71
rect -371 31 -283 37
rect -153 71 -65 77
rect -153 37 -141 71
rect -77 37 -65 71
rect -153 31 -65 37
rect 65 71 153 77
rect 65 37 77 71
rect 141 37 153 71
rect 65 31 153 37
rect 283 71 371 77
rect 283 37 295 71
rect 359 37 371 71
rect 283 31 371 37
rect 501 71 589 77
rect 501 37 513 71
rect 577 37 589 71
rect 501 31 589 37
rect 719 71 807 77
rect 719 37 731 71
rect 795 37 807 71
rect 719 31 807 37
rect 937 71 1025 77
rect 937 37 949 71
rect 1013 37 1025 71
rect 937 31 1025 37
rect -1025 -37 -937 -31
rect -1025 -71 -1013 -37
rect -949 -71 -937 -37
rect -1025 -77 -937 -71
rect -807 -37 -719 -31
rect -807 -71 -795 -37
rect -731 -71 -719 -37
rect -807 -77 -719 -71
rect -589 -37 -501 -31
rect -589 -71 -577 -37
rect -513 -71 -501 -37
rect -589 -77 -501 -71
rect -371 -37 -283 -31
rect -371 -71 -359 -37
rect -295 -71 -283 -37
rect -371 -77 -283 -71
rect -153 -37 -65 -31
rect -153 -71 -141 -37
rect -77 -71 -65 -37
rect -153 -77 -65 -71
rect 65 -37 153 -31
rect 65 -71 77 -37
rect 141 -71 153 -37
rect 65 -77 153 -71
rect 283 -37 371 -31
rect 283 -71 295 -37
rect 359 -71 371 -37
rect 283 -77 371 -71
rect 501 -37 589 -31
rect 501 -71 513 -37
rect 577 -71 589 -37
rect 501 -77 589 -71
rect 719 -37 807 -31
rect 719 -71 731 -37
rect 795 -71 807 -37
rect 719 -77 807 -71
rect 937 -37 1025 -31
rect 937 -71 949 -37
rect 1013 -71 1025 -37
rect 937 -77 1025 -71
rect -1113 -130 -1067 -118
rect -1113 -506 -1107 -130
rect -1073 -506 -1067 -130
rect -1113 -518 -1067 -506
rect -895 -130 -849 -118
rect -895 -506 -889 -130
rect -855 -506 -849 -130
rect -895 -518 -849 -506
rect -677 -130 -631 -118
rect -677 -506 -671 -130
rect -637 -506 -631 -130
rect -677 -518 -631 -506
rect -459 -130 -413 -118
rect -459 -506 -453 -130
rect -419 -506 -413 -130
rect -459 -518 -413 -506
rect -241 -130 -195 -118
rect -241 -506 -235 -130
rect -201 -506 -195 -130
rect -241 -518 -195 -506
rect -23 -130 23 -118
rect -23 -506 -17 -130
rect 17 -506 23 -130
rect -23 -518 23 -506
rect 195 -130 241 -118
rect 195 -506 201 -130
rect 235 -506 241 -130
rect 195 -518 241 -506
rect 413 -130 459 -118
rect 413 -506 419 -130
rect 453 -506 459 -130
rect 413 -518 459 -506
rect 631 -130 677 -118
rect 631 -506 637 -130
rect 671 -506 677 -130
rect 631 -518 677 -506
rect 849 -130 895 -118
rect 849 -506 855 -130
rect 889 -506 895 -130
rect 849 -518 895 -506
rect 1067 -130 1113 -118
rect 1067 -506 1073 -130
rect 1107 -506 1113 -130
rect 1067 -518 1113 -506
rect -1025 -565 -937 -559
rect -1025 -599 -1013 -565
rect -949 -599 -937 -565
rect -1025 -605 -937 -599
rect -807 -565 -719 -559
rect -807 -599 -795 -565
rect -731 -599 -719 -565
rect -807 -605 -719 -599
rect -589 -565 -501 -559
rect -589 -599 -577 -565
rect -513 -599 -501 -565
rect -589 -605 -501 -599
rect -371 -565 -283 -559
rect -371 -599 -359 -565
rect -295 -599 -283 -565
rect -371 -605 -283 -599
rect -153 -565 -65 -559
rect -153 -599 -141 -565
rect -77 -599 -65 -565
rect -153 -605 -65 -599
rect 65 -565 153 -559
rect 65 -599 77 -565
rect 141 -599 153 -565
rect 65 -605 153 -599
rect 283 -565 371 -559
rect 283 -599 295 -565
rect 359 -599 371 -565
rect 283 -605 371 -599
rect 501 -565 589 -559
rect 501 -599 513 -565
rect 577 -599 589 -565
rect 501 -605 589 -599
rect 719 -565 807 -559
rect 719 -599 731 -565
rect 795 -599 807 -565
rect 719 -605 807 -599
rect 937 -565 1025 -559
rect 937 -599 949 -565
rect 1013 -599 1025 -565
rect 937 -605 1025 -599
rect -1025 -673 -937 -667
rect -1025 -707 -1013 -673
rect -949 -707 -937 -673
rect -1025 -713 -937 -707
rect -807 -673 -719 -667
rect -807 -707 -795 -673
rect -731 -707 -719 -673
rect -807 -713 -719 -707
rect -589 -673 -501 -667
rect -589 -707 -577 -673
rect -513 -707 -501 -673
rect -589 -713 -501 -707
rect -371 -673 -283 -667
rect -371 -707 -359 -673
rect -295 -707 -283 -673
rect -371 -713 -283 -707
rect -153 -673 -65 -667
rect -153 -707 -141 -673
rect -77 -707 -65 -673
rect -153 -713 -65 -707
rect 65 -673 153 -667
rect 65 -707 77 -673
rect 141 -707 153 -673
rect 65 -713 153 -707
rect 283 -673 371 -667
rect 283 -707 295 -673
rect 359 -707 371 -673
rect 283 -713 371 -707
rect 501 -673 589 -667
rect 501 -707 513 -673
rect 577 -707 589 -673
rect 501 -713 589 -707
rect 719 -673 807 -667
rect 719 -707 731 -673
rect 795 -707 807 -673
rect 719 -713 807 -707
rect 937 -673 1025 -667
rect 937 -707 949 -673
rect 1013 -707 1025 -673
rect 937 -713 1025 -707
rect -1113 -766 -1067 -754
rect -1113 -1142 -1107 -766
rect -1073 -1142 -1067 -766
rect -1113 -1154 -1067 -1142
rect -895 -766 -849 -754
rect -895 -1142 -889 -766
rect -855 -1142 -849 -766
rect -895 -1154 -849 -1142
rect -677 -766 -631 -754
rect -677 -1142 -671 -766
rect -637 -1142 -631 -766
rect -677 -1154 -631 -1142
rect -459 -766 -413 -754
rect -459 -1142 -453 -766
rect -419 -1142 -413 -766
rect -459 -1154 -413 -1142
rect -241 -766 -195 -754
rect -241 -1142 -235 -766
rect -201 -1142 -195 -766
rect -241 -1154 -195 -1142
rect -23 -766 23 -754
rect -23 -1142 -17 -766
rect 17 -1142 23 -766
rect -23 -1154 23 -1142
rect 195 -766 241 -754
rect 195 -1142 201 -766
rect 235 -1142 241 -766
rect 195 -1154 241 -1142
rect 413 -766 459 -754
rect 413 -1142 419 -766
rect 453 -1142 459 -766
rect 413 -1154 459 -1142
rect 631 -766 677 -754
rect 631 -1142 637 -766
rect 671 -1142 677 -766
rect 631 -1154 677 -1142
rect 849 -766 895 -754
rect 849 -1142 855 -766
rect 889 -1142 895 -766
rect 849 -1154 895 -1142
rect 1067 -766 1113 -754
rect 1067 -1142 1073 -766
rect 1107 -1142 1113 -766
rect 1067 -1154 1113 -1142
rect -1025 -1201 -937 -1195
rect -1025 -1235 -1013 -1201
rect -949 -1235 -937 -1201
rect -1025 -1241 -937 -1235
rect -807 -1201 -719 -1195
rect -807 -1235 -795 -1201
rect -731 -1235 -719 -1201
rect -807 -1241 -719 -1235
rect -589 -1201 -501 -1195
rect -589 -1235 -577 -1201
rect -513 -1235 -501 -1201
rect -589 -1241 -501 -1235
rect -371 -1201 -283 -1195
rect -371 -1235 -359 -1201
rect -295 -1235 -283 -1201
rect -371 -1241 -283 -1235
rect -153 -1201 -65 -1195
rect -153 -1235 -141 -1201
rect -77 -1235 -65 -1201
rect -153 -1241 -65 -1235
rect 65 -1201 153 -1195
rect 65 -1235 77 -1201
rect 141 -1235 153 -1201
rect 65 -1241 153 -1235
rect 283 -1201 371 -1195
rect 283 -1235 295 -1201
rect 359 -1235 371 -1201
rect 283 -1241 371 -1235
rect 501 -1201 589 -1195
rect 501 -1235 513 -1201
rect 577 -1235 589 -1201
rect 501 -1241 589 -1235
rect 719 -1201 807 -1195
rect 719 -1235 731 -1201
rect 795 -1235 807 -1201
rect 719 -1241 807 -1235
rect 937 -1201 1025 -1195
rect 937 -1235 949 -1201
rect 1013 -1235 1025 -1201
rect 937 -1241 1025 -1235
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -1204 -1320 1204 1320
string parameters w 2 l 0.8 m 4 nf 10 diffcov 100 polycov 60 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viagl 0 viagr 0 viagt 0 viagb 0 viagate 50 viadrn 100 viasrc 100
string library sky130
<< end >>
