magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect -4660 -4274 4307 3538
<< nwell >>
rect -3358 -906 2840 2026
rect -3358 -2050 102 -906
rect -3358 -2066 -1014 -2050
rect 76 -2066 102 -2050
<< pwell >>
rect 866 -1502 2276 -1350
rect 866 -2608 1018 -1502
rect 2124 -2608 2276 -1502
rect 866 -2760 2276 -2608
<< psubdiff >>
rect 892 -1409 2250 -1376
rect 892 -1443 1087 -1409
rect 1121 -1443 1155 -1409
rect 1189 -1443 1223 -1409
rect 1257 -1443 1291 -1409
rect 1325 -1443 1359 -1409
rect 1393 -1443 1427 -1409
rect 1461 -1443 1495 -1409
rect 1529 -1443 1563 -1409
rect 1597 -1443 1631 -1409
rect 1665 -1443 1699 -1409
rect 1733 -1443 1767 -1409
rect 1801 -1443 1835 -1409
rect 1869 -1443 1903 -1409
rect 1937 -1443 1971 -1409
rect 2005 -1443 2250 -1409
rect 892 -1476 2250 -1443
rect 892 -1564 992 -1476
rect 892 -1598 925 -1564
rect 959 -1598 992 -1564
rect 892 -1632 992 -1598
rect 892 -1666 925 -1632
rect 959 -1666 992 -1632
rect 2150 -1568 2250 -1476
rect 2150 -1602 2183 -1568
rect 2217 -1602 2250 -1568
rect 2150 -1636 2250 -1602
rect 892 -1700 992 -1666
rect 892 -1734 925 -1700
rect 959 -1734 992 -1700
rect 892 -1768 992 -1734
rect 892 -1802 925 -1768
rect 959 -1802 992 -1768
rect 892 -1836 992 -1802
rect 892 -1870 925 -1836
rect 959 -1870 992 -1836
rect 2150 -1670 2183 -1636
rect 2217 -1670 2250 -1636
rect 2150 -1704 2250 -1670
rect 2150 -1738 2183 -1704
rect 2217 -1738 2250 -1704
rect 2150 -1772 2250 -1738
rect 2150 -1806 2183 -1772
rect 2217 -1806 2250 -1772
rect 2150 -1840 2250 -1806
rect 892 -1904 992 -1870
rect 892 -1938 925 -1904
rect 959 -1938 992 -1904
rect 892 -1972 992 -1938
rect 2150 -1874 2183 -1840
rect 2217 -1874 2250 -1840
rect 2150 -1908 2250 -1874
rect 2150 -1942 2183 -1908
rect 2217 -1942 2250 -1908
rect 892 -2006 925 -1972
rect 959 -2006 992 -1972
rect 892 -2040 992 -2006
rect 892 -2074 925 -2040
rect 959 -2074 992 -2040
rect 892 -2634 992 -2074
rect 2150 -1976 2250 -1942
rect 2150 -2010 2183 -1976
rect 2217 -2010 2250 -1976
rect 2150 -2044 2250 -2010
rect 2150 -2078 2183 -2044
rect 2217 -2078 2250 -2044
rect 2150 -2112 2250 -2078
rect 2150 -2146 2183 -2112
rect 2217 -2146 2250 -2112
rect 2150 -2634 2250 -2146
rect 892 -2667 2250 -2634
rect 892 -2701 1081 -2667
rect 1115 -2701 1149 -2667
rect 1183 -2701 1217 -2667
rect 1251 -2701 1285 -2667
rect 1319 -2701 1353 -2667
rect 1387 -2701 1421 -2667
rect 1455 -2701 1489 -2667
rect 1523 -2701 1557 -2667
rect 1591 -2701 1625 -2667
rect 1659 -2701 1693 -2667
rect 1727 -2701 1761 -2667
rect 1795 -2701 1829 -2667
rect 1863 -2701 1897 -2667
rect 1931 -2701 1965 -2667
rect 1999 -2701 2250 -2667
rect 892 -2734 2250 -2701
<< nsubdiff >>
rect -3322 1957 42 1990
rect -3322 1923 -3153 1957
rect -3119 1923 -3085 1957
rect -3051 1923 -3017 1957
rect -2983 1923 -2949 1957
rect -2915 1923 -2881 1957
rect -2847 1923 -2813 1957
rect -2779 1923 -2745 1957
rect -2711 1923 -2677 1957
rect -2643 1923 -2609 1957
rect -2575 1923 -2541 1957
rect -2507 1923 -2473 1957
rect -2439 1923 -2405 1957
rect -2371 1923 -2337 1957
rect -2303 1923 -2269 1957
rect -2235 1923 -2201 1957
rect -2167 1923 -2133 1957
rect -2099 1923 -2065 1957
rect -2031 1923 -1997 1957
rect -1963 1923 -1929 1957
rect -1895 1923 -1861 1957
rect -1827 1923 -1793 1957
rect -1759 1923 -1725 1957
rect -1691 1923 -1657 1957
rect -1623 1923 -1589 1957
rect -1555 1923 -1521 1957
rect -1487 1923 -1453 1957
rect -1419 1923 -1385 1957
rect -1351 1923 -1317 1957
rect -1283 1923 -1249 1957
rect -1215 1923 -1181 1957
rect -1147 1923 -1113 1957
rect -1079 1923 -1045 1957
rect -1011 1923 -977 1957
rect -943 1923 -909 1957
rect -875 1923 -841 1957
rect -807 1923 -773 1957
rect -739 1923 -705 1957
rect -671 1923 -637 1957
rect -603 1923 -569 1957
rect -535 1923 -501 1957
rect -467 1923 -433 1957
rect -399 1923 -365 1957
rect -331 1923 -297 1957
rect -263 1923 -229 1957
rect -195 1923 -161 1957
rect -127 1923 42 1957
rect -3322 1890 42 1923
rect -3322 1797 -3222 1890
rect -3322 1763 -3289 1797
rect -3255 1763 -3222 1797
rect -3322 1729 -3222 1763
rect -3322 1695 -3289 1729
rect -3255 1695 -3222 1729
rect -3322 1661 -3222 1695
rect -3322 1627 -3289 1661
rect -3255 1627 -3222 1661
rect -3322 1593 -3222 1627
rect -3322 1559 -3289 1593
rect -3255 1559 -3222 1593
rect -3322 1525 -3222 1559
rect -3322 1491 -3289 1525
rect -3255 1491 -3222 1525
rect -3322 1457 -3222 1491
rect -3322 1423 -3289 1457
rect -3255 1423 -3222 1457
rect -3322 1389 -3222 1423
rect -3322 1355 -3289 1389
rect -3255 1355 -3222 1389
rect -3322 1321 -3222 1355
rect -3322 1287 -3289 1321
rect -3255 1287 -3222 1321
rect -3322 1253 -3222 1287
rect -3322 1219 -3289 1253
rect -3255 1219 -3222 1253
rect -3322 1185 -3222 1219
rect -3322 1151 -3289 1185
rect -3255 1151 -3222 1185
rect -3322 1117 -3222 1151
rect -3322 1083 -3289 1117
rect -3255 1083 -3222 1117
rect -3322 1049 -3222 1083
rect -3322 1015 -3289 1049
rect -3255 1015 -3222 1049
rect -3322 981 -3222 1015
rect -3322 947 -3289 981
rect -3255 947 -3222 981
rect -3322 913 -3222 947
rect -3322 879 -3289 913
rect -3255 879 -3222 913
rect -3322 845 -3222 879
rect -3322 811 -3289 845
rect -3255 811 -3222 845
rect -3322 777 -3222 811
rect -3322 743 -3289 777
rect -3255 743 -3222 777
rect -3322 709 -3222 743
rect -3322 675 -3289 709
rect -3255 675 -3222 709
rect -3322 641 -3222 675
rect -3322 607 -3289 641
rect -3255 607 -3222 641
rect -3322 573 -3222 607
rect -3322 539 -3289 573
rect -3255 539 -3222 573
rect -3322 505 -3222 539
rect -3322 471 -3289 505
rect -3255 471 -3222 505
rect -3322 437 -3222 471
rect -3322 403 -3289 437
rect -3255 403 -3222 437
rect -3322 369 -3222 403
rect -3322 335 -3289 369
rect -3255 335 -3222 369
rect -3322 301 -3222 335
rect -3322 267 -3289 301
rect -3255 267 -3222 301
rect -3322 233 -3222 267
rect -3322 199 -3289 233
rect -3255 199 -3222 233
rect -3322 165 -3222 199
rect -3322 131 -3289 165
rect -3255 131 -3222 165
rect -3322 97 -3222 131
rect -3322 63 -3289 97
rect -3255 63 -3222 97
rect -3322 29 -3222 63
rect -3322 -5 -3289 29
rect -3255 -5 -3222 29
rect -3322 -39 -3222 -5
rect -3322 -73 -3289 -39
rect -3255 -73 -3222 -39
rect -3322 -107 -3222 -73
rect -3322 -141 -3289 -107
rect -3255 -141 -3222 -107
rect -3322 -175 -3222 -141
rect -3322 -209 -3289 -175
rect -3255 -209 -3222 -175
rect -3322 -243 -3222 -209
rect -3322 -277 -3289 -243
rect -3255 -277 -3222 -243
rect -3322 -311 -3222 -277
rect -3322 -345 -3289 -311
rect -3255 -345 -3222 -311
rect -3322 -379 -3222 -345
rect -3322 -413 -3289 -379
rect -3255 -413 -3222 -379
rect -3322 -447 -3222 -413
rect -3322 -481 -3289 -447
rect -3255 -481 -3222 -447
rect -3322 -515 -3222 -481
rect -3322 -549 -3289 -515
rect -3255 -549 -3222 -515
rect -3322 -583 -3222 -549
rect -3322 -617 -3289 -583
rect -3255 -617 -3222 -583
rect -3322 -651 -3222 -617
rect -3322 -685 -3289 -651
rect -3255 -685 -3222 -651
rect -3322 -719 -3222 -685
rect -3322 -753 -3289 -719
rect -3255 -753 -3222 -719
rect -3322 -787 -3222 -753
rect -3322 -821 -3289 -787
rect -3255 -821 -3222 -787
rect -3322 -855 -3222 -821
rect -3322 -889 -3289 -855
rect -3255 -889 -3222 -855
rect -3322 -923 -3222 -889
rect -3322 -957 -3289 -923
rect -3255 -957 -3222 -923
rect -3322 -991 -3222 -957
rect -3322 -1025 -3289 -991
rect -3255 -1025 -3222 -991
rect -3322 -1059 -3222 -1025
rect -3322 -1093 -3289 -1059
rect -3255 -1093 -3222 -1059
rect -3322 -1127 -3222 -1093
rect -3322 -1161 -3289 -1127
rect -3255 -1161 -3222 -1127
rect -3322 -1254 -3222 -1161
rect -58 1797 42 1890
rect -58 1763 -25 1797
rect 9 1763 42 1797
rect -58 1729 42 1763
rect -58 1695 -25 1729
rect 9 1695 42 1729
rect -58 1661 42 1695
rect -58 1627 -25 1661
rect 9 1627 42 1661
rect -58 1593 42 1627
rect -58 1559 -25 1593
rect 9 1559 42 1593
rect -58 1525 42 1559
rect -58 1491 -25 1525
rect 9 1491 42 1525
rect -58 1457 42 1491
rect -58 1423 -25 1457
rect 9 1423 42 1457
rect -58 1389 42 1423
rect -58 1355 -25 1389
rect 9 1355 42 1389
rect -58 1321 42 1355
rect -58 1287 -25 1321
rect 9 1287 42 1321
rect -58 1253 42 1287
rect -58 1219 -25 1253
rect 9 1219 42 1253
rect -58 1185 42 1219
rect -58 1151 -25 1185
rect 9 1151 42 1185
rect -58 1117 42 1151
rect -58 1083 -25 1117
rect 9 1083 42 1117
rect -58 1049 42 1083
rect -58 1015 -25 1049
rect 9 1015 42 1049
rect -58 981 42 1015
rect -58 947 -25 981
rect 9 947 42 981
rect -58 913 42 947
rect -58 879 -25 913
rect 9 879 42 913
rect -58 845 42 879
rect -58 811 -25 845
rect 9 811 42 845
rect -58 777 42 811
rect -58 743 -25 777
rect 9 743 42 777
rect -58 709 42 743
rect -58 675 -25 709
rect 9 675 42 709
rect -58 641 42 675
rect -58 607 -25 641
rect 9 607 42 641
rect -58 573 42 607
rect -58 539 -25 573
rect 9 539 42 573
rect -58 505 42 539
rect -58 471 -25 505
rect 9 471 42 505
rect -58 437 42 471
rect -58 403 -25 437
rect 9 403 42 437
rect -58 369 42 403
rect -58 335 -25 369
rect 9 335 42 369
rect -58 301 42 335
rect -58 267 -25 301
rect 9 267 42 301
rect -58 233 42 267
rect -58 199 -25 233
rect 9 199 42 233
rect -58 165 42 199
rect -58 131 -25 165
rect 9 131 42 165
rect -58 97 42 131
rect -58 63 -25 97
rect 9 63 42 97
rect -58 29 42 63
rect -58 -5 -25 29
rect 9 -5 42 29
rect -58 -39 42 -5
rect -58 -73 -25 -39
rect 9 -73 42 -39
rect -58 -107 42 -73
rect -58 -141 -25 -107
rect 9 -141 42 -107
rect -58 -175 42 -141
rect -58 -209 -25 -175
rect 9 -209 42 -175
rect -58 -243 42 -209
rect -58 -277 -25 -243
rect 9 -277 42 -243
rect -58 -311 42 -277
rect -58 -345 -25 -311
rect 9 -345 42 -311
rect -58 -379 42 -345
rect -58 -413 -25 -379
rect 9 -413 42 -379
rect -58 -447 42 -413
rect -58 -481 -25 -447
rect 9 -481 42 -447
rect -58 -515 42 -481
rect -58 -549 -25 -515
rect 9 -549 42 -515
rect -58 -583 42 -549
rect 380 1957 2784 1990
rect 380 1923 545 1957
rect 579 1923 613 1957
rect 647 1923 681 1957
rect 715 1923 749 1957
rect 783 1923 817 1957
rect 851 1923 885 1957
rect 919 1923 953 1957
rect 987 1923 1021 1957
rect 1055 1923 1089 1957
rect 1123 1923 1157 1957
rect 1191 1923 1225 1957
rect 1259 1923 1293 1957
rect 1327 1923 1361 1957
rect 1395 1923 1429 1957
rect 1463 1923 1497 1957
rect 1531 1923 1565 1957
rect 1599 1923 1633 1957
rect 1667 1923 1701 1957
rect 1735 1923 1769 1957
rect 1803 1923 1837 1957
rect 1871 1923 1905 1957
rect 1939 1923 1973 1957
rect 2007 1923 2041 1957
rect 2075 1923 2109 1957
rect 2143 1923 2177 1957
rect 2211 1923 2245 1957
rect 2279 1923 2313 1957
rect 2347 1923 2381 1957
rect 2415 1923 2449 1957
rect 2483 1923 2517 1957
rect 2551 1923 2585 1957
rect 2619 1923 2784 1957
rect 380 1890 2784 1923
rect 380 1820 480 1890
rect 380 1786 413 1820
rect 447 1786 480 1820
rect 380 1752 480 1786
rect 380 1718 413 1752
rect 447 1718 480 1752
rect 380 1684 480 1718
rect 380 1650 413 1684
rect 447 1650 480 1684
rect 380 1616 480 1650
rect 380 1582 413 1616
rect 447 1582 480 1616
rect 380 1548 480 1582
rect 380 1514 413 1548
rect 447 1514 480 1548
rect 380 1480 480 1514
rect 380 1446 413 1480
rect 447 1446 480 1480
rect 380 1412 480 1446
rect 380 1378 413 1412
rect 447 1378 480 1412
rect 380 1344 480 1378
rect 380 1310 413 1344
rect 447 1310 480 1344
rect 380 1276 480 1310
rect 380 1242 413 1276
rect 447 1242 480 1276
rect 380 1208 480 1242
rect 380 1174 413 1208
rect 447 1174 480 1208
rect 380 1140 480 1174
rect 380 1106 413 1140
rect 447 1106 480 1140
rect 380 1072 480 1106
rect 380 1038 413 1072
rect 447 1038 480 1072
rect 380 1004 480 1038
rect 380 970 413 1004
rect 447 970 480 1004
rect 380 936 480 970
rect 380 902 413 936
rect 447 902 480 936
rect 380 868 480 902
rect 380 834 413 868
rect 447 834 480 868
rect 380 800 480 834
rect 380 766 413 800
rect 447 766 480 800
rect 380 732 480 766
rect 380 698 413 732
rect 447 698 480 732
rect 380 664 480 698
rect 380 630 413 664
rect 447 630 480 664
rect 380 596 480 630
rect 380 562 413 596
rect 447 562 480 596
rect 380 528 480 562
rect 380 494 413 528
rect 447 494 480 528
rect 380 460 480 494
rect 380 426 413 460
rect 447 426 480 460
rect 380 392 480 426
rect 380 358 413 392
rect 447 358 480 392
rect 380 324 480 358
rect 380 290 413 324
rect 447 290 480 324
rect 380 256 480 290
rect 380 222 413 256
rect 447 222 480 256
rect 380 188 480 222
rect 380 154 413 188
rect 447 154 480 188
rect 380 120 480 154
rect 380 86 413 120
rect 447 86 480 120
rect 380 52 480 86
rect 380 18 413 52
rect 447 18 480 52
rect 380 -16 480 18
rect 380 -50 413 -16
rect 447 -50 480 -16
rect 380 -84 480 -50
rect 380 -118 413 -84
rect 447 -118 480 -84
rect 380 -152 480 -118
rect 380 -186 413 -152
rect 447 -186 480 -152
rect 380 -220 480 -186
rect 380 -254 413 -220
rect 447 -254 480 -220
rect 380 -288 480 -254
rect 380 -322 413 -288
rect 447 -322 480 -288
rect 380 -356 480 -322
rect 380 -390 413 -356
rect 447 -390 480 -356
rect 380 -460 480 -390
rect 2684 1820 2784 1890
rect 2684 1786 2717 1820
rect 2751 1786 2784 1820
rect 2684 1752 2784 1786
rect 2684 1718 2717 1752
rect 2751 1718 2784 1752
rect 2684 1684 2784 1718
rect 2684 1650 2717 1684
rect 2751 1650 2784 1684
rect 2684 1616 2784 1650
rect 2684 1582 2717 1616
rect 2751 1582 2784 1616
rect 2684 1548 2784 1582
rect 2684 1514 2717 1548
rect 2751 1514 2784 1548
rect 2684 1480 2784 1514
rect 2684 1446 2717 1480
rect 2751 1446 2784 1480
rect 2684 1412 2784 1446
rect 2684 1378 2717 1412
rect 2751 1378 2784 1412
rect 2684 1344 2784 1378
rect 2684 1310 2717 1344
rect 2751 1310 2784 1344
rect 2684 1276 2784 1310
rect 2684 1242 2717 1276
rect 2751 1242 2784 1276
rect 2684 1208 2784 1242
rect 2684 1174 2717 1208
rect 2751 1174 2784 1208
rect 2684 1140 2784 1174
rect 2684 1106 2717 1140
rect 2751 1106 2784 1140
rect 2684 1072 2784 1106
rect 2684 1038 2717 1072
rect 2751 1038 2784 1072
rect 2684 1004 2784 1038
rect 2684 970 2717 1004
rect 2751 970 2784 1004
rect 2684 936 2784 970
rect 2684 902 2717 936
rect 2751 902 2784 936
rect 2684 868 2784 902
rect 2684 834 2717 868
rect 2751 834 2784 868
rect 2684 800 2784 834
rect 2684 766 2717 800
rect 2751 766 2784 800
rect 2684 732 2784 766
rect 2684 698 2717 732
rect 2751 698 2784 732
rect 2684 664 2784 698
rect 2684 630 2717 664
rect 2751 630 2784 664
rect 2684 596 2784 630
rect 2684 562 2717 596
rect 2751 562 2784 596
rect 2684 528 2784 562
rect 2684 494 2717 528
rect 2751 494 2784 528
rect 2684 460 2784 494
rect 2684 426 2717 460
rect 2751 426 2784 460
rect 2684 392 2784 426
rect 2684 358 2717 392
rect 2751 358 2784 392
rect 2684 324 2784 358
rect 2684 290 2717 324
rect 2751 290 2784 324
rect 2684 256 2784 290
rect 2684 222 2717 256
rect 2751 222 2784 256
rect 2684 188 2784 222
rect 2684 154 2717 188
rect 2751 154 2784 188
rect 2684 120 2784 154
rect 2684 86 2717 120
rect 2751 86 2784 120
rect 2684 52 2784 86
rect 2684 18 2717 52
rect 2751 18 2784 52
rect 2684 -16 2784 18
rect 2684 -50 2717 -16
rect 2751 -50 2784 -16
rect 2684 -84 2784 -50
rect 2684 -118 2717 -84
rect 2751 -118 2784 -84
rect 2684 -152 2784 -118
rect 2684 -186 2717 -152
rect 2751 -186 2784 -152
rect 2684 -220 2784 -186
rect 2684 -254 2717 -220
rect 2751 -254 2784 -220
rect 2684 -288 2784 -254
rect 2684 -322 2717 -288
rect 2751 -322 2784 -288
rect 2684 -356 2784 -322
rect 2684 -390 2717 -356
rect 2751 -390 2784 -356
rect 2684 -460 2784 -390
rect 380 -493 2784 -460
rect 380 -527 545 -493
rect 579 -527 613 -493
rect 647 -527 681 -493
rect 715 -527 749 -493
rect 783 -527 817 -493
rect 851 -527 885 -493
rect 919 -527 953 -493
rect 987 -527 1021 -493
rect 1055 -527 1089 -493
rect 1123 -527 1157 -493
rect 1191 -527 1225 -493
rect 1259 -527 1293 -493
rect 1327 -527 1361 -493
rect 1395 -527 1429 -493
rect 1463 -527 1497 -493
rect 1531 -527 1565 -493
rect 1599 -527 1633 -493
rect 1667 -527 1701 -493
rect 1735 -527 1769 -493
rect 1803 -527 1837 -493
rect 1871 -527 1905 -493
rect 1939 -527 1973 -493
rect 2007 -527 2041 -493
rect 2075 -527 2109 -493
rect 2143 -527 2177 -493
rect 2211 -527 2245 -493
rect 2279 -527 2313 -493
rect 2347 -527 2381 -493
rect 2415 -527 2449 -493
rect 2483 -527 2517 -493
rect 2551 -527 2585 -493
rect 2619 -527 2784 -493
rect 380 -560 2784 -527
rect -58 -617 -25 -583
rect 9 -617 42 -583
rect -58 -651 42 -617
rect -58 -685 -25 -651
rect 9 -685 42 -651
rect -58 -719 42 -685
rect -58 -753 -25 -719
rect 9 -753 42 -719
rect -58 -787 42 -753
rect -58 -821 -25 -787
rect 9 -821 42 -787
rect -58 -855 42 -821
rect -58 -889 -25 -855
rect 9 -889 42 -855
rect -58 -923 42 -889
rect -58 -957 -25 -923
rect 9 -957 42 -923
rect -58 -991 42 -957
rect -58 -1025 -25 -991
rect 9 -1025 42 -991
rect -58 -1059 42 -1025
rect -58 -1093 -25 -1059
rect 9 -1093 42 -1059
rect -58 -1127 42 -1093
rect -58 -1161 -25 -1127
rect 9 -1161 42 -1127
rect -58 -1254 42 -1161
rect -3322 -1287 42 -1254
rect -3322 -1321 -3153 -1287
rect -3119 -1321 -3085 -1287
rect -3051 -1321 -3017 -1287
rect -2983 -1321 -2949 -1287
rect -2915 -1321 -2881 -1287
rect -2847 -1321 -2813 -1287
rect -2779 -1321 -2745 -1287
rect -2711 -1321 -2677 -1287
rect -2643 -1321 -2609 -1287
rect -2575 -1321 -2541 -1287
rect -2507 -1321 -2473 -1287
rect -2439 -1321 -2405 -1287
rect -2371 -1321 -2337 -1287
rect -2303 -1321 -2269 -1287
rect -2235 -1321 -2201 -1287
rect -2167 -1321 -2133 -1287
rect -2099 -1321 -2065 -1287
rect -2031 -1321 -1997 -1287
rect -1963 -1321 -1929 -1287
rect -1895 -1321 -1861 -1287
rect -1827 -1321 -1793 -1287
rect -1759 -1321 -1725 -1287
rect -1691 -1321 -1657 -1287
rect -1623 -1321 -1589 -1287
rect -1555 -1321 -1521 -1287
rect -1487 -1321 -1453 -1287
rect -1419 -1321 -1385 -1287
rect -1351 -1321 -1317 -1287
rect -1283 -1321 -1249 -1287
rect -1215 -1321 -1181 -1287
rect -1147 -1321 -1113 -1287
rect -1079 -1321 -1045 -1287
rect -1011 -1321 -977 -1287
rect -943 -1321 -909 -1287
rect -875 -1321 -841 -1287
rect -807 -1321 -773 -1287
rect -739 -1321 -705 -1287
rect -671 -1321 -637 -1287
rect -603 -1321 -569 -1287
rect -535 -1321 -501 -1287
rect -467 -1321 -433 -1287
rect -399 -1321 -365 -1287
rect -331 -1321 -297 -1287
rect -263 -1321 -229 -1287
rect -195 -1321 -161 -1287
rect -127 -1321 42 -1287
rect -3322 -1354 42 -1321
rect -1365 -1415 -7 -1414
rect -1365 -1448 40 -1415
rect -1365 -1449 -1340 -1448
rect -1344 -1450 -1340 -1449
rect 6 -1489 40 -1448
<< psubdiffcont >>
rect 1087 -1443 1121 -1409
rect 1155 -1443 1189 -1409
rect 1223 -1443 1257 -1409
rect 1291 -1443 1325 -1409
rect 1359 -1443 1393 -1409
rect 1427 -1443 1461 -1409
rect 1495 -1443 1529 -1409
rect 1563 -1443 1597 -1409
rect 1631 -1443 1665 -1409
rect 1699 -1443 1733 -1409
rect 1767 -1443 1801 -1409
rect 1835 -1443 1869 -1409
rect 1903 -1443 1937 -1409
rect 1971 -1443 2005 -1409
rect 925 -1598 959 -1564
rect 925 -1666 959 -1632
rect 2183 -1602 2217 -1568
rect 925 -1734 959 -1700
rect 925 -1802 959 -1768
rect 925 -1870 959 -1836
rect 2183 -1670 2217 -1636
rect 2183 -1738 2217 -1704
rect 2183 -1806 2217 -1772
rect 925 -1938 959 -1904
rect 2183 -1874 2217 -1840
rect 2183 -1942 2217 -1908
rect 925 -2006 959 -1972
rect 925 -2074 959 -2040
rect 2183 -2010 2217 -1976
rect 2183 -2078 2217 -2044
rect 2183 -2146 2217 -2112
rect 1081 -2701 1115 -2667
rect 1149 -2701 1183 -2667
rect 1217 -2701 1251 -2667
rect 1285 -2701 1319 -2667
rect 1353 -2701 1387 -2667
rect 1421 -2701 1455 -2667
rect 1489 -2701 1523 -2667
rect 1557 -2701 1591 -2667
rect 1625 -2701 1659 -2667
rect 1693 -2701 1727 -2667
rect 1761 -2701 1795 -2667
rect 1829 -2701 1863 -2667
rect 1897 -2701 1931 -2667
rect 1965 -2701 1999 -2667
<< nsubdiffcont >>
rect -3153 1923 -3119 1957
rect -3085 1923 -3051 1957
rect -3017 1923 -2983 1957
rect -2949 1923 -2915 1957
rect -2881 1923 -2847 1957
rect -2813 1923 -2779 1957
rect -2745 1923 -2711 1957
rect -2677 1923 -2643 1957
rect -2609 1923 -2575 1957
rect -2541 1923 -2507 1957
rect -2473 1923 -2439 1957
rect -2405 1923 -2371 1957
rect -2337 1923 -2303 1957
rect -2269 1923 -2235 1957
rect -2201 1923 -2167 1957
rect -2133 1923 -2099 1957
rect -2065 1923 -2031 1957
rect -1997 1923 -1963 1957
rect -1929 1923 -1895 1957
rect -1861 1923 -1827 1957
rect -1793 1923 -1759 1957
rect -1725 1923 -1691 1957
rect -1657 1923 -1623 1957
rect -1589 1923 -1555 1957
rect -1521 1923 -1487 1957
rect -1453 1923 -1419 1957
rect -1385 1923 -1351 1957
rect -1317 1923 -1283 1957
rect -1249 1923 -1215 1957
rect -1181 1923 -1147 1957
rect -1113 1923 -1079 1957
rect -1045 1923 -1011 1957
rect -977 1923 -943 1957
rect -909 1923 -875 1957
rect -841 1923 -807 1957
rect -773 1923 -739 1957
rect -705 1923 -671 1957
rect -637 1923 -603 1957
rect -569 1923 -535 1957
rect -501 1923 -467 1957
rect -433 1923 -399 1957
rect -365 1923 -331 1957
rect -297 1923 -263 1957
rect -229 1923 -195 1957
rect -161 1923 -127 1957
rect -3289 1763 -3255 1797
rect -3289 1695 -3255 1729
rect -3289 1627 -3255 1661
rect -3289 1559 -3255 1593
rect -3289 1491 -3255 1525
rect -3289 1423 -3255 1457
rect -3289 1355 -3255 1389
rect -3289 1287 -3255 1321
rect -3289 1219 -3255 1253
rect -3289 1151 -3255 1185
rect -3289 1083 -3255 1117
rect -3289 1015 -3255 1049
rect -3289 947 -3255 981
rect -3289 879 -3255 913
rect -3289 811 -3255 845
rect -3289 743 -3255 777
rect -3289 675 -3255 709
rect -3289 607 -3255 641
rect -3289 539 -3255 573
rect -3289 471 -3255 505
rect -3289 403 -3255 437
rect -3289 335 -3255 369
rect -3289 267 -3255 301
rect -3289 199 -3255 233
rect -3289 131 -3255 165
rect -3289 63 -3255 97
rect -3289 -5 -3255 29
rect -3289 -73 -3255 -39
rect -3289 -141 -3255 -107
rect -3289 -209 -3255 -175
rect -3289 -277 -3255 -243
rect -3289 -345 -3255 -311
rect -3289 -413 -3255 -379
rect -3289 -481 -3255 -447
rect -3289 -549 -3255 -515
rect -3289 -617 -3255 -583
rect -3289 -685 -3255 -651
rect -3289 -753 -3255 -719
rect -3289 -821 -3255 -787
rect -3289 -889 -3255 -855
rect -3289 -957 -3255 -923
rect -3289 -1025 -3255 -991
rect -3289 -1093 -3255 -1059
rect -3289 -1161 -3255 -1127
rect -25 1763 9 1797
rect -25 1695 9 1729
rect -25 1627 9 1661
rect -25 1559 9 1593
rect -25 1491 9 1525
rect -25 1423 9 1457
rect -25 1355 9 1389
rect -25 1287 9 1321
rect -25 1219 9 1253
rect -25 1151 9 1185
rect -25 1083 9 1117
rect -25 1015 9 1049
rect -25 947 9 981
rect -25 879 9 913
rect -25 811 9 845
rect -25 743 9 777
rect -25 675 9 709
rect -25 607 9 641
rect -25 539 9 573
rect -25 471 9 505
rect -25 403 9 437
rect -25 335 9 369
rect -25 267 9 301
rect -25 199 9 233
rect -25 131 9 165
rect -25 63 9 97
rect -25 -5 9 29
rect -25 -73 9 -39
rect -25 -141 9 -107
rect -25 -209 9 -175
rect -25 -277 9 -243
rect -25 -345 9 -311
rect -25 -413 9 -379
rect -25 -481 9 -447
rect -25 -549 9 -515
rect 545 1923 579 1957
rect 613 1923 647 1957
rect 681 1923 715 1957
rect 749 1923 783 1957
rect 817 1923 851 1957
rect 885 1923 919 1957
rect 953 1923 987 1957
rect 1021 1923 1055 1957
rect 1089 1923 1123 1957
rect 1157 1923 1191 1957
rect 1225 1923 1259 1957
rect 1293 1923 1327 1957
rect 1361 1923 1395 1957
rect 1429 1923 1463 1957
rect 1497 1923 1531 1957
rect 1565 1923 1599 1957
rect 1633 1923 1667 1957
rect 1701 1923 1735 1957
rect 1769 1923 1803 1957
rect 1837 1923 1871 1957
rect 1905 1923 1939 1957
rect 1973 1923 2007 1957
rect 2041 1923 2075 1957
rect 2109 1923 2143 1957
rect 2177 1923 2211 1957
rect 2245 1923 2279 1957
rect 2313 1923 2347 1957
rect 2381 1923 2415 1957
rect 2449 1923 2483 1957
rect 2517 1923 2551 1957
rect 2585 1923 2619 1957
rect 413 1786 447 1820
rect 413 1718 447 1752
rect 413 1650 447 1684
rect 413 1582 447 1616
rect 413 1514 447 1548
rect 413 1446 447 1480
rect 413 1378 447 1412
rect 413 1310 447 1344
rect 413 1242 447 1276
rect 413 1174 447 1208
rect 413 1106 447 1140
rect 413 1038 447 1072
rect 413 970 447 1004
rect 413 902 447 936
rect 413 834 447 868
rect 413 766 447 800
rect 413 698 447 732
rect 413 630 447 664
rect 413 562 447 596
rect 413 494 447 528
rect 413 426 447 460
rect 413 358 447 392
rect 413 290 447 324
rect 413 222 447 256
rect 413 154 447 188
rect 413 86 447 120
rect 413 18 447 52
rect 413 -50 447 -16
rect 413 -118 447 -84
rect 413 -186 447 -152
rect 413 -254 447 -220
rect 413 -322 447 -288
rect 413 -390 447 -356
rect 2717 1786 2751 1820
rect 2717 1718 2751 1752
rect 2717 1650 2751 1684
rect 2717 1582 2751 1616
rect 2717 1514 2751 1548
rect 2717 1446 2751 1480
rect 2717 1378 2751 1412
rect 2717 1310 2751 1344
rect 2717 1242 2751 1276
rect 2717 1174 2751 1208
rect 2717 1106 2751 1140
rect 2717 1038 2751 1072
rect 2717 970 2751 1004
rect 2717 902 2751 936
rect 2717 834 2751 868
rect 2717 766 2751 800
rect 2717 698 2751 732
rect 2717 630 2751 664
rect 2717 562 2751 596
rect 2717 494 2751 528
rect 2717 426 2751 460
rect 2717 358 2751 392
rect 2717 290 2751 324
rect 2717 222 2751 256
rect 2717 154 2751 188
rect 2717 86 2751 120
rect 2717 18 2751 52
rect 2717 -50 2751 -16
rect 2717 -118 2751 -84
rect 2717 -186 2751 -152
rect 2717 -254 2751 -220
rect 2717 -322 2751 -288
rect 2717 -390 2751 -356
rect 545 -527 579 -493
rect 613 -527 647 -493
rect 681 -527 715 -493
rect 749 -527 783 -493
rect 817 -527 851 -493
rect 885 -527 919 -493
rect 953 -527 987 -493
rect 1021 -527 1055 -493
rect 1089 -527 1123 -493
rect 1157 -527 1191 -493
rect 1225 -527 1259 -493
rect 1293 -527 1327 -493
rect 1361 -527 1395 -493
rect 1429 -527 1463 -493
rect 1497 -527 1531 -493
rect 1565 -527 1599 -493
rect 1633 -527 1667 -493
rect 1701 -527 1735 -493
rect 1769 -527 1803 -493
rect 1837 -527 1871 -493
rect 1905 -527 1939 -493
rect 1973 -527 2007 -493
rect 2041 -527 2075 -493
rect 2109 -527 2143 -493
rect 2177 -527 2211 -493
rect 2245 -527 2279 -493
rect 2313 -527 2347 -493
rect 2381 -527 2415 -493
rect 2449 -527 2483 -493
rect 2517 -527 2551 -493
rect 2585 -527 2619 -493
rect -25 -617 9 -583
rect -25 -685 9 -651
rect -25 -753 9 -719
rect -25 -821 9 -787
rect -25 -889 9 -855
rect -25 -957 9 -923
rect -25 -1025 9 -991
rect -25 -1093 9 -1059
rect -25 -1161 9 -1127
rect -3153 -1321 -3119 -1287
rect -3085 -1321 -3051 -1287
rect -3017 -1321 -2983 -1287
rect -2949 -1321 -2915 -1287
rect -2881 -1321 -2847 -1287
rect -2813 -1321 -2779 -1287
rect -2745 -1321 -2711 -1287
rect -2677 -1321 -2643 -1287
rect -2609 -1321 -2575 -1287
rect -2541 -1321 -2507 -1287
rect -2473 -1321 -2439 -1287
rect -2405 -1321 -2371 -1287
rect -2337 -1321 -2303 -1287
rect -2269 -1321 -2235 -1287
rect -2201 -1321 -2167 -1287
rect -2133 -1321 -2099 -1287
rect -2065 -1321 -2031 -1287
rect -1997 -1321 -1963 -1287
rect -1929 -1321 -1895 -1287
rect -1861 -1321 -1827 -1287
rect -1793 -1321 -1759 -1287
rect -1725 -1321 -1691 -1287
rect -1657 -1321 -1623 -1287
rect -1589 -1321 -1555 -1287
rect -1521 -1321 -1487 -1287
rect -1453 -1321 -1419 -1287
rect -1385 -1321 -1351 -1287
rect -1317 -1321 -1283 -1287
rect -1249 -1321 -1215 -1287
rect -1181 -1321 -1147 -1287
rect -1113 -1321 -1079 -1287
rect -1045 -1321 -1011 -1287
rect -977 -1321 -943 -1287
rect -909 -1321 -875 -1287
rect -841 -1321 -807 -1287
rect -773 -1321 -739 -1287
rect -705 -1321 -671 -1287
rect -637 -1321 -603 -1287
rect -569 -1321 -535 -1287
rect -501 -1321 -467 -1287
rect -433 -1321 -399 -1287
rect -365 -1321 -331 -1287
rect -297 -1321 -263 -1287
rect -229 -1321 -195 -1287
rect -161 -1321 -127 -1287
<< poly >>
rect -1092 -1525 -1010 -1507
rect -1092 -1559 -1068 -1525
rect -1034 -1559 -1010 -1525
rect -1092 -1577 -1010 -1559
rect -964 -1525 -882 -1507
rect -964 -1559 -940 -1525
rect -906 -1559 -882 -1525
rect -964 -1577 -882 -1559
rect -836 -1525 -754 -1507
rect -836 -1559 -812 -1525
rect -778 -1559 -754 -1525
rect -836 -1577 -754 -1559
rect -708 -1525 -626 -1507
rect -708 -1559 -684 -1525
rect -650 -1559 -626 -1525
rect -708 -1577 -626 -1559
rect -580 -1525 -498 -1507
rect -580 -1559 -556 -1525
rect -522 -1559 -498 -1525
rect -580 -1577 -498 -1559
rect -452 -1525 -370 -1507
rect -452 -1559 -428 -1525
rect -394 -1559 -370 -1525
rect -452 -1577 -370 -1559
rect -324 -1525 -242 -1507
rect -324 -1559 -300 -1525
rect -266 -1559 -242 -1525
rect -324 -1577 -242 -1559
rect -1086 -1624 -1016 -1577
rect -958 -1624 -888 -1577
rect -830 -1624 -760 -1577
rect -702 -1622 -632 -1577
rect -574 -1623 -504 -1577
rect -446 -1623 -376 -1577
rect -318 -1623 -248 -1577
rect 1248 -1545 1308 -1526
rect 1248 -1579 1261 -1545
rect 1295 -1579 1308 -1545
rect 1248 -1644 1308 -1579
rect 1478 -1545 1550 -1532
rect 1478 -1579 1497 -1545
rect 1531 -1579 1550 -1545
rect 1478 -1592 1550 -1579
rect 1596 -1545 1668 -1532
rect 1596 -1579 1615 -1545
rect 1649 -1579 1668 -1545
rect 1596 -1592 1668 -1579
rect 1832 -1545 1904 -1532
rect 1832 -1579 1851 -1545
rect 1885 -1579 1904 -1545
rect 1832 -1592 1904 -1579
rect 1484 -1646 1544 -1592
rect 1602 -1646 1662 -1592
rect 1838 -1644 1898 -1592
rect -1214 -1869 -1144 -1824
rect -190 -1869 -120 -1826
rect -1220 -1887 -1138 -1869
rect -1220 -1921 -1196 -1887
rect -1162 -1921 -1138 -1887
rect -1220 -1939 -1138 -1921
rect -196 -1887 -114 -1869
rect -196 -1921 -172 -1887
rect -138 -1921 -114 -1887
rect -196 -1939 -114 -1921
rect 1130 -1896 1190 -1848
rect 1064 -1909 1190 -1896
rect 1366 -1898 1426 -1846
rect 1720 -1898 1780 -1846
rect 1956 -1896 2016 -1848
rect 1064 -1943 1083 -1909
rect 1117 -1943 1190 -1909
rect 1064 -1956 1190 -1943
rect 1360 -1911 1432 -1898
rect 1360 -1945 1379 -1911
rect 1413 -1945 1432 -1911
rect 1360 -1958 1432 -1945
rect 1714 -1911 1786 -1898
rect 1714 -1945 1733 -1911
rect 1767 -1945 1786 -1911
rect 1714 -1958 1786 -1945
rect 1956 -1909 2084 -1896
rect 1956 -1943 2031 -1909
rect 2065 -1943 2084 -1909
rect 1956 -1956 2084 -1943
<< polycont >>
rect -1068 -1559 -1034 -1525
rect -940 -1559 -906 -1525
rect -812 -1559 -778 -1525
rect -684 -1559 -650 -1525
rect -556 -1559 -522 -1525
rect -428 -1559 -394 -1525
rect -300 -1559 -266 -1525
rect 1261 -1579 1295 -1545
rect 1497 -1579 1531 -1545
rect 1615 -1579 1649 -1545
rect 1851 -1579 1885 -1545
rect -1196 -1921 -1162 -1887
rect -172 -1921 -138 -1887
rect 1083 -1943 1117 -1909
rect 1379 -1945 1413 -1911
rect 1733 -1945 1767 -1911
rect 2031 -1943 2065 -1909
<< locali >>
rect -3322 1957 42 1990
rect -3322 1923 -3205 1957
rect -3171 1923 -3153 1957
rect -3099 1923 -3085 1957
rect -3027 1923 -3017 1957
rect -2955 1923 -2949 1957
rect -2883 1923 -2881 1957
rect -2847 1923 -2845 1957
rect -2779 1923 -2773 1957
rect -2711 1923 -2701 1957
rect -2643 1923 -2629 1957
rect -2575 1923 -2557 1957
rect -2507 1923 -2485 1957
rect -2439 1923 -2413 1957
rect -2371 1923 -2341 1957
rect -2303 1923 -2269 1957
rect -2235 1923 -2201 1957
rect -2163 1923 -2133 1957
rect -2091 1923 -2065 1957
rect -2019 1923 -1997 1957
rect -1947 1923 -1929 1957
rect -1875 1923 -1861 1957
rect -1803 1923 -1793 1957
rect -1731 1923 -1725 1957
rect -1659 1923 -1657 1957
rect -1623 1923 -1621 1957
rect -1555 1923 -1549 1957
rect -1487 1923 -1477 1957
rect -1419 1923 -1405 1957
rect -1351 1923 -1333 1957
rect -1283 1923 -1261 1957
rect -1215 1923 -1189 1957
rect -1147 1923 -1117 1957
rect -1079 1923 -1045 1957
rect -1011 1923 -977 1957
rect -939 1923 -909 1957
rect -867 1923 -841 1957
rect -795 1923 -773 1957
rect -723 1923 -705 1957
rect -651 1923 -637 1957
rect -579 1923 -569 1957
rect -507 1923 -501 1957
rect -435 1923 -433 1957
rect -399 1923 -397 1957
rect -331 1923 -325 1957
rect -263 1923 -253 1957
rect -195 1923 -181 1957
rect -127 1923 -109 1957
rect -75 1923 42 1957
rect -3322 1890 42 1923
rect -3322 1797 -3222 1890
rect -3322 1763 -3289 1797
rect -3255 1763 -3222 1797
rect -3322 1739 -3222 1763
rect -3322 1695 -3289 1739
rect -3255 1695 -3222 1739
rect -3322 1667 -3222 1695
rect -3322 1627 -3289 1667
rect -3255 1627 -3222 1667
rect -3322 1595 -3222 1627
rect -3322 1559 -3289 1595
rect -3255 1559 -3222 1595
rect -3322 1525 -3222 1559
rect -3322 1489 -3289 1525
rect -3255 1489 -3222 1525
rect -3322 1457 -3222 1489
rect -3322 1417 -3289 1457
rect -3255 1417 -3222 1457
rect -3322 1389 -3222 1417
rect -3322 1345 -3289 1389
rect -3255 1345 -3222 1389
rect -3322 1321 -3222 1345
rect -3322 1273 -3289 1321
rect -3255 1273 -3222 1321
rect -3322 1253 -3222 1273
rect -3322 1201 -3289 1253
rect -3255 1201 -3222 1253
rect -3322 1185 -3222 1201
rect -3322 1129 -3289 1185
rect -3255 1129 -3222 1185
rect -3322 1117 -3222 1129
rect -3322 1057 -3289 1117
rect -3255 1057 -3222 1117
rect -3322 1049 -3222 1057
rect -3322 985 -3289 1049
rect -3255 985 -3222 1049
rect -3322 981 -3222 985
rect -3322 879 -3289 981
rect -3255 879 -3222 981
rect -3322 875 -3222 879
rect -3322 811 -3289 875
rect -3255 811 -3222 875
rect -3322 803 -3222 811
rect -3322 743 -3289 803
rect -3255 743 -3222 803
rect -3322 731 -3222 743
rect -3322 675 -3289 731
rect -3255 675 -3222 731
rect -3322 659 -3222 675
rect -3322 607 -3289 659
rect -3255 607 -3222 659
rect -3322 587 -3222 607
rect -3322 539 -3289 587
rect -3255 539 -3222 587
rect -3322 515 -3222 539
rect -3322 471 -3289 515
rect -3255 471 -3222 515
rect -3322 443 -3222 471
rect -3322 403 -3289 443
rect -3255 403 -3222 443
rect -3322 371 -3222 403
rect -3322 335 -3289 371
rect -3255 335 -3222 371
rect -3322 301 -3222 335
rect -3322 265 -3289 301
rect -3255 265 -3222 301
rect -3322 233 -3222 265
rect -3322 193 -3289 233
rect -3255 193 -3222 233
rect -3322 165 -3222 193
rect -3322 121 -3289 165
rect -3255 121 -3222 165
rect -3322 97 -3222 121
rect -3322 49 -3289 97
rect -3255 49 -3222 97
rect -3322 29 -3222 49
rect -3322 -23 -3289 29
rect -3255 -23 -3222 29
rect -3322 -39 -3222 -23
rect -3322 -95 -3289 -39
rect -3255 -95 -3222 -39
rect -3322 -107 -3222 -95
rect -3322 -167 -3289 -107
rect -3255 -167 -3222 -107
rect -3322 -175 -3222 -167
rect -3322 -239 -3289 -175
rect -3255 -239 -3222 -175
rect -3322 -243 -3222 -239
rect -3322 -345 -3289 -243
rect -3255 -345 -3222 -243
rect -3322 -349 -3222 -345
rect -3322 -413 -3289 -349
rect -3255 -413 -3222 -349
rect -3322 -421 -3222 -413
rect -3322 -481 -3289 -421
rect -3255 -481 -3222 -421
rect -3322 -493 -3222 -481
rect -3322 -549 -3289 -493
rect -3255 -549 -3222 -493
rect -3322 -565 -3222 -549
rect -3322 -617 -3289 -565
rect -3255 -617 -3222 -565
rect -3322 -637 -3222 -617
rect -3322 -685 -3289 -637
rect -3255 -685 -3222 -637
rect -3322 -709 -3222 -685
rect -3322 -753 -3289 -709
rect -3255 -753 -3222 -709
rect -3322 -781 -3222 -753
rect -3322 -821 -3289 -781
rect -3255 -821 -3222 -781
rect -3322 -853 -3222 -821
rect -3322 -889 -3289 -853
rect -3255 -889 -3222 -853
rect -3322 -923 -3222 -889
rect -3322 -959 -3289 -923
rect -3255 -959 -3222 -923
rect -3322 -991 -3222 -959
rect -3322 -1031 -3289 -991
rect -3255 -1031 -3222 -991
rect -3322 -1059 -3222 -1031
rect -3322 -1103 -3289 -1059
rect -3255 -1103 -3222 -1059
rect -3322 -1127 -3222 -1103
rect -3322 -1161 -3289 -1127
rect -3255 -1161 -3222 -1127
rect -3322 -1254 -3222 -1161
rect -58 1797 42 1890
rect -58 1763 -25 1797
rect 9 1763 42 1797
rect -58 1739 42 1763
rect -58 1695 -25 1739
rect 9 1695 42 1739
rect -58 1667 42 1695
rect -58 1627 -25 1667
rect 9 1627 42 1667
rect -58 1595 42 1627
rect -58 1559 -25 1595
rect 9 1559 42 1595
rect -58 1525 42 1559
rect -58 1489 -25 1525
rect 9 1489 42 1525
rect -58 1457 42 1489
rect -58 1417 -25 1457
rect 9 1417 42 1457
rect -58 1389 42 1417
rect -58 1345 -25 1389
rect 9 1345 42 1389
rect -58 1321 42 1345
rect -58 1273 -25 1321
rect 9 1273 42 1321
rect -58 1253 42 1273
rect -58 1201 -25 1253
rect 9 1201 42 1253
rect -58 1185 42 1201
rect -58 1129 -25 1185
rect 9 1129 42 1185
rect -58 1117 42 1129
rect -58 1057 -25 1117
rect 9 1057 42 1117
rect -58 1049 42 1057
rect -58 985 -25 1049
rect 9 985 42 1049
rect -58 981 42 985
rect -58 879 -25 981
rect 9 879 42 981
rect -58 875 42 879
rect -58 811 -25 875
rect 9 811 42 875
rect -58 803 42 811
rect -58 743 -25 803
rect 9 743 42 803
rect -58 731 42 743
rect -58 675 -25 731
rect 9 675 42 731
rect -58 659 42 675
rect -58 607 -25 659
rect 9 607 42 659
rect -58 587 42 607
rect -58 539 -25 587
rect 9 539 42 587
rect -58 515 42 539
rect -58 471 -25 515
rect 9 471 42 515
rect -58 443 42 471
rect -58 403 -25 443
rect 9 403 42 443
rect -58 371 42 403
rect -58 335 -25 371
rect 9 335 42 371
rect -58 301 42 335
rect -58 265 -25 301
rect 9 265 42 301
rect -58 233 42 265
rect -58 193 -25 233
rect 9 193 42 233
rect -58 165 42 193
rect -58 121 -25 165
rect 9 121 42 165
rect -58 97 42 121
rect -58 49 -25 97
rect 9 49 42 97
rect -58 29 42 49
rect -58 -23 -25 29
rect 9 -23 42 29
rect -58 -39 42 -23
rect -58 -95 -25 -39
rect 9 -95 42 -39
rect -58 -107 42 -95
rect -58 -167 -25 -107
rect 9 -167 42 -107
rect -58 -175 42 -167
rect -58 -239 -25 -175
rect 9 -239 42 -175
rect -58 -243 42 -239
rect -58 -345 -25 -243
rect 9 -345 42 -243
rect -58 -349 42 -345
rect -58 -413 -25 -349
rect 9 -413 42 -349
rect -58 -421 42 -413
rect -58 -481 -25 -421
rect 9 -481 42 -421
rect -58 -493 42 -481
rect -58 -549 -25 -493
rect 9 -549 42 -493
rect -58 -565 42 -549
rect 380 1957 2784 1990
rect 380 1923 485 1957
rect 519 1923 545 1957
rect 591 1923 613 1957
rect 663 1923 681 1957
rect 735 1923 749 1957
rect 807 1923 817 1957
rect 879 1923 885 1957
rect 951 1923 953 1957
rect 987 1923 989 1957
rect 1055 1923 1061 1957
rect 1123 1923 1133 1957
rect 1191 1923 1205 1957
rect 1259 1923 1277 1957
rect 1327 1923 1349 1957
rect 1395 1923 1421 1957
rect 1463 1923 1493 1957
rect 1531 1923 1565 1957
rect 1599 1923 1633 1957
rect 1671 1923 1701 1957
rect 1743 1923 1769 1957
rect 1815 1923 1837 1957
rect 1887 1923 1905 1957
rect 1959 1923 1973 1957
rect 2031 1923 2041 1957
rect 2103 1923 2109 1957
rect 2175 1923 2177 1957
rect 2211 1923 2213 1957
rect 2279 1923 2285 1957
rect 2347 1923 2357 1957
rect 2415 1923 2429 1957
rect 2483 1923 2501 1957
rect 2551 1923 2573 1957
rect 2619 1923 2645 1957
rect 2679 1923 2784 1957
rect 380 1890 2784 1923
rect 380 1820 480 1890
rect 380 1786 413 1820
rect 447 1786 480 1820
rect 380 1776 480 1786
rect 380 1718 413 1776
rect 447 1718 480 1776
rect 380 1704 480 1718
rect 380 1650 413 1704
rect 447 1650 480 1704
rect 380 1632 480 1650
rect 380 1582 413 1632
rect 447 1582 480 1632
rect 380 1560 480 1582
rect 380 1514 413 1560
rect 447 1514 480 1560
rect 380 1488 480 1514
rect 380 1446 413 1488
rect 447 1446 480 1488
rect 380 1416 480 1446
rect 380 1378 413 1416
rect 447 1378 480 1416
rect 380 1344 480 1378
rect 380 1310 413 1344
rect 447 1310 480 1344
rect 380 1276 480 1310
rect 380 1238 413 1276
rect 447 1238 480 1276
rect 380 1208 480 1238
rect 380 1166 413 1208
rect 447 1166 480 1208
rect 380 1140 480 1166
rect 380 1094 413 1140
rect 447 1094 480 1140
rect 380 1072 480 1094
rect 380 1022 413 1072
rect 447 1022 480 1072
rect 380 1004 480 1022
rect 380 950 413 1004
rect 447 950 480 1004
rect 380 936 480 950
rect 380 878 413 936
rect 447 878 480 936
rect 380 868 480 878
rect 380 806 413 868
rect 447 806 480 868
rect 380 800 480 806
rect 380 734 413 800
rect 447 734 480 800
rect 380 732 480 734
rect 380 698 413 732
rect 447 698 480 732
rect 380 696 480 698
rect 380 630 413 696
rect 447 630 480 696
rect 380 624 480 630
rect 380 562 413 624
rect 447 562 480 624
rect 380 552 480 562
rect 380 494 413 552
rect 447 494 480 552
rect 380 480 480 494
rect 380 426 413 480
rect 447 426 480 480
rect 380 408 480 426
rect 380 358 413 408
rect 447 358 480 408
rect 380 336 480 358
rect 380 290 413 336
rect 447 290 480 336
rect 380 264 480 290
rect 380 222 413 264
rect 447 222 480 264
rect 380 192 480 222
rect 380 154 413 192
rect 447 154 480 192
rect 380 120 480 154
rect 380 86 413 120
rect 447 86 480 120
rect 380 52 480 86
rect 380 14 413 52
rect 447 14 480 52
rect 380 -16 480 14
rect 380 -58 413 -16
rect 447 -58 480 -16
rect 380 -84 480 -58
rect 380 -130 413 -84
rect 447 -130 480 -84
rect 380 -152 480 -130
rect 380 -202 413 -152
rect 447 -202 480 -152
rect 380 -220 480 -202
rect 380 -274 413 -220
rect 447 -274 480 -220
rect 380 -288 480 -274
rect 380 -346 413 -288
rect 447 -346 480 -288
rect 380 -356 480 -346
rect 380 -390 413 -356
rect 447 -390 480 -356
rect 380 -460 480 -390
rect 2684 1820 2784 1890
rect 2684 1786 2717 1820
rect 2751 1789 2784 1820
rect 2684 1755 2719 1786
rect 2753 1755 2784 1789
rect 2684 1752 2784 1755
rect 2684 1718 2717 1752
rect 2751 1718 2784 1752
rect 2684 1717 2784 1718
rect 2684 1684 2719 1717
rect 2684 1650 2717 1684
rect 2753 1683 2784 1717
rect 2751 1650 2784 1683
rect 2684 1645 2784 1650
rect 2684 1616 2719 1645
rect 2684 1582 2717 1616
rect 2753 1611 2784 1645
rect 2751 1582 2784 1611
rect 2684 1548 2784 1582
rect 2684 1514 2717 1548
rect 2751 1514 2784 1548
rect 2684 1496 2784 1514
rect 2684 1446 2717 1496
rect 2751 1446 2784 1496
rect 2684 1424 2784 1446
rect 2684 1378 2717 1424
rect 2751 1378 2784 1424
rect 2684 1352 2784 1378
rect 2684 1310 2717 1352
rect 2751 1310 2784 1352
rect 2684 1280 2784 1310
rect 2684 1242 2717 1280
rect 2751 1242 2784 1280
rect 2684 1208 2784 1242
rect 2684 1174 2717 1208
rect 2751 1174 2784 1208
rect 2684 1140 2784 1174
rect 2684 1102 2717 1140
rect 2751 1102 2784 1140
rect 2684 1072 2784 1102
rect 2684 1030 2717 1072
rect 2751 1030 2784 1072
rect 2684 1004 2784 1030
rect 2684 958 2717 1004
rect 2751 958 2784 1004
rect 2684 936 2784 958
rect 2684 886 2717 936
rect 2751 886 2784 936
rect 2684 868 2784 886
rect 2684 814 2717 868
rect 2751 814 2784 868
rect 2684 800 2784 814
rect 2684 742 2717 800
rect 2751 742 2784 800
rect 2684 732 2784 742
rect 2684 670 2717 732
rect 2751 670 2784 732
rect 2684 664 2784 670
rect 2684 598 2717 664
rect 2751 598 2784 664
rect 2684 596 2784 598
rect 2684 562 2717 596
rect 2751 562 2784 596
rect 2684 560 2784 562
rect 2684 494 2717 560
rect 2751 494 2784 560
rect 2684 488 2784 494
rect 2684 426 2717 488
rect 2751 426 2784 488
rect 2684 416 2784 426
rect 2684 358 2717 416
rect 2751 358 2784 416
rect 2684 344 2784 358
rect 2684 290 2717 344
rect 2751 290 2784 344
rect 2684 272 2784 290
rect 2684 222 2717 272
rect 2751 222 2784 272
rect 2684 200 2784 222
rect 2684 154 2717 200
rect 2751 154 2784 200
rect 2684 128 2784 154
rect 2684 86 2717 128
rect 2751 86 2784 128
rect 2684 56 2784 86
rect 2684 18 2717 56
rect 2751 18 2784 56
rect 2684 -16 2784 18
rect 2684 -50 2717 -16
rect 2751 -50 2784 -16
rect 2684 -84 2784 -50
rect 2684 -122 2717 -84
rect 2751 -122 2784 -84
rect 2684 -152 2784 -122
rect 2684 -194 2717 -152
rect 2751 -194 2784 -152
rect 2684 -220 2784 -194
rect 2684 -266 2717 -220
rect 2751 -266 2784 -220
rect 2684 -288 2784 -266
rect 2684 -338 2717 -288
rect 2751 -338 2784 -288
rect 2684 -356 2784 -338
rect 2684 -390 2717 -356
rect 2751 -390 2784 -356
rect 2684 -460 2784 -390
rect 380 -493 2784 -460
rect 380 -527 485 -493
rect 519 -527 545 -493
rect 591 -527 613 -493
rect 663 -527 681 -493
rect 735 -527 749 -493
rect 807 -527 817 -493
rect 879 -527 885 -493
rect 951 -527 953 -493
rect 987 -527 989 -493
rect 1055 -527 1061 -493
rect 1123 -527 1133 -493
rect 1191 -527 1205 -493
rect 1259 -527 1277 -493
rect 1327 -527 1349 -493
rect 1395 -527 1421 -493
rect 1463 -527 1493 -493
rect 1531 -527 1565 -493
rect 1599 -527 1633 -493
rect 1671 -527 1701 -493
rect 1743 -527 1769 -493
rect 1815 -527 1837 -493
rect 1887 -527 1905 -493
rect 1959 -527 1973 -493
rect 2031 -527 2041 -493
rect 2103 -527 2109 -493
rect 2175 -527 2177 -493
rect 2211 -527 2213 -493
rect 2279 -527 2285 -493
rect 2347 -527 2357 -493
rect 2415 -527 2429 -493
rect 2483 -527 2501 -493
rect 2551 -527 2573 -493
rect 2619 -527 2645 -493
rect 2679 -527 2784 -493
rect 380 -560 2784 -527
rect -58 -617 -25 -565
rect 9 -617 42 -565
rect -58 -637 42 -617
rect -58 -685 -25 -637
rect 9 -685 42 -637
rect 1353 -638 1480 -605
rect 1514 -638 1572 -605
rect 1606 -638 1667 -605
rect 1353 -639 1667 -638
rect -58 -709 42 -685
rect -58 -753 -25 -709
rect 9 -753 42 -709
rect -58 -781 42 -753
rect -58 -821 -25 -781
rect 9 -821 42 -781
rect -58 -853 42 -821
rect -58 -889 -25 -853
rect 9 -889 42 -853
rect -58 -923 42 -889
rect -58 -959 -25 -923
rect 9 -959 42 -923
rect 692 -909 740 -902
rect 692 -943 699 -909
rect 733 -943 740 -909
rect 692 -950 740 -943
rect 804 -909 852 -902
rect 804 -943 811 -909
rect 845 -943 852 -909
rect 804 -950 852 -943
rect 964 -909 1012 -902
rect 964 -943 971 -909
rect 1005 -943 1012 -909
rect 964 -950 1012 -943
rect 1072 -909 1120 -902
rect 1072 -943 1079 -909
rect 1113 -943 1120 -909
rect 1072 -950 1120 -943
rect 1204 -909 1252 -902
rect 1204 -943 1211 -909
rect 1245 -943 1252 -909
rect 1204 -950 1252 -943
rect 1378 -909 1426 -902
rect 1378 -943 1385 -909
rect 1419 -943 1426 -909
rect 1852 -911 1900 -904
rect 1378 -950 1426 -943
rect 1852 -945 1859 -911
rect 1893 -945 1900 -911
rect 1852 -952 1900 -945
rect 1966 -911 2014 -904
rect 1966 -945 1973 -911
rect 2007 -945 2014 -911
rect 1966 -952 2014 -945
rect 2082 -909 2130 -902
rect 2082 -943 2089 -909
rect 2123 -943 2130 -909
rect 2082 -950 2130 -943
rect 2242 -909 2290 -902
rect 2242 -943 2249 -909
rect 2283 -943 2290 -909
rect 2242 -950 2290 -943
rect 2354 -909 2402 -902
rect 2354 -943 2361 -909
rect 2395 -943 2402 -909
rect 2354 -950 2402 -943
rect -58 -991 42 -959
rect -58 -1031 -25 -991
rect 9 -1031 42 -991
rect -58 -1059 42 -1031
rect -58 -1103 -25 -1059
rect 9 -1103 42 -1059
rect 1384 -1027 1432 -1020
rect 1384 -1061 1391 -1027
rect 1425 -1061 1432 -1027
rect 1384 -1068 1432 -1061
rect 1664 -1027 1712 -1020
rect 1664 -1061 1671 -1027
rect 1705 -1061 1712 -1027
rect 1664 -1068 1712 -1061
rect -58 -1127 42 -1103
rect -58 -1161 -25 -1127
rect 9 -1161 42 -1127
rect -58 -1254 42 -1161
rect 1357 -1150 1572 -1149
rect 1357 -1183 1480 -1150
rect 1514 -1182 1572 -1150
rect 1606 -1182 1715 -1149
rect 1514 -1183 1715 -1182
rect -3322 -1287 42 -1254
rect -3322 -1321 -3205 -1287
rect -3171 -1321 -3153 -1287
rect -3099 -1321 -3085 -1287
rect -3027 -1321 -3017 -1287
rect -2955 -1321 -2949 -1287
rect -2883 -1321 -2881 -1287
rect -2847 -1321 -2845 -1287
rect -2779 -1321 -2773 -1287
rect -2711 -1321 -2701 -1287
rect -2643 -1321 -2629 -1287
rect -2575 -1321 -2557 -1287
rect -2507 -1321 -2485 -1287
rect -2439 -1321 -2413 -1287
rect -2371 -1321 -2341 -1287
rect -2303 -1321 -2269 -1287
rect -2235 -1321 -2201 -1287
rect -2163 -1321 -2133 -1287
rect -2091 -1321 -2065 -1287
rect -2019 -1321 -1997 -1287
rect -1947 -1321 -1929 -1287
rect -1875 -1321 -1861 -1287
rect -1803 -1321 -1793 -1287
rect -1731 -1321 -1725 -1287
rect -1659 -1321 -1657 -1287
rect -1623 -1321 -1621 -1287
rect -1555 -1321 -1549 -1287
rect -1487 -1321 -1477 -1287
rect -1419 -1321 -1405 -1287
rect -1351 -1321 -1333 -1287
rect -1283 -1321 -1261 -1287
rect -1215 -1321 -1189 -1287
rect -1147 -1321 -1117 -1287
rect -1079 -1321 -1045 -1287
rect -1011 -1321 -977 -1287
rect -939 -1321 -909 -1287
rect -867 -1321 -841 -1287
rect -795 -1321 -773 -1287
rect -723 -1321 -705 -1287
rect -651 -1321 -637 -1287
rect -579 -1321 -569 -1287
rect -507 -1321 -501 -1287
rect -435 -1321 -433 -1287
rect -399 -1321 -397 -1287
rect -331 -1321 -325 -1287
rect -263 -1321 -253 -1287
rect -195 -1321 -181 -1287
rect -127 -1321 -109 -1287
rect -75 -1321 42 -1287
rect -3322 -1354 42 -1321
rect 892 -1409 2250 -1376
rect -1347 -1448 -1259 -1414
rect -1225 -1448 -1187 -1414
rect -1153 -1448 -1115 -1414
rect -1081 -1448 -1043 -1414
rect -1009 -1448 -971 -1414
rect -937 -1448 -899 -1414
rect -865 -1448 -827 -1414
rect -793 -1448 -755 -1414
rect -721 -1448 -683 -1414
rect -649 -1448 -611 -1414
rect -577 -1448 -539 -1414
rect -505 -1448 -467 -1414
rect -433 -1448 -395 -1414
rect -361 -1448 -323 -1414
rect -289 -1448 -251 -1414
rect -217 -1448 -179 -1414
rect -145 -1448 -107 -1414
rect -73 -1415 -12 -1414
rect -73 -1448 40 -1415
rect -1347 -1449 -1340 -1448
rect -1344 -1450 -1340 -1449
rect -1374 -1485 -1340 -1484
rect 6 -1495 40 -1448
rect 892 -1443 1014 -1409
rect 1048 -1443 1086 -1409
rect 1121 -1443 1155 -1409
rect 1192 -1443 1223 -1409
rect 1264 -1443 1291 -1409
rect 1336 -1443 1359 -1409
rect 1408 -1443 1427 -1409
rect 1480 -1443 1495 -1409
rect 1552 -1443 1563 -1409
rect 1624 -1443 1631 -1409
rect 1696 -1443 1699 -1409
rect 1733 -1443 1734 -1409
rect 1801 -1443 1806 -1409
rect 1869 -1443 1878 -1409
rect 1937 -1443 1950 -1409
rect 2005 -1443 2022 -1409
rect 2056 -1443 2094 -1409
rect 2128 -1443 2250 -1409
rect 892 -1476 2250 -1443
rect -1076 -1512 -1026 -1501
rect -948 -1512 -898 -1501
rect -820 -1512 -770 -1501
rect -692 -1507 -642 -1501
rect -564 -1507 -514 -1501
rect -436 -1507 -386 -1501
rect -308 -1507 -258 -1501
rect -702 -1512 -119 -1507
rect -1374 -1557 -1340 -1519
rect -1272 -1525 -119 -1512
rect -1272 -1559 -1259 -1525
rect -1225 -1559 -1068 -1525
rect -1034 -1559 -940 -1525
rect -906 -1559 -812 -1525
rect -778 -1559 -684 -1525
rect -650 -1559 -556 -1525
rect -522 -1559 -428 -1525
rect -394 -1559 -300 -1525
rect -266 -1559 -171 -1525
rect -137 -1559 -119 -1525
rect -1272 -1572 -119 -1559
rect -1076 -1583 -1026 -1572
rect -948 -1583 -898 -1572
rect -820 -1583 -770 -1572
rect -702 -1577 -119 -1572
rect 6 -1532 40 -1506
rect -692 -1583 -642 -1577
rect -564 -1583 -514 -1577
rect -436 -1583 -386 -1577
rect -308 -1583 -258 -1577
rect -1374 -1629 -1340 -1591
rect -1374 -1701 -1340 -1663
rect -1374 -1773 -1340 -1735
rect 6 -1604 40 -1566
rect 6 -1676 40 -1638
rect 892 -1534 992 -1476
rect 1494 -1532 1652 -1526
rect 1848 -1532 1888 -1526
rect 892 -1598 925 -1534
rect 959 -1598 992 -1534
rect 1248 -1542 1308 -1532
rect 1242 -1545 1314 -1542
rect 1242 -1579 1261 -1545
rect 1295 -1579 1314 -1545
rect 1242 -1582 1314 -1579
rect 1484 -1545 1662 -1532
rect 1484 -1579 1497 -1545
rect 1531 -1579 1615 -1545
rect 1649 -1579 1662 -1545
rect 1248 -1592 1308 -1582
rect 1484 -1592 1662 -1579
rect 1838 -1545 1898 -1532
rect 1838 -1579 1851 -1545
rect 1885 -1579 1898 -1545
rect 1838 -1592 1898 -1579
rect 2150 -1534 2250 -1476
rect 1494 -1598 1652 -1592
rect 1848 -1598 1888 -1592
rect 892 -1606 992 -1598
rect 6 -1748 40 -1710
rect -1374 -1845 -1340 -1807
rect -1374 -1917 -1340 -1879
rect -1277 -1862 -1207 -1785
rect -125 -1862 -55 -1791
rect -1277 -1863 -1188 -1862
rect -132 -1863 -55 -1862
rect -1277 -1869 -1154 -1863
rect -180 -1869 -55 -1863
rect -1277 -1883 -1144 -1869
rect -1277 -1917 -1258 -1883
rect -1224 -1887 -1144 -1883
rect -1224 -1917 -1196 -1887
rect -1277 -1921 -1196 -1917
rect -1162 -1921 -1144 -1887
rect -1277 -1939 -1144 -1921
rect -190 -1883 -55 -1869
rect -190 -1887 -110 -1883
rect -190 -1921 -172 -1887
rect -138 -1917 -110 -1887
rect -76 -1917 -55 -1883
rect -138 -1921 -55 -1917
rect -190 -1939 -55 -1921
rect 6 -1820 40 -1782
rect 6 -1892 40 -1854
rect -1204 -1945 -1154 -1939
rect -180 -1945 -130 -1939
rect -1374 -1952 -1340 -1951
rect 6 -1952 40 -1926
rect 424 -1676 458 -1654
rect 424 -1748 458 -1710
rect 424 -1820 458 -1782
rect 424 -1892 458 -1854
rect 424 -1948 458 -1926
rect 770 -1676 804 -1654
rect 770 -1748 804 -1710
rect 770 -1820 804 -1782
rect 770 -1892 804 -1854
rect 770 -1948 804 -1926
rect 892 -1666 925 -1606
rect 959 -1666 992 -1606
rect 892 -1678 992 -1666
rect 892 -1734 925 -1678
rect 959 -1734 992 -1678
rect 1542 -1682 1602 -1598
rect 2150 -1602 2183 -1534
rect 2217 -1602 2250 -1534
rect 2150 -1606 2250 -1602
rect 2150 -1670 2183 -1606
rect 2217 -1670 2250 -1606
rect 2150 -1678 2250 -1670
rect 892 -1750 992 -1734
rect 892 -1802 925 -1750
rect 959 -1802 992 -1750
rect 892 -1822 992 -1802
rect 892 -1870 925 -1822
rect 959 -1870 992 -1822
rect 892 -1894 992 -1870
rect 2150 -1738 2183 -1678
rect 2217 -1738 2250 -1678
rect 2150 -1750 2250 -1738
rect 2150 -1806 2183 -1750
rect 2217 -1806 2250 -1750
rect 2150 -1822 2250 -1806
rect 2150 -1874 2183 -1822
rect 2217 -1874 2250 -1822
rect 892 -1938 925 -1894
rect 959 -1938 992 -1894
rect 1080 -1896 1120 -1890
rect 892 -1966 992 -1938
rect 1070 -1909 1130 -1896
rect 1376 -1898 1416 -1892
rect 1730 -1898 1770 -1892
rect 2028 -1896 2068 -1890
rect 2150 -1894 2250 -1874
rect 1070 -1943 1083 -1909
rect 1117 -1943 1130 -1909
rect 1070 -1956 1130 -1943
rect 1366 -1911 1500 -1898
rect 1366 -1945 1379 -1911
rect 1413 -1945 1453 -1911
rect 1487 -1945 1500 -1911
rect 1080 -1962 1120 -1956
rect 1366 -1958 1500 -1945
rect 1664 -1911 1780 -1898
rect 1664 -1945 1673 -1911
rect 1707 -1945 1733 -1911
rect 1767 -1945 1780 -1911
rect 1664 -1958 1780 -1945
rect 2018 -1909 2078 -1896
rect 2018 -1943 2031 -1909
rect 2065 -1943 2078 -1909
rect 2018 -1956 2078 -1943
rect 2150 -1942 2183 -1894
rect 2217 -1942 2250 -1894
rect 1376 -1964 1416 -1958
rect 1730 -1964 1770 -1958
rect 2028 -1962 2068 -1956
rect -1280 -2030 -1261 -1996
rect -1227 -2030 -1189 -1996
rect -1155 -2030 -1117 -1996
rect -1083 -2030 -1045 -1996
rect -1011 -2030 -973 -1996
rect -939 -2030 -901 -1996
rect -867 -2030 -829 -1996
rect -795 -2030 -757 -1996
rect -723 -2030 -685 -1996
rect -651 -2030 -613 -1996
rect -579 -2030 -541 -1996
rect -507 -2030 -469 -1996
rect -435 -2030 -397 -1996
rect -363 -2030 -325 -1996
rect -291 -2030 -253 -1996
rect -219 -2030 -181 -1996
rect -147 -2030 -109 -1996
rect -75 -2030 -56 -1996
rect 892 -2006 925 -1966
rect 959 -2006 992 -1966
rect 892 -2038 992 -2006
rect 892 -2074 925 -2038
rect 959 -2074 992 -2038
rect 892 -2110 992 -2074
rect 892 -2144 925 -2110
rect 959 -2144 992 -2110
rect 892 -2182 992 -2144
rect 892 -2216 925 -2182
rect 959 -2216 992 -2182
rect 892 -2254 992 -2216
rect 892 -2288 925 -2254
rect 959 -2288 992 -2254
rect 892 -2326 992 -2288
rect 892 -2360 925 -2326
rect 959 -2360 992 -2326
rect 892 -2398 992 -2360
rect 892 -2432 925 -2398
rect 959 -2432 992 -2398
rect 892 -2470 992 -2432
rect 892 -2504 925 -2470
rect 959 -2504 992 -2470
rect 892 -2542 992 -2504
rect 892 -2576 925 -2542
rect 959 -2576 992 -2542
rect 892 -2634 992 -2576
rect 2150 -1966 2250 -1942
rect 2328 -1676 2362 -1654
rect 2328 -1748 2362 -1710
rect 2328 -1820 2362 -1782
rect 2328 -1892 2362 -1854
rect 2328 -1948 2362 -1926
rect 2674 -1676 2708 -1654
rect 2674 -1748 2708 -1710
rect 2674 -1820 2708 -1782
rect 2674 -1892 2708 -1854
rect 2674 -1948 2708 -1926
rect 2150 -2010 2183 -1966
rect 2217 -2010 2250 -1966
rect 2150 -2038 2250 -2010
rect 2150 -2078 2183 -2038
rect 2217 -2078 2250 -2038
rect 2150 -2110 2250 -2078
rect 2150 -2146 2183 -2110
rect 2217 -2146 2250 -2110
rect 2150 -2182 2250 -2146
rect 2150 -2216 2183 -2182
rect 2217 -2216 2250 -2182
rect 2150 -2254 2250 -2216
rect 2150 -2288 2183 -2254
rect 2217 -2288 2250 -2254
rect 2150 -2326 2250 -2288
rect 2150 -2360 2183 -2326
rect 2217 -2360 2250 -2326
rect 2150 -2398 2250 -2360
rect 2150 -2432 2183 -2398
rect 2217 -2432 2250 -2398
rect 2150 -2470 2250 -2432
rect 2150 -2504 2183 -2470
rect 2217 -2504 2250 -2470
rect 2150 -2542 2250 -2504
rect 2150 -2576 2183 -2542
rect 2217 -2576 2250 -2542
rect 2150 -2634 2250 -2576
rect 892 -2667 2250 -2634
rect 892 -2701 1014 -2667
rect 1048 -2701 1081 -2667
rect 1120 -2701 1149 -2667
rect 1192 -2701 1217 -2667
rect 1264 -2701 1285 -2667
rect 1336 -2701 1353 -2667
rect 1408 -2701 1421 -2667
rect 1480 -2701 1489 -2667
rect 1552 -2701 1557 -2667
rect 1624 -2701 1625 -2667
rect 1659 -2701 1662 -2667
rect 1727 -2701 1734 -2667
rect 1795 -2701 1806 -2667
rect 1863 -2701 1878 -2667
rect 1931 -2701 1950 -2667
rect 1999 -2701 2022 -2667
rect 2056 -2701 2094 -2667
rect 2128 -2701 2250 -2667
rect 892 -2734 2250 -2701
<< viali >>
rect -3205 1923 -3171 1957
rect -3133 1923 -3119 1957
rect -3119 1923 -3099 1957
rect -3061 1923 -3051 1957
rect -3051 1923 -3027 1957
rect -2989 1923 -2983 1957
rect -2983 1923 -2955 1957
rect -2917 1923 -2915 1957
rect -2915 1923 -2883 1957
rect -2845 1923 -2813 1957
rect -2813 1923 -2811 1957
rect -2773 1923 -2745 1957
rect -2745 1923 -2739 1957
rect -2701 1923 -2677 1957
rect -2677 1923 -2667 1957
rect -2629 1923 -2609 1957
rect -2609 1923 -2595 1957
rect -2557 1923 -2541 1957
rect -2541 1923 -2523 1957
rect -2485 1923 -2473 1957
rect -2473 1923 -2451 1957
rect -2413 1923 -2405 1957
rect -2405 1923 -2379 1957
rect -2341 1923 -2337 1957
rect -2337 1923 -2307 1957
rect -2269 1923 -2235 1957
rect -2197 1923 -2167 1957
rect -2167 1923 -2163 1957
rect -2125 1923 -2099 1957
rect -2099 1923 -2091 1957
rect -2053 1923 -2031 1957
rect -2031 1923 -2019 1957
rect -1981 1923 -1963 1957
rect -1963 1923 -1947 1957
rect -1909 1923 -1895 1957
rect -1895 1923 -1875 1957
rect -1837 1923 -1827 1957
rect -1827 1923 -1803 1957
rect -1765 1923 -1759 1957
rect -1759 1923 -1731 1957
rect -1693 1923 -1691 1957
rect -1691 1923 -1659 1957
rect -1621 1923 -1589 1957
rect -1589 1923 -1587 1957
rect -1549 1923 -1521 1957
rect -1521 1923 -1515 1957
rect -1477 1923 -1453 1957
rect -1453 1923 -1443 1957
rect -1405 1923 -1385 1957
rect -1385 1923 -1371 1957
rect -1333 1923 -1317 1957
rect -1317 1923 -1299 1957
rect -1261 1923 -1249 1957
rect -1249 1923 -1227 1957
rect -1189 1923 -1181 1957
rect -1181 1923 -1155 1957
rect -1117 1923 -1113 1957
rect -1113 1923 -1083 1957
rect -1045 1923 -1011 1957
rect -973 1923 -943 1957
rect -943 1923 -939 1957
rect -901 1923 -875 1957
rect -875 1923 -867 1957
rect -829 1923 -807 1957
rect -807 1923 -795 1957
rect -757 1923 -739 1957
rect -739 1923 -723 1957
rect -685 1923 -671 1957
rect -671 1923 -651 1957
rect -613 1923 -603 1957
rect -603 1923 -579 1957
rect -541 1923 -535 1957
rect -535 1923 -507 1957
rect -469 1923 -467 1957
rect -467 1923 -435 1957
rect -397 1923 -365 1957
rect -365 1923 -363 1957
rect -325 1923 -297 1957
rect -297 1923 -291 1957
rect -253 1923 -229 1957
rect -229 1923 -219 1957
rect -181 1923 -161 1957
rect -161 1923 -147 1957
rect -109 1923 -75 1957
rect -3289 1729 -3255 1739
rect -3289 1705 -3255 1729
rect -3289 1661 -3255 1667
rect -3289 1633 -3255 1661
rect -3289 1593 -3255 1595
rect -3289 1561 -3255 1593
rect -3289 1491 -3255 1523
rect -3289 1489 -3255 1491
rect -3289 1423 -3255 1451
rect -3289 1417 -3255 1423
rect -3289 1355 -3255 1379
rect -3289 1345 -3255 1355
rect -3289 1287 -3255 1307
rect -3289 1273 -3255 1287
rect -3289 1219 -3255 1235
rect -3289 1201 -3255 1219
rect -3289 1151 -3255 1163
rect -3289 1129 -3255 1151
rect -3289 1083 -3255 1091
rect -3289 1057 -3255 1083
rect -3289 1015 -3255 1019
rect -3289 985 -3255 1015
rect -3289 913 -3255 947
rect -3289 845 -3255 875
rect -3289 841 -3255 845
rect -3289 777 -3255 803
rect -3289 769 -3255 777
rect -3289 709 -3255 731
rect -3289 697 -3255 709
rect -3289 641 -3255 659
rect -3289 625 -3255 641
rect -3289 573 -3255 587
rect -3289 553 -3255 573
rect -3289 505 -3255 515
rect -3289 481 -3255 505
rect -3289 437 -3255 443
rect -3289 409 -3255 437
rect -3289 369 -3255 371
rect -3289 337 -3255 369
rect -3289 267 -3255 299
rect -3289 265 -3255 267
rect -3289 199 -3255 227
rect -3289 193 -3255 199
rect -3289 131 -3255 155
rect -3289 121 -3255 131
rect -3289 63 -3255 83
rect -3289 49 -3255 63
rect -3289 -5 -3255 11
rect -3289 -23 -3255 -5
rect -3289 -73 -3255 -61
rect -3289 -95 -3255 -73
rect -3289 -141 -3255 -133
rect -3289 -167 -3255 -141
rect -3289 -209 -3255 -205
rect -3289 -239 -3255 -209
rect -3289 -311 -3255 -277
rect -3289 -379 -3255 -349
rect -3289 -383 -3255 -379
rect -3289 -447 -3255 -421
rect -3289 -455 -3255 -447
rect -3289 -515 -3255 -493
rect -3289 -527 -3255 -515
rect -3289 -583 -3255 -565
rect -3289 -599 -3255 -583
rect -3289 -651 -3255 -637
rect -3289 -671 -3255 -651
rect -3289 -719 -3255 -709
rect -3289 -743 -3255 -719
rect -3289 -787 -3255 -781
rect -3289 -815 -3255 -787
rect -3289 -855 -3255 -853
rect -3289 -887 -3255 -855
rect -3289 -957 -3255 -925
rect -3289 -959 -3255 -957
rect -3289 -1025 -3255 -997
rect -3289 -1031 -3255 -1025
rect -3289 -1093 -3255 -1069
rect -3289 -1103 -3255 -1093
rect -25 1729 9 1739
rect -25 1705 9 1729
rect -25 1661 9 1667
rect -25 1633 9 1661
rect -25 1593 9 1595
rect -25 1561 9 1593
rect -25 1491 9 1523
rect -25 1489 9 1491
rect -25 1423 9 1451
rect -25 1417 9 1423
rect -25 1355 9 1379
rect -25 1345 9 1355
rect -25 1287 9 1307
rect -25 1273 9 1287
rect -25 1219 9 1235
rect -25 1201 9 1219
rect -25 1151 9 1163
rect -25 1129 9 1151
rect -25 1083 9 1091
rect -25 1057 9 1083
rect -25 1015 9 1019
rect -25 985 9 1015
rect -25 913 9 947
rect -25 845 9 875
rect -25 841 9 845
rect -25 777 9 803
rect -25 769 9 777
rect -25 709 9 731
rect -25 697 9 709
rect -25 641 9 659
rect -25 625 9 641
rect -25 573 9 587
rect -25 553 9 573
rect -25 505 9 515
rect -25 481 9 505
rect -25 437 9 443
rect -25 409 9 437
rect -25 369 9 371
rect -25 337 9 369
rect -25 267 9 299
rect -25 265 9 267
rect -25 199 9 227
rect -25 193 9 199
rect -25 131 9 155
rect -25 121 9 131
rect -25 63 9 83
rect -25 49 9 63
rect -25 -5 9 11
rect -25 -23 9 -5
rect -25 -73 9 -61
rect -25 -95 9 -73
rect -25 -141 9 -133
rect -25 -167 9 -141
rect -25 -209 9 -205
rect -25 -239 9 -209
rect -25 -311 9 -277
rect -25 -379 9 -349
rect -25 -383 9 -379
rect -25 -447 9 -421
rect -25 -455 9 -447
rect -25 -515 9 -493
rect -25 -527 9 -515
rect 485 1923 519 1957
rect 557 1923 579 1957
rect 579 1923 591 1957
rect 629 1923 647 1957
rect 647 1923 663 1957
rect 701 1923 715 1957
rect 715 1923 735 1957
rect 773 1923 783 1957
rect 783 1923 807 1957
rect 845 1923 851 1957
rect 851 1923 879 1957
rect 917 1923 919 1957
rect 919 1923 951 1957
rect 989 1923 1021 1957
rect 1021 1923 1023 1957
rect 1061 1923 1089 1957
rect 1089 1923 1095 1957
rect 1133 1923 1157 1957
rect 1157 1923 1167 1957
rect 1205 1923 1225 1957
rect 1225 1923 1239 1957
rect 1277 1923 1293 1957
rect 1293 1923 1311 1957
rect 1349 1923 1361 1957
rect 1361 1923 1383 1957
rect 1421 1923 1429 1957
rect 1429 1923 1455 1957
rect 1493 1923 1497 1957
rect 1497 1923 1527 1957
rect 1565 1923 1599 1957
rect 1637 1923 1667 1957
rect 1667 1923 1671 1957
rect 1709 1923 1735 1957
rect 1735 1923 1743 1957
rect 1781 1923 1803 1957
rect 1803 1923 1815 1957
rect 1853 1923 1871 1957
rect 1871 1923 1887 1957
rect 1925 1923 1939 1957
rect 1939 1923 1959 1957
rect 1997 1923 2007 1957
rect 2007 1923 2031 1957
rect 2069 1923 2075 1957
rect 2075 1923 2103 1957
rect 2141 1923 2143 1957
rect 2143 1923 2175 1957
rect 2213 1923 2245 1957
rect 2245 1923 2247 1957
rect 2285 1923 2313 1957
rect 2313 1923 2319 1957
rect 2357 1923 2381 1957
rect 2381 1923 2391 1957
rect 2429 1923 2449 1957
rect 2449 1923 2463 1957
rect 2501 1923 2517 1957
rect 2517 1923 2535 1957
rect 2573 1923 2585 1957
rect 2585 1923 2607 1957
rect 2645 1923 2679 1957
rect 413 1752 447 1776
rect 413 1742 447 1752
rect 413 1684 447 1704
rect 413 1670 447 1684
rect 413 1616 447 1632
rect 413 1598 447 1616
rect 413 1548 447 1560
rect 413 1526 447 1548
rect 413 1480 447 1488
rect 413 1454 447 1480
rect 413 1412 447 1416
rect 413 1382 447 1412
rect 413 1310 447 1344
rect 413 1242 447 1272
rect 413 1238 447 1242
rect 413 1174 447 1200
rect 413 1166 447 1174
rect 413 1106 447 1128
rect 413 1094 447 1106
rect 413 1038 447 1056
rect 413 1022 447 1038
rect 413 970 447 984
rect 413 950 447 970
rect 413 902 447 912
rect 413 878 447 902
rect 413 834 447 840
rect 413 806 447 834
rect 413 766 447 768
rect 413 734 447 766
rect 413 664 447 696
rect 413 662 447 664
rect 413 596 447 624
rect 413 590 447 596
rect 413 528 447 552
rect 413 518 447 528
rect 413 460 447 480
rect 413 446 447 460
rect 413 392 447 408
rect 413 374 447 392
rect 413 324 447 336
rect 413 302 447 324
rect 413 256 447 264
rect 413 230 447 256
rect 413 188 447 192
rect 413 158 447 188
rect 413 86 447 120
rect 413 18 447 48
rect 413 14 447 18
rect 413 -50 447 -24
rect 413 -58 447 -50
rect 413 -118 447 -96
rect 413 -130 447 -118
rect 413 -186 447 -168
rect 413 -202 447 -186
rect 413 -254 447 -240
rect 413 -274 447 -254
rect 413 -322 447 -312
rect 413 -346 447 -322
rect 2719 1786 2751 1789
rect 2751 1786 2753 1789
rect 2719 1755 2753 1786
rect 2719 1684 2753 1717
rect 2719 1683 2751 1684
rect 2751 1683 2753 1684
rect 2719 1616 2753 1645
rect 2719 1611 2751 1616
rect 2751 1611 2753 1616
rect 2717 1480 2751 1496
rect 2717 1462 2751 1480
rect 2717 1412 2751 1424
rect 2717 1390 2751 1412
rect 2717 1344 2751 1352
rect 2717 1318 2751 1344
rect 2717 1276 2751 1280
rect 2717 1246 2751 1276
rect 2717 1174 2751 1208
rect 2717 1106 2751 1136
rect 2717 1102 2751 1106
rect 2717 1038 2751 1064
rect 2717 1030 2751 1038
rect 2717 970 2751 992
rect 2717 958 2751 970
rect 2717 902 2751 920
rect 2717 886 2751 902
rect 2717 834 2751 848
rect 2717 814 2751 834
rect 2717 766 2751 776
rect 2717 742 2751 766
rect 2717 698 2751 704
rect 2717 670 2751 698
rect 2717 630 2751 632
rect 2717 598 2751 630
rect 2717 528 2751 560
rect 2717 526 2751 528
rect 2717 460 2751 488
rect 2717 454 2751 460
rect 2717 392 2751 416
rect 2717 382 2751 392
rect 2717 324 2751 344
rect 2717 310 2751 324
rect 2717 256 2751 272
rect 2717 238 2751 256
rect 2717 188 2751 200
rect 2717 166 2751 188
rect 2717 120 2751 128
rect 2717 94 2751 120
rect 2717 52 2751 56
rect 2717 22 2751 52
rect 2717 -50 2751 -16
rect 2717 -118 2751 -88
rect 2717 -122 2751 -118
rect 2717 -186 2751 -160
rect 2717 -194 2751 -186
rect 2717 -254 2751 -232
rect 2717 -266 2751 -254
rect 2717 -322 2751 -304
rect 2717 -338 2751 -322
rect 485 -527 519 -493
rect 557 -527 579 -493
rect 579 -527 591 -493
rect 629 -527 647 -493
rect 647 -527 663 -493
rect 701 -527 715 -493
rect 715 -527 735 -493
rect 773 -527 783 -493
rect 783 -527 807 -493
rect 845 -527 851 -493
rect 851 -527 879 -493
rect 917 -527 919 -493
rect 919 -527 951 -493
rect 989 -527 1021 -493
rect 1021 -527 1023 -493
rect 1061 -527 1089 -493
rect 1089 -527 1095 -493
rect 1133 -527 1157 -493
rect 1157 -527 1167 -493
rect 1205 -527 1225 -493
rect 1225 -527 1239 -493
rect 1277 -527 1293 -493
rect 1293 -527 1311 -493
rect 1349 -527 1361 -493
rect 1361 -527 1383 -493
rect 1421 -527 1429 -493
rect 1429 -527 1455 -493
rect 1493 -527 1497 -493
rect 1497 -527 1527 -493
rect 1565 -527 1599 -493
rect 1637 -527 1667 -493
rect 1667 -527 1671 -493
rect 1709 -527 1735 -493
rect 1735 -527 1743 -493
rect 1781 -527 1803 -493
rect 1803 -527 1815 -493
rect 1853 -527 1871 -493
rect 1871 -527 1887 -493
rect 1925 -527 1939 -493
rect 1939 -527 1959 -493
rect 1997 -527 2007 -493
rect 2007 -527 2031 -493
rect 2069 -527 2075 -493
rect 2075 -527 2103 -493
rect 2141 -527 2143 -493
rect 2143 -527 2175 -493
rect 2213 -527 2245 -493
rect 2245 -527 2247 -493
rect 2285 -527 2313 -493
rect 2313 -527 2319 -493
rect 2357 -527 2381 -493
rect 2381 -527 2391 -493
rect 2429 -527 2449 -493
rect 2449 -527 2463 -493
rect 2501 -527 2517 -493
rect 2517 -527 2535 -493
rect 2573 -527 2585 -493
rect 2585 -527 2607 -493
rect 2645 -527 2679 -493
rect -25 -583 9 -565
rect -25 -599 9 -583
rect -25 -651 9 -637
rect -25 -671 9 -651
rect 1480 -638 1514 -604
rect 1572 -638 1606 -604
rect -25 -719 9 -709
rect -25 -743 9 -719
rect -25 -787 9 -781
rect -25 -815 9 -787
rect -25 -855 9 -853
rect -25 -887 9 -855
rect -25 -957 9 -925
rect -25 -959 9 -957
rect 699 -943 733 -909
rect 811 -943 845 -909
rect 971 -943 1005 -909
rect 1079 -943 1113 -909
rect 1211 -943 1245 -909
rect 1385 -943 1419 -909
rect 1674 -950 1708 -916
rect 1859 -945 1893 -911
rect 1973 -945 2007 -911
rect 2089 -943 2123 -909
rect 2249 -943 2283 -909
rect 2361 -943 2395 -909
rect -25 -1025 9 -997
rect -25 -1031 9 -1025
rect -25 -1093 9 -1069
rect -25 -1103 9 -1093
rect 1391 -1061 1425 -1027
rect 1671 -1061 1705 -1027
rect 1480 -1184 1514 -1150
rect 1572 -1182 1606 -1148
rect -3205 -1321 -3171 -1287
rect -3133 -1321 -3119 -1287
rect -3119 -1321 -3099 -1287
rect -3061 -1321 -3051 -1287
rect -3051 -1321 -3027 -1287
rect -2989 -1321 -2983 -1287
rect -2983 -1321 -2955 -1287
rect -2917 -1321 -2915 -1287
rect -2915 -1321 -2883 -1287
rect -2845 -1321 -2813 -1287
rect -2813 -1321 -2811 -1287
rect -2773 -1321 -2745 -1287
rect -2745 -1321 -2739 -1287
rect -2701 -1321 -2677 -1287
rect -2677 -1321 -2667 -1287
rect -2629 -1321 -2609 -1287
rect -2609 -1321 -2595 -1287
rect -2557 -1321 -2541 -1287
rect -2541 -1321 -2523 -1287
rect -2485 -1321 -2473 -1287
rect -2473 -1321 -2451 -1287
rect -2413 -1321 -2405 -1287
rect -2405 -1321 -2379 -1287
rect -2341 -1321 -2337 -1287
rect -2337 -1321 -2307 -1287
rect -2269 -1321 -2235 -1287
rect -2197 -1321 -2167 -1287
rect -2167 -1321 -2163 -1287
rect -2125 -1321 -2099 -1287
rect -2099 -1321 -2091 -1287
rect -2053 -1321 -2031 -1287
rect -2031 -1321 -2019 -1287
rect -1981 -1321 -1963 -1287
rect -1963 -1321 -1947 -1287
rect -1909 -1321 -1895 -1287
rect -1895 -1321 -1875 -1287
rect -1837 -1321 -1827 -1287
rect -1827 -1321 -1803 -1287
rect -1765 -1321 -1759 -1287
rect -1759 -1321 -1731 -1287
rect -1693 -1321 -1691 -1287
rect -1691 -1321 -1659 -1287
rect -1621 -1321 -1589 -1287
rect -1589 -1321 -1587 -1287
rect -1549 -1321 -1521 -1287
rect -1521 -1321 -1515 -1287
rect -1477 -1321 -1453 -1287
rect -1453 -1321 -1443 -1287
rect -1405 -1321 -1385 -1287
rect -1385 -1321 -1371 -1287
rect -1333 -1321 -1317 -1287
rect -1317 -1321 -1299 -1287
rect -1261 -1321 -1249 -1287
rect -1249 -1321 -1227 -1287
rect -1189 -1321 -1181 -1287
rect -1181 -1321 -1155 -1287
rect -1117 -1321 -1113 -1287
rect -1113 -1321 -1083 -1287
rect -1045 -1321 -1011 -1287
rect -973 -1321 -943 -1287
rect -943 -1321 -939 -1287
rect -901 -1321 -875 -1287
rect -875 -1321 -867 -1287
rect -829 -1321 -807 -1287
rect -807 -1321 -795 -1287
rect -757 -1321 -739 -1287
rect -739 -1321 -723 -1287
rect -685 -1321 -671 -1287
rect -671 -1321 -651 -1287
rect -613 -1321 -603 -1287
rect -603 -1321 -579 -1287
rect -541 -1321 -535 -1287
rect -535 -1321 -507 -1287
rect -469 -1321 -467 -1287
rect -467 -1321 -435 -1287
rect -397 -1321 -365 -1287
rect -365 -1321 -363 -1287
rect -325 -1321 -297 -1287
rect -297 -1321 -291 -1287
rect -253 -1321 -229 -1287
rect -229 -1321 -219 -1287
rect -181 -1321 -161 -1287
rect -161 -1321 -147 -1287
rect -109 -1321 -75 -1287
rect -1259 -1448 -1225 -1414
rect -1187 -1448 -1153 -1414
rect -1115 -1448 -1081 -1414
rect -1043 -1448 -1009 -1414
rect -971 -1448 -937 -1414
rect -899 -1448 -865 -1414
rect -827 -1448 -793 -1414
rect -755 -1448 -721 -1414
rect -683 -1448 -649 -1414
rect -611 -1448 -577 -1414
rect -539 -1448 -505 -1414
rect -467 -1448 -433 -1414
rect -395 -1448 -361 -1414
rect -323 -1448 -289 -1414
rect -251 -1448 -217 -1414
rect -179 -1448 -145 -1414
rect -107 -1448 -73 -1414
rect -1374 -1519 -1340 -1485
rect 1014 -1443 1048 -1409
rect 1086 -1443 1087 -1409
rect 1087 -1443 1120 -1409
rect 1158 -1443 1189 -1409
rect 1189 -1443 1192 -1409
rect 1230 -1443 1257 -1409
rect 1257 -1443 1264 -1409
rect 1302 -1443 1325 -1409
rect 1325 -1443 1336 -1409
rect 1374 -1443 1393 -1409
rect 1393 -1443 1408 -1409
rect 1446 -1443 1461 -1409
rect 1461 -1443 1480 -1409
rect 1518 -1443 1529 -1409
rect 1529 -1443 1552 -1409
rect 1590 -1443 1597 -1409
rect 1597 -1443 1624 -1409
rect 1662 -1443 1665 -1409
rect 1665 -1443 1696 -1409
rect 1734 -1443 1767 -1409
rect 1767 -1443 1768 -1409
rect 1806 -1443 1835 -1409
rect 1835 -1443 1840 -1409
rect 1878 -1443 1903 -1409
rect 1903 -1443 1912 -1409
rect 1950 -1443 1971 -1409
rect 1971 -1443 1984 -1409
rect 2022 -1443 2056 -1409
rect 2094 -1443 2128 -1409
rect -1374 -1591 -1340 -1557
rect -1259 -1559 -1225 -1525
rect -171 -1559 -137 -1525
rect 6 -1566 40 -1532
rect -1374 -1663 -1340 -1629
rect -1374 -1735 -1340 -1701
rect -1374 -1807 -1340 -1773
rect 6 -1638 40 -1604
rect 925 -1564 959 -1534
rect 925 -1568 959 -1564
rect 1261 -1579 1295 -1545
rect 1851 -1579 1885 -1545
rect 6 -1710 40 -1676
rect 6 -1782 40 -1748
rect -1374 -1879 -1340 -1845
rect -1374 -1951 -1340 -1917
rect -1258 -1917 -1224 -1883
rect -110 -1917 -76 -1883
rect 6 -1854 40 -1820
rect 6 -1926 40 -1892
rect 424 -1710 458 -1676
rect 424 -1782 458 -1748
rect 424 -1854 458 -1820
rect 424 -1926 458 -1892
rect 770 -1710 804 -1676
rect 770 -1782 804 -1748
rect 770 -1854 804 -1820
rect 770 -1926 804 -1892
rect 925 -1632 959 -1606
rect 925 -1640 959 -1632
rect 925 -1700 959 -1678
rect 925 -1712 959 -1700
rect 2183 -1568 2217 -1534
rect 2183 -1636 2217 -1606
rect 2183 -1640 2217 -1636
rect 925 -1768 959 -1750
rect 925 -1784 959 -1768
rect 925 -1836 959 -1822
rect 925 -1856 959 -1836
rect 2183 -1704 2217 -1678
rect 2183 -1712 2217 -1704
rect 2183 -1772 2217 -1750
rect 2183 -1784 2217 -1772
rect 2183 -1840 2217 -1822
rect 2183 -1856 2217 -1840
rect 925 -1904 959 -1894
rect 925 -1928 959 -1904
rect 1083 -1943 1117 -1909
rect 1453 -1945 1487 -1911
rect 1673 -1945 1707 -1911
rect 2031 -1943 2065 -1909
rect 2183 -1908 2217 -1894
rect 2183 -1928 2217 -1908
rect -1261 -2030 -1227 -1996
rect -1189 -2030 -1155 -1996
rect -1117 -2030 -1083 -1996
rect -1045 -2030 -1011 -1996
rect -973 -2030 -939 -1996
rect -901 -2030 -867 -1996
rect -829 -2030 -795 -1996
rect -757 -2030 -723 -1996
rect -685 -2030 -651 -1996
rect -613 -2030 -579 -1996
rect -541 -2030 -507 -1996
rect -469 -2030 -435 -1996
rect -397 -2030 -363 -1996
rect -325 -2030 -291 -1996
rect -253 -2030 -219 -1996
rect -181 -2030 -147 -1996
rect -109 -2030 -75 -1996
rect 925 -1972 959 -1966
rect 925 -2000 959 -1972
rect 925 -2040 959 -2038
rect 925 -2072 959 -2040
rect 925 -2144 959 -2110
rect 925 -2216 959 -2182
rect 925 -2288 959 -2254
rect 925 -2360 959 -2326
rect 925 -2432 959 -2398
rect 925 -2504 959 -2470
rect 925 -2576 959 -2542
rect 2328 -1710 2362 -1676
rect 2328 -1782 2362 -1748
rect 2328 -1854 2362 -1820
rect 2328 -1926 2362 -1892
rect 2674 -1710 2708 -1676
rect 2674 -1782 2708 -1748
rect 2674 -1854 2708 -1820
rect 2674 -1926 2708 -1892
rect 2183 -1976 2217 -1966
rect 2183 -2000 2217 -1976
rect 2183 -2044 2217 -2038
rect 2183 -2072 2217 -2044
rect 2183 -2112 2217 -2110
rect 2183 -2144 2217 -2112
rect 2183 -2216 2217 -2182
rect 2183 -2288 2217 -2254
rect 2183 -2360 2217 -2326
rect 2183 -2432 2217 -2398
rect 2183 -2504 2217 -2470
rect 2183 -2576 2217 -2542
rect 1014 -2701 1048 -2667
rect 1086 -2701 1115 -2667
rect 1115 -2701 1120 -2667
rect 1158 -2701 1183 -2667
rect 1183 -2701 1192 -2667
rect 1230 -2701 1251 -2667
rect 1251 -2701 1264 -2667
rect 1302 -2701 1319 -2667
rect 1319 -2701 1336 -2667
rect 1374 -2701 1387 -2667
rect 1387 -2701 1408 -2667
rect 1446 -2701 1455 -2667
rect 1455 -2701 1480 -2667
rect 1518 -2701 1523 -2667
rect 1523 -2701 1552 -2667
rect 1590 -2701 1591 -2667
rect 1591 -2701 1624 -2667
rect 1662 -2701 1693 -2667
rect 1693 -2701 1696 -2667
rect 1734 -2701 1761 -2667
rect 1761 -2701 1768 -2667
rect 1806 -2701 1829 -2667
rect 1829 -2701 1840 -2667
rect 1878 -2701 1897 -2667
rect 1897 -2701 1912 -2667
rect 1950 -2701 1965 -2667
rect 1965 -2701 1984 -2667
rect 2022 -2701 2056 -2667
rect 2094 -2701 2128 -2667
<< metal1 >>
rect -3328 1957 48 1996
rect -3328 1923 -3205 1957
rect -3171 1923 -3133 1957
rect -3099 1923 -3061 1957
rect -3027 1923 -2989 1957
rect -2955 1923 -2917 1957
rect -2883 1923 -2845 1957
rect -2811 1923 -2773 1957
rect -2739 1923 -2701 1957
rect -2667 1923 -2629 1957
rect -2595 1923 -2557 1957
rect -2523 1923 -2485 1957
rect -2451 1923 -2413 1957
rect -2379 1923 -2341 1957
rect -2307 1923 -2269 1957
rect -2235 1923 -2197 1957
rect -2163 1923 -2125 1957
rect -2091 1923 -2053 1957
rect -2019 1923 -1981 1957
rect -1947 1923 -1909 1957
rect -1875 1923 -1837 1957
rect -1803 1923 -1765 1957
rect -1731 1923 -1693 1957
rect -1659 1923 -1621 1957
rect -1587 1923 -1549 1957
rect -1515 1923 -1477 1957
rect -1443 1923 -1405 1957
rect -1371 1923 -1333 1957
rect -1299 1923 -1261 1957
rect -1227 1923 -1189 1957
rect -1155 1923 -1117 1957
rect -1083 1923 -1045 1957
rect -1011 1923 -973 1957
rect -939 1923 -901 1957
rect -867 1923 -829 1957
rect -795 1923 -757 1957
rect -723 1923 -685 1957
rect -651 1923 -613 1957
rect -579 1923 -541 1957
rect -507 1923 -469 1957
rect -435 1923 -397 1957
rect -363 1923 -325 1957
rect -291 1923 -253 1957
rect -219 1923 -181 1957
rect -147 1923 -109 1957
rect -75 1923 48 1957
rect -3328 1884 48 1923
rect -3328 1856 -330 1884
rect -3328 1739 -3216 1856
rect -3328 1705 -3289 1739
rect -3255 1705 -3216 1739
rect -3328 1667 -3216 1705
rect -3328 1633 -3289 1667
rect -3255 1633 -3216 1667
rect -3328 1612 -3216 1633
rect -348 1612 -330 1856
rect -3328 1595 -330 1612
rect -3328 1561 -3289 1595
rect -3255 1564 -330 1595
rect -64 1739 48 1884
rect -64 1705 -25 1739
rect 9 1705 48 1739
rect -64 1667 48 1705
rect -64 1633 -25 1667
rect 9 1633 48 1667
rect -64 1595 48 1633
rect -3255 1561 -3216 1564
rect -3328 1523 -3216 1561
rect -3328 1489 -3289 1523
rect -3255 1489 -3216 1523
rect -3328 1451 -3216 1489
rect -3328 1417 -3289 1451
rect -3255 1417 -3216 1451
rect -3328 1379 -3216 1417
rect -3328 1345 -3289 1379
rect -3255 1345 -3216 1379
rect -3328 1307 -3216 1345
rect -3328 1273 -3289 1307
rect -3255 1273 -3216 1307
rect -3328 1235 -3216 1273
rect -3328 1201 -3289 1235
rect -3255 1201 -3216 1235
rect -3328 1163 -3216 1201
rect -3328 1129 -3289 1163
rect -3255 1129 -3216 1163
rect -3328 1091 -3216 1129
rect -3328 1057 -3289 1091
rect -3255 1057 -3216 1091
rect -3328 1019 -3216 1057
rect -3328 985 -3289 1019
rect -3255 985 -3216 1019
rect -3328 947 -3216 985
rect -3328 913 -3289 947
rect -3255 913 -3216 947
rect -3328 875 -3216 913
rect -3328 841 -3289 875
rect -3255 841 -3216 875
rect -3328 803 -3216 841
rect -3328 769 -3289 803
rect -3255 769 -3216 803
rect -3328 731 -3216 769
rect -3328 697 -3289 731
rect -3255 697 -3216 731
rect -3328 659 -3216 697
rect -3328 625 -3289 659
rect -3255 625 -3216 659
rect -3166 710 -3106 1564
rect -2134 1242 -2074 1564
rect -1220 1250 -1160 1564
rect -64 1561 -25 1595
rect 9 1561 48 1595
rect -64 1523 48 1561
rect -64 1489 -25 1523
rect 9 1489 48 1523
rect -64 1451 48 1489
rect -64 1417 -25 1451
rect 9 1417 48 1451
rect -64 1379 48 1417
rect -64 1345 -25 1379
rect 9 1345 48 1379
rect -64 1307 48 1345
rect -64 1273 -25 1307
rect 9 1273 48 1307
rect -64 1235 48 1273
rect -64 1201 -25 1235
rect 9 1201 48 1235
rect -64 1163 48 1201
rect -3048 836 -2988 1122
rect -2820 836 -2760 1042
rect -2590 836 -2530 1144
rect -2364 953 -2304 1043
rect -1908 953 -1848 1044
rect -1676 953 -1616 1136
rect -1450 953 -1390 1040
rect -986 953 -926 1042
rect -2364 893 -926 953
rect -762 836 -702 1137
rect -530 836 -470 1044
rect -304 836 -244 1140
rect -3048 776 -244 836
rect -64 1129 -25 1163
rect 9 1129 48 1163
rect -64 1091 48 1129
rect -64 1057 -25 1091
rect 9 1057 48 1091
rect -64 1019 48 1057
rect -64 985 -25 1019
rect 9 985 48 1019
rect -64 947 48 985
rect -64 913 -25 947
rect 9 913 48 947
rect -64 875 48 913
rect -64 841 -25 875
rect 9 841 48 875
rect -64 803 48 841
rect -3166 650 -2802 710
rect -3328 587 -3216 625
rect -3328 553 -3289 587
rect -3255 553 -3216 587
rect -3328 515 -3216 553
rect -3104 592 -3032 596
rect -3104 540 -3094 592
rect -3042 540 -3032 592
rect -3104 536 -3032 540
rect -3328 481 -3289 515
rect -3255 481 -3216 515
rect -3328 443 -3216 481
rect -3328 409 -3289 443
rect -3255 409 -3216 443
rect -3328 371 -3216 409
rect -3328 337 -3289 371
rect -3255 337 -3216 371
rect -3328 299 -3216 337
rect -3328 265 -3289 299
rect -3255 265 -3216 299
rect -3328 227 -3216 265
rect -3328 193 -3289 227
rect -3255 193 -3216 227
rect -3328 155 -3216 193
rect -3328 121 -3289 155
rect -3255 121 -3216 155
rect -3328 83 -3216 121
rect -3328 49 -3289 83
rect -3255 49 -3216 83
rect -3328 11 -3216 49
rect -3328 -23 -3289 11
rect -3255 -23 -3216 11
rect -3328 -61 -3216 -23
rect -3328 -95 -3289 -61
rect -3255 -95 -3216 -61
rect -3328 -133 -3216 -95
rect -3328 -167 -3289 -133
rect -3255 -167 -3216 -133
rect -3328 -205 -3216 -167
rect -3328 -239 -3289 -205
rect -3255 -239 -3216 -205
rect -3328 -277 -3216 -239
rect -3328 -311 -3289 -277
rect -3255 -311 -3216 -277
rect -3328 -349 -3216 -311
rect -3328 -383 -3289 -349
rect -3255 -383 -3216 -349
rect -3328 -421 -3216 -383
rect -3328 -455 -3289 -421
rect -3255 -455 -3216 -421
rect -3328 -493 -3216 -455
rect -3328 -527 -3289 -493
rect -3255 -527 -3216 -493
rect -3328 -565 -3216 -527
rect -3328 -599 -3289 -565
rect -3255 -599 -3216 -565
rect -3328 -637 -3216 -599
rect -3328 -671 -3289 -637
rect -3255 -671 -3216 -637
rect -3328 -709 -3216 -671
rect -3328 -743 -3289 -709
rect -3255 -743 -3216 -709
rect -3328 -781 -3216 -743
rect -3328 -815 -3289 -781
rect -3255 -815 -3216 -781
rect -3328 -853 -3216 -815
rect -3328 -887 -3289 -853
rect -3255 -887 -3216 -853
rect -3328 -925 -3216 -887
rect -3328 -959 -3289 -925
rect -3255 -959 -3216 -925
rect -3328 -997 -3216 -959
rect -3098 -992 -3038 536
rect -2990 378 -2930 650
rect -2862 452 -2802 650
rect -2986 -192 -2926 50
rect -2862 -192 -2802 -38
rect -2986 -252 -2802 -192
rect -2986 -500 -2926 -252
rect -2862 -404 -2802 -252
rect -2730 -256 -2670 38
rect -2600 -136 -2540 -41
rect -2606 -140 -2534 -136
rect -2606 -192 -2596 -140
rect -2544 -192 -2534 -140
rect -2606 -196 -2534 -192
rect -2736 -260 -2664 -256
rect -2736 -312 -2726 -260
rect -2674 -312 -2664 -260
rect -2736 -316 -2664 -312
rect -2476 -528 -2416 776
rect -2220 710 -2148 714
rect -2220 658 -2210 710
rect -2158 658 -2148 710
rect -2220 654 -2148 658
rect -2350 592 -2278 596
rect -2350 540 -2340 592
rect -2288 540 -2278 592
rect -2350 536 -2278 540
rect -2344 460 -2284 536
rect -2214 336 -2154 654
rect -2092 592 -2020 596
rect -2092 540 -2082 592
rect -2030 540 -2020 592
rect -2092 536 -2020 540
rect -2086 460 -2026 536
rect -2352 -140 -2280 -136
rect -2352 -192 -2342 -140
rect -2290 -192 -2280 -140
rect -2352 -196 -2280 -192
rect -2092 -140 -2020 -136
rect -2092 -192 -2082 -140
rect -2030 -192 -2020 -140
rect -2092 -196 -2020 -192
rect -2346 -408 -2286 -196
rect -2222 -260 -2150 -256
rect -2222 -312 -2212 -260
rect -2160 -312 -2150 -260
rect -2222 -316 -2150 -312
rect -2216 -502 -2156 -316
rect -2086 -406 -2026 -196
rect -1958 -516 -1898 776
rect -1828 -136 -1768 -38
rect -1834 -140 -1762 -136
rect -1834 -192 -1824 -140
rect -1772 -192 -1762 -140
rect -1834 -196 -1762 -192
rect -1700 -256 -1640 60
rect -1570 -136 -1510 -42
rect -1576 -140 -1504 -136
rect -1576 -192 -1566 -140
rect -1514 -192 -1504 -140
rect -1576 -196 -1504 -192
rect -1706 -260 -1634 -256
rect -1706 -312 -1696 -260
rect -1644 -312 -1634 -260
rect -1706 -316 -1634 -312
rect -1442 -526 -1382 776
rect -1190 710 -1118 714
rect -1190 658 -1180 710
rect -1128 658 -1118 710
rect -1190 654 -1118 658
rect -1318 592 -1246 596
rect -1318 540 -1308 592
rect -1256 540 -1246 592
rect -1318 536 -1246 540
rect -1312 454 -1252 536
rect -1184 364 -1124 654
rect -1058 592 -986 596
rect -1058 540 -1048 592
rect -996 540 -986 592
rect -1058 536 -986 540
rect -1052 456 -992 536
rect -1318 -140 -1246 -136
rect -1318 -192 -1308 -140
rect -1256 -192 -1246 -140
rect -1318 -196 -1246 -192
rect -1060 -140 -988 -136
rect -1060 -192 -1050 -140
rect -998 -192 -988 -140
rect -1060 -196 -988 -192
rect -1312 -404 -1252 -196
rect -1190 -260 -1118 -256
rect -1190 -312 -1180 -260
rect -1128 -312 -1118 -260
rect -1190 -316 -1118 -312
rect -1184 -516 -1124 -316
rect -1054 -406 -994 -196
rect -928 -526 -868 776
rect -64 769 -25 803
rect 9 769 48 803
rect -64 731 48 769
rect -298 710 -226 714
rect -298 658 -288 710
rect -236 658 -226 710
rect -298 654 -226 658
rect -64 697 -25 731
rect 9 697 48 731
rect -64 659 48 697
rect -538 592 -350 596
rect -538 540 -470 592
rect -418 540 -350 592
rect -538 536 -350 540
rect -538 454 -478 536
rect -410 352 -350 536
rect -796 -136 -736 -42
rect -802 -140 -730 -136
rect -802 -192 -792 -140
rect -740 -192 -730 -140
rect -802 -196 -730 -192
rect -672 -256 -612 84
rect -538 -198 -478 -42
rect -410 -198 -350 64
rect -678 -260 -606 -256
rect -678 -312 -668 -260
rect -616 -312 -606 -260
rect -678 -316 -606 -312
rect -538 -258 -350 -198
rect -538 -404 -478 -258
rect -410 -504 -350 -258
rect -2990 -988 -2930 -792
rect -2860 -988 -2800 -900
rect -3328 -1031 -3289 -997
rect -3255 -1031 -3216 -997
rect -3328 -1069 -3216 -1031
rect -3104 -996 -3032 -992
rect -3104 -1048 -3094 -996
rect -3042 -1048 -3032 -996
rect -2990 -1048 -2800 -988
rect -2730 -1026 -2670 -810
rect -2604 -992 -2544 -901
rect -1828 -992 -1768 -902
rect -3104 -1052 -3032 -1048
rect -3328 -1103 -3289 -1069
rect -3255 -1103 -3216 -1069
rect -3328 -1248 -3216 -1103
rect -2732 -1108 -2670 -1026
rect -2610 -996 -2538 -992
rect -2610 -1048 -2600 -996
rect -2548 -1048 -2538 -996
rect -2610 -1052 -2538 -1048
rect -1834 -996 -1762 -992
rect -1834 -1048 -1824 -996
rect -1772 -1048 -1762 -996
rect -1834 -1052 -1762 -1048
rect -2738 -1112 -2666 -1108
rect -2738 -1164 -2728 -1112
rect -2676 -1164 -2666 -1112
rect -2738 -1168 -2666 -1164
rect -1700 -1114 -1640 -792
rect -1572 -992 -1512 -902
rect -800 -992 -740 -898
rect -1578 -996 -1506 -992
rect -1578 -1048 -1568 -996
rect -1516 -1048 -1506 -996
rect -1578 -1052 -1506 -1048
rect -806 -996 -734 -992
rect -806 -1048 -796 -996
rect -744 -1048 -734 -996
rect -806 -1052 -734 -1048
rect -1700 -1166 -1696 -1114
rect -1644 -1166 -1640 -1114
rect -1700 -1176 -1640 -1166
rect -670 -1114 -610 -798
rect -538 -990 -478 -904
rect -412 -990 -352 -800
rect -538 -1050 -352 -990
rect -670 -1166 -666 -1114
rect -614 -1166 -610 -1114
rect -670 -1176 -610 -1166
rect -292 -1114 -232 654
rect -292 -1166 -288 -1114
rect -236 -1166 -232 -1114
rect -292 -1176 -232 -1166
rect -64 625 -25 659
rect 9 625 48 659
rect -64 587 48 625
rect -64 553 -25 587
rect 9 553 48 587
rect -64 515 48 553
rect -64 481 -25 515
rect 9 481 48 515
rect -64 443 48 481
rect -64 409 -25 443
rect 9 409 48 443
rect 374 1957 2790 1996
rect 374 1923 485 1957
rect 519 1923 557 1957
rect 591 1923 629 1957
rect 663 1923 701 1957
rect 735 1923 773 1957
rect 807 1923 845 1957
rect 879 1923 917 1957
rect 951 1923 989 1957
rect 1023 1923 1061 1957
rect 1095 1923 1133 1957
rect 1167 1923 1205 1957
rect 1239 1923 1277 1957
rect 1311 1923 1349 1957
rect 1383 1923 1421 1957
rect 1455 1923 1493 1957
rect 1527 1923 1565 1957
rect 1599 1923 1637 1957
rect 1671 1923 1709 1957
rect 1743 1923 1781 1957
rect 1815 1923 1853 1957
rect 1887 1923 1925 1957
rect 1959 1923 1997 1957
rect 2031 1923 2069 1957
rect 2103 1923 2141 1957
rect 2175 1923 2213 1957
rect 2247 1923 2285 1957
rect 2319 1923 2357 1957
rect 2391 1923 2429 1957
rect 2463 1923 2501 1957
rect 2535 1923 2573 1957
rect 2607 1923 2645 1957
rect 2679 1923 2790 1957
rect 374 1884 2790 1923
rect 374 1776 486 1884
rect 374 1742 413 1776
rect 447 1742 486 1776
rect 374 1704 486 1742
rect 374 1670 413 1704
rect 447 1670 486 1704
rect 374 1632 486 1670
rect 374 1598 413 1632
rect 447 1598 486 1632
rect 374 1560 486 1598
rect 1038 1856 2790 1884
rect 1038 1612 1072 1856
rect 2660 1789 2790 1856
rect 2660 1755 2719 1789
rect 2753 1755 2790 1789
rect 2660 1717 2790 1755
rect 2660 1683 2719 1717
rect 2753 1683 2790 1717
rect 2660 1645 2790 1683
rect 2660 1612 2719 1645
rect 1038 1611 2719 1612
rect 2753 1611 2790 1645
rect 1038 1564 2790 1611
rect 374 1526 413 1560
rect 447 1526 486 1560
rect 374 1488 486 1526
rect 374 1454 413 1488
rect 447 1454 486 1488
rect 374 1416 486 1454
rect 374 1382 413 1416
rect 447 1382 486 1416
rect 1090 1414 1150 1564
rect 374 1344 486 1382
rect 374 1310 413 1344
rect 447 1310 486 1344
rect 374 1272 486 1310
rect 374 1238 413 1272
rect 447 1238 486 1272
rect 374 1200 486 1238
rect 374 1166 413 1200
rect 447 1166 486 1200
rect 374 1128 486 1166
rect 374 1094 413 1128
rect 447 1094 486 1128
rect 374 1056 486 1094
rect 374 1022 413 1056
rect 447 1022 486 1056
rect 578 1354 1150 1414
rect 578 1024 638 1354
rect 708 1146 768 1354
rect 834 1300 906 1304
rect 834 1248 844 1300
rect 896 1248 906 1300
rect 834 1244 906 1248
rect 840 1038 900 1244
rect 374 984 486 1022
rect 374 950 413 984
rect 447 950 486 984
rect 374 912 486 950
rect 374 878 413 912
rect 447 878 486 912
rect 374 840 486 878
rect 374 806 413 840
rect 447 806 486 840
rect 374 768 486 806
rect 374 734 413 768
rect 447 734 486 768
rect 374 696 486 734
rect 374 662 413 696
rect 447 662 486 696
rect 374 624 486 662
rect 374 590 413 624
rect 447 590 486 624
rect 374 552 486 590
rect 374 518 413 552
rect 447 518 486 552
rect 374 480 486 518
rect 374 446 413 480
rect 447 446 486 480
rect -64 371 48 409
rect -64 337 -25 371
rect 9 337 48 371
rect 248 422 320 426
rect 248 370 258 422
rect 310 370 320 422
rect 248 366 320 370
rect 374 408 486 446
rect 374 374 413 408
rect 447 374 486 408
rect -64 299 48 337
rect -64 265 -25 299
rect 9 265 48 299
rect -64 227 48 265
rect -64 193 -25 227
rect 9 193 48 227
rect -64 155 48 193
rect -64 121 -25 155
rect 9 121 48 155
rect -64 83 48 121
rect -64 49 -25 83
rect 9 49 48 83
rect -64 11 48 49
rect -64 -23 -25 11
rect 9 -23 48 11
rect -64 -61 48 -23
rect -64 -95 -25 -61
rect 9 -95 48 -61
rect -64 -133 48 -95
rect -64 -167 -25 -133
rect 9 -167 48 -133
rect -64 -205 48 -167
rect -64 -239 -25 -205
rect 9 -239 48 -205
rect -64 -277 48 -239
rect -64 -311 -25 -277
rect 9 -311 48 -277
rect -64 -349 48 -311
rect 102 -260 174 -256
rect 102 -312 112 -260
rect 164 -312 174 -260
rect 102 -316 174 -312
rect -64 -383 -25 -349
rect 9 -383 48 -349
rect -64 -421 48 -383
rect -64 -455 -25 -421
rect 9 -455 48 -421
rect -64 -493 48 -455
rect -64 -527 -25 -493
rect 9 -527 48 -493
rect -64 -565 48 -527
rect -64 -599 -25 -565
rect 9 -599 48 -565
rect -64 -637 48 -599
rect -64 -671 -25 -637
rect 9 -671 48 -637
rect -64 -709 48 -671
rect -64 -743 -25 -709
rect 9 -743 48 -709
rect -64 -781 48 -743
rect -64 -815 -25 -781
rect 9 -815 48 -781
rect -64 -853 48 -815
rect -64 -887 -25 -853
rect 9 -887 48 -853
rect -64 -925 48 -887
rect -64 -959 -25 -925
rect 9 -959 48 -925
rect -64 -997 48 -959
rect -64 -1031 -25 -997
rect 9 -1031 48 -997
rect -64 -1069 48 -1031
rect -64 -1103 -25 -1069
rect 9 -1103 48 -1069
rect -64 -1248 48 -1103
rect -3328 -1287 48 -1248
rect -3328 -1321 -3205 -1287
rect -3171 -1321 -3133 -1287
rect -3099 -1321 -3061 -1287
rect -3027 -1321 -2989 -1287
rect -2955 -1321 -2917 -1287
rect -2883 -1321 -2845 -1287
rect -2811 -1321 -2773 -1287
rect -2739 -1321 -2701 -1287
rect -2667 -1321 -2629 -1287
rect -2595 -1321 -2557 -1287
rect -2523 -1321 -2485 -1287
rect -2451 -1321 -2413 -1287
rect -2379 -1321 -2341 -1287
rect -2307 -1321 -2269 -1287
rect -2235 -1321 -2197 -1287
rect -2163 -1321 -2125 -1287
rect -2091 -1321 -2053 -1287
rect -2019 -1321 -1981 -1287
rect -1947 -1321 -1909 -1287
rect -1875 -1321 -1837 -1287
rect -1803 -1321 -1765 -1287
rect -1731 -1321 -1693 -1287
rect -1659 -1321 -1621 -1287
rect -1587 -1321 -1549 -1287
rect -1515 -1321 -1477 -1287
rect -1443 -1321 -1405 -1287
rect -1371 -1321 -1333 -1287
rect -1299 -1321 -1261 -1287
rect -1227 -1321 -1189 -1287
rect -1155 -1321 -1117 -1287
rect -1083 -1321 -1045 -1287
rect -1011 -1321 -973 -1287
rect -939 -1321 -901 -1287
rect -867 -1321 -829 -1287
rect -795 -1321 -757 -1287
rect -723 -1321 -685 -1287
rect -651 -1321 -613 -1287
rect -579 -1321 -541 -1287
rect -507 -1321 -469 -1287
rect -435 -1321 -397 -1287
rect -363 -1321 -325 -1287
rect -291 -1321 -253 -1287
rect -219 -1321 -181 -1287
rect -147 -1321 -109 -1287
rect -75 -1321 48 -1287
rect -3328 -1360 48 -1321
rect -1570 -1402 -1498 -1398
rect -1570 -1454 -1560 -1402
rect -1508 -1454 -1498 -1402
rect -1570 -1458 -1498 -1454
rect -1388 -1414 48 -1360
rect -1388 -1448 -1259 -1414
rect -1225 -1448 -1187 -1414
rect -1153 -1448 -1115 -1414
rect -1081 -1448 -1043 -1414
rect -1009 -1448 -971 -1414
rect -937 -1448 -899 -1414
rect -865 -1448 -827 -1414
rect -793 -1448 -755 -1414
rect -721 -1448 -683 -1414
rect -649 -1448 -611 -1414
rect -577 -1448 -539 -1414
rect -505 -1448 -467 -1414
rect -433 -1448 -395 -1414
rect -361 -1448 -323 -1414
rect -289 -1448 -251 -1414
rect -217 -1448 -179 -1414
rect -145 -1448 -107 -1414
rect -73 -1448 48 -1414
rect -1564 -2076 -1504 -1458
rect -1388 -1462 48 -1448
rect -1388 -1485 -1330 -1462
rect -1388 -1519 -1374 -1485
rect -1340 -1519 -1330 -1485
rect -1278 -1506 -1206 -1500
rect -1388 -1557 -1330 -1519
rect -1388 -1591 -1374 -1557
rect -1340 -1591 -1330 -1557
rect -1284 -1516 -1206 -1506
rect -1284 -1568 -1274 -1516
rect -1222 -1568 -1206 -1516
rect -1284 -1578 -1206 -1568
rect -1278 -1584 -1206 -1578
rect -195 -1501 -113 -1495
rect -195 -1516 -107 -1501
rect -195 -1568 -174 -1516
rect -122 -1568 -107 -1516
rect -195 -1583 -107 -1568
rect -10 -1532 48 -1462
rect -10 -1566 6 -1532
rect 40 -1566 48 -1532
rect -195 -1589 -113 -1583
rect -1388 -1629 -1330 -1591
rect -1388 -1663 -1374 -1629
rect -1340 -1663 -1330 -1629
rect -1388 -1701 -1330 -1663
rect -1388 -1735 -1374 -1701
rect -1340 -1735 -1330 -1701
rect -10 -1604 48 -1566
rect -10 -1638 6 -1604
rect 40 -1638 48 -1604
rect -10 -1676 48 -1638
rect -10 -1710 6 -1676
rect 40 -1710 48 -1676
rect -1388 -1773 -1330 -1735
rect -1388 -1807 -1374 -1773
rect -1340 -1807 -1330 -1773
rect -1152 -1770 -1080 -1766
rect -1388 -1845 -1330 -1807
rect -1388 -1879 -1374 -1845
rect -1340 -1879 -1330 -1845
rect -1276 -1857 -1203 -1786
rect -1152 -1822 -1142 -1770
rect -1090 -1822 -1080 -1770
rect -1152 -1826 -1080 -1822
rect -1388 -1917 -1330 -1879
rect -1388 -1951 -1374 -1917
rect -1340 -1951 -1330 -1917
rect -1289 -1883 -1192 -1857
rect -1289 -1917 -1258 -1883
rect -1224 -1917 -1192 -1883
rect -1289 -1942 -1192 -1917
rect -1016 -1874 -956 -1732
rect -638 -1750 -566 -1746
rect -896 -1760 -824 -1756
rect -896 -1812 -886 -1760
rect -834 -1812 -824 -1760
rect -896 -1816 -824 -1812
rect -762 -1874 -702 -1788
rect -638 -1802 -628 -1750
rect -576 -1802 -566 -1750
rect -386 -1752 -314 -1748
rect -638 -1806 -566 -1802
rect -506 -1874 -446 -1774
rect -386 -1804 -376 -1752
rect -324 -1804 -314 -1752
rect -386 -1808 -314 -1804
rect -252 -1750 -180 -1746
rect -252 -1802 -242 -1750
rect -190 -1802 -180 -1750
rect -10 -1748 48 -1710
rect -252 -1806 -180 -1802
rect -250 -1874 -190 -1806
rect -129 -1856 -54 -1759
rect -10 -1782 6 -1748
rect 40 -1782 48 -1748
rect -10 -1820 48 -1782
rect -10 -1854 6 -1820
rect 40 -1854 48 -1820
rect -1016 -1934 -190 -1874
rect -142 -1883 -43 -1856
rect -142 -1917 -110 -1883
rect -76 -1917 -43 -1883
rect -1388 -1979 -1330 -1951
rect -1276 -1979 -1203 -1942
rect -142 -1943 -43 -1917
rect -10 -1892 48 -1854
rect -10 -1926 6 -1892
rect 40 -1926 48 -1892
rect -129 -1979 -54 -1943
rect -10 -1979 48 -1926
rect -1388 -1996 48 -1979
rect -1388 -2030 -1261 -1996
rect -1227 -2030 -1189 -1996
rect -1155 -2030 -1117 -1996
rect -1083 -2030 -1045 -1996
rect -1011 -2030 -973 -1996
rect -939 -2030 -901 -1996
rect -867 -2030 -829 -1996
rect -795 -2030 -757 -1996
rect -723 -2030 -685 -1996
rect -651 -2030 -613 -1996
rect -579 -2030 -541 -1996
rect -507 -2030 -469 -1996
rect -435 -2030 -397 -1996
rect -363 -2030 -325 -1996
rect -291 -2030 -253 -1996
rect -219 -2030 -181 -1996
rect -147 -2030 -109 -1996
rect -75 -2030 48 -1996
rect -1388 -2038 48 -2030
rect -380 -2076 -320 -2070
rect -1564 -2080 -320 -2076
rect -1564 -2082 -886 -2080
rect -1564 -2134 -1142 -2082
rect -1090 -2132 -886 -2082
rect -834 -2132 -628 -2080
rect -576 -2132 -376 -2080
rect -324 -2132 -320 -2080
rect -1090 -2134 -320 -2132
rect -1564 -2136 -320 -2134
rect -1152 -2138 -1080 -2136
rect -380 -2142 -320 -2136
rect 108 -2100 168 -316
rect 254 -896 314 366
rect 374 336 486 374
rect 374 302 413 336
rect 447 302 486 336
rect 374 264 486 302
rect 374 230 413 264
rect 447 230 486 264
rect 374 192 486 230
rect 374 158 413 192
rect 447 158 486 192
rect 374 120 486 158
rect 374 86 413 120
rect 447 86 486 120
rect 374 48 486 86
rect 374 14 413 48
rect 447 14 486 48
rect 374 -24 486 14
rect 374 -58 413 -24
rect 447 -58 486 -24
rect 374 -96 486 -58
rect 374 -130 413 -96
rect 447 -130 486 -96
rect 374 -168 486 -130
rect 374 -202 413 -168
rect 447 -202 486 -168
rect 374 -240 486 -202
rect 374 -274 413 -240
rect 447 -274 486 -240
rect 374 -312 486 -274
rect 374 -346 413 -312
rect 447 -346 486 -312
rect 374 -454 486 -346
rect 574 492 634 850
rect 708 492 768 644
rect 574 432 768 492
rect 574 -312 634 432
rect 708 278 768 432
rect 964 426 1024 644
rect 834 422 906 426
rect 834 370 844 422
rect 896 370 906 422
rect 834 366 906 370
rect 958 422 1030 426
rect 958 370 968 422
rect 1020 370 1030 422
rect 958 366 1030 370
rect 840 64 900 366
rect 1090 150 1150 1354
rect 1220 1300 1292 1304
rect 1220 1248 1230 1300
rect 1282 1248 1292 1300
rect 1220 1244 1292 1248
rect 1478 1300 1550 1304
rect 1478 1248 1488 1300
rect 1540 1248 1550 1300
rect 1478 1244 1550 1248
rect 1226 1138 1286 1244
rect 1484 1134 1544 1244
rect 1354 426 1414 746
rect 1220 422 1292 426
rect 1220 370 1230 422
rect 1282 370 1292 422
rect 1220 366 1292 370
rect 1348 422 1420 426
rect 1348 370 1358 422
rect 1410 370 1420 422
rect 1348 366 1420 370
rect 1474 422 1546 426
rect 1474 370 1484 422
rect 1536 370 1546 422
rect 1474 366 1546 370
rect 1226 276 1286 366
rect 1480 276 1540 366
rect 1606 154 1666 1564
rect 1862 1300 1934 1304
rect 1862 1248 1872 1300
rect 1924 1248 1934 1300
rect 1862 1244 1934 1248
rect 1868 1046 1928 1244
rect 1738 426 1798 648
rect 1996 494 2056 645
rect 2124 498 2184 1564
rect 2260 498 2320 640
rect 2386 498 2446 1564
rect 2678 1496 2790 1564
rect 2678 1462 2717 1496
rect 2751 1462 2790 1496
rect 2678 1424 2790 1462
rect 2678 1390 2717 1424
rect 2751 1390 2790 1424
rect 2678 1352 2790 1390
rect 2678 1318 2717 1352
rect 2751 1318 2790 1352
rect 2502 1300 2574 1304
rect 2502 1248 2512 1300
rect 2564 1248 2574 1300
rect 2502 1244 2574 1248
rect 2678 1280 2790 1318
rect 2678 1246 2717 1280
rect 2751 1246 2790 1280
rect 1990 490 2062 494
rect 1990 438 2000 490
rect 2052 438 2062 490
rect 1990 434 2062 438
rect 2124 438 2446 498
rect 1732 422 1804 426
rect 1732 370 1742 422
rect 1794 370 1804 422
rect 1732 366 1804 370
rect 1862 422 1934 426
rect 1862 370 1872 422
rect 1924 370 1934 422
rect 1862 366 1934 370
rect 1868 172 1928 366
rect 1996 276 2056 434
rect 2124 172 2184 438
rect 2260 284 2320 438
rect 2386 176 2446 438
rect 712 -312 772 -218
rect 574 -372 772 -312
rect 960 -328 1020 -217
rect 1350 -328 1410 -112
rect 1738 -328 1798 -218
rect 2508 -328 2568 1244
rect 2678 1208 2790 1246
rect 2678 1174 2717 1208
rect 2751 1174 2790 1208
rect 2678 1136 2790 1174
rect 2678 1102 2717 1136
rect 2751 1102 2790 1136
rect 2678 1064 2790 1102
rect 2678 1030 2717 1064
rect 2751 1030 2790 1064
rect 2678 992 2790 1030
rect 2678 958 2717 992
rect 2751 958 2790 992
rect 2678 920 2790 958
rect 2678 886 2717 920
rect 2751 886 2790 920
rect 2678 848 2790 886
rect 2678 814 2717 848
rect 2751 814 2790 848
rect 2678 776 2790 814
rect 2678 742 2717 776
rect 2751 742 2790 776
rect 2678 704 2790 742
rect 2678 670 2717 704
rect 2751 670 2790 704
rect 2678 632 2790 670
rect 2678 598 2717 632
rect 2751 598 2790 632
rect 2678 560 2790 598
rect 2678 526 2717 560
rect 2751 526 2790 560
rect 2678 488 2790 526
rect 2678 454 2717 488
rect 2751 454 2790 488
rect 2678 416 2790 454
rect 2678 382 2717 416
rect 2751 382 2790 416
rect 2678 344 2790 382
rect 2678 310 2717 344
rect 2751 310 2790 344
rect 2678 272 2790 310
rect 2678 238 2717 272
rect 2751 238 2790 272
rect 2678 200 2790 238
rect 2678 166 2717 200
rect 2751 166 2790 200
rect 2678 128 2790 166
rect 2678 94 2717 128
rect 2751 94 2790 128
rect 2678 56 2790 94
rect 2678 22 2717 56
rect 2751 22 2790 56
rect 2678 -16 2790 22
rect 2678 -50 2717 -16
rect 2751 -50 2790 -16
rect 2678 -88 2790 -50
rect 2678 -122 2717 -88
rect 2751 -122 2790 -88
rect 2678 -160 2790 -122
rect 2678 -194 2717 -160
rect 2751 -194 2790 -160
rect 2678 -232 2790 -194
rect 2678 -266 2717 -232
rect 2751 -266 2790 -232
rect 2678 -304 2790 -266
rect 954 -332 1026 -328
rect 954 -384 964 -332
rect 1016 -384 1026 -332
rect 954 -388 1026 -384
rect 1344 -332 1416 -328
rect 1344 -384 1354 -332
rect 1406 -384 1416 -332
rect 1344 -388 1416 -384
rect 1732 -332 1804 -328
rect 1732 -384 1742 -332
rect 1794 -384 1804 -332
rect 1732 -388 1804 -384
rect 2502 -332 2574 -328
rect 2502 -384 2512 -332
rect 2564 -384 2574 -332
rect 2502 -388 2574 -384
rect 2678 -338 2717 -304
rect 2751 -338 2790 -304
rect 2678 -454 2790 -338
rect 374 -493 2790 -454
rect 374 -527 485 -493
rect 519 -527 557 -493
rect 591 -527 629 -493
rect 663 -527 701 -493
rect 735 -527 773 -493
rect 807 -527 845 -493
rect 879 -527 917 -493
rect 951 -527 989 -493
rect 1023 -527 1061 -493
rect 1095 -527 1133 -493
rect 1167 -527 1205 -493
rect 1239 -527 1277 -493
rect 1311 -527 1349 -493
rect 1383 -527 1421 -493
rect 1455 -527 1493 -493
rect 1527 -527 1565 -493
rect 1599 -527 1637 -493
rect 1671 -527 1709 -493
rect 1743 -527 1781 -493
rect 1815 -527 1853 -493
rect 1887 -527 1925 -493
rect 1959 -527 1997 -493
rect 2031 -527 2069 -493
rect 2103 -527 2141 -493
rect 2175 -527 2213 -493
rect 2247 -527 2285 -493
rect 2319 -527 2357 -493
rect 2391 -527 2429 -493
rect 2463 -527 2501 -493
rect 2535 -527 2573 -493
rect 2607 -527 2645 -493
rect 2679 -527 2790 -493
rect 374 -566 2790 -527
rect 626 -604 2470 -566
rect 626 -638 1480 -604
rect 1514 -638 1572 -604
rect 1606 -638 2470 -604
rect 626 -652 2470 -638
rect 2772 -624 2844 -620
rect 1418 -670 1658 -652
rect 2772 -676 2782 -624
rect 2834 -676 2844 -624
rect 2772 -680 2844 -676
rect 798 -896 858 -890
rect 958 -896 1018 -890
rect 254 -909 752 -896
rect 254 -943 699 -909
rect 733 -943 752 -909
rect 254 -956 752 -943
rect 798 -909 1018 -896
rect 798 -943 811 -909
rect 845 -943 971 -909
rect 1005 -943 1018 -909
rect 798 -956 1018 -943
rect 1060 -909 1264 -896
rect 1060 -943 1079 -909
rect 1113 -943 1211 -909
rect 1245 -943 1264 -909
rect 1060 -956 1264 -943
rect 1366 -909 1612 -896
rect 1846 -898 1906 -892
rect 1960 -898 2020 -892
rect 2076 -896 2136 -890
rect 2236 -896 2296 -890
rect 1366 -943 1385 -909
rect 1419 -943 1612 -909
rect 1366 -956 1612 -943
rect 254 -1988 314 -956
rect 798 -962 858 -956
rect 958 -962 1018 -956
rect 1378 -1014 1438 -1008
rect 1552 -1014 1612 -956
rect 1652 -908 1724 -904
rect 1652 -960 1662 -908
rect 1714 -960 1724 -908
rect 1652 -964 1724 -960
rect 1846 -911 2028 -898
rect 1846 -945 1859 -911
rect 1893 -945 1973 -911
rect 2007 -945 2028 -911
rect 1846 -958 2028 -945
rect 2076 -909 2296 -896
rect 2076 -943 2089 -909
rect 2123 -943 2249 -909
rect 2283 -943 2296 -909
rect 2076 -956 2296 -943
rect 1846 -964 1906 -958
rect 1960 -964 2020 -958
rect 2076 -962 2136 -956
rect 2236 -962 2296 -956
rect 2348 -896 2408 -890
rect 2778 -896 2838 -680
rect 2348 -909 2838 -896
rect 2348 -943 2361 -909
rect 2395 -943 2838 -909
rect 2348 -956 2838 -943
rect 2348 -962 2408 -956
rect 1658 -1014 1718 -1008
rect 1372 -1018 1444 -1014
rect 1372 -1070 1382 -1018
rect 1434 -1070 1444 -1018
rect 1372 -1074 1444 -1070
rect 1552 -1027 1718 -1014
rect 1552 -1061 1671 -1027
rect 1705 -1061 1718 -1027
rect 1552 -1074 1718 -1061
rect 1378 -1080 1438 -1074
rect 1658 -1080 1718 -1074
rect 1446 -1120 1686 -1118
rect 972 -1148 2110 -1120
rect 972 -1150 1572 -1148
rect 972 -1184 1480 -1150
rect 1514 -1182 1572 -1150
rect 1606 -1182 2110 -1148
rect 1514 -1184 2110 -1182
rect 972 -1202 2110 -1184
rect 886 -1409 2256 -1202
rect 886 -1443 1014 -1409
rect 1048 -1443 1086 -1409
rect 1120 -1443 1158 -1409
rect 1192 -1443 1230 -1409
rect 1264 -1443 1302 -1409
rect 1336 -1443 1374 -1409
rect 1408 -1443 1446 -1409
rect 1480 -1443 1518 -1409
rect 1552 -1443 1590 -1409
rect 1624 -1443 1662 -1409
rect 1696 -1443 1734 -1409
rect 1768 -1443 1806 -1409
rect 1840 -1443 1878 -1409
rect 1912 -1443 1950 -1409
rect 1984 -1443 2022 -1409
rect 2056 -1443 2094 -1409
rect 2128 -1443 2256 -1409
rect 886 -1482 2256 -1443
rect 886 -1534 998 -1482
rect 886 -1568 925 -1534
rect 959 -1568 998 -1534
rect 558 -1626 670 -1602
rect 412 -1676 472 -1640
rect 412 -1710 424 -1676
rect 458 -1710 472 -1676
rect 558 -1678 588 -1626
rect 640 -1678 670 -1626
rect 886 -1606 998 -1568
rect 1130 -1532 1190 -1526
rect 1242 -1532 1314 -1520
rect 1832 -1532 1904 -1520
rect 1130 -1536 1904 -1532
rect 1130 -1588 1134 -1536
rect 1186 -1545 1904 -1536
rect 1186 -1579 1261 -1545
rect 1295 -1579 1851 -1545
rect 1885 -1579 1904 -1545
rect 1186 -1588 1904 -1579
rect 1130 -1592 1904 -1588
rect 1130 -1598 1190 -1592
rect 1242 -1604 1314 -1592
rect 886 -1640 925 -1606
rect 959 -1640 998 -1606
rect 558 -1702 670 -1678
rect 756 -1676 820 -1642
rect 412 -1748 472 -1710
rect 756 -1710 770 -1676
rect 804 -1710 820 -1676
rect 412 -1782 424 -1748
rect 458 -1782 472 -1748
rect 412 -1820 472 -1782
rect 412 -1854 424 -1820
rect 458 -1854 472 -1820
rect 412 -1892 472 -1854
rect 412 -1926 424 -1892
rect 458 -1926 472 -1892
rect 248 -1992 320 -1988
rect 248 -2044 258 -1992
rect 310 -2044 320 -1992
rect 248 -2048 320 -2044
rect 108 -2152 112 -2100
rect 164 -2152 168 -2100
rect 108 -2162 168 -2152
rect 412 -2282 472 -1926
rect 526 -1988 586 -1764
rect 642 -1794 702 -1734
rect 756 -1748 820 -1710
rect 756 -1782 770 -1748
rect 804 -1782 820 -1748
rect 642 -1926 704 -1794
rect 756 -1820 820 -1782
rect 756 -1854 770 -1820
rect 804 -1854 820 -1820
rect 756 -1892 820 -1854
rect 756 -1926 770 -1892
rect 804 -1926 820 -1892
rect 642 -1988 702 -1926
rect 520 -1992 592 -1988
rect 520 -2044 530 -1992
rect 582 -2044 592 -1992
rect 520 -2048 592 -2044
rect 636 -1992 708 -1988
rect 636 -2044 646 -1992
rect 698 -2044 708 -1992
rect 636 -2048 708 -2044
rect 756 -2282 820 -1926
rect 886 -1678 998 -1640
rect 886 -1712 925 -1678
rect 959 -1712 998 -1678
rect 1424 -1680 1484 -1592
rect 1662 -1672 1722 -1592
rect 1832 -1604 1904 -1592
rect 2144 -1534 2256 -1482
rect 2144 -1568 2183 -1534
rect 2217 -1568 2256 -1534
rect 2144 -1606 2256 -1568
rect 2144 -1640 2183 -1606
rect 2217 -1640 2256 -1606
rect 2144 -1678 2256 -1640
rect 2462 -1628 2574 -1604
rect 886 -1750 998 -1712
rect 886 -1784 925 -1750
rect 959 -1784 998 -1750
rect 886 -1822 998 -1784
rect 2144 -1712 2183 -1678
rect 2217 -1712 2256 -1678
rect 2144 -1750 2256 -1712
rect 2144 -1784 2183 -1750
rect 2217 -1784 2256 -1750
rect 886 -1856 925 -1822
rect 959 -1856 998 -1822
rect 886 -1894 998 -1856
rect 1070 -1884 1130 -1814
rect 886 -1928 925 -1894
rect 959 -1928 998 -1894
rect 886 -1966 998 -1928
rect 886 -2000 925 -1966
rect 959 -2000 998 -1966
rect 1064 -1909 1136 -1884
rect 1064 -1943 1083 -1909
rect 1117 -1943 1136 -1909
rect 1064 -1968 1136 -1943
rect 886 -2038 998 -2000
rect 886 -2072 925 -2038
rect 959 -2072 998 -2038
rect 886 -2110 998 -2072
rect 886 -2144 925 -2110
rect 959 -2144 998 -2110
rect 886 -2182 998 -2144
rect 886 -2216 925 -2182
rect 959 -2216 998 -2182
rect 886 -2254 998 -2216
rect 886 -2282 925 -2254
rect 322 -2288 925 -2282
rect 959 -2280 998 -2254
rect 1070 -2280 1130 -1968
rect 1188 -2098 1248 -1814
rect 1182 -2102 1254 -2098
rect 1182 -2154 1192 -2102
rect 1244 -2154 1254 -2102
rect 1182 -2158 1254 -2154
rect 1310 -2280 1370 -1808
rect 1440 -1898 1500 -1892
rect 1434 -1902 1506 -1898
rect 1434 -1954 1444 -1902
rect 1496 -1954 1506 -1902
rect 1434 -1958 1506 -1954
rect 1440 -1964 1500 -1958
rect 1542 -2280 1602 -1822
rect 1660 -1898 1720 -1892
rect 1654 -1902 1726 -1898
rect 1654 -1954 1664 -1902
rect 1716 -1954 1726 -1902
rect 1654 -1958 1726 -1954
rect 1660 -1964 1720 -1958
rect 1778 -2280 1838 -1810
rect 1896 -2098 1956 -1810
rect 2018 -1884 2078 -1792
rect 2144 -1822 2256 -1784
rect 2144 -1856 2183 -1822
rect 2217 -1856 2256 -1822
rect 2012 -1909 2084 -1884
rect 2012 -1943 2031 -1909
rect 2065 -1943 2084 -1909
rect 2012 -1968 2084 -1943
rect 2144 -1894 2256 -1856
rect 2144 -1928 2183 -1894
rect 2217 -1928 2256 -1894
rect 2144 -1966 2256 -1928
rect 1890 -2102 1962 -2098
rect 1890 -2154 1900 -2102
rect 1952 -2154 1962 -2102
rect 1890 -2158 1962 -2154
rect 2018 -2280 2078 -1968
rect 2144 -2000 2183 -1966
rect 2217 -2000 2256 -1966
rect 2144 -2038 2256 -2000
rect 2144 -2072 2183 -2038
rect 2217 -2072 2256 -2038
rect 2144 -2110 2256 -2072
rect 2144 -2144 2183 -2110
rect 2217 -2144 2256 -2110
rect 2144 -2182 2256 -2144
rect 2144 -2216 2183 -2182
rect 2217 -2216 2256 -2182
rect 2144 -2254 2256 -2216
rect 2144 -2280 2183 -2254
rect 959 -2288 2183 -2280
rect 2217 -2280 2256 -2254
rect 2316 -1676 2376 -1642
rect 2316 -1710 2328 -1676
rect 2362 -1710 2376 -1676
rect 2462 -1680 2492 -1628
rect 2544 -1680 2574 -1628
rect 2462 -1704 2574 -1680
rect 2662 -1676 2722 -1644
rect 2316 -1748 2376 -1710
rect 2316 -1782 2328 -1748
rect 2362 -1782 2376 -1748
rect 2316 -1820 2376 -1782
rect 2316 -1854 2328 -1820
rect 2362 -1854 2376 -1820
rect 2316 -1892 2376 -1854
rect 2662 -1710 2674 -1676
rect 2708 -1710 2722 -1676
rect 2662 -1748 2722 -1710
rect 2662 -1782 2674 -1748
rect 2708 -1782 2722 -1748
rect 2662 -1820 2722 -1782
rect 2662 -1854 2674 -1820
rect 2708 -1854 2722 -1820
rect 2316 -1926 2328 -1892
rect 2362 -1926 2376 -1892
rect 2316 -2280 2376 -1926
rect 2426 -2098 2486 -1884
rect 2546 -1998 2606 -1878
rect 2662 -1892 2722 -1854
rect 2662 -1926 2674 -1892
rect 2708 -1926 2722 -1892
rect 2540 -2002 2612 -1998
rect 2540 -2054 2550 -2002
rect 2602 -2054 2612 -2002
rect 2540 -2058 2612 -2054
rect 2420 -2102 2492 -2098
rect 2420 -2154 2430 -2102
rect 2482 -2154 2492 -2102
rect 2420 -2158 2492 -2154
rect 2662 -2280 2722 -1926
rect 2778 -1998 2838 -956
rect 2772 -2002 2844 -1998
rect 2772 -2054 2782 -2002
rect 2834 -2054 2844 -2002
rect 2772 -2058 2844 -2054
rect 2217 -2288 2810 -2280
rect 322 -2326 2810 -2288
rect 322 -2339 925 -2326
rect 959 -2339 2183 -2326
rect 2217 -2339 2810 -2326
rect 322 -2583 358 -2339
rect 2778 -2583 2810 -2339
rect 322 -2632 2810 -2583
rect 886 -2667 2256 -2632
rect 886 -2701 1014 -2667
rect 1048 -2701 1086 -2667
rect 1120 -2701 1158 -2667
rect 1192 -2701 1230 -2667
rect 1264 -2701 1302 -2667
rect 1336 -2701 1374 -2667
rect 1408 -2701 1446 -2667
rect 1480 -2701 1518 -2667
rect 1552 -2701 1590 -2667
rect 1624 -2701 1662 -2667
rect 1696 -2701 1734 -2667
rect 1768 -2701 1806 -2667
rect 1840 -2701 1878 -2667
rect 1912 -2701 1950 -2667
rect 1984 -2701 2022 -2667
rect 2056 -2701 2094 -2667
rect 2128 -2701 2256 -2667
rect 886 -2740 2256 -2701
<< via1 >>
rect -3216 1612 -348 1856
rect -3094 540 -3042 592
rect -2596 -192 -2544 -140
rect -2726 -312 -2674 -260
rect -2210 658 -2158 710
rect -2340 540 -2288 592
rect -2082 540 -2030 592
rect -2342 -192 -2290 -140
rect -2082 -192 -2030 -140
rect -2212 -312 -2160 -260
rect -1824 -192 -1772 -140
rect -1566 -192 -1514 -140
rect -1696 -312 -1644 -260
rect -1180 658 -1128 710
rect -1308 540 -1256 592
rect -1048 540 -996 592
rect -1308 -192 -1256 -140
rect -1050 -192 -998 -140
rect -1180 -312 -1128 -260
rect -288 658 -236 710
rect -470 540 -418 592
rect -792 -192 -740 -140
rect -668 -312 -616 -260
rect -3094 -1048 -3042 -996
rect -2600 -1048 -2548 -996
rect -1824 -1048 -1772 -996
rect -2728 -1164 -2676 -1112
rect -1568 -1048 -1516 -996
rect -796 -1048 -744 -996
rect -1696 -1166 -1644 -1114
rect -666 -1166 -614 -1114
rect -288 -1166 -236 -1114
rect 1072 1612 2660 1856
rect 844 1248 896 1300
rect 258 370 310 422
rect 112 -312 164 -260
rect -1560 -1454 -1508 -1402
rect -1274 -1525 -1222 -1516
rect -1274 -1559 -1259 -1525
rect -1259 -1559 -1225 -1525
rect -1225 -1559 -1222 -1525
rect -1274 -1568 -1222 -1559
rect -174 -1525 -122 -1516
rect -174 -1559 -171 -1525
rect -171 -1559 -137 -1525
rect -137 -1559 -122 -1525
rect -174 -1568 -122 -1559
rect -1142 -1822 -1090 -1770
rect -886 -1812 -834 -1760
rect -628 -1802 -576 -1750
rect -376 -1804 -324 -1752
rect -242 -1802 -190 -1750
rect -1142 -2134 -1090 -2082
rect -886 -2132 -834 -2080
rect -628 -2132 -576 -2080
rect -376 -2132 -324 -2080
rect 844 370 896 422
rect 968 370 1020 422
rect 1230 1248 1282 1300
rect 1488 1248 1540 1300
rect 1230 370 1282 422
rect 1358 370 1410 422
rect 1484 370 1536 422
rect 1872 1248 1924 1300
rect 2512 1248 2564 1300
rect 2000 438 2052 490
rect 1742 370 1794 422
rect 1872 370 1924 422
rect 964 -384 1016 -332
rect 1354 -384 1406 -332
rect 1742 -384 1794 -332
rect 2512 -384 2564 -332
rect 2782 -676 2834 -624
rect 1662 -916 1714 -908
rect 1662 -950 1674 -916
rect 1674 -950 1708 -916
rect 1708 -950 1714 -916
rect 1662 -960 1714 -950
rect 1382 -1027 1434 -1018
rect 1382 -1061 1391 -1027
rect 1391 -1061 1425 -1027
rect 1425 -1061 1434 -1027
rect 1382 -1070 1434 -1061
rect 588 -1678 640 -1626
rect 1134 -1588 1186 -1536
rect 258 -2044 310 -1992
rect 112 -2152 164 -2100
rect 530 -2044 582 -1992
rect 646 -2044 698 -1992
rect 1192 -2154 1244 -2102
rect 1444 -1911 1496 -1902
rect 1444 -1945 1453 -1911
rect 1453 -1945 1487 -1911
rect 1487 -1945 1496 -1911
rect 1444 -1954 1496 -1945
rect 1664 -1911 1716 -1902
rect 1664 -1945 1673 -1911
rect 1673 -1945 1707 -1911
rect 1707 -1945 1716 -1911
rect 1664 -1954 1716 -1945
rect 1900 -2154 1952 -2102
rect 2492 -1680 2544 -1628
rect 2550 -2054 2602 -2002
rect 2430 -2154 2482 -2102
rect 2782 -2054 2834 -2002
rect 358 -2360 925 -2339
rect 925 -2360 959 -2339
rect 959 -2360 2183 -2339
rect 2183 -2360 2217 -2339
rect 2217 -2360 2778 -2339
rect 358 -2398 2778 -2360
rect 358 -2432 925 -2398
rect 925 -2432 959 -2398
rect 959 -2432 2183 -2398
rect 2183 -2432 2217 -2398
rect 2217 -2432 2778 -2398
rect 358 -2470 2778 -2432
rect 358 -2504 925 -2470
rect 925 -2504 959 -2470
rect 959 -2504 2183 -2470
rect 2183 -2504 2217 -2470
rect 2217 -2504 2778 -2470
rect 358 -2542 2778 -2504
rect 358 -2576 925 -2542
rect 925 -2576 959 -2542
rect 959 -2576 2183 -2542
rect 2183 -2576 2217 -2542
rect 2217 -2576 2778 -2542
rect 358 -2583 2778 -2576
<< metal2 >>
rect -3216 1882 -348 1894
rect -3216 1856 -3210 1882
rect -354 1856 -348 1882
rect 1056 1882 2676 1894
rect 1056 1856 1078 1882
rect 2654 1856 2676 1882
rect -348 1612 -112 1650
rect -3216 1586 -3210 1612
rect -354 1586 -112 1612
rect -3216 1574 -112 1586
rect 1056 1612 1072 1856
rect 2660 1612 2676 1856
rect 1056 1586 1078 1612
rect 2654 1586 2676 1612
rect 1056 1574 2676 1586
rect -2214 714 -2154 720
rect -1184 714 -1124 720
rect -292 714 -232 720
rect -2214 710 -232 714
rect -2214 658 -2210 710
rect -2158 658 -1180 710
rect -1128 658 -288 710
rect -236 658 -232 710
rect -2214 654 -232 658
rect -2214 648 -2154 654
rect -1184 648 -1124 654
rect -292 648 -232 654
rect -3098 596 -3038 602
rect -2344 596 -2284 602
rect -2086 596 -2026 602
rect -1312 596 -1252 602
rect -1052 596 -992 602
rect -3098 592 -992 596
rect -3098 540 -3094 592
rect -3042 540 -2340 592
rect -2288 540 -2082 592
rect -2030 540 -1308 592
rect -1256 540 -1048 592
rect -996 540 -992 592
rect -3098 536 -992 540
rect -3098 530 -3038 536
rect -2344 530 -2284 536
rect -2086 530 -2026 536
rect -1312 530 -1252 536
rect -1052 530 -992 536
rect -474 596 -414 602
rect -172 596 -112 1574
rect 840 1304 900 1310
rect 1226 1304 1286 1310
rect 1484 1304 1544 1310
rect 1868 1304 1928 1310
rect 2508 1304 2568 1310
rect 840 1300 2568 1304
rect 840 1248 844 1300
rect 896 1248 1230 1300
rect 1282 1248 1488 1300
rect 1540 1248 1872 1300
rect 1924 1248 2512 1300
rect 2564 1248 2568 1300
rect 840 1244 2568 1248
rect 840 1238 900 1244
rect 1226 1238 1286 1244
rect 1484 1238 1544 1244
rect 1868 1238 1928 1244
rect 2508 1238 2568 1244
rect -474 592 -112 596
rect -474 540 -470 592
rect -418 540 -112 592
rect -474 536 -112 540
rect -474 530 -414 536
rect 1996 494 2056 500
rect 1987 492 2065 494
rect 1987 436 1998 492
rect 2054 436 2065 492
rect 1987 434 2065 436
rect 254 426 314 432
rect 840 426 900 432
rect 964 426 1024 432
rect 1226 426 1286 432
rect 1354 426 1414 432
rect 1480 426 1540 432
rect 1738 426 1798 432
rect 1868 426 1928 432
rect 1996 428 2056 434
rect 254 422 1928 426
rect 254 370 258 422
rect 310 370 844 422
rect 896 370 968 422
rect 1020 370 1230 422
rect 1282 370 1358 422
rect 1410 370 1484 422
rect 1536 370 1742 422
rect 1794 370 1872 422
rect 1924 370 1928 422
rect 254 366 1928 370
rect 254 360 314 366
rect 840 360 900 366
rect 964 360 1024 366
rect 1226 360 1286 366
rect 1354 360 1414 366
rect 1480 360 1540 366
rect 1738 360 1798 366
rect 1868 360 1928 366
rect -2600 -136 -2540 -130
rect -2346 -136 -2286 -130
rect -2086 -136 -2026 -130
rect -1828 -136 -1768 -130
rect -1570 -136 -1510 -130
rect -1312 -136 -1252 -130
rect -1054 -136 -994 -130
rect -796 -136 -736 -130
rect -2600 -140 -736 -136
rect -2600 -192 -2596 -140
rect -2544 -192 -2342 -140
rect -2290 -192 -2082 -140
rect -2030 -192 -1824 -140
rect -1772 -192 -1566 -140
rect -1514 -192 -1308 -140
rect -1256 -192 -1050 -140
rect -998 -192 -792 -140
rect -740 -192 -736 -140
rect -2600 -196 -736 -192
rect -2600 -202 -2540 -196
rect -2346 -202 -2286 -196
rect -2086 -202 -2026 -196
rect -1828 -202 -1768 -196
rect -1570 -202 -1510 -196
rect -1312 -202 -1252 -196
rect -1054 -202 -994 -196
rect -796 -202 -736 -196
rect -2730 -256 -2670 -250
rect -2216 -256 -2156 -250
rect -1700 -256 -1640 -250
rect -1184 -256 -1124 -250
rect -672 -256 -612 -250
rect 108 -256 168 -250
rect -2730 -260 168 -256
rect -2730 -312 -2726 -260
rect -2674 -312 -2212 -260
rect -2160 -312 -1696 -260
rect -1644 -312 -1180 -260
rect -1128 -312 -668 -260
rect -616 -312 112 -260
rect 164 -312 168 -260
rect -2730 -316 168 -312
rect -2730 -322 -2670 -316
rect -2216 -322 -2156 -316
rect -1700 -322 -1640 -316
rect -1184 -322 -1124 -316
rect -672 -322 -612 -316
rect 108 -322 168 -316
rect 960 -328 1020 -322
rect 1350 -328 1410 -322
rect 1738 -328 1798 -322
rect 2508 -328 2568 -322
rect 960 -332 2838 -328
rect 960 -384 964 -332
rect 1016 -384 1354 -332
rect 1406 -384 1742 -332
rect 1794 -384 2512 -332
rect 2564 -384 2838 -332
rect 960 -388 2838 -384
rect 960 -394 1020 -388
rect 1350 -394 1410 -388
rect 1738 -394 1798 -388
rect 2508 -394 2568 -388
rect 1484 -570 2616 -510
rect 1484 -904 1544 -570
rect 1658 -904 1718 -898
rect 1484 -908 1718 -904
rect 1484 -960 1662 -908
rect 1714 -960 1718 -908
rect 1484 -964 1718 -960
rect -3098 -992 -3038 -986
rect -2604 -992 -2544 -986
rect -1828 -992 -1768 -986
rect -1572 -992 -1512 -986
rect -800 -992 -740 -986
rect -3098 -996 -740 -992
rect -3098 -1048 -3094 -996
rect -3042 -1048 -2600 -996
rect -2548 -1048 -1824 -996
rect -1772 -1048 -1568 -996
rect -1516 -1048 -796 -996
rect -744 -1048 -740 -996
rect -3098 -1052 -740 -1048
rect -3098 -1058 -3038 -1052
rect -2604 -1058 -2544 -1052
rect -1828 -1058 -1768 -1052
rect -1572 -1058 -1512 -1052
rect -800 -1058 -740 -1052
rect 1378 -1014 1438 -1008
rect 1484 -1014 1544 -964
rect 1658 -970 1718 -964
rect 2556 -962 2616 -570
rect 2778 -624 2838 -388
rect 2778 -676 2782 -624
rect 2834 -676 2838 -624
rect 2778 -686 2838 -676
rect 1378 -1018 1544 -1014
rect 1378 -1070 1382 -1018
rect 1434 -1070 1544 -1018
rect 2556 -1022 2844 -962
rect 1378 -1074 1544 -1070
rect 1378 -1080 1438 -1074
rect -2732 -1108 -2672 -1102
rect -2732 -1112 586 -1108
rect -2732 -1164 -2728 -1112
rect -2676 -1114 586 -1112
rect -2676 -1164 -1696 -1114
rect -2732 -1166 -1696 -1164
rect -1644 -1166 -666 -1114
rect -614 -1166 -288 -1114
rect -236 -1166 586 -1114
rect -2732 -1168 586 -1166
rect -2732 -1174 -2672 -1168
rect -1706 -1170 -1634 -1168
rect -1564 -1402 -1504 -1168
rect -676 -1170 -604 -1168
rect -298 -1170 -226 -1168
rect 526 -1208 586 -1168
rect 526 -1268 1018 -1208
rect -1564 -1454 -1560 -1402
rect -1508 -1454 -1504 -1402
rect -1564 -1464 -1504 -1454
rect -1278 -1506 -1218 -1500
rect -183 -1501 -113 -1495
rect -1287 -1514 -1209 -1506
rect -1287 -1570 -1276 -1514
rect -1220 -1570 -1209 -1514
rect -1287 -1578 -1209 -1570
rect -192 -1514 -104 -1501
rect -192 -1570 -176 -1514
rect -120 -1570 -104 -1514
rect -1278 -1584 -1218 -1578
rect -192 -1583 -104 -1570
rect 958 -1532 1018 -1268
rect 958 -1536 1196 -1532
rect -183 -1589 -113 -1583
rect 958 -1588 1134 -1536
rect 1186 -1588 1196 -1536
rect 958 -1592 1196 -1588
rect 564 -1607 664 -1596
rect 560 -1624 668 -1607
rect 560 -1680 586 -1624
rect 642 -1680 668 -1624
rect 560 -1697 668 -1680
rect 564 -1708 664 -1697
rect -632 -1750 -572 -1740
rect -890 -1760 -830 -1750
rect -1146 -1770 -1086 -1760
rect -1146 -1822 -1142 -1770
rect -1090 -1822 -1086 -1770
rect -1146 -2082 -1086 -1822
rect -1146 -2134 -1142 -2082
rect -1090 -2134 -1086 -2082
rect -1146 -2144 -1086 -2134
rect -890 -1812 -886 -1760
rect -834 -1812 -830 -1760
rect -890 -2080 -830 -1812
rect -890 -2132 -886 -2080
rect -834 -2132 -830 -2080
rect -890 -2142 -830 -2132
rect -632 -1802 -628 -1750
rect -576 -1802 -572 -1750
rect -632 -2080 -572 -1802
rect -380 -1752 -320 -1742
rect -380 -1804 -376 -1752
rect -324 -1804 -320 -1752
rect -380 -2076 -320 -1804
rect -246 -1750 -186 -1740
rect -246 -1802 -242 -1750
rect -190 -1802 -186 -1750
rect -632 -2132 -628 -2080
rect -576 -2132 -572 -2080
rect -632 -2142 -572 -2132
rect -386 -2080 -314 -2076
rect -386 -2132 -376 -2080
rect -324 -2132 -314 -2080
rect -386 -2136 -314 -2132
rect -246 -2098 -186 -1802
rect 254 -1988 314 -1982
rect 526 -1988 586 -1982
rect 642 -1988 702 -1982
rect 958 -1988 1018 -1592
rect 2468 -1609 2568 -1598
rect 2464 -1626 2572 -1609
rect 2464 -1682 2490 -1626
rect 2546 -1682 2572 -1626
rect 2464 -1699 2572 -1682
rect 2468 -1710 2568 -1699
rect 1434 -1902 1726 -1898
rect 1434 -1954 1444 -1902
rect 1496 -1954 1664 -1902
rect 1716 -1954 1726 -1902
rect 1434 -1958 1726 -1954
rect 254 -1992 586 -1988
rect 254 -2044 258 -1992
rect 310 -2044 530 -1992
rect 582 -2044 586 -1992
rect 254 -2048 586 -2044
rect 636 -1992 1018 -1988
rect 636 -2044 646 -1992
rect 698 -2044 1018 -1992
rect 636 -2048 1018 -2044
rect 254 -2054 314 -2048
rect 526 -2054 586 -2048
rect 642 -2054 702 -2048
rect 102 -2098 174 -2096
rect 1188 -2098 1248 -2092
rect 1542 -2098 1602 -1958
rect 2546 -1998 2606 -1992
rect 2778 -1998 2838 -1992
rect 2546 -2002 2838 -1998
rect 2546 -2054 2550 -2002
rect 2602 -2054 2782 -2002
rect 2834 -2054 2838 -2002
rect 2546 -2058 2838 -2054
rect 2546 -2064 2606 -2058
rect 2778 -2064 2838 -2058
rect 1896 -2098 1956 -2092
rect 2426 -2098 2486 -2092
rect -246 -2100 2486 -2098
rect -246 -2152 112 -2100
rect 164 -2102 2486 -2100
rect 164 -2152 1192 -2102
rect -246 -2154 1192 -2152
rect 1244 -2154 1900 -2102
rect 1952 -2154 2430 -2102
rect 2482 -2154 2486 -2102
rect -246 -2158 2486 -2154
rect 1188 -2164 1248 -2158
rect 2426 -2164 2486 -2158
rect 346 -2313 2790 -2298
rect 346 -2339 380 -2313
rect 2756 -2339 2790 -2313
rect 346 -2583 358 -2339
rect 2778 -2583 2790 -2339
rect 346 -2609 380 -2583
rect 2756 -2609 2790 -2583
rect 346 -2624 2790 -2609
<< via2 >>
rect -3210 1856 -354 1882
rect -3210 1612 -354 1856
rect 1078 1856 2654 1882
rect -3210 1586 -354 1612
rect 1078 1612 2654 1856
rect 1078 1586 2654 1612
rect 1998 490 2054 492
rect 1998 438 2000 490
rect 2000 438 2052 490
rect 2052 438 2054 490
rect 1998 436 2054 438
rect -1276 -1516 -1220 -1514
rect -1276 -1568 -1274 -1516
rect -1274 -1568 -1222 -1516
rect -1222 -1568 -1220 -1516
rect -1276 -1570 -1220 -1568
rect -176 -1516 -120 -1514
rect -176 -1568 -174 -1516
rect -174 -1568 -122 -1516
rect -122 -1568 -120 -1516
rect -176 -1570 -120 -1568
rect 586 -1626 642 -1624
rect 586 -1678 588 -1626
rect 588 -1678 640 -1626
rect 640 -1678 642 -1626
rect 586 -1680 642 -1678
rect 2490 -1628 2546 -1626
rect 2490 -1680 2492 -1628
rect 2492 -1680 2544 -1628
rect 2544 -1680 2546 -1628
rect 2490 -1682 2546 -1680
rect 380 -2339 2756 -2313
rect 380 -2583 2756 -2339
rect 380 -2609 2756 -2583
<< metal3 >>
rect -3226 1882 -338 1889
rect -3226 1846 -3210 1882
rect -354 1846 -338 1882
rect -3226 1622 -3214 1846
rect -350 1622 -338 1846
rect -3226 1586 -3210 1622
rect -354 1586 -338 1622
rect -3226 1579 -338 1586
rect 1046 1882 2686 1889
rect 1046 1846 1078 1882
rect 2654 1846 2686 1882
rect 1046 1622 1074 1846
rect 2658 1622 2686 1846
rect 1046 1586 1078 1622
rect 2654 1586 2686 1622
rect 1046 1579 2686 1586
rect 1978 496 2078 516
rect 1978 432 1997 496
rect 2061 432 2078 496
rect 1978 416 2078 432
rect 2946 -1256 3046 -1232
rect 2946 -1320 2964 -1256
rect 3028 -1320 3046 -1256
rect -2188 -1508 -2076 -1490
rect -2188 -1572 -2164 -1508
rect -2100 -1572 -2076 -1508
rect -2188 -1590 -2076 -1572
rect -1298 -1510 -1196 -1492
rect -1298 -1574 -1283 -1510
rect -1219 -1574 -1196 -1510
rect -2182 -2858 -2082 -1590
rect -1298 -1592 -1196 -1574
rect -202 -1510 -96 -1488
rect -202 -1514 -175 -1510
rect -202 -1570 -176 -1514
rect -202 -1574 -175 -1570
rect -111 -1574 -96 -1510
rect -202 -1596 -96 -1574
rect 564 -1603 664 -1602
rect 559 -1620 669 -1603
rect 2468 -1605 2568 -1604
rect 559 -1684 582 -1620
rect 646 -1684 669 -1620
rect 559 -1701 669 -1684
rect 2463 -1622 2573 -1605
rect 2463 -1686 2486 -1622
rect 2550 -1686 2573 -1622
rect 564 -1702 664 -1701
rect 2463 -1703 2573 -1686
rect 2468 -1704 2568 -1703
rect 336 -2309 2800 -2303
rect 336 -2613 376 -2309
rect 2760 -2613 2800 -2309
rect 336 -2619 2800 -2613
rect 2946 -2858 3046 -1320
rect -2182 -2958 3046 -2858
<< via3 >>
rect -3214 1622 -3210 1846
rect -3210 1622 -354 1846
rect -354 1622 -350 1846
rect 1074 1622 1078 1846
rect 1078 1622 2654 1846
rect 2654 1622 2658 1846
rect 1997 492 2061 496
rect 1997 436 1998 492
rect 1998 436 2054 492
rect 2054 436 2061 492
rect 1997 432 2061 436
rect 2964 -1320 3028 -1256
rect -2164 -1572 -2100 -1508
rect -1283 -1514 -1219 -1510
rect -1283 -1570 -1276 -1514
rect -1276 -1570 -1220 -1514
rect -1220 -1570 -1219 -1514
rect -1283 -1574 -1219 -1570
rect -175 -1514 -111 -1510
rect -175 -1570 -120 -1514
rect -120 -1570 -111 -1514
rect -175 -1574 -111 -1570
rect 582 -1624 646 -1620
rect 582 -1680 586 -1624
rect 586 -1680 642 -1624
rect 642 -1680 646 -1624
rect 582 -1684 646 -1680
rect 2486 -1626 2550 -1622
rect 2486 -1682 2490 -1626
rect 2490 -1682 2546 -1626
rect 2546 -1682 2550 -1626
rect 2486 -1686 2550 -1682
rect 376 -2313 2760 -2309
rect 376 -2609 380 -2313
rect 380 -2609 2756 -2313
rect 2756 -2609 2760 -2313
rect 376 -2613 2760 -2609
<< metal4 >>
rect -3400 1846 2890 2278
rect -3400 1622 -3214 1846
rect -350 1622 1074 1846
rect 2658 1622 2890 1846
rect -3400 1478 2890 1622
rect 1976 496 3044 516
rect 1976 432 1997 496
rect 2061 432 3044 496
rect 1976 416 3044 432
rect 2944 -1237 3044 416
rect 2944 -1244 3047 -1237
rect 2468 -1256 3047 -1244
rect 2468 -1320 2964 -1256
rect 3028 -1320 3047 -1256
rect 2468 -1339 3047 -1320
rect 2468 -1344 3044 -1339
rect -2183 -1492 -2081 -1489
rect -2190 -1508 668 -1492
rect -2190 -1572 -2164 -1508
rect -2100 -1510 668 -1508
rect -2100 -1572 -1283 -1510
rect -2190 -1574 -1283 -1572
rect -1219 -1574 -175 -1510
rect -111 -1574 668 -1510
rect -2190 -1592 668 -1574
rect 564 -1620 668 -1592
rect 564 -1684 582 -1620
rect 646 -1684 668 -1620
rect 564 -1702 668 -1684
rect 568 -1706 668 -1702
rect 2468 -1622 2568 -1344
rect 2468 -1686 2486 -1622
rect 2550 -1686 2568 -1622
rect 2468 -1704 2568 -1686
rect -3400 -2309 2890 -2214
rect -3400 -2613 376 -2309
rect 2760 -2613 2890 -2309
rect -3400 -3014 2890 -2613
use sky130_fd_pr__pfet_01v8_RCENQY  sky130_fd_pr__pfet_01v8_RCENQY_0
timestamp 1626486988
transform 1 0 -1645 0 1 1190
box -1439 -200 1439 200
use sky130_fd_pr__pfet_01v8_9JKHSP  sky130_fd_pr__pfet_01v8_9JKHSP_1
timestamp 1626486988
transform 1 0 1512 0 1 30
box -968 -300 968 300
use sky130_fd_pr__pfet_01v8_9JKHSP  sky130_fd_pr__pfet_01v8_9JKHSP_0
timestamp 1626486988
transform 1 0 1512 0 1 890
box -968 -300 968 300
use sky130_fd_pr__pfet_01v8_lvt_JN5RQF  sky130_fd_pr__pfet_01v8_lvt_JN5RQF_1
timestamp 1626486988
transform 1 0 -1670 0 1 -653
box -1355 -300 1355 300
use sky130_fd_pr__pfet_01v8_lvt_JN5RQF  sky130_fd_pr__pfet_01v8_lvt_JN5RQF_0
timestamp 1626486988
transform 1 0 -1670 0 1 207
box -1355 -300 1355 300
use sky130_fd_pr__nfet_01v8_BGQ2FN  sky130_fd_pr__nfet_01v8_BGQ2FN_1
timestamp 1626486988
transform 1 0 614 0 1 -1801
box -216 -269 216 269
use sky130_fd_pr__nfet_01v8_BGQ2FN  sky130_fd_pr__nfet_01v8_BGQ2FN_0
timestamp 1626486988
transform 1 0 2518 0 1 -1801
box -216 -269 216 269
use sky130_fd_pr__nfet_01v8_7DDHNL  sky130_fd_pr__nfet_01v8_7DDHNL_0
timestamp 1626486988
transform 1 0 1573 0 1 -1746
box -527 -126 527 126
use sky130_fd_pr__pfet_01v8_lvt_XJHVCG  sky130_fd_pr__pfet_01v8_lvt_XJHVCG_0
timestamp 1626486988
transform 1 0 -667 0 1 -1724
box -743 -342 743 344
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_0
timestamp 1626486988
transform 1 0 1178 0 1 -1166
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_1
timestamp 1626486988
transform -1 0 1916 0 1 -1166
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0
timestamp 1626486988
transform 1 0 626 0 1 -1166
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_1
timestamp 1626486988
transform 1 0 902 0 1 -1166
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_2
timestamp 1626486988
transform -1 0 2192 0 1 -1166
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_3
timestamp 1626486988
transform -1 0 2468 0 1 -1166
box -38 -48 314 592
<< labels >>
flabel metal4 s 324 2134 340 2140 1 FreeSans 600 0 0 0 VDD
flabel metal1 s -3086 -112 -3072 -100 1 FreeSans 600 0 0 0 vip
flabel metal1 s -2316 -232 -2306 -222 1 FreeSans 600 0 0 0 vim
flabel metal1 s -276 278 -262 298 1 FreeSans 600 0 0 0 vlatchm
flabel metal1 s -2710 -188 -2696 -178 1 FreeSans 600 0 0 0 vlatchp
flabel metal1 s -1664 800 -1646 814 1 FreeSans 600 0 0 0 vtailp
flabel metal1 s -1746 918 -1726 930 1 FreeSans 600 0 0 0 ibiasp
flabel metal2 s 862 368 878 384 1 FreeSans 600 0 0 0 vcompm
flabel metal1 s 2526 590 2546 614 1 FreeSans 600 0 0 0 vcompp
flabel metal4 s -186 -2534 -160 -2514 1 FreeSans 600 0 0 0 VSS
flabel metal1 s 1360 -1568 1366 -1562 1 FreeSans 600 0 0 0 vlatchm
flabel metal2 s 1448 -2134 1456 -2126 1 FreeSans 600 0 0 0 vlatchp
flabel metal1 s 1156 -934 1162 -928 1 FreeSans 200 0 0 0 vcompm_buf
flabel metal1 s 900 -934 906 -930 1 FreeSans 200 0 0 0 vcompmb
flabel metal1 s 1924 -930 1928 -926 1 FreeSans 200 0 0 0 vcompp_buf
flabel metal1 s 2178 -932 2184 -928 1 FreeSans 200 0 0 0 vcomppb
flabel metal2 s 2674 -990 2680 -984 1 FreeSans 600 0 0 0 vop
flabel metal1 s 1606 -1052 1612 -1044 1 FreeSans 600 0 0 0 vom
flabel metal4 s -1548 -1552 -1528 -1534 1 FreeSans 600 0 0 0 clk
<< properties >>
string FIXED_BBOX 308 88 2612 2032
<< end >>
