**.subckt inv4_stdcell VDD VSS A Y
*.ipin VDD
*.ipin VSS
*.ipin A
*.opin Y
x1 A VSS VSS VDD VDD Y sky130_fd_sc_hd__inv_4
**** begin user architecture code

.include ~/skywater-pdk/libraries/sky130_fd_sc_hd/latest/cells/inv/sky130_fd_sc_hd__inv_4.spice

**** end user architecture code
**.ends
** flattened .save nodes
.end
