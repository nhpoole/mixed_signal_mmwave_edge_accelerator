magic
tech sky130A
magscale 1 2
timestamp 1622096065
<< nwell >>
rect -194 -300 194 300
<< pmoslvt >>
rect -100 -200 100 200
<< pdiff >>
rect -158 188 -100 200
rect -158 -188 -146 188
rect -112 -188 -100 188
rect -158 -200 -100 -188
rect 100 188 158 200
rect 100 -188 112 188
rect 146 -188 158 188
rect 100 -200 158 -188
<< pdiffc >>
rect -146 -188 -112 188
rect 112 -188 146 188
<< poly >>
rect -66 281 66 297
rect -66 264 -50 281
rect -100 247 -50 264
rect 50 264 66 281
rect 50 247 100 264
rect -100 200 100 247
rect -100 -247 100 -200
rect -100 -264 -50 -247
rect -66 -281 -50 -264
rect 50 -264 100 -247
rect 50 -281 66 -264
rect -66 -297 66 -281
<< polycont >>
rect -50 247 50 281
rect -50 -281 50 -247
<< locali >>
rect -66 247 -50 281
rect 50 247 66 281
rect -146 188 -112 204
rect -146 -204 -112 -188
rect 112 188 146 204
rect 112 -204 146 -188
rect -66 -281 -50 -247
rect 50 -281 66 -247
<< viali >>
rect -42 247 42 281
rect -146 -188 -112 188
rect 112 -188 146 188
rect -42 -281 42 -247
<< metal1 >>
rect -54 281 54 287
rect -54 247 -42 281
rect 42 247 54 281
rect -54 241 54 247
rect -152 188 -106 200
rect -152 -188 -146 188
rect -112 -188 -106 188
rect -152 -200 -106 -188
rect 106 188 152 200
rect 106 -188 112 188
rect 146 -188 152 188
rect 106 -200 152 -188
rect -54 -247 54 -241
rect -54 -281 -42 -247
rect 42 -281 54 -247
rect -54 -287 54 -281
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string parameters w 2 l 1 m 1 nf 1 diffcov 100 polycov 60 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
