magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect -1801 -1260 2197 3516
<< nwell >>
rect -541 264 937 1614
<< pwell >>
rect 158 2135 356 2161
rect 158 1991 494 2135
rect 158 1845 356 1991
rect 70 1663 356 1845
rect 72 201 268 222
rect 72 57 424 201
rect 72 40 268 57
<< nmos >>
rect 242 2005 272 2135
rect 154 1689 184 1819
rect 242 1689 272 1819
rect 156 66 186 196
<< pmos >>
rect 154 1324 184 1576
rect 242 1324 272 1576
rect 154 702 184 1102
rect 346 702 376 1102
rect 156 302 186 554
<< ndiff >>
rect 184 2120 242 2135
rect 184 2086 196 2120
rect 230 2086 242 2120
rect 184 2052 242 2086
rect 184 2018 196 2052
rect 230 2018 242 2052
rect 184 2005 242 2018
rect 272 2122 330 2135
rect 272 2088 284 2122
rect 318 2088 330 2122
rect 272 2054 330 2088
rect 272 2020 284 2054
rect 318 2020 330 2054
rect 272 2005 330 2020
rect 96 1807 154 1819
rect 96 1773 108 1807
rect 142 1773 154 1807
rect 96 1739 154 1773
rect 96 1705 108 1739
rect 142 1705 154 1739
rect 96 1689 154 1705
rect 184 1807 242 1819
rect 184 1773 196 1807
rect 230 1773 242 1807
rect 184 1739 242 1773
rect 184 1705 196 1739
rect 230 1705 242 1739
rect 184 1689 242 1705
rect 272 1807 330 1819
rect 272 1773 284 1807
rect 318 1773 330 1807
rect 272 1739 330 1773
rect 272 1705 284 1739
rect 318 1705 330 1739
rect 272 1689 330 1705
rect 98 182 156 196
rect 98 148 110 182
rect 144 148 156 182
rect 98 114 156 148
rect 98 80 110 114
rect 144 80 156 114
rect 98 66 156 80
rect 186 182 242 196
rect 186 148 198 182
rect 232 148 242 182
rect 186 114 242 148
rect 186 80 198 114
rect 232 80 242 114
rect 186 66 242 80
<< pdiff >>
rect 100 1535 154 1576
rect 100 1501 108 1535
rect 142 1501 154 1535
rect 100 1467 154 1501
rect 100 1433 108 1467
rect 142 1433 154 1467
rect 100 1399 154 1433
rect 100 1365 108 1399
rect 142 1365 154 1399
rect 100 1324 154 1365
rect 184 1535 242 1576
rect 184 1501 196 1535
rect 230 1501 242 1535
rect 184 1467 242 1501
rect 184 1433 196 1467
rect 230 1433 242 1467
rect 184 1399 242 1433
rect 184 1365 196 1399
rect 230 1365 242 1399
rect 184 1324 242 1365
rect 272 1535 326 1576
rect 272 1501 284 1535
rect 318 1501 326 1535
rect 272 1467 326 1501
rect 272 1433 284 1467
rect 318 1433 326 1467
rect 272 1399 326 1433
rect 272 1365 284 1399
rect 318 1365 326 1399
rect 272 1324 326 1365
rect 100 1089 154 1102
rect 100 1055 108 1089
rect 142 1055 154 1089
rect 100 1021 154 1055
rect 100 987 108 1021
rect 142 987 154 1021
rect 100 953 154 987
rect 100 919 108 953
rect 142 919 154 953
rect 100 885 154 919
rect 100 851 108 885
rect 142 851 154 885
rect 100 817 154 851
rect 100 783 108 817
rect 142 783 154 817
rect 100 749 154 783
rect 100 715 108 749
rect 142 715 154 749
rect 100 702 154 715
rect 184 1089 238 1102
rect 184 1055 196 1089
rect 230 1055 238 1089
rect 184 1021 238 1055
rect 184 987 196 1021
rect 230 987 238 1021
rect 184 953 238 987
rect 184 919 196 953
rect 230 919 238 953
rect 184 885 238 919
rect 184 851 196 885
rect 230 851 238 885
rect 184 817 238 851
rect 184 783 196 817
rect 230 783 238 817
rect 184 749 238 783
rect 184 715 196 749
rect 230 715 238 749
rect 184 702 238 715
rect 292 1089 346 1102
rect 292 1055 300 1089
rect 334 1055 346 1089
rect 292 1021 346 1055
rect 292 987 300 1021
rect 334 987 346 1021
rect 292 953 346 987
rect 292 919 300 953
rect 334 919 346 953
rect 292 885 346 919
rect 292 851 300 885
rect 334 851 346 885
rect 292 817 346 851
rect 292 783 300 817
rect 334 783 346 817
rect 292 749 346 783
rect 292 715 300 749
rect 334 715 346 749
rect 292 702 346 715
rect 376 1089 430 1102
rect 376 1055 388 1089
rect 422 1055 430 1089
rect 376 1021 430 1055
rect 376 987 388 1021
rect 422 987 430 1021
rect 376 953 430 987
rect 376 919 388 953
rect 422 919 430 953
rect 376 885 430 919
rect 376 851 388 885
rect 422 851 430 885
rect 376 817 430 851
rect 376 783 388 817
rect 422 783 430 817
rect 376 749 430 783
rect 376 715 388 749
rect 422 715 430 749
rect 376 702 430 715
rect 98 513 156 554
rect 98 479 110 513
rect 144 479 156 513
rect 98 445 156 479
rect 98 411 110 445
rect 144 411 156 445
rect 98 377 156 411
rect 98 343 110 377
rect 144 343 156 377
rect 98 302 156 343
rect 186 513 240 554
rect 186 479 198 513
rect 232 479 240 513
rect 186 445 240 479
rect 186 411 198 445
rect 232 411 240 445
rect 186 377 240 411
rect 186 343 198 377
rect 232 343 240 377
rect 186 302 240 343
<< ndiffc >>
rect 196 2086 230 2120
rect 196 2018 230 2052
rect 284 2088 318 2122
rect 284 2020 318 2054
rect 108 1773 142 1807
rect 108 1705 142 1739
rect 196 1773 230 1807
rect 196 1705 230 1739
rect 284 1773 318 1807
rect 284 1705 318 1739
rect 110 148 144 182
rect 110 80 144 114
rect 198 148 232 182
rect 198 80 232 114
<< pdiffc >>
rect 108 1501 142 1535
rect 108 1433 142 1467
rect 108 1365 142 1399
rect 196 1501 230 1535
rect 196 1433 230 1467
rect 196 1365 230 1399
rect 284 1501 318 1535
rect 284 1433 318 1467
rect 284 1365 318 1399
rect 108 1055 142 1089
rect 108 987 142 1021
rect 108 919 142 953
rect 108 851 142 885
rect 108 783 142 817
rect 108 715 142 749
rect 196 1055 230 1089
rect 196 987 230 1021
rect 196 919 230 953
rect 196 851 230 885
rect 196 783 230 817
rect 196 715 230 749
rect 300 1055 334 1089
rect 300 987 334 1021
rect 300 919 334 953
rect 300 851 334 885
rect 300 783 334 817
rect 300 715 334 749
rect 388 1055 422 1089
rect 388 987 422 1021
rect 388 919 422 953
rect 388 851 422 885
rect 388 783 422 817
rect 388 715 422 749
rect 110 479 144 513
rect 110 411 144 445
rect 110 343 144 377
rect 198 479 232 513
rect 198 411 232 445
rect 198 343 232 377
<< psubdiff >>
rect 434 2085 468 2109
rect 434 2017 468 2051
rect 364 151 398 175
rect 364 83 398 117
<< nsubdiff >>
rect 388 1348 422 1376
rect 388 1290 422 1314
<< psubdiffcont >>
rect 434 2051 468 2085
rect 364 117 398 151
<< nsubdiffcont >>
rect 388 1314 422 1348
<< poly >>
rect 240 2220 274 2226
rect 230 2210 284 2220
rect 230 2176 240 2210
rect 274 2176 284 2210
rect 230 2166 284 2176
rect 240 2160 274 2166
rect 242 2135 272 2160
rect 242 1989 272 2005
rect 26 1959 272 1989
rect 26 1148 56 1959
rect 306 1917 372 1927
rect 154 1887 322 1917
rect 154 1819 184 1887
rect 306 1883 322 1887
rect 356 1883 372 1917
rect 306 1873 372 1883
rect 342 1862 372 1873
rect 242 1819 272 1845
rect 342 1828 376 1862
rect 154 1576 184 1689
rect 242 1576 272 1689
rect 345 1676 375 1828
rect 342 1642 376 1676
rect 154 1298 184 1324
rect 242 1256 272 1324
rect 98 1240 272 1256
rect 98 1206 108 1240
rect 142 1226 272 1240
rect 342 1232 372 1642
rect 142 1206 152 1226
rect 98 1196 152 1206
rect 342 1206 474 1232
rect 342 1202 430 1206
rect 108 1190 142 1196
rect 420 1172 430 1202
rect 464 1172 474 1206
rect 420 1158 474 1172
rect 430 1156 474 1158
rect 26 1118 184 1148
rect 154 1102 184 1118
rect 346 1102 376 1128
rect 154 686 184 702
rect 346 686 376 702
rect 154 656 376 686
rect 156 598 432 614
rect 156 584 388 598
rect 156 554 186 584
rect 378 564 388 584
rect 422 564 432 598
rect 378 548 432 564
rect 156 196 186 302
rect 156 36 186 66
<< polycont >>
rect 240 2176 274 2210
rect 322 1883 356 1917
rect 108 1206 142 1240
rect 430 1172 464 1206
rect 388 564 422 598
<< locali >>
rect 106 2211 140 2212
rect 140 2177 240 2210
rect 106 2176 240 2177
rect 274 2176 290 2210
rect 196 2120 230 2142
rect 196 2052 230 2086
rect 108 1807 142 1830
rect 108 1739 142 1773
rect 108 1535 142 1705
rect 196 1807 230 2018
rect 284 2122 318 2142
rect 284 2085 318 2088
rect 434 2085 468 2101
rect 284 2054 434 2085
rect 318 2051 434 2054
rect 284 2001 318 2020
rect 196 1739 230 1773
rect 196 1685 230 1705
rect 284 1883 322 1917
rect 356 1883 374 1917
rect 284 1807 318 1883
rect 284 1739 318 1773
rect 108 1467 142 1501
rect 108 1399 142 1433
rect 108 1240 142 1365
rect 196 1535 230 1580
rect 196 1467 230 1501
rect 196 1399 230 1433
rect 196 1286 230 1365
rect 284 1535 318 1705
rect 284 1467 318 1501
rect 284 1399 318 1433
rect 284 1320 318 1365
rect 352 1314 388 1348
rect 422 1314 438 1348
rect 352 1286 386 1314
rect 196 1252 352 1286
rect 108 1089 142 1206
rect 420 1206 474 1222
rect 420 1190 430 1206
rect 388 1172 430 1190
rect 464 1172 474 1206
rect 388 1156 474 1172
rect 108 1021 142 1055
rect 108 953 142 987
rect 108 885 142 919
rect 108 817 142 851
rect 108 749 142 783
rect 108 656 142 715
rect 196 1089 230 1090
rect 196 1021 230 1055
rect 196 953 230 987
rect 196 885 230 919
rect 196 817 230 851
rect 196 749 230 783
rect 196 694 230 715
rect 300 1089 334 1096
rect 300 1021 334 1055
rect 300 953 334 987
rect 300 885 334 919
rect 300 817 334 851
rect 300 749 334 783
rect 300 698 334 715
rect 388 1089 422 1156
rect 388 1021 422 1055
rect 388 953 422 987
rect 388 885 422 919
rect 388 817 422 851
rect 388 749 422 783
rect 388 598 422 715
rect 110 513 144 558
rect 110 445 144 479
rect 110 377 144 411
rect 110 242 144 343
rect 198 513 232 558
rect 388 548 422 564
rect 198 446 232 479
rect 198 445 364 446
rect 232 412 364 445
rect 198 377 232 411
rect 198 298 232 343
rect 110 182 144 208
rect 110 114 144 148
rect 110 60 144 80
rect 196 182 232 200
rect 196 148 198 182
rect 364 152 398 167
rect 232 151 398 152
rect 232 148 364 151
rect 196 116 364 148
rect 196 114 232 116
rect 196 80 198 114
rect 196 60 232 80
<< viali >>
rect 106 2177 140 2211
rect 434 2017 468 2051
rect 352 1252 386 1286
rect 196 1090 230 1124
rect 300 1096 334 1130
rect 364 412 398 446
rect 110 208 144 242
rect 364 83 398 117
<< metal1 >>
rect 94 2211 152 2224
rect 94 2177 106 2211
rect 140 2177 152 2211
rect 94 2164 152 2177
rect 196 1130 230 2256
rect 272 1142 300 2256
rect 428 2051 474 2079
rect 428 2017 434 2051
rect 468 2017 474 2051
rect 428 2005 474 2017
rect 338 1286 400 1302
rect 338 1252 352 1286
rect 386 1252 400 1286
rect 338 1234 400 1252
rect 272 1130 340 1142
rect 184 1124 242 1130
rect 184 1090 196 1124
rect 230 1090 242 1124
rect 184 1084 242 1090
rect 272 1096 300 1130
rect 334 1096 340 1130
rect 272 1084 340 1096
rect 104 242 150 254
rect 104 208 110 242
rect 144 208 150 242
rect 104 0 150 208
rect 196 0 230 1084
rect 272 0 300 1084
rect 358 446 404 468
rect 358 412 364 446
rect 398 412 404 446
rect 358 392 404 412
rect 358 117 404 145
rect 358 83 364 117
rect 398 83 404 117
rect 358 71 404 83
<< labels >>
rlabel metal1 s 196 1130 230 2256 4 BL
rlabel metal1 s 272 1142 300 2256 4 BR
rlabel metal1 s 104 0 150 254 4 DOUT
rlabel metal1 s 94 2164 152 2224 4 EN
rlabel metal1 s 428 2005 474 2079 4 GND
rlabel metal1 s 358 71 404 145 4 GND
rlabel metal1 s 338 1234 400 1302 4 VDD
rlabel metal1 s 358 392 404 468 4 VDD
rlabel metal1 s 213 1693 213 1693 4 bl
rlabel metal1 s 286 1699 286 1699 4 br
rlabel metal1 s 127 127 127 127 4 dout
rlabel metal1 s 123 2194 123 2194 4 en
rlabel metal1 s 369 1268 369 1268 4 vdd
rlabel metal1 s 381 430 381 430 4 vdd
rlabel metal1 s 451 2042 451 2042 4 gnd
rlabel metal1 s 381 108 381 108 4 gnd
<< properties >>
string FIXED_BBOX 0 0 500 2256
<< end >>
