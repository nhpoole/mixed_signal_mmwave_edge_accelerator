magic
tech sky130A
magscale 1 2
timestamp 1621559963
<< nwell >>
rect -3358 582 3358 3158
<< pwell >>
rect -3358 -3558 3358 418
<< nmos >>
rect 400 -584 600 -384
rect 658 -584 858 -384
rect 916 -584 1116 -384
rect 1174 -584 1374 -384
rect 1432 -584 1632 -384
rect 1690 -584 1890 -384
rect 2362 -758 2562 -358
rect -2517 -1815 -1717 -1615
rect -1659 -1815 -859 -1615
rect -801 -1815 -1 -1615
rect 57 -1815 857 -1615
rect 915 -1815 1715 -1615
rect 1773 -1815 2573 -1615
rect -2517 -2233 -1717 -2033
rect -1659 -2233 -859 -2033
rect -801 -2233 -1 -2033
rect 57 -2233 857 -2033
rect 915 -2233 1715 -2033
rect 1773 -2233 2573 -2033
<< pmos >>
rect -2597 1813 -2397 2013
rect -2339 1813 -2139 2013
rect -2081 1813 -1881 2013
rect -1823 1813 -1623 2013
rect -1565 1813 -1365 2013
rect -1307 1813 -1107 2013
rect -1049 1813 -849 2013
rect -791 1813 -591 2013
rect -533 1813 -333 2013
rect -275 1813 -75 2013
rect 402 1812 602 2012
rect 660 1812 860 2012
rect 918 1812 1118 2012
rect 1176 1812 1376 2012
rect 1434 1812 1634 2012
rect 1692 1812 1892 2012
rect -2597 1139 -2397 1339
rect -2339 1139 -2139 1339
rect -2081 1139 -1881 1339
rect -1823 1139 -1623 1339
rect -1565 1139 -1365 1339
rect -1307 1139 -1107 1339
rect -1049 1139 -849 1339
rect -791 1139 -591 1339
rect -533 1139 -333 1339
rect -275 1139 -75 1339
rect 402 1138 602 1338
rect 660 1138 860 1338
rect 918 1138 1118 1338
rect 1176 1138 1376 1338
rect 1434 1138 1634 1338
rect 1692 1138 1892 1338
<< pmoshvt >>
rect 2362 1138 2562 1938
<< nmoslvt >>
rect -2818 -622 -2618 -422
rect -2560 -622 -2360 -422
rect -2302 -622 -2102 -422
rect -2044 -622 -1844 -422
rect -1786 -622 -1586 -422
rect -1528 -622 -1328 -422
rect -1270 -622 -1070 -422
rect -1012 -622 -812 -422
rect -754 -622 -554 -422
rect -496 -622 -296 -422
<< ndiff >>
rect -2876 -434 -2818 -422
rect -2876 -610 -2864 -434
rect -2830 -610 -2818 -434
rect -2876 -622 -2818 -610
rect -2618 -434 -2560 -422
rect -2618 -610 -2606 -434
rect -2572 -610 -2560 -434
rect -2618 -622 -2560 -610
rect -2360 -434 -2302 -422
rect -2360 -610 -2348 -434
rect -2314 -610 -2302 -434
rect -2360 -622 -2302 -610
rect -2102 -434 -2044 -422
rect -2102 -610 -2090 -434
rect -2056 -610 -2044 -434
rect -2102 -622 -2044 -610
rect -1844 -434 -1786 -422
rect -1844 -610 -1832 -434
rect -1798 -610 -1786 -434
rect -1844 -622 -1786 -610
rect -1586 -434 -1528 -422
rect -1586 -610 -1574 -434
rect -1540 -610 -1528 -434
rect -1586 -622 -1528 -610
rect -1328 -434 -1270 -422
rect -1328 -610 -1316 -434
rect -1282 -610 -1270 -434
rect -1328 -622 -1270 -610
rect -1070 -434 -1012 -422
rect -1070 -610 -1058 -434
rect -1024 -610 -1012 -434
rect -1070 -622 -1012 -610
rect -812 -434 -754 -422
rect -812 -610 -800 -434
rect -766 -610 -754 -434
rect -812 -622 -754 -610
rect -554 -434 -496 -422
rect -554 -610 -542 -434
rect -508 -610 -496 -434
rect -554 -622 -496 -610
rect -296 -434 -238 -422
rect -296 -610 -284 -434
rect -250 -610 -238 -434
rect -296 -622 -238 -610
rect 2304 -370 2362 -358
rect 342 -396 400 -384
rect 342 -572 354 -396
rect 388 -572 400 -396
rect 342 -584 400 -572
rect 600 -396 658 -384
rect 600 -572 612 -396
rect 646 -572 658 -396
rect 600 -584 658 -572
rect 858 -396 916 -384
rect 858 -572 870 -396
rect 904 -572 916 -396
rect 858 -584 916 -572
rect 1116 -396 1174 -384
rect 1116 -572 1128 -396
rect 1162 -572 1174 -396
rect 1116 -584 1174 -572
rect 1374 -396 1432 -384
rect 1374 -572 1386 -396
rect 1420 -572 1432 -396
rect 1374 -584 1432 -572
rect 1632 -396 1690 -384
rect 1632 -572 1644 -396
rect 1678 -572 1690 -396
rect 1632 -584 1690 -572
rect 1890 -396 1948 -384
rect 1890 -572 1902 -396
rect 1936 -572 1948 -396
rect 1890 -584 1948 -572
rect 2304 -746 2316 -370
rect 2350 -746 2362 -370
rect 2304 -758 2362 -746
rect 2562 -370 2620 -358
rect 2562 -746 2574 -370
rect 2608 -746 2620 -370
rect 2562 -758 2620 -746
rect -2575 -1627 -2517 -1615
rect -2575 -1803 -2563 -1627
rect -2529 -1803 -2517 -1627
rect -2575 -1815 -2517 -1803
rect -1717 -1627 -1659 -1615
rect -1717 -1803 -1705 -1627
rect -1671 -1803 -1659 -1627
rect -1717 -1815 -1659 -1803
rect -859 -1627 -801 -1615
rect -859 -1803 -847 -1627
rect -813 -1803 -801 -1627
rect -859 -1815 -801 -1803
rect -1 -1627 57 -1615
rect -1 -1803 11 -1627
rect 45 -1803 57 -1627
rect -1 -1815 57 -1803
rect 857 -1627 915 -1615
rect 857 -1803 869 -1627
rect 903 -1803 915 -1627
rect 857 -1815 915 -1803
rect 1715 -1627 1773 -1615
rect 1715 -1803 1727 -1627
rect 1761 -1803 1773 -1627
rect 1715 -1815 1773 -1803
rect 2573 -1627 2631 -1615
rect 2573 -1803 2585 -1627
rect 2619 -1803 2631 -1627
rect 2573 -1815 2631 -1803
rect -2575 -2045 -2517 -2033
rect -2575 -2221 -2563 -2045
rect -2529 -2221 -2517 -2045
rect -2575 -2233 -2517 -2221
rect -1717 -2045 -1659 -2033
rect -1717 -2221 -1705 -2045
rect -1671 -2221 -1659 -2045
rect -1717 -2233 -1659 -2221
rect -859 -2045 -801 -2033
rect -859 -2221 -847 -2045
rect -813 -2221 -801 -2045
rect -859 -2233 -801 -2221
rect -1 -2045 57 -2033
rect -1 -2221 11 -2045
rect 45 -2221 57 -2045
rect -1 -2233 57 -2221
rect 857 -2045 915 -2033
rect 857 -2221 869 -2045
rect 903 -2221 915 -2045
rect 857 -2233 915 -2221
rect 1715 -2045 1773 -2033
rect 1715 -2221 1727 -2045
rect 1761 -2221 1773 -2045
rect 1715 -2233 1773 -2221
rect 2573 -2045 2631 -2033
rect 2573 -2221 2585 -2045
rect 2619 -2221 2631 -2045
rect 2573 -2233 2631 -2221
<< pdiff >>
rect -2655 2001 -2597 2013
rect -2655 1825 -2643 2001
rect -2609 1825 -2597 2001
rect -2655 1813 -2597 1825
rect -2397 2001 -2339 2013
rect -2397 1825 -2385 2001
rect -2351 1825 -2339 2001
rect -2397 1813 -2339 1825
rect -2139 2001 -2081 2013
rect -2139 1825 -2127 2001
rect -2093 1825 -2081 2001
rect -2139 1813 -2081 1825
rect -1881 2001 -1823 2013
rect -1881 1825 -1869 2001
rect -1835 1825 -1823 2001
rect -1881 1813 -1823 1825
rect -1623 2001 -1565 2013
rect -1623 1825 -1611 2001
rect -1577 1825 -1565 2001
rect -1623 1813 -1565 1825
rect -1365 2001 -1307 2013
rect -1365 1825 -1353 2001
rect -1319 1825 -1307 2001
rect -1365 1813 -1307 1825
rect -1107 2001 -1049 2013
rect -1107 1825 -1095 2001
rect -1061 1825 -1049 2001
rect -1107 1813 -1049 1825
rect -849 2001 -791 2013
rect -849 1825 -837 2001
rect -803 1825 -791 2001
rect -849 1813 -791 1825
rect -591 2001 -533 2013
rect -591 1825 -579 2001
rect -545 1825 -533 2001
rect -591 1813 -533 1825
rect -333 2001 -275 2013
rect -333 1825 -321 2001
rect -287 1825 -275 2001
rect -333 1813 -275 1825
rect -75 2001 -17 2013
rect -75 1825 -63 2001
rect -29 1825 -17 2001
rect -75 1813 -17 1825
rect 344 2000 402 2012
rect 344 1824 356 2000
rect 390 1824 402 2000
rect 344 1812 402 1824
rect 602 2000 660 2012
rect 602 1824 614 2000
rect 648 1824 660 2000
rect 602 1812 660 1824
rect 860 2000 918 2012
rect 860 1824 872 2000
rect 906 1824 918 2000
rect 860 1812 918 1824
rect 1118 2000 1176 2012
rect 1118 1824 1130 2000
rect 1164 1824 1176 2000
rect 1118 1812 1176 1824
rect 1376 2000 1434 2012
rect 1376 1824 1388 2000
rect 1422 1824 1434 2000
rect 1376 1812 1434 1824
rect 1634 2000 1692 2012
rect 1634 1824 1646 2000
rect 1680 1824 1692 2000
rect 1634 1812 1692 1824
rect 1892 2000 1950 2012
rect 1892 1824 1904 2000
rect 1938 1824 1950 2000
rect 1892 1812 1950 1824
rect 2304 1926 2362 1938
rect -2655 1327 -2597 1339
rect -2655 1151 -2643 1327
rect -2609 1151 -2597 1327
rect -2655 1139 -2597 1151
rect -2397 1327 -2339 1339
rect -2397 1151 -2385 1327
rect -2351 1151 -2339 1327
rect -2397 1139 -2339 1151
rect -2139 1327 -2081 1339
rect -2139 1151 -2127 1327
rect -2093 1151 -2081 1327
rect -2139 1139 -2081 1151
rect -1881 1327 -1823 1339
rect -1881 1151 -1869 1327
rect -1835 1151 -1823 1327
rect -1881 1139 -1823 1151
rect -1623 1327 -1565 1339
rect -1623 1151 -1611 1327
rect -1577 1151 -1565 1327
rect -1623 1139 -1565 1151
rect -1365 1327 -1307 1339
rect -1365 1151 -1353 1327
rect -1319 1151 -1307 1327
rect -1365 1139 -1307 1151
rect -1107 1327 -1049 1339
rect -1107 1151 -1095 1327
rect -1061 1151 -1049 1327
rect -1107 1139 -1049 1151
rect -849 1327 -791 1339
rect -849 1151 -837 1327
rect -803 1151 -791 1327
rect -849 1139 -791 1151
rect -591 1327 -533 1339
rect -591 1151 -579 1327
rect -545 1151 -533 1327
rect -591 1139 -533 1151
rect -333 1327 -275 1339
rect -333 1151 -321 1327
rect -287 1151 -275 1327
rect -333 1139 -275 1151
rect -75 1327 -17 1339
rect -75 1151 -63 1327
rect -29 1151 -17 1327
rect -75 1139 -17 1151
rect 344 1326 402 1338
rect 344 1150 356 1326
rect 390 1150 402 1326
rect 344 1138 402 1150
rect 602 1326 660 1338
rect 602 1150 614 1326
rect 648 1150 660 1326
rect 602 1138 660 1150
rect 860 1326 918 1338
rect 860 1150 872 1326
rect 906 1150 918 1326
rect 860 1138 918 1150
rect 1118 1326 1176 1338
rect 1118 1150 1130 1326
rect 1164 1150 1176 1326
rect 1118 1138 1176 1150
rect 1376 1326 1434 1338
rect 1376 1150 1388 1326
rect 1422 1150 1434 1326
rect 1376 1138 1434 1150
rect 1634 1326 1692 1338
rect 1634 1150 1646 1326
rect 1680 1150 1692 1326
rect 1634 1138 1692 1150
rect 1892 1326 1950 1338
rect 1892 1150 1904 1326
rect 1938 1150 1950 1326
rect 1892 1138 1950 1150
rect 2304 1150 2316 1926
rect 2350 1150 2362 1926
rect 2304 1138 2362 1150
rect 2562 1926 2620 1938
rect 2562 1150 2574 1926
rect 2608 1150 2620 1926
rect 2562 1138 2620 1150
<< ndiffc >>
rect -2864 -610 -2830 -434
rect -2606 -610 -2572 -434
rect -2348 -610 -2314 -434
rect -2090 -610 -2056 -434
rect -1832 -610 -1798 -434
rect -1574 -610 -1540 -434
rect -1316 -610 -1282 -434
rect -1058 -610 -1024 -434
rect -800 -610 -766 -434
rect -542 -610 -508 -434
rect -284 -610 -250 -434
rect 354 -572 388 -396
rect 612 -572 646 -396
rect 870 -572 904 -396
rect 1128 -572 1162 -396
rect 1386 -572 1420 -396
rect 1644 -572 1678 -396
rect 1902 -572 1936 -396
rect 2316 -746 2350 -370
rect 2574 -746 2608 -370
rect -2563 -1803 -2529 -1627
rect -1705 -1803 -1671 -1627
rect -847 -1803 -813 -1627
rect 11 -1803 45 -1627
rect 869 -1803 903 -1627
rect 1727 -1803 1761 -1627
rect 2585 -1803 2619 -1627
rect -2563 -2221 -2529 -2045
rect -1705 -2221 -1671 -2045
rect -847 -2221 -813 -2045
rect 11 -2221 45 -2045
rect 869 -2221 903 -2045
rect 1727 -2221 1761 -2045
rect 2585 -2221 2619 -2045
<< pdiffc >>
rect -2643 1825 -2609 2001
rect -2385 1825 -2351 2001
rect -2127 1825 -2093 2001
rect -1869 1825 -1835 2001
rect -1611 1825 -1577 2001
rect -1353 1825 -1319 2001
rect -1095 1825 -1061 2001
rect -837 1825 -803 2001
rect -579 1825 -545 2001
rect -321 1825 -287 2001
rect -63 1825 -29 2001
rect 356 1824 390 2000
rect 614 1824 648 2000
rect 872 1824 906 2000
rect 1130 1824 1164 2000
rect 1388 1824 1422 2000
rect 1646 1824 1680 2000
rect 1904 1824 1938 2000
rect -2643 1151 -2609 1327
rect -2385 1151 -2351 1327
rect -2127 1151 -2093 1327
rect -1869 1151 -1835 1327
rect -1611 1151 -1577 1327
rect -1353 1151 -1319 1327
rect -1095 1151 -1061 1327
rect -837 1151 -803 1327
rect -579 1151 -545 1327
rect -321 1151 -287 1327
rect -63 1151 -29 1327
rect 356 1150 390 1326
rect 614 1150 648 1326
rect 872 1150 906 1326
rect 1130 1150 1164 1326
rect 1388 1150 1422 1326
rect 1646 1150 1680 1326
rect 1904 1150 1938 1326
rect 2316 1150 2350 1926
rect 2574 1150 2608 1926
<< psubdiff >>
rect -3322 282 -3160 382
rect 3160 282 3322 382
rect -3322 220 -3222 282
rect 3222 220 3322 282
rect -3122 82 -2960 182
rect -240 82 -78 182
rect -3122 20 -3022 82
rect -178 20 -78 82
rect -3122 -1002 -3022 -940
rect -178 -1002 -78 -940
rect -3122 -1102 -2960 -1002
rect -240 -1102 -78 -1002
rect -3122 -1318 -2960 -1218
rect 2960 -1318 3122 -1218
rect -3122 -1380 -3022 -1318
rect 3022 -1380 3122 -1318
rect -3122 -2642 -3022 -2580
rect 3022 -2642 3122 -2580
rect -3122 -2742 -2960 -2642
rect 2960 -2742 3122 -2642
rect -3322 -3422 -3222 -3360
rect 3222 -3422 3322 -3360
rect -3322 -3522 -3160 -3422
rect 3160 -3522 3322 -3422
<< nsubdiff >>
rect -3322 3022 -3160 3122
rect 3160 3022 3322 3122
rect -3322 2960 -3222 3022
rect 3222 2960 3322 3022
rect -3322 718 -3222 780
rect 3222 718 3322 780
rect -3322 618 -3160 718
rect 3160 618 3322 718
<< psubdiffcont >>
rect -3160 282 3160 382
rect -3322 -3360 -3222 220
rect -2960 82 -240 182
rect -3122 -940 -3022 20
rect -178 -940 -78 20
rect -2960 -1102 -240 -1002
rect -2960 -1318 2960 -1218
rect -3122 -2580 -3022 -1380
rect 3022 -2580 3122 -1380
rect -2960 -2742 2960 -2642
rect 3222 -3360 3322 220
rect -3160 -3522 3160 -3422
<< nsubdiffcont >>
rect -3160 3022 3160 3122
rect -3322 780 -3222 2960
rect 3222 780 3322 2960
rect -3160 618 3160 718
<< poly >>
rect -2597 2094 -2397 2110
rect -2597 2060 -2581 2094
rect -2413 2060 -2397 2094
rect -2597 2013 -2397 2060
rect -2339 2094 -2139 2110
rect -2339 2060 -2323 2094
rect -2155 2060 -2139 2094
rect -2339 2013 -2139 2060
rect -2081 2094 -1881 2110
rect -2081 2060 -2065 2094
rect -1897 2060 -1881 2094
rect -2081 2013 -1881 2060
rect -1823 2094 -1623 2110
rect -1823 2060 -1807 2094
rect -1639 2060 -1623 2094
rect -1823 2013 -1623 2060
rect -1565 2094 -1365 2110
rect -1565 2060 -1549 2094
rect -1381 2060 -1365 2094
rect -1565 2013 -1365 2060
rect -1307 2094 -1107 2110
rect -1307 2060 -1291 2094
rect -1123 2060 -1107 2094
rect -1307 2013 -1107 2060
rect -1049 2094 -849 2110
rect -1049 2060 -1033 2094
rect -865 2060 -849 2094
rect -1049 2013 -849 2060
rect -791 2094 -591 2110
rect -791 2060 -775 2094
rect -607 2060 -591 2094
rect -791 2013 -591 2060
rect -533 2094 -333 2110
rect -533 2060 -517 2094
rect -349 2060 -333 2094
rect -533 2013 -333 2060
rect -275 2094 -75 2110
rect -275 2060 -259 2094
rect -91 2060 -75 2094
rect 436 2093 568 2109
rect 436 2076 452 2093
rect -275 2013 -75 2060
rect 402 2059 452 2076
rect 552 2076 568 2093
rect 694 2093 826 2109
rect 694 2076 710 2093
rect 552 2059 602 2076
rect 402 2012 602 2059
rect 660 2059 710 2076
rect 810 2076 826 2093
rect 952 2093 1084 2109
rect 952 2076 968 2093
rect 810 2059 860 2076
rect 660 2012 860 2059
rect 918 2059 968 2076
rect 1068 2076 1084 2093
rect 1210 2093 1342 2109
rect 1210 2076 1226 2093
rect 1068 2059 1118 2076
rect 918 2012 1118 2059
rect 1176 2059 1226 2076
rect 1326 2076 1342 2093
rect 1468 2093 1600 2109
rect 1468 2076 1484 2093
rect 1326 2059 1376 2076
rect 1176 2012 1376 2059
rect 1434 2059 1484 2076
rect 1584 2076 1600 2093
rect 1726 2093 1858 2109
rect 1726 2076 1742 2093
rect 1584 2059 1634 2076
rect 1434 2012 1634 2059
rect 1692 2059 1742 2076
rect 1842 2076 1858 2093
rect 1842 2059 1892 2076
rect 1692 2012 1892 2059
rect 2396 2019 2528 2035
rect -2597 1766 -2397 1813
rect -2597 1732 -2581 1766
rect -2413 1732 -2397 1766
rect -2597 1716 -2397 1732
rect -2339 1766 -2139 1813
rect -2339 1732 -2323 1766
rect -2155 1732 -2139 1766
rect -2339 1716 -2139 1732
rect -2081 1766 -1881 1813
rect -2081 1732 -2065 1766
rect -1897 1732 -1881 1766
rect -2081 1716 -1881 1732
rect -1823 1766 -1623 1813
rect -1823 1732 -1807 1766
rect -1639 1732 -1623 1766
rect -1823 1716 -1623 1732
rect -1565 1766 -1365 1813
rect -1565 1732 -1549 1766
rect -1381 1732 -1365 1766
rect -1565 1716 -1365 1732
rect -1307 1766 -1107 1813
rect -1307 1732 -1291 1766
rect -1123 1732 -1107 1766
rect -1307 1716 -1107 1732
rect -1049 1766 -849 1813
rect -1049 1732 -1033 1766
rect -865 1732 -849 1766
rect -1049 1716 -849 1732
rect -791 1766 -591 1813
rect -791 1732 -775 1766
rect -607 1732 -591 1766
rect -791 1716 -591 1732
rect -533 1766 -333 1813
rect -533 1732 -517 1766
rect -349 1732 -333 1766
rect -533 1716 -333 1732
rect -275 1766 -75 1813
rect 2396 2002 2412 2019
rect 2362 1985 2412 2002
rect 2512 2002 2528 2019
rect 2512 1985 2562 2002
rect 2362 1938 2562 1985
rect -275 1732 -259 1766
rect -91 1732 -75 1766
rect 402 1765 602 1812
rect 402 1748 452 1765
rect -275 1716 -75 1732
rect 436 1731 452 1748
rect 552 1748 602 1765
rect 660 1765 860 1812
rect 660 1748 710 1765
rect 552 1731 568 1748
rect 436 1715 568 1731
rect 694 1731 710 1748
rect 810 1748 860 1765
rect 918 1765 1118 1812
rect 918 1748 968 1765
rect 810 1731 826 1748
rect 694 1715 826 1731
rect 952 1731 968 1748
rect 1068 1748 1118 1765
rect 1176 1765 1376 1812
rect 1176 1748 1226 1765
rect 1068 1731 1084 1748
rect 952 1715 1084 1731
rect 1210 1731 1226 1748
rect 1326 1748 1376 1765
rect 1434 1765 1634 1812
rect 1434 1748 1484 1765
rect 1326 1731 1342 1748
rect 1210 1715 1342 1731
rect 1468 1731 1484 1748
rect 1584 1748 1634 1765
rect 1692 1765 1892 1812
rect 1692 1748 1742 1765
rect 1584 1731 1600 1748
rect 1468 1715 1600 1731
rect 1726 1731 1742 1748
rect 1842 1748 1892 1765
rect 1842 1731 1858 1748
rect 1726 1715 1858 1731
rect -2597 1420 -2397 1436
rect -2597 1386 -2581 1420
rect -2413 1386 -2397 1420
rect -2597 1339 -2397 1386
rect -2339 1420 -2139 1436
rect -2339 1386 -2323 1420
rect -2155 1386 -2139 1420
rect -2339 1339 -2139 1386
rect -2081 1420 -1881 1436
rect -2081 1386 -2065 1420
rect -1897 1386 -1881 1420
rect -2081 1339 -1881 1386
rect -1823 1420 -1623 1436
rect -1823 1386 -1807 1420
rect -1639 1386 -1623 1420
rect -1823 1339 -1623 1386
rect -1565 1420 -1365 1436
rect -1565 1386 -1549 1420
rect -1381 1386 -1365 1420
rect -1565 1339 -1365 1386
rect -1307 1420 -1107 1436
rect -1307 1386 -1291 1420
rect -1123 1386 -1107 1420
rect -1307 1339 -1107 1386
rect -1049 1420 -849 1436
rect -1049 1386 -1033 1420
rect -865 1386 -849 1420
rect -1049 1339 -849 1386
rect -791 1420 -591 1436
rect -791 1386 -775 1420
rect -607 1386 -591 1420
rect -791 1339 -591 1386
rect -533 1420 -333 1436
rect -533 1386 -517 1420
rect -349 1386 -333 1420
rect -533 1339 -333 1386
rect -275 1420 -75 1436
rect -275 1386 -259 1420
rect -91 1386 -75 1420
rect 436 1419 568 1435
rect 436 1402 452 1419
rect -275 1339 -75 1386
rect 402 1385 452 1402
rect 552 1402 568 1419
rect 694 1419 826 1435
rect 694 1402 710 1419
rect 552 1385 602 1402
rect 402 1338 602 1385
rect 660 1385 710 1402
rect 810 1402 826 1419
rect 952 1419 1084 1435
rect 952 1402 968 1419
rect 810 1385 860 1402
rect 660 1338 860 1385
rect 918 1385 968 1402
rect 1068 1402 1084 1419
rect 1210 1419 1342 1435
rect 1210 1402 1226 1419
rect 1068 1385 1118 1402
rect 918 1338 1118 1385
rect 1176 1385 1226 1402
rect 1326 1402 1342 1419
rect 1468 1419 1600 1435
rect 1468 1402 1484 1419
rect 1326 1385 1376 1402
rect 1176 1338 1376 1385
rect 1434 1385 1484 1402
rect 1584 1402 1600 1419
rect 1726 1419 1858 1435
rect 1726 1402 1742 1419
rect 1584 1385 1634 1402
rect 1434 1338 1634 1385
rect 1692 1385 1742 1402
rect 1842 1402 1858 1419
rect 1842 1385 1892 1402
rect 1692 1338 1892 1385
rect -2597 1092 -2397 1139
rect -2597 1058 -2581 1092
rect -2413 1058 -2397 1092
rect -2597 1042 -2397 1058
rect -2339 1092 -2139 1139
rect -2339 1058 -2323 1092
rect -2155 1058 -2139 1092
rect -2339 1042 -2139 1058
rect -2081 1092 -1881 1139
rect -2081 1058 -2065 1092
rect -1897 1058 -1881 1092
rect -2081 1042 -1881 1058
rect -1823 1092 -1623 1139
rect -1823 1058 -1807 1092
rect -1639 1058 -1623 1092
rect -1823 1042 -1623 1058
rect -1565 1092 -1365 1139
rect -1565 1058 -1549 1092
rect -1381 1058 -1365 1092
rect -1565 1042 -1365 1058
rect -1307 1092 -1107 1139
rect -1307 1058 -1291 1092
rect -1123 1058 -1107 1092
rect -1307 1042 -1107 1058
rect -1049 1092 -849 1139
rect -1049 1058 -1033 1092
rect -865 1058 -849 1092
rect -1049 1042 -849 1058
rect -791 1092 -591 1139
rect -791 1058 -775 1092
rect -607 1058 -591 1092
rect -791 1042 -591 1058
rect -533 1092 -333 1139
rect -533 1058 -517 1092
rect -349 1058 -333 1092
rect -533 1042 -333 1058
rect -275 1092 -75 1139
rect -275 1058 -259 1092
rect -91 1058 -75 1092
rect 402 1091 602 1138
rect 402 1074 452 1091
rect -275 1042 -75 1058
rect 436 1057 452 1074
rect 552 1074 602 1091
rect 660 1091 860 1138
rect 660 1074 710 1091
rect 552 1057 568 1074
rect 436 1041 568 1057
rect 694 1057 710 1074
rect 810 1074 860 1091
rect 918 1091 1118 1138
rect 918 1074 968 1091
rect 810 1057 826 1074
rect 694 1041 826 1057
rect 952 1057 968 1074
rect 1068 1074 1118 1091
rect 1176 1091 1376 1138
rect 1176 1074 1226 1091
rect 1068 1057 1084 1074
rect 952 1041 1084 1057
rect 1210 1057 1226 1074
rect 1326 1074 1376 1091
rect 1434 1091 1634 1138
rect 1434 1074 1484 1091
rect 1326 1057 1342 1074
rect 1210 1041 1342 1057
rect 1468 1057 1484 1074
rect 1584 1074 1634 1091
rect 1692 1091 1892 1138
rect 1692 1074 1742 1091
rect 1584 1057 1600 1074
rect 1468 1041 1600 1057
rect 1726 1057 1742 1074
rect 1842 1074 1892 1091
rect 2362 1091 2562 1138
rect 2362 1074 2412 1091
rect 1842 1057 1858 1074
rect 1726 1041 1858 1057
rect 2396 1057 2412 1074
rect 2512 1074 2562 1091
rect 2512 1057 2528 1074
rect 2396 1041 2528 1057
rect -2784 -350 -2652 -334
rect -2784 -367 -2768 -350
rect -2818 -384 -2768 -367
rect -2668 -367 -2652 -350
rect -2526 -350 -2394 -334
rect -2526 -367 -2510 -350
rect -2668 -384 -2618 -367
rect -2818 -422 -2618 -384
rect -2560 -384 -2510 -367
rect -2410 -367 -2394 -350
rect -2268 -350 -2136 -334
rect -2268 -367 -2252 -350
rect -2410 -384 -2360 -367
rect -2560 -422 -2360 -384
rect -2302 -384 -2252 -367
rect -2152 -367 -2136 -350
rect -2010 -350 -1878 -334
rect -2010 -367 -1994 -350
rect -2152 -384 -2102 -367
rect -2302 -422 -2102 -384
rect -2044 -384 -1994 -367
rect -1894 -367 -1878 -350
rect -1752 -350 -1620 -334
rect -1752 -367 -1736 -350
rect -1894 -384 -1844 -367
rect -2044 -422 -1844 -384
rect -1786 -384 -1736 -367
rect -1636 -367 -1620 -350
rect -1494 -350 -1362 -334
rect -1494 -367 -1478 -350
rect -1636 -384 -1586 -367
rect -1786 -422 -1586 -384
rect -1528 -384 -1478 -367
rect -1378 -367 -1362 -350
rect -1236 -350 -1104 -334
rect -1236 -367 -1220 -350
rect -1378 -384 -1328 -367
rect -1528 -422 -1328 -384
rect -1270 -384 -1220 -367
rect -1120 -367 -1104 -350
rect -978 -350 -846 -334
rect -978 -367 -962 -350
rect -1120 -384 -1070 -367
rect -1270 -422 -1070 -384
rect -1012 -384 -962 -367
rect -862 -367 -846 -350
rect -720 -350 -588 -334
rect -720 -367 -704 -350
rect -862 -384 -812 -367
rect -1012 -422 -812 -384
rect -754 -384 -704 -367
rect -604 -367 -588 -350
rect -462 -350 -330 -334
rect -462 -367 -446 -350
rect -604 -384 -554 -367
rect -754 -422 -554 -384
rect -496 -384 -446 -367
rect -346 -367 -330 -350
rect -346 -384 -296 -367
rect -496 -422 -296 -384
rect -2818 -660 -2618 -622
rect -2818 -677 -2768 -660
rect -2784 -694 -2768 -677
rect -2668 -677 -2618 -660
rect -2560 -660 -2360 -622
rect -2560 -677 -2510 -660
rect -2668 -694 -2652 -677
rect -2784 -710 -2652 -694
rect -2526 -694 -2510 -677
rect -2410 -677 -2360 -660
rect -2302 -660 -2102 -622
rect -2302 -677 -2252 -660
rect -2410 -694 -2394 -677
rect -2526 -710 -2394 -694
rect -2268 -694 -2252 -677
rect -2152 -677 -2102 -660
rect -2044 -660 -1844 -622
rect -2044 -677 -1994 -660
rect -2152 -694 -2136 -677
rect -2268 -710 -2136 -694
rect -2010 -694 -1994 -677
rect -1894 -677 -1844 -660
rect -1786 -660 -1586 -622
rect -1786 -677 -1736 -660
rect -1894 -694 -1878 -677
rect -2010 -710 -1878 -694
rect -1752 -694 -1736 -677
rect -1636 -677 -1586 -660
rect -1528 -660 -1328 -622
rect -1528 -677 -1478 -660
rect -1636 -694 -1620 -677
rect -1752 -710 -1620 -694
rect -1494 -694 -1478 -677
rect -1378 -677 -1328 -660
rect -1270 -660 -1070 -622
rect -1270 -677 -1220 -660
rect -1378 -694 -1362 -677
rect -1494 -710 -1362 -694
rect -1236 -694 -1220 -677
rect -1120 -677 -1070 -660
rect -1012 -660 -812 -622
rect -1012 -677 -962 -660
rect -1120 -694 -1104 -677
rect -1236 -710 -1104 -694
rect -978 -694 -962 -677
rect -862 -677 -812 -660
rect -754 -660 -554 -622
rect -754 -677 -704 -660
rect -862 -694 -846 -677
rect -978 -710 -846 -694
rect -720 -694 -704 -677
rect -604 -677 -554 -660
rect -496 -660 -296 -622
rect -496 -677 -446 -660
rect -604 -694 -588 -677
rect -720 -710 -588 -694
rect -462 -694 -446 -677
rect -346 -677 -296 -660
rect -346 -694 -330 -677
rect -462 -710 -330 -694
rect 2396 -286 2528 -270
rect 442 -312 558 -296
rect 442 -329 458 -312
rect 400 -346 458 -329
rect 542 -329 558 -312
rect 700 -312 816 -296
rect 700 -329 716 -312
rect 542 -346 600 -329
rect 400 -384 600 -346
rect 658 -346 716 -329
rect 800 -329 816 -312
rect 958 -312 1074 -296
rect 958 -329 974 -312
rect 800 -346 858 -329
rect 658 -384 858 -346
rect 916 -346 974 -329
rect 1058 -329 1074 -312
rect 1216 -312 1332 -296
rect 1216 -329 1232 -312
rect 1058 -346 1116 -329
rect 916 -384 1116 -346
rect 1174 -346 1232 -329
rect 1316 -329 1332 -312
rect 1474 -312 1590 -296
rect 1474 -329 1490 -312
rect 1316 -346 1374 -329
rect 1174 -384 1374 -346
rect 1432 -346 1490 -329
rect 1574 -329 1590 -312
rect 1732 -312 1848 -296
rect 2396 -303 2412 -286
rect 1732 -329 1748 -312
rect 1574 -346 1632 -329
rect 1432 -384 1632 -346
rect 1690 -346 1748 -329
rect 1832 -329 1848 -312
rect 2362 -320 2412 -303
rect 2512 -303 2528 -286
rect 2512 -320 2562 -303
rect 1832 -346 1890 -329
rect 1690 -384 1890 -346
rect 2362 -358 2562 -320
rect 400 -622 600 -584
rect 400 -639 458 -622
rect 442 -656 458 -639
rect 542 -639 600 -622
rect 658 -622 858 -584
rect 658 -639 716 -622
rect 542 -656 558 -639
rect 442 -672 558 -656
rect 700 -656 716 -639
rect 800 -639 858 -622
rect 916 -622 1116 -584
rect 916 -639 974 -622
rect 800 -656 816 -639
rect 700 -672 816 -656
rect 958 -656 974 -639
rect 1058 -639 1116 -622
rect 1174 -622 1374 -584
rect 1174 -639 1232 -622
rect 1058 -656 1074 -639
rect 958 -672 1074 -656
rect 1216 -656 1232 -639
rect 1316 -639 1374 -622
rect 1432 -622 1632 -584
rect 1432 -639 1490 -622
rect 1316 -656 1332 -639
rect 1216 -672 1332 -656
rect 1474 -656 1490 -639
rect 1574 -639 1632 -622
rect 1690 -622 1890 -584
rect 1690 -639 1748 -622
rect 1574 -656 1590 -639
rect 1474 -672 1590 -656
rect 1732 -656 1748 -639
rect 1832 -639 1890 -622
rect 1832 -656 1848 -639
rect 1732 -672 1848 -656
rect 2362 -796 2562 -758
rect 2362 -813 2412 -796
rect 2396 -830 2412 -813
rect 2512 -813 2562 -796
rect 2512 -830 2528 -813
rect 2396 -846 2528 -830
rect -2363 -1543 -1871 -1527
rect -2363 -1560 -2347 -1543
rect -2517 -1577 -2347 -1560
rect -1887 -1560 -1871 -1543
rect -1505 -1543 -1013 -1527
rect -1505 -1560 -1489 -1543
rect -1887 -1577 -1717 -1560
rect -2517 -1615 -1717 -1577
rect -1659 -1577 -1489 -1560
rect -1029 -1560 -1013 -1543
rect -647 -1543 -155 -1527
rect -647 -1560 -631 -1543
rect -1029 -1577 -859 -1560
rect -1659 -1615 -859 -1577
rect -801 -1577 -631 -1560
rect -171 -1560 -155 -1543
rect 211 -1543 703 -1527
rect 211 -1560 227 -1543
rect -171 -1577 -1 -1560
rect -801 -1615 -1 -1577
rect 57 -1577 227 -1560
rect 687 -1560 703 -1543
rect 1069 -1543 1561 -1527
rect 1069 -1560 1085 -1543
rect 687 -1577 857 -1560
rect 57 -1615 857 -1577
rect 915 -1577 1085 -1560
rect 1545 -1560 1561 -1543
rect 1927 -1543 2419 -1527
rect 1927 -1560 1943 -1543
rect 1545 -1577 1715 -1560
rect 915 -1615 1715 -1577
rect 1773 -1577 1943 -1560
rect 2403 -1560 2419 -1543
rect 2403 -1577 2573 -1560
rect 1773 -1615 2573 -1577
rect -2517 -1853 -1717 -1815
rect -2517 -1870 -2347 -1853
rect -2363 -1887 -2347 -1870
rect -1887 -1870 -1717 -1853
rect -1659 -1853 -859 -1815
rect -1659 -1870 -1489 -1853
rect -1887 -1887 -1871 -1870
rect -2363 -1903 -1871 -1887
rect -1505 -1887 -1489 -1870
rect -1029 -1870 -859 -1853
rect -801 -1853 -1 -1815
rect -801 -1870 -631 -1853
rect -1029 -1887 -1013 -1870
rect -1505 -1903 -1013 -1887
rect -647 -1887 -631 -1870
rect -171 -1870 -1 -1853
rect 57 -1853 857 -1815
rect 57 -1870 227 -1853
rect -171 -1887 -155 -1870
rect -647 -1903 -155 -1887
rect 211 -1887 227 -1870
rect 687 -1870 857 -1853
rect 915 -1853 1715 -1815
rect 915 -1870 1085 -1853
rect 687 -1887 703 -1870
rect 211 -1903 703 -1887
rect 1069 -1887 1085 -1870
rect 1545 -1870 1715 -1853
rect 1773 -1853 2573 -1815
rect 1773 -1870 1943 -1853
rect 1545 -1887 1561 -1870
rect 1069 -1903 1561 -1887
rect 1927 -1887 1943 -1870
rect 2403 -1870 2573 -1853
rect 2403 -1887 2419 -1870
rect 1927 -1903 2419 -1887
rect -2363 -1961 -1871 -1945
rect -2363 -1978 -2347 -1961
rect -2517 -1995 -2347 -1978
rect -1887 -1978 -1871 -1961
rect -1505 -1961 -1013 -1945
rect -1505 -1978 -1489 -1961
rect -1887 -1995 -1717 -1978
rect -2517 -2033 -1717 -1995
rect -1659 -1995 -1489 -1978
rect -1029 -1978 -1013 -1961
rect -647 -1961 -155 -1945
rect -647 -1978 -631 -1961
rect -1029 -1995 -859 -1978
rect -1659 -2033 -859 -1995
rect -801 -1995 -631 -1978
rect -171 -1978 -155 -1961
rect 211 -1961 703 -1945
rect 211 -1978 227 -1961
rect -171 -1995 -1 -1978
rect -801 -2033 -1 -1995
rect 57 -1995 227 -1978
rect 687 -1978 703 -1961
rect 1069 -1961 1561 -1945
rect 1069 -1978 1085 -1961
rect 687 -1995 857 -1978
rect 57 -2033 857 -1995
rect 915 -1995 1085 -1978
rect 1545 -1978 1561 -1961
rect 1927 -1961 2419 -1945
rect 1927 -1978 1943 -1961
rect 1545 -1995 1715 -1978
rect 915 -2033 1715 -1995
rect 1773 -1995 1943 -1978
rect 2403 -1978 2419 -1961
rect 2403 -1995 2573 -1978
rect 1773 -2033 2573 -1995
rect -2517 -2271 -1717 -2233
rect -2517 -2288 -2347 -2271
rect -2363 -2305 -2347 -2288
rect -1887 -2288 -1717 -2271
rect -1659 -2271 -859 -2233
rect -1659 -2288 -1489 -2271
rect -1887 -2305 -1871 -2288
rect -2363 -2321 -1871 -2305
rect -1505 -2305 -1489 -2288
rect -1029 -2288 -859 -2271
rect -801 -2271 -1 -2233
rect -801 -2288 -631 -2271
rect -1029 -2305 -1013 -2288
rect -1505 -2321 -1013 -2305
rect -647 -2305 -631 -2288
rect -171 -2288 -1 -2271
rect 57 -2271 857 -2233
rect 57 -2288 227 -2271
rect -171 -2305 -155 -2288
rect -647 -2321 -155 -2305
rect 211 -2305 227 -2288
rect 687 -2288 857 -2271
rect 915 -2271 1715 -2233
rect 915 -2288 1085 -2271
rect 687 -2305 703 -2288
rect 211 -2321 703 -2305
rect 1069 -2305 1085 -2288
rect 1545 -2288 1715 -2271
rect 1773 -2271 2573 -2233
rect 1773 -2288 1943 -2271
rect 1545 -2305 1561 -2288
rect 1069 -2321 1561 -2305
rect 1927 -2305 1943 -2288
rect 2403 -2288 2573 -2271
rect 2403 -2305 2419 -2288
rect 1927 -2321 2419 -2305
<< polycont >>
rect -2581 2060 -2413 2094
rect -2323 2060 -2155 2094
rect -2065 2060 -1897 2094
rect -1807 2060 -1639 2094
rect -1549 2060 -1381 2094
rect -1291 2060 -1123 2094
rect -1033 2060 -865 2094
rect -775 2060 -607 2094
rect -517 2060 -349 2094
rect -259 2060 -91 2094
rect 452 2059 552 2093
rect 710 2059 810 2093
rect 968 2059 1068 2093
rect 1226 2059 1326 2093
rect 1484 2059 1584 2093
rect 1742 2059 1842 2093
rect -2581 1732 -2413 1766
rect -2323 1732 -2155 1766
rect -2065 1732 -1897 1766
rect -1807 1732 -1639 1766
rect -1549 1732 -1381 1766
rect -1291 1732 -1123 1766
rect -1033 1732 -865 1766
rect -775 1732 -607 1766
rect -517 1732 -349 1766
rect 2412 1985 2512 2019
rect -259 1732 -91 1766
rect 452 1731 552 1765
rect 710 1731 810 1765
rect 968 1731 1068 1765
rect 1226 1731 1326 1765
rect 1484 1731 1584 1765
rect 1742 1731 1842 1765
rect -2581 1386 -2413 1420
rect -2323 1386 -2155 1420
rect -2065 1386 -1897 1420
rect -1807 1386 -1639 1420
rect -1549 1386 -1381 1420
rect -1291 1386 -1123 1420
rect -1033 1386 -865 1420
rect -775 1386 -607 1420
rect -517 1386 -349 1420
rect -259 1386 -91 1420
rect 452 1385 552 1419
rect 710 1385 810 1419
rect 968 1385 1068 1419
rect 1226 1385 1326 1419
rect 1484 1385 1584 1419
rect 1742 1385 1842 1419
rect -2581 1058 -2413 1092
rect -2323 1058 -2155 1092
rect -2065 1058 -1897 1092
rect -1807 1058 -1639 1092
rect -1549 1058 -1381 1092
rect -1291 1058 -1123 1092
rect -1033 1058 -865 1092
rect -775 1058 -607 1092
rect -517 1058 -349 1092
rect -259 1058 -91 1092
rect 452 1057 552 1091
rect 710 1057 810 1091
rect 968 1057 1068 1091
rect 1226 1057 1326 1091
rect 1484 1057 1584 1091
rect 1742 1057 1842 1091
rect 2412 1057 2512 1091
rect -2768 -384 -2668 -350
rect -2510 -384 -2410 -350
rect -2252 -384 -2152 -350
rect -1994 -384 -1894 -350
rect -1736 -384 -1636 -350
rect -1478 -384 -1378 -350
rect -1220 -384 -1120 -350
rect -962 -384 -862 -350
rect -704 -384 -604 -350
rect -446 -384 -346 -350
rect -2768 -694 -2668 -660
rect -2510 -694 -2410 -660
rect -2252 -694 -2152 -660
rect -1994 -694 -1894 -660
rect -1736 -694 -1636 -660
rect -1478 -694 -1378 -660
rect -1220 -694 -1120 -660
rect -962 -694 -862 -660
rect -704 -694 -604 -660
rect -446 -694 -346 -660
rect 458 -346 542 -312
rect 716 -346 800 -312
rect 974 -346 1058 -312
rect 1232 -346 1316 -312
rect 1490 -346 1574 -312
rect 1748 -346 1832 -312
rect 2412 -320 2512 -286
rect 458 -656 542 -622
rect 716 -656 800 -622
rect 974 -656 1058 -622
rect 1232 -656 1316 -622
rect 1490 -656 1574 -622
rect 1748 -656 1832 -622
rect 2412 -830 2512 -796
rect -2347 -1577 -1887 -1543
rect -1489 -1577 -1029 -1543
rect -631 -1577 -171 -1543
rect 227 -1577 687 -1543
rect 1085 -1577 1545 -1543
rect 1943 -1577 2403 -1543
rect -2347 -1887 -1887 -1853
rect -1489 -1887 -1029 -1853
rect -631 -1887 -171 -1853
rect 227 -1887 687 -1853
rect 1085 -1887 1545 -1853
rect 1943 -1887 2403 -1853
rect -2347 -1995 -1887 -1961
rect -1489 -1995 -1029 -1961
rect -631 -1995 -171 -1961
rect 227 -1995 687 -1961
rect 1085 -1995 1545 -1961
rect 1943 -1995 2403 -1961
rect -2347 -2305 -1887 -2271
rect -1489 -2305 -1029 -2271
rect -631 -2305 -171 -2271
rect 227 -2305 687 -2271
rect 1085 -2305 1545 -2271
rect 1943 -2305 2403 -2271
<< locali >>
rect -3322 2960 -3222 3122
rect 3222 2960 3322 3122
rect -2597 2060 -2581 2094
rect -2413 2060 -2397 2094
rect -2339 2060 -2323 2094
rect -2155 2060 -2139 2094
rect -2081 2060 -2065 2094
rect -1897 2060 -1881 2094
rect -1823 2060 -1807 2094
rect -1639 2060 -1623 2094
rect -1565 2060 -1549 2094
rect -1381 2060 -1365 2094
rect -1307 2060 -1291 2094
rect -1123 2060 -1107 2094
rect -1049 2060 -1033 2094
rect -865 2060 -849 2094
rect -791 2060 -775 2094
rect -607 2060 -591 2094
rect -533 2060 -517 2094
rect -349 2060 -333 2094
rect -275 2060 -259 2094
rect -91 2060 -75 2094
rect 436 2059 452 2093
rect 552 2059 568 2093
rect 694 2059 710 2093
rect 810 2059 826 2093
rect 952 2059 968 2093
rect 1068 2059 1084 2093
rect 1210 2059 1226 2093
rect 1326 2059 1342 2093
rect 1468 2059 1484 2093
rect 1584 2059 1600 2093
rect 1726 2059 1742 2093
rect 1842 2059 1858 2093
rect -2643 2001 -2609 2017
rect -2643 1809 -2609 1825
rect -2385 2001 -2351 2017
rect -2385 1809 -2351 1825
rect -2127 2001 -2093 2017
rect -2127 1809 -2093 1825
rect -1869 2001 -1835 2017
rect -1869 1809 -1835 1825
rect -1611 2001 -1577 2017
rect -1611 1809 -1577 1825
rect -1353 2001 -1319 2017
rect -1353 1809 -1319 1825
rect -1095 2001 -1061 2017
rect -1095 1809 -1061 1825
rect -837 2001 -803 2017
rect -837 1809 -803 1825
rect -579 2001 -545 2017
rect -579 1809 -545 1825
rect -321 2001 -287 2017
rect -321 1809 -287 1825
rect -63 2001 -29 2017
rect -63 1809 -29 1825
rect 356 2000 390 2016
rect 356 1808 390 1824
rect 614 2000 648 2016
rect 614 1808 648 1824
rect 872 2000 906 2016
rect 872 1808 906 1824
rect 1130 2000 1164 2016
rect 1130 1808 1164 1824
rect 1388 2000 1422 2016
rect 1388 1808 1422 1824
rect 1646 2000 1680 2016
rect 1646 1808 1680 1824
rect 1904 2000 1938 2016
rect 2396 1985 2412 2019
rect 2512 1985 2528 2019
rect 1904 1808 1938 1824
rect 2316 1926 2350 1942
rect -2597 1732 -2581 1766
rect -2413 1732 -2397 1766
rect -2339 1732 -2323 1766
rect -2155 1732 -2139 1766
rect -2081 1732 -2065 1766
rect -1897 1732 -1881 1766
rect -1823 1732 -1807 1766
rect -1639 1732 -1623 1766
rect -1565 1732 -1549 1766
rect -1381 1732 -1365 1766
rect -1307 1732 -1291 1766
rect -1123 1732 -1107 1766
rect -1049 1732 -1033 1766
rect -865 1732 -849 1766
rect -791 1732 -775 1766
rect -607 1732 -591 1766
rect -533 1732 -517 1766
rect -349 1732 -333 1766
rect -275 1732 -259 1766
rect -91 1732 -75 1766
rect 436 1731 452 1765
rect 552 1731 568 1765
rect 694 1731 710 1765
rect 810 1731 826 1765
rect 952 1731 968 1765
rect 1068 1731 1084 1765
rect 1210 1731 1226 1765
rect 1326 1731 1342 1765
rect 1468 1731 1484 1765
rect 1584 1731 1600 1765
rect 1726 1731 1742 1765
rect 1842 1731 1858 1765
rect -2597 1386 -2581 1420
rect -2413 1386 -2397 1420
rect -2339 1386 -2323 1420
rect -2155 1386 -2139 1420
rect -2081 1386 -2065 1420
rect -1897 1386 -1881 1420
rect -1823 1386 -1807 1420
rect -1639 1386 -1623 1420
rect -1565 1386 -1549 1420
rect -1381 1386 -1365 1420
rect -1307 1386 -1291 1420
rect -1123 1386 -1107 1420
rect -1049 1386 -1033 1420
rect -865 1386 -849 1420
rect -791 1386 -775 1420
rect -607 1386 -591 1420
rect -533 1386 -517 1420
rect -349 1386 -333 1420
rect -275 1386 -259 1420
rect -91 1386 -75 1420
rect 436 1385 452 1419
rect 552 1385 568 1419
rect 694 1385 710 1419
rect 810 1385 826 1419
rect 952 1385 968 1419
rect 1068 1385 1084 1419
rect 1210 1385 1226 1419
rect 1326 1385 1342 1419
rect 1468 1385 1484 1419
rect 1584 1385 1600 1419
rect 1726 1385 1742 1419
rect 1842 1385 1858 1419
rect -2643 1327 -2609 1343
rect -2643 1135 -2609 1151
rect -2385 1327 -2351 1343
rect -2385 1135 -2351 1151
rect -2127 1327 -2093 1343
rect -2127 1135 -2093 1151
rect -1869 1327 -1835 1343
rect -1869 1135 -1835 1151
rect -1611 1327 -1577 1343
rect -1611 1135 -1577 1151
rect -1353 1327 -1319 1343
rect -1353 1135 -1319 1151
rect -1095 1327 -1061 1343
rect -1095 1135 -1061 1151
rect -837 1327 -803 1343
rect -837 1135 -803 1151
rect -579 1327 -545 1343
rect -579 1135 -545 1151
rect -321 1327 -287 1343
rect -321 1135 -287 1151
rect -63 1327 -29 1343
rect -63 1135 -29 1151
rect 356 1326 390 1342
rect 356 1134 390 1150
rect 614 1326 648 1342
rect 614 1134 648 1150
rect 872 1326 906 1342
rect 872 1134 906 1150
rect 1130 1326 1164 1342
rect 1130 1134 1164 1150
rect 1388 1326 1422 1342
rect 1388 1134 1422 1150
rect 1646 1326 1680 1342
rect 1646 1134 1680 1150
rect 1904 1326 1938 1342
rect 1904 1134 1938 1150
rect 2316 1134 2350 1150
rect 2574 1926 2608 1942
rect 2574 1134 2608 1150
rect -2597 1058 -2581 1092
rect -2413 1058 -2397 1092
rect -2339 1058 -2323 1092
rect -2155 1058 -2139 1092
rect -2081 1058 -2065 1092
rect -1897 1058 -1881 1092
rect -1823 1058 -1807 1092
rect -1639 1058 -1623 1092
rect -1565 1058 -1549 1092
rect -1381 1058 -1365 1092
rect -1307 1058 -1291 1092
rect -1123 1058 -1107 1092
rect -1049 1058 -1033 1092
rect -865 1058 -849 1092
rect -791 1058 -775 1092
rect -607 1058 -591 1092
rect -533 1058 -517 1092
rect -349 1058 -333 1092
rect -275 1058 -259 1092
rect -91 1058 -75 1092
rect 436 1057 452 1091
rect 552 1057 568 1091
rect 694 1057 710 1091
rect 810 1057 826 1091
rect 952 1057 968 1091
rect 1068 1057 1084 1091
rect 1210 1057 1226 1091
rect 1326 1057 1342 1091
rect 1468 1057 1484 1091
rect 1584 1057 1600 1091
rect 1726 1057 1742 1091
rect 1842 1057 1858 1091
rect 2396 1057 2412 1091
rect 2512 1057 2528 1091
rect -3322 618 -3222 780
rect 3222 618 3322 780
rect -3322 220 -3222 382
rect 3222 220 3322 382
rect -3122 28 -3022 182
rect -178 28 -78 182
rect -2784 -384 -2768 -350
rect -2668 -384 -2652 -350
rect -2526 -384 -2510 -350
rect -2410 -384 -2394 -350
rect -2268 -384 -2252 -350
rect -2152 -384 -2136 -350
rect -2010 -384 -1994 -350
rect -1894 -384 -1878 -350
rect -1752 -384 -1736 -350
rect -1636 -384 -1620 -350
rect -1494 -384 -1478 -350
rect -1378 -384 -1362 -350
rect -1236 -384 -1220 -350
rect -1120 -384 -1104 -350
rect -978 -384 -962 -350
rect -862 -384 -846 -350
rect -720 -384 -704 -350
rect -604 -384 -588 -350
rect -462 -384 -446 -350
rect -346 -384 -330 -350
rect -2864 -434 -2830 -418
rect -2864 -626 -2830 -610
rect -2606 -434 -2572 -418
rect -2606 -626 -2572 -610
rect -2348 -434 -2314 -418
rect -2348 -626 -2314 -610
rect -2090 -434 -2056 -418
rect -2090 -626 -2056 -610
rect -1832 -434 -1798 -418
rect -1832 -626 -1798 -610
rect -1574 -434 -1540 -418
rect -1574 -626 -1540 -610
rect -1316 -434 -1282 -418
rect -1316 -626 -1282 -610
rect -1058 -434 -1024 -418
rect -1058 -626 -1024 -610
rect -800 -434 -766 -418
rect -800 -626 -766 -610
rect -542 -434 -508 -418
rect -542 -626 -508 -610
rect -284 -434 -250 -418
rect -284 -626 -250 -610
rect -2784 -694 -2768 -660
rect -2668 -694 -2652 -660
rect -2526 -694 -2510 -660
rect -2410 -694 -2394 -660
rect -2268 -694 -2252 -660
rect -2152 -694 -2136 -660
rect -2010 -694 -1994 -660
rect -1894 -694 -1878 -660
rect -1752 -694 -1736 -660
rect -1636 -694 -1620 -660
rect -1494 -694 -1478 -660
rect -1378 -694 -1362 -660
rect -1236 -694 -1220 -660
rect -1120 -694 -1104 -660
rect -978 -694 -962 -660
rect -862 -694 -846 -660
rect -720 -694 -704 -660
rect -604 -694 -588 -660
rect -462 -694 -446 -660
rect -346 -694 -330 -660
rect -3122 -1102 -3022 -948
rect 442 -346 458 -312
rect 542 -346 558 -312
rect 700 -346 716 -312
rect 800 -346 816 -312
rect 958 -346 974 -312
rect 1058 -346 1074 -312
rect 1216 -346 1232 -312
rect 1316 -346 1332 -312
rect 1474 -346 1490 -312
rect 1574 -346 1590 -312
rect 1732 -346 1748 -312
rect 1832 -346 1848 -312
rect 2396 -320 2412 -286
rect 2512 -320 2528 -286
rect 2316 -370 2350 -354
rect 354 -396 388 -380
rect 354 -588 388 -572
rect 612 -396 646 -380
rect 612 -588 646 -572
rect 870 -396 904 -380
rect 870 -588 904 -572
rect 1128 -396 1162 -380
rect 1128 -588 1162 -572
rect 1386 -396 1420 -380
rect 1386 -588 1420 -572
rect 1644 -396 1678 -380
rect 1644 -588 1678 -572
rect 1902 -396 1936 -380
rect 1902 -588 1936 -572
rect 442 -656 458 -622
rect 542 -656 558 -622
rect 700 -656 716 -622
rect 800 -656 816 -622
rect 958 -656 974 -622
rect 1058 -656 1074 -622
rect 1216 -656 1232 -622
rect 1316 -656 1332 -622
rect 1474 -656 1490 -622
rect 1574 -656 1590 -622
rect 1732 -656 1748 -622
rect 1832 -656 1848 -622
rect 2316 -762 2350 -746
rect 2574 -370 2608 -354
rect 2574 -762 2608 -746
rect 2396 -830 2412 -796
rect 2512 -830 2528 -796
rect -178 -1102 -78 -948
rect -3122 -1380 -3022 -1218
rect 3022 -1380 3122 -1218
rect -2363 -1577 -2347 -1543
rect -1887 -1577 -1871 -1543
rect -1505 -1577 -1489 -1543
rect -1029 -1577 -1013 -1543
rect -647 -1577 -631 -1543
rect -171 -1577 -155 -1543
rect 211 -1577 227 -1543
rect 687 -1577 703 -1543
rect 1069 -1577 1085 -1543
rect 1545 -1577 1561 -1543
rect 1927 -1577 1943 -1543
rect 2403 -1577 2419 -1543
rect -2563 -1627 -2529 -1611
rect -2563 -1819 -2529 -1803
rect -1705 -1627 -1671 -1611
rect -1705 -1819 -1671 -1803
rect -847 -1627 -813 -1611
rect -847 -1819 -813 -1803
rect 11 -1627 45 -1611
rect 11 -1819 45 -1803
rect 869 -1627 903 -1611
rect 869 -1819 903 -1803
rect 1727 -1627 1761 -1611
rect 1727 -1819 1761 -1803
rect 2585 -1627 2619 -1611
rect 2585 -1819 2619 -1803
rect -2363 -1887 -2347 -1853
rect -1887 -1887 -1871 -1853
rect -1505 -1887 -1489 -1853
rect -1029 -1887 -1013 -1853
rect -647 -1887 -631 -1853
rect -171 -1887 -155 -1853
rect 211 -1887 227 -1853
rect 687 -1887 703 -1853
rect 1069 -1887 1085 -1853
rect 1545 -1887 1561 -1853
rect 1927 -1887 1943 -1853
rect 2403 -1887 2419 -1853
rect -2363 -1995 -2347 -1961
rect -1887 -1995 -1871 -1961
rect -1505 -1995 -1489 -1961
rect -1029 -1995 -1013 -1961
rect -647 -1995 -631 -1961
rect -171 -1995 -155 -1961
rect 211 -1995 227 -1961
rect 687 -1995 703 -1961
rect 1069 -1995 1085 -1961
rect 1545 -1995 1561 -1961
rect 1927 -1995 1943 -1961
rect 2403 -1995 2419 -1961
rect -2563 -2045 -2529 -2029
rect -2563 -2237 -2529 -2221
rect -1705 -2045 -1671 -2029
rect -1705 -2237 -1671 -2221
rect -847 -2045 -813 -2029
rect -847 -2237 -813 -2221
rect 11 -2045 45 -2029
rect 11 -2237 45 -2221
rect 869 -2045 903 -2029
rect 869 -2237 903 -2221
rect 1727 -2045 1761 -2029
rect 1727 -2237 1761 -2221
rect 2585 -2045 2619 -2029
rect 2585 -2237 2619 -2221
rect -2363 -2305 -2347 -2271
rect -1887 -2305 -1871 -2271
rect -1505 -2305 -1489 -2271
rect -1029 -2305 -1013 -2271
rect -647 -2305 -631 -2271
rect -171 -2305 -155 -2271
rect 211 -2305 227 -2271
rect 687 -2305 703 -2271
rect 1069 -2305 1085 -2271
rect 1545 -2305 1561 -2271
rect 1927 -2305 1943 -2271
rect 2403 -2305 2419 -2271
rect -3122 -2742 -3022 -2580
rect 3022 -2742 3122 -2580
rect -3322 -3522 -3222 -3360
rect 3222 -3522 3322 -3360
<< viali >>
rect -3222 3022 -3160 3122
rect -3160 3022 3160 3122
rect 3160 3022 3222 3122
rect -3322 833 -3222 2907
rect -2539 2060 -2455 2094
rect -2281 2060 -2197 2094
rect -2023 2060 -1939 2094
rect -1765 2060 -1681 2094
rect -1507 2060 -1423 2094
rect -1249 2060 -1165 2094
rect -991 2060 -907 2094
rect -733 2060 -649 2094
rect -475 2060 -391 2094
rect -217 2060 -133 2094
rect 460 2059 544 2093
rect 718 2059 802 2093
rect 976 2059 1060 2093
rect 1234 2059 1318 2093
rect 1492 2059 1576 2093
rect 1750 2059 1834 2093
rect -2643 1825 -2609 2001
rect -2385 1825 -2351 2001
rect -2127 1825 -2093 2001
rect -1869 1825 -1835 2001
rect -1611 1825 -1577 2001
rect -1353 1825 -1319 2001
rect -1095 1825 -1061 2001
rect -837 1825 -803 2001
rect -579 1825 -545 2001
rect -321 1825 -287 2001
rect -63 1825 -29 2001
rect 356 1824 390 2000
rect 614 1824 648 2000
rect 872 1824 906 2000
rect 1130 1824 1164 2000
rect 1388 1824 1422 2000
rect 1646 1824 1680 2000
rect 1904 1824 1938 2000
rect 2420 1985 2504 2019
rect -2539 1732 -2455 1766
rect -2281 1732 -2197 1766
rect -2023 1732 -1939 1766
rect -1765 1732 -1681 1766
rect -1507 1732 -1423 1766
rect -1249 1732 -1165 1766
rect -991 1732 -907 1766
rect -733 1732 -649 1766
rect -475 1732 -391 1766
rect -217 1732 -133 1766
rect 460 1731 544 1765
rect 718 1731 802 1765
rect 976 1731 1060 1765
rect 1234 1731 1318 1765
rect 1492 1731 1576 1765
rect 1750 1731 1834 1765
rect -2539 1386 -2455 1420
rect -2281 1386 -2197 1420
rect -2023 1386 -1939 1420
rect -1765 1386 -1681 1420
rect -1507 1386 -1423 1420
rect -1249 1386 -1165 1420
rect -991 1386 -907 1420
rect -733 1386 -649 1420
rect -475 1386 -391 1420
rect -217 1386 -133 1420
rect 460 1385 544 1419
rect 718 1385 802 1419
rect 976 1385 1060 1419
rect 1234 1385 1318 1419
rect 1492 1385 1576 1419
rect 1750 1385 1834 1419
rect -2643 1151 -2609 1327
rect -2385 1151 -2351 1327
rect -2127 1151 -2093 1327
rect -1869 1151 -1835 1327
rect -1611 1151 -1577 1327
rect -1353 1151 -1319 1327
rect -1095 1151 -1061 1327
rect -837 1151 -803 1327
rect -579 1151 -545 1327
rect -321 1151 -287 1327
rect -63 1151 -29 1327
rect 356 1150 390 1326
rect 614 1150 648 1326
rect 872 1150 906 1326
rect 1130 1150 1164 1326
rect 1388 1150 1422 1326
rect 1646 1150 1680 1326
rect 1904 1150 1938 1326
rect 2316 1150 2350 1926
rect 2574 1150 2608 1926
rect -2539 1058 -2455 1092
rect -2281 1058 -2197 1092
rect -2023 1058 -1939 1092
rect -1765 1058 -1681 1092
rect -1507 1058 -1423 1092
rect -1249 1058 -1165 1092
rect -991 1058 -907 1092
rect -733 1058 -649 1092
rect -475 1058 -391 1092
rect -217 1058 -133 1092
rect 460 1057 544 1091
rect 718 1057 802 1091
rect 976 1057 1060 1091
rect 1234 1057 1318 1091
rect 1492 1057 1576 1091
rect 1750 1057 1834 1091
rect 2420 1057 2504 1091
rect 3222 833 3322 2907
rect -3222 618 -3160 718
rect -3160 618 3160 718
rect 3160 618 3222 718
rect -3222 282 -3160 382
rect -3160 282 3160 382
rect 3160 282 3222 382
rect -3322 -3237 -3222 97
rect -3022 82 -2960 182
rect -2960 82 -240 182
rect -240 82 -178 182
rect -3122 20 -3022 28
rect -3122 -940 -3022 20
rect -178 20 -78 28
rect -2760 -384 -2676 -350
rect -2502 -384 -2418 -350
rect -2244 -384 -2160 -350
rect -1986 -384 -1902 -350
rect -1728 -384 -1644 -350
rect -1470 -384 -1386 -350
rect -1212 -384 -1128 -350
rect -954 -384 -870 -350
rect -696 -384 -612 -350
rect -438 -384 -354 -350
rect -2864 -610 -2830 -434
rect -2606 -610 -2572 -434
rect -2348 -610 -2314 -434
rect -2090 -610 -2056 -434
rect -1832 -610 -1798 -434
rect -1574 -610 -1540 -434
rect -1316 -610 -1282 -434
rect -1058 -610 -1024 -434
rect -800 -610 -766 -434
rect -542 -610 -508 -434
rect -284 -610 -250 -434
rect -2760 -694 -2676 -660
rect -2502 -694 -2418 -660
rect -2244 -694 -2160 -660
rect -1986 -694 -1902 -660
rect -1728 -694 -1644 -660
rect -1470 -694 -1386 -660
rect -1212 -694 -1128 -660
rect -954 -694 -870 -660
rect -696 -694 -612 -660
rect -438 -694 -354 -660
rect -3122 -948 -3022 -940
rect -178 -940 -78 20
rect 458 -346 542 -312
rect 716 -346 800 -312
rect 974 -346 1058 -312
rect 1232 -346 1316 -312
rect 1490 -346 1574 -312
rect 1748 -346 1832 -312
rect 2420 -320 2504 -286
rect 354 -572 388 -396
rect 612 -572 646 -396
rect 870 -572 904 -396
rect 1128 -572 1162 -396
rect 1386 -572 1420 -396
rect 1644 -572 1678 -396
rect 1902 -572 1936 -396
rect 458 -656 542 -622
rect 716 -656 800 -622
rect 974 -656 1058 -622
rect 1232 -656 1316 -622
rect 1490 -656 1574 -622
rect 1748 -656 1832 -622
rect 2316 -746 2350 -370
rect 2574 -746 2608 -370
rect 2420 -830 2504 -796
rect -178 -948 -78 -940
rect -3022 -1102 -2960 -1002
rect -2960 -1102 -240 -1002
rect -240 -1102 -178 -1002
rect -3022 -1318 -2960 -1218
rect -2960 -1318 2960 -1218
rect 2960 -1318 3022 -1218
rect -3122 -2576 -3022 -1384
rect -2309 -1577 -1925 -1543
rect -1451 -1577 -1067 -1543
rect -593 -1577 -209 -1543
rect 265 -1577 649 -1543
rect 1123 -1577 1507 -1543
rect 1981 -1577 2365 -1543
rect -2563 -1803 -2529 -1627
rect -1705 -1803 -1671 -1627
rect -847 -1803 -813 -1627
rect 11 -1803 45 -1627
rect 869 -1803 903 -1627
rect 1727 -1803 1761 -1627
rect 2585 -1803 2619 -1627
rect -2309 -1887 -1925 -1853
rect -1451 -1887 -1067 -1853
rect -593 -1887 -209 -1853
rect 265 -1887 649 -1853
rect 1123 -1887 1507 -1853
rect 1981 -1887 2365 -1853
rect -2309 -1995 -1925 -1961
rect -1451 -1995 -1067 -1961
rect -593 -1995 -209 -1961
rect 265 -1995 649 -1961
rect 1123 -1995 1507 -1961
rect 1981 -1995 2365 -1961
rect -2563 -2221 -2529 -2045
rect -1705 -2221 -1671 -2045
rect -847 -2221 -813 -2045
rect 11 -2221 45 -2045
rect 869 -2221 903 -2045
rect 1727 -2221 1761 -2045
rect 2585 -2221 2619 -2045
rect -2309 -2305 -1925 -2271
rect -1451 -2305 -1067 -2271
rect -593 -2305 -209 -2271
rect 265 -2305 649 -2271
rect 1123 -2305 1507 -2271
rect 1981 -2305 2365 -2271
rect 3022 -2576 3122 -1384
rect -3022 -2742 -2960 -2642
rect -2960 -2742 2960 -2642
rect 2960 -2742 3022 -2642
rect 3222 -3237 3322 97
rect -3222 -3522 -3160 -3422
rect -3160 -3522 3160 -3422
rect 3160 -3522 3222 -3422
<< metal1 >>
rect -3328 3122 3328 3128
rect -3328 3022 -3222 3122
rect 3222 3022 3328 3122
rect -3328 3016 3328 3022
rect -3328 2907 -3216 3016
rect -3328 833 -3322 2907
rect -3222 833 -3216 2907
rect -2616 2716 -2606 3016
rect 2606 2716 2616 3016
rect 3216 2907 3328 3016
rect -2674 2528 2566 2562
rect -2674 2456 -2646 2528
rect 2544 2456 2566 2528
rect -2674 2430 2566 2456
rect -2782 2146 -2776 2206
rect -2716 2146 -2710 2206
rect -2776 978 -2716 2146
rect -2654 2001 -2594 2430
rect -2551 2094 -2443 2100
rect -2551 2060 -2539 2094
rect -2455 2060 -2443 2094
rect -2551 2054 -2443 2060
rect -2654 1825 -2643 2001
rect -2609 1825 -2594 2001
rect -2654 1602 -2594 1825
rect -2400 2001 -2340 2430
rect -2272 2146 -2266 2206
rect -2206 2146 -2200 2206
rect -2266 2100 -2206 2146
rect -2293 2094 -2185 2100
rect -2293 2060 -2281 2094
rect -2197 2060 -2185 2094
rect -2293 2054 -2185 2060
rect -2035 2094 -1927 2100
rect -2035 2060 -2023 2094
rect -1939 2060 -1927 2094
rect -2035 2054 -1927 2060
rect -2400 1825 -2385 2001
rect -2351 1825 -2340 2001
rect -2133 2001 -2087 2013
rect -2133 1890 -2127 2001
rect -2551 1766 -2443 1772
rect -2551 1732 -2539 1766
rect -2455 1732 -2443 1766
rect -2551 1726 -2443 1732
rect -2528 1602 -2468 1726
rect -2400 1602 -2340 1825
rect -2138 1825 -2127 1890
rect -2093 1890 -2087 2001
rect -1880 2001 -1820 2430
rect -1628 2146 -1622 2206
rect -1562 2146 -1556 2206
rect -1502 2146 -1496 2206
rect -1436 2146 -1430 2206
rect -1777 2094 -1669 2100
rect -1777 2060 -1765 2094
rect -1681 2060 -1669 2094
rect -1777 2054 -1669 2060
rect -2093 1825 -2078 1890
rect -2293 1766 -2185 1772
rect -2293 1732 -2281 1766
rect -2197 1732 -2185 1766
rect -2293 1726 -2185 1732
rect -2270 1664 -2210 1726
rect -2276 1604 -2270 1664
rect -2210 1604 -2204 1664
rect -2654 1542 -2340 1602
rect -2654 1327 -2594 1542
rect -2528 1426 -2468 1542
rect -2551 1420 -2443 1426
rect -2551 1386 -2539 1420
rect -2455 1386 -2443 1420
rect -2551 1380 -2443 1386
rect -2654 1318 -2643 1327
rect -2649 1151 -2643 1318
rect -2609 1318 -2594 1327
rect -2400 1327 -2340 1542
rect -2270 1426 -2210 1604
rect -2138 1530 -2078 1825
rect -1880 1825 -1869 2001
rect -1835 1825 -1820 2001
rect -1622 2001 -1562 2146
rect -1496 2100 -1436 2146
rect -1519 2094 -1411 2100
rect -1519 2060 -1507 2094
rect -1423 2060 -1411 2094
rect -1519 2054 -1411 2060
rect -1622 1966 -1611 2001
rect -2035 1766 -1927 1772
rect -2035 1732 -2023 1766
rect -1939 1732 -1927 1766
rect -2035 1726 -1927 1732
rect -2008 1530 -1948 1726
rect -2144 1470 -2138 1530
rect -2078 1470 -2072 1530
rect -2014 1470 -2008 1530
rect -1948 1470 -1942 1530
rect -2008 1426 -1948 1470
rect -2293 1420 -2185 1426
rect -2293 1386 -2281 1420
rect -2197 1386 -2185 1420
rect -2293 1380 -2185 1386
rect -2035 1420 -1927 1426
rect -2035 1386 -2023 1420
rect -1939 1386 -1927 1420
rect -2035 1380 -1927 1386
rect -2609 1151 -2603 1318
rect -2400 1284 -2385 1327
rect -2649 1139 -2603 1151
rect -2391 1151 -2385 1284
rect -2351 1284 -2340 1327
rect -2133 1327 -2087 1339
rect -2351 1151 -2345 1284
rect -2133 1198 -2127 1327
rect -2391 1139 -2345 1151
rect -2142 1151 -2127 1198
rect -2093 1198 -2087 1327
rect -1880 1327 -1820 1825
rect -1617 1825 -1611 1966
rect -1577 1966 -1562 2001
rect -1366 2001 -1306 2430
rect -1238 2146 -1232 2206
rect -1172 2146 -1166 2206
rect -1232 2100 -1172 2146
rect -1261 2094 -1153 2100
rect -1261 2060 -1249 2094
rect -1165 2060 -1153 2094
rect -1261 2054 -1153 2060
rect -1003 2094 -895 2100
rect -1003 2060 -991 2094
rect -907 2060 -895 2094
rect -1003 2054 -895 2060
rect -1577 1825 -1571 1966
rect -1617 1813 -1571 1825
rect -1366 1825 -1353 2001
rect -1319 1825 -1306 2001
rect -1101 2001 -1055 2013
rect -1101 1872 -1095 2001
rect -1777 1766 -1669 1772
rect -1777 1732 -1765 1766
rect -1681 1732 -1669 1766
rect -1777 1726 -1669 1732
rect -1519 1766 -1411 1772
rect -1519 1732 -1507 1766
rect -1423 1732 -1411 1766
rect -1519 1726 -1411 1732
rect -1750 1530 -1690 1726
rect -1494 1664 -1434 1726
rect -1500 1604 -1494 1664
rect -1434 1604 -1428 1664
rect -1756 1470 -1750 1530
rect -1690 1470 -1684 1530
rect -1634 1470 -1628 1530
rect -1568 1470 -1562 1530
rect -1750 1426 -1690 1470
rect -1777 1420 -1669 1426
rect -1777 1386 -1765 1420
rect -1681 1386 -1669 1420
rect -1777 1380 -1669 1386
rect -1880 1292 -1869 1327
rect -2093 1151 -2082 1198
rect -2551 1092 -2443 1098
rect -2551 1058 -2539 1092
rect -2455 1058 -2443 1092
rect -2551 1052 -2443 1058
rect -2293 1092 -2185 1098
rect -2293 1058 -2281 1092
rect -2197 1058 -2185 1092
rect -2293 1052 -2185 1058
rect -2274 978 -2214 1052
rect -2142 978 -2082 1151
rect -1875 1151 -1869 1292
rect -1835 1292 -1820 1327
rect -1628 1327 -1568 1470
rect -1494 1426 -1434 1604
rect -1519 1420 -1411 1426
rect -1519 1386 -1507 1420
rect -1423 1386 -1411 1420
rect -1519 1380 -1411 1386
rect -1835 1151 -1829 1292
rect -1628 1280 -1611 1327
rect -1875 1139 -1829 1151
rect -1617 1151 -1611 1280
rect -1577 1280 -1568 1327
rect -1366 1327 -1306 1825
rect -1112 1825 -1095 1872
rect -1061 1872 -1055 2001
rect -846 2001 -786 2430
rect -602 2146 -596 2206
rect -536 2146 -530 2206
rect -470 2146 -464 2206
rect -404 2146 -398 2206
rect -745 2094 -637 2100
rect -745 2060 -733 2094
rect -649 2060 -637 2094
rect -745 2054 -637 2060
rect -1061 1825 -1052 1872
rect -1261 1766 -1153 1772
rect -1261 1732 -1249 1766
rect -1165 1732 -1153 1766
rect -1261 1726 -1153 1732
rect -1240 1664 -1180 1726
rect -1246 1604 -1240 1664
rect -1180 1604 -1174 1664
rect -1240 1426 -1180 1604
rect -1112 1530 -1052 1825
rect -846 1825 -837 2001
rect -803 1825 -786 2001
rect -596 2001 -536 2146
rect -464 2100 -404 2146
rect -487 2094 -379 2100
rect -487 2060 -475 2094
rect -391 2060 -379 2094
rect -487 2054 -379 2060
rect -596 1940 -579 2001
rect -1003 1766 -895 1772
rect -1003 1732 -991 1766
rect -907 1732 -895 1766
rect -1003 1726 -895 1732
rect -980 1530 -920 1726
rect -1118 1470 -1112 1530
rect -1052 1470 -1046 1530
rect -986 1470 -980 1530
rect -920 1470 -914 1530
rect -980 1426 -920 1470
rect -1261 1420 -1153 1426
rect -1261 1386 -1249 1420
rect -1165 1386 -1153 1420
rect -1261 1380 -1153 1386
rect -1003 1420 -895 1426
rect -1003 1386 -991 1420
rect -907 1386 -895 1420
rect -1003 1380 -895 1386
rect -1366 1298 -1353 1327
rect -1577 1151 -1571 1280
rect -1617 1139 -1571 1151
rect -1359 1151 -1353 1298
rect -1319 1298 -1306 1327
rect -1101 1327 -1055 1339
rect -1319 1151 -1313 1298
rect -1101 1190 -1095 1327
rect -1359 1139 -1313 1151
rect -1108 1151 -1095 1190
rect -1061 1190 -1055 1327
rect -846 1327 -786 1825
rect -585 1825 -579 1940
rect -545 1940 -536 2001
rect -334 2001 -274 2430
rect -229 2094 -121 2100
rect -229 2060 -217 2094
rect -133 2060 -121 2094
rect -229 2054 -121 2060
rect -545 1825 -539 1940
rect -585 1813 -539 1825
rect -334 1825 -321 2001
rect -287 1825 -274 2001
rect -745 1766 -637 1772
rect -745 1732 -733 1766
rect -649 1732 -637 1766
rect -745 1726 -637 1732
rect -487 1766 -379 1772
rect -487 1732 -475 1766
rect -391 1732 -379 1766
rect -487 1726 -379 1732
rect -720 1530 -660 1726
rect -464 1664 -404 1726
rect -470 1604 -464 1664
rect -404 1604 -398 1664
rect -726 1470 -720 1530
rect -660 1470 -654 1530
rect -602 1470 -596 1530
rect -536 1470 -530 1530
rect -720 1426 -660 1470
rect -745 1420 -637 1426
rect -745 1386 -733 1420
rect -649 1386 -637 1420
rect -745 1380 -637 1386
rect -846 1284 -837 1327
rect -1061 1151 -1048 1190
rect -2035 1092 -1927 1098
rect -2035 1058 -2023 1092
rect -1939 1058 -1927 1092
rect -2035 1052 -1927 1058
rect -1777 1092 -1669 1098
rect -1777 1058 -1765 1092
rect -1681 1058 -1669 1092
rect -1777 1052 -1669 1058
rect -1519 1092 -1411 1098
rect -1519 1058 -1507 1092
rect -1423 1058 -1411 1092
rect -1519 1052 -1411 1058
rect -1261 1092 -1153 1098
rect -1261 1058 -1249 1092
rect -1165 1058 -1153 1092
rect -1261 1052 -1153 1058
rect -2782 918 -2776 978
rect -2716 918 -2710 978
rect -2280 918 -2274 978
rect -2214 918 -2208 978
rect -2148 918 -2142 978
rect -2082 918 -2076 978
rect -2014 874 -1954 1052
rect -1500 978 -1440 1052
rect -1240 978 -1180 1052
rect -1108 978 -1048 1151
rect -843 1151 -837 1284
rect -803 1284 -786 1327
rect -596 1327 -536 1470
rect -464 1426 -404 1604
rect -334 1598 -274 1825
rect -76 2001 -16 2430
rect 210 2258 216 2318
rect 276 2258 282 2318
rect 594 2258 600 2318
rect 660 2258 666 2318
rect -76 1825 -63 2001
rect -29 1825 -16 2001
rect -229 1766 -121 1772
rect -229 1732 -217 1766
rect -133 1732 -121 1766
rect -229 1726 -121 1732
rect -210 1598 -150 1726
rect -76 1598 -16 1825
rect -334 1538 -16 1598
rect -487 1420 -379 1426
rect -487 1386 -475 1420
rect -391 1386 -379 1420
rect -487 1380 -379 1386
rect -803 1151 -797 1284
rect -596 1272 -579 1327
rect -843 1139 -797 1151
rect -585 1151 -579 1272
rect -545 1272 -536 1327
rect -334 1327 -274 1538
rect -210 1426 -150 1538
rect -229 1420 -121 1426
rect -229 1386 -217 1420
rect -133 1386 -121 1420
rect -229 1380 -121 1386
rect -334 1276 -321 1327
rect -545 1151 -539 1272
rect -585 1139 -539 1151
rect -327 1151 -321 1276
rect -287 1276 -274 1327
rect -76 1327 -16 1538
rect -76 1302 -63 1327
rect -287 1151 -281 1276
rect -327 1139 -281 1151
rect -69 1151 -63 1302
rect -29 1302 -16 1327
rect -29 1151 -23 1302
rect -69 1139 -23 1151
rect -1003 1092 -895 1098
rect -1003 1058 -991 1092
rect -907 1058 -895 1092
rect -1003 1052 -895 1058
rect -745 1092 -637 1098
rect -745 1058 -733 1092
rect -649 1058 -637 1092
rect -745 1052 -637 1058
rect -487 1092 -379 1098
rect -487 1058 -475 1092
rect -391 1058 -379 1092
rect -487 1052 -379 1058
rect -229 1092 -121 1098
rect -229 1058 -217 1092
rect -133 1058 -121 1092
rect -229 1052 -121 1058
rect -1506 918 -1500 978
rect -1440 918 -1434 978
rect -1246 918 -1240 978
rect -1180 918 -1174 978
rect -1114 918 -1108 978
rect -1048 918 -1042 978
rect -3328 724 -3216 833
rect -2020 814 -2014 874
rect -1954 814 -1948 874
rect -724 866 -664 1052
rect -464 978 -404 1052
rect -470 918 -464 978
rect -404 918 -398 978
rect 216 874 276 2258
rect 448 2093 556 2099
rect 448 2059 460 2093
rect 544 2059 556 2093
rect 448 2053 556 2059
rect 350 2000 396 2012
rect 350 1858 356 2000
rect 344 1824 356 1858
rect 390 1858 396 2000
rect 600 2000 660 2258
rect 706 2093 814 2099
rect 706 2059 718 2093
rect 802 2059 814 2093
rect 706 2053 814 2059
rect 390 1824 404 1858
rect 344 1664 404 1824
rect 600 1824 614 2000
rect 648 1824 660 2000
rect 448 1765 556 1771
rect 448 1731 460 1765
rect 544 1731 556 1765
rect 448 1725 556 1731
rect 474 1664 534 1725
rect 600 1664 660 1824
rect 856 2000 916 2430
rect 982 2146 988 2206
rect 1048 2146 1054 2206
rect 1238 2146 1244 2206
rect 1304 2146 1310 2206
rect 988 2099 1048 2146
rect 1244 2099 1304 2146
rect 964 2093 1072 2099
rect 964 2059 976 2093
rect 1060 2059 1072 2093
rect 964 2053 1072 2059
rect 1222 2093 1330 2099
rect 1222 2059 1234 2093
rect 1318 2059 1330 2093
rect 1222 2053 1330 2059
rect 856 1824 872 2000
rect 906 1824 916 2000
rect 1124 2000 1170 2012
rect 1124 1854 1130 2000
rect 706 1765 814 1771
rect 706 1731 718 1765
rect 802 1731 814 1765
rect 706 1725 814 1731
rect 344 1604 660 1664
rect 730 1662 790 1725
rect 724 1602 730 1662
rect 790 1602 796 1662
rect 592 1478 598 1538
rect 658 1478 664 1538
rect 448 1419 556 1425
rect 448 1385 460 1419
rect 544 1385 556 1419
rect 448 1379 556 1385
rect 350 1326 396 1338
rect 350 1192 356 1326
rect 342 1150 356 1192
rect 390 1192 396 1326
rect 598 1326 658 1478
rect 706 1419 814 1425
rect 706 1385 718 1419
rect 802 1385 814 1419
rect 706 1379 814 1385
rect 390 1150 402 1192
rect 342 988 402 1150
rect 598 1150 614 1326
rect 648 1150 658 1326
rect 856 1326 916 1824
rect 1116 1824 1130 1854
rect 1164 1854 1170 2000
rect 1374 2000 1434 2430
rect 1626 2258 1632 2318
rect 1692 2258 1698 2318
rect 1480 2093 1588 2099
rect 1480 2059 1492 2093
rect 1576 2059 1588 2093
rect 1480 2053 1588 2059
rect 1164 1824 1176 1854
rect 964 1765 1072 1771
rect 964 1731 976 1765
rect 1060 1731 1072 1765
rect 964 1725 1072 1731
rect 982 1602 988 1662
rect 1048 1602 1054 1662
rect 988 1425 1048 1602
rect 1116 1538 1176 1824
rect 1374 1824 1388 2000
rect 1422 1824 1434 2000
rect 1222 1765 1330 1771
rect 1222 1731 1234 1765
rect 1318 1731 1330 1765
rect 1222 1725 1330 1731
rect 1240 1602 1246 1662
rect 1306 1602 1312 1662
rect 1110 1478 1116 1538
rect 1176 1478 1182 1538
rect 1246 1425 1306 1602
rect 964 1419 1072 1425
rect 964 1385 976 1419
rect 1060 1385 1072 1419
rect 964 1379 1072 1385
rect 1222 1419 1330 1425
rect 1222 1385 1234 1419
rect 1318 1385 1330 1419
rect 1222 1379 1330 1385
rect 856 1292 872 1326
rect 448 1091 556 1097
rect 448 1057 460 1091
rect 544 1057 556 1091
rect 448 1051 556 1057
rect 474 988 534 1051
rect 598 988 658 1150
rect 866 1150 872 1292
rect 906 1292 916 1326
rect 1124 1326 1170 1338
rect 906 1150 912 1292
rect 1124 1186 1130 1326
rect 866 1138 912 1150
rect 1114 1150 1130 1186
rect 1164 1186 1170 1326
rect 1374 1326 1434 1824
rect 1632 2000 1692 2258
rect 1996 2146 2002 2206
rect 2062 2146 2068 2206
rect 1738 2093 1846 2099
rect 1738 2059 1750 2093
rect 1834 2059 1846 2093
rect 1738 2053 1846 2059
rect 1632 1824 1646 2000
rect 1680 1824 1692 2000
rect 1898 2000 1944 2012
rect 1898 1872 1904 2000
rect 1480 1765 1588 1771
rect 1480 1731 1492 1765
rect 1576 1731 1588 1765
rect 1480 1725 1588 1731
rect 1500 1662 1560 1725
rect 1632 1662 1692 1824
rect 1892 1824 1904 1872
rect 1938 1872 1944 2000
rect 1938 1824 1952 1872
rect 1738 1765 1846 1771
rect 1738 1731 1750 1765
rect 1834 1731 1846 1765
rect 1738 1725 1846 1731
rect 1762 1662 1822 1725
rect 1892 1662 1952 1824
rect 1494 1602 1500 1662
rect 1560 1602 1566 1662
rect 1632 1602 1952 1662
rect 1624 1478 1630 1538
rect 1690 1478 1950 1538
rect 1480 1419 1588 1425
rect 1480 1385 1492 1419
rect 1576 1385 1588 1419
rect 1480 1379 1588 1385
rect 1374 1310 1388 1326
rect 1164 1150 1174 1186
rect 706 1091 814 1097
rect 706 1057 718 1091
rect 802 1057 814 1091
rect 706 1051 814 1057
rect 964 1091 1072 1097
rect 964 1057 976 1091
rect 1060 1057 1072 1091
rect 964 1051 1072 1057
rect 342 928 658 988
rect 728 986 788 1051
rect 722 926 728 986
rect 788 926 794 986
rect 1114 874 1174 1150
rect 1382 1150 1388 1310
rect 1422 1310 1434 1326
rect 1630 1326 1690 1478
rect 1762 1425 1822 1478
rect 1738 1419 1846 1425
rect 1738 1385 1750 1419
rect 1834 1385 1846 1419
rect 1738 1379 1846 1385
rect 1422 1150 1428 1310
rect 1630 1300 1646 1326
rect 1382 1138 1428 1150
rect 1640 1150 1646 1300
rect 1680 1300 1690 1326
rect 1890 1326 1950 1478
rect 1680 1150 1686 1300
rect 1890 1288 1904 1326
rect 1640 1138 1686 1150
rect 1898 1150 1904 1288
rect 1938 1288 1950 1326
rect 1938 1150 1944 1288
rect 1898 1138 1944 1150
rect 1222 1091 1330 1097
rect 1222 1057 1234 1091
rect 1318 1057 1330 1091
rect 1222 1051 1330 1057
rect 1480 1091 1588 1097
rect 1480 1057 1492 1091
rect 1576 1057 1588 1091
rect 1480 1051 1588 1057
rect 1738 1091 1846 1097
rect 1738 1057 1750 1091
rect 1834 1057 1846 1091
rect 1738 1051 1846 1057
rect 1502 986 1562 1051
rect 2002 986 2062 2146
rect 2304 1926 2364 2430
rect 2426 2094 2432 2154
rect 2492 2094 2498 2154
rect 2432 2025 2492 2094
rect 2408 2019 2516 2025
rect 2408 1985 2420 2019
rect 2504 1985 2516 2019
rect 2408 1979 2516 1985
rect 2304 1888 2316 1926
rect 2310 1150 2316 1888
rect 2350 1888 2364 1926
rect 2568 1926 2614 1938
rect 2350 1150 2356 1888
rect 2568 1196 2574 1926
rect 2310 1138 2356 1150
rect 2556 1150 2574 1196
rect 2608 1196 2614 1926
rect 2608 1150 2616 1196
rect 2408 1091 2516 1097
rect 2408 1057 2420 1091
rect 2504 1057 2516 1091
rect 2408 1051 2516 1057
rect 1496 926 1502 986
rect 1562 926 1568 986
rect 1996 926 2002 986
rect 2062 926 2068 986
rect 2432 984 2492 1051
rect 2556 976 2616 1150
rect 2432 918 2492 924
rect 2550 916 2556 976
rect 2616 916 2622 976
rect 210 814 216 874
rect 276 814 282 874
rect 1108 814 1114 874
rect 1174 814 1180 874
rect 3216 833 3222 2907
rect 3322 833 3328 2907
rect -724 800 -664 806
rect 3216 724 3328 833
rect -3328 718 3328 724
rect -3328 618 -3222 718
rect 3222 618 3328 718
rect -3328 612 3328 618
rect -3328 382 3328 388
rect -3328 282 -3222 382
rect 3222 282 3328 382
rect -3328 276 3328 282
rect -3328 97 -3216 276
rect -3328 -3237 -3322 97
rect -3222 -3237 -3216 97
rect -3128 182 -72 188
rect -3128 82 -3022 182
rect -178 82 -72 182
rect -3128 76 -72 82
rect -3128 28 -3016 76
rect -3128 -948 -3122 28
rect -3022 -948 -3016 28
rect -184 28 -72 76
rect -2112 -46 -2106 14
rect -2046 -46 -2040 14
rect -1078 -46 -1072 14
rect -1012 -46 -1006 14
rect -2628 -162 -2622 -102
rect -2562 -162 -2556 -102
rect -2622 -220 -2562 -162
rect -2876 -280 -2562 -220
rect -2496 -280 -2490 -220
rect -2430 -280 -2424 -220
rect -2876 -434 -2816 -280
rect -2750 -344 -2690 -280
rect -2772 -350 -2664 -344
rect -2772 -384 -2760 -350
rect -2676 -384 -2664 -350
rect -2772 -390 -2664 -384
rect -2876 -462 -2864 -434
rect -2870 -610 -2864 -462
rect -2830 -462 -2816 -434
rect -2622 -434 -2562 -280
rect -2490 -344 -2430 -280
rect -2514 -350 -2406 -344
rect -2514 -384 -2502 -350
rect -2418 -384 -2406 -350
rect -2514 -390 -2406 -384
rect -2256 -350 -2148 -344
rect -2256 -384 -2244 -350
rect -2160 -384 -2148 -350
rect -2256 -390 -2148 -384
rect -2830 -610 -2824 -462
rect -2622 -486 -2606 -434
rect -2870 -622 -2824 -610
rect -2612 -610 -2606 -486
rect -2572 -486 -2562 -434
rect -2354 -434 -2308 -422
rect -2572 -610 -2566 -486
rect -2354 -580 -2348 -434
rect -2612 -622 -2566 -610
rect -2362 -610 -2348 -580
rect -2314 -580 -2308 -434
rect -2106 -434 -2046 -46
rect -1592 -162 -1586 -102
rect -1526 -162 -1520 -102
rect -1720 -280 -1714 -220
rect -1654 -280 -1648 -220
rect -1714 -344 -1654 -280
rect -1998 -350 -1890 -344
rect -1998 -384 -1986 -350
rect -1902 -384 -1890 -350
rect -1998 -390 -1890 -384
rect -1740 -350 -1632 -344
rect -1740 -384 -1728 -350
rect -1644 -384 -1632 -350
rect -1740 -390 -1632 -384
rect -2106 -474 -2090 -434
rect -2314 -610 -2302 -580
rect -2772 -660 -2664 -654
rect -2772 -694 -2760 -660
rect -2676 -694 -2664 -660
rect -2772 -700 -2664 -694
rect -2514 -660 -2406 -654
rect -2514 -694 -2502 -660
rect -2418 -694 -2406 -660
rect -2514 -700 -2406 -694
rect -2362 -874 -2302 -610
rect -2096 -610 -2090 -474
rect -2056 -474 -2046 -434
rect -1838 -434 -1792 -422
rect -2056 -610 -2050 -474
rect -1838 -570 -1832 -434
rect -2096 -622 -2050 -610
rect -1846 -610 -1832 -570
rect -1798 -570 -1792 -434
rect -1586 -434 -1526 -162
rect -1466 -280 -1460 -220
rect -1400 -280 -1394 -220
rect -1460 -344 -1400 -280
rect -1482 -350 -1374 -344
rect -1482 -384 -1470 -350
rect -1386 -384 -1374 -350
rect -1482 -390 -1374 -384
rect -1224 -350 -1116 -344
rect -1224 -384 -1212 -350
rect -1128 -384 -1116 -350
rect -1224 -390 -1116 -384
rect -1586 -474 -1574 -434
rect -1798 -610 -1786 -570
rect -2256 -660 -2148 -654
rect -2256 -694 -2244 -660
rect -2160 -694 -2148 -660
rect -2256 -700 -2148 -694
rect -1998 -660 -1890 -654
rect -1998 -694 -1986 -660
rect -1902 -694 -1890 -660
rect -1998 -700 -1890 -694
rect -2230 -756 -2170 -700
rect -1974 -756 -1914 -700
rect -2236 -816 -2230 -756
rect -2170 -816 -2164 -756
rect -1980 -816 -1974 -756
rect -1914 -816 -1908 -756
rect -1846 -874 -1786 -610
rect -1580 -610 -1574 -474
rect -1540 -474 -1526 -434
rect -1322 -434 -1276 -422
rect -1540 -610 -1534 -474
rect -1322 -580 -1316 -434
rect -1580 -622 -1534 -610
rect -1326 -610 -1316 -580
rect -1282 -580 -1276 -434
rect -1072 -434 -1012 -46
rect -562 -162 -556 -102
rect -496 -162 -490 -102
rect -556 -220 -496 -162
rect -686 -280 -680 -220
rect -620 -280 -614 -220
rect -556 -280 -236 -220
rect -680 -344 -620 -280
rect -966 -350 -858 -344
rect -966 -384 -954 -350
rect -870 -384 -858 -350
rect -966 -390 -858 -384
rect -708 -350 -600 -344
rect -708 -384 -696 -350
rect -612 -384 -600 -350
rect -708 -390 -600 -384
rect -1072 -472 -1058 -434
rect -1282 -610 -1266 -580
rect -1740 -660 -1632 -654
rect -1740 -694 -1728 -660
rect -1644 -694 -1632 -660
rect -1740 -700 -1632 -694
rect -1482 -660 -1374 -654
rect -1482 -694 -1470 -660
rect -1386 -694 -1374 -660
rect -1482 -700 -1374 -694
rect -1326 -874 -1266 -610
rect -1064 -610 -1058 -472
rect -1024 -472 -1012 -434
rect -806 -434 -760 -422
rect -1024 -610 -1018 -472
rect -806 -576 -800 -434
rect -1064 -622 -1018 -610
rect -814 -610 -800 -576
rect -766 -576 -760 -434
rect -556 -434 -496 -280
rect -426 -344 -366 -280
rect -450 -350 -342 -344
rect -450 -384 -438 -350
rect -354 -384 -342 -350
rect -450 -390 -342 -384
rect -556 -480 -542 -434
rect -766 -610 -754 -576
rect -1224 -660 -1116 -654
rect -1224 -694 -1212 -660
rect -1128 -694 -1116 -660
rect -1224 -700 -1116 -694
rect -966 -660 -858 -654
rect -966 -694 -954 -660
rect -870 -694 -858 -660
rect -966 -700 -858 -694
rect -1200 -756 -1140 -700
rect -942 -756 -882 -700
rect -1206 -816 -1200 -756
rect -1140 -816 -1134 -756
rect -948 -816 -942 -756
rect -882 -816 -876 -756
rect -814 -874 -754 -610
rect -548 -610 -542 -480
rect -508 -480 -496 -434
rect -296 -434 -236 -280
rect -296 -480 -284 -434
rect -508 -610 -502 -480
rect -548 -622 -502 -610
rect -290 -610 -284 -480
rect -250 -480 -236 -434
rect -250 -610 -244 -480
rect -290 -622 -244 -610
rect -708 -660 -600 -654
rect -708 -694 -696 -660
rect -612 -694 -600 -660
rect -708 -700 -600 -694
rect -450 -660 -342 -654
rect -450 -694 -438 -660
rect -354 -694 -342 -660
rect -450 -700 -342 -694
rect -2368 -934 -2362 -874
rect -2302 -934 -2296 -874
rect -1852 -934 -1846 -874
rect -1786 -934 -1780 -874
rect -1332 -934 -1326 -874
rect -1266 -934 -1260 -874
rect -820 -934 -814 -874
rect -754 -934 -748 -874
rect -3128 -996 -3016 -948
rect -184 -948 -178 28
rect -78 -948 -72 28
rect 3216 97 3328 276
rect 1114 -66 1174 -60
rect 2426 -124 2432 -64
rect 2492 -124 2498 -64
rect 2556 -72 2616 -66
rect 1114 -182 1174 -126
rect 726 -242 1560 -182
rect 726 -306 786 -242
rect 988 -306 1048 -242
rect 446 -312 554 -306
rect 446 -346 458 -312
rect 542 -346 554 -312
rect 446 -352 554 -346
rect 704 -312 812 -306
rect 704 -346 716 -312
rect 800 -346 812 -312
rect 704 -352 812 -346
rect 962 -312 1070 -306
rect 962 -346 974 -312
rect 1058 -346 1070 -312
rect 962 -352 1070 -346
rect 348 -396 394 -384
rect 348 -542 354 -396
rect 344 -572 354 -542
rect 388 -542 394 -396
rect 606 -396 652 -384
rect 606 -524 612 -396
rect 388 -572 404 -542
rect 344 -702 404 -572
rect 596 -572 612 -524
rect 646 -524 652 -396
rect 864 -396 910 -384
rect 646 -572 656 -524
rect 864 -526 870 -396
rect 446 -622 554 -616
rect 446 -656 458 -622
rect 542 -656 554 -622
rect 446 -662 554 -656
rect 470 -702 530 -662
rect 596 -702 656 -572
rect 854 -572 870 -526
rect 904 -526 910 -396
rect 1114 -396 1174 -242
rect 1242 -306 1302 -242
rect 1500 -306 1560 -242
rect 2432 -280 2492 -124
rect 2408 -286 2516 -280
rect 1220 -312 1328 -306
rect 1220 -346 1232 -312
rect 1316 -346 1328 -312
rect 1220 -352 1328 -346
rect 1478 -312 1586 -306
rect 1478 -346 1490 -312
rect 1574 -346 1586 -312
rect 1478 -352 1586 -346
rect 1736 -312 1844 -306
rect 1736 -346 1748 -312
rect 1832 -346 1844 -312
rect 2408 -320 2420 -286
rect 2504 -320 2516 -286
rect 2408 -326 2516 -320
rect 1736 -352 1844 -346
rect 2310 -370 2356 -358
rect 904 -572 914 -526
rect 1114 -558 1128 -396
rect 704 -622 812 -616
rect 704 -656 716 -622
rect 800 -656 812 -622
rect 704 -662 812 -656
rect 344 -762 596 -702
rect 656 -762 662 -702
rect -184 -996 -72 -948
rect -3128 -1002 -72 -996
rect -3128 -1102 -3022 -1002
rect -178 -1102 -72 -1002
rect -3128 -1108 -72 -1102
rect 854 -850 914 -572
rect 1122 -572 1128 -558
rect 1162 -558 1174 -396
rect 1380 -396 1426 -384
rect 1380 -526 1386 -396
rect 1162 -572 1168 -558
rect 1122 -584 1168 -572
rect 1370 -572 1386 -526
rect 1420 -526 1426 -396
rect 1638 -396 1684 -384
rect 1420 -572 1430 -526
rect 1638 -530 1644 -396
rect 962 -622 1070 -616
rect 962 -656 974 -622
rect 1058 -656 1070 -622
rect 962 -662 1070 -656
rect 1220 -622 1328 -616
rect 1220 -656 1232 -622
rect 1316 -656 1328 -622
rect 1220 -662 1328 -656
rect 1370 -850 1430 -572
rect 1630 -572 1644 -530
rect 1678 -530 1684 -396
rect 1896 -396 1942 -384
rect 1678 -572 1690 -530
rect 1896 -546 1902 -396
rect 1478 -622 1586 -616
rect 1478 -656 1490 -622
rect 1574 -656 1586 -622
rect 1478 -662 1586 -656
rect 1630 -702 1690 -572
rect 1888 -572 1902 -546
rect 1936 -546 1942 -396
rect 1936 -572 1948 -546
rect 1736 -622 1844 -616
rect 1736 -656 1748 -622
rect 1832 -656 1844 -622
rect 1736 -662 1844 -656
rect 1760 -702 1820 -662
rect 1888 -702 1948 -572
rect 2310 -690 2316 -370
rect 1624 -762 1630 -702
rect 1690 -762 1948 -702
rect 2296 -746 2316 -690
rect 2350 -746 2356 -370
rect 2556 -370 2616 -132
rect 2556 -422 2574 -370
rect 2296 -850 2356 -746
rect 2568 -746 2574 -422
rect 2608 -422 2616 -370
rect 2608 -746 2614 -422
rect 2568 -758 2614 -746
rect 2408 -796 2516 -790
rect 2408 -830 2420 -796
rect 2504 -830 2516 -796
rect 2408 -836 2516 -830
rect 854 -910 2356 -850
rect 2432 -888 2492 -836
rect 854 -1212 914 -910
rect 2296 -1212 2356 -910
rect 2426 -948 2432 -888
rect 2492 -948 2498 -888
rect -3128 -1218 3128 -1212
rect -3128 -1318 -3022 -1218
rect 3022 -1318 3128 -1218
rect -3128 -1324 3128 -1318
rect -3128 -1384 -3016 -1324
rect -3128 -2576 -3122 -1384
rect -3022 -2576 -3016 -1384
rect -2728 -1468 -2722 -1408
rect -2662 -1468 -2656 -1408
rect -2722 -2356 -2662 -1468
rect -2576 -1489 -1660 -1429
rect -1302 -1468 -1296 -1408
rect -1236 -1468 -1230 -1408
rect -434 -1468 -428 -1408
rect -368 -1468 -362 -1408
rect -8 -1468 -2 -1408
rect 58 -1468 64 -1408
rect 418 -1468 424 -1408
rect 484 -1468 490 -1408
rect -2576 -1627 -2516 -1489
rect -2138 -1537 -2078 -1489
rect -2321 -1543 -1913 -1537
rect -2321 -1577 -2309 -1543
rect -1925 -1577 -1913 -1543
rect -2321 -1583 -1913 -1577
rect -2576 -1672 -2563 -1627
rect -2569 -1742 -2563 -1672
rect -2582 -1803 -2563 -1742
rect -2529 -1672 -2516 -1627
rect -1720 -1627 -1660 -1489
rect -1296 -1537 -1236 -1468
rect -428 -1537 -368 -1468
rect -1463 -1543 -1055 -1537
rect -1463 -1577 -1451 -1543
rect -1067 -1577 -1055 -1543
rect -1463 -1583 -1055 -1577
rect -605 -1543 -197 -1537
rect -605 -1577 -593 -1543
rect -209 -1577 -197 -1543
rect -605 -1583 -197 -1577
rect -1296 -1588 -1236 -1583
rect -2529 -1742 -2523 -1672
rect -1720 -1676 -1705 -1627
rect -2529 -1803 -2522 -1742
rect -2582 -1892 -2522 -1803
rect -1711 -1803 -1705 -1676
rect -1671 -1676 -1660 -1627
rect -853 -1627 -807 -1615
rect -1671 -1803 -1665 -1676
rect -853 -1765 -847 -1627
rect -1711 -1815 -1665 -1803
rect -860 -1803 -847 -1765
rect -813 -1765 -807 -1627
rect -2 -1627 58 -1468
rect 424 -1537 484 -1468
rect 253 -1543 661 -1537
rect 253 -1577 265 -1543
rect 649 -1577 661 -1543
rect 253 -1583 661 -1577
rect 424 -1586 484 -1583
rect -2 -1674 11 -1627
rect -813 -1803 -800 -1765
rect -2321 -1853 -1913 -1847
rect -2321 -1887 -2309 -1853
rect -1925 -1887 -1913 -1853
rect -2588 -1952 -2582 -1892
rect -2522 -1952 -2516 -1892
rect -2321 -1893 -1913 -1887
rect -1463 -1853 -1055 -1847
rect -1463 -1887 -1451 -1853
rect -1067 -1887 -1055 -1853
rect -1463 -1893 -1055 -1887
rect -1286 -1955 -1226 -1893
rect -2321 -1961 -1913 -1955
rect -2321 -1995 -2309 -1961
rect -1925 -1995 -1913 -1961
rect -2321 -2001 -1913 -1995
rect -1463 -1961 -1055 -1955
rect -1463 -1995 -1451 -1961
rect -1067 -1995 -1055 -1961
rect -1463 -2001 -1055 -1995
rect -2569 -2045 -2523 -2033
rect -2569 -2160 -2563 -2045
rect -2576 -2221 -2563 -2160
rect -2529 -2160 -2523 -2045
rect -1711 -2045 -1665 -2033
rect -2529 -2221 -2516 -2160
rect -1711 -2166 -1705 -2045
rect -2576 -2356 -2516 -2221
rect -1720 -2221 -1705 -2166
rect -1671 -2166 -1665 -2045
rect -860 -2045 -800 -1803
rect 5 -1803 11 -1674
rect 45 -1674 58 -1627
rect 854 -1627 914 -1324
rect 3016 -1384 3128 -1324
rect 1290 -1468 1296 -1408
rect 1356 -1468 1362 -1408
rect 1296 -1537 1356 -1468
rect 1712 -1489 2768 -1429
rect 1111 -1543 1519 -1537
rect 1111 -1577 1123 -1543
rect 1507 -1577 1519 -1543
rect 1111 -1583 1519 -1577
rect 45 -1803 51 -1674
rect 854 -1680 869 -1627
rect 863 -1761 869 -1680
rect 5 -1815 51 -1803
rect 852 -1803 869 -1761
rect 903 -1680 914 -1627
rect 1712 -1627 1772 -1489
rect 2132 -1537 2192 -1489
rect 1969 -1543 2377 -1537
rect 1969 -1577 1981 -1543
rect 2365 -1577 2377 -1543
rect 1969 -1583 2377 -1577
rect 1712 -1660 1727 -1627
rect 903 -1761 909 -1680
rect 903 -1803 912 -1761
rect -605 -1853 -197 -1847
rect -605 -1887 -593 -1853
rect -209 -1887 -197 -1853
rect -605 -1893 -197 -1887
rect 253 -1853 661 -1847
rect 253 -1887 265 -1853
rect 649 -1887 661 -1853
rect 253 -1893 661 -1887
rect -424 -1955 -364 -1893
rect 432 -1955 492 -1893
rect -605 -1961 -197 -1955
rect -605 -1995 -593 -1961
rect -209 -1995 -197 -1961
rect -605 -2001 -197 -1995
rect 253 -1961 661 -1955
rect 253 -1995 265 -1961
rect 649 -1995 661 -1961
rect 253 -2001 661 -1995
rect -1671 -2221 -1660 -2166
rect -2321 -2271 -1913 -2265
rect -2321 -2305 -2309 -2271
rect -1925 -2305 -1913 -2271
rect -2321 -2311 -1913 -2305
rect -2138 -2356 -2078 -2311
rect -1720 -2356 -1660 -2221
rect -860 -2221 -847 -2045
rect -813 -2221 -800 -2045
rect 5 -2045 51 -2033
rect 5 -2178 11 -2045
rect -1463 -2271 -1055 -2265
rect -1463 -2305 -1451 -2271
rect -1067 -2305 -1055 -2271
rect -1463 -2311 -1055 -2305
rect -2722 -2416 -1660 -2356
rect -860 -2372 -800 -2221
rect -2 -2221 11 -2178
rect 45 -2178 51 -2045
rect 852 -2045 912 -1803
rect 1721 -1803 1727 -1660
rect 1761 -1660 1772 -1627
rect 2568 -1627 2628 -1489
rect 1761 -1803 1767 -1660
rect 2568 -1694 2585 -1627
rect 1721 -1815 1767 -1803
rect 2579 -1803 2585 -1694
rect 2619 -1694 2628 -1627
rect 2619 -1803 2625 -1694
rect 2579 -1815 2625 -1803
rect 1111 -1853 1519 -1847
rect 1111 -1887 1123 -1853
rect 1507 -1887 1519 -1853
rect 1111 -1893 1519 -1887
rect 1969 -1853 2377 -1847
rect 1969 -1887 1981 -1853
rect 2365 -1887 2377 -1853
rect 1969 -1893 2377 -1887
rect 1284 -1955 1344 -1893
rect 1111 -1961 1519 -1955
rect 1111 -1995 1123 -1961
rect 1507 -1995 1519 -1961
rect 1111 -2001 1519 -1995
rect 1969 -1961 2377 -1955
rect 2562 -1958 2568 -1898
rect 2628 -1958 2634 -1898
rect 1969 -1995 1981 -1961
rect 2365 -1995 2377 -1961
rect 1969 -2001 2377 -1995
rect 1284 -2002 1344 -2001
rect 852 -2088 869 -2045
rect 863 -2162 869 -2088
rect 45 -2221 58 -2178
rect -605 -2271 -197 -2265
rect -605 -2305 -593 -2271
rect -209 -2305 -197 -2271
rect -605 -2311 -197 -2305
rect -866 -2432 -860 -2372
rect -800 -2432 -794 -2372
rect -3128 -2636 -3016 -2576
rect -860 -2636 -800 -2432
rect -2 -2486 58 -2221
rect 850 -2221 869 -2162
rect 903 -2088 912 -2045
rect 1721 -2045 1767 -2033
rect 903 -2162 909 -2088
rect 1721 -2160 1727 -2045
rect 903 -2221 910 -2162
rect 253 -2271 661 -2265
rect 253 -2305 265 -2271
rect 649 -2305 661 -2271
rect 253 -2311 661 -2305
rect 850 -2372 910 -2221
rect 1712 -2221 1727 -2160
rect 1761 -2160 1767 -2045
rect 2568 -2045 2628 -1958
rect 1761 -2221 1772 -2160
rect 1111 -2271 1519 -2265
rect 1111 -2305 1123 -2271
rect 1507 -2305 1519 -2271
rect 1111 -2311 1519 -2305
rect 1712 -2356 1772 -2221
rect 2568 -2221 2585 -2045
rect 2619 -2221 2628 -2045
rect 1969 -2271 2377 -2265
rect 1969 -2305 1981 -2271
rect 2365 -2305 2377 -2271
rect 1969 -2311 2377 -2305
rect 2150 -2356 2210 -2311
rect 2568 -2356 2628 -2221
rect 844 -2432 850 -2372
rect 910 -2432 916 -2372
rect 1712 -2416 2628 -2356
rect -8 -2546 -2 -2486
rect 58 -2546 64 -2486
rect 850 -2636 910 -2432
rect 2708 -2486 2768 -1489
rect 2702 -2546 2708 -2486
rect 2768 -2546 2774 -2486
rect 3016 -2576 3022 -1384
rect 3122 -2576 3128 -1384
rect 3016 -2636 3128 -2576
rect -3128 -2642 3128 -2636
rect -3128 -2742 -3022 -2642
rect 3022 -2742 3128 -2642
rect -3128 -2748 3128 -2742
rect -860 -2836 -800 -2748
rect 850 -2836 910 -2748
rect -928 -2864 970 -2836
rect -928 -2974 -898 -2864
rect 942 -2974 970 -2864
rect -928 -3002 970 -2974
rect -3328 -3416 -3216 -3237
rect -2616 -3416 -2606 -3116
rect 2606 -3416 2616 -3116
rect 3216 -3237 3222 97
rect 3322 -3237 3328 97
rect 3216 -3416 3328 -3237
rect -3328 -3422 3328 -3416
rect -3328 -3522 -3222 -3422
rect 3222 -3522 3328 -3422
rect -3328 -3528 3328 -3522
<< via1 >>
rect -3216 2716 -2616 3016
rect 2616 2716 3216 3016
rect -2646 2456 2544 2528
rect -2776 2146 -2716 2206
rect -2266 2146 -2206 2206
rect -1622 2146 -1562 2206
rect -1496 2146 -1436 2206
rect -2270 1604 -2210 1664
rect -2138 1470 -2078 1530
rect -2008 1470 -1948 1530
rect -1232 2146 -1172 2206
rect -1494 1604 -1434 1664
rect -1750 1470 -1690 1530
rect -1628 1470 -1568 1530
rect -596 2146 -536 2206
rect -464 2146 -404 2206
rect -1240 1604 -1180 1664
rect -1112 1470 -1052 1530
rect -980 1470 -920 1530
rect -464 1604 -404 1664
rect -720 1470 -660 1530
rect -596 1470 -536 1530
rect -2776 918 -2716 978
rect -2274 918 -2214 978
rect -2142 918 -2082 978
rect 216 2258 276 2318
rect 600 2258 660 2318
rect -1500 918 -1440 978
rect -1240 918 -1180 978
rect -1108 918 -1048 978
rect -2014 814 -1954 874
rect -464 918 -404 978
rect 988 2146 1048 2206
rect 1244 2146 1304 2206
rect 730 1602 790 1662
rect 598 1478 658 1538
rect 1632 2258 1692 2318
rect 988 1602 1048 1662
rect 1246 1602 1306 1662
rect 1116 1478 1176 1538
rect 2002 2146 2062 2206
rect 1500 1602 1560 1662
rect 1630 1478 1690 1538
rect 728 926 788 986
rect 2432 2094 2492 2154
rect 1502 926 1562 986
rect 2002 926 2062 986
rect 2432 924 2492 984
rect 2556 916 2616 976
rect -724 806 -664 866
rect 216 814 276 874
rect 1114 814 1174 874
rect -2106 -46 -2046 14
rect -1072 -46 -1012 14
rect -2622 -162 -2562 -102
rect -2490 -280 -2430 -220
rect -1586 -162 -1526 -102
rect -1714 -280 -1654 -220
rect -1460 -280 -1400 -220
rect -2230 -816 -2170 -756
rect -1974 -816 -1914 -756
rect -556 -162 -496 -102
rect -680 -280 -620 -220
rect -1200 -816 -1140 -756
rect -942 -816 -882 -756
rect -2362 -934 -2302 -874
rect -1846 -934 -1786 -874
rect -1326 -934 -1266 -874
rect -814 -934 -754 -874
rect 1114 -126 1174 -66
rect 2432 -124 2492 -64
rect 2556 -132 2616 -72
rect 596 -762 656 -702
rect 1630 -762 1690 -702
rect 2432 -948 2492 -888
rect -2722 -1468 -2662 -1408
rect -1296 -1468 -1236 -1408
rect -428 -1468 -368 -1408
rect -2 -1468 58 -1408
rect 424 -1468 484 -1408
rect -2582 -1952 -2522 -1892
rect 1296 -1468 1356 -1408
rect 2568 -1958 2628 -1898
rect -860 -2432 -800 -2372
rect 850 -2432 910 -2372
rect -2 -2546 58 -2486
rect 2708 -2546 2768 -2486
rect -898 -2974 942 -2864
rect -3216 -3416 -2616 -3116
rect 2616 -3416 3216 -3116
<< metal2 >>
rect -3216 3016 -2616 3026
rect -3216 2706 -2616 2716
rect 2616 3016 3216 3026
rect 2616 2706 3216 2716
rect -2674 2528 2566 2562
rect -2674 2456 -2646 2528
rect 2544 2456 2566 2528
rect -2674 2430 2566 2456
rect 216 2318 276 2324
rect 600 2318 660 2324
rect 1632 2318 1692 2324
rect 276 2258 600 2318
rect 660 2258 1632 2318
rect 216 2252 276 2258
rect 600 2252 660 2258
rect 1632 2252 1692 2258
rect -2776 2206 -2716 2212
rect -2266 2206 -2206 2212
rect -1622 2206 -1562 2212
rect -1496 2206 -1436 2212
rect -1232 2206 -1172 2212
rect -596 2206 -536 2212
rect -464 2206 -404 2212
rect 988 2206 1048 2212
rect 1244 2206 1304 2212
rect 2002 2206 2062 2212
rect -2716 2146 -2266 2206
rect -2206 2146 -1622 2206
rect -1562 2146 -1496 2206
rect -1436 2146 -1232 2206
rect -1172 2146 -596 2206
rect -536 2146 -464 2206
rect -404 2146 988 2206
rect 1048 2146 1244 2206
rect 1304 2146 2002 2206
rect 2432 2154 2492 2160
rect -2776 2140 -2716 2146
rect -2266 2140 -2206 2146
rect -1622 2140 -1562 2146
rect -1496 2140 -1436 2146
rect -1232 2140 -1172 2146
rect -596 2140 -536 2146
rect -464 2140 -404 2146
rect 988 2140 1048 2146
rect 1244 2140 1304 2146
rect 2002 2140 2062 2146
rect 2132 2094 2432 2154
rect -2270 1664 -2210 1670
rect -1494 1664 -1434 1670
rect -1240 1664 -1180 1670
rect -464 1664 -404 1670
rect -2210 1604 -1494 1664
rect -1434 1604 -1240 1664
rect -1180 1604 -464 1664
rect 730 1662 790 1668
rect 988 1662 1048 1668
rect 1246 1662 1306 1668
rect 1500 1662 1560 1668
rect -2270 1598 -2210 1604
rect -1494 1598 -1434 1604
rect -1240 1598 -1180 1604
rect -464 1598 -404 1604
rect 72 1602 730 1662
rect 790 1602 988 1662
rect 1048 1602 1246 1662
rect 1306 1602 1500 1662
rect -2138 1530 -2078 1536
rect -2008 1530 -1948 1536
rect -1750 1530 -1690 1536
rect -1628 1530 -1568 1536
rect -1112 1530 -1052 1536
rect -980 1530 -920 1536
rect -720 1530 -660 1536
rect -596 1530 -536 1536
rect 72 1530 132 1602
rect 730 1596 790 1602
rect 988 1596 1048 1602
rect 1246 1596 1306 1602
rect 1500 1596 1560 1602
rect -2078 1470 -2008 1530
rect -1948 1470 -1750 1530
rect -1690 1470 -1628 1530
rect -1568 1470 -1112 1530
rect -1052 1470 -980 1530
rect -920 1470 -720 1530
rect -660 1470 -596 1530
rect -536 1470 132 1530
rect 598 1538 658 1544
rect 1116 1538 1176 1544
rect 1630 1538 1690 1544
rect 2132 1538 2192 2094
rect 2432 2088 2492 2094
rect 658 1478 1116 1538
rect 1176 1478 1630 1538
rect 1690 1478 2192 1538
rect 598 1472 658 1478
rect 1116 1472 1176 1478
rect 1630 1472 1690 1478
rect -2138 1464 -2078 1470
rect -2008 1464 -1948 1470
rect -1750 1464 -1690 1470
rect -1628 1464 -1568 1470
rect -1112 1464 -1052 1470
rect -980 1464 -920 1470
rect -720 1464 -660 1470
rect -596 1464 -536 1470
rect 728 986 788 992
rect 1502 986 1562 992
rect 2002 986 2062 992
rect -2776 978 -2716 984
rect -2274 978 -2214 984
rect -2142 978 -2082 984
rect -1500 978 -1440 984
rect -1240 978 -1180 984
rect -1108 978 -1048 984
rect -464 978 -404 984
rect -2716 918 -2274 978
rect -2214 918 -2142 978
rect -2082 918 -1500 978
rect -1440 918 -1240 978
rect -1180 918 -1108 978
rect -1048 918 -464 978
rect 788 926 1502 986
rect 1562 926 2002 986
rect 728 920 788 926
rect 1502 920 1562 926
rect 2002 920 2062 926
rect -2776 912 -2716 918
rect -2274 912 -2214 918
rect -2142 912 -2082 918
rect -2014 874 -1954 880
rect -2014 534 -1954 814
rect -2234 474 -1954 534
rect -2622 -102 -2562 -96
rect -2234 -102 -2174 474
rect -2106 14 -2046 20
rect -1748 14 -1688 918
rect -1500 912 -1440 918
rect -1370 14 -1310 918
rect -1240 912 -1180 918
rect -1108 912 -1048 918
rect -464 912 -404 918
rect 216 874 276 880
rect 1114 874 1174 880
rect -730 806 -724 866
rect -664 806 -658 866
rect 276 814 1114 874
rect 216 808 276 814
rect -1072 14 -1012 20
rect -2046 -46 -1072 14
rect -2106 -52 -2046 -46
rect -1072 -52 -1012 -46
rect -1586 -102 -1526 -96
rect -724 -102 -664 806
rect 1114 -66 1174 814
rect 2132 254 2192 1478
rect 2426 924 2432 984
rect 2492 924 2498 984
rect 2556 976 2616 982
rect 2432 254 2492 924
rect 2132 194 2492 254
rect -556 -102 -496 -96
rect -2562 -162 -1586 -102
rect -1526 -162 -556 -102
rect 1108 -126 1114 -66
rect 1174 -126 1180 -66
rect -2622 -168 -2562 -162
rect -1586 -168 -1526 -162
rect -556 -168 -496 -162
rect -2490 -220 -2430 -214
rect -1714 -220 -1654 -214
rect -1460 -220 -1400 -214
rect -680 -220 -620 -214
rect -2430 -280 -1714 -220
rect -1654 -280 -1460 -220
rect -1400 -280 -680 -220
rect -2490 -286 -2430 -280
rect -1714 -286 -1654 -280
rect -1460 -286 -1400 -280
rect -680 -286 -620 -280
rect 596 -702 656 -696
rect 1630 -702 1690 -696
rect 2132 -702 2192 194
rect 2432 -64 2492 194
rect 2556 -72 2616 916
rect 2432 -130 2492 -124
rect 2550 -132 2556 -72
rect 2616 -132 2622 -72
rect -2230 -756 -2170 -750
rect -1974 -756 -1914 -750
rect -1200 -756 -1140 -750
rect -942 -756 -882 -750
rect -2170 -816 -1974 -756
rect -1914 -816 -1200 -756
rect -1140 -816 -942 -756
rect 656 -762 1630 -702
rect 1690 -762 2192 -702
rect 596 -768 656 -762
rect 1630 -768 1690 -762
rect -2230 -822 -2170 -816
rect -1974 -822 -1914 -816
rect -1200 -822 -1140 -816
rect -942 -822 -882 -816
rect -2362 -874 -2302 -868
rect -1846 -874 -1786 -868
rect -1326 -874 -1266 -868
rect -814 -874 -754 -868
rect -2852 -934 -2362 -874
rect -2302 -934 -1846 -874
rect -1786 -934 -1326 -874
rect -1266 -934 -814 -874
rect -2852 -1892 -2792 -934
rect -2362 -940 -2302 -934
rect -1846 -940 -1786 -934
rect -1326 -940 -1266 -934
rect -814 -940 -754 -934
rect 2132 -888 2192 -762
rect 2432 -888 2492 -882
rect 2132 -948 2432 -888
rect 2432 -954 2492 -948
rect -2722 -1408 -2662 -1402
rect -1296 -1408 -1236 -1402
rect -428 -1408 -368 -1402
rect -2 -1408 58 -1402
rect 424 -1408 484 -1402
rect 1296 -1408 1356 -1402
rect -2662 -1468 -1296 -1408
rect -1236 -1468 -428 -1408
rect -368 -1468 -2 -1408
rect 58 -1468 424 -1408
rect 484 -1468 1296 -1408
rect 1356 -1468 2908 -1408
rect -2722 -1474 -2662 -1468
rect -1296 -1474 -1236 -1468
rect -428 -1474 -368 -1468
rect -2 -1474 58 -1468
rect 424 -1474 484 -1468
rect 1296 -1474 1356 -1468
rect -2582 -1892 -2522 -1886
rect -2852 -1952 -2582 -1892
rect -2852 -2486 -2792 -1952
rect -2582 -1958 -2522 -1952
rect 2568 -1898 2628 -1892
rect 2848 -1898 2908 -1468
rect 2628 -1958 2908 -1898
rect 2568 -1964 2628 -1958
rect -860 -2372 -800 -2366
rect 850 -2372 910 -2366
rect -800 -2432 850 -2372
rect -860 -2438 -800 -2432
rect 850 -2438 910 -2432
rect -2 -2486 58 -2480
rect 2708 -2486 2768 -2480
rect -2852 -2546 -2 -2486
rect 58 -2546 2708 -2486
rect -2 -2552 58 -2546
rect 2708 -2552 2768 -2546
rect -928 -2864 970 -2836
rect -928 -2974 -898 -2864
rect 942 -2974 970 -2864
rect -928 -3002 970 -2974
rect -3216 -3116 -2616 -3106
rect -3216 -3426 -2616 -3416
rect 2616 -3116 3216 -3106
rect 2616 -3426 3216 -3416
<< via2 >>
rect -3216 2716 -2616 3016
rect 2616 2716 3216 3016
rect -2646 2456 2544 2528
rect -898 -2974 942 -2864
rect -3216 -3416 -2616 -3116
rect 2616 -3416 3216 -3116
<< metal3 >>
rect -3226 3016 -2606 3021
rect -3226 2716 -3216 3016
rect -2616 2716 -2606 3016
rect -3226 2711 -2606 2716
rect 2606 3016 3226 3021
rect 2606 2716 2616 3016
rect 3216 2716 3226 3016
rect 2606 2711 3226 2716
rect -2674 2528 2566 2562
rect -2674 2456 -2646 2528
rect 2544 2456 2566 2528
rect -2674 2430 2566 2456
rect -928 -2864 970 -2836
rect -928 -2974 -898 -2864
rect 942 -2974 970 -2864
rect -928 -3002 970 -2974
rect -3226 -3116 -2606 -3111
rect -3226 -3416 -3216 -3116
rect -2616 -3416 -2606 -3116
rect -3226 -3421 -2606 -3416
rect 2606 -3116 3226 -3111
rect 2606 -3416 2616 -3116
rect 3216 -3416 3226 -3116
rect 2606 -3421 3226 -3416
<< via3 >>
rect -3216 2716 -2616 3016
rect 2616 2716 3216 3016
rect -2646 2456 2544 2528
rect -898 -2974 942 -2864
rect -3216 -3416 -2616 -3116
rect 2616 -3416 3216 -3116
<< metal4 >>
rect -3400 3016 3400 3200
rect -3400 2716 -3216 3016
rect -2616 2716 2616 3016
rect 3216 2716 3400 3016
rect -3400 2528 3400 2716
rect -3400 2456 -2646 2528
rect 2544 2456 3400 2528
rect -3400 2400 3400 2456
rect -3400 -2864 3400 -2800
rect -3400 -2974 -898 -2864
rect 942 -2974 3400 -2864
rect -3400 -3116 3400 -2974
rect -3400 -3416 -3216 -3116
rect -2616 -3416 2616 -3116
rect 3216 -3416 3400 -3116
rect -3400 -3600 3400 -3416
<< labels >>
flabel metal1 886 -216 900 -202 1 FreeSans 480 0 0 0 vmirror
flabel metal1 436 -744 448 -730 1 FreeSans 480 0 0 0 vo1
flabel metal1 2726 -2168 2748 -2144 1 FreeSans 480 0 0 0 vtail
flabel metal2 -820 -1444 -780 -1426 1 FreeSans 480 0 0 0 ibiasn
port 4 n
flabel metal2 -452 -2416 -440 -2394 1 FreeSans 480 0 0 0 VSS
port 6 n ground bidirectional
flabel metal1 -2766 -264 -2732 -234 1 FreeSans 480 0 0 0 vcompm
flabel metal2 -2292 -262 -2260 -238 1 FreeSans 480 0 0 0 vip
port 1 n
flabel metal2 -1592 -802 -1560 -774 1 FreeSans 480 0 0 0 vim
port 2 n
flabel metal2 -1592 -914 -1566 -890 1 FreeSans 480 0 0 0 vtail
flabel metal2 -1654 -28 -1634 -4 1 FreeSans 480 0 0 0 vcompp
flabel metal1 2026 1582 2042 1600 1 FreeSans 480 0 0 0 vcompp
flabel metal1 1522 1686 1534 1696 1 FreeSans 480 0 0 0 vcompm
flabel metal2 1500 1502 1516 1514 1 FreeSans 480 0 0 0 vo1
flabel metal2 824 832 836 848 1 FreeSans 480 0 0 0 vmirror
flabel metal1 -2122 1544 -2104 1566 1 FreeSans 480 0 0 0 vcompm
flabel metal2 2586 472 2596 480 1 FreeSans 480 0 0 0 vo
port 3 n
flabel metal2 -720 2168 -702 2188 1 FreeSans 480 0 0 0 vcompp
flabel metal4 -1674 2724 -1612 2786 1 FreeSans 480 0 0 0 VDD
port 5 n power bidirectional
<< end >>
