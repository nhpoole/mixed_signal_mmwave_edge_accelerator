magic
tech sky130A
magscale 1 2
timestamp 1624494425
<< error_s >>
rect 38 102322 80 102331
rect 38 102305 113 102322
rect 30 102293 38 102305
rect 42 102288 76 102305
rect 79 102288 113 102305
rect 42 102209 46 102243
rect 72 102209 76 102243
rect -25 102172 25 102174
rect -8 102164 14 102171
rect -8 102163 17 102164
rect 25 102163 27 102172
rect -12 102156 38 102163
rect -12 102155 34 102156
rect -12 102151 8 102155
rect 0 102139 8 102151
rect 14 102139 34 102155
rect 0 102138 34 102139
rect 0 102131 38 102138
rect 14 102130 17 102131
rect 25 102122 27 102131
rect 42 102102 45 102192
rect 71 102161 80 102189
rect 69 102123 80 102161
rect 144 102151 148 102305
rect 151 102288 156 102322
rect 180 102291 185 102322
rect 400 102305 442 102331
rect 174 102283 246 102291
rect 256 102283 328 102291
rect 332 102289 336 102305
rect 392 102297 438 102305
rect 392 102293 408 102297
rect 400 102290 408 102293
rect 434 102290 438 102297
rect 442 102293 450 102305
rect 388 102289 454 102290
rect 224 102253 226 102269
rect 196 102245 226 102253
rect 196 102241 232 102245
rect 196 102211 204 102241
rect 216 102211 232 102241
rect 224 102164 226 102211
rect 300 102184 308 102253
rect 332 102251 342 102289
rect 400 102281 404 102289
rect 454 102275 504 102277
rect 494 102271 548 102275
rect 494 102266 514 102271
rect 504 102251 506 102266
rect 336 102239 342 102251
rect 289 102174 308 102184
rect 300 102168 308 102174
rect 332 102205 342 102239
rect 400 102243 404 102251
rect 400 102209 408 102243
rect 434 102209 438 102243
rect 498 102241 506 102251
rect 514 102241 515 102261
rect 504 102225 506 102241
rect 525 102232 528 102266
rect 547 102241 548 102261
rect 557 102241 564 102251
rect 514 102225 530 102231
rect 532 102225 548 102231
rect 332 102177 373 102205
rect 332 102171 351 102177
rect 107 102117 119 102151
rect 129 102117 149 102151
rect 196 102130 204 102164
rect 216 102130 232 102164
rect 244 102158 257 102164
rect 278 102158 291 102168
rect 244 102134 291 102158
rect 300 102158 321 102168
rect 336 102161 351 102171
rect 300 102134 329 102158
rect 332 102143 351 102161
rect 361 102171 375 102177
rect 400 102171 411 102209
rect 562 102172 612 102174
rect 361 102143 381 102171
rect 400 102143 409 102171
rect 466 102163 497 102171
rect 565 102163 596 102171
rect 442 102156 500 102163
rect 466 102155 500 102156
rect 565 102155 599 102163
rect 244 102130 257 102134
rect 42 102051 46 102085
rect 72 102051 76 102085
rect 42 102004 76 102008
rect 42 101989 46 102004
rect 72 101989 76 102004
rect 38 101971 80 101989
rect 16 101965 102 101971
rect 144 101965 148 102117
rect 174 102093 181 102121
rect 224 102083 226 102130
rect 300 102121 308 102134
rect 278 102110 305 102121
rect 332 102093 342 102143
rect 400 102123 404 102143
rect 497 102139 500 102155
rect 596 102139 599 102155
rect 466 102138 500 102139
rect 442 102131 500 102138
rect 565 102131 599 102139
rect 612 102122 614 102172
rect 256 102083 328 102091
rect 336 102085 342 102093
rect 400 102085 404 102093
rect 196 102053 204 102083
rect 216 102053 232 102083
rect 196 102049 232 102053
rect 196 102041 226 102049
rect 224 102025 226 102041
rect 332 102013 336 102081
rect 400 102051 408 102085
rect 434 102051 438 102085
rect 454 102069 504 102071
rect 504 102053 506 102069
rect 514 102063 530 102069
rect 532 102063 548 102069
rect 525 102053 548 102062
rect 400 102043 404 102051
rect 498 102043 506 102053
rect 504 102019 506 102043
rect 514 102033 515 102053
rect 525 102028 528 102053
rect 547 102033 548 102053
rect 557 102043 564 102053
rect 514 102019 548 102023
rect 400 102013 442 102014
rect 174 102003 246 102011
rect 400 102006 404 102013
rect 295 101972 300 102006
rect 324 101972 329 102006
rect 367 101989 438 102006
rect 367 101972 442 101989
rect 400 101971 442 101972
rect 378 101965 464 101971
rect 38 101949 80 101965
rect 400 101949 442 101965
rect -25 101935 25 101937
rect 42 101935 76 101949
rect 404 101935 438 101949
rect 455 101935 505 101937
rect 557 101935 607 101937
rect 16 101927 102 101935
rect 378 101927 464 101935
rect 8 101893 17 101927
rect 18 101925 51 101927
rect 80 101925 100 101927
rect 18 101893 100 101925
rect 380 101925 404 101927
rect 429 101925 438 101927
rect 442 101925 462 101927
rect 16 101885 102 101893
rect 42 101869 76 101885
rect 16 101849 38 101855
rect 42 101846 76 101850
rect 80 101849 102 101855
rect 42 101816 46 101846
rect 72 101816 76 101846
rect 42 101735 46 101769
rect 72 101735 76 101769
rect -25 101698 25 101700
rect -8 101690 14 101697
rect -8 101689 17 101690
rect 25 101689 27 101698
rect -12 101682 38 101689
rect -12 101681 34 101682
rect -12 101677 8 101681
rect 0 101665 8 101677
rect 14 101665 34 101681
rect 0 101664 34 101665
rect 0 101657 38 101664
rect 14 101656 17 101657
rect 25 101648 27 101657
rect 42 101628 45 101718
rect 69 101703 80 101735
rect 107 101703 143 101731
rect 144 101703 148 101923
rect 332 101855 336 101923
rect 380 101893 462 101925
rect 463 101893 472 101927
rect 480 101893 497 101927
rect 378 101885 464 101893
rect 505 101885 507 101935
rect 514 101893 548 101927
rect 565 101893 582 101927
rect 607 101885 609 101935
rect 404 101869 438 101885
rect 400 101855 442 101856
rect 378 101849 404 101855
rect 442 101849 464 101855
rect 400 101848 404 101849
rect 174 101809 246 101817
rect 295 101814 300 101848
rect 324 101814 329 101848
rect 224 101779 226 101795
rect 196 101771 226 101779
rect 332 101777 336 101845
rect 367 101814 438 101848
rect 400 101807 404 101814
rect 454 101801 504 101803
rect 494 101797 548 101801
rect 494 101792 514 101797
rect 504 101777 506 101792
rect 196 101767 232 101771
rect 196 101737 204 101767
rect 216 101737 232 101767
rect 400 101769 404 101777
rect 107 101697 119 101703
rect 109 101669 119 101697
rect 129 101669 149 101703
rect 174 101699 181 101729
rect 224 101690 226 101737
rect 256 101729 328 101737
rect 332 101735 336 101765
rect 400 101735 408 101769
rect 434 101735 438 101769
rect 498 101767 506 101777
rect 514 101767 515 101787
rect 504 101751 506 101767
rect 525 101758 528 101792
rect 547 101767 548 101787
rect 557 101767 564 101777
rect 514 101751 530 101757
rect 532 101751 548 101757
rect 278 101699 305 101710
rect 42 101577 46 101611
rect 72 101577 76 101611
rect 38 101539 80 101540
rect 42 101498 76 101532
rect 79 101498 113 101532
rect 42 101419 46 101453
rect 72 101419 76 101453
rect -25 101382 25 101384
rect -8 101374 14 101381
rect -8 101373 17 101374
rect 25 101373 27 101382
rect -12 101366 38 101373
rect -12 101365 34 101366
rect -12 101361 8 101365
rect 0 101349 8 101361
rect 14 101349 34 101365
rect 0 101348 34 101349
rect 0 101341 38 101348
rect 14 101340 17 101341
rect 25 101332 27 101341
rect 42 101312 45 101402
rect 71 101371 80 101399
rect 69 101333 80 101371
rect 144 101361 148 101669
rect 196 101656 204 101690
rect 216 101656 232 101690
rect 244 101686 257 101690
rect 300 101686 308 101699
rect 332 101697 342 101735
rect 400 101727 404 101735
rect 336 101687 342 101697
rect 244 101662 291 101686
rect 244 101656 257 101662
rect 224 101609 226 101656
rect 278 101652 291 101662
rect 300 101662 329 101686
rect 332 101677 342 101687
rect 400 101687 409 101715
rect 562 101698 612 101700
rect 466 101689 497 101697
rect 565 101689 596 101697
rect 300 101652 321 101662
rect 300 101646 308 101652
rect 289 101636 308 101646
rect 196 101579 204 101609
rect 216 101579 232 101609
rect 196 101575 232 101579
rect 196 101567 226 101575
rect 300 101567 308 101636
rect 332 101643 351 101677
rect 361 101649 381 101677
rect 361 101643 375 101649
rect 400 101643 411 101687
rect 442 101682 500 101689
rect 466 101681 500 101682
rect 565 101681 599 101689
rect 497 101665 500 101681
rect 596 101665 599 101681
rect 466 101664 500 101665
rect 442 101657 500 101664
rect 565 101657 599 101665
rect 612 101648 614 101698
rect 332 101619 342 101643
rect 336 101607 342 101619
rect 224 101551 226 101567
rect 332 101539 342 101607
rect 400 101611 404 101619
rect 400 101577 408 101611
rect 434 101577 438 101611
rect 454 101595 504 101597
rect 504 101579 506 101595
rect 514 101589 530 101595
rect 532 101589 548 101595
rect 525 101579 548 101588
rect 400 101569 404 101577
rect 498 101569 506 101579
rect 504 101545 506 101569
rect 514 101559 515 101579
rect 525 101554 528 101579
rect 547 101559 548 101579
rect 557 101569 564 101579
rect 514 101545 548 101549
rect 151 101498 156 101532
rect 174 101529 246 101537
rect 256 101529 328 101537
rect 336 101531 342 101539
rect 400 101534 404 101539
rect 180 101501 185 101529
rect 174 101493 246 101501
rect 256 101493 328 101501
rect 332 101499 336 101529
rect 400 101500 438 101534
rect 224 101463 226 101479
rect 196 101455 226 101463
rect 196 101451 232 101455
rect 196 101421 204 101451
rect 216 101421 232 101451
rect 224 101374 226 101421
rect 300 101394 308 101463
rect 332 101461 342 101499
rect 400 101491 404 101500
rect 454 101485 504 101487
rect 494 101481 548 101485
rect 494 101476 514 101481
rect 504 101461 506 101476
rect 336 101449 342 101461
rect 289 101384 308 101394
rect 300 101378 308 101384
rect 332 101415 342 101449
rect 400 101453 404 101461
rect 400 101419 408 101453
rect 434 101419 438 101453
rect 498 101451 506 101461
rect 514 101451 515 101471
rect 504 101435 506 101451
rect 525 101442 528 101476
rect 547 101451 548 101471
rect 557 101451 564 101461
rect 514 101435 530 101441
rect 532 101435 548 101441
rect 332 101387 373 101415
rect 332 101381 351 101387
rect 107 101327 119 101361
rect 129 101327 149 101361
rect 196 101340 204 101374
rect 216 101340 232 101374
rect 244 101368 257 101374
rect 278 101368 291 101378
rect 244 101344 291 101368
rect 300 101368 321 101378
rect 336 101371 351 101381
rect 300 101344 329 101368
rect 332 101353 351 101371
rect 361 101381 375 101387
rect 400 101381 411 101419
rect 562 101382 612 101384
rect 361 101353 381 101381
rect 400 101353 409 101381
rect 466 101373 497 101381
rect 565 101373 596 101381
rect 442 101366 500 101373
rect 466 101365 500 101366
rect 565 101365 599 101373
rect 244 101340 257 101344
rect 42 101261 46 101295
rect 72 101261 76 101295
rect 42 101214 76 101218
rect 42 101199 46 101214
rect 72 101199 76 101214
rect 38 101181 80 101199
rect 16 101175 102 101181
rect 144 101175 148 101327
rect 174 101303 181 101331
rect 224 101293 226 101340
rect 300 101331 308 101344
rect 278 101320 305 101331
rect 332 101303 342 101353
rect 400 101333 404 101353
rect 497 101349 500 101365
rect 596 101349 599 101365
rect 466 101348 500 101349
rect 442 101341 500 101348
rect 565 101341 599 101349
rect 612 101332 614 101382
rect 256 101293 328 101301
rect 336 101295 342 101303
rect 400 101295 404 101303
rect 196 101263 204 101293
rect 216 101263 232 101293
rect 196 101259 232 101263
rect 196 101251 226 101259
rect 224 101235 226 101251
rect 332 101223 336 101291
rect 400 101261 408 101295
rect 434 101261 438 101295
rect 454 101279 504 101281
rect 504 101263 506 101279
rect 514 101273 530 101279
rect 532 101273 548 101279
rect 525 101263 548 101272
rect 400 101253 404 101261
rect 498 101253 506 101263
rect 504 101229 506 101253
rect 514 101243 515 101263
rect 525 101238 528 101263
rect 547 101243 548 101263
rect 557 101253 564 101263
rect 514 101229 548 101233
rect 400 101223 442 101224
rect 174 101213 246 101221
rect 400 101216 404 101223
rect 295 101182 300 101216
rect 324 101182 329 101216
rect 367 101199 438 101216
rect 367 101182 442 101199
rect 400 101181 442 101182
rect 378 101175 464 101181
rect 38 101159 80 101175
rect 400 101159 442 101175
rect -25 101145 25 101147
rect 42 101145 76 101159
rect 404 101145 438 101159
rect 455 101145 505 101147
rect 557 101145 607 101147
rect 16 101137 102 101145
rect 378 101137 464 101145
rect 8 101103 17 101137
rect 18 101135 51 101137
rect 80 101135 100 101137
rect 18 101103 100 101135
rect 380 101135 404 101137
rect 429 101135 438 101137
rect 442 101135 462 101137
rect 16 101095 102 101103
rect 42 101079 76 101095
rect 16 101059 38 101065
rect 42 101056 76 101060
rect 80 101059 102 101065
rect 42 101026 46 101056
rect 72 101026 76 101056
rect 42 100945 46 100979
rect 72 100945 76 100979
rect -25 100908 25 100910
rect -8 100900 14 100907
rect -8 100899 17 100900
rect 25 100899 27 100908
rect -12 100892 38 100899
rect -12 100891 34 100892
rect -12 100887 8 100891
rect 0 100875 8 100887
rect 14 100875 34 100891
rect 0 100874 34 100875
rect 0 100867 38 100874
rect 14 100866 17 100867
rect 25 100858 27 100867
rect 42 100838 45 100928
rect 69 100913 80 100945
rect 107 100913 143 100941
rect 144 100913 148 101133
rect 332 101065 336 101133
rect 380 101103 462 101135
rect 463 101103 472 101137
rect 480 101103 497 101137
rect 378 101095 464 101103
rect 505 101095 507 101145
rect 514 101103 548 101137
rect 565 101103 582 101137
rect 607 101095 609 101145
rect 404 101079 438 101095
rect 400 101065 442 101066
rect 378 101059 404 101065
rect 442 101059 464 101065
rect 400 101058 404 101059
rect 174 101019 246 101027
rect 295 101024 300 101058
rect 324 101024 329 101058
rect 224 100989 226 101005
rect 196 100981 226 100989
rect 332 100987 336 101055
rect 367 101024 438 101058
rect 400 101017 404 101024
rect 454 101011 504 101013
rect 494 101007 548 101011
rect 494 101002 514 101007
rect 504 100987 506 101002
rect 196 100977 232 100981
rect 196 100947 204 100977
rect 216 100947 232 100977
rect 400 100979 404 100987
rect 107 100907 119 100913
rect 109 100879 119 100907
rect 129 100879 149 100913
rect 174 100909 181 100939
rect 224 100900 226 100947
rect 256 100939 328 100947
rect 332 100945 336 100975
rect 400 100945 408 100979
rect 434 100945 438 100979
rect 498 100977 506 100987
rect 514 100977 515 100997
rect 504 100961 506 100977
rect 525 100968 528 101002
rect 547 100977 548 100997
rect 557 100977 564 100987
rect 514 100961 530 100967
rect 532 100961 548 100967
rect 278 100909 305 100920
rect 42 100787 46 100821
rect 72 100787 76 100821
rect 38 100749 80 100750
rect 42 100708 76 100742
rect 79 100708 113 100742
rect 42 100629 46 100663
rect 72 100629 76 100663
rect -25 100592 25 100594
rect -8 100584 14 100591
rect -8 100583 17 100584
rect 25 100583 27 100592
rect -12 100576 38 100583
rect -12 100575 34 100576
rect -12 100571 8 100575
rect 0 100559 8 100571
rect 14 100559 34 100575
rect 0 100558 34 100559
rect 0 100551 38 100558
rect 14 100550 17 100551
rect 25 100542 27 100551
rect 42 100522 45 100612
rect 71 100581 80 100609
rect 69 100543 80 100581
rect 144 100571 148 100879
rect 196 100866 204 100900
rect 216 100866 232 100900
rect 244 100896 257 100900
rect 300 100896 308 100909
rect 332 100907 342 100945
rect 400 100937 404 100945
rect 336 100897 342 100907
rect 244 100872 291 100896
rect 244 100866 257 100872
rect 224 100819 226 100866
rect 278 100862 291 100872
rect 300 100872 329 100896
rect 332 100887 342 100897
rect 400 100897 409 100925
rect 562 100908 612 100910
rect 466 100899 497 100907
rect 565 100899 596 100907
rect 300 100862 321 100872
rect 300 100856 308 100862
rect 289 100846 308 100856
rect 196 100789 204 100819
rect 216 100789 232 100819
rect 196 100785 232 100789
rect 196 100777 226 100785
rect 300 100777 308 100846
rect 332 100853 351 100887
rect 361 100859 381 100887
rect 361 100853 375 100859
rect 400 100853 411 100897
rect 442 100892 500 100899
rect 466 100891 500 100892
rect 565 100891 599 100899
rect 497 100875 500 100891
rect 596 100875 599 100891
rect 466 100874 500 100875
rect 442 100867 500 100874
rect 565 100867 599 100875
rect 612 100858 614 100908
rect 332 100829 342 100853
rect 336 100800 342 100829
rect 224 100761 226 100777
rect 332 100749 342 100800
rect 400 100821 404 100829
rect 400 100787 408 100821
rect 434 100787 438 100821
rect 454 100805 504 100807
rect 504 100789 506 100805
rect 514 100799 530 100805
rect 532 100799 548 100805
rect 525 100789 548 100798
rect 400 100779 404 100787
rect 498 100779 506 100789
rect 504 100755 506 100779
rect 514 100769 515 100789
rect 525 100764 528 100789
rect 547 100769 548 100789
rect 557 100779 564 100789
rect 514 100755 548 100759
rect 151 100708 156 100742
rect 174 100739 246 100747
rect 256 100739 328 100747
rect 336 100741 342 100749
rect 400 100744 404 100749
rect 180 100711 185 100739
rect 174 100703 246 100711
rect 256 100703 328 100711
rect 332 100709 336 100739
rect 400 100710 438 100744
rect 224 100673 226 100689
rect 196 100665 226 100673
rect 196 100661 232 100665
rect 196 100631 204 100661
rect 216 100631 232 100661
rect 224 100584 226 100631
rect 300 100604 308 100673
rect 332 100671 342 100709
rect 400 100701 404 100710
rect 454 100695 504 100697
rect 494 100691 548 100695
rect 494 100686 514 100691
rect 504 100671 506 100686
rect 336 100659 342 100671
rect 289 100594 308 100604
rect 300 100588 308 100594
rect 332 100625 342 100659
rect 400 100663 404 100671
rect 400 100629 408 100663
rect 434 100629 438 100663
rect 498 100661 506 100671
rect 514 100661 515 100681
rect 504 100645 506 100661
rect 525 100652 528 100686
rect 547 100661 548 100681
rect 557 100661 564 100671
rect 514 100645 530 100651
rect 532 100645 548 100651
rect 332 100597 373 100625
rect 332 100591 351 100597
rect 107 100537 119 100571
rect 129 100537 149 100571
rect 196 100550 204 100584
rect 216 100550 232 100584
rect 244 100578 257 100584
rect 278 100578 291 100588
rect 244 100554 291 100578
rect 300 100578 321 100588
rect 336 100581 351 100591
rect 300 100554 329 100578
rect 332 100563 351 100581
rect 361 100591 375 100597
rect 400 100591 411 100629
rect 562 100592 612 100594
rect 361 100563 381 100591
rect 400 100563 409 100591
rect 466 100583 497 100591
rect 565 100583 596 100591
rect 442 100576 500 100583
rect 466 100575 500 100576
rect 565 100575 599 100583
rect 244 100550 257 100554
rect 42 100471 46 100505
rect 72 100471 76 100505
rect 42 100424 76 100428
rect 42 100409 46 100424
rect 72 100409 76 100424
rect 38 100391 80 100409
rect 16 100385 102 100391
rect 144 100385 148 100537
rect 174 100513 181 100541
rect 224 100503 226 100550
rect 300 100541 308 100554
rect 278 100530 305 100541
rect 332 100513 342 100563
rect 400 100543 404 100563
rect 497 100559 500 100575
rect 596 100559 599 100575
rect 466 100558 500 100559
rect 442 100551 500 100558
rect 565 100551 599 100559
rect 612 100542 614 100592
rect 256 100503 328 100511
rect 336 100505 342 100513
rect 400 100505 404 100513
rect 196 100473 204 100503
rect 216 100473 232 100503
rect 196 100469 232 100473
rect 196 100461 226 100469
rect 224 100445 226 100461
rect 332 100433 336 100501
rect 400 100471 408 100505
rect 434 100471 438 100505
rect 454 100489 504 100491
rect 504 100473 506 100489
rect 514 100483 530 100489
rect 532 100483 548 100489
rect 525 100473 548 100482
rect 400 100463 404 100471
rect 498 100463 506 100473
rect 504 100439 506 100463
rect 514 100453 515 100473
rect 525 100448 528 100473
rect 547 100453 548 100473
rect 557 100463 564 100473
rect 514 100439 548 100443
rect 400 100433 442 100434
rect 174 100423 246 100431
rect 400 100426 404 100433
rect 295 100392 300 100426
rect 324 100392 329 100426
rect 367 100409 438 100426
rect 367 100392 442 100409
rect 400 100391 442 100392
rect 378 100385 464 100391
rect 38 100369 80 100385
rect 400 100369 442 100385
rect -25 100355 25 100357
rect 42 100355 76 100369
rect 404 100355 438 100369
rect 455 100355 505 100357
rect 557 100355 607 100357
rect 16 100347 102 100355
rect 378 100347 464 100355
rect 8 100313 17 100347
rect 18 100345 51 100347
rect 80 100345 100 100347
rect 18 100313 100 100345
rect 380 100345 404 100347
rect 429 100345 438 100347
rect 442 100345 462 100347
rect 16 100305 102 100313
rect 42 100289 76 100305
rect 16 100269 38 100275
rect 42 100266 76 100270
rect 80 100269 102 100275
rect 42 100236 46 100266
rect 72 100236 76 100266
rect 42 100155 46 100189
rect 72 100155 76 100189
rect -25 100118 25 100120
rect -8 100110 14 100117
rect -8 100109 17 100110
rect 25 100109 27 100118
rect -12 100102 38 100109
rect -12 100101 34 100102
rect -12 100097 8 100101
rect 0 100085 8 100097
rect 14 100085 34 100101
rect 0 100084 34 100085
rect 0 100077 38 100084
rect 14 100076 17 100077
rect 25 100068 27 100077
rect 42 100048 45 100138
rect 69 100123 80 100155
rect 107 100123 143 100151
rect 144 100123 148 100343
rect 332 100275 336 100343
rect 380 100313 462 100345
rect 463 100313 472 100347
rect 480 100313 497 100347
rect 378 100305 464 100313
rect 505 100305 507 100355
rect 514 100313 548 100347
rect 565 100313 582 100347
rect 607 100305 609 100355
rect 404 100289 438 100305
rect 400 100275 442 100276
rect 378 100269 404 100275
rect 442 100269 464 100275
rect 400 100268 404 100269
rect 174 100229 246 100237
rect 295 100234 300 100268
rect 324 100234 329 100268
rect 224 100199 226 100215
rect 196 100191 226 100199
rect 332 100197 336 100265
rect 367 100234 438 100268
rect 400 100227 404 100234
rect 454 100221 504 100223
rect 494 100217 548 100221
rect 494 100212 514 100217
rect 504 100197 506 100212
rect 196 100187 232 100191
rect 196 100157 204 100187
rect 216 100157 232 100187
rect 400 100189 404 100197
rect 107 100117 119 100123
rect 109 100089 119 100117
rect 129 100089 149 100123
rect 174 100119 181 100149
rect 224 100110 226 100157
rect 256 100149 328 100157
rect 332 100155 336 100185
rect 400 100155 408 100189
rect 434 100155 438 100189
rect 498 100187 506 100197
rect 514 100187 515 100207
rect 504 100171 506 100187
rect 525 100178 528 100212
rect 547 100187 548 100207
rect 557 100187 564 100197
rect 514 100171 530 100177
rect 532 100171 548 100177
rect 278 100119 305 100130
rect 42 99997 46 100031
rect 72 99997 76 100031
rect 38 99959 80 99960
rect 42 99918 76 99952
rect 79 99918 113 99952
rect 42 99839 46 99873
rect 72 99839 76 99873
rect -25 99802 25 99804
rect -8 99794 14 99801
rect -8 99793 17 99794
rect 25 99793 27 99802
rect -12 99786 38 99793
rect -12 99785 34 99786
rect -12 99781 8 99785
rect 0 99769 8 99781
rect 14 99769 34 99785
rect 0 99768 34 99769
rect 0 99761 38 99768
rect 14 99760 17 99761
rect 25 99752 27 99761
rect 42 99732 45 99822
rect 71 99791 80 99819
rect 69 99753 80 99791
rect 144 99781 148 100089
rect 196 100076 204 100110
rect 216 100076 232 100110
rect 244 100106 257 100110
rect 300 100106 308 100119
rect 332 100117 342 100155
rect 400 100147 404 100155
rect 336 100107 342 100117
rect 244 100082 291 100106
rect 244 100076 257 100082
rect 224 100029 226 100076
rect 278 100072 291 100082
rect 300 100082 329 100106
rect 332 100097 342 100107
rect 400 100107 409 100135
rect 562 100118 612 100120
rect 466 100109 497 100117
rect 565 100109 596 100117
rect 300 100072 321 100082
rect 300 100066 308 100072
rect 289 100056 308 100066
rect 196 99999 204 100029
rect 216 99999 232 100029
rect 196 99995 232 99999
rect 196 99987 226 99995
rect 300 99987 308 100056
rect 332 100063 351 100097
rect 361 100069 381 100097
rect 361 100063 375 100069
rect 400 100063 411 100107
rect 442 100102 500 100109
rect 466 100101 500 100102
rect 565 100101 599 100109
rect 497 100085 500 100101
rect 596 100085 599 100101
rect 466 100084 500 100085
rect 442 100077 500 100084
rect 565 100077 599 100085
rect 612 100068 614 100118
rect 332 100039 342 100063
rect 336 100027 342 100039
rect 224 99971 226 99987
rect 332 99959 342 100027
rect 400 100031 404 100039
rect 400 99997 408 100031
rect 434 99997 438 100031
rect 454 100015 504 100017
rect 504 99999 506 100015
rect 514 100009 530 100015
rect 532 100009 548 100015
rect 525 99999 548 100008
rect 400 99989 404 99997
rect 498 99989 506 99999
rect 504 99965 506 99989
rect 514 99979 515 99999
rect 525 99974 528 99999
rect 547 99979 548 99999
rect 557 99989 564 99999
rect 514 99965 548 99969
rect 151 99918 156 99952
rect 174 99949 246 99957
rect 256 99949 328 99957
rect 336 99951 342 99959
rect 400 99954 404 99959
rect 180 99921 185 99949
rect 174 99913 246 99921
rect 256 99913 328 99921
rect 332 99919 336 99949
rect 400 99920 438 99954
rect 224 99883 226 99899
rect 196 99875 226 99883
rect 196 99871 232 99875
rect 196 99841 204 99871
rect 216 99841 232 99871
rect 224 99794 226 99841
rect 300 99814 308 99883
rect 332 99881 342 99919
rect 400 99911 404 99920
rect 454 99905 504 99907
rect 494 99901 548 99905
rect 494 99896 514 99901
rect 504 99881 506 99896
rect 336 99869 342 99881
rect 289 99804 308 99814
rect 300 99798 308 99804
rect 332 99835 342 99869
rect 400 99873 404 99881
rect 400 99839 408 99873
rect 434 99839 438 99873
rect 498 99871 506 99881
rect 514 99871 515 99891
rect 504 99855 506 99871
rect 525 99862 528 99896
rect 547 99871 548 99891
rect 557 99871 564 99881
rect 514 99855 530 99861
rect 532 99855 548 99861
rect 332 99807 373 99835
rect 332 99801 351 99807
rect 107 99747 119 99781
rect 129 99747 149 99781
rect 196 99760 204 99794
rect 216 99760 232 99794
rect 244 99788 257 99794
rect 278 99788 291 99798
rect 244 99764 291 99788
rect 300 99788 321 99798
rect 336 99791 351 99801
rect 300 99764 329 99788
rect 332 99773 351 99791
rect 361 99801 375 99807
rect 400 99801 411 99839
rect 562 99802 612 99804
rect 361 99773 381 99801
rect 400 99773 409 99801
rect 466 99793 497 99801
rect 565 99793 596 99801
rect 442 99786 500 99793
rect 466 99785 500 99786
rect 565 99785 599 99793
rect 244 99760 257 99764
rect 42 99681 46 99715
rect 72 99681 76 99715
rect 42 99634 76 99638
rect 42 99619 46 99634
rect 72 99619 76 99634
rect 38 99601 80 99619
rect 16 99595 102 99601
rect 144 99595 148 99747
rect 174 99723 181 99751
rect 224 99713 226 99760
rect 300 99751 308 99764
rect 278 99740 305 99751
rect 332 99723 342 99773
rect 400 99753 404 99773
rect 497 99769 500 99785
rect 596 99769 599 99785
rect 466 99768 500 99769
rect 442 99761 500 99768
rect 565 99761 599 99769
rect 612 99752 614 99802
rect 256 99713 328 99721
rect 336 99715 342 99723
rect 400 99715 404 99723
rect 196 99683 204 99713
rect 216 99683 232 99713
rect 196 99679 232 99683
rect 196 99671 226 99679
rect 224 99655 226 99671
rect 332 99643 336 99711
rect 400 99681 408 99715
rect 434 99681 438 99715
rect 454 99699 504 99701
rect 504 99683 506 99699
rect 514 99693 530 99699
rect 532 99693 548 99699
rect 525 99683 548 99692
rect 400 99673 404 99681
rect 498 99673 506 99683
rect 504 99649 506 99673
rect 514 99663 515 99683
rect 525 99658 528 99683
rect 547 99663 548 99683
rect 557 99673 564 99683
rect 514 99649 548 99653
rect 400 99643 442 99644
rect 174 99633 246 99641
rect 400 99636 404 99643
rect 295 99602 300 99636
rect 324 99602 329 99636
rect 367 99619 438 99636
rect 367 99602 442 99619
rect 400 99601 442 99602
rect 378 99595 464 99601
rect 38 99579 80 99595
rect 400 99579 442 99595
rect -25 99565 25 99567
rect 42 99565 76 99579
rect 404 99565 438 99579
rect 455 99565 505 99567
rect 557 99565 607 99567
rect 16 99557 102 99565
rect 378 99557 464 99565
rect 8 99523 17 99557
rect 18 99555 51 99557
rect 80 99555 100 99557
rect 18 99523 100 99555
rect 380 99555 404 99557
rect 429 99555 438 99557
rect 442 99555 462 99557
rect 16 99515 102 99523
rect 42 99499 76 99515
rect 16 99479 38 99485
rect 42 99476 76 99480
rect 80 99479 102 99485
rect 42 99446 46 99476
rect 72 99446 76 99476
rect 42 99365 46 99399
rect 72 99365 76 99399
rect -25 99328 25 99330
rect -8 99320 14 99327
rect -8 99319 17 99320
rect 25 99319 27 99328
rect -12 99312 38 99319
rect -12 99311 34 99312
rect -12 99307 8 99311
rect 0 99295 8 99307
rect 14 99295 34 99311
rect 0 99294 34 99295
rect 0 99287 38 99294
rect 14 99286 17 99287
rect 25 99278 27 99287
rect 42 99258 45 99348
rect 69 99333 80 99365
rect 107 99333 143 99361
rect 144 99333 148 99553
rect 332 99485 336 99553
rect 380 99523 462 99555
rect 463 99523 472 99557
rect 480 99523 497 99557
rect 378 99515 464 99523
rect 505 99515 507 99565
rect 514 99523 548 99557
rect 565 99523 582 99557
rect 607 99515 609 99565
rect 404 99499 438 99515
rect 400 99485 442 99486
rect 378 99479 404 99485
rect 442 99479 464 99485
rect 400 99478 404 99479
rect 174 99439 246 99447
rect 295 99444 300 99478
rect 324 99444 329 99478
rect 224 99409 226 99425
rect 196 99401 226 99409
rect 332 99407 336 99475
rect 367 99444 438 99478
rect 400 99437 404 99444
rect 454 99431 504 99433
rect 494 99427 548 99431
rect 494 99422 514 99427
rect 504 99407 506 99422
rect 196 99397 232 99401
rect 196 99367 204 99397
rect 216 99367 232 99397
rect 400 99399 404 99407
rect 107 99327 119 99333
rect 109 99299 119 99327
rect 129 99299 149 99333
rect 174 99329 181 99359
rect 224 99320 226 99367
rect 256 99359 328 99367
rect 332 99365 336 99395
rect 400 99365 408 99399
rect 434 99365 438 99399
rect 498 99397 506 99407
rect 514 99397 515 99417
rect 504 99381 506 99397
rect 525 99388 528 99422
rect 547 99397 548 99417
rect 557 99397 564 99407
rect 514 99381 530 99387
rect 532 99381 548 99387
rect 278 99329 305 99340
rect 42 99207 46 99241
rect 72 99207 76 99241
rect 38 99169 80 99170
rect 42 99128 76 99162
rect 79 99128 113 99162
rect 42 99049 46 99083
rect 72 99049 76 99083
rect -25 99012 25 99014
rect -8 99004 14 99011
rect -8 99003 17 99004
rect 25 99003 27 99012
rect -12 98996 38 99003
rect -12 98995 34 98996
rect -12 98991 8 98995
rect 0 98979 8 98991
rect 14 98979 34 98995
rect 0 98978 34 98979
rect 0 98971 38 98978
rect 14 98970 17 98971
rect 25 98962 27 98971
rect 42 98942 45 99032
rect 71 99001 80 99029
rect 69 98963 80 99001
rect 144 98991 148 99299
rect 196 99286 204 99320
rect 216 99286 232 99320
rect 244 99316 257 99320
rect 300 99316 308 99329
rect 332 99327 342 99365
rect 400 99357 404 99365
rect 336 99317 342 99327
rect 244 99292 291 99316
rect 244 99286 257 99292
rect 224 99239 226 99286
rect 278 99282 291 99292
rect 300 99292 329 99316
rect 332 99307 342 99317
rect 400 99317 409 99345
rect 562 99328 612 99330
rect 466 99319 497 99327
rect 565 99319 596 99327
rect 300 99282 321 99292
rect 300 99276 308 99282
rect 289 99266 308 99276
rect 196 99209 204 99239
rect 216 99209 232 99239
rect 196 99205 232 99209
rect 196 99197 226 99205
rect 300 99197 308 99266
rect 332 99273 351 99307
rect 361 99279 381 99307
rect 361 99273 375 99279
rect 400 99273 411 99317
rect 442 99312 500 99319
rect 466 99311 500 99312
rect 565 99311 599 99319
rect 497 99295 500 99311
rect 596 99295 599 99311
rect 466 99294 500 99295
rect 442 99287 500 99294
rect 565 99287 599 99295
rect 612 99278 614 99328
rect 332 99249 342 99273
rect 336 99237 342 99249
rect 224 99181 226 99197
rect 332 99169 342 99237
rect 400 99241 404 99249
rect 400 99207 408 99241
rect 434 99207 438 99241
rect 454 99225 504 99227
rect 504 99209 506 99225
rect 514 99219 530 99225
rect 532 99219 548 99225
rect 525 99209 548 99218
rect 400 99199 404 99207
rect 498 99199 506 99209
rect 504 99175 506 99199
rect 514 99189 515 99209
rect 525 99184 528 99209
rect 547 99189 548 99209
rect 557 99199 564 99209
rect 514 99175 548 99179
rect 151 99128 156 99162
rect 174 99159 246 99167
rect 256 99159 328 99167
rect 336 99161 342 99169
rect 400 99164 404 99169
rect 180 99131 185 99159
rect 174 99123 246 99131
rect 256 99123 328 99131
rect 332 99129 336 99159
rect 400 99130 438 99164
rect 224 99093 226 99109
rect 196 99085 226 99093
rect 196 99081 232 99085
rect 196 99051 204 99081
rect 216 99051 232 99081
rect 224 99004 226 99051
rect 300 99024 308 99093
rect 332 99091 342 99129
rect 400 99121 404 99130
rect 454 99115 504 99117
rect 494 99111 548 99115
rect 494 99106 514 99111
rect 504 99091 506 99106
rect 336 99079 342 99091
rect 289 99014 308 99024
rect 300 99008 308 99014
rect 332 99045 342 99079
rect 400 99083 404 99091
rect 400 99049 408 99083
rect 434 99049 438 99083
rect 498 99081 506 99091
rect 514 99081 515 99101
rect 504 99065 506 99081
rect 525 99072 528 99106
rect 547 99081 548 99101
rect 557 99081 564 99091
rect 514 99065 530 99071
rect 532 99065 548 99071
rect 332 99017 373 99045
rect 332 99011 351 99017
rect 107 98957 119 98991
rect 129 98957 149 98991
rect 196 98970 204 99004
rect 216 98970 232 99004
rect 244 98998 257 99004
rect 278 98998 291 99008
rect 244 98974 291 98998
rect 300 98998 321 99008
rect 336 99001 351 99011
rect 300 98974 329 98998
rect 332 98983 351 99001
rect 361 99011 375 99017
rect 400 99011 411 99049
rect 562 99012 612 99014
rect 361 98983 381 99011
rect 400 98983 409 99011
rect 466 99003 497 99011
rect 565 99003 596 99011
rect 442 98996 500 99003
rect 466 98995 500 98996
rect 565 98995 599 99003
rect 244 98970 257 98974
rect 42 98891 46 98925
rect 72 98891 76 98925
rect 42 98844 76 98848
rect 42 98829 46 98844
rect 72 98829 76 98844
rect 38 98811 80 98829
rect 16 98805 102 98811
rect 144 98805 148 98957
rect 174 98933 181 98961
rect 224 98923 226 98970
rect 300 98961 308 98974
rect 278 98950 305 98961
rect 332 98933 342 98983
rect 400 98963 404 98983
rect 497 98979 500 98995
rect 596 98979 599 98995
rect 466 98978 500 98979
rect 442 98971 500 98978
rect 565 98971 599 98979
rect 612 98962 614 99012
rect 256 98923 328 98931
rect 336 98925 342 98933
rect 400 98925 404 98933
rect 196 98893 204 98923
rect 216 98893 232 98923
rect 196 98889 232 98893
rect 196 98881 226 98889
rect 224 98865 226 98881
rect 332 98853 336 98921
rect 400 98891 408 98925
rect 434 98891 438 98925
rect 454 98909 504 98911
rect 504 98893 506 98909
rect 514 98903 530 98909
rect 532 98903 548 98909
rect 525 98893 548 98902
rect 400 98883 404 98891
rect 498 98883 506 98893
rect 504 98859 506 98883
rect 514 98873 515 98893
rect 525 98868 528 98893
rect 547 98873 548 98893
rect 557 98883 564 98893
rect 514 98859 548 98863
rect 400 98853 442 98854
rect 174 98843 246 98851
rect 400 98846 404 98853
rect 295 98812 300 98846
rect 324 98812 329 98846
rect 367 98829 438 98846
rect 367 98812 442 98829
rect 400 98811 442 98812
rect 378 98805 464 98811
rect 38 98789 80 98805
rect 400 98789 442 98805
rect -25 98775 25 98777
rect 42 98775 76 98789
rect 404 98775 438 98789
rect 455 98775 505 98777
rect 557 98775 607 98777
rect 16 98767 102 98775
rect 378 98767 464 98775
rect 8 98733 17 98767
rect 18 98765 51 98767
rect 80 98765 100 98767
rect 18 98733 100 98765
rect 380 98765 404 98767
rect 429 98765 438 98767
rect 442 98765 462 98767
rect 16 98725 102 98733
rect 42 98709 76 98725
rect 16 98689 38 98695
rect 42 98686 76 98690
rect 80 98689 102 98695
rect 42 98656 46 98686
rect 72 98656 76 98686
rect 42 98575 46 98609
rect 72 98575 76 98609
rect -25 98538 25 98540
rect -8 98530 14 98537
rect -8 98529 17 98530
rect 25 98529 27 98538
rect -12 98522 38 98529
rect -12 98521 34 98522
rect -12 98517 8 98521
rect 0 98505 8 98517
rect 14 98505 34 98521
rect 0 98504 34 98505
rect 0 98497 38 98504
rect 14 98496 17 98497
rect 25 98488 27 98497
rect 42 98468 45 98558
rect 69 98543 80 98575
rect 107 98543 143 98571
rect 144 98543 148 98763
rect 332 98695 336 98763
rect 380 98733 462 98765
rect 463 98733 472 98767
rect 480 98733 497 98767
rect 378 98725 464 98733
rect 505 98725 507 98775
rect 514 98733 548 98767
rect 565 98733 582 98767
rect 607 98725 609 98775
rect 404 98709 438 98725
rect 400 98695 442 98696
rect 378 98689 404 98695
rect 442 98689 464 98695
rect 400 98688 404 98689
rect 174 98649 246 98657
rect 295 98654 300 98688
rect 324 98654 329 98688
rect 224 98619 226 98635
rect 196 98611 226 98619
rect 332 98617 336 98685
rect 367 98654 438 98688
rect 400 98647 404 98654
rect 454 98641 504 98643
rect 494 98637 548 98641
rect 494 98632 514 98637
rect 504 98617 506 98632
rect 196 98607 232 98611
rect 196 98577 204 98607
rect 216 98577 232 98607
rect 400 98609 404 98617
rect 107 98537 119 98543
rect 109 98509 119 98537
rect 129 98509 149 98543
rect 174 98539 181 98569
rect 224 98530 226 98577
rect 256 98569 328 98577
rect 332 98575 336 98605
rect 400 98575 408 98609
rect 434 98575 438 98609
rect 498 98607 506 98617
rect 514 98607 515 98627
rect 504 98591 506 98607
rect 525 98598 528 98632
rect 547 98607 548 98627
rect 557 98607 564 98617
rect 514 98591 530 98597
rect 532 98591 548 98597
rect 278 98539 305 98550
rect 42 98417 46 98451
rect 72 98417 76 98451
rect 38 98379 80 98380
rect 42 98338 76 98372
rect 79 98338 113 98372
rect 42 98259 46 98293
rect 72 98259 76 98293
rect -25 98222 25 98224
rect -8 98214 14 98221
rect -8 98213 17 98214
rect 25 98213 27 98222
rect -12 98206 38 98213
rect -12 98205 34 98206
rect -12 98201 8 98205
rect 0 98189 8 98201
rect 14 98189 34 98205
rect 0 98188 34 98189
rect 0 98181 38 98188
rect 14 98180 17 98181
rect 25 98172 27 98181
rect 42 98152 45 98242
rect 71 98211 80 98239
rect 69 98173 80 98211
rect 144 98201 148 98509
rect 196 98496 204 98530
rect 216 98496 232 98530
rect 244 98526 257 98530
rect 300 98526 308 98539
rect 332 98537 342 98575
rect 400 98567 404 98575
rect 336 98527 342 98537
rect 244 98502 291 98526
rect 244 98496 257 98502
rect 224 98449 226 98496
rect 278 98492 291 98502
rect 300 98502 329 98526
rect 332 98517 342 98527
rect 400 98527 409 98555
rect 562 98538 612 98540
rect 466 98529 497 98537
rect 565 98529 596 98537
rect 300 98492 321 98502
rect 300 98486 308 98492
rect 289 98476 308 98486
rect 196 98419 204 98449
rect 216 98419 232 98449
rect 196 98415 232 98419
rect 196 98407 226 98415
rect 300 98407 308 98476
rect 332 98483 351 98517
rect 361 98489 381 98517
rect 361 98483 375 98489
rect 400 98483 411 98527
rect 442 98522 500 98529
rect 466 98521 500 98522
rect 565 98521 599 98529
rect 497 98505 500 98521
rect 596 98505 599 98521
rect 466 98504 500 98505
rect 442 98497 500 98504
rect 565 98497 599 98505
rect 612 98488 614 98538
rect 332 98459 342 98483
rect 336 98447 342 98459
rect 224 98391 226 98407
rect 332 98379 342 98447
rect 400 98451 404 98459
rect 400 98417 408 98451
rect 434 98417 438 98451
rect 454 98435 504 98437
rect 504 98419 506 98435
rect 514 98429 530 98435
rect 532 98429 548 98435
rect 525 98419 548 98428
rect 400 98409 404 98417
rect 498 98409 506 98419
rect 504 98385 506 98409
rect 514 98399 515 98419
rect 525 98394 528 98419
rect 547 98399 548 98419
rect 557 98409 564 98419
rect 514 98385 548 98389
rect 151 98338 156 98372
rect 174 98369 246 98377
rect 256 98369 328 98377
rect 336 98371 342 98379
rect 400 98374 404 98379
rect 180 98341 185 98369
rect 174 98333 246 98341
rect 256 98333 328 98341
rect 332 98339 336 98369
rect 400 98340 438 98374
rect 224 98303 226 98319
rect 196 98295 226 98303
rect 196 98291 232 98295
rect 196 98261 204 98291
rect 216 98261 232 98291
rect 224 98214 226 98261
rect 300 98234 308 98303
rect 332 98301 342 98339
rect 400 98331 404 98340
rect 454 98325 504 98327
rect 494 98321 548 98325
rect 494 98316 514 98321
rect 504 98301 506 98316
rect 336 98289 342 98301
rect 289 98224 308 98234
rect 300 98218 308 98224
rect 332 98255 342 98289
rect 400 98293 404 98301
rect 400 98259 408 98293
rect 434 98259 438 98293
rect 498 98291 506 98301
rect 514 98291 515 98311
rect 504 98275 506 98291
rect 525 98282 528 98316
rect 547 98291 548 98311
rect 557 98291 564 98301
rect 514 98275 530 98281
rect 532 98275 548 98281
rect 332 98227 373 98255
rect 332 98221 351 98227
rect 107 98167 119 98201
rect 129 98167 149 98201
rect 196 98180 204 98214
rect 216 98180 232 98214
rect 244 98208 257 98214
rect 278 98208 291 98218
rect 244 98184 291 98208
rect 300 98208 321 98218
rect 336 98211 351 98221
rect 300 98184 329 98208
rect 332 98193 351 98211
rect 361 98221 375 98227
rect 400 98221 411 98259
rect 562 98222 612 98224
rect 361 98193 381 98221
rect 400 98193 409 98221
rect 466 98213 497 98221
rect 565 98213 596 98221
rect 442 98206 500 98213
rect 466 98205 500 98206
rect 565 98205 599 98213
rect 244 98180 257 98184
rect 42 98101 46 98135
rect 72 98101 76 98135
rect 42 98054 76 98058
rect 42 98039 46 98054
rect 72 98039 76 98054
rect 38 98021 80 98039
rect 16 98015 102 98021
rect 144 98015 148 98167
rect 174 98143 181 98171
rect 224 98133 226 98180
rect 300 98171 308 98184
rect 278 98160 305 98171
rect 332 98143 342 98193
rect 400 98173 404 98193
rect 497 98189 500 98205
rect 596 98189 599 98205
rect 466 98188 500 98189
rect 442 98181 500 98188
rect 565 98181 599 98189
rect 612 98172 614 98222
rect 256 98133 328 98141
rect 336 98135 342 98143
rect 400 98135 404 98143
rect 196 98103 204 98133
rect 216 98103 232 98133
rect 196 98099 232 98103
rect 196 98091 226 98099
rect 224 98075 226 98091
rect 332 98063 336 98131
rect 400 98101 408 98135
rect 434 98101 438 98135
rect 454 98119 504 98121
rect 504 98103 506 98119
rect 514 98113 530 98119
rect 532 98113 548 98119
rect 525 98103 548 98112
rect 400 98093 404 98101
rect 498 98093 506 98103
rect 504 98069 506 98093
rect 514 98083 515 98103
rect 525 98078 528 98103
rect 547 98083 548 98103
rect 557 98093 564 98103
rect 514 98069 548 98073
rect 400 98063 442 98064
rect 174 98053 246 98061
rect 400 98056 404 98063
rect 295 98022 300 98056
rect 324 98022 329 98056
rect 367 98039 438 98056
rect 367 98022 442 98039
rect 400 98021 442 98022
rect 378 98015 464 98021
rect 38 97999 80 98015
rect 400 97999 442 98015
rect -25 97985 25 97987
rect 42 97985 76 97999
rect 404 97985 438 97999
rect 455 97985 505 97987
rect 557 97985 607 97987
rect 16 97977 102 97985
rect 378 97977 464 97985
rect 8 97943 17 97977
rect 18 97975 51 97977
rect 80 97975 100 97977
rect 18 97943 100 97975
rect 380 97975 404 97977
rect 429 97975 438 97977
rect 442 97975 462 97977
rect 16 97935 102 97943
rect 42 97919 76 97935
rect 16 97899 38 97905
rect 42 97896 76 97900
rect 80 97899 102 97905
rect 42 97866 46 97896
rect 72 97866 76 97896
rect 42 97785 46 97819
rect 72 97785 76 97819
rect -25 97748 25 97750
rect -8 97740 14 97747
rect -8 97739 17 97740
rect 25 97739 27 97748
rect -12 97732 38 97739
rect -12 97731 34 97732
rect -12 97727 8 97731
rect 0 97715 8 97727
rect 14 97715 34 97731
rect 0 97714 34 97715
rect 0 97707 38 97714
rect 14 97706 17 97707
rect 25 97698 27 97707
rect 42 97678 45 97768
rect 69 97753 80 97785
rect 107 97753 143 97781
rect 144 97753 148 97973
rect 332 97905 336 97973
rect 380 97943 462 97975
rect 463 97943 472 97977
rect 480 97943 497 97977
rect 378 97935 464 97943
rect 505 97935 507 97985
rect 514 97943 548 97977
rect 565 97943 582 97977
rect 607 97935 609 97985
rect 404 97919 438 97935
rect 400 97905 442 97906
rect 378 97899 404 97905
rect 442 97899 464 97905
rect 400 97898 404 97899
rect 174 97859 246 97867
rect 295 97864 300 97898
rect 324 97864 329 97898
rect 224 97829 226 97845
rect 196 97821 226 97829
rect 332 97827 336 97895
rect 367 97864 438 97898
rect 400 97857 404 97864
rect 454 97851 504 97853
rect 494 97847 548 97851
rect 494 97842 514 97847
rect 504 97827 506 97842
rect 196 97817 232 97821
rect 196 97787 204 97817
rect 216 97787 232 97817
rect 400 97819 404 97827
rect 107 97747 119 97753
rect 109 97719 119 97747
rect 129 97719 149 97753
rect 174 97749 181 97779
rect 224 97740 226 97787
rect 256 97779 328 97787
rect 332 97785 336 97815
rect 400 97785 408 97819
rect 434 97785 438 97819
rect 498 97817 506 97827
rect 514 97817 515 97837
rect 504 97801 506 97817
rect 525 97808 528 97842
rect 547 97817 548 97837
rect 557 97817 564 97827
rect 514 97801 530 97807
rect 532 97801 548 97807
rect 278 97749 305 97760
rect 42 97627 46 97661
rect 72 97627 76 97661
rect 38 97589 80 97590
rect 42 97548 76 97582
rect 79 97548 113 97582
rect 42 97469 46 97503
rect 72 97469 76 97503
rect -25 97432 25 97434
rect -8 97424 14 97431
rect -8 97423 17 97424
rect 25 97423 27 97432
rect -12 97416 38 97423
rect -12 97415 34 97416
rect -12 97411 8 97415
rect 0 97399 8 97411
rect 14 97399 34 97415
rect 0 97398 34 97399
rect 0 97391 38 97398
rect 14 97390 17 97391
rect 25 97382 27 97391
rect 42 97362 45 97452
rect 71 97421 80 97449
rect 69 97383 80 97421
rect 144 97411 148 97719
rect 196 97706 204 97740
rect 216 97706 232 97740
rect 244 97736 257 97740
rect 300 97736 308 97749
rect 332 97747 342 97785
rect 400 97777 404 97785
rect 336 97737 342 97747
rect 244 97712 291 97736
rect 244 97706 257 97712
rect 224 97659 226 97706
rect 278 97702 291 97712
rect 300 97712 329 97736
rect 332 97727 342 97737
rect 400 97737 409 97765
rect 562 97748 612 97750
rect 466 97739 497 97747
rect 565 97739 596 97747
rect 300 97702 321 97712
rect 300 97696 308 97702
rect 289 97686 308 97696
rect 196 97629 204 97659
rect 216 97629 232 97659
rect 196 97625 232 97629
rect 196 97617 226 97625
rect 300 97617 308 97686
rect 332 97693 351 97727
rect 361 97699 381 97727
rect 361 97693 375 97699
rect 400 97693 411 97737
rect 442 97732 500 97739
rect 466 97731 500 97732
rect 565 97731 599 97739
rect 497 97715 500 97731
rect 596 97715 599 97731
rect 466 97714 500 97715
rect 442 97707 500 97714
rect 565 97707 599 97715
rect 612 97698 614 97748
rect 332 97669 342 97693
rect 336 97657 342 97669
rect 224 97601 226 97617
rect 332 97589 342 97657
rect 400 97661 404 97669
rect 400 97627 408 97661
rect 434 97627 438 97661
rect 454 97645 504 97647
rect 504 97629 506 97645
rect 514 97639 530 97645
rect 532 97639 548 97645
rect 525 97629 548 97638
rect 400 97619 404 97627
rect 498 97619 506 97629
rect 504 97595 506 97619
rect 514 97609 515 97629
rect 525 97604 528 97629
rect 547 97609 548 97629
rect 557 97619 564 97629
rect 514 97595 548 97599
rect 151 97548 156 97582
rect 174 97579 246 97587
rect 256 97579 328 97587
rect 336 97581 342 97589
rect 400 97584 404 97589
rect 180 97551 185 97579
rect 174 97543 246 97551
rect 256 97543 328 97551
rect 332 97549 336 97579
rect 400 97550 438 97584
rect 224 97513 226 97529
rect 196 97505 226 97513
rect 196 97501 232 97505
rect 196 97471 204 97501
rect 216 97471 232 97501
rect 224 97424 226 97471
rect 300 97444 308 97513
rect 332 97511 342 97549
rect 400 97541 404 97550
rect 454 97535 504 97537
rect 494 97531 548 97535
rect 494 97526 514 97531
rect 504 97511 506 97526
rect 336 97499 342 97511
rect 289 97434 308 97444
rect 300 97428 308 97434
rect 332 97465 342 97499
rect 400 97503 404 97511
rect 400 97469 408 97503
rect 434 97469 438 97503
rect 498 97501 506 97511
rect 514 97501 515 97521
rect 504 97485 506 97501
rect 525 97492 528 97526
rect 547 97501 548 97521
rect 557 97501 564 97511
rect 514 97485 530 97491
rect 532 97485 548 97491
rect 332 97437 373 97465
rect 332 97431 351 97437
rect 107 97377 119 97411
rect 129 97377 149 97411
rect 196 97390 204 97424
rect 216 97390 232 97424
rect 244 97418 257 97424
rect 278 97418 291 97428
rect 244 97394 291 97418
rect 300 97418 321 97428
rect 336 97421 351 97431
rect 300 97394 329 97418
rect 332 97403 351 97421
rect 361 97431 375 97437
rect 400 97431 411 97469
rect 562 97432 612 97434
rect 361 97403 381 97431
rect 400 97403 409 97431
rect 466 97423 497 97431
rect 565 97423 596 97431
rect 442 97416 500 97423
rect 466 97415 500 97416
rect 565 97415 599 97423
rect 244 97390 257 97394
rect 42 97311 46 97345
rect 72 97311 76 97345
rect 42 97264 76 97268
rect 42 97249 46 97264
rect 72 97249 76 97264
rect 38 97231 80 97249
rect 16 97225 102 97231
rect 144 97225 148 97377
rect 174 97353 181 97381
rect 224 97343 226 97390
rect 300 97381 308 97394
rect 278 97370 305 97381
rect 332 97353 342 97403
rect 400 97383 404 97403
rect 497 97399 500 97415
rect 596 97399 599 97415
rect 466 97398 500 97399
rect 442 97391 500 97398
rect 565 97391 599 97399
rect 612 97382 614 97432
rect 256 97343 328 97351
rect 336 97345 342 97353
rect 400 97345 404 97353
rect 196 97313 204 97343
rect 216 97313 232 97343
rect 196 97309 232 97313
rect 196 97301 226 97309
rect 224 97285 226 97301
rect 332 97273 336 97341
rect 400 97311 408 97345
rect 434 97311 438 97345
rect 454 97329 504 97331
rect 504 97313 506 97329
rect 514 97323 530 97329
rect 532 97323 548 97329
rect 525 97313 548 97322
rect 400 97303 404 97311
rect 498 97303 506 97313
rect 504 97279 506 97303
rect 514 97293 515 97313
rect 525 97288 528 97313
rect 547 97293 548 97313
rect 557 97303 564 97313
rect 514 97279 548 97283
rect 400 97273 442 97274
rect 174 97263 246 97271
rect 400 97266 404 97273
rect 295 97232 300 97266
rect 324 97232 329 97266
rect 367 97249 438 97266
rect 367 97232 442 97249
rect 400 97231 442 97232
rect 378 97225 464 97231
rect 38 97209 80 97225
rect 400 97209 442 97225
rect -25 97195 25 97197
rect 42 97195 76 97209
rect 404 97195 438 97209
rect 455 97195 505 97197
rect 557 97195 607 97197
rect 16 97187 102 97195
rect 378 97187 464 97195
rect 8 97153 17 97187
rect 18 97185 51 97187
rect 80 97185 100 97187
rect 18 97153 100 97185
rect 380 97185 404 97187
rect 429 97185 438 97187
rect 442 97185 462 97187
rect 16 97145 102 97153
rect 42 97129 76 97145
rect 16 97109 38 97115
rect 42 97106 76 97110
rect 80 97109 102 97115
rect 42 97076 46 97106
rect 72 97076 76 97106
rect 42 96995 46 97029
rect 72 96995 76 97029
rect -25 96958 25 96960
rect -8 96950 14 96957
rect -8 96949 17 96950
rect 25 96949 27 96958
rect -12 96942 38 96949
rect -12 96941 34 96942
rect -12 96937 8 96941
rect 0 96925 8 96937
rect 14 96925 34 96941
rect 0 96924 34 96925
rect 0 96917 38 96924
rect 14 96916 17 96917
rect 25 96908 27 96917
rect 42 96888 45 96978
rect 69 96963 80 96995
rect 107 96963 143 96991
rect 144 96963 148 97183
rect 332 97115 336 97183
rect 380 97153 462 97185
rect 463 97153 472 97187
rect 480 97153 497 97187
rect 378 97145 464 97153
rect 505 97145 507 97195
rect 514 97153 548 97187
rect 565 97153 582 97187
rect 607 97145 609 97195
rect 404 97129 438 97145
rect 400 97115 442 97116
rect 378 97109 404 97115
rect 442 97109 464 97115
rect 400 97108 404 97109
rect 174 97069 246 97077
rect 295 97074 300 97108
rect 324 97074 329 97108
rect 224 97039 226 97055
rect 196 97031 226 97039
rect 332 97037 336 97105
rect 367 97074 438 97108
rect 400 97067 404 97074
rect 454 97061 504 97063
rect 494 97057 548 97061
rect 494 97052 514 97057
rect 504 97037 506 97052
rect 196 97027 232 97031
rect 196 96997 204 97027
rect 216 96997 232 97027
rect 400 97029 404 97037
rect 107 96957 119 96963
rect 109 96929 119 96957
rect 129 96929 149 96963
rect 174 96959 181 96989
rect 224 96950 226 96997
rect 256 96989 328 96997
rect 332 96995 336 97025
rect 400 96995 408 97029
rect 434 96995 438 97029
rect 498 97027 506 97037
rect 514 97027 515 97047
rect 504 97011 506 97027
rect 525 97018 528 97052
rect 547 97027 548 97047
rect 557 97027 564 97037
rect 514 97011 530 97017
rect 532 97011 548 97017
rect 278 96959 305 96970
rect 42 96837 46 96871
rect 72 96837 76 96871
rect 38 96799 80 96800
rect 42 96758 76 96792
rect 79 96758 113 96792
rect 42 96679 46 96713
rect 72 96679 76 96713
rect -25 96642 25 96644
rect -8 96634 14 96641
rect -8 96633 17 96634
rect 25 96633 27 96642
rect -12 96626 38 96633
rect -12 96625 34 96626
rect -12 96621 8 96625
rect 0 96609 8 96621
rect 14 96609 34 96625
rect 0 96608 34 96609
rect 0 96601 38 96608
rect 14 96600 17 96601
rect 25 96592 27 96601
rect 42 96572 45 96662
rect 71 96631 80 96659
rect 69 96593 80 96631
rect 144 96621 148 96929
rect 196 96916 204 96950
rect 216 96916 232 96950
rect 244 96946 257 96950
rect 300 96946 308 96959
rect 332 96957 342 96995
rect 400 96987 404 96995
rect 336 96947 342 96957
rect 244 96922 291 96946
rect 244 96916 257 96922
rect 224 96869 226 96916
rect 278 96912 291 96922
rect 300 96922 329 96946
rect 332 96937 342 96947
rect 400 96947 409 96975
rect 562 96958 612 96960
rect 466 96949 497 96957
rect 565 96949 596 96957
rect 300 96912 321 96922
rect 300 96906 308 96912
rect 289 96896 308 96906
rect 196 96839 204 96869
rect 216 96839 232 96869
rect 196 96835 232 96839
rect 196 96827 226 96835
rect 300 96827 308 96896
rect 332 96903 351 96937
rect 361 96909 381 96937
rect 361 96903 375 96909
rect 400 96903 411 96947
rect 442 96942 500 96949
rect 466 96941 500 96942
rect 565 96941 599 96949
rect 497 96925 500 96941
rect 596 96925 599 96941
rect 466 96924 500 96925
rect 442 96917 500 96924
rect 565 96917 599 96925
rect 612 96908 614 96958
rect 332 96879 342 96903
rect 336 96867 342 96879
rect 224 96811 226 96827
rect 332 96799 342 96867
rect 400 96871 404 96879
rect 400 96837 408 96871
rect 434 96837 438 96871
rect 454 96855 504 96857
rect 504 96839 506 96855
rect 514 96849 530 96855
rect 532 96849 548 96855
rect 525 96839 548 96848
rect 400 96829 404 96837
rect 498 96829 506 96839
rect 504 96805 506 96829
rect 514 96819 515 96839
rect 525 96814 528 96839
rect 547 96819 548 96839
rect 557 96829 564 96839
rect 514 96805 548 96809
rect 151 96758 156 96792
rect 174 96789 246 96797
rect 256 96789 328 96797
rect 336 96791 342 96799
rect 400 96794 404 96799
rect 180 96761 185 96789
rect 174 96753 246 96761
rect 256 96753 328 96761
rect 332 96759 336 96789
rect 400 96760 438 96794
rect 224 96723 226 96739
rect 196 96715 226 96723
rect 196 96711 232 96715
rect 196 96681 204 96711
rect 216 96681 232 96711
rect 224 96634 226 96681
rect 300 96654 308 96723
rect 332 96721 342 96759
rect 400 96751 404 96760
rect 454 96745 504 96747
rect 494 96741 548 96745
rect 494 96736 514 96741
rect 504 96721 506 96736
rect 336 96709 342 96721
rect 289 96644 308 96654
rect 300 96638 308 96644
rect 332 96675 342 96709
rect 400 96713 404 96721
rect 400 96679 408 96713
rect 434 96679 438 96713
rect 498 96711 506 96721
rect 514 96711 515 96731
rect 504 96695 506 96711
rect 525 96702 528 96736
rect 547 96711 548 96731
rect 557 96711 564 96721
rect 514 96695 530 96701
rect 532 96695 548 96701
rect 332 96647 373 96675
rect 332 96641 351 96647
rect 107 96587 119 96621
rect 129 96587 149 96621
rect 196 96600 204 96634
rect 216 96600 232 96634
rect 244 96628 257 96634
rect 278 96628 291 96638
rect 244 96604 291 96628
rect 300 96628 321 96638
rect 336 96631 351 96641
rect 300 96604 329 96628
rect 332 96613 351 96631
rect 361 96641 375 96647
rect 400 96641 411 96679
rect 562 96642 612 96644
rect 361 96613 381 96641
rect 400 96613 409 96641
rect 466 96633 497 96641
rect 565 96633 596 96641
rect 442 96626 500 96633
rect 466 96625 500 96626
rect 565 96625 599 96633
rect 244 96600 257 96604
rect 42 96521 46 96555
rect 72 96521 76 96555
rect 42 96474 76 96478
rect 42 96459 46 96474
rect 72 96459 76 96474
rect 38 96441 80 96459
rect 16 96435 102 96441
rect 144 96435 148 96587
rect 174 96563 181 96591
rect 224 96553 226 96600
rect 300 96591 308 96604
rect 278 96580 305 96591
rect 332 96563 342 96613
rect 400 96593 404 96613
rect 497 96609 500 96625
rect 596 96609 599 96625
rect 466 96608 500 96609
rect 442 96601 500 96608
rect 565 96601 599 96609
rect 612 96592 614 96642
rect 256 96553 328 96561
rect 336 96555 342 96563
rect 400 96555 404 96563
rect 196 96523 204 96553
rect 216 96523 232 96553
rect 196 96519 232 96523
rect 196 96511 226 96519
rect 224 96495 226 96511
rect 332 96483 336 96551
rect 400 96521 408 96555
rect 434 96521 438 96555
rect 454 96539 504 96541
rect 504 96523 506 96539
rect 514 96533 530 96539
rect 532 96533 548 96539
rect 525 96523 548 96532
rect 400 96513 404 96521
rect 498 96513 506 96523
rect 504 96489 506 96513
rect 514 96503 515 96523
rect 525 96498 528 96523
rect 547 96503 548 96523
rect 557 96513 564 96523
rect 514 96489 548 96493
rect 400 96483 442 96484
rect 174 96473 246 96481
rect 400 96476 404 96483
rect 295 96442 300 96476
rect 324 96442 329 96476
rect 367 96459 438 96476
rect 367 96442 442 96459
rect 400 96441 442 96442
rect 378 96435 464 96441
rect 38 96419 80 96435
rect 400 96419 442 96435
rect -25 96405 25 96407
rect 42 96405 76 96419
rect 404 96405 438 96419
rect 455 96405 505 96407
rect 557 96405 607 96407
rect 16 96397 102 96405
rect 378 96397 464 96405
rect 8 96363 17 96397
rect 18 96395 51 96397
rect 80 96395 100 96397
rect 18 96363 100 96395
rect 380 96395 404 96397
rect 429 96395 438 96397
rect 442 96395 462 96397
rect 16 96355 102 96363
rect 42 96339 76 96355
rect 16 96319 38 96325
rect 42 96316 76 96320
rect 80 96319 102 96325
rect 42 96286 46 96316
rect 72 96286 76 96316
rect 42 96205 46 96239
rect 72 96205 76 96239
rect -25 96168 25 96170
rect -8 96160 14 96167
rect -8 96159 17 96160
rect 25 96159 27 96168
rect -12 96152 38 96159
rect -12 96151 34 96152
rect -12 96147 8 96151
rect 0 96135 8 96147
rect 14 96135 34 96151
rect 0 96134 34 96135
rect 0 96127 38 96134
rect 14 96126 17 96127
rect 25 96118 27 96127
rect 42 96098 45 96188
rect 69 96173 80 96205
rect 107 96173 143 96201
rect 144 96173 148 96393
rect 332 96325 336 96393
rect 380 96363 462 96395
rect 463 96363 472 96397
rect 480 96363 497 96397
rect 378 96355 464 96363
rect 505 96355 507 96405
rect 514 96363 548 96397
rect 565 96363 582 96397
rect 607 96355 609 96405
rect 404 96339 438 96355
rect 400 96325 442 96326
rect 378 96319 404 96325
rect 442 96319 464 96325
rect 400 96318 404 96319
rect 174 96279 246 96287
rect 295 96284 300 96318
rect 324 96284 329 96318
rect 224 96249 226 96265
rect 196 96241 226 96249
rect 332 96247 336 96315
rect 367 96284 438 96318
rect 400 96277 404 96284
rect 454 96271 504 96273
rect 494 96267 548 96271
rect 494 96262 514 96267
rect 504 96247 506 96262
rect 196 96237 232 96241
rect 196 96207 204 96237
rect 216 96207 232 96237
rect 400 96239 404 96247
rect 107 96167 119 96173
rect 109 96139 119 96167
rect 129 96139 149 96173
rect 174 96169 181 96199
rect 224 96160 226 96207
rect 256 96199 328 96207
rect 332 96205 336 96235
rect 400 96205 408 96239
rect 434 96205 438 96239
rect 498 96237 506 96247
rect 514 96237 515 96257
rect 504 96221 506 96237
rect 525 96228 528 96262
rect 547 96237 548 96257
rect 557 96237 564 96247
rect 514 96221 530 96227
rect 532 96221 548 96227
rect 278 96169 305 96180
rect 42 96047 46 96081
rect 72 96047 76 96081
rect 38 96009 80 96010
rect 42 95968 76 96002
rect 79 95968 113 96002
rect 42 95889 46 95923
rect 72 95889 76 95923
rect -25 95852 25 95854
rect -8 95844 14 95851
rect -8 95843 17 95844
rect 25 95843 27 95852
rect -12 95836 38 95843
rect -12 95835 34 95836
rect -12 95831 8 95835
rect 0 95819 8 95831
rect 14 95819 34 95835
rect 0 95818 34 95819
rect 0 95811 38 95818
rect 14 95810 17 95811
rect 25 95802 27 95811
rect 42 95782 45 95872
rect 71 95841 80 95869
rect 69 95803 80 95841
rect 144 95831 148 96139
rect 196 96126 204 96160
rect 216 96126 232 96160
rect 244 96156 257 96160
rect 300 96156 308 96169
rect 332 96167 342 96205
rect 400 96197 404 96205
rect 336 96157 342 96167
rect 244 96132 291 96156
rect 244 96126 257 96132
rect 224 96079 226 96126
rect 278 96122 291 96132
rect 300 96132 329 96156
rect 332 96147 342 96157
rect 400 96157 409 96185
rect 562 96168 612 96170
rect 466 96159 497 96167
rect 565 96159 596 96167
rect 300 96122 321 96132
rect 300 96116 308 96122
rect 289 96106 308 96116
rect 196 96049 204 96079
rect 216 96049 232 96079
rect 196 96045 232 96049
rect 196 96037 226 96045
rect 300 96037 308 96106
rect 332 96113 351 96147
rect 361 96119 381 96147
rect 361 96113 375 96119
rect 400 96113 411 96157
rect 442 96152 500 96159
rect 466 96151 500 96152
rect 565 96151 599 96159
rect 497 96135 500 96151
rect 596 96135 599 96151
rect 466 96134 500 96135
rect 442 96127 500 96134
rect 565 96127 599 96135
rect 612 96118 614 96168
rect 332 96089 342 96113
rect 336 96077 342 96089
rect 224 96021 226 96037
rect 332 96009 342 96077
rect 400 96081 404 96089
rect 400 96047 408 96081
rect 434 96047 438 96081
rect 454 96065 504 96067
rect 504 96049 506 96065
rect 514 96059 530 96065
rect 532 96059 548 96065
rect 525 96049 548 96058
rect 400 96039 404 96047
rect 498 96039 506 96049
rect 504 96015 506 96039
rect 514 96029 515 96049
rect 525 96024 528 96049
rect 547 96029 548 96049
rect 557 96039 564 96049
rect 514 96015 548 96019
rect 151 95968 156 96002
rect 174 95999 246 96007
rect 256 95999 328 96007
rect 336 96001 342 96009
rect 400 96004 404 96009
rect 180 95971 185 95999
rect 174 95963 246 95971
rect 256 95963 328 95971
rect 332 95969 336 95999
rect 400 95970 438 96004
rect 224 95933 226 95949
rect 196 95925 226 95933
rect 196 95921 232 95925
rect 196 95891 204 95921
rect 216 95891 232 95921
rect 224 95844 226 95891
rect 300 95864 308 95933
rect 332 95931 342 95969
rect 400 95961 404 95970
rect 454 95955 504 95957
rect 494 95951 548 95955
rect 494 95946 514 95951
rect 504 95931 506 95946
rect 336 95919 342 95931
rect 289 95854 308 95864
rect 300 95848 308 95854
rect 332 95885 342 95919
rect 400 95923 404 95931
rect 400 95889 408 95923
rect 434 95889 438 95923
rect 498 95921 506 95931
rect 514 95921 515 95941
rect 504 95905 506 95921
rect 525 95912 528 95946
rect 547 95921 548 95941
rect 557 95921 564 95931
rect 514 95905 530 95911
rect 532 95905 548 95911
rect 332 95857 373 95885
rect 332 95851 351 95857
rect 107 95797 119 95831
rect 129 95797 149 95831
rect 196 95810 204 95844
rect 216 95810 232 95844
rect 244 95838 257 95844
rect 278 95838 291 95848
rect 244 95814 291 95838
rect 300 95838 321 95848
rect 336 95841 351 95851
rect 300 95814 329 95838
rect 332 95823 351 95841
rect 361 95851 375 95857
rect 400 95851 411 95889
rect 562 95852 612 95854
rect 361 95823 381 95851
rect 400 95823 409 95851
rect 466 95843 497 95851
rect 565 95843 596 95851
rect 442 95836 500 95843
rect 466 95835 500 95836
rect 565 95835 599 95843
rect 244 95810 257 95814
rect 42 95731 46 95765
rect 72 95731 76 95765
rect 42 95684 76 95688
rect 42 95669 46 95684
rect 72 95669 76 95684
rect 38 95651 80 95669
rect 16 95645 102 95651
rect 144 95645 148 95797
rect 174 95773 181 95801
rect 224 95763 226 95810
rect 300 95801 308 95814
rect 278 95790 305 95801
rect 332 95773 342 95823
rect 400 95803 404 95823
rect 497 95819 500 95835
rect 596 95819 599 95835
rect 466 95818 500 95819
rect 442 95811 500 95818
rect 565 95811 599 95819
rect 612 95802 614 95852
rect 256 95763 328 95771
rect 336 95765 342 95773
rect 400 95765 404 95773
rect 196 95733 204 95763
rect 216 95733 232 95763
rect 196 95729 232 95733
rect 196 95721 226 95729
rect 224 95705 226 95721
rect 332 95693 336 95761
rect 400 95731 408 95765
rect 434 95731 438 95765
rect 454 95749 504 95751
rect 504 95733 506 95749
rect 514 95743 530 95749
rect 532 95743 548 95749
rect 525 95733 548 95742
rect 400 95723 404 95731
rect 498 95723 506 95733
rect 504 95699 506 95723
rect 514 95713 515 95733
rect 525 95708 528 95733
rect 547 95713 548 95733
rect 557 95723 564 95733
rect 514 95699 548 95703
rect 400 95693 442 95694
rect 174 95683 246 95691
rect 400 95686 404 95693
rect 295 95652 300 95686
rect 324 95652 329 95686
rect 367 95669 438 95686
rect 367 95652 442 95669
rect 400 95651 442 95652
rect 378 95645 464 95651
rect 38 95629 80 95645
rect 400 95629 442 95645
rect -25 95615 25 95617
rect 42 95615 76 95629
rect 404 95615 438 95629
rect 455 95615 505 95617
rect 557 95615 607 95617
rect 16 95607 102 95615
rect 378 95607 464 95615
rect 8 95573 17 95607
rect 18 95605 51 95607
rect 80 95605 100 95607
rect 18 95573 100 95605
rect 380 95605 404 95607
rect 429 95605 438 95607
rect 442 95605 462 95607
rect 16 95565 102 95573
rect 42 95549 76 95565
rect 16 95529 38 95535
rect 42 95526 76 95530
rect 80 95529 102 95535
rect 42 95496 46 95526
rect 72 95496 76 95526
rect 42 95415 46 95449
rect 72 95415 76 95449
rect -25 95378 25 95380
rect -8 95370 14 95377
rect -8 95369 17 95370
rect 25 95369 27 95378
rect -12 95362 38 95369
rect -12 95361 34 95362
rect -12 95357 8 95361
rect 0 95345 8 95357
rect 14 95345 34 95361
rect 0 95344 34 95345
rect 0 95337 38 95344
rect 14 95336 17 95337
rect 25 95328 27 95337
rect 42 95308 45 95398
rect 69 95383 80 95415
rect 107 95383 143 95411
rect 144 95383 148 95603
rect 332 95535 336 95603
rect 380 95573 462 95605
rect 463 95573 472 95607
rect 480 95573 497 95607
rect 378 95565 464 95573
rect 505 95565 507 95615
rect 514 95573 548 95607
rect 565 95573 582 95607
rect 607 95565 609 95615
rect 404 95549 438 95565
rect 400 95535 442 95536
rect 378 95529 404 95535
rect 442 95529 464 95535
rect 400 95528 404 95529
rect 174 95489 246 95497
rect 295 95494 300 95528
rect 324 95494 329 95528
rect 224 95459 226 95475
rect 196 95451 226 95459
rect 332 95457 336 95525
rect 367 95494 438 95528
rect 400 95487 404 95494
rect 454 95481 504 95483
rect 494 95477 548 95481
rect 494 95472 514 95477
rect 504 95457 506 95472
rect 196 95447 232 95451
rect 196 95417 204 95447
rect 216 95417 232 95447
rect 400 95449 404 95457
rect 107 95377 119 95383
rect 109 95349 119 95377
rect 129 95349 149 95383
rect 174 95379 181 95409
rect 224 95370 226 95417
rect 256 95409 328 95417
rect 332 95415 336 95445
rect 400 95415 408 95449
rect 434 95415 438 95449
rect 498 95447 506 95457
rect 514 95447 515 95467
rect 504 95431 506 95447
rect 525 95438 528 95472
rect 547 95447 548 95467
rect 557 95447 564 95457
rect 514 95431 530 95437
rect 532 95431 548 95437
rect 278 95379 305 95390
rect 42 95257 46 95291
rect 72 95257 76 95291
rect 38 95219 80 95220
rect 42 95178 76 95212
rect 79 95178 113 95212
rect 42 95099 46 95133
rect 72 95099 76 95133
rect -25 95062 25 95064
rect -8 95054 14 95061
rect -8 95053 17 95054
rect 25 95053 27 95062
rect -12 95046 38 95053
rect -12 95045 34 95046
rect -12 95041 8 95045
rect 0 95029 8 95041
rect 14 95029 34 95045
rect 0 95028 34 95029
rect 0 95021 38 95028
rect 14 95020 17 95021
rect 25 95012 27 95021
rect 42 94992 45 95082
rect 71 95051 80 95079
rect 69 95013 80 95051
rect 144 95041 148 95349
rect 196 95336 204 95370
rect 216 95336 232 95370
rect 244 95366 257 95370
rect 300 95366 308 95379
rect 332 95377 342 95415
rect 400 95407 404 95415
rect 336 95367 342 95377
rect 244 95342 291 95366
rect 244 95336 257 95342
rect 224 95289 226 95336
rect 278 95332 291 95342
rect 300 95342 329 95366
rect 332 95357 342 95367
rect 400 95367 409 95395
rect 562 95378 612 95380
rect 466 95369 497 95377
rect 565 95369 596 95377
rect 300 95332 321 95342
rect 300 95326 308 95332
rect 289 95316 308 95326
rect 196 95259 204 95289
rect 216 95259 232 95289
rect 196 95255 232 95259
rect 196 95247 226 95255
rect 300 95247 308 95316
rect 332 95323 351 95357
rect 361 95329 381 95357
rect 361 95323 375 95329
rect 400 95323 411 95367
rect 442 95362 500 95369
rect 466 95361 500 95362
rect 565 95361 599 95369
rect 497 95345 500 95361
rect 596 95345 599 95361
rect 466 95344 500 95345
rect 442 95337 500 95344
rect 565 95337 599 95345
rect 612 95328 614 95378
rect 332 95299 342 95323
rect 336 95287 342 95299
rect 224 95231 226 95247
rect 332 95219 342 95287
rect 400 95291 404 95299
rect 400 95257 408 95291
rect 434 95257 438 95291
rect 454 95275 504 95277
rect 504 95259 506 95275
rect 514 95269 530 95275
rect 532 95269 548 95275
rect 525 95259 548 95268
rect 400 95249 404 95257
rect 498 95249 506 95259
rect 504 95225 506 95249
rect 514 95239 515 95259
rect 525 95234 528 95259
rect 547 95239 548 95259
rect 557 95249 564 95259
rect 514 95225 548 95229
rect 151 95178 156 95212
rect 174 95209 246 95217
rect 256 95209 328 95217
rect 336 95211 342 95219
rect 400 95214 404 95219
rect 180 95181 185 95209
rect 174 95173 246 95181
rect 256 95173 328 95181
rect 332 95179 336 95209
rect 400 95180 438 95214
rect 224 95143 226 95159
rect 196 95135 226 95143
rect 196 95131 232 95135
rect 196 95101 204 95131
rect 216 95101 232 95131
rect 224 95054 226 95101
rect 300 95074 308 95143
rect 332 95141 342 95179
rect 400 95171 404 95180
rect 454 95165 504 95167
rect 494 95161 548 95165
rect 494 95156 514 95161
rect 504 95141 506 95156
rect 336 95129 342 95141
rect 289 95064 308 95074
rect 300 95058 308 95064
rect 332 95095 342 95129
rect 400 95133 404 95141
rect 400 95099 408 95133
rect 434 95099 438 95133
rect 498 95131 506 95141
rect 514 95131 515 95151
rect 504 95115 506 95131
rect 525 95122 528 95156
rect 547 95131 548 95151
rect 557 95131 564 95141
rect 514 95115 530 95121
rect 532 95115 548 95121
rect 332 95067 373 95095
rect 332 95061 351 95067
rect 107 95007 119 95041
rect 129 95007 149 95041
rect 196 95020 204 95054
rect 216 95020 232 95054
rect 244 95048 257 95054
rect 278 95048 291 95058
rect 244 95024 291 95048
rect 300 95048 321 95058
rect 336 95051 351 95061
rect 300 95024 329 95048
rect 332 95033 351 95051
rect 361 95061 375 95067
rect 400 95061 411 95099
rect 562 95062 612 95064
rect 361 95033 381 95061
rect 400 95033 409 95061
rect 466 95053 497 95061
rect 565 95053 596 95061
rect 442 95046 500 95053
rect 466 95045 500 95046
rect 565 95045 599 95053
rect 244 95020 257 95024
rect 42 94941 46 94975
rect 72 94941 76 94975
rect 42 94894 76 94898
rect 42 94879 46 94894
rect 72 94879 76 94894
rect 38 94861 80 94879
rect 16 94855 102 94861
rect 144 94855 148 95007
rect 174 94983 181 95011
rect 224 94973 226 95020
rect 300 95011 308 95024
rect 278 95000 305 95011
rect 332 94983 342 95033
rect 400 95013 404 95033
rect 497 95029 500 95045
rect 596 95029 599 95045
rect 466 95028 500 95029
rect 442 95021 500 95028
rect 565 95021 599 95029
rect 612 95012 614 95062
rect 256 94973 328 94981
rect 336 94975 342 94983
rect 400 94975 404 94983
rect 196 94943 204 94973
rect 216 94943 232 94973
rect 196 94939 232 94943
rect 196 94931 226 94939
rect 224 94915 226 94931
rect 332 94903 336 94971
rect 400 94941 408 94975
rect 434 94941 438 94975
rect 454 94959 504 94961
rect 504 94943 506 94959
rect 514 94953 530 94959
rect 532 94953 548 94959
rect 525 94943 548 94952
rect 400 94933 404 94941
rect 498 94933 506 94943
rect 504 94909 506 94933
rect 514 94923 515 94943
rect 525 94918 528 94943
rect 547 94923 548 94943
rect 557 94933 564 94943
rect 514 94909 548 94913
rect 400 94903 442 94904
rect 174 94893 246 94901
rect 400 94896 404 94903
rect 295 94862 300 94896
rect 324 94862 329 94896
rect 367 94879 438 94896
rect 367 94862 442 94879
rect 400 94861 442 94862
rect 378 94855 464 94861
rect 38 94839 80 94855
rect 400 94839 442 94855
rect -25 94825 25 94827
rect 42 94825 76 94839
rect 404 94825 438 94839
rect 455 94825 505 94827
rect 557 94825 607 94827
rect 16 94817 102 94825
rect 378 94817 464 94825
rect 8 94783 17 94817
rect 18 94815 51 94817
rect 80 94815 100 94817
rect 18 94783 100 94815
rect 380 94815 404 94817
rect 429 94815 438 94817
rect 442 94815 462 94817
rect 16 94775 102 94783
rect 42 94759 76 94775
rect 16 94739 38 94745
rect 42 94736 76 94740
rect 80 94739 102 94745
rect 42 94706 46 94736
rect 72 94706 76 94736
rect 42 94625 46 94659
rect 72 94625 76 94659
rect -25 94588 25 94590
rect -8 94580 14 94587
rect -8 94579 17 94580
rect 25 94579 27 94588
rect -12 94572 38 94579
rect -12 94571 34 94572
rect -12 94567 8 94571
rect 0 94555 8 94567
rect 14 94555 34 94571
rect 0 94554 34 94555
rect 0 94547 38 94554
rect 14 94546 17 94547
rect 25 94538 27 94547
rect 42 94518 45 94608
rect 69 94593 80 94625
rect 107 94593 143 94621
rect 144 94593 148 94813
rect 332 94745 336 94813
rect 380 94783 462 94815
rect 463 94783 472 94817
rect 480 94783 497 94817
rect 378 94775 464 94783
rect 505 94775 507 94825
rect 514 94783 548 94817
rect 565 94783 582 94817
rect 607 94775 609 94825
rect 404 94759 438 94775
rect 400 94745 442 94746
rect 378 94739 404 94745
rect 442 94739 464 94745
rect 400 94738 404 94739
rect 174 94699 246 94707
rect 295 94704 300 94738
rect 324 94704 329 94738
rect 224 94669 226 94685
rect 196 94661 226 94669
rect 332 94667 336 94735
rect 367 94704 438 94738
rect 400 94697 404 94704
rect 454 94691 504 94693
rect 494 94687 548 94691
rect 494 94682 514 94687
rect 504 94667 506 94682
rect 196 94657 232 94661
rect 196 94627 204 94657
rect 216 94627 232 94657
rect 400 94659 404 94667
rect 107 94587 119 94593
rect 109 94559 119 94587
rect 129 94559 149 94593
rect 174 94589 181 94619
rect 224 94580 226 94627
rect 256 94619 328 94627
rect 332 94625 336 94655
rect 400 94625 408 94659
rect 434 94625 438 94659
rect 498 94657 506 94667
rect 514 94657 515 94677
rect 504 94641 506 94657
rect 525 94648 528 94682
rect 547 94657 548 94677
rect 557 94657 564 94667
rect 514 94641 530 94647
rect 532 94641 548 94647
rect 278 94589 305 94600
rect 42 94467 46 94501
rect 72 94467 76 94501
rect 38 94429 80 94430
rect 42 94388 76 94422
rect 79 94388 113 94422
rect 42 94309 46 94343
rect 72 94309 76 94343
rect -25 94272 25 94274
rect -8 94264 14 94271
rect -8 94263 17 94264
rect 25 94263 27 94272
rect -12 94256 38 94263
rect -12 94255 34 94256
rect -12 94251 8 94255
rect 0 94239 8 94251
rect 14 94239 34 94255
rect 0 94238 34 94239
rect 0 94231 38 94238
rect 14 94230 17 94231
rect 25 94222 27 94231
rect 42 94202 45 94292
rect 71 94261 80 94289
rect 69 94223 80 94261
rect 144 94251 148 94559
rect 196 94546 204 94580
rect 216 94546 232 94580
rect 244 94576 257 94580
rect 300 94576 308 94589
rect 332 94587 342 94625
rect 400 94617 404 94625
rect 336 94577 342 94587
rect 244 94552 291 94576
rect 244 94546 257 94552
rect 224 94499 226 94546
rect 278 94542 291 94552
rect 300 94552 329 94576
rect 332 94567 342 94577
rect 400 94577 409 94605
rect 562 94588 612 94590
rect 466 94579 497 94587
rect 565 94579 596 94587
rect 300 94542 321 94552
rect 300 94536 308 94542
rect 289 94526 308 94536
rect 196 94469 204 94499
rect 216 94469 232 94499
rect 196 94465 232 94469
rect 196 94457 226 94465
rect 300 94457 308 94526
rect 332 94533 351 94567
rect 361 94539 381 94567
rect 361 94533 375 94539
rect 400 94533 411 94577
rect 442 94572 500 94579
rect 466 94571 500 94572
rect 565 94571 599 94579
rect 497 94555 500 94571
rect 596 94555 599 94571
rect 466 94554 500 94555
rect 442 94547 500 94554
rect 565 94547 599 94555
rect 612 94538 614 94588
rect 332 94509 342 94533
rect 336 94497 342 94509
rect 224 94441 226 94457
rect 332 94429 342 94497
rect 400 94501 404 94509
rect 400 94467 408 94501
rect 434 94467 438 94501
rect 454 94485 504 94487
rect 504 94469 506 94485
rect 514 94479 530 94485
rect 532 94479 548 94485
rect 525 94469 548 94478
rect 400 94459 404 94467
rect 498 94459 506 94469
rect 504 94435 506 94459
rect 514 94449 515 94469
rect 525 94444 528 94469
rect 547 94449 548 94469
rect 557 94459 564 94469
rect 514 94435 548 94439
rect 151 94388 156 94422
rect 174 94419 246 94427
rect 256 94419 328 94427
rect 336 94421 342 94429
rect 400 94424 404 94429
rect 180 94391 185 94419
rect 174 94383 246 94391
rect 256 94383 328 94391
rect 332 94389 336 94419
rect 400 94390 438 94424
rect 224 94353 226 94369
rect 196 94345 226 94353
rect 196 94341 232 94345
rect 196 94311 204 94341
rect 216 94311 232 94341
rect 224 94264 226 94311
rect 300 94284 308 94353
rect 332 94351 342 94389
rect 400 94381 404 94390
rect 454 94375 504 94377
rect 494 94371 548 94375
rect 494 94366 514 94371
rect 504 94351 506 94366
rect 336 94339 342 94351
rect 289 94274 308 94284
rect 300 94268 308 94274
rect 332 94305 342 94339
rect 400 94343 404 94351
rect 400 94309 408 94343
rect 434 94309 438 94343
rect 498 94341 506 94351
rect 514 94341 515 94361
rect 504 94325 506 94341
rect 525 94332 528 94366
rect 547 94341 548 94361
rect 557 94341 564 94351
rect 514 94325 530 94331
rect 532 94325 548 94331
rect 332 94277 373 94305
rect 332 94271 351 94277
rect 107 94217 119 94251
rect 129 94217 149 94251
rect 196 94230 204 94264
rect 216 94230 232 94264
rect 244 94258 257 94264
rect 278 94258 291 94268
rect 244 94234 291 94258
rect 300 94258 321 94268
rect 336 94261 351 94271
rect 300 94234 329 94258
rect 332 94243 351 94261
rect 361 94271 375 94277
rect 400 94271 411 94309
rect 562 94272 612 94274
rect 361 94243 381 94271
rect 400 94243 409 94271
rect 466 94263 497 94271
rect 565 94263 596 94271
rect 442 94256 500 94263
rect 466 94255 500 94256
rect 565 94255 599 94263
rect 244 94230 257 94234
rect 42 94151 46 94185
rect 72 94151 76 94185
rect 42 94104 76 94108
rect 42 94089 46 94104
rect 72 94089 76 94104
rect 38 94071 80 94089
rect 16 94065 102 94071
rect 144 94065 148 94217
rect 174 94193 181 94221
rect 224 94183 226 94230
rect 300 94221 308 94234
rect 278 94210 305 94221
rect 332 94193 342 94243
rect 400 94223 404 94243
rect 497 94239 500 94255
rect 596 94239 599 94255
rect 466 94238 500 94239
rect 442 94231 500 94238
rect 565 94231 599 94239
rect 612 94222 614 94272
rect 256 94183 328 94191
rect 336 94185 342 94193
rect 400 94185 404 94193
rect 196 94153 204 94183
rect 216 94153 232 94183
rect 196 94149 232 94153
rect 196 94141 226 94149
rect 224 94125 226 94141
rect 332 94113 336 94181
rect 400 94151 408 94185
rect 434 94151 438 94185
rect 454 94169 504 94171
rect 504 94153 506 94169
rect 514 94163 530 94169
rect 532 94163 548 94169
rect 525 94153 548 94162
rect 400 94143 404 94151
rect 498 94143 506 94153
rect 504 94119 506 94143
rect 514 94133 515 94153
rect 525 94128 528 94153
rect 547 94133 548 94153
rect 557 94143 564 94153
rect 514 94119 548 94123
rect 400 94113 442 94114
rect 174 94103 246 94111
rect 400 94106 404 94113
rect 295 94072 300 94106
rect 324 94072 329 94106
rect 367 94089 438 94106
rect 367 94072 442 94089
rect 400 94071 442 94072
rect 378 94065 464 94071
rect 38 94049 80 94065
rect 400 94049 442 94065
rect -25 94035 25 94037
rect 42 94035 76 94049
rect 404 94035 438 94049
rect 455 94035 505 94037
rect 557 94035 607 94037
rect 16 94027 102 94035
rect 378 94027 464 94035
rect 8 93993 17 94027
rect 18 94025 51 94027
rect 80 94025 100 94027
rect 18 93993 100 94025
rect 380 94025 404 94027
rect 429 94025 438 94027
rect 442 94025 462 94027
rect 16 93985 102 93993
rect 42 93969 76 93985
rect 16 93949 38 93955
rect 42 93946 76 93950
rect 80 93949 102 93955
rect 42 93916 46 93946
rect 72 93916 76 93946
rect 42 93835 46 93869
rect 72 93835 76 93869
rect -25 93798 25 93800
rect -8 93790 14 93797
rect -8 93789 17 93790
rect 25 93789 27 93798
rect -12 93782 38 93789
rect -12 93781 34 93782
rect -12 93777 8 93781
rect 0 93765 8 93777
rect 14 93765 34 93781
rect 0 93764 34 93765
rect 0 93757 38 93764
rect 14 93756 17 93757
rect 25 93748 27 93757
rect 42 93728 45 93818
rect 69 93803 80 93835
rect 107 93803 143 93831
rect 144 93803 148 94023
rect 332 93955 336 94023
rect 380 93993 462 94025
rect 463 93993 472 94027
rect 480 93993 497 94027
rect 378 93985 464 93993
rect 505 93985 507 94035
rect 514 93993 548 94027
rect 565 93993 582 94027
rect 607 93985 609 94035
rect 404 93969 438 93985
rect 400 93955 442 93956
rect 378 93949 404 93955
rect 442 93949 464 93955
rect 400 93948 404 93949
rect 174 93909 246 93917
rect 295 93914 300 93948
rect 324 93914 329 93948
rect 224 93879 226 93895
rect 196 93871 226 93879
rect 332 93877 336 93945
rect 367 93914 438 93948
rect 400 93907 404 93914
rect 454 93901 504 93903
rect 494 93897 548 93901
rect 494 93892 514 93897
rect 504 93877 506 93892
rect 196 93867 232 93871
rect 196 93837 204 93867
rect 216 93837 232 93867
rect 400 93869 404 93877
rect 107 93797 119 93803
rect 109 93769 119 93797
rect 129 93769 149 93803
rect 174 93799 181 93829
rect 224 93790 226 93837
rect 256 93829 328 93837
rect 332 93835 336 93865
rect 400 93835 408 93869
rect 434 93835 438 93869
rect 498 93867 506 93877
rect 514 93867 515 93887
rect 504 93851 506 93867
rect 525 93858 528 93892
rect 547 93867 548 93887
rect 557 93867 564 93877
rect 514 93851 530 93857
rect 532 93851 548 93857
rect 278 93799 305 93810
rect 42 93677 46 93711
rect 72 93677 76 93711
rect 38 93639 80 93640
rect 42 93598 76 93632
rect 79 93598 113 93632
rect 42 93519 46 93553
rect 72 93519 76 93553
rect -25 93482 25 93484
rect -8 93474 14 93481
rect -8 93473 17 93474
rect 25 93473 27 93482
rect -12 93466 38 93473
rect -12 93465 34 93466
rect -12 93461 8 93465
rect 0 93449 8 93461
rect 14 93449 34 93465
rect 0 93448 34 93449
rect 0 93441 38 93448
rect 14 93440 17 93441
rect 25 93432 27 93441
rect 42 93412 45 93502
rect 71 93471 80 93499
rect 69 93433 80 93471
rect 144 93461 148 93769
rect 196 93756 204 93790
rect 216 93756 232 93790
rect 244 93786 257 93790
rect 300 93786 308 93799
rect 332 93797 342 93835
rect 400 93827 404 93835
rect 336 93787 342 93797
rect 244 93762 291 93786
rect 244 93756 257 93762
rect 224 93709 226 93756
rect 278 93752 291 93762
rect 300 93762 329 93786
rect 332 93777 342 93787
rect 400 93787 409 93815
rect 562 93798 612 93800
rect 466 93789 497 93797
rect 565 93789 596 93797
rect 300 93752 321 93762
rect 300 93746 308 93752
rect 289 93736 308 93746
rect 196 93679 204 93709
rect 216 93679 232 93709
rect 196 93675 232 93679
rect 196 93667 226 93675
rect 300 93667 308 93736
rect 332 93743 351 93777
rect 361 93749 381 93777
rect 361 93743 375 93749
rect 400 93743 411 93787
rect 442 93782 500 93789
rect 466 93781 500 93782
rect 565 93781 599 93789
rect 497 93765 500 93781
rect 596 93765 599 93781
rect 466 93764 500 93765
rect 442 93757 500 93764
rect 565 93757 599 93765
rect 612 93748 614 93798
rect 332 93719 342 93743
rect 336 93707 342 93719
rect 224 93651 226 93667
rect 332 93639 342 93707
rect 400 93711 404 93719
rect 400 93677 408 93711
rect 434 93677 438 93711
rect 454 93695 504 93697
rect 504 93679 506 93695
rect 514 93689 530 93695
rect 532 93689 548 93695
rect 525 93679 548 93688
rect 400 93669 404 93677
rect 498 93669 506 93679
rect 504 93645 506 93669
rect 514 93659 515 93679
rect 525 93654 528 93679
rect 547 93659 548 93679
rect 557 93669 564 93679
rect 514 93645 548 93649
rect 151 93598 156 93632
rect 174 93629 246 93637
rect 256 93629 328 93637
rect 336 93631 342 93639
rect 400 93634 404 93639
rect 180 93601 185 93629
rect 174 93593 246 93601
rect 256 93593 328 93601
rect 332 93599 336 93629
rect 400 93600 438 93634
rect 224 93563 226 93579
rect 196 93555 226 93563
rect 196 93551 232 93555
rect 196 93521 204 93551
rect 216 93521 232 93551
rect 224 93474 226 93521
rect 300 93494 308 93563
rect 332 93561 342 93599
rect 400 93591 404 93600
rect 454 93585 504 93587
rect 494 93581 548 93585
rect 494 93576 514 93581
rect 504 93561 506 93576
rect 336 93549 342 93561
rect 289 93484 308 93494
rect 300 93478 308 93484
rect 332 93515 342 93549
rect 400 93553 404 93561
rect 400 93519 408 93553
rect 434 93519 438 93553
rect 498 93551 506 93561
rect 514 93551 515 93571
rect 504 93535 506 93551
rect 525 93542 528 93576
rect 547 93551 548 93571
rect 557 93551 564 93561
rect 514 93535 530 93541
rect 532 93535 548 93541
rect 332 93487 373 93515
rect 332 93481 351 93487
rect 107 93427 119 93461
rect 129 93427 149 93461
rect 196 93440 204 93474
rect 216 93440 232 93474
rect 244 93468 257 93474
rect 278 93468 291 93478
rect 244 93444 291 93468
rect 300 93468 321 93478
rect 336 93471 351 93481
rect 300 93444 329 93468
rect 332 93453 351 93471
rect 361 93481 375 93487
rect 400 93481 411 93519
rect 562 93482 612 93484
rect 361 93453 381 93481
rect 400 93453 409 93481
rect 466 93473 497 93481
rect 565 93473 596 93481
rect 442 93466 500 93473
rect 466 93465 500 93466
rect 565 93465 599 93473
rect 244 93440 257 93444
rect 42 93361 46 93395
rect 72 93361 76 93395
rect 42 93314 76 93318
rect 42 93299 46 93314
rect 72 93299 76 93314
rect 38 93281 80 93299
rect 16 93275 102 93281
rect 144 93275 148 93427
rect 174 93403 181 93431
rect 224 93393 226 93440
rect 300 93431 308 93444
rect 278 93420 305 93431
rect 332 93403 342 93453
rect 400 93433 404 93453
rect 497 93449 500 93465
rect 596 93449 599 93465
rect 466 93448 500 93449
rect 442 93441 500 93448
rect 565 93441 599 93449
rect 612 93432 614 93482
rect 256 93393 328 93401
rect 336 93395 342 93403
rect 400 93395 404 93403
rect 196 93363 204 93393
rect 216 93363 232 93393
rect 196 93359 232 93363
rect 196 93351 226 93359
rect 224 93335 226 93351
rect 332 93323 336 93391
rect 400 93361 408 93395
rect 434 93361 438 93395
rect 454 93379 504 93381
rect 504 93363 506 93379
rect 514 93373 530 93379
rect 532 93373 548 93379
rect 525 93363 548 93372
rect 400 93353 404 93361
rect 498 93353 506 93363
rect 504 93329 506 93353
rect 514 93343 515 93363
rect 525 93338 528 93363
rect 547 93343 548 93363
rect 557 93353 564 93363
rect 514 93329 548 93333
rect 400 93323 442 93324
rect 174 93313 246 93321
rect 400 93316 404 93323
rect 295 93282 300 93316
rect 324 93282 329 93316
rect 367 93299 438 93316
rect 367 93282 442 93299
rect 400 93281 442 93282
rect 378 93275 464 93281
rect 38 93259 80 93275
rect 400 93259 442 93275
rect -25 93245 25 93247
rect 42 93245 76 93259
rect 404 93245 438 93259
rect 455 93245 505 93247
rect 557 93245 607 93247
rect 16 93237 102 93245
rect 378 93237 464 93245
rect 8 93203 17 93237
rect 18 93235 51 93237
rect 80 93235 100 93237
rect 18 93203 100 93235
rect 380 93235 404 93237
rect 429 93235 438 93237
rect 442 93235 462 93237
rect 16 93195 102 93203
rect 42 93179 76 93195
rect 16 93159 38 93165
rect 42 93156 76 93160
rect 80 93159 102 93165
rect 42 93126 46 93156
rect 72 93126 76 93156
rect 42 93045 46 93079
rect 72 93045 76 93079
rect -25 93008 25 93010
rect -8 93000 14 93007
rect -8 92999 17 93000
rect 25 92999 27 93008
rect -12 92992 38 92999
rect -12 92991 34 92992
rect -12 92987 8 92991
rect 0 92975 8 92987
rect 14 92975 34 92991
rect 0 92974 34 92975
rect 0 92967 38 92974
rect 14 92966 17 92967
rect 25 92958 27 92967
rect 42 92938 45 93028
rect 69 93013 80 93045
rect 107 93013 143 93041
rect 144 93013 148 93233
rect 332 93165 336 93233
rect 380 93203 462 93235
rect 463 93203 472 93237
rect 480 93203 497 93237
rect 378 93195 464 93203
rect 505 93195 507 93245
rect 514 93203 548 93237
rect 565 93203 582 93237
rect 607 93195 609 93245
rect 404 93179 438 93195
rect 400 93165 442 93166
rect 378 93159 404 93165
rect 442 93159 464 93165
rect 400 93158 404 93159
rect 174 93119 246 93127
rect 295 93124 300 93158
rect 324 93124 329 93158
rect 224 93089 226 93105
rect 196 93081 226 93089
rect 332 93087 336 93155
rect 367 93124 438 93158
rect 400 93117 404 93124
rect 454 93111 504 93113
rect 494 93107 548 93111
rect 494 93102 514 93107
rect 504 93087 506 93102
rect 196 93077 232 93081
rect 196 93047 204 93077
rect 216 93047 232 93077
rect 400 93079 404 93087
rect 107 93007 119 93013
rect 109 92979 119 93007
rect 129 92979 149 93013
rect 174 93009 181 93039
rect 224 93000 226 93047
rect 256 93039 328 93047
rect 332 93045 336 93075
rect 400 93045 408 93079
rect 434 93045 438 93079
rect 498 93077 506 93087
rect 514 93077 515 93097
rect 504 93061 506 93077
rect 525 93068 528 93102
rect 547 93077 548 93097
rect 557 93077 564 93087
rect 514 93061 530 93067
rect 532 93061 548 93067
rect 278 93009 305 93020
rect 42 92887 46 92921
rect 72 92887 76 92921
rect 38 92849 80 92850
rect 42 92808 76 92842
rect 79 92808 113 92842
rect 42 92729 46 92763
rect 72 92729 76 92763
rect -25 92692 25 92694
rect -8 92684 14 92691
rect -8 92683 17 92684
rect 25 92683 27 92692
rect -12 92676 38 92683
rect -12 92675 34 92676
rect -12 92671 8 92675
rect 0 92659 8 92671
rect 14 92659 34 92675
rect 0 92658 34 92659
rect 0 92651 38 92658
rect 14 92650 17 92651
rect 25 92642 27 92651
rect 42 92622 45 92712
rect 71 92681 80 92709
rect 69 92643 80 92681
rect 144 92671 148 92979
rect 196 92966 204 93000
rect 216 92966 232 93000
rect 244 92996 257 93000
rect 300 92996 308 93009
rect 332 93007 342 93045
rect 400 93037 404 93045
rect 336 92997 342 93007
rect 244 92972 291 92996
rect 244 92966 257 92972
rect 224 92919 226 92966
rect 278 92962 291 92972
rect 300 92972 329 92996
rect 332 92987 342 92997
rect 400 92997 409 93025
rect 562 93008 612 93010
rect 466 92999 497 93007
rect 565 92999 596 93007
rect 300 92962 321 92972
rect 300 92956 308 92962
rect 289 92946 308 92956
rect 196 92889 204 92919
rect 216 92889 232 92919
rect 196 92885 232 92889
rect 196 92877 226 92885
rect 300 92877 308 92946
rect 332 92953 351 92987
rect 361 92959 381 92987
rect 361 92953 375 92959
rect 400 92953 411 92997
rect 442 92992 500 92999
rect 466 92991 500 92992
rect 565 92991 599 92999
rect 497 92975 500 92991
rect 596 92975 599 92991
rect 466 92974 500 92975
rect 442 92967 500 92974
rect 565 92967 599 92975
rect 612 92958 614 93008
rect 332 92929 342 92953
rect 336 92917 342 92929
rect 224 92861 226 92877
rect 332 92849 342 92917
rect 400 92921 404 92929
rect 400 92887 408 92921
rect 434 92887 438 92921
rect 454 92905 504 92907
rect 504 92889 506 92905
rect 514 92899 530 92905
rect 532 92899 548 92905
rect 525 92889 548 92898
rect 400 92879 404 92887
rect 498 92879 506 92889
rect 504 92855 506 92879
rect 514 92869 515 92889
rect 525 92864 528 92889
rect 547 92869 548 92889
rect 557 92879 564 92889
rect 514 92855 548 92859
rect 151 92808 156 92842
rect 174 92839 246 92847
rect 256 92839 328 92847
rect 336 92841 342 92849
rect 400 92844 404 92849
rect 180 92811 185 92839
rect 174 92803 246 92811
rect 256 92803 328 92811
rect 332 92809 336 92839
rect 400 92810 438 92844
rect 224 92773 226 92789
rect 196 92765 226 92773
rect 196 92761 232 92765
rect 196 92731 204 92761
rect 216 92731 232 92761
rect 224 92684 226 92731
rect 300 92704 308 92773
rect 332 92771 342 92809
rect 400 92801 404 92810
rect 454 92795 504 92797
rect 494 92791 548 92795
rect 494 92786 514 92791
rect 504 92771 506 92786
rect 336 92759 342 92771
rect 289 92694 308 92704
rect 300 92688 308 92694
rect 332 92725 342 92759
rect 400 92763 404 92771
rect 400 92729 408 92763
rect 434 92729 438 92763
rect 498 92761 506 92771
rect 514 92761 515 92781
rect 504 92745 506 92761
rect 525 92752 528 92786
rect 547 92761 548 92781
rect 557 92761 564 92771
rect 514 92745 530 92751
rect 532 92745 548 92751
rect 332 92697 373 92725
rect 332 92691 351 92697
rect 107 92637 119 92671
rect 129 92637 149 92671
rect 196 92650 204 92684
rect 216 92650 232 92684
rect 244 92678 257 92684
rect 278 92678 291 92688
rect 244 92654 291 92678
rect 300 92678 321 92688
rect 336 92681 351 92691
rect 300 92654 329 92678
rect 332 92663 351 92681
rect 361 92691 375 92697
rect 400 92691 411 92729
rect 562 92692 612 92694
rect 361 92663 381 92691
rect 400 92663 409 92691
rect 466 92683 497 92691
rect 565 92683 596 92691
rect 442 92676 500 92683
rect 466 92675 500 92676
rect 565 92675 599 92683
rect 244 92650 257 92654
rect 42 92571 46 92605
rect 72 92571 76 92605
rect 42 92524 76 92528
rect 42 92509 46 92524
rect 72 92509 76 92524
rect 38 92491 80 92509
rect 16 92485 102 92491
rect 144 92485 148 92637
rect 174 92613 181 92641
rect 224 92603 226 92650
rect 300 92641 308 92654
rect 278 92630 305 92641
rect 332 92613 342 92663
rect 400 92643 404 92663
rect 497 92659 500 92675
rect 596 92659 599 92675
rect 466 92658 500 92659
rect 442 92651 500 92658
rect 565 92651 599 92659
rect 612 92642 614 92692
rect 256 92603 328 92611
rect 336 92605 342 92613
rect 400 92605 404 92613
rect 196 92573 204 92603
rect 216 92573 232 92603
rect 196 92569 232 92573
rect 196 92561 226 92569
rect 224 92545 226 92561
rect 332 92533 336 92601
rect 400 92571 408 92605
rect 434 92571 438 92605
rect 454 92589 504 92591
rect 504 92573 506 92589
rect 514 92583 530 92589
rect 532 92583 548 92589
rect 525 92573 548 92582
rect 400 92563 404 92571
rect 498 92563 506 92573
rect 504 92539 506 92563
rect 514 92553 515 92573
rect 525 92548 528 92573
rect 547 92553 548 92573
rect 557 92563 564 92573
rect 514 92539 548 92543
rect 400 92533 442 92534
rect 174 92523 246 92531
rect 400 92526 404 92533
rect 295 92492 300 92526
rect 324 92492 329 92526
rect 367 92509 438 92526
rect 367 92492 442 92509
rect 400 92491 442 92492
rect 378 92485 464 92491
rect 38 92469 80 92485
rect 400 92469 442 92485
rect -25 92455 25 92457
rect 42 92455 76 92469
rect 404 92455 438 92469
rect 455 92455 505 92457
rect 557 92455 607 92457
rect 16 92447 102 92455
rect 378 92447 464 92455
rect 8 92413 17 92447
rect 18 92445 51 92447
rect 80 92445 100 92447
rect 18 92413 100 92445
rect 380 92445 404 92447
rect 429 92445 438 92447
rect 442 92445 462 92447
rect 16 92405 102 92413
rect 42 92389 76 92405
rect 16 92369 38 92375
rect 42 92366 76 92370
rect 80 92369 102 92375
rect 42 92336 46 92366
rect 72 92336 76 92366
rect 42 92255 46 92289
rect 72 92255 76 92289
rect -25 92218 25 92220
rect -8 92210 14 92217
rect -8 92209 17 92210
rect 25 92209 27 92218
rect -12 92202 38 92209
rect -12 92201 34 92202
rect -12 92197 8 92201
rect 0 92185 8 92197
rect 14 92185 34 92201
rect 0 92184 34 92185
rect 0 92177 38 92184
rect 14 92176 17 92177
rect 25 92168 27 92177
rect 42 92148 45 92238
rect 69 92223 80 92255
rect 107 92223 143 92251
rect 144 92223 148 92443
rect 332 92375 336 92443
rect 380 92413 462 92445
rect 463 92413 472 92447
rect 480 92413 497 92447
rect 378 92405 464 92413
rect 505 92405 507 92455
rect 514 92413 548 92447
rect 565 92413 582 92447
rect 607 92405 609 92455
rect 404 92389 438 92405
rect 400 92375 442 92376
rect 378 92369 404 92375
rect 442 92369 464 92375
rect 400 92368 404 92369
rect 174 92329 246 92337
rect 295 92334 300 92368
rect 324 92334 329 92368
rect 224 92299 226 92315
rect 196 92291 226 92299
rect 332 92297 336 92365
rect 367 92334 438 92368
rect 400 92327 404 92334
rect 454 92321 504 92323
rect 494 92317 548 92321
rect 494 92312 514 92317
rect 504 92297 506 92312
rect 196 92287 232 92291
rect 196 92257 204 92287
rect 216 92257 232 92287
rect 400 92289 404 92297
rect 107 92217 119 92223
rect 109 92189 119 92217
rect 129 92189 149 92223
rect 174 92219 181 92249
rect 224 92210 226 92257
rect 256 92249 328 92257
rect 332 92255 336 92285
rect 400 92255 408 92289
rect 434 92255 438 92289
rect 498 92287 506 92297
rect 514 92287 515 92307
rect 504 92271 506 92287
rect 525 92278 528 92312
rect 547 92287 548 92307
rect 557 92287 564 92297
rect 514 92271 530 92277
rect 532 92271 548 92277
rect 278 92219 305 92230
rect 42 92097 46 92131
rect 72 92097 76 92131
rect 38 92059 80 92060
rect 42 92018 76 92052
rect 79 92018 113 92052
rect 42 91939 46 91973
rect 72 91939 76 91973
rect -25 91902 25 91904
rect -8 91894 14 91901
rect -8 91893 17 91894
rect 25 91893 27 91902
rect -12 91886 38 91893
rect -12 91885 34 91886
rect -12 91881 8 91885
rect 0 91869 8 91881
rect 14 91869 34 91885
rect 0 91868 34 91869
rect 0 91861 38 91868
rect 14 91860 17 91861
rect 25 91852 27 91861
rect 42 91832 45 91922
rect 71 91891 80 91919
rect 69 91853 80 91891
rect 144 91881 148 92189
rect 196 92176 204 92210
rect 216 92176 232 92210
rect 244 92206 257 92210
rect 300 92206 308 92219
rect 332 92217 342 92255
rect 400 92247 404 92255
rect 336 92207 342 92217
rect 244 92182 291 92206
rect 244 92176 257 92182
rect 224 92129 226 92176
rect 278 92172 291 92182
rect 300 92182 329 92206
rect 332 92197 342 92207
rect 400 92207 409 92235
rect 562 92218 612 92220
rect 466 92209 497 92217
rect 565 92209 596 92217
rect 300 92172 321 92182
rect 300 92166 308 92172
rect 289 92156 308 92166
rect 196 92099 204 92129
rect 216 92099 232 92129
rect 196 92095 232 92099
rect 196 92087 226 92095
rect 300 92087 308 92156
rect 332 92163 351 92197
rect 361 92169 381 92197
rect 361 92163 375 92169
rect 400 92163 411 92207
rect 442 92202 500 92209
rect 466 92201 500 92202
rect 565 92201 599 92209
rect 497 92185 500 92201
rect 596 92185 599 92201
rect 466 92184 500 92185
rect 442 92177 500 92184
rect 565 92177 599 92185
rect 612 92168 614 92218
rect 332 92139 342 92163
rect 336 92127 342 92139
rect 224 92071 226 92087
rect 332 92059 342 92127
rect 400 92131 404 92139
rect 400 92097 408 92131
rect 434 92097 438 92131
rect 454 92115 504 92117
rect 504 92099 506 92115
rect 514 92109 530 92115
rect 532 92109 548 92115
rect 525 92099 548 92108
rect 400 92089 404 92097
rect 498 92089 506 92099
rect 504 92065 506 92089
rect 514 92079 515 92099
rect 525 92074 528 92099
rect 547 92079 548 92099
rect 557 92089 564 92099
rect 514 92065 548 92069
rect 151 92018 156 92052
rect 174 92049 246 92057
rect 256 92049 328 92057
rect 336 92051 342 92059
rect 400 92054 404 92059
rect 180 92021 185 92049
rect 174 92013 246 92021
rect 256 92013 328 92021
rect 332 92019 336 92049
rect 400 92020 438 92054
rect 224 91983 226 91999
rect 196 91975 226 91983
rect 196 91971 232 91975
rect 196 91941 204 91971
rect 216 91941 232 91971
rect 224 91894 226 91941
rect 300 91914 308 91983
rect 332 91981 342 92019
rect 400 92011 404 92020
rect 454 92005 504 92007
rect 494 92001 548 92005
rect 494 91996 514 92001
rect 504 91981 506 91996
rect 336 91969 342 91981
rect 289 91904 308 91914
rect 300 91898 308 91904
rect 332 91935 342 91969
rect 400 91973 404 91981
rect 400 91939 408 91973
rect 434 91939 438 91973
rect 498 91971 506 91981
rect 514 91971 515 91991
rect 504 91955 506 91971
rect 525 91962 528 91996
rect 547 91971 548 91991
rect 557 91971 564 91981
rect 514 91955 530 91961
rect 532 91955 548 91961
rect 332 91907 373 91935
rect 332 91901 351 91907
rect 107 91847 119 91881
rect 129 91847 149 91881
rect 196 91860 204 91894
rect 216 91860 232 91894
rect 244 91888 257 91894
rect 278 91888 291 91898
rect 244 91864 291 91888
rect 300 91888 321 91898
rect 336 91891 351 91901
rect 300 91864 329 91888
rect 332 91873 351 91891
rect 361 91901 375 91907
rect 400 91901 411 91939
rect 562 91902 612 91904
rect 361 91873 381 91901
rect 400 91873 409 91901
rect 466 91893 497 91901
rect 565 91893 596 91901
rect 442 91886 500 91893
rect 466 91885 500 91886
rect 565 91885 599 91893
rect 244 91860 257 91864
rect 42 91781 46 91815
rect 72 91781 76 91815
rect 42 91734 76 91738
rect 42 91719 46 91734
rect 72 91719 76 91734
rect 38 91701 80 91719
rect 16 91695 102 91701
rect 144 91695 148 91847
rect 174 91823 181 91851
rect 224 91813 226 91860
rect 300 91851 308 91864
rect 278 91840 305 91851
rect 332 91823 342 91873
rect 400 91853 404 91873
rect 497 91869 500 91885
rect 596 91869 599 91885
rect 466 91868 500 91869
rect 442 91861 500 91868
rect 565 91861 599 91869
rect 612 91852 614 91902
rect 256 91813 328 91821
rect 336 91815 342 91823
rect 400 91815 404 91823
rect 196 91783 204 91813
rect 216 91783 232 91813
rect 196 91779 232 91783
rect 196 91771 226 91779
rect 224 91755 226 91771
rect 332 91743 336 91811
rect 400 91781 408 91815
rect 434 91781 438 91815
rect 454 91799 504 91801
rect 504 91783 506 91799
rect 514 91793 530 91799
rect 532 91793 548 91799
rect 525 91783 548 91792
rect 400 91773 404 91781
rect 498 91773 506 91783
rect 504 91749 506 91773
rect 514 91763 515 91783
rect 525 91758 528 91783
rect 547 91763 548 91783
rect 557 91773 564 91783
rect 514 91749 548 91753
rect 400 91743 442 91744
rect 174 91733 246 91741
rect 400 91736 404 91743
rect 295 91702 300 91736
rect 324 91702 329 91736
rect 367 91719 438 91736
rect 367 91702 442 91719
rect 400 91701 442 91702
rect 378 91695 464 91701
rect 38 91679 80 91695
rect 400 91679 442 91695
rect -25 91665 25 91667
rect 42 91665 76 91679
rect 404 91665 438 91679
rect 455 91665 505 91667
rect 557 91665 607 91667
rect 16 91657 102 91665
rect 378 91657 464 91665
rect 8 91623 17 91657
rect 18 91655 51 91657
rect 80 91655 100 91657
rect 18 91623 100 91655
rect 380 91655 404 91657
rect 429 91655 438 91657
rect 442 91655 462 91657
rect 16 91615 102 91623
rect 42 91599 76 91615
rect 16 91579 38 91585
rect 42 91576 76 91580
rect 80 91579 102 91585
rect 42 91546 46 91576
rect 72 91546 76 91576
rect 42 91465 46 91499
rect 72 91465 76 91499
rect -25 91428 25 91430
rect -8 91420 14 91427
rect -8 91419 17 91420
rect 25 91419 27 91428
rect -12 91412 38 91419
rect -12 91411 34 91412
rect -12 91407 8 91411
rect 0 91395 8 91407
rect 14 91395 34 91411
rect 0 91394 34 91395
rect 0 91387 38 91394
rect 14 91386 17 91387
rect 25 91378 27 91387
rect 42 91358 45 91448
rect 69 91433 80 91465
rect 107 91433 143 91461
rect 144 91433 148 91653
rect 332 91585 336 91653
rect 380 91623 462 91655
rect 463 91623 472 91657
rect 480 91623 497 91657
rect 378 91615 464 91623
rect 505 91615 507 91665
rect 514 91623 548 91657
rect 565 91623 582 91657
rect 607 91615 609 91665
rect 404 91599 438 91615
rect 400 91585 442 91586
rect 378 91579 404 91585
rect 442 91579 464 91585
rect 400 91578 404 91579
rect 174 91539 246 91547
rect 295 91544 300 91578
rect 324 91544 329 91578
rect 224 91509 226 91525
rect 196 91501 226 91509
rect 332 91507 336 91575
rect 367 91544 438 91578
rect 400 91537 404 91544
rect 454 91531 504 91533
rect 494 91527 548 91531
rect 494 91522 514 91527
rect 504 91507 506 91522
rect 196 91497 232 91501
rect 196 91467 204 91497
rect 216 91467 232 91497
rect 400 91499 404 91507
rect 107 91427 119 91433
rect 109 91399 119 91427
rect 129 91399 149 91433
rect 174 91429 181 91459
rect 224 91420 226 91467
rect 256 91459 328 91467
rect 332 91465 336 91495
rect 400 91465 408 91499
rect 434 91465 438 91499
rect 498 91497 506 91507
rect 514 91497 515 91517
rect 504 91481 506 91497
rect 525 91488 528 91522
rect 547 91497 548 91517
rect 557 91497 564 91507
rect 514 91481 530 91487
rect 532 91481 548 91487
rect 278 91429 305 91440
rect 42 91307 46 91341
rect 72 91307 76 91341
rect 38 91269 80 91270
rect 42 91228 76 91262
rect 79 91228 113 91262
rect 42 91149 46 91183
rect 72 91149 76 91183
rect -25 91112 25 91114
rect -8 91104 14 91111
rect -8 91103 17 91104
rect 25 91103 27 91112
rect -12 91096 38 91103
rect -12 91095 34 91096
rect -12 91091 8 91095
rect 0 91079 8 91091
rect 14 91079 34 91095
rect 0 91078 34 91079
rect 0 91071 38 91078
rect 14 91070 17 91071
rect 25 91062 27 91071
rect 42 91042 45 91132
rect 71 91101 80 91129
rect 69 91063 80 91101
rect 144 91091 148 91399
rect 196 91386 204 91420
rect 216 91386 232 91420
rect 244 91416 257 91420
rect 300 91416 308 91429
rect 332 91427 342 91465
rect 400 91457 404 91465
rect 336 91417 342 91427
rect 244 91392 291 91416
rect 244 91386 257 91392
rect 224 91339 226 91386
rect 278 91382 291 91392
rect 300 91392 329 91416
rect 332 91407 342 91417
rect 400 91417 409 91445
rect 562 91428 612 91430
rect 466 91419 497 91427
rect 565 91419 596 91427
rect 300 91382 321 91392
rect 300 91376 308 91382
rect 289 91366 308 91376
rect 196 91309 204 91339
rect 216 91309 232 91339
rect 196 91305 232 91309
rect 196 91297 226 91305
rect 300 91297 308 91366
rect 332 91373 351 91407
rect 361 91379 381 91407
rect 361 91373 375 91379
rect 400 91373 411 91417
rect 442 91412 500 91419
rect 466 91411 500 91412
rect 565 91411 599 91419
rect 497 91395 500 91411
rect 596 91395 599 91411
rect 466 91394 500 91395
rect 442 91387 500 91394
rect 565 91387 599 91395
rect 612 91378 614 91428
rect 332 91349 342 91373
rect 336 91337 342 91349
rect 224 91281 226 91297
rect 332 91269 342 91337
rect 400 91341 404 91349
rect 400 91307 408 91341
rect 434 91307 438 91341
rect 454 91325 504 91327
rect 504 91309 506 91325
rect 514 91319 530 91325
rect 532 91319 548 91325
rect 525 91309 548 91318
rect 400 91299 404 91307
rect 498 91299 506 91309
rect 504 91275 506 91299
rect 514 91289 515 91309
rect 525 91284 528 91309
rect 547 91289 548 91309
rect 557 91299 564 91309
rect 514 91275 548 91279
rect 151 91228 156 91262
rect 174 91259 246 91267
rect 256 91259 328 91267
rect 336 91261 342 91269
rect 400 91264 404 91269
rect 180 91231 185 91259
rect 174 91223 246 91231
rect 256 91223 328 91231
rect 332 91229 336 91259
rect 400 91230 438 91264
rect 224 91193 226 91209
rect 196 91185 226 91193
rect 196 91181 232 91185
rect 196 91151 204 91181
rect 216 91151 232 91181
rect 224 91104 226 91151
rect 300 91124 308 91193
rect 332 91191 342 91229
rect 400 91221 404 91230
rect 454 91215 504 91217
rect 494 91211 548 91215
rect 494 91206 514 91211
rect 504 91191 506 91206
rect 336 91179 342 91191
rect 289 91114 308 91124
rect 300 91108 308 91114
rect 332 91145 342 91179
rect 400 91183 404 91191
rect 400 91149 408 91183
rect 434 91149 438 91183
rect 498 91181 506 91191
rect 514 91181 515 91201
rect 504 91165 506 91181
rect 525 91172 528 91206
rect 547 91181 548 91201
rect 557 91181 564 91191
rect 514 91165 530 91171
rect 532 91165 548 91171
rect 332 91117 373 91145
rect 332 91111 351 91117
rect 107 91057 119 91091
rect 129 91057 149 91091
rect 196 91070 204 91104
rect 216 91070 232 91104
rect 244 91098 257 91104
rect 278 91098 291 91108
rect 244 91074 291 91098
rect 300 91098 321 91108
rect 336 91101 351 91111
rect 300 91074 329 91098
rect 332 91083 351 91101
rect 361 91111 375 91117
rect 400 91111 411 91149
rect 562 91112 612 91114
rect 361 91083 381 91111
rect 400 91083 409 91111
rect 466 91103 497 91111
rect 565 91103 596 91111
rect 442 91096 500 91103
rect 466 91095 500 91096
rect 565 91095 599 91103
rect 244 91070 257 91074
rect 42 90991 46 91025
rect 72 90991 76 91025
rect 42 90944 76 90948
rect 42 90929 46 90944
rect 72 90929 76 90944
rect 38 90911 80 90929
rect 16 90905 102 90911
rect 144 90905 148 91057
rect 174 91033 181 91061
rect 224 91023 226 91070
rect 300 91061 308 91074
rect 278 91050 305 91061
rect 332 91033 342 91083
rect 400 91063 404 91083
rect 497 91079 500 91095
rect 596 91079 599 91095
rect 466 91078 500 91079
rect 442 91071 500 91078
rect 565 91071 599 91079
rect 612 91062 614 91112
rect 256 91023 328 91031
rect 336 91025 342 91033
rect 400 91025 404 91033
rect 196 90993 204 91023
rect 216 90993 232 91023
rect 196 90989 232 90993
rect 196 90981 226 90989
rect 224 90965 226 90981
rect 332 90953 336 91021
rect 400 90991 408 91025
rect 434 90991 438 91025
rect 454 91009 504 91011
rect 504 90993 506 91009
rect 514 91003 530 91009
rect 532 91003 548 91009
rect 525 90993 548 91002
rect 400 90983 404 90991
rect 498 90983 506 90993
rect 504 90959 506 90983
rect 514 90973 515 90993
rect 525 90968 528 90993
rect 547 90973 548 90993
rect 557 90983 564 90993
rect 514 90959 548 90963
rect 400 90953 442 90954
rect 174 90943 246 90951
rect 400 90946 404 90953
rect 295 90912 300 90946
rect 324 90912 329 90946
rect 367 90929 438 90946
rect 367 90912 442 90929
rect 400 90911 442 90912
rect 378 90905 464 90911
rect 38 90889 80 90905
rect 400 90889 442 90905
rect -25 90875 25 90877
rect 42 90875 76 90889
rect 404 90875 438 90889
rect 455 90875 505 90877
rect 557 90875 607 90877
rect 16 90867 102 90875
rect 378 90867 464 90875
rect 8 90833 17 90867
rect 18 90865 51 90867
rect 80 90865 100 90867
rect 18 90833 100 90865
rect 380 90865 404 90867
rect 429 90865 438 90867
rect 442 90865 462 90867
rect 16 90825 102 90833
rect 42 90809 76 90825
rect 16 90789 38 90795
rect 42 90786 76 90790
rect 80 90789 102 90795
rect 42 90756 46 90786
rect 72 90756 76 90786
rect 42 90675 46 90709
rect 72 90675 76 90709
rect -25 90638 25 90640
rect -8 90630 14 90637
rect -8 90629 17 90630
rect 25 90629 27 90638
rect -12 90622 38 90629
rect -12 90621 34 90622
rect -12 90617 8 90621
rect 0 90605 8 90617
rect 14 90605 34 90621
rect 0 90604 34 90605
rect 0 90597 38 90604
rect 14 90596 17 90597
rect 25 90588 27 90597
rect 42 90568 45 90658
rect 69 90643 80 90675
rect 107 90643 143 90671
rect 144 90643 148 90863
rect 332 90795 336 90863
rect 380 90833 462 90865
rect 463 90833 472 90867
rect 480 90833 497 90867
rect 378 90825 464 90833
rect 505 90825 507 90875
rect 514 90833 548 90867
rect 565 90833 582 90867
rect 607 90825 609 90875
rect 404 90809 438 90825
rect 400 90795 442 90796
rect 378 90789 404 90795
rect 442 90789 464 90795
rect 400 90788 404 90789
rect 174 90749 246 90757
rect 295 90754 300 90788
rect 324 90754 329 90788
rect 224 90719 226 90735
rect 196 90711 226 90719
rect 332 90717 336 90785
rect 367 90754 438 90788
rect 400 90747 404 90754
rect 454 90741 504 90743
rect 494 90737 548 90741
rect 494 90732 514 90737
rect 504 90717 506 90732
rect 196 90707 232 90711
rect 196 90677 204 90707
rect 216 90677 232 90707
rect 400 90709 404 90717
rect 107 90637 119 90643
rect 109 90609 119 90637
rect 129 90609 149 90643
rect 174 90639 181 90669
rect 224 90630 226 90677
rect 256 90669 328 90677
rect 332 90675 336 90705
rect 400 90675 408 90709
rect 434 90675 438 90709
rect 498 90707 506 90717
rect 514 90707 515 90727
rect 504 90691 506 90707
rect 525 90698 528 90732
rect 547 90707 548 90727
rect 557 90707 564 90717
rect 514 90691 530 90697
rect 532 90691 548 90697
rect 278 90639 305 90650
rect 42 90517 46 90551
rect 72 90517 76 90551
rect 38 90479 80 90480
rect 42 90438 76 90472
rect 79 90438 113 90472
rect 42 90359 46 90393
rect 72 90359 76 90393
rect -25 90322 25 90324
rect -8 90314 14 90321
rect -8 90313 17 90314
rect 25 90313 27 90322
rect -12 90306 38 90313
rect -12 90305 34 90306
rect -12 90301 8 90305
rect 0 90289 8 90301
rect 14 90289 34 90305
rect 0 90288 34 90289
rect 0 90281 38 90288
rect 14 90280 17 90281
rect 25 90272 27 90281
rect 42 90252 45 90342
rect 71 90311 80 90339
rect 69 90273 80 90311
rect 144 90301 148 90609
rect 196 90596 204 90630
rect 216 90596 232 90630
rect 244 90626 257 90630
rect 300 90626 308 90639
rect 332 90637 342 90675
rect 400 90667 404 90675
rect 336 90627 342 90637
rect 244 90602 291 90626
rect 244 90596 257 90602
rect 224 90549 226 90596
rect 278 90592 291 90602
rect 300 90602 329 90626
rect 332 90617 342 90627
rect 400 90627 409 90655
rect 562 90638 612 90640
rect 466 90629 497 90637
rect 565 90629 596 90637
rect 300 90592 321 90602
rect 300 90586 308 90592
rect 289 90576 308 90586
rect 196 90519 204 90549
rect 216 90519 232 90549
rect 196 90515 232 90519
rect 196 90507 226 90515
rect 300 90507 308 90576
rect 332 90583 351 90617
rect 361 90589 381 90617
rect 361 90583 375 90589
rect 400 90583 411 90627
rect 442 90622 500 90629
rect 466 90621 500 90622
rect 565 90621 599 90629
rect 497 90605 500 90621
rect 596 90605 599 90621
rect 466 90604 500 90605
rect 442 90597 500 90604
rect 565 90597 599 90605
rect 612 90588 614 90638
rect 332 90559 342 90583
rect 336 90547 342 90559
rect 224 90491 226 90507
rect 332 90479 342 90547
rect 400 90551 404 90559
rect 400 90517 408 90551
rect 434 90517 438 90551
rect 454 90535 504 90537
rect 504 90519 506 90535
rect 514 90529 530 90535
rect 532 90529 548 90535
rect 525 90519 548 90528
rect 400 90509 404 90517
rect 498 90509 506 90519
rect 504 90485 506 90509
rect 514 90499 515 90519
rect 525 90494 528 90519
rect 547 90499 548 90519
rect 557 90509 564 90519
rect 514 90485 548 90489
rect 151 90438 156 90472
rect 174 90469 246 90477
rect 256 90469 328 90477
rect 336 90471 342 90479
rect 400 90474 404 90479
rect 180 90441 185 90469
rect 174 90433 246 90441
rect 256 90433 328 90441
rect 332 90439 336 90469
rect 400 90440 438 90474
rect 224 90403 226 90419
rect 196 90395 226 90403
rect 196 90391 232 90395
rect 196 90361 204 90391
rect 216 90361 232 90391
rect 224 90314 226 90361
rect 300 90334 308 90403
rect 332 90401 342 90439
rect 400 90431 404 90440
rect 454 90425 504 90427
rect 494 90421 548 90425
rect 494 90416 514 90421
rect 504 90401 506 90416
rect 336 90389 342 90401
rect 289 90324 308 90334
rect 300 90318 308 90324
rect 332 90355 342 90389
rect 400 90393 404 90401
rect 400 90359 408 90393
rect 434 90359 438 90393
rect 498 90391 506 90401
rect 514 90391 515 90411
rect 504 90375 506 90391
rect 525 90382 528 90416
rect 547 90391 548 90411
rect 557 90391 564 90401
rect 514 90375 530 90381
rect 532 90375 548 90381
rect 332 90327 373 90355
rect 332 90321 351 90327
rect 107 90267 119 90301
rect 129 90267 149 90301
rect 196 90280 204 90314
rect 216 90280 232 90314
rect 244 90308 257 90314
rect 278 90308 291 90318
rect 244 90284 291 90308
rect 300 90308 321 90318
rect 336 90311 351 90321
rect 300 90284 329 90308
rect 332 90293 351 90311
rect 361 90321 375 90327
rect 400 90321 411 90359
rect 562 90322 612 90324
rect 361 90293 381 90321
rect 400 90293 409 90321
rect 466 90313 497 90321
rect 565 90313 596 90321
rect 442 90306 500 90313
rect 466 90305 500 90306
rect 565 90305 599 90313
rect 244 90280 257 90284
rect 42 90201 46 90235
rect 72 90201 76 90235
rect 42 90154 76 90158
rect 42 90139 46 90154
rect 72 90139 76 90154
rect 38 90121 80 90139
rect 16 90115 102 90121
rect 144 90115 148 90267
rect 174 90243 181 90271
rect 224 90233 226 90280
rect 300 90271 308 90284
rect 278 90260 305 90271
rect 332 90243 342 90293
rect 400 90273 404 90293
rect 497 90289 500 90305
rect 596 90289 599 90305
rect 466 90288 500 90289
rect 442 90281 500 90288
rect 565 90281 599 90289
rect 612 90272 614 90322
rect 256 90233 328 90241
rect 336 90235 342 90243
rect 400 90235 404 90243
rect 196 90203 204 90233
rect 216 90203 232 90233
rect 196 90199 232 90203
rect 196 90191 226 90199
rect 224 90175 226 90191
rect 332 90163 336 90231
rect 400 90201 408 90235
rect 434 90201 438 90235
rect 454 90219 504 90221
rect 504 90203 506 90219
rect 514 90213 530 90219
rect 532 90213 548 90219
rect 525 90203 548 90212
rect 400 90193 404 90201
rect 498 90193 506 90203
rect 504 90169 506 90193
rect 514 90183 515 90203
rect 525 90178 528 90203
rect 547 90183 548 90203
rect 557 90193 564 90203
rect 514 90169 548 90173
rect 400 90163 442 90164
rect 174 90153 246 90161
rect 400 90156 404 90163
rect 295 90122 300 90156
rect 324 90122 329 90156
rect 367 90139 438 90156
rect 367 90122 442 90139
rect 400 90121 442 90122
rect 378 90115 464 90121
rect 38 90099 80 90115
rect 400 90099 442 90115
rect -25 90085 25 90087
rect 42 90085 76 90099
rect 404 90085 438 90099
rect 455 90085 505 90087
rect 557 90085 607 90087
rect 16 90077 102 90085
rect 378 90077 464 90085
rect 8 90043 17 90077
rect 18 90075 51 90077
rect 80 90075 100 90077
rect 18 90043 100 90075
rect 380 90075 404 90077
rect 429 90075 438 90077
rect 442 90075 462 90077
rect 16 90035 102 90043
rect 42 90019 76 90035
rect 16 89999 38 90005
rect 42 89996 76 90000
rect 80 89999 102 90005
rect 42 89966 46 89996
rect 72 89966 76 89996
rect 42 89885 46 89919
rect 72 89885 76 89919
rect -25 89848 25 89850
rect -8 89840 14 89847
rect -8 89839 17 89840
rect 25 89839 27 89848
rect -12 89832 38 89839
rect -12 89831 34 89832
rect -12 89827 8 89831
rect 0 89815 8 89827
rect 14 89815 34 89831
rect 0 89814 34 89815
rect 0 89807 38 89814
rect 14 89806 17 89807
rect 25 89798 27 89807
rect 42 89778 45 89868
rect 69 89853 80 89885
rect 107 89853 143 89881
rect 144 89853 148 90073
rect 332 90005 336 90073
rect 380 90043 462 90075
rect 463 90043 472 90077
rect 480 90043 497 90077
rect 378 90035 464 90043
rect 505 90035 507 90085
rect 514 90043 548 90077
rect 565 90043 582 90077
rect 607 90035 609 90085
rect 404 90019 438 90035
rect 400 90005 442 90006
rect 378 89999 404 90005
rect 442 89999 464 90005
rect 400 89998 404 89999
rect 174 89959 246 89967
rect 295 89964 300 89998
rect 324 89964 329 89998
rect 224 89929 226 89945
rect 196 89921 226 89929
rect 332 89927 336 89995
rect 367 89964 438 89998
rect 400 89957 404 89964
rect 454 89951 504 89953
rect 494 89947 548 89951
rect 494 89942 514 89947
rect 504 89927 506 89942
rect 196 89917 232 89921
rect 196 89887 204 89917
rect 216 89887 232 89917
rect 400 89919 404 89927
rect 107 89847 119 89853
rect 109 89819 119 89847
rect 129 89819 149 89853
rect 174 89849 181 89879
rect 224 89840 226 89887
rect 256 89879 328 89887
rect 332 89885 336 89915
rect 400 89885 408 89919
rect 434 89885 438 89919
rect 498 89917 506 89927
rect 514 89917 515 89937
rect 504 89901 506 89917
rect 525 89908 528 89942
rect 547 89917 548 89937
rect 557 89917 564 89927
rect 514 89901 530 89907
rect 532 89901 548 89907
rect 278 89849 305 89860
rect 42 89727 46 89761
rect 72 89727 76 89761
rect 38 89689 80 89690
rect 42 89648 76 89682
rect 79 89648 113 89682
rect 42 89569 46 89603
rect 72 89569 76 89603
rect -25 89532 25 89534
rect -8 89524 14 89531
rect -8 89523 17 89524
rect 25 89523 27 89532
rect -12 89516 38 89523
rect -12 89515 34 89516
rect -12 89511 8 89515
rect 0 89499 8 89511
rect 14 89499 34 89515
rect 0 89498 34 89499
rect 0 89491 38 89498
rect 14 89490 17 89491
rect 25 89482 27 89491
rect 42 89462 45 89552
rect 71 89521 80 89549
rect 69 89483 80 89521
rect 144 89511 148 89819
rect 196 89806 204 89840
rect 216 89806 232 89840
rect 244 89836 257 89840
rect 300 89836 308 89849
rect 332 89847 342 89885
rect 400 89877 404 89885
rect 336 89837 342 89847
rect 244 89812 291 89836
rect 244 89806 257 89812
rect 224 89759 226 89806
rect 278 89802 291 89812
rect 300 89812 329 89836
rect 332 89827 342 89837
rect 400 89837 409 89865
rect 562 89848 612 89850
rect 466 89839 497 89847
rect 565 89839 596 89847
rect 300 89802 321 89812
rect 300 89796 308 89802
rect 289 89786 308 89796
rect 196 89729 204 89759
rect 216 89729 232 89759
rect 196 89725 232 89729
rect 196 89717 226 89725
rect 300 89717 308 89786
rect 332 89793 351 89827
rect 361 89799 381 89827
rect 361 89793 375 89799
rect 400 89793 411 89837
rect 442 89832 500 89839
rect 466 89831 500 89832
rect 565 89831 599 89839
rect 497 89815 500 89831
rect 596 89815 599 89831
rect 466 89814 500 89815
rect 442 89807 500 89814
rect 565 89807 599 89815
rect 612 89798 614 89848
rect 332 89769 342 89793
rect 336 89757 342 89769
rect 224 89701 226 89717
rect 332 89689 342 89757
rect 400 89761 404 89769
rect 400 89727 408 89761
rect 434 89727 438 89761
rect 454 89745 504 89747
rect 504 89729 506 89745
rect 514 89739 530 89745
rect 532 89739 548 89745
rect 525 89729 548 89738
rect 400 89719 404 89727
rect 498 89719 506 89729
rect 504 89695 506 89719
rect 514 89709 515 89729
rect 525 89704 528 89729
rect 547 89709 548 89729
rect 557 89719 564 89729
rect 514 89695 548 89699
rect 151 89648 156 89682
rect 174 89679 246 89687
rect 256 89679 328 89687
rect 336 89681 342 89689
rect 400 89684 404 89689
rect 180 89651 185 89679
rect 174 89643 246 89651
rect 256 89643 328 89651
rect 332 89649 336 89679
rect 400 89650 438 89684
rect 224 89613 226 89629
rect 196 89605 226 89613
rect 196 89601 232 89605
rect 196 89571 204 89601
rect 216 89571 232 89601
rect 224 89524 226 89571
rect 300 89544 308 89613
rect 332 89611 342 89649
rect 400 89641 404 89650
rect 454 89635 504 89637
rect 494 89631 548 89635
rect 494 89626 514 89631
rect 504 89611 506 89626
rect 336 89599 342 89611
rect 289 89534 308 89544
rect 300 89528 308 89534
rect 332 89565 342 89599
rect 400 89603 404 89611
rect 400 89569 408 89603
rect 434 89569 438 89603
rect 498 89601 506 89611
rect 514 89601 515 89621
rect 504 89585 506 89601
rect 525 89592 528 89626
rect 547 89601 548 89621
rect 557 89601 564 89611
rect 514 89585 530 89591
rect 532 89585 548 89591
rect 332 89537 373 89565
rect 332 89531 351 89537
rect 107 89477 119 89511
rect 129 89477 149 89511
rect 196 89490 204 89524
rect 216 89490 232 89524
rect 244 89518 257 89524
rect 278 89518 291 89528
rect 244 89494 291 89518
rect 300 89518 321 89528
rect 336 89521 351 89531
rect 300 89494 329 89518
rect 332 89503 351 89521
rect 361 89531 375 89537
rect 400 89531 411 89569
rect 562 89532 612 89534
rect 361 89503 381 89531
rect 400 89503 409 89531
rect 466 89523 497 89531
rect 565 89523 596 89531
rect 442 89516 500 89523
rect 466 89515 500 89516
rect 565 89515 599 89523
rect 244 89490 257 89494
rect 42 89411 46 89445
rect 72 89411 76 89445
rect 42 89364 76 89368
rect 42 89349 46 89364
rect 72 89349 76 89364
rect 38 89331 80 89349
rect 16 89325 102 89331
rect 144 89325 148 89477
rect 174 89453 181 89481
rect 224 89443 226 89490
rect 300 89481 308 89494
rect 278 89470 305 89481
rect 332 89453 342 89503
rect 400 89483 404 89503
rect 497 89499 500 89515
rect 596 89499 599 89515
rect 466 89498 500 89499
rect 442 89491 500 89498
rect 565 89491 599 89499
rect 612 89482 614 89532
rect 256 89443 328 89451
rect 336 89445 342 89453
rect 400 89445 404 89453
rect 196 89413 204 89443
rect 216 89413 232 89443
rect 196 89409 232 89413
rect 196 89401 226 89409
rect 224 89385 226 89401
rect 332 89373 336 89441
rect 400 89411 408 89445
rect 434 89411 438 89445
rect 454 89429 504 89431
rect 504 89413 506 89429
rect 514 89423 530 89429
rect 532 89423 548 89429
rect 525 89413 548 89422
rect 400 89403 404 89411
rect 498 89403 506 89413
rect 504 89379 506 89403
rect 514 89393 515 89413
rect 525 89388 528 89413
rect 547 89393 548 89413
rect 557 89403 564 89413
rect 514 89379 548 89383
rect 400 89373 442 89374
rect 174 89363 246 89371
rect 400 89366 404 89373
rect 295 89332 300 89366
rect 324 89332 329 89366
rect 367 89349 438 89366
rect 367 89332 442 89349
rect 400 89331 442 89332
rect 378 89325 464 89331
rect 38 89309 80 89325
rect 400 89309 442 89325
rect -25 89295 25 89297
rect 42 89295 76 89309
rect 404 89295 438 89309
rect 455 89295 505 89297
rect 557 89295 607 89297
rect 16 89287 102 89295
rect 378 89287 464 89295
rect 8 89253 17 89287
rect 18 89285 51 89287
rect 80 89285 100 89287
rect 18 89253 100 89285
rect 380 89285 404 89287
rect 429 89285 438 89287
rect 442 89285 462 89287
rect 16 89245 102 89253
rect 42 89229 76 89245
rect 16 89209 38 89215
rect 42 89206 76 89210
rect 80 89209 102 89215
rect 42 89176 46 89206
rect 72 89176 76 89206
rect 42 89095 46 89129
rect 72 89095 76 89129
rect -25 89058 25 89060
rect -8 89050 14 89057
rect -8 89049 17 89050
rect 25 89049 27 89058
rect -12 89042 38 89049
rect -12 89041 34 89042
rect -12 89037 8 89041
rect 0 89025 8 89037
rect 14 89025 34 89041
rect 0 89024 34 89025
rect 0 89017 38 89024
rect 14 89016 17 89017
rect 25 89008 27 89017
rect 42 88988 45 89078
rect 69 89063 80 89095
rect 107 89063 143 89091
rect 144 89063 148 89283
rect 332 89215 336 89283
rect 380 89253 462 89285
rect 463 89253 472 89287
rect 480 89253 497 89287
rect 378 89245 464 89253
rect 505 89245 507 89295
rect 514 89253 548 89287
rect 565 89253 582 89287
rect 607 89245 609 89295
rect 404 89229 438 89245
rect 400 89215 442 89216
rect 378 89209 404 89215
rect 442 89209 464 89215
rect 400 89208 404 89209
rect 174 89169 246 89177
rect 295 89174 300 89208
rect 324 89174 329 89208
rect 224 89139 226 89155
rect 196 89131 226 89139
rect 332 89137 336 89205
rect 367 89174 438 89208
rect 400 89167 404 89174
rect 454 89161 504 89163
rect 494 89157 548 89161
rect 494 89152 514 89157
rect 504 89137 506 89152
rect 196 89127 232 89131
rect 196 89097 204 89127
rect 216 89097 232 89127
rect 400 89129 404 89137
rect 107 89057 119 89063
rect 109 89029 119 89057
rect 129 89029 149 89063
rect 174 89059 181 89089
rect 224 89050 226 89097
rect 256 89089 328 89097
rect 332 89095 336 89125
rect 400 89095 408 89129
rect 434 89095 438 89129
rect 498 89127 506 89137
rect 514 89127 515 89147
rect 504 89111 506 89127
rect 525 89118 528 89152
rect 547 89127 548 89147
rect 557 89127 564 89137
rect 514 89111 530 89117
rect 532 89111 548 89117
rect 278 89059 305 89070
rect 42 88937 46 88971
rect 72 88937 76 88971
rect 38 88899 80 88900
rect 42 88858 76 88892
rect 79 88858 113 88892
rect 42 88779 46 88813
rect 72 88779 76 88813
rect -25 88742 25 88744
rect -8 88734 14 88741
rect -8 88733 17 88734
rect 25 88733 27 88742
rect -12 88726 38 88733
rect -12 88725 34 88726
rect -12 88721 8 88725
rect 0 88709 8 88721
rect 14 88709 34 88725
rect 0 88708 34 88709
rect 0 88701 38 88708
rect 14 88700 17 88701
rect 25 88692 27 88701
rect 42 88672 45 88762
rect 71 88731 80 88759
rect 69 88693 80 88731
rect 144 88721 148 89029
rect 196 89016 204 89050
rect 216 89016 232 89050
rect 244 89046 257 89050
rect 300 89046 308 89059
rect 332 89057 342 89095
rect 400 89087 404 89095
rect 336 89047 342 89057
rect 244 89022 291 89046
rect 244 89016 257 89022
rect 224 88969 226 89016
rect 278 89012 291 89022
rect 300 89022 329 89046
rect 332 89037 342 89047
rect 400 89047 409 89075
rect 562 89058 612 89060
rect 466 89049 497 89057
rect 565 89049 596 89057
rect 300 89012 321 89022
rect 300 89006 308 89012
rect 289 88996 308 89006
rect 196 88939 204 88969
rect 216 88939 232 88969
rect 196 88935 232 88939
rect 196 88927 226 88935
rect 300 88927 308 88996
rect 332 89003 351 89037
rect 361 89009 381 89037
rect 361 89003 375 89009
rect 400 89003 411 89047
rect 442 89042 500 89049
rect 466 89041 500 89042
rect 565 89041 599 89049
rect 497 89025 500 89041
rect 596 89025 599 89041
rect 466 89024 500 89025
rect 442 89017 500 89024
rect 565 89017 599 89025
rect 612 89008 614 89058
rect 332 88979 342 89003
rect 336 88967 342 88979
rect 224 88911 226 88927
rect 332 88899 342 88967
rect 400 88971 404 88979
rect 400 88937 408 88971
rect 434 88937 438 88971
rect 454 88955 504 88957
rect 504 88939 506 88955
rect 514 88949 530 88955
rect 532 88949 548 88955
rect 525 88939 548 88948
rect 400 88929 404 88937
rect 498 88929 506 88939
rect 504 88905 506 88929
rect 514 88919 515 88939
rect 525 88914 528 88939
rect 547 88919 548 88939
rect 557 88929 564 88939
rect 514 88905 548 88909
rect 151 88858 156 88892
rect 174 88889 246 88897
rect 256 88889 328 88897
rect 336 88891 342 88899
rect 400 88894 404 88899
rect 180 88861 185 88889
rect 174 88853 246 88861
rect 256 88853 328 88861
rect 332 88859 336 88889
rect 400 88860 438 88894
rect 224 88823 226 88839
rect 196 88815 226 88823
rect 196 88811 232 88815
rect 196 88781 204 88811
rect 216 88781 232 88811
rect 224 88734 226 88781
rect 300 88754 308 88823
rect 332 88821 342 88859
rect 400 88851 404 88860
rect 454 88845 504 88847
rect 494 88841 548 88845
rect 494 88836 514 88841
rect 504 88821 506 88836
rect 336 88809 342 88821
rect 289 88744 308 88754
rect 300 88738 308 88744
rect 332 88775 342 88809
rect 400 88813 404 88821
rect 400 88779 408 88813
rect 434 88779 438 88813
rect 498 88811 506 88821
rect 514 88811 515 88831
rect 504 88795 506 88811
rect 525 88802 528 88836
rect 547 88811 548 88831
rect 557 88811 564 88821
rect 514 88795 530 88801
rect 532 88795 548 88801
rect 332 88747 373 88775
rect 332 88741 351 88747
rect 107 88687 119 88721
rect 129 88687 149 88721
rect 196 88700 204 88734
rect 216 88700 232 88734
rect 244 88728 257 88734
rect 278 88728 291 88738
rect 244 88704 291 88728
rect 300 88728 321 88738
rect 336 88731 351 88741
rect 300 88704 329 88728
rect 332 88713 351 88731
rect 361 88741 375 88747
rect 400 88741 411 88779
rect 562 88742 612 88744
rect 361 88713 381 88741
rect 400 88713 409 88741
rect 466 88733 497 88741
rect 565 88733 596 88741
rect 442 88726 500 88733
rect 466 88725 500 88726
rect 565 88725 599 88733
rect 244 88700 257 88704
rect 42 88621 46 88655
rect 72 88621 76 88655
rect 42 88574 76 88578
rect 42 88559 46 88574
rect 72 88559 76 88574
rect 38 88541 80 88559
rect 16 88535 102 88541
rect 144 88535 148 88687
rect 174 88663 181 88691
rect 224 88653 226 88700
rect 300 88691 308 88704
rect 278 88680 305 88691
rect 332 88663 342 88713
rect 400 88693 404 88713
rect 497 88709 500 88725
rect 596 88709 599 88725
rect 466 88708 500 88709
rect 442 88701 500 88708
rect 565 88701 599 88709
rect 612 88692 614 88742
rect 256 88653 328 88661
rect 336 88655 342 88663
rect 400 88655 404 88663
rect 196 88623 204 88653
rect 216 88623 232 88653
rect 196 88619 232 88623
rect 196 88611 226 88619
rect 224 88595 226 88611
rect 332 88583 336 88651
rect 400 88621 408 88655
rect 434 88621 438 88655
rect 454 88639 504 88641
rect 504 88623 506 88639
rect 514 88633 530 88639
rect 532 88633 548 88639
rect 525 88623 548 88632
rect 400 88613 404 88621
rect 498 88613 506 88623
rect 504 88589 506 88613
rect 514 88603 515 88623
rect 525 88598 528 88623
rect 547 88603 548 88623
rect 557 88613 564 88623
rect 514 88589 548 88593
rect 400 88583 442 88584
rect 174 88573 246 88581
rect 400 88576 404 88583
rect 295 88542 300 88576
rect 324 88542 329 88576
rect 367 88559 438 88576
rect 367 88542 442 88559
rect 400 88541 442 88542
rect 378 88535 464 88541
rect 38 88519 80 88535
rect 400 88519 442 88535
rect -25 88505 25 88507
rect 42 88505 76 88519
rect 404 88505 438 88519
rect 455 88505 505 88507
rect 557 88505 607 88507
rect 16 88497 102 88505
rect 378 88497 464 88505
rect 8 88463 17 88497
rect 18 88495 51 88497
rect 80 88495 100 88497
rect 18 88463 100 88495
rect 380 88495 404 88497
rect 429 88495 438 88497
rect 442 88495 462 88497
rect 16 88455 102 88463
rect 42 88439 76 88455
rect 16 88419 38 88425
rect 42 88416 76 88420
rect 80 88419 102 88425
rect 42 88386 46 88416
rect 72 88386 76 88416
rect 42 88305 46 88339
rect 72 88305 76 88339
rect -25 88268 25 88270
rect -8 88260 14 88267
rect -8 88259 17 88260
rect 25 88259 27 88268
rect -12 88252 38 88259
rect -12 88251 34 88252
rect -12 88247 8 88251
rect 0 88235 8 88247
rect 14 88235 34 88251
rect 0 88234 34 88235
rect 0 88227 38 88234
rect 14 88226 17 88227
rect 25 88218 27 88227
rect 42 88198 45 88288
rect 69 88273 80 88305
rect 107 88273 143 88301
rect 144 88273 148 88493
rect 332 88425 336 88493
rect 380 88463 462 88495
rect 463 88463 472 88497
rect 480 88463 497 88497
rect 378 88455 464 88463
rect 505 88455 507 88505
rect 514 88463 548 88497
rect 565 88463 582 88497
rect 607 88455 609 88505
rect 404 88439 438 88455
rect 400 88425 442 88426
rect 378 88419 404 88425
rect 442 88419 464 88425
rect 400 88418 404 88419
rect 174 88379 246 88387
rect 295 88384 300 88418
rect 324 88384 329 88418
rect 224 88349 226 88365
rect 196 88341 226 88349
rect 332 88347 336 88415
rect 367 88384 438 88418
rect 400 88377 404 88384
rect 454 88371 504 88373
rect 494 88367 548 88371
rect 494 88362 514 88367
rect 504 88347 506 88362
rect 196 88337 232 88341
rect 196 88307 204 88337
rect 216 88307 232 88337
rect 400 88339 404 88347
rect 107 88267 119 88273
rect 109 88239 119 88267
rect 129 88239 149 88273
rect 174 88269 181 88299
rect 224 88260 226 88307
rect 256 88299 328 88307
rect 332 88305 336 88335
rect 400 88305 408 88339
rect 434 88305 438 88339
rect 498 88337 506 88347
rect 514 88337 515 88357
rect 504 88321 506 88337
rect 525 88328 528 88362
rect 547 88337 548 88357
rect 557 88337 564 88347
rect 514 88321 530 88327
rect 532 88321 548 88327
rect 278 88269 305 88280
rect 42 88147 46 88181
rect 72 88147 76 88181
rect 38 88109 80 88110
rect 42 88068 76 88102
rect 79 88068 113 88102
rect 42 87989 46 88023
rect 72 87989 76 88023
rect -25 87952 25 87954
rect -8 87944 14 87951
rect -8 87943 17 87944
rect 25 87943 27 87952
rect -12 87936 38 87943
rect -12 87935 34 87936
rect -12 87931 8 87935
rect 0 87919 8 87931
rect 14 87919 34 87935
rect 0 87918 34 87919
rect 0 87911 38 87918
rect 14 87910 17 87911
rect 25 87902 27 87911
rect 42 87882 45 87972
rect 71 87941 80 87969
rect 69 87903 80 87941
rect 144 87931 148 88239
rect 196 88226 204 88260
rect 216 88226 232 88260
rect 244 88256 257 88260
rect 300 88256 308 88269
rect 332 88267 342 88305
rect 400 88297 404 88305
rect 336 88257 342 88267
rect 244 88232 291 88256
rect 244 88226 257 88232
rect 224 88179 226 88226
rect 278 88222 291 88232
rect 300 88232 329 88256
rect 332 88247 342 88257
rect 400 88257 409 88285
rect 562 88268 612 88270
rect 466 88259 497 88267
rect 565 88259 596 88267
rect 300 88222 321 88232
rect 300 88216 308 88222
rect 289 88206 308 88216
rect 196 88149 204 88179
rect 216 88149 232 88179
rect 196 88145 232 88149
rect 196 88137 226 88145
rect 300 88137 308 88206
rect 332 88213 351 88247
rect 361 88219 381 88247
rect 361 88213 375 88219
rect 400 88213 411 88257
rect 442 88252 500 88259
rect 466 88251 500 88252
rect 565 88251 599 88259
rect 497 88235 500 88251
rect 596 88235 599 88251
rect 466 88234 500 88235
rect 442 88227 500 88234
rect 565 88227 599 88235
rect 612 88218 614 88268
rect 332 88189 342 88213
rect 336 88177 342 88189
rect 224 88121 226 88137
rect 332 88109 342 88177
rect 400 88181 404 88189
rect 400 88147 408 88181
rect 434 88147 438 88181
rect 454 88165 504 88167
rect 504 88149 506 88165
rect 514 88159 530 88165
rect 532 88159 548 88165
rect 525 88149 548 88158
rect 400 88139 404 88147
rect 498 88139 506 88149
rect 504 88115 506 88139
rect 514 88129 515 88149
rect 525 88124 528 88149
rect 547 88129 548 88149
rect 557 88139 564 88149
rect 514 88115 548 88119
rect 151 88068 156 88102
rect 174 88099 246 88107
rect 256 88099 328 88107
rect 336 88101 342 88109
rect 400 88104 404 88109
rect 180 88071 185 88099
rect 174 88063 246 88071
rect 256 88063 328 88071
rect 332 88069 336 88099
rect 400 88070 438 88104
rect 224 88033 226 88049
rect 196 88025 226 88033
rect 196 88021 232 88025
rect 196 87991 204 88021
rect 216 87991 232 88021
rect 224 87944 226 87991
rect 300 87964 308 88033
rect 332 88031 342 88069
rect 400 88061 404 88070
rect 454 88055 504 88057
rect 494 88051 548 88055
rect 494 88046 514 88051
rect 504 88031 506 88046
rect 336 88019 342 88031
rect 289 87954 308 87964
rect 300 87948 308 87954
rect 332 87985 342 88019
rect 400 88023 404 88031
rect 400 87989 408 88023
rect 434 87989 438 88023
rect 498 88021 506 88031
rect 514 88021 515 88041
rect 504 88005 506 88021
rect 525 88012 528 88046
rect 547 88021 548 88041
rect 557 88021 564 88031
rect 514 88005 530 88011
rect 532 88005 548 88011
rect 332 87957 373 87985
rect 332 87951 351 87957
rect 107 87897 119 87931
rect 129 87897 149 87931
rect 196 87910 204 87944
rect 216 87910 232 87944
rect 244 87938 257 87944
rect 278 87938 291 87948
rect 244 87914 291 87938
rect 300 87938 321 87948
rect 336 87941 351 87951
rect 300 87914 329 87938
rect 332 87923 351 87941
rect 361 87951 375 87957
rect 400 87951 411 87989
rect 562 87952 612 87954
rect 361 87923 381 87951
rect 400 87923 409 87951
rect 466 87943 497 87951
rect 565 87943 596 87951
rect 442 87936 500 87943
rect 466 87935 500 87936
rect 565 87935 599 87943
rect 244 87910 257 87914
rect 42 87831 46 87865
rect 72 87831 76 87865
rect 42 87784 76 87788
rect 42 87769 46 87784
rect 72 87769 76 87784
rect 38 87751 80 87769
rect 16 87745 102 87751
rect 144 87745 148 87897
rect 174 87873 181 87901
rect 224 87863 226 87910
rect 300 87901 308 87914
rect 278 87890 305 87901
rect 332 87873 342 87923
rect 400 87903 404 87923
rect 497 87919 500 87935
rect 596 87919 599 87935
rect 466 87918 500 87919
rect 442 87911 500 87918
rect 565 87911 599 87919
rect 612 87902 614 87952
rect 256 87863 328 87871
rect 336 87865 342 87873
rect 400 87865 404 87873
rect 196 87833 204 87863
rect 216 87833 232 87863
rect 196 87829 232 87833
rect 196 87821 226 87829
rect 224 87805 226 87821
rect 332 87793 336 87861
rect 400 87831 408 87865
rect 434 87831 438 87865
rect 454 87849 504 87851
rect 504 87833 506 87849
rect 514 87843 530 87849
rect 532 87843 548 87849
rect 525 87833 548 87842
rect 400 87823 404 87831
rect 498 87823 506 87833
rect 504 87799 506 87823
rect 514 87813 515 87833
rect 525 87808 528 87833
rect 547 87813 548 87833
rect 557 87823 564 87833
rect 514 87799 548 87803
rect 400 87793 442 87794
rect 174 87783 246 87791
rect 400 87786 404 87793
rect 295 87752 300 87786
rect 324 87752 329 87786
rect 367 87769 438 87786
rect 367 87752 442 87769
rect 400 87751 442 87752
rect 378 87745 464 87751
rect 38 87729 80 87745
rect 400 87729 442 87745
rect -25 87715 25 87717
rect 42 87715 76 87729
rect 404 87715 438 87729
rect 455 87715 505 87717
rect 557 87715 607 87717
rect 16 87707 102 87715
rect 378 87707 464 87715
rect 8 87673 17 87707
rect 18 87705 51 87707
rect 80 87705 100 87707
rect 18 87673 100 87705
rect 380 87705 404 87707
rect 429 87705 438 87707
rect 442 87705 462 87707
rect 16 87665 102 87673
rect 42 87649 76 87665
rect 16 87629 38 87635
rect 42 87626 76 87630
rect 80 87629 102 87635
rect 42 87596 46 87626
rect 72 87596 76 87626
rect 42 87515 46 87549
rect 72 87515 76 87549
rect -25 87478 25 87480
rect -8 87470 14 87477
rect -8 87469 17 87470
rect 25 87469 27 87478
rect -12 87462 38 87469
rect -12 87461 34 87462
rect -12 87457 8 87461
rect 0 87445 8 87457
rect 14 87445 34 87461
rect 0 87444 34 87445
rect 0 87437 38 87444
rect 14 87436 17 87437
rect 25 87428 27 87437
rect 42 87408 45 87498
rect 69 87483 80 87515
rect 107 87483 143 87511
rect 144 87483 148 87703
rect 332 87635 336 87703
rect 380 87673 462 87705
rect 463 87673 472 87707
rect 480 87673 497 87707
rect 378 87665 464 87673
rect 505 87665 507 87715
rect 514 87673 548 87707
rect 565 87673 582 87707
rect 607 87665 609 87715
rect 404 87649 438 87665
rect 400 87635 442 87636
rect 378 87629 404 87635
rect 442 87629 464 87635
rect 400 87628 404 87629
rect 174 87589 246 87597
rect 295 87594 300 87628
rect 324 87594 329 87628
rect 224 87559 226 87575
rect 196 87551 226 87559
rect 332 87557 336 87625
rect 367 87594 438 87628
rect 400 87587 404 87594
rect 454 87581 504 87583
rect 494 87577 548 87581
rect 494 87572 514 87577
rect 504 87557 506 87572
rect 196 87547 232 87551
rect 196 87517 204 87547
rect 216 87517 232 87547
rect 400 87549 404 87557
rect 107 87477 119 87483
rect 109 87449 119 87477
rect 129 87449 149 87483
rect 174 87479 181 87509
rect 224 87470 226 87517
rect 256 87509 328 87517
rect 332 87515 336 87545
rect 400 87515 408 87549
rect 434 87515 438 87549
rect 498 87547 506 87557
rect 514 87547 515 87567
rect 504 87531 506 87547
rect 525 87538 528 87572
rect 547 87547 548 87567
rect 557 87547 564 87557
rect 514 87531 530 87537
rect 532 87531 548 87537
rect 278 87479 305 87490
rect 42 87357 46 87391
rect 72 87357 76 87391
rect 38 87319 80 87320
rect 42 87278 76 87312
rect 79 87278 113 87312
rect 42 87199 46 87233
rect 72 87199 76 87233
rect -25 87162 25 87164
rect -8 87154 14 87161
rect -8 87153 17 87154
rect 25 87153 27 87162
rect -12 87146 38 87153
rect -12 87145 34 87146
rect -12 87141 8 87145
rect 0 87129 8 87141
rect 14 87129 34 87145
rect 0 87128 34 87129
rect 0 87121 38 87128
rect 14 87120 17 87121
rect 25 87112 27 87121
rect 42 87092 45 87182
rect 71 87151 80 87179
rect 69 87113 80 87151
rect 144 87141 148 87449
rect 196 87436 204 87470
rect 216 87436 232 87470
rect 244 87466 257 87470
rect 300 87466 308 87479
rect 332 87477 342 87515
rect 400 87507 404 87515
rect 336 87467 342 87477
rect 244 87442 291 87466
rect 244 87436 257 87442
rect 224 87389 226 87436
rect 278 87432 291 87442
rect 300 87442 329 87466
rect 332 87457 342 87467
rect 400 87467 409 87495
rect 562 87478 612 87480
rect 466 87469 497 87477
rect 565 87469 596 87477
rect 300 87432 321 87442
rect 300 87426 308 87432
rect 289 87416 308 87426
rect 196 87359 204 87389
rect 216 87359 232 87389
rect 196 87355 232 87359
rect 196 87347 226 87355
rect 300 87347 308 87416
rect 332 87423 351 87457
rect 361 87429 381 87457
rect 361 87423 375 87429
rect 400 87423 411 87467
rect 442 87462 500 87469
rect 466 87461 500 87462
rect 565 87461 599 87469
rect 497 87445 500 87461
rect 596 87445 599 87461
rect 466 87444 500 87445
rect 442 87437 500 87444
rect 565 87437 599 87445
rect 612 87428 614 87478
rect 332 87399 342 87423
rect 336 87387 342 87399
rect 224 87331 226 87347
rect 332 87319 342 87387
rect 400 87391 404 87399
rect 400 87357 408 87391
rect 434 87357 438 87391
rect 454 87375 504 87377
rect 504 87359 506 87375
rect 514 87369 530 87375
rect 532 87369 548 87375
rect 525 87359 548 87368
rect 400 87349 404 87357
rect 498 87349 506 87359
rect 504 87325 506 87349
rect 514 87339 515 87359
rect 525 87334 528 87359
rect 547 87339 548 87359
rect 557 87349 564 87359
rect 514 87325 548 87329
rect 151 87278 156 87312
rect 174 87309 246 87317
rect 256 87309 328 87317
rect 336 87311 342 87319
rect 400 87314 404 87319
rect 180 87281 185 87309
rect 174 87273 246 87281
rect 256 87273 328 87281
rect 332 87279 336 87309
rect 400 87280 438 87314
rect 224 87243 226 87259
rect 196 87235 226 87243
rect 196 87231 232 87235
rect 196 87201 204 87231
rect 216 87201 232 87231
rect 224 87154 226 87201
rect 300 87174 308 87243
rect 332 87241 342 87279
rect 400 87271 404 87280
rect 454 87265 504 87267
rect 494 87261 548 87265
rect 494 87256 514 87261
rect 504 87241 506 87256
rect 336 87229 342 87241
rect 289 87164 308 87174
rect 300 87158 308 87164
rect 332 87195 342 87229
rect 400 87233 404 87241
rect 400 87199 408 87233
rect 434 87199 438 87233
rect 498 87231 506 87241
rect 514 87231 515 87251
rect 504 87215 506 87231
rect 525 87222 528 87256
rect 547 87231 548 87251
rect 557 87231 564 87241
rect 514 87215 530 87221
rect 532 87215 548 87221
rect 332 87167 373 87195
rect 332 87161 351 87167
rect 107 87107 119 87141
rect 129 87107 149 87141
rect 196 87120 204 87154
rect 216 87120 232 87154
rect 244 87148 257 87154
rect 278 87148 291 87158
rect 244 87124 291 87148
rect 300 87148 321 87158
rect 336 87151 351 87161
rect 300 87124 329 87148
rect 332 87133 351 87151
rect 361 87161 375 87167
rect 400 87161 411 87199
rect 562 87162 612 87164
rect 361 87133 381 87161
rect 400 87133 409 87161
rect 466 87153 497 87161
rect 565 87153 596 87161
rect 442 87146 500 87153
rect 466 87145 500 87146
rect 565 87145 599 87153
rect 244 87120 257 87124
rect 42 87041 46 87075
rect 72 87041 76 87075
rect 42 86994 76 86998
rect 42 86979 46 86994
rect 72 86979 76 86994
rect 38 86961 80 86979
rect 16 86955 102 86961
rect 144 86955 148 87107
rect 174 87083 181 87111
rect 224 87073 226 87120
rect 300 87111 308 87124
rect 278 87100 305 87111
rect 332 87083 342 87133
rect 400 87113 404 87133
rect 497 87129 500 87145
rect 596 87129 599 87145
rect 466 87128 500 87129
rect 442 87121 500 87128
rect 565 87121 599 87129
rect 612 87112 614 87162
rect 256 87073 328 87081
rect 336 87075 342 87083
rect 400 87075 404 87083
rect 196 87043 204 87073
rect 216 87043 232 87073
rect 196 87039 232 87043
rect 196 87031 226 87039
rect 224 87015 226 87031
rect 332 87003 336 87071
rect 400 87041 408 87075
rect 434 87041 438 87075
rect 454 87059 504 87061
rect 504 87043 506 87059
rect 514 87053 530 87059
rect 532 87053 548 87059
rect 525 87043 548 87052
rect 400 87033 404 87041
rect 498 87033 506 87043
rect 504 87009 506 87033
rect 514 87023 515 87043
rect 525 87018 528 87043
rect 547 87023 548 87043
rect 557 87033 564 87043
rect 514 87009 548 87013
rect 400 87003 442 87004
rect 174 86993 246 87001
rect 400 86996 404 87003
rect 295 86962 300 86996
rect 324 86962 329 86996
rect 367 86979 438 86996
rect 367 86962 442 86979
rect 400 86961 442 86962
rect 378 86955 464 86961
rect 38 86939 80 86955
rect 400 86939 442 86955
rect -25 86925 25 86927
rect 42 86925 76 86939
rect 404 86925 438 86939
rect 455 86925 505 86927
rect 557 86925 607 86927
rect 16 86917 102 86925
rect 378 86917 464 86925
rect 8 86883 17 86917
rect 18 86915 51 86917
rect 80 86915 100 86917
rect 18 86883 100 86915
rect 380 86915 404 86917
rect 429 86915 438 86917
rect 442 86915 462 86917
rect 16 86875 102 86883
rect 42 86859 76 86875
rect 16 86839 38 86845
rect 42 86836 76 86840
rect 80 86839 102 86845
rect 42 86806 46 86836
rect 72 86806 76 86836
rect 42 86725 46 86759
rect 72 86725 76 86759
rect -25 86688 25 86690
rect -8 86680 14 86687
rect -8 86679 17 86680
rect 25 86679 27 86688
rect -12 86672 38 86679
rect -12 86671 34 86672
rect -12 86667 8 86671
rect 0 86655 8 86667
rect 14 86655 34 86671
rect 0 86654 34 86655
rect 0 86647 38 86654
rect 14 86646 17 86647
rect 25 86638 27 86647
rect 42 86618 45 86708
rect 69 86693 80 86725
rect 107 86693 143 86721
rect 144 86693 148 86913
rect 332 86845 336 86913
rect 380 86883 462 86915
rect 463 86883 472 86917
rect 480 86883 497 86917
rect 378 86875 464 86883
rect 505 86875 507 86925
rect 514 86883 548 86917
rect 565 86883 582 86917
rect 607 86875 609 86925
rect 404 86859 438 86875
rect 400 86845 442 86846
rect 378 86839 404 86845
rect 442 86839 464 86845
rect 400 86838 404 86839
rect 174 86799 246 86807
rect 295 86804 300 86838
rect 324 86804 329 86838
rect 224 86769 226 86785
rect 196 86761 226 86769
rect 332 86767 336 86835
rect 367 86804 438 86838
rect 400 86797 404 86804
rect 454 86791 504 86793
rect 494 86787 548 86791
rect 494 86782 514 86787
rect 504 86767 506 86782
rect 196 86757 232 86761
rect 196 86727 204 86757
rect 216 86727 232 86757
rect 400 86759 404 86767
rect 107 86687 119 86693
rect 109 86659 119 86687
rect 129 86659 149 86693
rect 174 86689 181 86719
rect 224 86680 226 86727
rect 256 86719 328 86727
rect 332 86725 336 86755
rect 400 86725 408 86759
rect 434 86725 438 86759
rect 498 86757 506 86767
rect 514 86757 515 86777
rect 504 86741 506 86757
rect 525 86748 528 86782
rect 547 86757 548 86777
rect 557 86757 564 86767
rect 514 86741 530 86747
rect 532 86741 548 86747
rect 278 86689 305 86700
rect 42 86567 46 86601
rect 72 86567 76 86601
rect 38 86529 80 86530
rect 42 86488 76 86522
rect 79 86488 113 86522
rect 42 86409 46 86443
rect 72 86409 76 86443
rect -25 86372 25 86374
rect -8 86364 14 86371
rect -8 86363 17 86364
rect 25 86363 27 86372
rect -12 86356 38 86363
rect -12 86355 34 86356
rect -12 86351 8 86355
rect 0 86339 8 86351
rect 14 86339 34 86355
rect 0 86338 34 86339
rect 0 86331 38 86338
rect 14 86330 17 86331
rect 25 86322 27 86331
rect 42 86302 45 86392
rect 71 86361 80 86389
rect 69 86323 80 86361
rect 144 86351 148 86659
rect 196 86646 204 86680
rect 216 86646 232 86680
rect 244 86676 257 86680
rect 300 86676 308 86689
rect 332 86687 342 86725
rect 400 86717 404 86725
rect 336 86677 342 86687
rect 244 86652 291 86676
rect 244 86646 257 86652
rect 224 86599 226 86646
rect 278 86642 291 86652
rect 300 86652 329 86676
rect 332 86667 342 86677
rect 400 86677 409 86705
rect 562 86688 612 86690
rect 466 86679 497 86687
rect 565 86679 596 86687
rect 300 86642 321 86652
rect 300 86636 308 86642
rect 289 86626 308 86636
rect 196 86569 204 86599
rect 216 86569 232 86599
rect 196 86565 232 86569
rect 196 86557 226 86565
rect 300 86557 308 86626
rect 332 86633 351 86667
rect 361 86639 381 86667
rect 361 86633 375 86639
rect 400 86633 411 86677
rect 442 86672 500 86679
rect 466 86671 500 86672
rect 565 86671 599 86679
rect 497 86655 500 86671
rect 596 86655 599 86671
rect 466 86654 500 86655
rect 442 86647 500 86654
rect 565 86647 599 86655
rect 612 86638 614 86688
rect 332 86609 342 86633
rect 336 86597 342 86609
rect 224 86541 226 86557
rect 332 86529 342 86597
rect 400 86601 404 86609
rect 400 86567 408 86601
rect 434 86567 438 86601
rect 454 86585 504 86587
rect 504 86569 506 86585
rect 514 86579 530 86585
rect 532 86579 548 86585
rect 525 86569 548 86578
rect 400 86559 404 86567
rect 498 86559 506 86569
rect 504 86535 506 86559
rect 514 86549 515 86569
rect 525 86544 528 86569
rect 547 86549 548 86569
rect 557 86559 564 86569
rect 514 86535 548 86539
rect 151 86488 156 86522
rect 174 86519 246 86527
rect 256 86519 328 86527
rect 336 86521 342 86529
rect 400 86524 404 86529
rect 180 86491 185 86519
rect 174 86483 246 86491
rect 256 86483 328 86491
rect 332 86489 336 86519
rect 400 86490 438 86524
rect 224 86453 226 86469
rect 196 86445 226 86453
rect 196 86441 232 86445
rect 196 86411 204 86441
rect 216 86411 232 86441
rect 224 86364 226 86411
rect 300 86384 308 86453
rect 332 86451 342 86489
rect 400 86481 404 86490
rect 454 86475 504 86477
rect 494 86471 548 86475
rect 494 86466 514 86471
rect 504 86451 506 86466
rect 336 86439 342 86451
rect 289 86374 308 86384
rect 300 86368 308 86374
rect 332 86405 342 86439
rect 400 86443 404 86451
rect 400 86409 408 86443
rect 434 86409 438 86443
rect 498 86441 506 86451
rect 514 86441 515 86461
rect 504 86425 506 86441
rect 525 86432 528 86466
rect 547 86441 548 86461
rect 557 86441 564 86451
rect 514 86425 530 86431
rect 532 86425 548 86431
rect 332 86377 373 86405
rect 332 86371 351 86377
rect 107 86317 119 86351
rect 129 86317 149 86351
rect 196 86330 204 86364
rect 216 86330 232 86364
rect 244 86358 257 86364
rect 278 86358 291 86368
rect 244 86334 291 86358
rect 300 86358 321 86368
rect 336 86361 351 86371
rect 300 86334 329 86358
rect 332 86343 351 86361
rect 361 86371 375 86377
rect 400 86371 411 86409
rect 562 86372 612 86374
rect 361 86343 381 86371
rect 400 86343 409 86371
rect 466 86363 497 86371
rect 565 86363 596 86371
rect 442 86356 500 86363
rect 466 86355 500 86356
rect 565 86355 599 86363
rect 244 86330 257 86334
rect 42 86251 46 86285
rect 72 86251 76 86285
rect 42 86204 76 86208
rect 42 86189 46 86204
rect 72 86189 76 86204
rect 38 86171 80 86189
rect 16 86165 102 86171
rect 144 86165 148 86317
rect 174 86293 181 86321
rect 224 86283 226 86330
rect 300 86321 308 86334
rect 278 86310 305 86321
rect 332 86293 342 86343
rect 400 86323 404 86343
rect 497 86339 500 86355
rect 596 86339 599 86355
rect 466 86338 500 86339
rect 442 86331 500 86338
rect 565 86331 599 86339
rect 612 86322 614 86372
rect 256 86283 328 86291
rect 336 86285 342 86293
rect 400 86285 404 86293
rect 196 86253 204 86283
rect 216 86253 232 86283
rect 196 86249 232 86253
rect 196 86241 226 86249
rect 224 86225 226 86241
rect 332 86213 336 86281
rect 400 86251 408 86285
rect 434 86251 438 86285
rect 454 86269 504 86271
rect 504 86253 506 86269
rect 514 86263 530 86269
rect 532 86263 548 86269
rect 525 86253 548 86262
rect 400 86243 404 86251
rect 498 86243 506 86253
rect 504 86219 506 86243
rect 514 86233 515 86253
rect 525 86228 528 86253
rect 547 86233 548 86253
rect 557 86243 564 86253
rect 514 86219 548 86223
rect 400 86213 442 86214
rect 174 86203 246 86211
rect 400 86206 404 86213
rect 295 86172 300 86206
rect 324 86172 329 86206
rect 367 86189 438 86206
rect 367 86172 442 86189
rect 400 86171 442 86172
rect 378 86165 464 86171
rect 38 86149 80 86165
rect 400 86149 442 86165
rect -25 86135 25 86137
rect 42 86135 76 86149
rect 404 86135 438 86149
rect 455 86135 505 86137
rect 557 86135 607 86137
rect 16 86127 102 86135
rect 378 86127 464 86135
rect 8 86093 17 86127
rect 18 86125 51 86127
rect 80 86125 100 86127
rect 18 86093 100 86125
rect 380 86125 404 86127
rect 429 86125 438 86127
rect 442 86125 462 86127
rect 16 86085 102 86093
rect 42 86069 76 86085
rect 16 86049 38 86055
rect 42 86046 76 86050
rect 80 86049 102 86055
rect 42 86016 46 86046
rect 72 86016 76 86046
rect 42 85935 46 85969
rect 72 85935 76 85969
rect -25 85898 25 85900
rect -8 85890 14 85897
rect -8 85889 17 85890
rect 25 85889 27 85898
rect -12 85882 38 85889
rect -12 85881 34 85882
rect -12 85877 8 85881
rect 0 85865 8 85877
rect 14 85865 34 85881
rect 0 85864 34 85865
rect 0 85857 38 85864
rect 14 85856 17 85857
rect 25 85848 27 85857
rect 42 85828 45 85918
rect 69 85903 80 85935
rect 107 85903 143 85931
rect 144 85903 148 86123
rect 332 86055 336 86123
rect 380 86093 462 86125
rect 463 86093 472 86127
rect 480 86093 497 86127
rect 378 86085 464 86093
rect 505 86085 507 86135
rect 514 86093 548 86127
rect 565 86093 582 86127
rect 607 86085 609 86135
rect 404 86069 438 86085
rect 400 86055 442 86056
rect 378 86049 404 86055
rect 442 86049 464 86055
rect 400 86048 404 86049
rect 174 86009 246 86017
rect 295 86014 300 86048
rect 324 86014 329 86048
rect 224 85979 226 85995
rect 196 85971 226 85979
rect 332 85977 336 86045
rect 367 86014 438 86048
rect 400 86007 404 86014
rect 454 86001 504 86003
rect 494 85997 548 86001
rect 494 85992 514 85997
rect 504 85977 506 85992
rect 196 85967 232 85971
rect 196 85937 204 85967
rect 216 85937 232 85967
rect 400 85969 404 85977
rect 107 85897 119 85903
rect 109 85869 119 85897
rect 129 85869 149 85903
rect 174 85899 181 85929
rect 224 85890 226 85937
rect 256 85929 328 85937
rect 332 85935 336 85965
rect 400 85935 408 85969
rect 434 85935 438 85969
rect 498 85967 506 85977
rect 514 85967 515 85987
rect 504 85951 506 85967
rect 525 85958 528 85992
rect 547 85967 548 85987
rect 557 85967 564 85977
rect 514 85951 530 85957
rect 532 85951 548 85957
rect 278 85899 305 85910
rect 42 85777 46 85811
rect 72 85777 76 85811
rect 38 85739 80 85740
rect 42 85698 76 85732
rect 79 85698 113 85732
rect 42 85619 46 85653
rect 72 85619 76 85653
rect -25 85582 25 85584
rect -8 85574 14 85581
rect -8 85573 17 85574
rect 25 85573 27 85582
rect -12 85566 38 85573
rect -12 85565 34 85566
rect -12 85561 8 85565
rect 0 85549 8 85561
rect 14 85549 34 85565
rect 0 85548 34 85549
rect 0 85541 38 85548
rect 14 85540 17 85541
rect 25 85532 27 85541
rect 42 85512 45 85602
rect 71 85571 80 85599
rect 69 85533 80 85571
rect 144 85561 148 85869
rect 196 85856 204 85890
rect 216 85856 232 85890
rect 244 85886 257 85890
rect 300 85886 308 85899
rect 332 85897 342 85935
rect 400 85927 404 85935
rect 336 85887 342 85897
rect 244 85862 291 85886
rect 244 85856 257 85862
rect 224 85809 226 85856
rect 278 85852 291 85862
rect 300 85862 329 85886
rect 332 85877 342 85887
rect 400 85887 409 85915
rect 562 85898 612 85900
rect 466 85889 497 85897
rect 565 85889 596 85897
rect 300 85852 321 85862
rect 300 85846 308 85852
rect 289 85836 308 85846
rect 196 85779 204 85809
rect 216 85779 232 85809
rect 196 85775 232 85779
rect 196 85767 226 85775
rect 300 85767 308 85836
rect 332 85843 351 85877
rect 361 85849 381 85877
rect 361 85843 375 85849
rect 400 85843 411 85887
rect 442 85882 500 85889
rect 466 85881 500 85882
rect 565 85881 599 85889
rect 497 85865 500 85881
rect 596 85865 599 85881
rect 466 85864 500 85865
rect 442 85857 500 85864
rect 565 85857 599 85865
rect 612 85848 614 85898
rect 332 85819 342 85843
rect 336 85807 342 85819
rect 224 85751 226 85767
rect 332 85739 342 85807
rect 400 85811 404 85819
rect 400 85777 408 85811
rect 434 85777 438 85811
rect 454 85795 504 85797
rect 504 85779 506 85795
rect 514 85789 530 85795
rect 532 85789 548 85795
rect 525 85779 548 85788
rect 400 85769 404 85777
rect 498 85769 506 85779
rect 504 85745 506 85769
rect 514 85759 515 85779
rect 525 85754 528 85779
rect 547 85759 548 85779
rect 557 85769 564 85779
rect 514 85745 548 85749
rect 151 85698 156 85732
rect 174 85729 246 85737
rect 256 85729 328 85737
rect 336 85731 342 85739
rect 400 85734 404 85739
rect 180 85701 185 85729
rect 174 85693 246 85701
rect 256 85693 328 85701
rect 332 85699 336 85729
rect 400 85700 438 85734
rect 224 85663 226 85679
rect 196 85655 226 85663
rect 196 85651 232 85655
rect 196 85621 204 85651
rect 216 85621 232 85651
rect 224 85574 226 85621
rect 300 85594 308 85663
rect 332 85661 342 85699
rect 400 85691 404 85700
rect 454 85685 504 85687
rect 494 85681 548 85685
rect 494 85676 514 85681
rect 504 85661 506 85676
rect 336 85649 342 85661
rect 289 85584 308 85594
rect 300 85578 308 85584
rect 332 85615 342 85649
rect 400 85653 404 85661
rect 400 85619 408 85653
rect 434 85619 438 85653
rect 498 85651 506 85661
rect 514 85651 515 85671
rect 504 85635 506 85651
rect 525 85642 528 85676
rect 547 85651 548 85671
rect 557 85651 564 85661
rect 514 85635 530 85641
rect 532 85635 548 85641
rect 332 85587 373 85615
rect 332 85581 351 85587
rect 107 85527 119 85561
rect 129 85527 149 85561
rect 196 85540 204 85574
rect 216 85540 232 85574
rect 244 85568 257 85574
rect 278 85568 291 85578
rect 244 85544 291 85568
rect 300 85568 321 85578
rect 336 85571 351 85581
rect 300 85544 329 85568
rect 332 85553 351 85571
rect 361 85581 375 85587
rect 400 85581 411 85619
rect 562 85582 612 85584
rect 361 85553 381 85581
rect 400 85553 409 85581
rect 466 85573 497 85581
rect 565 85573 596 85581
rect 442 85566 500 85573
rect 466 85565 500 85566
rect 565 85565 599 85573
rect 244 85540 257 85544
rect 42 85461 46 85495
rect 72 85461 76 85495
rect 42 85414 76 85418
rect 42 85399 46 85414
rect 72 85399 76 85414
rect 38 85381 80 85399
rect 16 85375 102 85381
rect 144 85375 148 85527
rect 174 85503 181 85531
rect 224 85493 226 85540
rect 300 85531 308 85544
rect 278 85520 305 85531
rect 332 85503 342 85553
rect 400 85533 404 85553
rect 497 85549 500 85565
rect 596 85549 599 85565
rect 466 85548 500 85549
rect 442 85541 500 85548
rect 565 85541 599 85549
rect 612 85532 614 85582
rect 256 85493 328 85501
rect 336 85495 342 85503
rect 400 85495 404 85503
rect 196 85463 204 85493
rect 216 85463 232 85493
rect 196 85459 232 85463
rect 196 85451 226 85459
rect 224 85435 226 85451
rect 332 85423 336 85491
rect 400 85461 408 85495
rect 434 85461 438 85495
rect 454 85479 504 85481
rect 504 85463 506 85479
rect 514 85473 530 85479
rect 532 85473 548 85479
rect 525 85463 548 85472
rect 400 85453 404 85461
rect 498 85453 506 85463
rect 504 85429 506 85453
rect 514 85443 515 85463
rect 525 85438 528 85463
rect 547 85443 548 85463
rect 557 85453 564 85463
rect 514 85429 548 85433
rect 400 85423 442 85424
rect 174 85413 246 85421
rect 400 85416 404 85423
rect 295 85382 300 85416
rect 324 85382 329 85416
rect 367 85399 438 85416
rect 367 85382 442 85399
rect 400 85381 442 85382
rect 378 85375 464 85381
rect 38 85359 80 85375
rect 400 85359 442 85375
rect -25 85345 25 85347
rect 42 85345 76 85359
rect 404 85345 438 85359
rect 455 85345 505 85347
rect 557 85345 607 85347
rect 16 85337 102 85345
rect 378 85337 464 85345
rect 8 85303 17 85337
rect 18 85335 51 85337
rect 80 85335 100 85337
rect 18 85303 100 85335
rect 380 85335 404 85337
rect 429 85335 438 85337
rect 442 85335 462 85337
rect 16 85295 102 85303
rect 42 85279 76 85295
rect 16 85259 38 85265
rect 42 85256 76 85260
rect 80 85259 102 85265
rect 42 85226 46 85256
rect 72 85226 76 85256
rect 42 85145 46 85179
rect 72 85145 76 85179
rect -25 85108 25 85110
rect -8 85100 14 85107
rect -8 85099 17 85100
rect 25 85099 27 85108
rect -12 85092 38 85099
rect -12 85091 34 85092
rect -12 85087 8 85091
rect 0 85075 8 85087
rect 14 85075 34 85091
rect 0 85074 34 85075
rect 0 85067 38 85074
rect 14 85066 17 85067
rect 25 85058 27 85067
rect 42 85038 45 85128
rect 69 85113 80 85145
rect 107 85113 143 85141
rect 144 85113 148 85333
rect 332 85265 336 85333
rect 380 85303 462 85335
rect 463 85303 472 85337
rect 480 85303 497 85337
rect 378 85295 464 85303
rect 505 85295 507 85345
rect 514 85303 548 85337
rect 565 85303 582 85337
rect 607 85295 609 85345
rect 404 85279 438 85295
rect 400 85265 442 85266
rect 378 85259 404 85265
rect 442 85259 464 85265
rect 400 85258 404 85259
rect 174 85219 246 85227
rect 295 85224 300 85258
rect 324 85224 329 85258
rect 224 85189 226 85205
rect 196 85181 226 85189
rect 332 85187 336 85255
rect 367 85224 438 85258
rect 400 85217 404 85224
rect 454 85211 504 85213
rect 494 85207 548 85211
rect 494 85202 514 85207
rect 504 85187 506 85202
rect 196 85177 232 85181
rect 196 85147 204 85177
rect 216 85147 232 85177
rect 400 85179 404 85187
rect 107 85107 119 85113
rect 109 85079 119 85107
rect 129 85079 149 85113
rect 174 85109 181 85139
rect 224 85100 226 85147
rect 256 85139 328 85147
rect 332 85145 336 85175
rect 400 85145 408 85179
rect 434 85145 438 85179
rect 498 85177 506 85187
rect 514 85177 515 85197
rect 504 85161 506 85177
rect 525 85168 528 85202
rect 547 85177 548 85197
rect 557 85177 564 85187
rect 514 85161 530 85167
rect 532 85161 548 85167
rect 278 85109 305 85120
rect 42 84987 46 85021
rect 72 84987 76 85021
rect 38 84949 80 84950
rect 42 84908 76 84942
rect 79 84908 113 84942
rect 42 84829 46 84863
rect 72 84829 76 84863
rect -25 84792 25 84794
rect -8 84784 14 84791
rect -8 84783 17 84784
rect 25 84783 27 84792
rect -12 84776 38 84783
rect -12 84775 34 84776
rect -12 84771 8 84775
rect 0 84759 8 84771
rect 14 84759 34 84775
rect 0 84758 34 84759
rect 0 84751 38 84758
rect 14 84750 17 84751
rect 25 84742 27 84751
rect 42 84722 45 84812
rect 71 84781 80 84809
rect 69 84743 80 84781
rect 144 84771 148 85079
rect 196 85066 204 85100
rect 216 85066 232 85100
rect 244 85096 257 85100
rect 300 85096 308 85109
rect 332 85107 342 85145
rect 400 85137 404 85145
rect 336 85097 342 85107
rect 244 85072 291 85096
rect 244 85066 257 85072
rect 224 85019 226 85066
rect 278 85062 291 85072
rect 300 85072 329 85096
rect 332 85087 342 85097
rect 400 85097 409 85125
rect 562 85108 612 85110
rect 466 85099 497 85107
rect 565 85099 596 85107
rect 300 85062 321 85072
rect 300 85056 308 85062
rect 289 85046 308 85056
rect 196 84989 204 85019
rect 216 84989 232 85019
rect 196 84985 232 84989
rect 196 84977 226 84985
rect 300 84977 308 85046
rect 332 85053 351 85087
rect 361 85059 381 85087
rect 361 85053 375 85059
rect 400 85053 411 85097
rect 442 85092 500 85099
rect 466 85091 500 85092
rect 565 85091 599 85099
rect 497 85075 500 85091
rect 596 85075 599 85091
rect 466 85074 500 85075
rect 442 85067 500 85074
rect 565 85067 599 85075
rect 612 85058 614 85108
rect 332 85029 342 85053
rect 336 85017 342 85029
rect 224 84961 226 84977
rect 332 84949 342 85017
rect 400 85021 404 85029
rect 400 84987 408 85021
rect 434 84987 438 85021
rect 454 85005 504 85007
rect 504 84989 506 85005
rect 514 84999 530 85005
rect 532 84999 548 85005
rect 525 84989 548 84998
rect 400 84979 404 84987
rect 498 84979 506 84989
rect 504 84955 506 84979
rect 514 84969 515 84989
rect 525 84964 528 84989
rect 547 84969 548 84989
rect 557 84979 564 84989
rect 514 84955 548 84959
rect 151 84908 156 84942
rect 174 84939 246 84947
rect 256 84939 328 84947
rect 336 84941 342 84949
rect 400 84944 404 84949
rect 180 84911 185 84939
rect 174 84903 246 84911
rect 256 84903 328 84911
rect 332 84909 336 84939
rect 400 84910 438 84944
rect 224 84873 226 84889
rect 196 84865 226 84873
rect 196 84861 232 84865
rect 196 84831 204 84861
rect 216 84831 232 84861
rect 224 84784 226 84831
rect 300 84804 308 84873
rect 332 84871 342 84909
rect 400 84901 404 84910
rect 454 84895 504 84897
rect 494 84891 548 84895
rect 494 84886 514 84891
rect 504 84871 506 84886
rect 336 84859 342 84871
rect 289 84794 308 84804
rect 300 84788 308 84794
rect 332 84825 342 84859
rect 400 84863 404 84871
rect 400 84829 408 84863
rect 434 84829 438 84863
rect 498 84861 506 84871
rect 514 84861 515 84881
rect 504 84845 506 84861
rect 525 84852 528 84886
rect 547 84861 548 84881
rect 557 84861 564 84871
rect 514 84845 530 84851
rect 532 84845 548 84851
rect 332 84797 373 84825
rect 332 84791 351 84797
rect 107 84737 119 84771
rect 129 84737 149 84771
rect 196 84750 204 84784
rect 216 84750 232 84784
rect 244 84778 257 84784
rect 278 84778 291 84788
rect 244 84754 291 84778
rect 300 84778 321 84788
rect 336 84781 351 84791
rect 300 84754 329 84778
rect 332 84763 351 84781
rect 361 84791 375 84797
rect 400 84791 411 84829
rect 562 84792 612 84794
rect 361 84763 381 84791
rect 400 84763 409 84791
rect 466 84783 497 84791
rect 565 84783 596 84791
rect 442 84776 500 84783
rect 466 84775 500 84776
rect 565 84775 599 84783
rect 244 84750 257 84754
rect 42 84671 46 84705
rect 72 84671 76 84705
rect 42 84624 76 84628
rect 42 84609 46 84624
rect 72 84609 76 84624
rect 38 84591 80 84609
rect 16 84585 102 84591
rect 144 84585 148 84737
rect 174 84713 181 84741
rect 224 84703 226 84750
rect 300 84741 308 84754
rect 278 84730 305 84741
rect 332 84713 342 84763
rect 400 84743 404 84763
rect 497 84759 500 84775
rect 596 84759 599 84775
rect 466 84758 500 84759
rect 442 84751 500 84758
rect 565 84751 599 84759
rect 612 84742 614 84792
rect 256 84703 328 84711
rect 336 84705 342 84713
rect 400 84705 404 84713
rect 196 84673 204 84703
rect 216 84673 232 84703
rect 196 84669 232 84673
rect 196 84661 226 84669
rect 224 84645 226 84661
rect 332 84633 336 84701
rect 400 84671 408 84705
rect 434 84671 438 84705
rect 454 84689 504 84691
rect 504 84673 506 84689
rect 514 84683 530 84689
rect 532 84683 548 84689
rect 525 84673 548 84682
rect 400 84663 404 84671
rect 498 84663 506 84673
rect 504 84639 506 84663
rect 514 84653 515 84673
rect 525 84648 528 84673
rect 547 84653 548 84673
rect 557 84663 564 84673
rect 514 84639 548 84643
rect 400 84633 442 84634
rect 174 84623 246 84631
rect 400 84626 404 84633
rect 295 84592 300 84626
rect 324 84592 329 84626
rect 367 84609 438 84626
rect 367 84592 442 84609
rect 400 84591 442 84592
rect 378 84585 464 84591
rect 38 84569 80 84585
rect 400 84569 442 84585
rect -25 84555 25 84557
rect 42 84555 76 84569
rect 404 84555 438 84569
rect 455 84555 505 84557
rect 557 84555 607 84557
rect 16 84547 102 84555
rect 378 84547 464 84555
rect 8 84513 17 84547
rect 18 84545 51 84547
rect 80 84545 100 84547
rect 18 84513 100 84545
rect 380 84545 404 84547
rect 429 84545 438 84547
rect 442 84545 462 84547
rect 16 84505 102 84513
rect 42 84489 76 84505
rect 16 84469 38 84475
rect 42 84466 76 84470
rect 80 84469 102 84475
rect 42 84436 46 84466
rect 72 84436 76 84466
rect 42 84355 46 84389
rect 72 84355 76 84389
rect -25 84318 25 84320
rect -8 84310 14 84317
rect -8 84309 17 84310
rect 25 84309 27 84318
rect -12 84302 38 84309
rect -12 84301 34 84302
rect -12 84297 8 84301
rect 0 84285 8 84297
rect 14 84285 34 84301
rect 0 84284 34 84285
rect 0 84277 38 84284
rect 14 84276 17 84277
rect 25 84268 27 84277
rect 42 84248 45 84338
rect 69 84323 80 84355
rect 107 84323 143 84351
rect 144 84323 148 84543
rect 332 84475 336 84543
rect 380 84513 462 84545
rect 463 84513 472 84547
rect 480 84513 497 84547
rect 378 84505 464 84513
rect 505 84505 507 84555
rect 514 84513 548 84547
rect 565 84513 582 84547
rect 607 84505 609 84555
rect 404 84489 438 84505
rect 400 84475 442 84476
rect 378 84469 404 84475
rect 442 84469 464 84475
rect 400 84468 404 84469
rect 174 84429 246 84437
rect 295 84434 300 84468
rect 324 84434 329 84468
rect 224 84399 226 84415
rect 196 84391 226 84399
rect 332 84397 336 84465
rect 367 84434 438 84468
rect 400 84427 404 84434
rect 454 84421 504 84423
rect 494 84417 548 84421
rect 494 84412 514 84417
rect 504 84397 506 84412
rect 196 84387 232 84391
rect 196 84357 204 84387
rect 216 84357 232 84387
rect 400 84389 404 84397
rect 107 84317 119 84323
rect 109 84289 119 84317
rect 129 84289 149 84323
rect 174 84319 181 84349
rect 224 84310 226 84357
rect 256 84349 328 84357
rect 332 84355 336 84385
rect 400 84355 408 84389
rect 434 84355 438 84389
rect 498 84387 506 84397
rect 514 84387 515 84407
rect 504 84371 506 84387
rect 525 84378 528 84412
rect 547 84387 548 84407
rect 557 84387 564 84397
rect 514 84371 530 84377
rect 532 84371 548 84377
rect 278 84319 305 84330
rect 42 84197 46 84231
rect 72 84197 76 84231
rect 38 84159 80 84160
rect 42 84118 76 84152
rect 79 84118 113 84152
rect 42 84039 46 84073
rect 72 84039 76 84073
rect -25 84002 25 84004
rect -8 83994 14 84001
rect -8 83993 17 83994
rect 25 83993 27 84002
rect -12 83986 38 83993
rect -12 83985 34 83986
rect -12 83981 8 83985
rect 0 83969 8 83981
rect 14 83969 34 83985
rect 0 83968 34 83969
rect 0 83961 38 83968
rect 14 83960 17 83961
rect 25 83952 27 83961
rect 42 83932 45 84022
rect 71 83991 80 84019
rect 69 83953 80 83991
rect 144 83981 148 84289
rect 196 84276 204 84310
rect 216 84276 232 84310
rect 244 84306 257 84310
rect 300 84306 308 84319
rect 332 84317 342 84355
rect 400 84347 404 84355
rect 336 84307 342 84317
rect 244 84282 291 84306
rect 244 84276 257 84282
rect 224 84229 226 84276
rect 278 84272 291 84282
rect 300 84282 329 84306
rect 332 84297 342 84307
rect 400 84307 409 84335
rect 562 84318 612 84320
rect 466 84309 497 84317
rect 565 84309 596 84317
rect 300 84272 321 84282
rect 300 84266 308 84272
rect 289 84256 308 84266
rect 196 84199 204 84229
rect 216 84199 232 84229
rect 196 84195 232 84199
rect 196 84187 226 84195
rect 300 84187 308 84256
rect 332 84263 351 84297
rect 361 84269 381 84297
rect 361 84263 375 84269
rect 400 84263 411 84307
rect 442 84302 500 84309
rect 466 84301 500 84302
rect 565 84301 599 84309
rect 497 84285 500 84301
rect 596 84285 599 84301
rect 466 84284 500 84285
rect 442 84277 500 84284
rect 565 84277 599 84285
rect 612 84268 614 84318
rect 332 84239 342 84263
rect 336 84227 342 84239
rect 224 84171 226 84187
rect 332 84159 342 84227
rect 400 84231 404 84239
rect 400 84197 408 84231
rect 434 84197 438 84231
rect 454 84215 504 84217
rect 504 84199 506 84215
rect 514 84209 530 84215
rect 532 84209 548 84215
rect 525 84199 548 84208
rect 400 84189 404 84197
rect 498 84189 506 84199
rect 504 84165 506 84189
rect 514 84179 515 84199
rect 525 84174 528 84199
rect 547 84179 548 84199
rect 557 84189 564 84199
rect 514 84165 548 84169
rect 151 84118 156 84152
rect 174 84149 246 84157
rect 256 84149 328 84157
rect 336 84151 342 84159
rect 400 84154 404 84159
rect 180 84121 185 84149
rect 174 84113 246 84121
rect 256 84113 328 84121
rect 332 84119 336 84149
rect 400 84120 438 84154
rect 224 84083 226 84099
rect 196 84075 226 84083
rect 196 84071 232 84075
rect 196 84041 204 84071
rect 216 84041 232 84071
rect 224 83994 226 84041
rect 300 84014 308 84083
rect 332 84081 342 84119
rect 400 84111 404 84120
rect 454 84105 504 84107
rect 494 84101 548 84105
rect 494 84096 514 84101
rect 504 84081 506 84096
rect 336 84069 342 84081
rect 289 84004 308 84014
rect 300 83998 308 84004
rect 332 84035 342 84069
rect 400 84073 404 84081
rect 400 84039 408 84073
rect 434 84039 438 84073
rect 498 84071 506 84081
rect 514 84071 515 84091
rect 504 84055 506 84071
rect 525 84062 528 84096
rect 547 84071 548 84091
rect 557 84071 564 84081
rect 514 84055 530 84061
rect 532 84055 548 84061
rect 332 84007 373 84035
rect 332 84001 351 84007
rect 107 83947 119 83981
rect 129 83947 149 83981
rect 196 83960 204 83994
rect 216 83960 232 83994
rect 244 83988 257 83994
rect 278 83988 291 83998
rect 244 83964 291 83988
rect 300 83988 321 83998
rect 336 83991 351 84001
rect 300 83964 329 83988
rect 332 83973 351 83991
rect 361 84001 375 84007
rect 400 84001 411 84039
rect 562 84002 612 84004
rect 361 83973 381 84001
rect 400 83973 409 84001
rect 466 83993 497 84001
rect 565 83993 596 84001
rect 442 83986 500 83993
rect 466 83985 500 83986
rect 565 83985 599 83993
rect 244 83960 257 83964
rect 42 83881 46 83915
rect 72 83881 76 83915
rect 42 83834 76 83838
rect 42 83819 46 83834
rect 72 83819 76 83834
rect 38 83801 80 83819
rect 16 83795 102 83801
rect 144 83795 148 83947
rect 174 83923 181 83951
rect 224 83913 226 83960
rect 300 83951 308 83964
rect 278 83940 305 83951
rect 332 83923 342 83973
rect 400 83953 404 83973
rect 497 83969 500 83985
rect 596 83969 599 83985
rect 466 83968 500 83969
rect 442 83961 500 83968
rect 565 83961 599 83969
rect 612 83952 614 84002
rect 256 83913 328 83921
rect 336 83915 342 83923
rect 400 83915 404 83923
rect 196 83883 204 83913
rect 216 83883 232 83913
rect 196 83879 232 83883
rect 196 83871 226 83879
rect 224 83855 226 83871
rect 332 83843 336 83911
rect 400 83881 408 83915
rect 434 83881 438 83915
rect 454 83899 504 83901
rect 504 83883 506 83899
rect 514 83893 530 83899
rect 532 83893 548 83899
rect 525 83883 548 83892
rect 400 83873 404 83881
rect 498 83873 506 83883
rect 504 83849 506 83873
rect 514 83863 515 83883
rect 525 83858 528 83883
rect 547 83863 548 83883
rect 557 83873 564 83883
rect 514 83849 548 83853
rect 400 83843 442 83844
rect 174 83833 246 83841
rect 400 83836 404 83843
rect 295 83802 300 83836
rect 324 83802 329 83836
rect 367 83819 438 83836
rect 367 83802 442 83819
rect 400 83801 442 83802
rect 378 83795 464 83801
rect 38 83779 80 83795
rect 400 83779 442 83795
rect -25 83765 25 83767
rect 42 83765 76 83779
rect 404 83765 438 83779
rect 455 83765 505 83767
rect 557 83765 607 83767
rect 16 83757 102 83765
rect 378 83757 464 83765
rect 8 83723 17 83757
rect 18 83755 51 83757
rect 80 83755 100 83757
rect 18 83723 100 83755
rect 380 83755 404 83757
rect 429 83755 438 83757
rect 442 83755 462 83757
rect 16 83715 102 83723
rect 42 83699 76 83715
rect 16 83679 38 83685
rect 42 83676 76 83680
rect 80 83679 102 83685
rect 42 83646 46 83676
rect 72 83646 76 83676
rect 42 83565 46 83599
rect 72 83565 76 83599
rect -25 83528 25 83530
rect -8 83520 14 83527
rect -8 83519 17 83520
rect 25 83519 27 83528
rect -12 83512 38 83519
rect -12 83511 34 83512
rect -12 83507 8 83511
rect 0 83495 8 83507
rect 14 83495 34 83511
rect 0 83494 34 83495
rect 0 83487 38 83494
rect 14 83486 17 83487
rect 25 83478 27 83487
rect 42 83458 45 83548
rect 69 83533 80 83565
rect 107 83533 143 83561
rect 144 83533 148 83753
rect 332 83685 336 83753
rect 380 83723 462 83755
rect 463 83723 472 83757
rect 480 83723 497 83757
rect 378 83715 464 83723
rect 505 83715 507 83765
rect 514 83723 548 83757
rect 565 83723 582 83757
rect 607 83715 609 83765
rect 404 83699 438 83715
rect 400 83685 442 83686
rect 378 83679 404 83685
rect 442 83679 464 83685
rect 400 83678 404 83679
rect 174 83639 246 83647
rect 295 83644 300 83678
rect 324 83644 329 83678
rect 224 83609 226 83625
rect 196 83601 226 83609
rect 332 83607 336 83675
rect 367 83644 438 83678
rect 400 83637 404 83644
rect 454 83631 504 83633
rect 494 83627 548 83631
rect 494 83622 514 83627
rect 504 83607 506 83622
rect 196 83597 232 83601
rect 196 83567 204 83597
rect 216 83567 232 83597
rect 400 83599 404 83607
rect 107 83527 119 83533
rect 109 83499 119 83527
rect 129 83499 149 83533
rect 174 83529 181 83559
rect 224 83520 226 83567
rect 256 83559 328 83567
rect 332 83565 336 83595
rect 400 83565 408 83599
rect 434 83565 438 83599
rect 498 83597 506 83607
rect 514 83597 515 83617
rect 504 83581 506 83597
rect 525 83588 528 83622
rect 547 83597 548 83617
rect 557 83597 564 83607
rect 514 83581 530 83587
rect 532 83581 548 83587
rect 278 83529 305 83540
rect 42 83407 46 83441
rect 72 83407 76 83441
rect 38 83369 80 83370
rect 42 83328 76 83362
rect 79 83328 113 83362
rect 42 83249 46 83283
rect 72 83249 76 83283
rect -25 83212 25 83214
rect -8 83204 14 83211
rect -8 83203 17 83204
rect 25 83203 27 83212
rect -12 83196 38 83203
rect -12 83195 34 83196
rect -12 83191 8 83195
rect 0 83179 8 83191
rect 14 83179 34 83195
rect 0 83178 34 83179
rect 0 83171 38 83178
rect 14 83170 17 83171
rect 25 83162 27 83171
rect 42 83142 45 83232
rect 71 83201 80 83229
rect 69 83163 80 83201
rect 144 83191 148 83499
rect 196 83486 204 83520
rect 216 83486 232 83520
rect 244 83516 257 83520
rect 300 83516 308 83529
rect 332 83527 342 83565
rect 400 83557 404 83565
rect 336 83517 342 83527
rect 244 83492 291 83516
rect 244 83486 257 83492
rect 224 83439 226 83486
rect 278 83482 291 83492
rect 300 83492 329 83516
rect 332 83507 342 83517
rect 400 83517 409 83545
rect 562 83528 612 83530
rect 466 83519 497 83527
rect 565 83519 596 83527
rect 300 83482 321 83492
rect 300 83476 308 83482
rect 289 83466 308 83476
rect 196 83409 204 83439
rect 216 83409 232 83439
rect 196 83405 232 83409
rect 196 83397 226 83405
rect 300 83397 308 83466
rect 332 83473 351 83507
rect 361 83479 381 83507
rect 361 83473 375 83479
rect 400 83473 411 83517
rect 442 83512 500 83519
rect 466 83511 500 83512
rect 565 83511 599 83519
rect 497 83495 500 83511
rect 596 83495 599 83511
rect 466 83494 500 83495
rect 442 83487 500 83494
rect 565 83487 599 83495
rect 612 83478 614 83528
rect 332 83449 342 83473
rect 336 83437 342 83449
rect 224 83381 226 83397
rect 332 83369 342 83437
rect 400 83441 404 83449
rect 400 83407 408 83441
rect 434 83407 438 83441
rect 454 83425 504 83427
rect 504 83409 506 83425
rect 514 83419 530 83425
rect 532 83419 548 83425
rect 525 83409 548 83418
rect 400 83399 404 83407
rect 498 83399 506 83409
rect 504 83375 506 83399
rect 514 83389 515 83409
rect 525 83384 528 83409
rect 547 83389 548 83409
rect 557 83399 564 83409
rect 514 83375 548 83379
rect 151 83328 156 83362
rect 174 83359 246 83367
rect 256 83359 328 83367
rect 336 83361 342 83369
rect 400 83364 404 83369
rect 180 83331 185 83359
rect 174 83323 246 83331
rect 256 83323 328 83331
rect 332 83329 336 83359
rect 400 83330 438 83364
rect 224 83293 226 83309
rect 196 83285 226 83293
rect 196 83281 232 83285
rect 196 83251 204 83281
rect 216 83251 232 83281
rect 224 83204 226 83251
rect 300 83224 308 83293
rect 332 83291 342 83329
rect 400 83321 404 83330
rect 454 83315 504 83317
rect 494 83311 548 83315
rect 494 83306 514 83311
rect 504 83291 506 83306
rect 336 83279 342 83291
rect 289 83214 308 83224
rect 300 83208 308 83214
rect 332 83245 342 83279
rect 400 83283 404 83291
rect 400 83249 408 83283
rect 434 83249 438 83283
rect 498 83281 506 83291
rect 514 83281 515 83301
rect 504 83265 506 83281
rect 525 83272 528 83306
rect 547 83281 548 83301
rect 557 83281 564 83291
rect 514 83265 530 83271
rect 532 83265 548 83271
rect 332 83217 373 83245
rect 332 83211 351 83217
rect 107 83157 119 83191
rect 129 83157 149 83191
rect 196 83170 204 83204
rect 216 83170 232 83204
rect 244 83198 257 83204
rect 278 83198 291 83208
rect 244 83174 291 83198
rect 300 83198 321 83208
rect 336 83201 351 83211
rect 300 83174 329 83198
rect 332 83183 351 83201
rect 361 83211 375 83217
rect 400 83211 411 83249
rect 562 83212 612 83214
rect 361 83183 381 83211
rect 400 83183 409 83211
rect 466 83203 497 83211
rect 565 83203 596 83211
rect 442 83196 500 83203
rect 466 83195 500 83196
rect 565 83195 599 83203
rect 244 83170 257 83174
rect 42 83091 46 83125
rect 72 83091 76 83125
rect 42 83044 76 83048
rect 42 83029 46 83044
rect 72 83029 76 83044
rect 38 83011 80 83029
rect 16 83005 102 83011
rect 144 83005 148 83157
rect 174 83133 181 83161
rect 224 83123 226 83170
rect 300 83161 308 83174
rect 278 83150 305 83161
rect 332 83133 342 83183
rect 400 83163 404 83183
rect 497 83179 500 83195
rect 596 83179 599 83195
rect 466 83178 500 83179
rect 442 83171 500 83178
rect 565 83171 599 83179
rect 612 83162 614 83212
rect 256 83123 328 83131
rect 336 83125 342 83133
rect 400 83125 404 83133
rect 196 83093 204 83123
rect 216 83093 232 83123
rect 196 83089 232 83093
rect 196 83081 226 83089
rect 224 83065 226 83081
rect 332 83053 336 83121
rect 400 83091 408 83125
rect 434 83091 438 83125
rect 454 83109 504 83111
rect 504 83093 506 83109
rect 514 83103 530 83109
rect 532 83103 548 83109
rect 525 83093 548 83102
rect 400 83083 404 83091
rect 498 83083 506 83093
rect 504 83059 506 83083
rect 514 83073 515 83093
rect 525 83068 528 83093
rect 547 83073 548 83093
rect 557 83083 564 83093
rect 514 83059 548 83063
rect 400 83053 442 83054
rect 174 83043 246 83051
rect 400 83046 404 83053
rect 295 83012 300 83046
rect 324 83012 329 83046
rect 367 83029 438 83046
rect 367 83012 442 83029
rect 400 83011 442 83012
rect 378 83005 464 83011
rect 38 82989 80 83005
rect 400 82989 442 83005
rect -25 82975 25 82977
rect 42 82975 76 82989
rect 404 82975 438 82989
rect 455 82975 505 82977
rect 557 82975 607 82977
rect 16 82967 102 82975
rect 378 82967 464 82975
rect 8 82933 17 82967
rect 18 82965 51 82967
rect 80 82965 100 82967
rect 18 82933 100 82965
rect 380 82965 404 82967
rect 429 82965 438 82967
rect 442 82965 462 82967
rect 16 82925 102 82933
rect 42 82909 76 82925
rect 16 82889 38 82895
rect 42 82886 76 82890
rect 80 82889 102 82895
rect 42 82856 46 82886
rect 72 82856 76 82886
rect 42 82775 46 82809
rect 72 82775 76 82809
rect -25 82738 25 82740
rect -8 82730 14 82737
rect -8 82729 17 82730
rect 25 82729 27 82738
rect -12 82722 38 82729
rect -12 82721 34 82722
rect -12 82717 8 82721
rect 0 82705 8 82717
rect 14 82705 34 82721
rect 0 82704 34 82705
rect 0 82697 38 82704
rect 14 82696 17 82697
rect 25 82688 27 82697
rect 42 82668 45 82758
rect 69 82743 80 82775
rect 107 82743 143 82771
rect 144 82743 148 82963
rect 332 82895 336 82963
rect 380 82933 462 82965
rect 463 82933 472 82967
rect 480 82933 497 82967
rect 378 82925 464 82933
rect 505 82925 507 82975
rect 514 82933 548 82967
rect 565 82933 582 82967
rect 607 82925 609 82975
rect 404 82909 438 82925
rect 400 82895 442 82896
rect 378 82889 404 82895
rect 442 82889 464 82895
rect 400 82888 404 82889
rect 174 82849 246 82857
rect 295 82854 300 82888
rect 324 82854 329 82888
rect 224 82819 226 82835
rect 196 82811 226 82819
rect 332 82817 336 82885
rect 367 82854 438 82888
rect 400 82847 404 82854
rect 454 82841 504 82843
rect 494 82837 548 82841
rect 494 82832 514 82837
rect 504 82817 506 82832
rect 196 82807 232 82811
rect 196 82777 204 82807
rect 216 82777 232 82807
rect 400 82809 404 82817
rect 107 82737 119 82743
rect 109 82709 119 82737
rect 129 82709 149 82743
rect 174 82739 181 82769
rect 224 82730 226 82777
rect 256 82769 328 82777
rect 332 82775 336 82805
rect 400 82775 408 82809
rect 434 82775 438 82809
rect 498 82807 506 82817
rect 514 82807 515 82827
rect 504 82791 506 82807
rect 525 82798 528 82832
rect 547 82807 548 82827
rect 557 82807 564 82817
rect 514 82791 530 82797
rect 532 82791 548 82797
rect 278 82739 305 82750
rect 42 82617 46 82651
rect 72 82617 76 82651
rect 38 82579 80 82580
rect 42 82538 76 82572
rect 79 82538 113 82572
rect 42 82459 46 82493
rect 72 82459 76 82493
rect -25 82422 25 82424
rect -8 82414 14 82421
rect -8 82413 17 82414
rect 25 82413 27 82422
rect -12 82406 38 82413
rect -12 82405 34 82406
rect -12 82401 8 82405
rect 0 82389 8 82401
rect 14 82389 34 82405
rect 0 82388 34 82389
rect 0 82381 38 82388
rect 14 82380 17 82381
rect 25 82372 27 82381
rect 42 82352 45 82442
rect 71 82411 80 82439
rect 69 82373 80 82411
rect 144 82401 148 82709
rect 196 82696 204 82730
rect 216 82696 232 82730
rect 244 82726 257 82730
rect 300 82726 308 82739
rect 332 82737 342 82775
rect 400 82767 404 82775
rect 336 82727 342 82737
rect 244 82702 291 82726
rect 244 82696 257 82702
rect 224 82649 226 82696
rect 278 82692 291 82702
rect 300 82702 329 82726
rect 332 82717 342 82727
rect 400 82727 409 82755
rect 562 82738 612 82740
rect 466 82729 497 82737
rect 565 82729 596 82737
rect 300 82692 321 82702
rect 300 82686 308 82692
rect 289 82676 308 82686
rect 196 82619 204 82649
rect 216 82619 232 82649
rect 196 82615 232 82619
rect 196 82607 226 82615
rect 300 82607 308 82676
rect 332 82683 351 82717
rect 361 82689 381 82717
rect 361 82683 375 82689
rect 400 82683 411 82727
rect 442 82722 500 82729
rect 466 82721 500 82722
rect 565 82721 599 82729
rect 497 82705 500 82721
rect 596 82705 599 82721
rect 466 82704 500 82705
rect 442 82697 500 82704
rect 565 82697 599 82705
rect 612 82688 614 82738
rect 332 82659 342 82683
rect 336 82647 342 82659
rect 224 82591 226 82607
rect 332 82579 342 82647
rect 400 82651 404 82659
rect 400 82617 408 82651
rect 434 82617 438 82651
rect 454 82635 504 82637
rect 504 82619 506 82635
rect 514 82629 530 82635
rect 532 82629 548 82635
rect 525 82619 548 82628
rect 400 82609 404 82617
rect 498 82609 506 82619
rect 504 82585 506 82609
rect 514 82599 515 82619
rect 525 82594 528 82619
rect 547 82599 548 82619
rect 557 82609 564 82619
rect 514 82585 548 82589
rect 151 82538 156 82572
rect 174 82569 246 82577
rect 256 82569 328 82577
rect 336 82571 342 82579
rect 400 82574 404 82579
rect 180 82541 185 82569
rect 174 82533 246 82541
rect 256 82533 328 82541
rect 332 82539 336 82569
rect 400 82540 438 82574
rect 224 82503 226 82519
rect 196 82495 226 82503
rect 196 82491 232 82495
rect 196 82461 204 82491
rect 216 82461 232 82491
rect 224 82414 226 82461
rect 300 82434 308 82503
rect 332 82501 342 82539
rect 400 82531 404 82540
rect 454 82525 504 82527
rect 494 82521 548 82525
rect 494 82516 514 82521
rect 504 82501 506 82516
rect 336 82489 342 82501
rect 289 82424 308 82434
rect 300 82418 308 82424
rect 332 82455 342 82489
rect 400 82493 404 82501
rect 400 82459 408 82493
rect 434 82459 438 82493
rect 498 82491 506 82501
rect 514 82491 515 82511
rect 504 82475 506 82491
rect 525 82482 528 82516
rect 547 82491 548 82511
rect 557 82491 564 82501
rect 514 82475 530 82481
rect 532 82475 548 82481
rect 332 82427 373 82455
rect 332 82421 351 82427
rect 107 82367 119 82401
rect 129 82367 149 82401
rect 196 82380 204 82414
rect 216 82380 232 82414
rect 244 82408 257 82414
rect 278 82408 291 82418
rect 244 82384 291 82408
rect 300 82408 321 82418
rect 336 82411 351 82421
rect 300 82384 329 82408
rect 332 82393 351 82411
rect 361 82421 375 82427
rect 400 82421 411 82459
rect 562 82422 612 82424
rect 361 82393 381 82421
rect 400 82393 409 82421
rect 466 82413 497 82421
rect 565 82413 596 82421
rect 442 82406 500 82413
rect 466 82405 500 82406
rect 565 82405 599 82413
rect 244 82380 257 82384
rect 42 82301 46 82335
rect 72 82301 76 82335
rect 42 82254 76 82258
rect 42 82239 46 82254
rect 72 82239 76 82254
rect 38 82221 80 82239
rect 16 82215 102 82221
rect 144 82215 148 82367
rect 174 82343 181 82371
rect 224 82333 226 82380
rect 300 82371 308 82384
rect 278 82360 305 82371
rect 332 82343 342 82393
rect 400 82373 404 82393
rect 497 82389 500 82405
rect 596 82389 599 82405
rect 466 82388 500 82389
rect 442 82381 500 82388
rect 565 82381 599 82389
rect 612 82372 614 82422
rect 256 82333 328 82341
rect 336 82335 342 82343
rect 400 82335 404 82343
rect 196 82303 204 82333
rect 216 82303 232 82333
rect 196 82299 232 82303
rect 196 82291 226 82299
rect 224 82275 226 82291
rect 332 82263 336 82331
rect 400 82301 408 82335
rect 434 82301 438 82335
rect 454 82319 504 82321
rect 504 82303 506 82319
rect 514 82313 530 82319
rect 532 82313 548 82319
rect 525 82303 548 82312
rect 400 82293 404 82301
rect 498 82293 506 82303
rect 504 82269 506 82293
rect 514 82283 515 82303
rect 525 82278 528 82303
rect 547 82283 548 82303
rect 557 82293 564 82303
rect 514 82269 548 82273
rect 400 82263 442 82264
rect 174 82253 246 82261
rect 400 82256 404 82263
rect 295 82222 300 82256
rect 324 82222 329 82256
rect 367 82239 438 82256
rect 367 82222 442 82239
rect 400 82221 442 82222
rect 378 82215 464 82221
rect 38 82199 80 82215
rect 400 82199 442 82215
rect -25 82185 25 82187
rect 42 82185 76 82199
rect 404 82185 438 82199
rect 455 82185 505 82187
rect 557 82185 607 82187
rect 16 82177 102 82185
rect 378 82177 464 82185
rect 8 82143 17 82177
rect 18 82175 51 82177
rect 80 82175 100 82177
rect 18 82143 100 82175
rect 380 82175 404 82177
rect 429 82175 438 82177
rect 442 82175 462 82177
rect 16 82135 102 82143
rect 42 82119 76 82135
rect 16 82099 38 82105
rect 42 82096 76 82100
rect 80 82099 102 82105
rect 42 82066 46 82096
rect 72 82066 76 82096
rect 42 81985 46 82019
rect 72 81985 76 82019
rect -25 81948 25 81950
rect -8 81940 14 81947
rect -8 81939 17 81940
rect 25 81939 27 81948
rect -12 81932 38 81939
rect -12 81931 34 81932
rect -12 81927 8 81931
rect 0 81915 8 81927
rect 14 81915 34 81931
rect 0 81914 34 81915
rect 0 81907 38 81914
rect 14 81906 17 81907
rect 25 81898 27 81907
rect 42 81878 45 81968
rect 69 81953 80 81985
rect 107 81953 143 81981
rect 144 81953 148 82173
rect 332 82105 336 82173
rect 380 82143 462 82175
rect 463 82143 472 82177
rect 480 82143 497 82177
rect 378 82135 464 82143
rect 505 82135 507 82185
rect 514 82143 548 82177
rect 565 82143 582 82177
rect 607 82135 609 82185
rect 404 82119 438 82135
rect 400 82105 442 82106
rect 378 82099 404 82105
rect 442 82099 464 82105
rect 400 82098 404 82099
rect 174 82059 246 82067
rect 295 82064 300 82098
rect 324 82064 329 82098
rect 224 82029 226 82045
rect 196 82021 226 82029
rect 332 82027 336 82095
rect 367 82064 438 82098
rect 400 82057 404 82064
rect 454 82051 504 82053
rect 494 82047 548 82051
rect 494 82042 514 82047
rect 504 82027 506 82042
rect 196 82017 232 82021
rect 196 81987 204 82017
rect 216 81987 232 82017
rect 400 82019 404 82027
rect 107 81947 119 81953
rect 109 81919 119 81947
rect 129 81919 149 81953
rect 174 81949 181 81979
rect 224 81940 226 81987
rect 256 81979 328 81987
rect 332 81985 336 82015
rect 400 81985 408 82019
rect 434 81985 438 82019
rect 498 82017 506 82027
rect 514 82017 515 82037
rect 504 82001 506 82017
rect 525 82008 528 82042
rect 547 82017 548 82037
rect 557 82017 564 82027
rect 514 82001 530 82007
rect 532 82001 548 82007
rect 278 81949 305 81960
rect 42 81827 46 81861
rect 72 81827 76 81861
rect 38 81789 80 81790
rect 42 81748 76 81782
rect 79 81748 113 81782
rect 42 81669 46 81703
rect 72 81669 76 81703
rect -25 81632 25 81634
rect -8 81624 14 81631
rect -8 81623 17 81624
rect 25 81623 27 81632
rect -12 81616 38 81623
rect -12 81615 34 81616
rect -12 81611 8 81615
rect 0 81599 8 81611
rect 14 81599 34 81615
rect 0 81598 34 81599
rect 0 81591 38 81598
rect 14 81590 17 81591
rect 25 81582 27 81591
rect 42 81562 45 81652
rect 71 81621 80 81649
rect 69 81583 80 81621
rect 144 81611 148 81919
rect 196 81906 204 81940
rect 216 81906 232 81940
rect 244 81936 257 81940
rect 300 81936 308 81949
rect 332 81947 342 81985
rect 400 81977 404 81985
rect 336 81937 342 81947
rect 244 81912 291 81936
rect 244 81906 257 81912
rect 224 81859 226 81906
rect 278 81902 291 81912
rect 300 81912 329 81936
rect 332 81927 342 81937
rect 400 81937 409 81965
rect 562 81948 612 81950
rect 466 81939 497 81947
rect 565 81939 596 81947
rect 300 81902 321 81912
rect 300 81896 308 81902
rect 289 81886 308 81896
rect 196 81829 204 81859
rect 216 81829 232 81859
rect 196 81825 232 81829
rect 196 81817 226 81825
rect 300 81817 308 81886
rect 332 81893 351 81927
rect 361 81899 381 81927
rect 361 81893 375 81899
rect 400 81893 411 81937
rect 442 81932 500 81939
rect 466 81931 500 81932
rect 565 81931 599 81939
rect 497 81915 500 81931
rect 596 81915 599 81931
rect 466 81914 500 81915
rect 442 81907 500 81914
rect 565 81907 599 81915
rect 612 81898 614 81948
rect 332 81869 342 81893
rect 336 81857 342 81869
rect 224 81801 226 81817
rect 332 81789 342 81857
rect 400 81861 404 81869
rect 400 81827 408 81861
rect 434 81827 438 81861
rect 454 81845 504 81847
rect 504 81829 506 81845
rect 514 81839 530 81845
rect 532 81839 548 81845
rect 525 81829 548 81838
rect 400 81819 404 81827
rect 498 81819 506 81829
rect 504 81795 506 81819
rect 514 81809 515 81829
rect 525 81804 528 81829
rect 547 81809 548 81829
rect 557 81819 564 81829
rect 514 81795 548 81799
rect 151 81748 156 81782
rect 174 81779 246 81787
rect 256 81779 328 81787
rect 336 81781 342 81789
rect 400 81784 404 81789
rect 180 81751 185 81779
rect 174 81743 246 81751
rect 256 81743 328 81751
rect 332 81749 336 81779
rect 400 81750 438 81784
rect 224 81713 226 81729
rect 196 81705 226 81713
rect 196 81701 232 81705
rect 196 81671 204 81701
rect 216 81671 232 81701
rect 224 81624 226 81671
rect 300 81644 308 81713
rect 332 81711 342 81749
rect 400 81741 404 81750
rect 454 81735 504 81737
rect 494 81731 548 81735
rect 494 81726 514 81731
rect 504 81711 506 81726
rect 336 81699 342 81711
rect 289 81634 308 81644
rect 300 81628 308 81634
rect 332 81665 342 81699
rect 400 81703 404 81711
rect 400 81669 408 81703
rect 434 81669 438 81703
rect 498 81701 506 81711
rect 514 81701 515 81721
rect 504 81685 506 81701
rect 525 81692 528 81726
rect 547 81701 548 81721
rect 557 81701 564 81711
rect 514 81685 530 81691
rect 532 81685 548 81691
rect 332 81637 373 81665
rect 332 81631 351 81637
rect 107 81577 119 81611
rect 129 81577 149 81611
rect 196 81590 204 81624
rect 216 81590 232 81624
rect 244 81618 257 81624
rect 278 81618 291 81628
rect 244 81594 291 81618
rect 300 81618 321 81628
rect 336 81621 351 81631
rect 300 81594 329 81618
rect 332 81603 351 81621
rect 361 81631 375 81637
rect 400 81631 411 81669
rect 562 81632 612 81634
rect 361 81603 381 81631
rect 400 81603 409 81631
rect 466 81623 497 81631
rect 565 81623 596 81631
rect 442 81616 500 81623
rect 466 81615 500 81616
rect 565 81615 599 81623
rect 244 81590 257 81594
rect 42 81511 46 81545
rect 72 81511 76 81545
rect 42 81464 76 81468
rect 42 81449 46 81464
rect 72 81449 76 81464
rect 38 81431 80 81449
rect 16 81425 102 81431
rect 144 81425 148 81577
rect 174 81553 181 81581
rect 224 81543 226 81590
rect 300 81581 308 81594
rect 278 81570 305 81581
rect 332 81553 342 81603
rect 400 81583 404 81603
rect 497 81599 500 81615
rect 596 81599 599 81615
rect 466 81598 500 81599
rect 442 81591 500 81598
rect 565 81591 599 81599
rect 612 81582 614 81632
rect 256 81543 328 81551
rect 336 81545 342 81553
rect 400 81545 404 81553
rect 196 81513 204 81543
rect 216 81513 232 81543
rect 196 81509 232 81513
rect 196 81501 226 81509
rect 224 81485 226 81501
rect 332 81473 336 81541
rect 400 81511 408 81545
rect 434 81511 438 81545
rect 454 81529 504 81531
rect 504 81513 506 81529
rect 514 81523 530 81529
rect 532 81523 548 81529
rect 525 81513 548 81522
rect 400 81503 404 81511
rect 498 81503 506 81513
rect 504 81479 506 81503
rect 514 81493 515 81513
rect 525 81488 528 81513
rect 547 81493 548 81513
rect 557 81503 564 81513
rect 514 81479 548 81483
rect 400 81473 442 81474
rect 174 81463 246 81471
rect 400 81466 404 81473
rect 295 81432 300 81466
rect 324 81432 329 81466
rect 367 81449 438 81466
rect 367 81432 442 81449
rect 400 81431 442 81432
rect 378 81425 464 81431
rect 38 81409 80 81425
rect 400 81409 442 81425
rect -25 81395 25 81397
rect 42 81395 76 81409
rect 404 81395 438 81409
rect 455 81395 505 81397
rect 557 81395 607 81397
rect 16 81387 102 81395
rect 378 81387 464 81395
rect 8 81353 17 81387
rect 18 81385 51 81387
rect 80 81385 100 81387
rect 18 81353 100 81385
rect 380 81385 404 81387
rect 429 81385 438 81387
rect 442 81385 462 81387
rect 16 81345 102 81353
rect 42 81329 76 81345
rect 16 81309 38 81315
rect 42 81306 76 81310
rect 80 81309 102 81315
rect 42 81276 46 81306
rect 72 81276 76 81306
rect 42 81195 46 81229
rect 72 81195 76 81229
rect -25 81158 25 81160
rect -8 81150 14 81157
rect -8 81149 17 81150
rect 25 81149 27 81158
rect -12 81142 38 81149
rect -12 81141 34 81142
rect -12 81137 8 81141
rect 0 81125 8 81137
rect 14 81125 34 81141
rect 0 81124 34 81125
rect 0 81117 38 81124
rect 14 81116 17 81117
rect 25 81108 27 81117
rect 42 81088 45 81178
rect 69 81163 80 81195
rect 107 81163 143 81191
rect 144 81163 148 81383
rect 332 81315 336 81383
rect 380 81353 462 81385
rect 463 81353 472 81387
rect 480 81353 497 81387
rect 378 81345 464 81353
rect 505 81345 507 81395
rect 514 81353 548 81387
rect 565 81353 582 81387
rect 607 81345 609 81395
rect 404 81329 438 81345
rect 400 81315 442 81316
rect 378 81309 404 81315
rect 442 81309 464 81315
rect 400 81308 404 81309
rect 174 81269 246 81277
rect 295 81274 300 81308
rect 324 81274 329 81308
rect 224 81239 226 81255
rect 196 81231 226 81239
rect 332 81237 336 81305
rect 367 81274 438 81308
rect 400 81267 404 81274
rect 454 81261 504 81263
rect 494 81257 548 81261
rect 494 81252 514 81257
rect 504 81237 506 81252
rect 196 81227 232 81231
rect 196 81197 204 81227
rect 216 81197 232 81227
rect 400 81229 404 81237
rect 107 81157 119 81163
rect 109 81129 119 81157
rect 129 81129 149 81163
rect 174 81159 181 81189
rect 224 81150 226 81197
rect 256 81189 328 81197
rect 332 81195 336 81225
rect 400 81195 408 81229
rect 434 81195 438 81229
rect 498 81227 506 81237
rect 514 81227 515 81247
rect 504 81211 506 81227
rect 525 81218 528 81252
rect 547 81227 548 81247
rect 557 81227 564 81237
rect 514 81211 530 81217
rect 532 81211 548 81217
rect 278 81159 305 81170
rect 42 81037 46 81071
rect 72 81037 76 81071
rect 38 80999 80 81000
rect 42 80958 76 80992
rect 79 80958 113 80992
rect 42 80879 46 80913
rect 72 80879 76 80913
rect -25 80842 25 80844
rect -8 80834 14 80841
rect -8 80833 17 80834
rect 25 80833 27 80842
rect -12 80826 38 80833
rect -12 80825 34 80826
rect -12 80821 8 80825
rect 0 80809 8 80821
rect 14 80809 34 80825
rect 0 80808 34 80809
rect 0 80801 38 80808
rect 14 80800 17 80801
rect 25 80792 27 80801
rect 42 80772 45 80862
rect 71 80831 80 80859
rect 69 80793 80 80831
rect 144 80821 148 81129
rect 196 81116 204 81150
rect 216 81116 232 81150
rect 244 81146 257 81150
rect 300 81146 308 81159
rect 332 81157 342 81195
rect 400 81187 404 81195
rect 336 81147 342 81157
rect 244 81122 291 81146
rect 244 81116 257 81122
rect 224 81069 226 81116
rect 278 81112 291 81122
rect 300 81122 329 81146
rect 332 81137 342 81147
rect 400 81147 409 81175
rect 562 81158 612 81160
rect 466 81149 497 81157
rect 565 81149 596 81157
rect 300 81112 321 81122
rect 300 81106 308 81112
rect 289 81096 308 81106
rect 196 81039 204 81069
rect 216 81039 232 81069
rect 196 81035 232 81039
rect 196 81027 226 81035
rect 300 81027 308 81096
rect 332 81103 351 81137
rect 361 81109 381 81137
rect 361 81103 375 81109
rect 400 81103 411 81147
rect 442 81142 500 81149
rect 466 81141 500 81142
rect 565 81141 599 81149
rect 497 81125 500 81141
rect 596 81125 599 81141
rect 466 81124 500 81125
rect 442 81117 500 81124
rect 565 81117 599 81125
rect 612 81108 614 81158
rect 332 81079 342 81103
rect 336 81067 342 81079
rect 224 81011 226 81027
rect 332 80999 342 81067
rect 400 81071 404 81079
rect 400 81037 408 81071
rect 434 81037 438 81071
rect 454 81055 504 81057
rect 504 81039 506 81055
rect 514 81049 530 81055
rect 532 81049 548 81055
rect 525 81039 548 81048
rect 400 81029 404 81037
rect 498 81029 506 81039
rect 504 81005 506 81029
rect 514 81019 515 81039
rect 525 81014 528 81039
rect 547 81019 548 81039
rect 557 81029 564 81039
rect 514 81005 548 81009
rect 151 80958 156 80992
rect 174 80989 246 80997
rect 256 80989 328 80997
rect 336 80991 342 80999
rect 400 80994 404 80999
rect 180 80961 185 80989
rect 174 80953 246 80961
rect 256 80953 328 80961
rect 332 80959 336 80989
rect 400 80960 438 80994
rect 224 80923 226 80939
rect 196 80915 226 80923
rect 196 80911 232 80915
rect 196 80881 204 80911
rect 216 80881 232 80911
rect 224 80834 226 80881
rect 300 80854 308 80923
rect 332 80921 342 80959
rect 400 80951 404 80960
rect 454 80945 504 80947
rect 494 80941 548 80945
rect 494 80936 514 80941
rect 504 80921 506 80936
rect 336 80909 342 80921
rect 289 80844 308 80854
rect 300 80838 308 80844
rect 332 80875 342 80909
rect 400 80913 404 80921
rect 400 80879 408 80913
rect 434 80879 438 80913
rect 498 80911 506 80921
rect 514 80911 515 80931
rect 504 80895 506 80911
rect 525 80902 528 80936
rect 547 80911 548 80931
rect 557 80911 564 80921
rect 514 80895 530 80901
rect 532 80895 548 80901
rect 332 80847 373 80875
rect 332 80841 351 80847
rect 107 80787 119 80821
rect 129 80787 149 80821
rect 196 80800 204 80834
rect 216 80800 232 80834
rect 244 80828 257 80834
rect 278 80828 291 80838
rect 244 80804 291 80828
rect 300 80828 321 80838
rect 336 80831 351 80841
rect 300 80804 329 80828
rect 332 80813 351 80831
rect 361 80841 375 80847
rect 400 80841 411 80879
rect 562 80842 612 80844
rect 361 80813 381 80841
rect 400 80813 409 80841
rect 466 80833 497 80841
rect 565 80833 596 80841
rect 442 80826 500 80833
rect 466 80825 500 80826
rect 565 80825 599 80833
rect 244 80800 257 80804
rect 42 80721 46 80755
rect 72 80721 76 80755
rect 42 80674 76 80678
rect 42 80659 46 80674
rect 72 80659 76 80674
rect 38 80641 80 80659
rect 16 80635 102 80641
rect 144 80635 148 80787
rect 174 80763 181 80791
rect 224 80753 226 80800
rect 300 80791 308 80804
rect 278 80780 305 80791
rect 332 80763 342 80813
rect 400 80793 404 80813
rect 497 80809 500 80825
rect 596 80809 599 80825
rect 466 80808 500 80809
rect 442 80801 500 80808
rect 565 80801 599 80809
rect 612 80792 614 80842
rect 256 80753 328 80761
rect 336 80755 342 80763
rect 400 80755 404 80763
rect 196 80723 204 80753
rect 216 80723 232 80753
rect 196 80719 232 80723
rect 196 80711 226 80719
rect 224 80695 226 80711
rect 332 80683 336 80751
rect 400 80721 408 80755
rect 434 80721 438 80755
rect 454 80739 504 80741
rect 504 80723 506 80739
rect 514 80733 530 80739
rect 532 80733 548 80739
rect 525 80723 548 80732
rect 400 80713 404 80721
rect 498 80713 506 80723
rect 504 80689 506 80713
rect 514 80703 515 80723
rect 525 80698 528 80723
rect 547 80703 548 80723
rect 557 80713 564 80723
rect 514 80689 548 80693
rect 400 80683 442 80684
rect 174 80673 246 80681
rect 400 80676 404 80683
rect 295 80642 300 80676
rect 324 80642 329 80676
rect 367 80659 438 80676
rect 367 80642 442 80659
rect 400 80641 442 80642
rect 378 80635 464 80641
rect 38 80619 80 80635
rect 400 80619 442 80635
rect -25 80605 25 80607
rect 42 80605 76 80619
rect 404 80605 438 80619
rect 455 80605 505 80607
rect 557 80605 607 80607
rect 16 80597 102 80605
rect 378 80597 464 80605
rect 8 80563 17 80597
rect 18 80595 51 80597
rect 80 80595 100 80597
rect 18 80563 100 80595
rect 380 80595 404 80597
rect 429 80595 438 80597
rect 442 80595 462 80597
rect 16 80555 102 80563
rect 42 80539 76 80555
rect 16 80519 38 80525
rect 42 80516 76 80520
rect 80 80519 102 80525
rect 42 80486 46 80516
rect 72 80486 76 80516
rect 42 80405 46 80439
rect 72 80405 76 80439
rect -25 80368 25 80370
rect -8 80360 14 80367
rect -8 80359 17 80360
rect 25 80359 27 80368
rect -12 80352 38 80359
rect -12 80351 34 80352
rect -12 80347 8 80351
rect 0 80335 8 80347
rect 14 80335 34 80351
rect 0 80334 34 80335
rect 0 80327 38 80334
rect 14 80326 17 80327
rect 25 80318 27 80327
rect 42 80298 45 80388
rect 69 80373 80 80405
rect 107 80373 143 80401
rect 144 80373 148 80593
rect 332 80525 336 80593
rect 380 80563 462 80595
rect 463 80563 472 80597
rect 480 80563 497 80597
rect 378 80555 464 80563
rect 505 80555 507 80605
rect 514 80563 548 80597
rect 565 80563 582 80597
rect 607 80555 609 80605
rect 404 80539 438 80555
rect 400 80525 442 80526
rect 378 80519 404 80525
rect 442 80519 464 80525
rect 400 80518 404 80519
rect 174 80479 246 80487
rect 295 80484 300 80518
rect 324 80484 329 80518
rect 224 80449 226 80465
rect 196 80441 226 80449
rect 332 80447 336 80515
rect 367 80484 438 80518
rect 400 80477 404 80484
rect 454 80471 504 80473
rect 494 80467 548 80471
rect 494 80462 514 80467
rect 504 80447 506 80462
rect 196 80437 232 80441
rect 196 80407 204 80437
rect 216 80407 232 80437
rect 400 80439 404 80447
rect 107 80367 119 80373
rect 109 80339 119 80367
rect 129 80339 149 80373
rect 174 80369 181 80399
rect 224 80360 226 80407
rect 256 80399 328 80407
rect 332 80405 336 80435
rect 400 80405 408 80439
rect 434 80405 438 80439
rect 498 80437 506 80447
rect 514 80437 515 80457
rect 504 80421 506 80437
rect 525 80428 528 80462
rect 547 80437 548 80457
rect 557 80437 564 80447
rect 514 80421 530 80427
rect 532 80421 548 80427
rect 278 80369 305 80380
rect 42 80247 46 80281
rect 72 80247 76 80281
rect 38 80209 80 80210
rect 42 80168 76 80202
rect 79 80168 113 80202
rect 42 80089 46 80123
rect 72 80089 76 80123
rect -25 80052 25 80054
rect -8 80044 14 80051
rect -8 80043 17 80044
rect 25 80043 27 80052
rect -12 80036 38 80043
rect -12 80035 34 80036
rect -12 80031 8 80035
rect 0 80019 8 80031
rect 14 80019 34 80035
rect 0 80018 34 80019
rect 0 80011 38 80018
rect 14 80010 17 80011
rect 25 80002 27 80011
rect 42 79982 45 80072
rect 71 80041 80 80069
rect 69 80003 80 80041
rect 144 80031 148 80339
rect 196 80326 204 80360
rect 216 80326 232 80360
rect 244 80356 257 80360
rect 300 80356 308 80369
rect 332 80367 342 80405
rect 400 80397 404 80405
rect 336 80357 342 80367
rect 244 80332 291 80356
rect 244 80326 257 80332
rect 224 80279 226 80326
rect 278 80322 291 80332
rect 300 80332 329 80356
rect 332 80347 342 80357
rect 400 80357 409 80385
rect 562 80368 612 80370
rect 466 80359 497 80367
rect 565 80359 596 80367
rect 300 80322 321 80332
rect 300 80316 308 80322
rect 289 80306 308 80316
rect 196 80249 204 80279
rect 216 80249 232 80279
rect 196 80245 232 80249
rect 196 80237 226 80245
rect 300 80237 308 80306
rect 332 80313 351 80347
rect 361 80319 381 80347
rect 361 80313 375 80319
rect 400 80313 411 80357
rect 442 80352 500 80359
rect 466 80351 500 80352
rect 565 80351 599 80359
rect 497 80335 500 80351
rect 596 80335 599 80351
rect 466 80334 500 80335
rect 442 80327 500 80334
rect 565 80327 599 80335
rect 612 80318 614 80368
rect 332 80289 342 80313
rect 336 80277 342 80289
rect 224 80221 226 80237
rect 332 80209 342 80277
rect 400 80281 404 80289
rect 400 80247 408 80281
rect 434 80247 438 80281
rect 454 80265 504 80267
rect 504 80249 506 80265
rect 514 80259 530 80265
rect 532 80259 548 80265
rect 525 80249 548 80258
rect 400 80239 404 80247
rect 498 80239 506 80249
rect 504 80215 506 80239
rect 514 80229 515 80249
rect 525 80224 528 80249
rect 547 80229 548 80249
rect 557 80239 564 80249
rect 514 80215 548 80219
rect 151 80168 156 80202
rect 174 80199 246 80207
rect 256 80199 328 80207
rect 336 80201 342 80209
rect 400 80204 404 80209
rect 180 80171 185 80199
rect 174 80163 246 80171
rect 256 80163 328 80171
rect 332 80169 336 80199
rect 400 80170 438 80204
rect 224 80133 226 80149
rect 196 80125 226 80133
rect 196 80121 232 80125
rect 196 80091 204 80121
rect 216 80091 232 80121
rect 224 80044 226 80091
rect 300 80064 308 80133
rect 332 80131 342 80169
rect 400 80161 404 80170
rect 454 80155 504 80157
rect 494 80151 548 80155
rect 494 80146 514 80151
rect 504 80131 506 80146
rect 336 80119 342 80131
rect 289 80054 308 80064
rect 300 80048 308 80054
rect 332 80085 342 80119
rect 400 80123 404 80131
rect 400 80089 408 80123
rect 434 80089 438 80123
rect 498 80121 506 80131
rect 514 80121 515 80141
rect 504 80105 506 80121
rect 525 80112 528 80146
rect 547 80121 548 80141
rect 557 80121 564 80131
rect 514 80105 530 80111
rect 532 80105 548 80111
rect 332 80057 373 80085
rect 332 80051 351 80057
rect 107 79997 119 80031
rect 129 79997 149 80031
rect 196 80010 204 80044
rect 216 80010 232 80044
rect 244 80038 257 80044
rect 278 80038 291 80048
rect 244 80014 291 80038
rect 300 80038 321 80048
rect 336 80041 351 80051
rect 300 80014 329 80038
rect 332 80023 351 80041
rect 361 80051 375 80057
rect 400 80051 411 80089
rect 562 80052 612 80054
rect 361 80023 381 80051
rect 400 80023 409 80051
rect 466 80043 497 80051
rect 565 80043 596 80051
rect 442 80036 500 80043
rect 466 80035 500 80036
rect 565 80035 599 80043
rect 244 80010 257 80014
rect 42 79931 46 79965
rect 72 79931 76 79965
rect 42 79884 76 79888
rect 42 79869 46 79884
rect 72 79869 76 79884
rect 38 79851 80 79869
rect 16 79845 102 79851
rect 144 79845 148 79997
rect 174 79973 181 80001
rect 224 79963 226 80010
rect 300 80001 308 80014
rect 278 79990 305 80001
rect 332 79973 342 80023
rect 400 80003 404 80023
rect 497 80019 500 80035
rect 596 80019 599 80035
rect 466 80018 500 80019
rect 442 80011 500 80018
rect 565 80011 599 80019
rect 612 80002 614 80052
rect 256 79963 328 79971
rect 336 79965 342 79973
rect 400 79965 404 79973
rect 196 79933 204 79963
rect 216 79933 232 79963
rect 196 79929 232 79933
rect 196 79921 226 79929
rect 224 79905 226 79921
rect 332 79893 336 79961
rect 400 79931 408 79965
rect 434 79931 438 79965
rect 454 79949 504 79951
rect 504 79933 506 79949
rect 514 79943 530 79949
rect 532 79943 548 79949
rect 525 79933 548 79942
rect 400 79923 404 79931
rect 498 79923 506 79933
rect 504 79899 506 79923
rect 514 79913 515 79933
rect 525 79908 528 79933
rect 547 79913 548 79933
rect 557 79923 564 79933
rect 514 79899 548 79903
rect 400 79893 442 79894
rect 174 79883 246 79891
rect 400 79886 404 79893
rect 295 79852 300 79886
rect 324 79852 329 79886
rect 367 79869 438 79886
rect 367 79852 442 79869
rect 400 79851 442 79852
rect 378 79845 464 79851
rect 38 79829 80 79845
rect 400 79829 442 79845
rect -25 79815 25 79817
rect 42 79815 76 79829
rect 404 79815 438 79829
rect 455 79815 505 79817
rect 557 79815 607 79817
rect 16 79807 102 79815
rect 378 79807 464 79815
rect 8 79773 17 79807
rect 18 79805 51 79807
rect 80 79805 100 79807
rect 18 79773 100 79805
rect 380 79805 404 79807
rect 429 79805 438 79807
rect 442 79805 462 79807
rect 16 79765 102 79773
rect 42 79749 76 79765
rect 16 79729 38 79735
rect 42 79726 76 79730
rect 80 79729 102 79735
rect 42 79696 46 79726
rect 72 79696 76 79726
rect 42 79615 46 79649
rect 72 79615 76 79649
rect -25 79578 25 79580
rect -8 79570 14 79577
rect -8 79569 17 79570
rect 25 79569 27 79578
rect -12 79562 38 79569
rect -12 79561 34 79562
rect -12 79557 8 79561
rect 0 79545 8 79557
rect 14 79545 34 79561
rect 0 79544 34 79545
rect 0 79537 38 79544
rect 14 79536 17 79537
rect 25 79528 27 79537
rect 42 79508 45 79598
rect 69 79583 80 79615
rect 107 79583 143 79611
rect 144 79583 148 79803
rect 332 79735 336 79803
rect 380 79773 462 79805
rect 463 79773 472 79807
rect 480 79773 497 79807
rect 378 79765 464 79773
rect 505 79765 507 79815
rect 514 79773 548 79807
rect 565 79773 582 79807
rect 607 79765 609 79815
rect 404 79749 438 79765
rect 400 79735 442 79736
rect 378 79729 404 79735
rect 442 79729 464 79735
rect 400 79728 404 79729
rect 174 79689 246 79697
rect 295 79694 300 79728
rect 324 79694 329 79728
rect 224 79659 226 79675
rect 196 79651 226 79659
rect 332 79657 336 79725
rect 367 79694 438 79728
rect 400 79687 404 79694
rect 454 79681 504 79683
rect 494 79677 548 79681
rect 494 79672 514 79677
rect 504 79657 506 79672
rect 196 79647 232 79651
rect 196 79617 204 79647
rect 216 79617 232 79647
rect 400 79649 404 79657
rect 107 79577 119 79583
rect 109 79549 119 79577
rect 129 79549 149 79583
rect 174 79579 181 79609
rect 224 79570 226 79617
rect 256 79609 328 79617
rect 332 79615 336 79645
rect 400 79615 408 79649
rect 434 79615 438 79649
rect 498 79647 506 79657
rect 514 79647 515 79667
rect 504 79631 506 79647
rect 525 79638 528 79672
rect 547 79647 548 79667
rect 557 79647 564 79657
rect 514 79631 530 79637
rect 532 79631 548 79637
rect 278 79579 305 79590
rect 42 79457 46 79491
rect 72 79457 76 79491
rect 38 79419 80 79420
rect 42 79378 76 79412
rect 79 79378 113 79412
rect 42 79299 46 79333
rect 72 79299 76 79333
rect -25 79262 25 79264
rect -8 79254 14 79261
rect -8 79253 17 79254
rect 25 79253 27 79262
rect -12 79246 38 79253
rect -12 79245 34 79246
rect -12 79241 8 79245
rect 0 79229 8 79241
rect 14 79229 34 79245
rect 0 79228 34 79229
rect 0 79221 38 79228
rect 14 79220 17 79221
rect 25 79212 27 79221
rect 42 79192 45 79282
rect 71 79251 80 79279
rect 69 79213 80 79251
rect 144 79241 148 79549
rect 196 79536 204 79570
rect 216 79536 232 79570
rect 244 79566 257 79570
rect 300 79566 308 79579
rect 332 79577 342 79615
rect 400 79607 404 79615
rect 336 79567 342 79577
rect 244 79542 291 79566
rect 244 79536 257 79542
rect 224 79489 226 79536
rect 278 79532 291 79542
rect 300 79542 329 79566
rect 332 79557 342 79567
rect 400 79567 409 79595
rect 562 79578 612 79580
rect 466 79569 497 79577
rect 565 79569 596 79577
rect 300 79532 321 79542
rect 300 79526 308 79532
rect 289 79516 308 79526
rect 196 79459 204 79489
rect 216 79459 232 79489
rect 196 79455 232 79459
rect 196 79447 226 79455
rect 300 79447 308 79516
rect 332 79523 351 79557
rect 361 79529 381 79557
rect 361 79523 375 79529
rect 400 79523 411 79567
rect 442 79562 500 79569
rect 466 79561 500 79562
rect 565 79561 599 79569
rect 497 79545 500 79561
rect 596 79545 599 79561
rect 466 79544 500 79545
rect 442 79537 500 79544
rect 565 79537 599 79545
rect 612 79528 614 79578
rect 332 79499 342 79523
rect 336 79487 342 79499
rect 224 79431 226 79447
rect 332 79419 342 79487
rect 400 79491 404 79499
rect 400 79457 408 79491
rect 434 79457 438 79491
rect 454 79475 504 79477
rect 504 79459 506 79475
rect 514 79469 530 79475
rect 532 79469 548 79475
rect 525 79459 548 79468
rect 400 79449 404 79457
rect 498 79449 506 79459
rect 504 79425 506 79449
rect 514 79439 515 79459
rect 525 79434 528 79459
rect 547 79439 548 79459
rect 557 79449 564 79459
rect 514 79425 548 79429
rect 151 79378 156 79412
rect 174 79409 246 79417
rect 256 79409 328 79417
rect 336 79411 342 79419
rect 400 79414 404 79419
rect 180 79381 185 79409
rect 174 79373 246 79381
rect 256 79373 328 79381
rect 332 79379 336 79409
rect 400 79380 438 79414
rect 224 79343 226 79359
rect 196 79335 226 79343
rect 196 79331 232 79335
rect 196 79301 204 79331
rect 216 79301 232 79331
rect 224 79254 226 79301
rect 300 79274 308 79343
rect 332 79341 342 79379
rect 400 79371 404 79380
rect 454 79365 504 79367
rect 494 79361 548 79365
rect 494 79356 514 79361
rect 504 79341 506 79356
rect 336 79329 342 79341
rect 289 79264 308 79274
rect 300 79258 308 79264
rect 332 79295 342 79329
rect 400 79333 404 79341
rect 400 79299 408 79333
rect 434 79299 438 79333
rect 498 79331 506 79341
rect 514 79331 515 79351
rect 504 79315 506 79331
rect 525 79322 528 79356
rect 547 79331 548 79351
rect 557 79331 564 79341
rect 514 79315 530 79321
rect 532 79315 548 79321
rect 332 79267 373 79295
rect 332 79261 351 79267
rect 107 79207 119 79241
rect 129 79207 149 79241
rect 196 79220 204 79254
rect 216 79220 232 79254
rect 244 79248 257 79254
rect 278 79248 291 79258
rect 244 79224 291 79248
rect 300 79248 321 79258
rect 336 79251 351 79261
rect 300 79224 329 79248
rect 332 79233 351 79251
rect 361 79261 375 79267
rect 400 79261 411 79299
rect 562 79262 612 79264
rect 361 79233 381 79261
rect 400 79233 409 79261
rect 466 79253 497 79261
rect 565 79253 596 79261
rect 442 79246 500 79253
rect 466 79245 500 79246
rect 565 79245 599 79253
rect 244 79220 257 79224
rect 42 79141 46 79175
rect 72 79141 76 79175
rect 42 79094 76 79098
rect 42 79079 46 79094
rect 72 79079 76 79094
rect 38 79061 80 79079
rect 16 79055 102 79061
rect 144 79055 148 79207
rect 174 79183 181 79211
rect 224 79173 226 79220
rect 300 79211 308 79224
rect 278 79200 305 79211
rect 332 79183 342 79233
rect 400 79213 404 79233
rect 497 79229 500 79245
rect 596 79229 599 79245
rect 466 79228 500 79229
rect 442 79221 500 79228
rect 565 79221 599 79229
rect 612 79212 614 79262
rect 256 79173 328 79181
rect 336 79175 342 79183
rect 400 79175 404 79183
rect 196 79143 204 79173
rect 216 79143 232 79173
rect 196 79139 232 79143
rect 196 79131 226 79139
rect 224 79115 226 79131
rect 332 79103 336 79171
rect 400 79141 408 79175
rect 434 79141 438 79175
rect 454 79159 504 79161
rect 504 79143 506 79159
rect 514 79153 530 79159
rect 532 79153 548 79159
rect 525 79143 548 79152
rect 400 79133 404 79141
rect 498 79133 506 79143
rect 504 79109 506 79133
rect 514 79123 515 79143
rect 525 79118 528 79143
rect 547 79123 548 79143
rect 557 79133 564 79143
rect 514 79109 548 79113
rect 400 79103 442 79104
rect 174 79093 246 79101
rect 400 79096 404 79103
rect 295 79062 300 79096
rect 324 79062 329 79096
rect 367 79079 438 79096
rect 367 79062 442 79079
rect 400 79061 442 79062
rect 378 79055 464 79061
rect 38 79039 80 79055
rect 400 79039 442 79055
rect -25 79025 25 79027
rect 42 79025 76 79039
rect 404 79025 438 79039
rect 455 79025 505 79027
rect 557 79025 607 79027
rect 16 79017 102 79025
rect 378 79017 464 79025
rect 8 78983 17 79017
rect 18 79015 51 79017
rect 80 79015 100 79017
rect 18 78983 100 79015
rect 380 79015 404 79017
rect 429 79015 438 79017
rect 442 79015 462 79017
rect 16 78975 102 78983
rect 42 78959 76 78975
rect 16 78939 38 78945
rect 42 78936 76 78940
rect 80 78939 102 78945
rect 42 78906 46 78936
rect 72 78906 76 78936
rect 42 78825 46 78859
rect 72 78825 76 78859
rect -25 78788 25 78790
rect -8 78780 14 78787
rect -8 78779 17 78780
rect 25 78779 27 78788
rect -12 78772 38 78779
rect -12 78771 34 78772
rect -12 78767 8 78771
rect 0 78755 8 78767
rect 14 78755 34 78771
rect 0 78754 34 78755
rect 0 78747 38 78754
rect 14 78746 17 78747
rect 25 78738 27 78747
rect 42 78718 45 78808
rect 69 78793 80 78825
rect 107 78793 143 78821
rect 144 78793 148 79013
rect 332 78945 336 79013
rect 380 78983 462 79015
rect 463 78983 472 79017
rect 480 78983 497 79017
rect 378 78975 464 78983
rect 505 78975 507 79025
rect 514 78983 548 79017
rect 565 78983 582 79017
rect 607 78975 609 79025
rect 404 78959 438 78975
rect 400 78945 442 78946
rect 378 78939 404 78945
rect 442 78939 464 78945
rect 400 78938 404 78939
rect 174 78899 246 78907
rect 295 78904 300 78938
rect 324 78904 329 78938
rect 224 78869 226 78885
rect 196 78861 226 78869
rect 332 78867 336 78935
rect 367 78904 438 78938
rect 400 78897 404 78904
rect 454 78891 504 78893
rect 494 78887 548 78891
rect 494 78882 514 78887
rect 504 78867 506 78882
rect 196 78857 232 78861
rect 196 78827 204 78857
rect 216 78827 232 78857
rect 400 78859 404 78867
rect 107 78787 119 78793
rect 109 78759 119 78787
rect 129 78759 149 78793
rect 174 78789 181 78819
rect 224 78780 226 78827
rect 256 78819 328 78827
rect 332 78825 336 78855
rect 400 78825 408 78859
rect 434 78825 438 78859
rect 498 78857 506 78867
rect 514 78857 515 78877
rect 504 78841 506 78857
rect 525 78848 528 78882
rect 547 78857 548 78877
rect 557 78857 564 78867
rect 514 78841 530 78847
rect 532 78841 548 78847
rect 278 78789 305 78800
rect 42 78667 46 78701
rect 72 78667 76 78701
rect 38 78629 80 78630
rect 42 78588 76 78622
rect 79 78588 113 78622
rect 42 78509 46 78543
rect 72 78509 76 78543
rect -25 78472 25 78474
rect -8 78464 14 78471
rect -8 78463 17 78464
rect 25 78463 27 78472
rect -12 78456 38 78463
rect -12 78455 34 78456
rect -12 78451 8 78455
rect 0 78439 8 78451
rect 14 78439 34 78455
rect 0 78438 34 78439
rect 0 78431 38 78438
rect 14 78430 17 78431
rect 25 78422 27 78431
rect 42 78402 45 78492
rect 71 78461 80 78489
rect 69 78423 80 78461
rect 144 78451 148 78759
rect 196 78746 204 78780
rect 216 78746 232 78780
rect 244 78776 257 78780
rect 300 78776 308 78789
rect 332 78787 342 78825
rect 400 78817 404 78825
rect 336 78777 342 78787
rect 244 78752 291 78776
rect 244 78746 257 78752
rect 224 78699 226 78746
rect 278 78742 291 78752
rect 300 78752 329 78776
rect 332 78767 342 78777
rect 400 78777 409 78805
rect 562 78788 612 78790
rect 466 78779 497 78787
rect 565 78779 596 78787
rect 300 78742 321 78752
rect 300 78736 308 78742
rect 289 78726 308 78736
rect 196 78669 204 78699
rect 216 78669 232 78699
rect 196 78665 232 78669
rect 196 78657 226 78665
rect 300 78657 308 78726
rect 332 78733 351 78767
rect 361 78739 381 78767
rect 361 78733 375 78739
rect 400 78733 411 78777
rect 442 78772 500 78779
rect 466 78771 500 78772
rect 565 78771 599 78779
rect 497 78755 500 78771
rect 596 78755 599 78771
rect 466 78754 500 78755
rect 442 78747 500 78754
rect 565 78747 599 78755
rect 612 78738 614 78788
rect 332 78709 342 78733
rect 336 78697 342 78709
rect 224 78641 226 78657
rect 332 78629 342 78697
rect 400 78701 404 78709
rect 400 78667 408 78701
rect 434 78667 438 78701
rect 454 78685 504 78687
rect 504 78669 506 78685
rect 514 78679 530 78685
rect 532 78679 548 78685
rect 525 78669 548 78678
rect 400 78659 404 78667
rect 498 78659 506 78669
rect 504 78635 506 78659
rect 514 78649 515 78669
rect 525 78644 528 78669
rect 547 78649 548 78669
rect 557 78659 564 78669
rect 514 78635 548 78639
rect 151 78588 156 78622
rect 174 78619 246 78627
rect 256 78619 328 78627
rect 336 78621 342 78629
rect 400 78624 404 78629
rect 180 78591 185 78619
rect 174 78583 246 78591
rect 256 78583 328 78591
rect 332 78589 336 78619
rect 400 78590 438 78624
rect 224 78553 226 78569
rect 196 78545 226 78553
rect 196 78541 232 78545
rect 196 78511 204 78541
rect 216 78511 232 78541
rect 224 78464 226 78511
rect 300 78484 308 78553
rect 332 78551 342 78589
rect 400 78581 404 78590
rect 454 78575 504 78577
rect 494 78571 548 78575
rect 494 78566 514 78571
rect 504 78551 506 78566
rect 336 78539 342 78551
rect 289 78474 308 78484
rect 300 78468 308 78474
rect 332 78505 342 78539
rect 400 78543 404 78551
rect 400 78509 408 78543
rect 434 78509 438 78543
rect 498 78541 506 78551
rect 514 78541 515 78561
rect 504 78525 506 78541
rect 525 78532 528 78566
rect 547 78541 548 78561
rect 557 78541 564 78551
rect 514 78525 530 78531
rect 532 78525 548 78531
rect 332 78477 373 78505
rect 332 78471 351 78477
rect 107 78417 119 78451
rect 129 78417 149 78451
rect 196 78430 204 78464
rect 216 78430 232 78464
rect 244 78458 257 78464
rect 278 78458 291 78468
rect 244 78434 291 78458
rect 300 78458 321 78468
rect 336 78461 351 78471
rect 300 78434 329 78458
rect 332 78443 351 78461
rect 361 78471 375 78477
rect 400 78471 411 78509
rect 562 78472 612 78474
rect 361 78443 381 78471
rect 400 78443 409 78471
rect 466 78463 497 78471
rect 565 78463 596 78471
rect 442 78456 500 78463
rect 466 78455 500 78456
rect 565 78455 599 78463
rect 244 78430 257 78434
rect 42 78351 46 78385
rect 72 78351 76 78385
rect 42 78304 76 78308
rect 42 78289 46 78304
rect 72 78289 76 78304
rect 38 78271 80 78289
rect 16 78265 102 78271
rect 144 78265 148 78417
rect 174 78393 181 78421
rect 224 78383 226 78430
rect 300 78421 308 78434
rect 278 78410 305 78421
rect 332 78393 342 78443
rect 400 78423 404 78443
rect 497 78439 500 78455
rect 596 78439 599 78455
rect 466 78438 500 78439
rect 442 78431 500 78438
rect 565 78431 599 78439
rect 612 78422 614 78472
rect 256 78383 328 78391
rect 336 78385 342 78393
rect 400 78385 404 78393
rect 196 78353 204 78383
rect 216 78353 232 78383
rect 196 78349 232 78353
rect 196 78341 226 78349
rect 224 78325 226 78341
rect 332 78313 336 78381
rect 400 78351 408 78385
rect 434 78351 438 78385
rect 454 78369 504 78371
rect 504 78353 506 78369
rect 514 78363 530 78369
rect 532 78363 548 78369
rect 525 78353 548 78362
rect 400 78343 404 78351
rect 498 78343 506 78353
rect 504 78319 506 78343
rect 514 78333 515 78353
rect 525 78328 528 78353
rect 547 78333 548 78353
rect 557 78343 564 78353
rect 514 78319 548 78323
rect 400 78313 442 78314
rect 174 78303 246 78311
rect 400 78306 404 78313
rect 295 78272 300 78306
rect 324 78272 329 78306
rect 367 78289 438 78306
rect 367 78272 442 78289
rect 400 78271 442 78272
rect 378 78265 464 78271
rect 38 78249 80 78265
rect 400 78249 442 78265
rect -25 78235 25 78237
rect 42 78235 76 78249
rect 404 78235 438 78249
rect 455 78235 505 78237
rect 557 78235 607 78237
rect 16 78227 102 78235
rect 378 78227 464 78235
rect 8 78193 17 78227
rect 18 78225 51 78227
rect 80 78225 100 78227
rect 18 78193 100 78225
rect 380 78225 404 78227
rect 429 78225 438 78227
rect 442 78225 462 78227
rect 16 78185 102 78193
rect 42 78169 76 78185
rect 16 78149 38 78155
rect 42 78146 76 78150
rect 80 78149 102 78155
rect 42 78116 46 78146
rect 72 78116 76 78146
rect 42 78035 46 78069
rect 72 78035 76 78069
rect -25 77998 25 78000
rect -8 77990 14 77997
rect -8 77989 17 77990
rect 25 77989 27 77998
rect -12 77982 38 77989
rect -12 77981 34 77982
rect -12 77977 8 77981
rect 0 77965 8 77977
rect 14 77965 34 77981
rect 0 77964 34 77965
rect 0 77957 38 77964
rect 14 77956 17 77957
rect 25 77948 27 77957
rect 42 77928 45 78018
rect 69 78003 80 78035
rect 107 78003 143 78031
rect 144 78003 148 78223
rect 332 78155 336 78223
rect 380 78193 462 78225
rect 463 78193 472 78227
rect 480 78193 497 78227
rect 378 78185 464 78193
rect 505 78185 507 78235
rect 514 78193 548 78227
rect 565 78193 582 78227
rect 607 78185 609 78235
rect 404 78169 438 78185
rect 400 78155 442 78156
rect 378 78149 404 78155
rect 442 78149 464 78155
rect 400 78148 404 78149
rect 174 78109 246 78117
rect 295 78114 300 78148
rect 324 78114 329 78148
rect 224 78079 226 78095
rect 196 78071 226 78079
rect 332 78077 336 78145
rect 367 78114 438 78148
rect 400 78107 404 78114
rect 454 78101 504 78103
rect 494 78097 548 78101
rect 494 78092 514 78097
rect 504 78077 506 78092
rect 196 78067 232 78071
rect 196 78037 204 78067
rect 216 78037 232 78067
rect 400 78069 404 78077
rect 107 77997 119 78003
rect 109 77969 119 77997
rect 129 77969 149 78003
rect 174 77999 181 78029
rect 224 77990 226 78037
rect 256 78029 328 78037
rect 332 78035 336 78065
rect 400 78035 408 78069
rect 434 78035 438 78069
rect 498 78067 506 78077
rect 514 78067 515 78087
rect 504 78051 506 78067
rect 525 78058 528 78092
rect 547 78067 548 78087
rect 557 78067 564 78077
rect 514 78051 530 78057
rect 532 78051 548 78057
rect 278 77999 305 78010
rect 42 77877 46 77911
rect 72 77877 76 77911
rect 38 77839 80 77840
rect 42 77798 76 77832
rect 79 77798 113 77832
rect 42 77719 46 77753
rect 72 77719 76 77753
rect -25 77682 25 77684
rect -8 77674 14 77681
rect -8 77673 17 77674
rect 25 77673 27 77682
rect -12 77666 38 77673
rect -12 77665 34 77666
rect -12 77661 8 77665
rect 0 77649 8 77661
rect 14 77649 34 77665
rect 0 77648 34 77649
rect 0 77641 38 77648
rect 14 77640 17 77641
rect 25 77632 27 77641
rect 42 77612 45 77702
rect 71 77671 80 77699
rect 69 77633 80 77671
rect 144 77661 148 77969
rect 196 77956 204 77990
rect 216 77956 232 77990
rect 244 77986 257 77990
rect 300 77986 308 77999
rect 332 77997 342 78035
rect 400 78027 404 78035
rect 336 77987 342 77997
rect 244 77962 291 77986
rect 244 77956 257 77962
rect 224 77909 226 77956
rect 278 77952 291 77962
rect 300 77962 329 77986
rect 332 77977 342 77987
rect 400 77987 409 78015
rect 562 77998 612 78000
rect 466 77989 497 77997
rect 565 77989 596 77997
rect 300 77952 321 77962
rect 300 77946 308 77952
rect 289 77936 308 77946
rect 196 77879 204 77909
rect 216 77879 232 77909
rect 196 77875 232 77879
rect 196 77867 226 77875
rect 300 77867 308 77936
rect 332 77943 351 77977
rect 361 77949 381 77977
rect 361 77943 375 77949
rect 400 77943 411 77987
rect 442 77982 500 77989
rect 466 77981 500 77982
rect 565 77981 599 77989
rect 497 77965 500 77981
rect 596 77965 599 77981
rect 466 77964 500 77965
rect 442 77957 500 77964
rect 565 77957 599 77965
rect 612 77948 614 77998
rect 332 77919 342 77943
rect 336 77907 342 77919
rect 224 77851 226 77867
rect 332 77839 342 77907
rect 400 77911 404 77919
rect 400 77877 408 77911
rect 434 77877 438 77911
rect 454 77895 504 77897
rect 504 77879 506 77895
rect 514 77889 530 77895
rect 532 77889 548 77895
rect 525 77879 548 77888
rect 400 77869 404 77877
rect 498 77869 506 77879
rect 504 77845 506 77869
rect 514 77859 515 77879
rect 525 77854 528 77879
rect 547 77859 548 77879
rect 557 77869 564 77879
rect 514 77845 548 77849
rect 151 77798 156 77832
rect 174 77829 246 77837
rect 256 77829 328 77837
rect 336 77831 342 77839
rect 400 77834 404 77839
rect 180 77801 185 77829
rect 174 77793 246 77801
rect 256 77793 328 77801
rect 332 77799 336 77829
rect 400 77800 438 77834
rect 224 77763 226 77779
rect 196 77755 226 77763
rect 196 77751 232 77755
rect 196 77721 204 77751
rect 216 77721 232 77751
rect 224 77674 226 77721
rect 300 77694 308 77763
rect 332 77761 342 77799
rect 400 77791 404 77800
rect 454 77785 504 77787
rect 494 77781 548 77785
rect 494 77776 514 77781
rect 504 77761 506 77776
rect 336 77749 342 77761
rect 289 77684 308 77694
rect 300 77678 308 77684
rect 332 77715 342 77749
rect 400 77753 404 77761
rect 400 77719 408 77753
rect 434 77719 438 77753
rect 498 77751 506 77761
rect 514 77751 515 77771
rect 504 77735 506 77751
rect 525 77742 528 77776
rect 547 77751 548 77771
rect 557 77751 564 77761
rect 514 77735 530 77741
rect 532 77735 548 77741
rect 332 77687 373 77715
rect 332 77681 351 77687
rect 107 77627 119 77661
rect 129 77627 149 77661
rect 196 77640 204 77674
rect 216 77640 232 77674
rect 244 77668 257 77674
rect 278 77668 291 77678
rect 244 77644 291 77668
rect 300 77668 321 77678
rect 336 77671 351 77681
rect 300 77644 329 77668
rect 332 77653 351 77671
rect 361 77681 375 77687
rect 400 77681 411 77719
rect 562 77682 612 77684
rect 361 77653 381 77681
rect 400 77653 409 77681
rect 466 77673 497 77681
rect 565 77673 596 77681
rect 442 77666 500 77673
rect 466 77665 500 77666
rect 565 77665 599 77673
rect 244 77640 257 77644
rect 42 77561 46 77595
rect 72 77561 76 77595
rect 42 77514 76 77518
rect 42 77499 46 77514
rect 72 77499 76 77514
rect 38 77481 80 77499
rect 16 77475 102 77481
rect 144 77475 148 77627
rect 174 77603 181 77631
rect 224 77593 226 77640
rect 300 77631 308 77644
rect 278 77620 305 77631
rect 332 77603 342 77653
rect 400 77633 404 77653
rect 497 77649 500 77665
rect 596 77649 599 77665
rect 466 77648 500 77649
rect 442 77641 500 77648
rect 565 77641 599 77649
rect 612 77632 614 77682
rect 256 77593 328 77601
rect 336 77595 342 77603
rect 400 77595 404 77603
rect 196 77563 204 77593
rect 216 77563 232 77593
rect 196 77559 232 77563
rect 196 77551 226 77559
rect 224 77535 226 77551
rect 332 77523 336 77591
rect 400 77561 408 77595
rect 434 77561 438 77595
rect 454 77579 504 77581
rect 504 77563 506 77579
rect 514 77573 530 77579
rect 532 77573 548 77579
rect 525 77563 548 77572
rect 400 77553 404 77561
rect 498 77553 506 77563
rect 504 77529 506 77553
rect 514 77543 515 77563
rect 525 77538 528 77563
rect 547 77543 548 77563
rect 557 77553 564 77563
rect 514 77529 548 77533
rect 400 77523 442 77524
rect 174 77513 246 77521
rect 400 77516 404 77523
rect 295 77482 300 77516
rect 324 77482 329 77516
rect 367 77499 438 77516
rect 367 77482 442 77499
rect 400 77481 442 77482
rect 378 77475 464 77481
rect 38 77459 80 77475
rect 400 77459 442 77475
rect -25 77445 25 77447
rect 42 77445 76 77459
rect 404 77445 438 77459
rect 455 77445 505 77447
rect 557 77445 607 77447
rect 16 77437 102 77445
rect 378 77437 464 77445
rect 8 77403 17 77437
rect 18 77435 51 77437
rect 80 77435 100 77437
rect 18 77403 100 77435
rect 380 77435 404 77437
rect 429 77435 438 77437
rect 442 77435 462 77437
rect 16 77395 102 77403
rect 42 77379 76 77395
rect 16 77359 38 77365
rect 42 77356 76 77360
rect 80 77359 102 77365
rect 42 77326 46 77356
rect 72 77326 76 77356
rect 42 77245 46 77279
rect 72 77245 76 77279
rect -25 77208 25 77210
rect -8 77200 14 77207
rect -8 77199 17 77200
rect 25 77199 27 77208
rect -12 77192 38 77199
rect -12 77191 34 77192
rect -12 77187 8 77191
rect 0 77175 8 77187
rect 14 77175 34 77191
rect 0 77174 34 77175
rect 0 77167 38 77174
rect 14 77166 17 77167
rect 25 77158 27 77167
rect 42 77138 45 77228
rect 69 77213 80 77245
rect 107 77213 143 77241
rect 144 77213 148 77433
rect 332 77365 336 77433
rect 380 77403 462 77435
rect 463 77403 472 77437
rect 480 77403 497 77437
rect 378 77395 464 77403
rect 505 77395 507 77445
rect 514 77403 548 77437
rect 565 77403 582 77437
rect 607 77395 609 77445
rect 404 77379 438 77395
rect 400 77365 442 77366
rect 378 77359 404 77365
rect 442 77359 464 77365
rect 400 77358 404 77359
rect 174 77319 246 77327
rect 295 77324 300 77358
rect 324 77324 329 77358
rect 224 77289 226 77305
rect 196 77281 226 77289
rect 332 77287 336 77355
rect 367 77324 438 77358
rect 400 77317 404 77324
rect 454 77311 504 77313
rect 494 77307 548 77311
rect 494 77302 514 77307
rect 504 77287 506 77302
rect 196 77277 232 77281
rect 196 77247 204 77277
rect 216 77247 232 77277
rect 400 77279 404 77287
rect 107 77207 119 77213
rect 109 77179 119 77207
rect 129 77179 149 77213
rect 174 77209 181 77239
rect 224 77200 226 77247
rect 256 77239 328 77247
rect 332 77245 336 77275
rect 400 77245 408 77279
rect 434 77245 438 77279
rect 498 77277 506 77287
rect 514 77277 515 77297
rect 504 77261 506 77277
rect 525 77268 528 77302
rect 547 77277 548 77297
rect 557 77277 564 77287
rect 514 77261 530 77267
rect 532 77261 548 77267
rect 278 77209 305 77220
rect 42 77087 46 77121
rect 72 77087 76 77121
rect 38 77049 80 77050
rect 42 77008 76 77042
rect 79 77008 113 77042
rect 42 76929 46 76963
rect 72 76929 76 76963
rect -25 76892 25 76894
rect -8 76884 14 76891
rect -8 76883 17 76884
rect 25 76883 27 76892
rect -12 76876 38 76883
rect -12 76875 34 76876
rect -12 76871 8 76875
rect 0 76859 8 76871
rect 14 76859 34 76875
rect 0 76858 34 76859
rect 0 76851 38 76858
rect 14 76850 17 76851
rect 25 76842 27 76851
rect 42 76822 45 76912
rect 71 76881 80 76909
rect 69 76843 80 76881
rect 144 76871 148 77179
rect 196 77166 204 77200
rect 216 77166 232 77200
rect 244 77196 257 77200
rect 300 77196 308 77209
rect 332 77207 342 77245
rect 400 77237 404 77245
rect 336 77197 342 77207
rect 244 77172 291 77196
rect 244 77166 257 77172
rect 224 77119 226 77166
rect 278 77162 291 77172
rect 300 77172 329 77196
rect 332 77187 342 77197
rect 400 77197 409 77225
rect 562 77208 612 77210
rect 466 77199 497 77207
rect 565 77199 596 77207
rect 300 77162 321 77172
rect 300 77156 308 77162
rect 289 77146 308 77156
rect 196 77089 204 77119
rect 216 77089 232 77119
rect 196 77085 232 77089
rect 196 77077 226 77085
rect 300 77077 308 77146
rect 332 77153 351 77187
rect 361 77159 381 77187
rect 361 77153 375 77159
rect 400 77153 411 77197
rect 442 77192 500 77199
rect 466 77191 500 77192
rect 565 77191 599 77199
rect 497 77175 500 77191
rect 596 77175 599 77191
rect 466 77174 500 77175
rect 442 77167 500 77174
rect 565 77167 599 77175
rect 612 77158 614 77208
rect 332 77129 342 77153
rect 336 77117 342 77129
rect 224 77061 226 77077
rect 332 77049 342 77117
rect 400 77121 404 77129
rect 400 77087 408 77121
rect 434 77087 438 77121
rect 454 77105 504 77107
rect 504 77089 506 77105
rect 514 77099 530 77105
rect 532 77099 548 77105
rect 525 77089 548 77098
rect 400 77079 404 77087
rect 498 77079 506 77089
rect 504 77055 506 77079
rect 514 77069 515 77089
rect 525 77064 528 77089
rect 547 77069 548 77089
rect 557 77079 564 77089
rect 514 77055 548 77059
rect 151 77008 156 77042
rect 174 77039 246 77047
rect 256 77039 328 77047
rect 336 77041 342 77049
rect 400 77044 404 77049
rect 180 77011 185 77039
rect 174 77003 246 77011
rect 256 77003 328 77011
rect 332 77009 336 77039
rect 400 77010 438 77044
rect 224 76973 226 76989
rect 196 76965 226 76973
rect 196 76961 232 76965
rect 196 76931 204 76961
rect 216 76931 232 76961
rect 224 76884 226 76931
rect 300 76904 308 76973
rect 332 76971 342 77009
rect 400 77001 404 77010
rect 454 76995 504 76997
rect 494 76991 548 76995
rect 494 76986 514 76991
rect 504 76971 506 76986
rect 336 76959 342 76971
rect 289 76894 308 76904
rect 300 76888 308 76894
rect 332 76925 342 76959
rect 400 76963 404 76971
rect 400 76929 408 76963
rect 434 76929 438 76963
rect 498 76961 506 76971
rect 514 76961 515 76981
rect 504 76945 506 76961
rect 525 76952 528 76986
rect 547 76961 548 76981
rect 557 76961 564 76971
rect 514 76945 530 76951
rect 532 76945 548 76951
rect 332 76897 373 76925
rect 332 76891 351 76897
rect 107 76837 119 76871
rect 129 76837 149 76871
rect 196 76850 204 76884
rect 216 76850 232 76884
rect 244 76878 257 76884
rect 278 76878 291 76888
rect 244 76854 291 76878
rect 300 76878 321 76888
rect 336 76881 351 76891
rect 300 76854 329 76878
rect 332 76863 351 76881
rect 361 76891 375 76897
rect 400 76891 411 76929
rect 562 76892 612 76894
rect 361 76863 381 76891
rect 400 76863 409 76891
rect 466 76883 497 76891
rect 565 76883 596 76891
rect 442 76876 500 76883
rect 466 76875 500 76876
rect 565 76875 599 76883
rect 244 76850 257 76854
rect 42 76771 46 76805
rect 72 76771 76 76805
rect 42 76724 76 76728
rect 42 76709 46 76724
rect 72 76709 76 76724
rect 38 76691 80 76709
rect 16 76685 102 76691
rect 144 76685 148 76837
rect 174 76813 181 76841
rect 224 76803 226 76850
rect 300 76841 308 76854
rect 278 76830 305 76841
rect 332 76813 342 76863
rect 400 76843 404 76863
rect 497 76859 500 76875
rect 596 76859 599 76875
rect 466 76858 500 76859
rect 442 76851 500 76858
rect 565 76851 599 76859
rect 612 76842 614 76892
rect 256 76803 328 76811
rect 336 76805 342 76813
rect 400 76805 404 76813
rect 196 76773 204 76803
rect 216 76773 232 76803
rect 196 76769 232 76773
rect 196 76761 226 76769
rect 224 76745 226 76761
rect 332 76733 336 76801
rect 400 76771 408 76805
rect 434 76771 438 76805
rect 454 76789 504 76791
rect 504 76773 506 76789
rect 514 76783 530 76789
rect 532 76783 548 76789
rect 525 76773 548 76782
rect 400 76763 404 76771
rect 498 76763 506 76773
rect 504 76739 506 76763
rect 514 76753 515 76773
rect 525 76748 528 76773
rect 547 76753 548 76773
rect 557 76763 564 76773
rect 514 76739 548 76743
rect 400 76733 442 76734
rect 174 76723 246 76731
rect 400 76726 404 76733
rect 295 76692 300 76726
rect 324 76692 329 76726
rect 367 76709 438 76726
rect 367 76692 442 76709
rect 400 76691 442 76692
rect 378 76685 464 76691
rect 38 76669 80 76685
rect 400 76669 442 76685
rect -25 76655 25 76657
rect 42 76655 76 76669
rect 404 76655 438 76669
rect 455 76655 505 76657
rect 557 76655 607 76657
rect 16 76647 102 76655
rect 378 76647 464 76655
rect 8 76613 17 76647
rect 18 76645 51 76647
rect 80 76645 100 76647
rect 18 76613 100 76645
rect 380 76645 404 76647
rect 429 76645 438 76647
rect 442 76645 462 76647
rect 16 76605 102 76613
rect 42 76589 76 76605
rect 16 76569 38 76575
rect 42 76566 76 76570
rect 80 76569 102 76575
rect 42 76536 46 76566
rect 72 76536 76 76566
rect 42 76455 46 76489
rect 72 76455 76 76489
rect -25 76418 25 76420
rect -8 76410 14 76417
rect -8 76409 17 76410
rect 25 76409 27 76418
rect -12 76402 38 76409
rect -12 76401 34 76402
rect -12 76397 8 76401
rect 0 76385 8 76397
rect 14 76385 34 76401
rect 0 76384 34 76385
rect 0 76377 38 76384
rect 14 76376 17 76377
rect 25 76368 27 76377
rect 42 76348 45 76438
rect 69 76423 80 76455
rect 107 76423 143 76451
rect 144 76423 148 76643
rect 332 76575 336 76643
rect 380 76613 462 76645
rect 463 76613 472 76647
rect 480 76613 497 76647
rect 378 76605 464 76613
rect 505 76605 507 76655
rect 514 76613 548 76647
rect 565 76613 582 76647
rect 607 76605 609 76655
rect 404 76589 438 76605
rect 400 76575 442 76576
rect 378 76569 404 76575
rect 442 76569 464 76575
rect 400 76568 404 76569
rect 174 76529 246 76537
rect 295 76534 300 76568
rect 324 76534 329 76568
rect 224 76499 226 76515
rect 196 76491 226 76499
rect 332 76497 336 76565
rect 367 76534 438 76568
rect 400 76527 404 76534
rect 454 76521 504 76523
rect 494 76517 548 76521
rect 494 76512 514 76517
rect 504 76497 506 76512
rect 196 76487 232 76491
rect 196 76457 204 76487
rect 216 76457 232 76487
rect 400 76489 404 76497
rect 107 76417 119 76423
rect 109 76389 119 76417
rect 129 76389 149 76423
rect 174 76419 181 76449
rect 224 76410 226 76457
rect 256 76449 328 76457
rect 332 76455 336 76485
rect 400 76455 408 76489
rect 434 76455 438 76489
rect 498 76487 506 76497
rect 514 76487 515 76507
rect 504 76471 506 76487
rect 525 76478 528 76512
rect 547 76487 548 76507
rect 557 76487 564 76497
rect 514 76471 530 76477
rect 532 76471 548 76477
rect 278 76419 305 76430
rect 42 76297 46 76331
rect 72 76297 76 76331
rect 38 76259 80 76260
rect 42 76218 76 76252
rect 79 76218 113 76252
rect 42 76139 46 76173
rect 72 76139 76 76173
rect -25 76102 25 76104
rect -8 76094 14 76101
rect -8 76093 17 76094
rect 25 76093 27 76102
rect -12 76086 38 76093
rect -12 76085 34 76086
rect -12 76081 8 76085
rect 0 76069 8 76081
rect 14 76069 34 76085
rect 0 76068 34 76069
rect 0 76061 38 76068
rect 14 76060 17 76061
rect 25 76052 27 76061
rect 42 76032 45 76122
rect 71 76091 80 76119
rect 69 76053 80 76091
rect 144 76081 148 76389
rect 196 76376 204 76410
rect 216 76376 232 76410
rect 244 76406 257 76410
rect 300 76406 308 76419
rect 332 76417 342 76455
rect 400 76447 404 76455
rect 336 76407 342 76417
rect 244 76382 291 76406
rect 244 76376 257 76382
rect 224 76329 226 76376
rect 278 76372 291 76382
rect 300 76382 329 76406
rect 332 76397 342 76407
rect 400 76407 409 76435
rect 562 76418 612 76420
rect 466 76409 497 76417
rect 565 76409 596 76417
rect 300 76372 321 76382
rect 300 76366 308 76372
rect 289 76356 308 76366
rect 196 76299 204 76329
rect 216 76299 232 76329
rect 196 76295 232 76299
rect 196 76287 226 76295
rect 300 76287 308 76356
rect 332 76363 351 76397
rect 361 76369 381 76397
rect 361 76363 375 76369
rect 400 76363 411 76407
rect 442 76402 500 76409
rect 466 76401 500 76402
rect 565 76401 599 76409
rect 497 76385 500 76401
rect 596 76385 599 76401
rect 466 76384 500 76385
rect 442 76377 500 76384
rect 565 76377 599 76385
rect 612 76368 614 76418
rect 332 76339 342 76363
rect 336 76327 342 76339
rect 224 76271 226 76287
rect 332 76259 342 76327
rect 400 76331 404 76339
rect 400 76297 408 76331
rect 434 76297 438 76331
rect 454 76315 504 76317
rect 504 76299 506 76315
rect 514 76309 530 76315
rect 532 76309 548 76315
rect 525 76299 548 76308
rect 400 76289 404 76297
rect 498 76289 506 76299
rect 504 76265 506 76289
rect 514 76279 515 76299
rect 525 76274 528 76299
rect 547 76279 548 76299
rect 557 76289 564 76299
rect 514 76265 548 76269
rect 151 76218 156 76252
rect 174 76249 246 76257
rect 256 76249 328 76257
rect 336 76251 342 76259
rect 400 76254 404 76259
rect 180 76221 185 76249
rect 174 76213 246 76221
rect 256 76213 328 76221
rect 332 76219 336 76249
rect 400 76220 438 76254
rect 224 76183 226 76199
rect 196 76175 226 76183
rect 196 76171 232 76175
rect 196 76141 204 76171
rect 216 76141 232 76171
rect 224 76094 226 76141
rect 300 76114 308 76183
rect 332 76181 342 76219
rect 400 76211 404 76220
rect 454 76205 504 76207
rect 494 76201 548 76205
rect 494 76196 514 76201
rect 504 76181 506 76196
rect 336 76169 342 76181
rect 289 76104 308 76114
rect 300 76098 308 76104
rect 332 76135 342 76169
rect 400 76173 404 76181
rect 400 76139 408 76173
rect 434 76139 438 76173
rect 498 76171 506 76181
rect 514 76171 515 76191
rect 504 76155 506 76171
rect 525 76162 528 76196
rect 547 76171 548 76191
rect 557 76171 564 76181
rect 514 76155 530 76161
rect 532 76155 548 76161
rect 332 76107 373 76135
rect 332 76101 351 76107
rect 107 76047 119 76081
rect 129 76047 149 76081
rect 196 76060 204 76094
rect 216 76060 232 76094
rect 244 76088 257 76094
rect 278 76088 291 76098
rect 244 76064 291 76088
rect 300 76088 321 76098
rect 336 76091 351 76101
rect 300 76064 329 76088
rect 332 76073 351 76091
rect 361 76101 375 76107
rect 400 76101 411 76139
rect 562 76102 612 76104
rect 361 76073 381 76101
rect 400 76073 409 76101
rect 466 76093 497 76101
rect 565 76093 596 76101
rect 442 76086 500 76093
rect 466 76085 500 76086
rect 565 76085 599 76093
rect 244 76060 257 76064
rect 42 75981 46 76015
rect 72 75981 76 76015
rect 42 75934 76 75938
rect 42 75919 46 75934
rect 72 75919 76 75934
rect 38 75901 80 75919
rect 16 75895 102 75901
rect 144 75895 148 76047
rect 174 76023 181 76051
rect 224 76013 226 76060
rect 300 76051 308 76064
rect 278 76040 305 76051
rect 332 76023 342 76073
rect 400 76053 404 76073
rect 497 76069 500 76085
rect 596 76069 599 76085
rect 466 76068 500 76069
rect 442 76061 500 76068
rect 565 76061 599 76069
rect 612 76052 614 76102
rect 256 76013 328 76021
rect 336 76015 342 76023
rect 400 76015 404 76023
rect 196 75983 204 76013
rect 216 75983 232 76013
rect 196 75979 232 75983
rect 196 75971 226 75979
rect 224 75955 226 75971
rect 332 75943 336 76011
rect 400 75981 408 76015
rect 434 75981 438 76015
rect 454 75999 504 76001
rect 504 75983 506 75999
rect 514 75993 530 75999
rect 532 75993 548 75999
rect 525 75983 548 75992
rect 400 75973 404 75981
rect 498 75973 506 75983
rect 504 75949 506 75973
rect 514 75963 515 75983
rect 525 75958 528 75983
rect 547 75963 548 75983
rect 557 75973 564 75983
rect 514 75949 548 75953
rect 400 75943 442 75944
rect 174 75933 246 75941
rect 400 75936 404 75943
rect 295 75902 300 75936
rect 324 75902 329 75936
rect 367 75919 438 75936
rect 367 75902 442 75919
rect 400 75901 442 75902
rect 378 75895 464 75901
rect 38 75879 80 75895
rect 400 75879 442 75895
rect -25 75865 25 75867
rect 42 75865 76 75879
rect 404 75865 438 75879
rect 455 75865 505 75867
rect 557 75865 607 75867
rect 16 75857 102 75865
rect 378 75857 464 75865
rect 8 75823 17 75857
rect 18 75855 51 75857
rect 80 75855 100 75857
rect 18 75823 100 75855
rect 380 75855 404 75857
rect 429 75855 438 75857
rect 442 75855 462 75857
rect 16 75815 102 75823
rect 42 75799 76 75815
rect 16 75779 38 75785
rect 42 75776 76 75780
rect 80 75779 102 75785
rect 42 75746 46 75776
rect 72 75746 76 75776
rect 42 75665 46 75699
rect 72 75665 76 75699
rect -25 75628 25 75630
rect -8 75620 14 75627
rect -8 75619 17 75620
rect 25 75619 27 75628
rect -12 75612 38 75619
rect -12 75611 34 75612
rect -12 75607 8 75611
rect 0 75595 8 75607
rect 14 75595 34 75611
rect 0 75594 34 75595
rect 0 75587 38 75594
rect 14 75586 17 75587
rect 25 75578 27 75587
rect 42 75558 45 75648
rect 69 75633 80 75665
rect 107 75633 143 75661
rect 144 75633 148 75853
rect 332 75785 336 75853
rect 380 75823 462 75855
rect 463 75823 472 75857
rect 480 75823 497 75857
rect 378 75815 464 75823
rect 505 75815 507 75865
rect 514 75823 548 75857
rect 565 75823 582 75857
rect 607 75815 609 75865
rect 404 75799 438 75815
rect 400 75785 442 75786
rect 378 75779 404 75785
rect 442 75779 464 75785
rect 400 75778 404 75779
rect 174 75739 246 75747
rect 295 75744 300 75778
rect 324 75744 329 75778
rect 224 75709 226 75725
rect 196 75701 226 75709
rect 332 75707 336 75775
rect 367 75744 438 75778
rect 400 75737 404 75744
rect 454 75731 504 75733
rect 494 75727 548 75731
rect 494 75722 514 75727
rect 504 75707 506 75722
rect 196 75697 232 75701
rect 196 75667 204 75697
rect 216 75667 232 75697
rect 400 75699 404 75707
rect 107 75627 119 75633
rect 109 75599 119 75627
rect 129 75599 149 75633
rect 174 75629 181 75659
rect 224 75620 226 75667
rect 256 75659 328 75667
rect 332 75665 336 75695
rect 400 75665 408 75699
rect 434 75665 438 75699
rect 498 75697 506 75707
rect 514 75697 515 75717
rect 504 75681 506 75697
rect 525 75688 528 75722
rect 547 75697 548 75717
rect 557 75697 564 75707
rect 514 75681 530 75687
rect 532 75681 548 75687
rect 278 75629 305 75640
rect 42 75507 46 75541
rect 72 75507 76 75541
rect 38 75469 80 75470
rect 42 75428 76 75462
rect 79 75428 113 75462
rect 42 75349 46 75383
rect 72 75349 76 75383
rect -25 75312 25 75314
rect -8 75304 14 75311
rect -8 75303 17 75304
rect 25 75303 27 75312
rect -12 75296 38 75303
rect -12 75295 34 75296
rect -12 75291 8 75295
rect 0 75279 8 75291
rect 14 75279 34 75295
rect 0 75278 34 75279
rect 0 75271 38 75278
rect 14 75270 17 75271
rect 25 75262 27 75271
rect 42 75242 45 75332
rect 71 75301 80 75329
rect 69 75263 80 75301
rect 144 75291 148 75599
rect 196 75586 204 75620
rect 216 75586 232 75620
rect 244 75616 257 75620
rect 300 75616 308 75629
rect 332 75627 342 75665
rect 400 75657 404 75665
rect 336 75617 342 75627
rect 244 75592 291 75616
rect 244 75586 257 75592
rect 224 75539 226 75586
rect 278 75582 291 75592
rect 300 75592 329 75616
rect 332 75607 342 75617
rect 400 75617 409 75645
rect 562 75628 612 75630
rect 466 75619 497 75627
rect 565 75619 596 75627
rect 300 75582 321 75592
rect 300 75576 308 75582
rect 289 75566 308 75576
rect 196 75509 204 75539
rect 216 75509 232 75539
rect 196 75505 232 75509
rect 196 75497 226 75505
rect 300 75497 308 75566
rect 332 75573 351 75607
rect 361 75579 381 75607
rect 361 75573 375 75579
rect 400 75573 411 75617
rect 442 75612 500 75619
rect 466 75611 500 75612
rect 565 75611 599 75619
rect 497 75595 500 75611
rect 596 75595 599 75611
rect 466 75594 500 75595
rect 442 75587 500 75594
rect 565 75587 599 75595
rect 612 75578 614 75628
rect 332 75549 342 75573
rect 336 75537 342 75549
rect 224 75481 226 75497
rect 332 75469 342 75537
rect 400 75541 404 75549
rect 400 75507 408 75541
rect 434 75507 438 75541
rect 454 75525 504 75527
rect 504 75509 506 75525
rect 514 75519 530 75525
rect 532 75519 548 75525
rect 525 75509 548 75518
rect 400 75499 404 75507
rect 498 75499 506 75509
rect 504 75475 506 75499
rect 514 75489 515 75509
rect 525 75484 528 75509
rect 547 75489 548 75509
rect 557 75499 564 75509
rect 514 75475 548 75479
rect 151 75428 156 75462
rect 174 75459 246 75467
rect 256 75459 328 75467
rect 336 75461 342 75469
rect 400 75464 404 75469
rect 180 75431 185 75459
rect 174 75423 246 75431
rect 256 75423 328 75431
rect 332 75429 336 75459
rect 400 75430 438 75464
rect 224 75393 226 75409
rect 196 75385 226 75393
rect 196 75381 232 75385
rect 196 75351 204 75381
rect 216 75351 232 75381
rect 224 75304 226 75351
rect 300 75324 308 75393
rect 332 75391 342 75429
rect 400 75421 404 75430
rect 454 75415 504 75417
rect 494 75411 548 75415
rect 494 75406 514 75411
rect 504 75391 506 75406
rect 336 75379 342 75391
rect 289 75314 308 75324
rect 300 75308 308 75314
rect 332 75345 342 75379
rect 400 75383 404 75391
rect 400 75349 408 75383
rect 434 75349 438 75383
rect 498 75381 506 75391
rect 514 75381 515 75401
rect 504 75365 506 75381
rect 525 75372 528 75406
rect 547 75381 548 75401
rect 557 75381 564 75391
rect 514 75365 530 75371
rect 532 75365 548 75371
rect 332 75317 373 75345
rect 332 75311 351 75317
rect 107 75257 119 75291
rect 129 75257 149 75291
rect 196 75270 204 75304
rect 216 75270 232 75304
rect 244 75298 257 75304
rect 278 75298 291 75308
rect 244 75274 291 75298
rect 300 75298 321 75308
rect 336 75301 351 75311
rect 300 75274 329 75298
rect 332 75283 351 75301
rect 361 75311 375 75317
rect 400 75311 411 75349
rect 562 75312 612 75314
rect 361 75283 381 75311
rect 400 75283 409 75311
rect 466 75303 497 75311
rect 565 75303 596 75311
rect 442 75296 500 75303
rect 466 75295 500 75296
rect 565 75295 599 75303
rect 244 75270 257 75274
rect 42 75191 46 75225
rect 72 75191 76 75225
rect 42 75144 76 75148
rect 42 75129 46 75144
rect 72 75129 76 75144
rect 38 75111 80 75129
rect 16 75105 102 75111
rect 144 75105 148 75257
rect 174 75233 181 75261
rect 224 75223 226 75270
rect 300 75261 308 75274
rect 278 75250 305 75261
rect 332 75233 342 75283
rect 400 75263 404 75283
rect 497 75279 500 75295
rect 596 75279 599 75295
rect 466 75278 500 75279
rect 442 75271 500 75278
rect 565 75271 599 75279
rect 612 75262 614 75312
rect 256 75223 328 75231
rect 336 75225 342 75233
rect 400 75225 404 75233
rect 196 75193 204 75223
rect 216 75193 232 75223
rect 196 75189 232 75193
rect 196 75181 226 75189
rect 224 75165 226 75181
rect 332 75153 336 75221
rect 400 75191 408 75225
rect 434 75191 438 75225
rect 454 75209 504 75211
rect 504 75193 506 75209
rect 514 75203 530 75209
rect 532 75203 548 75209
rect 525 75193 548 75202
rect 400 75183 404 75191
rect 498 75183 506 75193
rect 504 75159 506 75183
rect 514 75173 515 75193
rect 525 75168 528 75193
rect 547 75173 548 75193
rect 557 75183 564 75193
rect 514 75159 548 75163
rect 400 75153 442 75154
rect 174 75143 246 75151
rect 400 75146 404 75153
rect 295 75112 300 75146
rect 324 75112 329 75146
rect 367 75129 438 75146
rect 367 75112 442 75129
rect 400 75111 442 75112
rect 378 75105 464 75111
rect 38 75089 80 75105
rect 400 75089 442 75105
rect -25 75075 25 75077
rect 42 75075 76 75089
rect 404 75075 438 75089
rect 455 75075 505 75077
rect 557 75075 607 75077
rect 16 75067 102 75075
rect 378 75067 464 75075
rect 8 75033 17 75067
rect 18 75065 51 75067
rect 80 75065 100 75067
rect 18 75033 100 75065
rect 380 75065 404 75067
rect 429 75065 438 75067
rect 442 75065 462 75067
rect 16 75025 102 75033
rect 42 75009 76 75025
rect 16 74989 38 74995
rect 42 74986 76 74990
rect 80 74989 102 74995
rect 42 74956 46 74986
rect 72 74956 76 74986
rect 42 74875 46 74909
rect 72 74875 76 74909
rect -25 74838 25 74840
rect -8 74830 14 74837
rect -8 74829 17 74830
rect 25 74829 27 74838
rect -12 74822 38 74829
rect -12 74821 34 74822
rect -12 74817 8 74821
rect 0 74805 8 74817
rect 14 74805 34 74821
rect 0 74804 34 74805
rect 0 74797 38 74804
rect 14 74796 17 74797
rect 25 74788 27 74797
rect 42 74768 45 74858
rect 69 74843 80 74875
rect 107 74843 143 74871
rect 144 74843 148 75063
rect 332 74995 336 75063
rect 380 75033 462 75065
rect 463 75033 472 75067
rect 480 75033 497 75067
rect 378 75025 464 75033
rect 505 75025 507 75075
rect 514 75033 548 75067
rect 565 75033 582 75067
rect 607 75025 609 75075
rect 404 75009 438 75025
rect 400 74995 442 74996
rect 378 74989 404 74995
rect 442 74989 464 74995
rect 400 74988 404 74989
rect 174 74949 246 74957
rect 295 74954 300 74988
rect 324 74954 329 74988
rect 224 74919 226 74935
rect 196 74911 226 74919
rect 332 74917 336 74985
rect 367 74954 438 74988
rect 400 74947 404 74954
rect 454 74941 504 74943
rect 494 74937 548 74941
rect 494 74932 514 74937
rect 504 74917 506 74932
rect 196 74907 232 74911
rect 196 74877 204 74907
rect 216 74877 232 74907
rect 400 74909 404 74917
rect 107 74837 119 74843
rect 109 74809 119 74837
rect 129 74809 149 74843
rect 174 74839 181 74869
rect 224 74830 226 74877
rect 256 74869 328 74877
rect 332 74875 336 74905
rect 400 74875 408 74909
rect 434 74875 438 74909
rect 498 74907 506 74917
rect 514 74907 515 74927
rect 504 74891 506 74907
rect 525 74898 528 74932
rect 547 74907 548 74927
rect 557 74907 564 74917
rect 514 74891 530 74897
rect 532 74891 548 74897
rect 278 74839 305 74850
rect 42 74717 46 74751
rect 72 74717 76 74751
rect 38 74679 80 74680
rect 42 74638 76 74672
rect 79 74638 113 74672
rect 42 74559 46 74593
rect 72 74559 76 74593
rect -25 74522 25 74524
rect -8 74514 14 74521
rect -8 74513 17 74514
rect 25 74513 27 74522
rect -12 74506 38 74513
rect -12 74505 34 74506
rect -12 74501 8 74505
rect 0 74489 8 74501
rect 14 74489 34 74505
rect 0 74488 34 74489
rect 0 74481 38 74488
rect 14 74480 17 74481
rect 25 74472 27 74481
rect 42 74452 45 74542
rect 71 74511 80 74539
rect 69 74473 80 74511
rect 144 74501 148 74809
rect 196 74796 204 74830
rect 216 74796 232 74830
rect 244 74826 257 74830
rect 300 74826 308 74839
rect 332 74837 342 74875
rect 400 74867 404 74875
rect 336 74827 342 74837
rect 244 74802 291 74826
rect 244 74796 257 74802
rect 224 74749 226 74796
rect 278 74792 291 74802
rect 300 74802 329 74826
rect 332 74817 342 74827
rect 400 74827 409 74855
rect 562 74838 612 74840
rect 466 74829 497 74837
rect 565 74829 596 74837
rect 300 74792 321 74802
rect 300 74786 308 74792
rect 289 74776 308 74786
rect 196 74719 204 74749
rect 216 74719 232 74749
rect 196 74715 232 74719
rect 196 74707 226 74715
rect 300 74707 308 74776
rect 332 74783 351 74817
rect 361 74789 381 74817
rect 361 74783 375 74789
rect 400 74783 411 74827
rect 442 74822 500 74829
rect 466 74821 500 74822
rect 565 74821 599 74829
rect 497 74805 500 74821
rect 596 74805 599 74821
rect 466 74804 500 74805
rect 442 74797 500 74804
rect 565 74797 599 74805
rect 612 74788 614 74838
rect 332 74759 342 74783
rect 336 74747 342 74759
rect 224 74691 226 74707
rect 332 74679 342 74747
rect 400 74751 404 74759
rect 400 74717 408 74751
rect 434 74717 438 74751
rect 454 74735 504 74737
rect 504 74719 506 74735
rect 514 74729 530 74735
rect 532 74729 548 74735
rect 525 74719 548 74728
rect 400 74709 404 74717
rect 498 74709 506 74719
rect 504 74685 506 74709
rect 514 74699 515 74719
rect 525 74694 528 74719
rect 547 74699 548 74719
rect 557 74709 564 74719
rect 514 74685 548 74689
rect 151 74638 156 74672
rect 174 74669 246 74677
rect 256 74669 328 74677
rect 336 74671 342 74679
rect 400 74674 404 74679
rect 180 74641 185 74669
rect 174 74633 246 74641
rect 256 74633 328 74641
rect 332 74639 336 74669
rect 400 74640 438 74674
rect 224 74603 226 74619
rect 196 74595 226 74603
rect 196 74591 232 74595
rect 196 74561 204 74591
rect 216 74561 232 74591
rect 224 74514 226 74561
rect 300 74534 308 74603
rect 332 74601 342 74639
rect 400 74631 404 74640
rect 454 74625 504 74627
rect 494 74621 548 74625
rect 494 74616 514 74621
rect 504 74601 506 74616
rect 336 74589 342 74601
rect 289 74524 308 74534
rect 300 74518 308 74524
rect 332 74555 342 74589
rect 400 74593 404 74601
rect 400 74559 408 74593
rect 434 74559 438 74593
rect 498 74591 506 74601
rect 514 74591 515 74611
rect 504 74575 506 74591
rect 525 74582 528 74616
rect 547 74591 548 74611
rect 557 74591 564 74601
rect 514 74575 530 74581
rect 532 74575 548 74581
rect 332 74527 373 74555
rect 332 74521 351 74527
rect 107 74467 119 74501
rect 129 74467 149 74501
rect 196 74480 204 74514
rect 216 74480 232 74514
rect 244 74508 257 74514
rect 278 74508 291 74518
rect 244 74484 291 74508
rect 300 74508 321 74518
rect 336 74511 351 74521
rect 300 74484 329 74508
rect 332 74493 351 74511
rect 361 74521 375 74527
rect 400 74521 411 74559
rect 562 74522 612 74524
rect 361 74493 381 74521
rect 400 74493 409 74521
rect 466 74513 497 74521
rect 565 74513 596 74521
rect 442 74506 500 74513
rect 466 74505 500 74506
rect 565 74505 599 74513
rect 244 74480 257 74484
rect 42 74401 46 74435
rect 72 74401 76 74435
rect 42 74354 76 74358
rect 42 74339 46 74354
rect 72 74339 76 74354
rect 38 74321 80 74339
rect 16 74315 102 74321
rect 144 74315 148 74467
rect 174 74443 181 74471
rect 224 74433 226 74480
rect 300 74471 308 74484
rect 278 74460 305 74471
rect 332 74443 342 74493
rect 400 74473 404 74493
rect 497 74489 500 74505
rect 596 74489 599 74505
rect 466 74488 500 74489
rect 442 74481 500 74488
rect 565 74481 599 74489
rect 612 74472 614 74522
rect 256 74433 328 74441
rect 336 74435 342 74443
rect 400 74435 404 74443
rect 196 74403 204 74433
rect 216 74403 232 74433
rect 196 74399 232 74403
rect 196 74391 226 74399
rect 224 74375 226 74391
rect 332 74363 336 74431
rect 400 74401 408 74435
rect 434 74401 438 74435
rect 454 74419 504 74421
rect 504 74403 506 74419
rect 514 74413 530 74419
rect 532 74413 548 74419
rect 525 74403 548 74412
rect 400 74393 404 74401
rect 498 74393 506 74403
rect 504 74369 506 74393
rect 514 74383 515 74403
rect 525 74378 528 74403
rect 547 74383 548 74403
rect 557 74393 564 74403
rect 514 74369 548 74373
rect 400 74363 442 74364
rect 174 74353 246 74361
rect 400 74356 404 74363
rect 295 74322 300 74356
rect 324 74322 329 74356
rect 367 74339 438 74356
rect 367 74322 442 74339
rect 400 74321 442 74322
rect 378 74315 464 74321
rect 38 74299 80 74315
rect 400 74299 442 74315
rect -25 74285 25 74287
rect 42 74285 76 74299
rect 404 74285 438 74299
rect 455 74285 505 74287
rect 557 74285 607 74287
rect 16 74277 102 74285
rect 378 74277 464 74285
rect 8 74243 17 74277
rect 18 74275 51 74277
rect 80 74275 100 74277
rect 18 74243 100 74275
rect 380 74275 404 74277
rect 429 74275 438 74277
rect 442 74275 462 74277
rect 16 74235 102 74243
rect 42 74219 76 74235
rect 16 74199 38 74205
rect 42 74196 76 74200
rect 80 74199 102 74205
rect 42 74166 46 74196
rect 72 74166 76 74196
rect 42 74085 46 74119
rect 72 74085 76 74119
rect -25 74048 25 74050
rect -8 74040 14 74047
rect -8 74039 17 74040
rect 25 74039 27 74048
rect -12 74032 38 74039
rect -12 74031 34 74032
rect -12 74027 8 74031
rect 0 74015 8 74027
rect 14 74015 34 74031
rect 0 74014 34 74015
rect 0 74007 38 74014
rect 14 74006 17 74007
rect 25 73998 27 74007
rect 42 73978 45 74068
rect 69 74053 80 74085
rect 107 74053 143 74081
rect 144 74053 148 74273
rect 332 74205 336 74273
rect 380 74243 462 74275
rect 463 74243 472 74277
rect 480 74243 497 74277
rect 378 74235 464 74243
rect 505 74235 507 74285
rect 514 74243 548 74277
rect 565 74243 582 74277
rect 607 74235 609 74285
rect 404 74219 438 74235
rect 400 74205 442 74206
rect 378 74199 404 74205
rect 442 74199 464 74205
rect 400 74198 404 74199
rect 174 74159 246 74167
rect 295 74164 300 74198
rect 324 74164 329 74198
rect 224 74129 226 74145
rect 196 74121 226 74129
rect 332 74127 336 74195
rect 367 74164 438 74198
rect 400 74157 404 74164
rect 454 74151 504 74153
rect 494 74147 548 74151
rect 494 74142 514 74147
rect 504 74127 506 74142
rect 196 74117 232 74121
rect 196 74087 204 74117
rect 216 74087 232 74117
rect 400 74119 404 74127
rect 107 74047 119 74053
rect 109 74019 119 74047
rect 129 74019 149 74053
rect 174 74049 181 74079
rect 224 74040 226 74087
rect 256 74079 328 74087
rect 332 74085 336 74115
rect 400 74085 408 74119
rect 434 74085 438 74119
rect 498 74117 506 74127
rect 514 74117 515 74137
rect 504 74101 506 74117
rect 525 74108 528 74142
rect 547 74117 548 74137
rect 557 74117 564 74127
rect 514 74101 530 74107
rect 532 74101 548 74107
rect 278 74049 305 74060
rect 42 73927 46 73961
rect 72 73927 76 73961
rect 38 73889 80 73890
rect 42 73848 76 73882
rect 79 73848 113 73882
rect 42 73769 46 73803
rect 72 73769 76 73803
rect -25 73732 25 73734
rect -8 73724 14 73731
rect -8 73723 17 73724
rect 25 73723 27 73732
rect -12 73716 38 73723
rect -12 73715 34 73716
rect -12 73711 8 73715
rect 0 73699 8 73711
rect 14 73699 34 73715
rect 0 73698 34 73699
rect 0 73691 38 73698
rect 14 73690 17 73691
rect 25 73682 27 73691
rect 42 73662 45 73752
rect 71 73721 80 73749
rect 69 73683 80 73721
rect 144 73711 148 74019
rect 196 74006 204 74040
rect 216 74006 232 74040
rect 244 74036 257 74040
rect 300 74036 308 74049
rect 332 74047 342 74085
rect 400 74077 404 74085
rect 336 74037 342 74047
rect 244 74012 291 74036
rect 244 74006 257 74012
rect 224 73959 226 74006
rect 278 74002 291 74012
rect 300 74012 329 74036
rect 332 74027 342 74037
rect 400 74037 409 74065
rect 562 74048 612 74050
rect 466 74039 497 74047
rect 565 74039 596 74047
rect 300 74002 321 74012
rect 300 73996 308 74002
rect 289 73986 308 73996
rect 196 73929 204 73959
rect 216 73929 232 73959
rect 196 73925 232 73929
rect 196 73917 226 73925
rect 300 73917 308 73986
rect 332 73993 351 74027
rect 361 73999 381 74027
rect 361 73993 375 73999
rect 400 73993 411 74037
rect 442 74032 500 74039
rect 466 74031 500 74032
rect 565 74031 599 74039
rect 497 74015 500 74031
rect 596 74015 599 74031
rect 466 74014 500 74015
rect 442 74007 500 74014
rect 565 74007 599 74015
rect 612 73998 614 74048
rect 332 73969 342 73993
rect 336 73957 342 73969
rect 224 73901 226 73917
rect 332 73889 342 73957
rect 400 73961 404 73969
rect 400 73927 408 73961
rect 434 73927 438 73961
rect 454 73945 504 73947
rect 504 73929 506 73945
rect 514 73939 530 73945
rect 532 73939 548 73945
rect 525 73929 548 73938
rect 400 73919 404 73927
rect 498 73919 506 73929
rect 504 73895 506 73919
rect 514 73909 515 73929
rect 525 73904 528 73929
rect 547 73909 548 73929
rect 557 73919 564 73929
rect 514 73895 548 73899
rect 151 73848 156 73882
rect 174 73879 246 73887
rect 256 73879 328 73887
rect 336 73881 342 73889
rect 400 73884 404 73889
rect 180 73851 185 73879
rect 174 73843 246 73851
rect 256 73843 328 73851
rect 332 73849 336 73879
rect 400 73850 438 73884
rect 224 73813 226 73829
rect 196 73805 226 73813
rect 196 73801 232 73805
rect 196 73771 204 73801
rect 216 73771 232 73801
rect 224 73724 226 73771
rect 300 73744 308 73813
rect 332 73811 342 73849
rect 400 73841 404 73850
rect 454 73835 504 73837
rect 494 73831 548 73835
rect 494 73826 514 73831
rect 504 73811 506 73826
rect 336 73799 342 73811
rect 289 73734 308 73744
rect 300 73728 308 73734
rect 332 73765 342 73799
rect 400 73803 404 73811
rect 400 73769 408 73803
rect 434 73769 438 73803
rect 498 73801 506 73811
rect 514 73801 515 73821
rect 504 73785 506 73801
rect 525 73792 528 73826
rect 547 73801 548 73821
rect 557 73801 564 73811
rect 514 73785 530 73791
rect 532 73785 548 73791
rect 332 73737 373 73765
rect 332 73731 351 73737
rect 107 73677 119 73711
rect 129 73677 149 73711
rect 196 73690 204 73724
rect 216 73690 232 73724
rect 244 73718 257 73724
rect 278 73718 291 73728
rect 244 73694 291 73718
rect 300 73718 321 73728
rect 336 73721 351 73731
rect 300 73694 329 73718
rect 332 73703 351 73721
rect 361 73731 375 73737
rect 400 73731 411 73769
rect 562 73732 612 73734
rect 361 73703 381 73731
rect 400 73703 409 73731
rect 466 73723 497 73731
rect 565 73723 596 73731
rect 442 73716 500 73723
rect 466 73715 500 73716
rect 565 73715 599 73723
rect 244 73690 257 73694
rect 42 73611 46 73645
rect 72 73611 76 73645
rect 42 73564 76 73568
rect 42 73549 46 73564
rect 72 73549 76 73564
rect 38 73531 80 73549
rect 16 73525 102 73531
rect 144 73525 148 73677
rect 174 73653 181 73681
rect 224 73643 226 73690
rect 300 73681 308 73694
rect 278 73670 305 73681
rect 332 73653 342 73703
rect 400 73683 404 73703
rect 497 73699 500 73715
rect 596 73699 599 73715
rect 466 73698 500 73699
rect 442 73691 500 73698
rect 565 73691 599 73699
rect 612 73682 614 73732
rect 256 73643 328 73651
rect 336 73645 342 73653
rect 400 73645 404 73653
rect 196 73613 204 73643
rect 216 73613 232 73643
rect 196 73609 232 73613
rect 196 73601 226 73609
rect 224 73585 226 73601
rect 332 73573 336 73641
rect 400 73611 408 73645
rect 434 73611 438 73645
rect 454 73629 504 73631
rect 504 73613 506 73629
rect 514 73623 530 73629
rect 532 73623 548 73629
rect 525 73613 548 73622
rect 400 73603 404 73611
rect 498 73603 506 73613
rect 504 73579 506 73603
rect 514 73593 515 73613
rect 525 73588 528 73613
rect 547 73593 548 73613
rect 557 73603 564 73613
rect 514 73579 548 73583
rect 400 73573 442 73574
rect 174 73563 246 73571
rect 400 73566 404 73573
rect 295 73532 300 73566
rect 324 73532 329 73566
rect 367 73549 438 73566
rect 367 73532 442 73549
rect 400 73531 442 73532
rect 378 73525 464 73531
rect 38 73509 80 73525
rect 400 73509 442 73525
rect -25 73495 25 73497
rect 42 73495 76 73509
rect 404 73495 438 73509
rect 455 73495 505 73497
rect 557 73495 607 73497
rect 16 73487 102 73495
rect 378 73487 464 73495
rect 8 73453 17 73487
rect 18 73485 51 73487
rect 80 73485 100 73487
rect 18 73453 100 73485
rect 380 73485 404 73487
rect 429 73485 438 73487
rect 442 73485 462 73487
rect 16 73445 102 73453
rect 42 73429 76 73445
rect 16 73409 38 73415
rect 42 73406 76 73410
rect 80 73409 102 73415
rect 42 73376 46 73406
rect 72 73376 76 73406
rect 42 73295 46 73329
rect 72 73295 76 73329
rect -25 73258 25 73260
rect -8 73250 14 73257
rect -8 73249 17 73250
rect 25 73249 27 73258
rect -12 73242 38 73249
rect -12 73241 34 73242
rect -12 73237 8 73241
rect 0 73225 8 73237
rect 14 73225 34 73241
rect 0 73224 34 73225
rect 0 73217 38 73224
rect 14 73216 17 73217
rect 25 73208 27 73217
rect 42 73188 45 73278
rect 69 73263 80 73295
rect 107 73263 143 73291
rect 144 73263 148 73483
rect 332 73415 336 73483
rect 380 73453 462 73485
rect 463 73453 472 73487
rect 480 73453 497 73487
rect 378 73445 464 73453
rect 505 73445 507 73495
rect 514 73453 548 73487
rect 565 73453 582 73487
rect 607 73445 609 73495
rect 404 73429 438 73445
rect 400 73415 442 73416
rect 378 73409 404 73415
rect 442 73409 464 73415
rect 400 73408 404 73409
rect 174 73369 246 73377
rect 295 73374 300 73408
rect 324 73374 329 73408
rect 224 73339 226 73355
rect 196 73331 226 73339
rect 332 73337 336 73405
rect 367 73374 438 73408
rect 400 73367 404 73374
rect 454 73361 504 73363
rect 494 73357 548 73361
rect 494 73352 514 73357
rect 504 73337 506 73352
rect 196 73327 232 73331
rect 196 73297 204 73327
rect 216 73297 232 73327
rect 400 73329 404 73337
rect 107 73257 119 73263
rect 109 73229 119 73257
rect 129 73229 149 73263
rect 174 73259 181 73289
rect 224 73250 226 73297
rect 256 73289 328 73297
rect 332 73295 336 73325
rect 400 73295 408 73329
rect 434 73295 438 73329
rect 498 73327 506 73337
rect 514 73327 515 73347
rect 504 73311 506 73327
rect 525 73318 528 73352
rect 547 73327 548 73347
rect 557 73327 564 73337
rect 514 73311 530 73317
rect 532 73311 548 73317
rect 278 73259 305 73270
rect 42 73137 46 73171
rect 72 73137 76 73171
rect 38 73099 80 73100
rect 42 73058 76 73092
rect 79 73058 113 73092
rect 42 72979 46 73013
rect 72 72979 76 73013
rect -25 72942 25 72944
rect -8 72934 14 72941
rect -8 72933 17 72934
rect 25 72933 27 72942
rect -12 72926 38 72933
rect -12 72925 34 72926
rect -12 72921 8 72925
rect 0 72909 8 72921
rect 14 72909 34 72925
rect 0 72908 34 72909
rect 0 72901 38 72908
rect 14 72900 17 72901
rect 25 72892 27 72901
rect 42 72872 45 72962
rect 71 72931 80 72959
rect 69 72893 80 72931
rect 144 72921 148 73229
rect 196 73216 204 73250
rect 216 73216 232 73250
rect 244 73246 257 73250
rect 300 73246 308 73259
rect 332 73257 342 73295
rect 400 73287 404 73295
rect 336 73247 342 73257
rect 244 73222 291 73246
rect 244 73216 257 73222
rect 224 73169 226 73216
rect 278 73212 291 73222
rect 300 73222 329 73246
rect 332 73237 342 73247
rect 400 73247 409 73275
rect 562 73258 612 73260
rect 466 73249 497 73257
rect 565 73249 596 73257
rect 300 73212 321 73222
rect 300 73206 308 73212
rect 289 73196 308 73206
rect 196 73139 204 73169
rect 216 73139 232 73169
rect 196 73135 232 73139
rect 196 73127 226 73135
rect 300 73127 308 73196
rect 332 73203 351 73237
rect 361 73209 381 73237
rect 361 73203 375 73209
rect 400 73203 411 73247
rect 442 73242 500 73249
rect 466 73241 500 73242
rect 565 73241 599 73249
rect 497 73225 500 73241
rect 596 73225 599 73241
rect 466 73224 500 73225
rect 442 73217 500 73224
rect 565 73217 599 73225
rect 612 73208 614 73258
rect 332 73179 342 73203
rect 336 73167 342 73179
rect 224 73111 226 73127
rect 332 73099 342 73167
rect 400 73171 404 73179
rect 400 73137 408 73171
rect 434 73137 438 73171
rect 454 73155 504 73157
rect 504 73139 506 73155
rect 514 73149 530 73155
rect 532 73149 548 73155
rect 525 73139 548 73148
rect 400 73129 404 73137
rect 498 73129 506 73139
rect 504 73105 506 73129
rect 514 73119 515 73139
rect 525 73114 528 73139
rect 547 73119 548 73139
rect 557 73129 564 73139
rect 514 73105 548 73109
rect 151 73058 156 73092
rect 174 73089 246 73097
rect 256 73089 328 73097
rect 336 73091 342 73099
rect 400 73094 404 73099
rect 180 73061 185 73089
rect 174 73053 246 73061
rect 256 73053 328 73061
rect 332 73059 336 73089
rect 400 73060 438 73094
rect 224 73023 226 73039
rect 196 73015 226 73023
rect 196 73011 232 73015
rect 196 72981 204 73011
rect 216 72981 232 73011
rect 224 72934 226 72981
rect 300 72954 308 73023
rect 332 73021 342 73059
rect 400 73051 404 73060
rect 454 73045 504 73047
rect 494 73041 548 73045
rect 494 73036 514 73041
rect 504 73021 506 73036
rect 336 73009 342 73021
rect 289 72944 308 72954
rect 300 72938 308 72944
rect 332 72975 342 73009
rect 400 73013 404 73021
rect 400 72979 408 73013
rect 434 72979 438 73013
rect 498 73011 506 73021
rect 514 73011 515 73031
rect 504 72995 506 73011
rect 525 73002 528 73036
rect 547 73011 548 73031
rect 557 73011 564 73021
rect 514 72995 530 73001
rect 532 72995 548 73001
rect 332 72947 373 72975
rect 332 72941 351 72947
rect 107 72887 119 72921
rect 129 72887 149 72921
rect 196 72900 204 72934
rect 216 72900 232 72934
rect 244 72928 257 72934
rect 278 72928 291 72938
rect 244 72904 291 72928
rect 300 72928 321 72938
rect 336 72931 351 72941
rect 300 72904 329 72928
rect 332 72913 351 72931
rect 361 72941 375 72947
rect 400 72941 411 72979
rect 562 72942 612 72944
rect 361 72913 381 72941
rect 400 72913 409 72941
rect 466 72933 497 72941
rect 565 72933 596 72941
rect 442 72926 500 72933
rect 466 72925 500 72926
rect 565 72925 599 72933
rect 244 72900 257 72904
rect 42 72821 46 72855
rect 72 72821 76 72855
rect 42 72774 76 72778
rect 42 72759 46 72774
rect 72 72759 76 72774
rect 38 72741 80 72759
rect 16 72735 102 72741
rect 144 72735 148 72887
rect 174 72863 181 72891
rect 224 72853 226 72900
rect 300 72891 308 72904
rect 278 72880 305 72891
rect 332 72863 342 72913
rect 400 72893 404 72913
rect 497 72909 500 72925
rect 596 72909 599 72925
rect 466 72908 500 72909
rect 442 72901 500 72908
rect 565 72901 599 72909
rect 612 72892 614 72942
rect 256 72853 328 72861
rect 336 72855 342 72863
rect 400 72855 404 72863
rect 196 72823 204 72853
rect 216 72823 232 72853
rect 196 72819 232 72823
rect 196 72811 226 72819
rect 224 72795 226 72811
rect 332 72783 336 72851
rect 400 72821 408 72855
rect 434 72821 438 72855
rect 454 72839 504 72841
rect 504 72823 506 72839
rect 514 72833 530 72839
rect 532 72833 548 72839
rect 525 72823 548 72832
rect 400 72813 404 72821
rect 498 72813 506 72823
rect 504 72789 506 72813
rect 514 72803 515 72823
rect 525 72798 528 72823
rect 547 72803 548 72823
rect 557 72813 564 72823
rect 514 72789 548 72793
rect 400 72783 442 72784
rect 174 72773 246 72781
rect 400 72776 404 72783
rect 295 72742 300 72776
rect 324 72742 329 72776
rect 367 72759 438 72776
rect 367 72742 442 72759
rect 400 72741 442 72742
rect 378 72735 464 72741
rect 38 72719 80 72735
rect 400 72719 442 72735
rect -25 72705 25 72707
rect 42 72705 76 72719
rect 404 72705 438 72719
rect 455 72705 505 72707
rect 557 72705 607 72707
rect 16 72697 102 72705
rect 378 72697 464 72705
rect 8 72663 17 72697
rect 18 72695 51 72697
rect 80 72695 100 72697
rect 18 72663 100 72695
rect 380 72695 404 72697
rect 429 72695 438 72697
rect 442 72695 462 72697
rect 16 72655 102 72663
rect 42 72639 76 72655
rect 16 72619 38 72625
rect 42 72616 76 72620
rect 80 72619 102 72625
rect 42 72586 46 72616
rect 72 72586 76 72616
rect 42 72505 46 72539
rect 72 72505 76 72539
rect -25 72468 25 72470
rect -8 72460 14 72467
rect -8 72459 17 72460
rect 25 72459 27 72468
rect -12 72452 38 72459
rect -12 72451 34 72452
rect -12 72447 8 72451
rect 0 72435 8 72447
rect 14 72435 34 72451
rect 0 72434 34 72435
rect 0 72427 38 72434
rect 14 72426 17 72427
rect 25 72418 27 72427
rect 42 72398 45 72488
rect 69 72473 80 72505
rect 107 72473 143 72501
rect 144 72473 148 72693
rect 332 72625 336 72693
rect 380 72663 462 72695
rect 463 72663 472 72697
rect 480 72663 497 72697
rect 378 72655 464 72663
rect 505 72655 507 72705
rect 514 72663 548 72697
rect 565 72663 582 72697
rect 607 72655 609 72705
rect 404 72639 438 72655
rect 400 72625 442 72626
rect 378 72619 404 72625
rect 442 72619 464 72625
rect 400 72618 404 72619
rect 174 72579 246 72587
rect 295 72584 300 72618
rect 324 72584 329 72618
rect 224 72549 226 72565
rect 196 72541 226 72549
rect 332 72547 336 72615
rect 367 72584 438 72618
rect 400 72577 404 72584
rect 454 72571 504 72573
rect 494 72567 548 72571
rect 494 72562 514 72567
rect 504 72547 506 72562
rect 196 72537 232 72541
rect 196 72507 204 72537
rect 216 72507 232 72537
rect 400 72539 404 72547
rect 107 72467 119 72473
rect 109 72439 119 72467
rect 129 72439 149 72473
rect 174 72469 181 72499
rect 224 72460 226 72507
rect 256 72499 328 72507
rect 332 72505 336 72535
rect 400 72505 408 72539
rect 434 72505 438 72539
rect 498 72537 506 72547
rect 514 72537 515 72557
rect 504 72521 506 72537
rect 525 72528 528 72562
rect 547 72537 548 72557
rect 557 72537 564 72547
rect 514 72521 530 72527
rect 532 72521 548 72527
rect 278 72469 305 72480
rect 42 72347 46 72381
rect 72 72347 76 72381
rect 38 72309 80 72310
rect 42 72268 76 72302
rect 79 72268 113 72302
rect 42 72189 46 72223
rect 72 72189 76 72223
rect -25 72152 25 72154
rect -8 72144 14 72151
rect -8 72143 17 72144
rect 25 72143 27 72152
rect -12 72136 38 72143
rect -12 72135 34 72136
rect -12 72131 8 72135
rect 0 72119 8 72131
rect 14 72119 34 72135
rect 0 72118 34 72119
rect 0 72111 38 72118
rect 14 72110 17 72111
rect 25 72102 27 72111
rect 42 72082 45 72172
rect 71 72141 80 72169
rect 69 72103 80 72141
rect 144 72131 148 72439
rect 196 72426 204 72460
rect 216 72426 232 72460
rect 244 72456 257 72460
rect 300 72456 308 72469
rect 332 72467 342 72505
rect 400 72497 404 72505
rect 336 72457 342 72467
rect 244 72432 291 72456
rect 244 72426 257 72432
rect 224 72379 226 72426
rect 278 72422 291 72432
rect 300 72432 329 72456
rect 332 72447 342 72457
rect 400 72457 409 72485
rect 562 72468 612 72470
rect 466 72459 497 72467
rect 565 72459 596 72467
rect 300 72422 321 72432
rect 300 72416 308 72422
rect 289 72406 308 72416
rect 196 72349 204 72379
rect 216 72349 232 72379
rect 196 72345 232 72349
rect 196 72337 226 72345
rect 300 72337 308 72406
rect 332 72413 351 72447
rect 361 72419 381 72447
rect 361 72413 375 72419
rect 400 72413 411 72457
rect 442 72452 500 72459
rect 466 72451 500 72452
rect 565 72451 599 72459
rect 497 72435 500 72451
rect 596 72435 599 72451
rect 466 72434 500 72435
rect 442 72427 500 72434
rect 565 72427 599 72435
rect 612 72418 614 72468
rect 332 72389 342 72413
rect 336 72377 342 72389
rect 224 72321 226 72337
rect 332 72309 342 72377
rect 400 72381 404 72389
rect 400 72347 408 72381
rect 434 72347 438 72381
rect 454 72365 504 72367
rect 504 72349 506 72365
rect 514 72359 530 72365
rect 532 72359 548 72365
rect 525 72349 548 72358
rect 400 72339 404 72347
rect 498 72339 506 72349
rect 504 72315 506 72339
rect 514 72329 515 72349
rect 525 72324 528 72349
rect 547 72329 548 72349
rect 557 72339 564 72349
rect 514 72315 548 72319
rect 151 72268 156 72302
rect 174 72299 246 72307
rect 256 72299 328 72307
rect 336 72301 342 72309
rect 400 72304 404 72309
rect 180 72271 185 72299
rect 174 72263 246 72271
rect 256 72263 328 72271
rect 332 72269 336 72299
rect 400 72270 438 72304
rect 224 72233 226 72249
rect 196 72225 226 72233
rect 196 72221 232 72225
rect 196 72191 204 72221
rect 216 72191 232 72221
rect 224 72144 226 72191
rect 300 72164 308 72233
rect 332 72231 342 72269
rect 400 72261 404 72270
rect 454 72255 504 72257
rect 494 72251 548 72255
rect 494 72246 514 72251
rect 504 72231 506 72246
rect 336 72219 342 72231
rect 289 72154 308 72164
rect 300 72148 308 72154
rect 332 72185 342 72219
rect 400 72223 404 72231
rect 400 72189 408 72223
rect 434 72189 438 72223
rect 498 72221 506 72231
rect 514 72221 515 72241
rect 504 72205 506 72221
rect 525 72212 528 72246
rect 547 72221 548 72241
rect 557 72221 564 72231
rect 514 72205 530 72211
rect 532 72205 548 72211
rect 332 72157 373 72185
rect 332 72151 351 72157
rect 107 72097 119 72131
rect 129 72097 149 72131
rect 196 72110 204 72144
rect 216 72110 232 72144
rect 244 72138 257 72144
rect 278 72138 291 72148
rect 244 72114 291 72138
rect 300 72138 321 72148
rect 336 72141 351 72151
rect 300 72114 329 72138
rect 332 72123 351 72141
rect 361 72151 375 72157
rect 400 72151 411 72189
rect 562 72152 612 72154
rect 361 72123 381 72151
rect 400 72123 409 72151
rect 466 72143 497 72151
rect 565 72143 596 72151
rect 442 72136 500 72143
rect 466 72135 500 72136
rect 565 72135 599 72143
rect 244 72110 257 72114
rect 42 72031 46 72065
rect 72 72031 76 72065
rect 42 71984 76 71988
rect 42 71969 46 71984
rect 72 71969 76 71984
rect 38 71951 80 71969
rect 16 71945 102 71951
rect 144 71945 148 72097
rect 174 72073 181 72101
rect 224 72063 226 72110
rect 300 72101 308 72114
rect 278 72090 305 72101
rect 332 72073 342 72123
rect 400 72103 404 72123
rect 497 72119 500 72135
rect 596 72119 599 72135
rect 466 72118 500 72119
rect 442 72111 500 72118
rect 565 72111 599 72119
rect 612 72102 614 72152
rect 256 72063 328 72071
rect 336 72065 342 72073
rect 400 72065 404 72073
rect 196 72033 204 72063
rect 216 72033 232 72063
rect 196 72029 232 72033
rect 196 72021 226 72029
rect 224 72005 226 72021
rect 332 71993 336 72061
rect 400 72031 408 72065
rect 434 72031 438 72065
rect 454 72049 504 72051
rect 504 72033 506 72049
rect 514 72043 530 72049
rect 532 72043 548 72049
rect 525 72033 548 72042
rect 400 72023 404 72031
rect 498 72023 506 72033
rect 504 71999 506 72023
rect 514 72013 515 72033
rect 525 72008 528 72033
rect 547 72013 548 72033
rect 557 72023 564 72033
rect 514 71999 548 72003
rect 400 71993 442 71994
rect 174 71983 246 71991
rect 400 71986 404 71993
rect 295 71952 300 71986
rect 324 71952 329 71986
rect 367 71969 438 71986
rect 367 71952 442 71969
rect 400 71951 442 71952
rect 378 71945 464 71951
rect 38 71929 80 71945
rect 400 71929 442 71945
rect -25 71915 25 71917
rect 42 71915 76 71929
rect 404 71915 438 71929
rect 455 71915 505 71917
rect 557 71915 607 71917
rect 16 71907 102 71915
rect 378 71907 464 71915
rect 8 71873 17 71907
rect 18 71905 51 71907
rect 80 71905 100 71907
rect 18 71873 100 71905
rect 380 71905 404 71907
rect 429 71905 438 71907
rect 442 71905 462 71907
rect 16 71865 102 71873
rect 42 71849 76 71865
rect 16 71829 38 71835
rect 42 71826 76 71830
rect 80 71829 102 71835
rect 42 71796 46 71826
rect 72 71796 76 71826
rect 42 71715 46 71749
rect 72 71715 76 71749
rect -25 71678 25 71680
rect -8 71670 14 71677
rect -8 71669 17 71670
rect 25 71669 27 71678
rect -12 71662 38 71669
rect -12 71661 34 71662
rect -12 71657 8 71661
rect 0 71645 8 71657
rect 14 71645 34 71661
rect 0 71644 34 71645
rect 0 71637 38 71644
rect 14 71636 17 71637
rect 25 71628 27 71637
rect 42 71608 45 71698
rect 69 71683 80 71715
rect 107 71683 143 71711
rect 144 71683 148 71903
rect 332 71835 336 71903
rect 380 71873 462 71905
rect 463 71873 472 71907
rect 480 71873 497 71907
rect 378 71865 464 71873
rect 505 71865 507 71915
rect 514 71873 548 71907
rect 565 71873 582 71907
rect 607 71865 609 71915
rect 404 71849 438 71865
rect 400 71835 442 71836
rect 378 71829 404 71835
rect 442 71829 464 71835
rect 400 71828 404 71829
rect 174 71789 246 71797
rect 295 71794 300 71828
rect 324 71794 329 71828
rect 224 71759 226 71775
rect 196 71751 226 71759
rect 332 71757 336 71825
rect 367 71794 438 71828
rect 400 71787 404 71794
rect 454 71781 504 71783
rect 494 71777 548 71781
rect 494 71772 514 71777
rect 504 71757 506 71772
rect 196 71747 232 71751
rect 196 71717 204 71747
rect 216 71717 232 71747
rect 400 71749 404 71757
rect 107 71677 119 71683
rect 109 71649 119 71677
rect 129 71649 149 71683
rect 174 71679 181 71709
rect 224 71670 226 71717
rect 256 71709 328 71717
rect 332 71715 336 71745
rect 400 71715 408 71749
rect 434 71715 438 71749
rect 498 71747 506 71757
rect 514 71747 515 71767
rect 504 71731 506 71747
rect 525 71738 528 71772
rect 547 71747 548 71767
rect 557 71747 564 71757
rect 514 71731 530 71737
rect 532 71731 548 71737
rect 278 71679 305 71690
rect 42 71557 46 71591
rect 72 71557 76 71591
rect 38 71519 80 71520
rect 42 71478 76 71512
rect 79 71478 113 71512
rect 42 71399 46 71433
rect 72 71399 76 71433
rect -25 71362 25 71364
rect -8 71354 14 71361
rect -8 71353 17 71354
rect 25 71353 27 71362
rect -12 71346 38 71353
rect -12 71345 34 71346
rect -12 71341 8 71345
rect 0 71329 8 71341
rect 14 71329 34 71345
rect 0 71328 34 71329
rect 0 71321 38 71328
rect 14 71320 17 71321
rect 25 71312 27 71321
rect 42 71292 45 71382
rect 71 71351 80 71379
rect 69 71313 80 71351
rect 144 71341 148 71649
rect 196 71636 204 71670
rect 216 71636 232 71670
rect 244 71666 257 71670
rect 300 71666 308 71679
rect 332 71677 342 71715
rect 400 71707 404 71715
rect 336 71667 342 71677
rect 244 71642 291 71666
rect 244 71636 257 71642
rect 224 71589 226 71636
rect 278 71632 291 71642
rect 300 71642 329 71666
rect 332 71657 342 71667
rect 400 71667 409 71695
rect 562 71678 612 71680
rect 466 71669 497 71677
rect 565 71669 596 71677
rect 300 71632 321 71642
rect 300 71626 308 71632
rect 289 71616 308 71626
rect 196 71559 204 71589
rect 216 71559 232 71589
rect 196 71555 232 71559
rect 196 71547 226 71555
rect 300 71547 308 71616
rect 332 71623 351 71657
rect 361 71629 381 71657
rect 361 71623 375 71629
rect 400 71623 411 71667
rect 442 71662 500 71669
rect 466 71661 500 71662
rect 565 71661 599 71669
rect 497 71645 500 71661
rect 596 71645 599 71661
rect 466 71644 500 71645
rect 442 71637 500 71644
rect 565 71637 599 71645
rect 612 71628 614 71678
rect 332 71599 342 71623
rect 336 71587 342 71599
rect 224 71531 226 71547
rect 332 71519 342 71587
rect 400 71591 404 71599
rect 400 71557 408 71591
rect 434 71557 438 71591
rect 454 71575 504 71577
rect 504 71559 506 71575
rect 514 71569 530 71575
rect 532 71569 548 71575
rect 525 71559 548 71568
rect 400 71549 404 71557
rect 498 71549 506 71559
rect 504 71525 506 71549
rect 514 71539 515 71559
rect 525 71534 528 71559
rect 547 71539 548 71559
rect 557 71549 564 71559
rect 514 71525 548 71529
rect 151 71478 156 71512
rect 174 71509 246 71517
rect 256 71509 328 71517
rect 336 71511 342 71519
rect 400 71514 404 71519
rect 180 71481 185 71509
rect 174 71473 246 71481
rect 256 71473 328 71481
rect 332 71479 336 71509
rect 400 71480 438 71514
rect 224 71443 226 71459
rect 196 71435 226 71443
rect 196 71431 232 71435
rect 196 71401 204 71431
rect 216 71401 232 71431
rect 224 71354 226 71401
rect 300 71374 308 71443
rect 332 71441 342 71479
rect 400 71471 404 71480
rect 454 71465 504 71467
rect 494 71461 548 71465
rect 494 71456 514 71461
rect 504 71441 506 71456
rect 336 71429 342 71441
rect 289 71364 308 71374
rect 300 71358 308 71364
rect 332 71395 342 71429
rect 400 71433 404 71441
rect 400 71399 408 71433
rect 434 71399 438 71433
rect 498 71431 506 71441
rect 514 71431 515 71451
rect 504 71415 506 71431
rect 525 71422 528 71456
rect 547 71431 548 71451
rect 557 71431 564 71441
rect 514 71415 530 71421
rect 532 71415 548 71421
rect 332 71367 373 71395
rect 332 71361 351 71367
rect 107 71307 119 71341
rect 129 71307 149 71341
rect 196 71320 204 71354
rect 216 71320 232 71354
rect 244 71348 257 71354
rect 278 71348 291 71358
rect 244 71324 291 71348
rect 300 71348 321 71358
rect 336 71351 351 71361
rect 300 71324 329 71348
rect 332 71333 351 71351
rect 361 71361 375 71367
rect 400 71361 411 71399
rect 562 71362 612 71364
rect 361 71333 381 71361
rect 400 71333 409 71361
rect 466 71353 497 71361
rect 565 71353 596 71361
rect 442 71346 500 71353
rect 466 71345 500 71346
rect 565 71345 599 71353
rect 244 71320 257 71324
rect 42 71241 46 71275
rect 72 71241 76 71275
rect 42 71194 76 71198
rect 42 71179 46 71194
rect 72 71179 76 71194
rect 38 71161 80 71179
rect 16 71155 102 71161
rect 144 71155 148 71307
rect 174 71283 181 71311
rect 224 71273 226 71320
rect 300 71311 308 71324
rect 278 71300 305 71311
rect 332 71283 342 71333
rect 400 71313 404 71333
rect 497 71329 500 71345
rect 596 71329 599 71345
rect 466 71328 500 71329
rect 442 71321 500 71328
rect 565 71321 599 71329
rect 612 71312 614 71362
rect 256 71273 328 71281
rect 336 71275 342 71283
rect 400 71275 404 71283
rect 196 71243 204 71273
rect 216 71243 232 71273
rect 196 71239 232 71243
rect 196 71231 226 71239
rect 224 71215 226 71231
rect 332 71203 336 71271
rect 400 71241 408 71275
rect 434 71241 438 71275
rect 454 71259 504 71261
rect 504 71243 506 71259
rect 514 71253 530 71259
rect 532 71253 548 71259
rect 525 71243 548 71252
rect 400 71233 404 71241
rect 498 71233 506 71243
rect 504 71209 506 71233
rect 514 71223 515 71243
rect 525 71218 528 71243
rect 547 71223 548 71243
rect 557 71233 564 71243
rect 514 71209 548 71213
rect 400 71203 442 71204
rect 174 71193 246 71201
rect 400 71196 404 71203
rect 295 71162 300 71196
rect 324 71162 329 71196
rect 367 71179 438 71196
rect 367 71162 442 71179
rect 400 71161 442 71162
rect 378 71155 464 71161
rect 38 71139 80 71155
rect 400 71139 442 71155
rect -25 71125 25 71127
rect 42 71125 76 71139
rect 404 71125 438 71139
rect 455 71125 505 71127
rect 557 71125 607 71127
rect 16 71117 102 71125
rect 378 71117 464 71125
rect 8 71083 17 71117
rect 18 71115 51 71117
rect 80 71115 100 71117
rect 18 71083 100 71115
rect 380 71115 404 71117
rect 429 71115 438 71117
rect 442 71115 462 71117
rect 16 71075 102 71083
rect 42 71059 76 71075
rect 16 71039 38 71045
rect 42 71036 76 71040
rect 80 71039 102 71045
rect 42 71006 46 71036
rect 72 71006 76 71036
rect 42 70925 46 70959
rect 72 70925 76 70959
rect -25 70888 25 70890
rect -8 70880 14 70887
rect -8 70879 17 70880
rect 25 70879 27 70888
rect -12 70872 38 70879
rect -12 70871 34 70872
rect -12 70867 8 70871
rect 0 70855 8 70867
rect 14 70855 34 70871
rect 0 70854 34 70855
rect 0 70847 38 70854
rect 14 70846 17 70847
rect 25 70838 27 70847
rect 42 70818 45 70908
rect 69 70893 80 70925
rect 107 70893 143 70921
rect 144 70893 148 71113
rect 332 71045 336 71113
rect 380 71083 462 71115
rect 463 71083 472 71117
rect 480 71083 497 71117
rect 378 71075 464 71083
rect 505 71075 507 71125
rect 514 71083 548 71117
rect 565 71083 582 71117
rect 607 71075 609 71125
rect 404 71059 438 71075
rect 400 71045 442 71046
rect 378 71039 404 71045
rect 442 71039 464 71045
rect 400 71038 404 71039
rect 174 70999 246 71007
rect 295 71004 300 71038
rect 324 71004 329 71038
rect 224 70969 226 70985
rect 196 70961 226 70969
rect 332 70967 336 71035
rect 367 71004 438 71038
rect 400 70997 404 71004
rect 454 70991 504 70993
rect 494 70987 548 70991
rect 494 70982 514 70987
rect 504 70967 506 70982
rect 196 70957 232 70961
rect 196 70927 204 70957
rect 216 70927 232 70957
rect 400 70959 404 70967
rect 107 70887 119 70893
rect 109 70859 119 70887
rect 129 70859 149 70893
rect 174 70889 181 70919
rect 224 70880 226 70927
rect 256 70919 328 70927
rect 332 70925 336 70955
rect 400 70925 408 70959
rect 434 70925 438 70959
rect 498 70957 506 70967
rect 514 70957 515 70977
rect 504 70941 506 70957
rect 525 70948 528 70982
rect 547 70957 548 70977
rect 557 70957 564 70967
rect 514 70941 530 70947
rect 532 70941 548 70947
rect 278 70889 305 70900
rect 42 70767 46 70801
rect 72 70767 76 70801
rect 38 70729 80 70730
rect 42 70688 76 70722
rect 79 70688 113 70722
rect 42 70609 46 70643
rect 72 70609 76 70643
rect -25 70572 25 70574
rect -8 70564 14 70571
rect -8 70563 17 70564
rect 25 70563 27 70572
rect -12 70556 38 70563
rect -12 70555 34 70556
rect -12 70551 8 70555
rect 0 70539 8 70551
rect 14 70539 34 70555
rect 0 70538 34 70539
rect 0 70531 38 70538
rect 14 70530 17 70531
rect 25 70522 27 70531
rect 42 70502 45 70592
rect 71 70561 80 70589
rect 69 70523 80 70561
rect 144 70551 148 70859
rect 196 70846 204 70880
rect 216 70846 232 70880
rect 244 70876 257 70880
rect 300 70876 308 70889
rect 332 70887 342 70925
rect 400 70917 404 70925
rect 336 70877 342 70887
rect 244 70852 291 70876
rect 244 70846 257 70852
rect 224 70799 226 70846
rect 278 70842 291 70852
rect 300 70852 329 70876
rect 332 70867 342 70877
rect 400 70877 409 70905
rect 562 70888 612 70890
rect 466 70879 497 70887
rect 565 70879 596 70887
rect 300 70842 321 70852
rect 300 70836 308 70842
rect 289 70826 308 70836
rect 196 70769 204 70799
rect 216 70769 232 70799
rect 196 70765 232 70769
rect 196 70757 226 70765
rect 300 70757 308 70826
rect 332 70833 351 70867
rect 361 70839 381 70867
rect 361 70833 375 70839
rect 400 70833 411 70877
rect 442 70872 500 70879
rect 466 70871 500 70872
rect 565 70871 599 70879
rect 497 70855 500 70871
rect 596 70855 599 70871
rect 466 70854 500 70855
rect 442 70847 500 70854
rect 565 70847 599 70855
rect 612 70838 614 70888
rect 332 70809 342 70833
rect 336 70797 342 70809
rect 224 70741 226 70757
rect 332 70729 342 70797
rect 400 70801 404 70809
rect 400 70767 408 70801
rect 434 70767 438 70801
rect 454 70785 504 70787
rect 504 70769 506 70785
rect 514 70779 530 70785
rect 532 70779 548 70785
rect 525 70769 548 70778
rect 400 70759 404 70767
rect 498 70759 506 70769
rect 504 70735 506 70759
rect 514 70749 515 70769
rect 525 70744 528 70769
rect 547 70749 548 70769
rect 557 70759 564 70769
rect 514 70735 548 70739
rect 151 70688 156 70722
rect 174 70719 246 70727
rect 256 70719 328 70727
rect 336 70721 342 70729
rect 400 70724 404 70729
rect 180 70691 185 70719
rect 174 70683 246 70691
rect 256 70683 328 70691
rect 332 70689 336 70719
rect 400 70690 438 70724
rect 224 70653 226 70669
rect 196 70645 226 70653
rect 196 70641 232 70645
rect 196 70611 204 70641
rect 216 70611 232 70641
rect 224 70564 226 70611
rect 300 70584 308 70653
rect 332 70651 342 70689
rect 400 70681 404 70690
rect 454 70675 504 70677
rect 494 70671 548 70675
rect 494 70666 514 70671
rect 504 70651 506 70666
rect 336 70639 342 70651
rect 289 70574 308 70584
rect 300 70568 308 70574
rect 332 70605 342 70639
rect 400 70643 404 70651
rect 400 70609 408 70643
rect 434 70609 438 70643
rect 498 70641 506 70651
rect 514 70641 515 70661
rect 504 70625 506 70641
rect 525 70632 528 70666
rect 547 70641 548 70661
rect 557 70641 564 70651
rect 514 70625 530 70631
rect 532 70625 548 70631
rect 332 70577 373 70605
rect 332 70571 351 70577
rect 107 70517 119 70551
rect 129 70517 149 70551
rect 196 70530 204 70564
rect 216 70530 232 70564
rect 244 70558 257 70564
rect 278 70558 291 70568
rect 244 70534 291 70558
rect 300 70558 321 70568
rect 336 70561 351 70571
rect 300 70534 329 70558
rect 332 70543 351 70561
rect 361 70571 375 70577
rect 400 70571 411 70609
rect 562 70572 612 70574
rect 361 70543 381 70571
rect 400 70543 409 70571
rect 466 70563 497 70571
rect 565 70563 596 70571
rect 442 70556 500 70563
rect 466 70555 500 70556
rect 565 70555 599 70563
rect 244 70530 257 70534
rect 42 70451 46 70485
rect 72 70451 76 70485
rect 42 70404 76 70408
rect 42 70389 46 70404
rect 72 70389 76 70404
rect 38 70371 80 70389
rect 16 70365 102 70371
rect 144 70365 148 70517
rect 174 70493 181 70521
rect 224 70483 226 70530
rect 300 70521 308 70534
rect 278 70510 305 70521
rect 332 70493 342 70543
rect 400 70523 404 70543
rect 497 70539 500 70555
rect 596 70539 599 70555
rect 466 70538 500 70539
rect 442 70531 500 70538
rect 565 70531 599 70539
rect 612 70522 614 70572
rect 256 70483 328 70491
rect 336 70485 342 70493
rect 400 70485 404 70493
rect 196 70453 204 70483
rect 216 70453 232 70483
rect 196 70449 232 70453
rect 196 70441 226 70449
rect 224 70425 226 70441
rect 332 70413 336 70481
rect 400 70451 408 70485
rect 434 70451 438 70485
rect 454 70469 504 70471
rect 504 70453 506 70469
rect 514 70463 530 70469
rect 532 70463 548 70469
rect 525 70453 548 70462
rect 400 70443 404 70451
rect 498 70443 506 70453
rect 504 70419 506 70443
rect 514 70433 515 70453
rect 525 70428 528 70453
rect 547 70433 548 70453
rect 557 70443 564 70453
rect 514 70419 548 70423
rect 400 70413 442 70414
rect 174 70403 246 70411
rect 400 70406 404 70413
rect 295 70372 300 70406
rect 324 70372 329 70406
rect 367 70389 438 70406
rect 367 70372 442 70389
rect 400 70371 442 70372
rect 378 70365 464 70371
rect 38 70349 80 70365
rect 400 70349 442 70365
rect -25 70335 25 70337
rect 42 70335 76 70349
rect 404 70335 438 70349
rect 455 70335 505 70337
rect 557 70335 607 70337
rect 16 70327 102 70335
rect 378 70327 464 70335
rect 8 70293 17 70327
rect 18 70325 51 70327
rect 80 70325 100 70327
rect 18 70293 100 70325
rect 380 70325 404 70327
rect 429 70325 438 70327
rect 442 70325 462 70327
rect 16 70285 102 70293
rect 42 70269 76 70285
rect 16 70249 38 70255
rect 42 70246 76 70250
rect 80 70249 102 70255
rect 42 70216 46 70246
rect 72 70216 76 70246
rect 42 70135 46 70169
rect 72 70135 76 70169
rect -25 70098 25 70100
rect -8 70090 14 70097
rect -8 70089 17 70090
rect 25 70089 27 70098
rect -12 70082 38 70089
rect -12 70081 34 70082
rect -12 70077 8 70081
rect 0 70065 8 70077
rect 14 70065 34 70081
rect 0 70064 34 70065
rect 0 70057 38 70064
rect 14 70056 17 70057
rect 25 70048 27 70057
rect 42 70028 45 70118
rect 69 70103 80 70135
rect 107 70103 143 70131
rect 144 70103 148 70323
rect 332 70255 336 70323
rect 380 70293 462 70325
rect 463 70293 472 70327
rect 480 70293 497 70327
rect 378 70285 464 70293
rect 505 70285 507 70335
rect 514 70293 548 70327
rect 565 70293 582 70327
rect 607 70285 609 70335
rect 404 70269 438 70285
rect 400 70255 442 70256
rect 378 70249 404 70255
rect 442 70249 464 70255
rect 400 70248 404 70249
rect 174 70209 246 70217
rect 295 70214 300 70248
rect 324 70214 329 70248
rect 224 70179 226 70195
rect 196 70171 226 70179
rect 332 70177 336 70245
rect 367 70214 438 70248
rect 400 70207 404 70214
rect 454 70201 504 70203
rect 494 70197 548 70201
rect 494 70192 514 70197
rect 504 70177 506 70192
rect 196 70167 232 70171
rect 196 70137 204 70167
rect 216 70137 232 70167
rect 400 70169 404 70177
rect 107 70097 119 70103
rect 109 70069 119 70097
rect 129 70069 149 70103
rect 174 70099 181 70129
rect 224 70090 226 70137
rect 256 70129 328 70137
rect 332 70135 336 70165
rect 400 70135 408 70169
rect 434 70135 438 70169
rect 498 70167 506 70177
rect 514 70167 515 70187
rect 504 70151 506 70167
rect 525 70158 528 70192
rect 547 70167 548 70187
rect 557 70167 564 70177
rect 514 70151 530 70157
rect 532 70151 548 70157
rect 278 70099 305 70110
rect 42 69977 46 70011
rect 72 69977 76 70011
rect 38 69939 80 69940
rect 42 69898 76 69932
rect 79 69898 113 69932
rect 42 69819 46 69853
rect 72 69819 76 69853
rect -25 69782 25 69784
rect -8 69774 14 69781
rect -8 69773 17 69774
rect 25 69773 27 69782
rect -12 69766 38 69773
rect -12 69765 34 69766
rect -12 69761 8 69765
rect 0 69749 8 69761
rect 14 69749 34 69765
rect 0 69748 34 69749
rect 0 69741 38 69748
rect 14 69740 17 69741
rect 25 69732 27 69741
rect 42 69712 45 69802
rect 71 69771 80 69799
rect 69 69733 80 69771
rect 144 69761 148 70069
rect 196 70056 204 70090
rect 216 70056 232 70090
rect 244 70086 257 70090
rect 300 70086 308 70099
rect 332 70097 342 70135
rect 400 70127 404 70135
rect 336 70087 342 70097
rect 244 70062 291 70086
rect 244 70056 257 70062
rect 224 70009 226 70056
rect 278 70052 291 70062
rect 300 70062 329 70086
rect 332 70077 342 70087
rect 400 70087 409 70115
rect 562 70098 612 70100
rect 466 70089 497 70097
rect 565 70089 596 70097
rect 300 70052 321 70062
rect 300 70046 308 70052
rect 289 70036 308 70046
rect 196 69979 204 70009
rect 216 69979 232 70009
rect 196 69975 232 69979
rect 196 69967 226 69975
rect 300 69967 308 70036
rect 332 70043 351 70077
rect 361 70049 381 70077
rect 361 70043 375 70049
rect 400 70043 411 70087
rect 442 70082 500 70089
rect 466 70081 500 70082
rect 565 70081 599 70089
rect 497 70065 500 70081
rect 596 70065 599 70081
rect 466 70064 500 70065
rect 442 70057 500 70064
rect 565 70057 599 70065
rect 612 70048 614 70098
rect 332 70019 342 70043
rect 336 70007 342 70019
rect 224 69951 226 69967
rect 332 69939 342 70007
rect 400 70011 404 70019
rect 400 69977 408 70011
rect 434 69977 438 70011
rect 454 69995 504 69997
rect 504 69979 506 69995
rect 514 69989 530 69995
rect 532 69989 548 69995
rect 525 69979 548 69988
rect 400 69969 404 69977
rect 498 69969 506 69979
rect 504 69945 506 69969
rect 514 69959 515 69979
rect 525 69954 528 69979
rect 547 69959 548 69979
rect 557 69969 564 69979
rect 514 69945 548 69949
rect 151 69898 156 69932
rect 174 69929 246 69937
rect 256 69929 328 69937
rect 336 69931 342 69939
rect 400 69934 404 69939
rect 180 69901 185 69929
rect 174 69893 246 69901
rect 256 69893 328 69901
rect 332 69899 336 69929
rect 400 69900 438 69934
rect 224 69863 226 69879
rect 196 69855 226 69863
rect 196 69851 232 69855
rect 196 69821 204 69851
rect 216 69821 232 69851
rect 224 69774 226 69821
rect 300 69794 308 69863
rect 332 69861 342 69899
rect 400 69891 404 69900
rect 454 69885 504 69887
rect 494 69881 548 69885
rect 494 69876 514 69881
rect 504 69861 506 69876
rect 336 69849 342 69861
rect 289 69784 308 69794
rect 300 69778 308 69784
rect 332 69815 342 69849
rect 400 69853 404 69861
rect 400 69819 408 69853
rect 434 69819 438 69853
rect 498 69851 506 69861
rect 514 69851 515 69871
rect 504 69835 506 69851
rect 525 69842 528 69876
rect 547 69851 548 69871
rect 557 69851 564 69861
rect 514 69835 530 69841
rect 532 69835 548 69841
rect 332 69787 373 69815
rect 332 69781 351 69787
rect 107 69727 119 69761
rect 129 69727 149 69761
rect 196 69740 204 69774
rect 216 69740 232 69774
rect 244 69768 257 69774
rect 278 69768 291 69778
rect 244 69744 291 69768
rect 300 69768 321 69778
rect 336 69771 351 69781
rect 300 69744 329 69768
rect 332 69753 351 69771
rect 361 69781 375 69787
rect 400 69781 411 69819
rect 562 69782 612 69784
rect 361 69753 381 69781
rect 400 69753 409 69781
rect 466 69773 497 69781
rect 565 69773 596 69781
rect 442 69766 500 69773
rect 466 69765 500 69766
rect 565 69765 599 69773
rect 244 69740 257 69744
rect 42 69661 46 69695
rect 72 69661 76 69695
rect 42 69614 76 69618
rect 42 69599 46 69614
rect 72 69599 76 69614
rect 38 69581 80 69599
rect 16 69575 102 69581
rect 144 69575 148 69727
rect 174 69703 181 69731
rect 224 69693 226 69740
rect 300 69731 308 69744
rect 278 69720 305 69731
rect 332 69703 342 69753
rect 400 69733 404 69753
rect 497 69749 500 69765
rect 596 69749 599 69765
rect 466 69748 500 69749
rect 442 69741 500 69748
rect 565 69741 599 69749
rect 612 69732 614 69782
rect 256 69693 328 69701
rect 336 69695 342 69703
rect 400 69695 404 69703
rect 196 69663 204 69693
rect 216 69663 232 69693
rect 196 69659 232 69663
rect 196 69651 226 69659
rect 224 69635 226 69651
rect 332 69623 336 69691
rect 400 69661 408 69695
rect 434 69661 438 69695
rect 454 69679 504 69681
rect 504 69663 506 69679
rect 514 69673 530 69679
rect 532 69673 548 69679
rect 525 69663 548 69672
rect 400 69653 404 69661
rect 498 69653 506 69663
rect 504 69629 506 69653
rect 514 69643 515 69663
rect 525 69638 528 69663
rect 547 69643 548 69663
rect 557 69653 564 69663
rect 514 69629 548 69633
rect 400 69623 442 69624
rect 174 69613 246 69621
rect 400 69616 404 69623
rect 295 69582 300 69616
rect 324 69582 329 69616
rect 367 69599 438 69616
rect 367 69582 442 69599
rect 400 69581 442 69582
rect 378 69575 464 69581
rect 38 69559 80 69575
rect 400 69559 442 69575
rect -25 69545 25 69547
rect 42 69545 76 69559
rect 404 69545 438 69559
rect 455 69545 505 69547
rect 557 69545 607 69547
rect 16 69537 102 69545
rect 378 69537 464 69545
rect 8 69503 17 69537
rect 18 69535 51 69537
rect 80 69535 100 69537
rect 18 69503 100 69535
rect 380 69535 404 69537
rect 429 69535 438 69537
rect 442 69535 462 69537
rect 16 69495 102 69503
rect 42 69479 76 69495
rect 16 69459 38 69465
rect 42 69456 76 69460
rect 80 69459 102 69465
rect 42 69426 46 69456
rect 72 69426 76 69456
rect 42 69345 46 69379
rect 72 69345 76 69379
rect -25 69308 25 69310
rect -8 69300 14 69307
rect -8 69299 17 69300
rect 25 69299 27 69308
rect -12 69292 38 69299
rect -12 69291 34 69292
rect -12 69287 8 69291
rect 0 69275 8 69287
rect 14 69275 34 69291
rect 0 69274 34 69275
rect 0 69267 38 69274
rect 14 69266 17 69267
rect 25 69258 27 69267
rect 42 69238 45 69328
rect 69 69313 80 69345
rect 107 69313 143 69341
rect 144 69313 148 69533
rect 332 69465 336 69533
rect 380 69503 462 69535
rect 463 69503 472 69537
rect 480 69503 497 69537
rect 378 69495 464 69503
rect 505 69495 507 69545
rect 514 69503 548 69537
rect 565 69503 582 69537
rect 607 69495 609 69545
rect 404 69479 438 69495
rect 400 69465 442 69466
rect 378 69459 404 69465
rect 442 69459 464 69465
rect 400 69458 404 69459
rect 174 69419 246 69427
rect 295 69424 300 69458
rect 324 69424 329 69458
rect 224 69389 226 69405
rect 196 69381 226 69389
rect 332 69387 336 69455
rect 367 69424 438 69458
rect 400 69417 404 69424
rect 454 69411 504 69413
rect 494 69407 548 69411
rect 494 69402 514 69407
rect 504 69387 506 69402
rect 196 69377 232 69381
rect 196 69347 204 69377
rect 216 69347 232 69377
rect 400 69379 404 69387
rect 107 69307 119 69313
rect 109 69279 119 69307
rect 129 69279 149 69313
rect 174 69309 181 69339
rect 224 69300 226 69347
rect 256 69339 328 69347
rect 332 69345 336 69375
rect 400 69345 408 69379
rect 434 69345 438 69379
rect 498 69377 506 69387
rect 514 69377 515 69397
rect 504 69361 506 69377
rect 525 69368 528 69402
rect 547 69377 548 69397
rect 557 69377 564 69387
rect 514 69361 530 69367
rect 532 69361 548 69367
rect 278 69309 305 69320
rect 42 69187 46 69221
rect 72 69187 76 69221
rect 38 69149 80 69150
rect 42 69108 76 69142
rect 79 69108 113 69142
rect 42 69029 46 69063
rect 72 69029 76 69063
rect -25 68992 25 68994
rect -8 68984 14 68991
rect -8 68983 17 68984
rect 25 68983 27 68992
rect -12 68976 38 68983
rect -12 68975 34 68976
rect -12 68971 8 68975
rect 0 68959 8 68971
rect 14 68959 34 68975
rect 0 68958 34 68959
rect 0 68951 38 68958
rect 14 68950 17 68951
rect 25 68942 27 68951
rect 42 68922 45 69012
rect 71 68981 80 69009
rect 69 68943 80 68981
rect 144 68971 148 69279
rect 196 69266 204 69300
rect 216 69266 232 69300
rect 244 69296 257 69300
rect 300 69296 308 69309
rect 332 69307 342 69345
rect 400 69337 404 69345
rect 336 69297 342 69307
rect 244 69272 291 69296
rect 244 69266 257 69272
rect 224 69219 226 69266
rect 278 69262 291 69272
rect 300 69272 329 69296
rect 332 69287 342 69297
rect 400 69297 409 69325
rect 562 69308 612 69310
rect 466 69299 497 69307
rect 565 69299 596 69307
rect 300 69262 321 69272
rect 300 69256 308 69262
rect 289 69246 308 69256
rect 196 69189 204 69219
rect 216 69189 232 69219
rect 196 69185 232 69189
rect 196 69177 226 69185
rect 300 69177 308 69246
rect 332 69253 351 69287
rect 361 69259 381 69287
rect 361 69253 375 69259
rect 400 69253 411 69297
rect 442 69292 500 69299
rect 466 69291 500 69292
rect 565 69291 599 69299
rect 497 69275 500 69291
rect 596 69275 599 69291
rect 466 69274 500 69275
rect 442 69267 500 69274
rect 565 69267 599 69275
rect 612 69258 614 69308
rect 332 69229 342 69253
rect 336 69217 342 69229
rect 224 69161 226 69177
rect 332 69149 342 69217
rect 400 69221 404 69229
rect 400 69187 408 69221
rect 434 69187 438 69221
rect 454 69205 504 69207
rect 504 69189 506 69205
rect 514 69199 530 69205
rect 532 69199 548 69205
rect 525 69189 548 69198
rect 400 69179 404 69187
rect 498 69179 506 69189
rect 504 69155 506 69179
rect 514 69169 515 69189
rect 525 69164 528 69189
rect 547 69169 548 69189
rect 557 69179 564 69189
rect 514 69155 548 69159
rect 151 69108 156 69142
rect 174 69139 246 69147
rect 256 69139 328 69147
rect 336 69141 342 69149
rect 400 69144 404 69149
rect 180 69111 185 69139
rect 174 69103 246 69111
rect 256 69103 328 69111
rect 332 69109 336 69139
rect 400 69110 438 69144
rect 224 69073 226 69089
rect 196 69065 226 69073
rect 196 69061 232 69065
rect 196 69031 204 69061
rect 216 69031 232 69061
rect 224 68984 226 69031
rect 300 69004 308 69073
rect 332 69071 342 69109
rect 400 69101 404 69110
rect 454 69095 504 69097
rect 494 69091 548 69095
rect 494 69086 514 69091
rect 504 69071 506 69086
rect 336 69059 342 69071
rect 289 68994 308 69004
rect 300 68988 308 68994
rect 332 69025 342 69059
rect 400 69063 404 69071
rect 400 69029 408 69063
rect 434 69029 438 69063
rect 498 69061 506 69071
rect 514 69061 515 69081
rect 504 69045 506 69061
rect 525 69052 528 69086
rect 547 69061 548 69081
rect 557 69061 564 69071
rect 514 69045 530 69051
rect 532 69045 548 69051
rect 332 68997 373 69025
rect 332 68991 351 68997
rect 107 68937 119 68971
rect 129 68937 149 68971
rect 196 68950 204 68984
rect 216 68950 232 68984
rect 244 68978 257 68984
rect 278 68978 291 68988
rect 244 68954 291 68978
rect 300 68978 321 68988
rect 336 68981 351 68991
rect 300 68954 329 68978
rect 332 68963 351 68981
rect 361 68991 375 68997
rect 400 68991 411 69029
rect 562 68992 612 68994
rect 361 68963 381 68991
rect 400 68963 409 68991
rect 466 68983 497 68991
rect 565 68983 596 68991
rect 442 68976 500 68983
rect 466 68975 500 68976
rect 565 68975 599 68983
rect 244 68950 257 68954
rect 42 68871 46 68905
rect 72 68871 76 68905
rect 42 68824 76 68828
rect 42 68809 46 68824
rect 72 68809 76 68824
rect 38 68791 80 68809
rect 16 68785 102 68791
rect 144 68785 148 68937
rect 174 68913 181 68941
rect 224 68903 226 68950
rect 300 68941 308 68954
rect 278 68930 305 68941
rect 332 68913 342 68963
rect 400 68943 404 68963
rect 497 68959 500 68975
rect 596 68959 599 68975
rect 466 68958 500 68959
rect 442 68951 500 68958
rect 565 68951 599 68959
rect 612 68942 614 68992
rect 256 68903 328 68911
rect 336 68905 342 68913
rect 400 68905 404 68913
rect 196 68873 204 68903
rect 216 68873 232 68903
rect 196 68869 232 68873
rect 196 68861 226 68869
rect 224 68845 226 68861
rect 332 68833 336 68901
rect 400 68871 408 68905
rect 434 68871 438 68905
rect 454 68889 504 68891
rect 504 68873 506 68889
rect 514 68883 530 68889
rect 532 68883 548 68889
rect 525 68873 548 68882
rect 400 68863 404 68871
rect 498 68863 506 68873
rect 504 68839 506 68863
rect 514 68853 515 68873
rect 525 68848 528 68873
rect 547 68853 548 68873
rect 557 68863 564 68873
rect 514 68839 548 68843
rect 400 68833 442 68834
rect 174 68823 246 68831
rect 400 68826 404 68833
rect 295 68792 300 68826
rect 324 68792 329 68826
rect 367 68809 438 68826
rect 367 68792 442 68809
rect 400 68791 442 68792
rect 378 68785 464 68791
rect 38 68769 80 68785
rect 400 68769 442 68785
rect -25 68755 25 68757
rect 42 68755 76 68769
rect 404 68755 438 68769
rect 455 68755 505 68757
rect 557 68755 607 68757
rect 16 68747 102 68755
rect 378 68747 464 68755
rect 8 68713 17 68747
rect 18 68745 51 68747
rect 80 68745 100 68747
rect 18 68713 100 68745
rect 380 68745 404 68747
rect 429 68745 438 68747
rect 442 68745 462 68747
rect 16 68705 102 68713
rect 42 68689 76 68705
rect 16 68669 38 68675
rect 42 68666 76 68670
rect 80 68669 102 68675
rect 42 68636 46 68666
rect 72 68636 76 68666
rect 42 68555 46 68589
rect 72 68555 76 68589
rect -25 68518 25 68520
rect -8 68510 14 68517
rect -8 68509 17 68510
rect 25 68509 27 68518
rect -12 68502 38 68509
rect -12 68501 34 68502
rect -12 68497 8 68501
rect 0 68485 8 68497
rect 14 68485 34 68501
rect 0 68484 34 68485
rect 0 68477 38 68484
rect 14 68476 17 68477
rect 25 68468 27 68477
rect 42 68448 45 68538
rect 69 68523 80 68555
rect 107 68523 143 68551
rect 144 68523 148 68743
rect 332 68675 336 68743
rect 380 68713 462 68745
rect 463 68713 472 68747
rect 480 68713 497 68747
rect 378 68705 464 68713
rect 505 68705 507 68755
rect 514 68713 548 68747
rect 565 68713 582 68747
rect 607 68705 609 68755
rect 404 68689 438 68705
rect 400 68675 442 68676
rect 378 68669 404 68675
rect 442 68669 464 68675
rect 400 68668 404 68669
rect 174 68629 246 68637
rect 295 68634 300 68668
rect 324 68634 329 68668
rect 224 68599 226 68615
rect 196 68591 226 68599
rect 332 68597 336 68665
rect 367 68634 438 68668
rect 400 68627 404 68634
rect 454 68621 504 68623
rect 494 68617 548 68621
rect 494 68612 514 68617
rect 504 68597 506 68612
rect 196 68587 232 68591
rect 196 68557 204 68587
rect 216 68557 232 68587
rect 400 68589 404 68597
rect 107 68517 119 68523
rect 109 68489 119 68517
rect 129 68489 149 68523
rect 174 68519 181 68549
rect 224 68510 226 68557
rect 256 68549 328 68557
rect 332 68555 336 68585
rect 400 68555 408 68589
rect 434 68555 438 68589
rect 498 68587 506 68597
rect 514 68587 515 68607
rect 504 68571 506 68587
rect 525 68578 528 68612
rect 547 68587 548 68607
rect 557 68587 564 68597
rect 514 68571 530 68577
rect 532 68571 548 68577
rect 278 68519 305 68530
rect 42 68397 46 68431
rect 72 68397 76 68431
rect 38 68359 80 68360
rect 42 68318 76 68352
rect 79 68318 113 68352
rect 42 68239 46 68273
rect 72 68239 76 68273
rect -25 68202 25 68204
rect -8 68194 14 68201
rect -8 68193 17 68194
rect 25 68193 27 68202
rect -12 68186 38 68193
rect -12 68185 34 68186
rect -12 68181 8 68185
rect 0 68169 8 68181
rect 14 68169 34 68185
rect 0 68168 34 68169
rect 0 68161 38 68168
rect 14 68160 17 68161
rect 25 68152 27 68161
rect 42 68132 45 68222
rect 71 68191 80 68219
rect 69 68153 80 68191
rect 144 68181 148 68489
rect 196 68476 204 68510
rect 216 68476 232 68510
rect 244 68506 257 68510
rect 300 68506 308 68519
rect 332 68517 342 68555
rect 400 68547 404 68555
rect 336 68507 342 68517
rect 244 68482 291 68506
rect 244 68476 257 68482
rect 224 68429 226 68476
rect 278 68472 291 68482
rect 300 68482 329 68506
rect 332 68497 342 68507
rect 400 68507 409 68535
rect 562 68518 612 68520
rect 466 68509 497 68517
rect 565 68509 596 68517
rect 300 68472 321 68482
rect 300 68466 308 68472
rect 289 68456 308 68466
rect 196 68399 204 68429
rect 216 68399 232 68429
rect 196 68395 232 68399
rect 196 68387 226 68395
rect 300 68387 308 68456
rect 332 68463 351 68497
rect 361 68469 381 68497
rect 361 68463 375 68469
rect 400 68463 411 68507
rect 442 68502 500 68509
rect 466 68501 500 68502
rect 565 68501 599 68509
rect 497 68485 500 68501
rect 596 68485 599 68501
rect 466 68484 500 68485
rect 442 68477 500 68484
rect 565 68477 599 68485
rect 612 68468 614 68518
rect 332 68439 342 68463
rect 336 68427 342 68439
rect 224 68371 226 68387
rect 332 68359 342 68427
rect 400 68431 404 68439
rect 400 68397 408 68431
rect 434 68397 438 68431
rect 454 68415 504 68417
rect 504 68399 506 68415
rect 514 68409 530 68415
rect 532 68409 548 68415
rect 525 68399 548 68408
rect 400 68389 404 68397
rect 498 68389 506 68399
rect 504 68365 506 68389
rect 514 68379 515 68399
rect 525 68374 528 68399
rect 547 68379 548 68399
rect 557 68389 564 68399
rect 514 68365 548 68369
rect 151 68318 156 68352
rect 174 68349 246 68357
rect 256 68349 328 68357
rect 336 68351 342 68359
rect 400 68354 404 68359
rect 180 68321 185 68349
rect 174 68313 246 68321
rect 256 68313 328 68321
rect 332 68319 336 68349
rect 400 68320 438 68354
rect 224 68283 226 68299
rect 196 68275 226 68283
rect 196 68271 232 68275
rect 196 68241 204 68271
rect 216 68241 232 68271
rect 224 68194 226 68241
rect 300 68214 308 68283
rect 332 68281 342 68319
rect 400 68311 404 68320
rect 454 68305 504 68307
rect 494 68301 548 68305
rect 494 68296 514 68301
rect 504 68281 506 68296
rect 336 68269 342 68281
rect 289 68204 308 68214
rect 300 68198 308 68204
rect 332 68235 342 68269
rect 400 68273 404 68281
rect 400 68239 408 68273
rect 434 68239 438 68273
rect 498 68271 506 68281
rect 514 68271 515 68291
rect 504 68255 506 68271
rect 525 68262 528 68296
rect 547 68271 548 68291
rect 557 68271 564 68281
rect 514 68255 530 68261
rect 532 68255 548 68261
rect 332 68207 373 68235
rect 332 68201 351 68207
rect 107 68147 119 68181
rect 129 68147 149 68181
rect 196 68160 204 68194
rect 216 68160 232 68194
rect 244 68188 257 68194
rect 278 68188 291 68198
rect 244 68164 291 68188
rect 300 68188 321 68198
rect 336 68191 351 68201
rect 300 68164 329 68188
rect 332 68173 351 68191
rect 361 68201 375 68207
rect 400 68201 411 68239
rect 562 68202 612 68204
rect 361 68173 381 68201
rect 400 68173 409 68201
rect 466 68193 497 68201
rect 565 68193 596 68201
rect 442 68186 500 68193
rect 466 68185 500 68186
rect 565 68185 599 68193
rect 244 68160 257 68164
rect 42 68081 46 68115
rect 72 68081 76 68115
rect 42 68034 76 68038
rect 42 68019 46 68034
rect 72 68019 76 68034
rect 38 68001 80 68019
rect 16 67995 102 68001
rect 144 67995 148 68147
rect 174 68123 181 68151
rect 224 68113 226 68160
rect 300 68151 308 68164
rect 278 68140 305 68151
rect 332 68123 342 68173
rect 400 68153 404 68173
rect 497 68169 500 68185
rect 596 68169 599 68185
rect 466 68168 500 68169
rect 442 68161 500 68168
rect 565 68161 599 68169
rect 612 68152 614 68202
rect 256 68113 328 68121
rect 336 68115 342 68123
rect 400 68115 404 68123
rect 196 68083 204 68113
rect 216 68083 232 68113
rect 196 68079 232 68083
rect 196 68071 226 68079
rect 224 68055 226 68071
rect 332 68043 336 68111
rect 400 68081 408 68115
rect 434 68081 438 68115
rect 454 68099 504 68101
rect 504 68083 506 68099
rect 514 68093 530 68099
rect 532 68093 548 68099
rect 525 68083 548 68092
rect 400 68073 404 68081
rect 498 68073 506 68083
rect 504 68049 506 68073
rect 514 68063 515 68083
rect 525 68058 528 68083
rect 547 68063 548 68083
rect 557 68073 564 68083
rect 514 68049 548 68053
rect 400 68043 442 68044
rect 174 68033 246 68041
rect 400 68036 404 68043
rect 295 68002 300 68036
rect 324 68002 329 68036
rect 367 68019 438 68036
rect 367 68002 442 68019
rect 400 68001 442 68002
rect 378 67995 464 68001
rect 38 67979 80 67995
rect 400 67979 442 67995
rect -25 67965 25 67967
rect 42 67965 76 67979
rect 404 67965 438 67979
rect 455 67965 505 67967
rect 557 67965 607 67967
rect 16 67957 102 67965
rect 378 67957 464 67965
rect 8 67923 17 67957
rect 18 67955 51 67957
rect 80 67955 100 67957
rect 18 67923 100 67955
rect 380 67955 404 67957
rect 429 67955 438 67957
rect 442 67955 462 67957
rect 16 67915 102 67923
rect 42 67899 76 67915
rect 16 67879 38 67885
rect 42 67876 76 67880
rect 80 67879 102 67885
rect 42 67846 46 67876
rect 72 67846 76 67876
rect 42 67765 46 67799
rect 72 67765 76 67799
rect -25 67728 25 67730
rect -8 67720 14 67727
rect -8 67719 17 67720
rect 25 67719 27 67728
rect -12 67712 38 67719
rect -12 67711 34 67712
rect -12 67707 8 67711
rect 0 67695 8 67707
rect 14 67695 34 67711
rect 0 67694 34 67695
rect 0 67687 38 67694
rect 14 67686 17 67687
rect 25 67678 27 67687
rect 42 67658 45 67748
rect 69 67733 80 67765
rect 107 67733 143 67761
rect 144 67733 148 67953
rect 332 67885 336 67953
rect 380 67923 462 67955
rect 463 67923 472 67957
rect 480 67923 497 67957
rect 378 67915 464 67923
rect 505 67915 507 67965
rect 514 67923 548 67957
rect 565 67923 582 67957
rect 607 67915 609 67965
rect 404 67899 438 67915
rect 400 67885 442 67886
rect 378 67879 404 67885
rect 442 67879 464 67885
rect 400 67878 404 67879
rect 174 67839 246 67847
rect 295 67844 300 67878
rect 324 67844 329 67878
rect 224 67809 226 67825
rect 196 67801 226 67809
rect 332 67807 336 67875
rect 367 67844 438 67878
rect 400 67837 404 67844
rect 454 67831 504 67833
rect 494 67827 548 67831
rect 494 67822 514 67827
rect 504 67807 506 67822
rect 196 67797 232 67801
rect 196 67767 204 67797
rect 216 67767 232 67797
rect 400 67799 404 67807
rect 107 67727 119 67733
rect 109 67699 119 67727
rect 129 67699 149 67733
rect 174 67729 181 67759
rect 224 67720 226 67767
rect 256 67759 328 67767
rect 332 67765 336 67795
rect 400 67765 408 67799
rect 434 67765 438 67799
rect 498 67797 506 67807
rect 514 67797 515 67817
rect 504 67781 506 67797
rect 525 67788 528 67822
rect 547 67797 548 67817
rect 557 67797 564 67807
rect 514 67781 530 67787
rect 532 67781 548 67787
rect 278 67729 305 67740
rect 42 67607 46 67641
rect 72 67607 76 67641
rect 38 67569 80 67570
rect 42 67528 76 67562
rect 79 67528 113 67562
rect 42 67449 46 67483
rect 72 67449 76 67483
rect -25 67412 25 67414
rect -8 67404 14 67411
rect -8 67403 17 67404
rect 25 67403 27 67412
rect -12 67396 38 67403
rect -12 67395 34 67396
rect -12 67391 8 67395
rect 0 67379 8 67391
rect 14 67379 34 67395
rect 0 67378 34 67379
rect 0 67371 38 67378
rect 14 67370 17 67371
rect 25 67362 27 67371
rect 42 67342 45 67432
rect 71 67401 80 67429
rect 69 67363 80 67401
rect 144 67391 148 67699
rect 196 67686 204 67720
rect 216 67686 232 67720
rect 244 67716 257 67720
rect 300 67716 308 67729
rect 332 67727 342 67765
rect 400 67757 404 67765
rect 336 67717 342 67727
rect 244 67692 291 67716
rect 244 67686 257 67692
rect 224 67639 226 67686
rect 278 67682 291 67692
rect 300 67692 329 67716
rect 332 67707 342 67717
rect 400 67717 409 67745
rect 562 67728 612 67730
rect 466 67719 497 67727
rect 565 67719 596 67727
rect 300 67682 321 67692
rect 300 67676 308 67682
rect 289 67666 308 67676
rect 196 67609 204 67639
rect 216 67609 232 67639
rect 196 67605 232 67609
rect 196 67597 226 67605
rect 300 67597 308 67666
rect 332 67673 351 67707
rect 361 67679 381 67707
rect 361 67673 375 67679
rect 400 67673 411 67717
rect 442 67712 500 67719
rect 466 67711 500 67712
rect 565 67711 599 67719
rect 497 67695 500 67711
rect 596 67695 599 67711
rect 466 67694 500 67695
rect 442 67687 500 67694
rect 565 67687 599 67695
rect 612 67678 614 67728
rect 332 67649 342 67673
rect 336 67637 342 67649
rect 224 67581 226 67597
rect 332 67569 342 67637
rect 400 67641 404 67649
rect 400 67607 408 67641
rect 434 67607 438 67641
rect 454 67625 504 67627
rect 504 67609 506 67625
rect 514 67619 530 67625
rect 532 67619 548 67625
rect 525 67609 548 67618
rect 400 67599 404 67607
rect 498 67599 506 67609
rect 504 67575 506 67599
rect 514 67589 515 67609
rect 525 67584 528 67609
rect 547 67589 548 67609
rect 557 67599 564 67609
rect 514 67575 548 67579
rect 151 67528 156 67562
rect 174 67559 246 67567
rect 256 67559 328 67567
rect 336 67561 342 67569
rect 400 67564 404 67569
rect 180 67531 185 67559
rect 174 67523 246 67531
rect 256 67523 328 67531
rect 332 67529 336 67559
rect 400 67530 438 67564
rect 224 67493 226 67509
rect 196 67485 226 67493
rect 196 67481 232 67485
rect 196 67451 204 67481
rect 216 67451 232 67481
rect 224 67404 226 67451
rect 300 67424 308 67493
rect 332 67491 342 67529
rect 400 67521 404 67530
rect 454 67515 504 67517
rect 494 67511 548 67515
rect 494 67506 514 67511
rect 504 67491 506 67506
rect 336 67479 342 67491
rect 289 67414 308 67424
rect 300 67408 308 67414
rect 332 67445 342 67479
rect 400 67483 404 67491
rect 400 67449 408 67483
rect 434 67449 438 67483
rect 498 67481 506 67491
rect 514 67481 515 67501
rect 504 67465 506 67481
rect 525 67472 528 67506
rect 547 67481 548 67501
rect 557 67481 564 67491
rect 514 67465 530 67471
rect 532 67465 548 67471
rect 332 67417 373 67445
rect 332 67411 351 67417
rect 107 67357 119 67391
rect 129 67357 149 67391
rect 196 67370 204 67404
rect 216 67370 232 67404
rect 244 67398 257 67404
rect 278 67398 291 67408
rect 244 67374 291 67398
rect 300 67398 321 67408
rect 336 67401 351 67411
rect 300 67374 329 67398
rect 332 67383 351 67401
rect 361 67411 375 67417
rect 400 67411 411 67449
rect 562 67412 612 67414
rect 361 67383 381 67411
rect 400 67383 409 67411
rect 466 67403 497 67411
rect 565 67403 596 67411
rect 442 67396 500 67403
rect 466 67395 500 67396
rect 565 67395 599 67403
rect 244 67370 257 67374
rect 42 67291 46 67325
rect 72 67291 76 67325
rect 42 67244 76 67248
rect 42 67229 46 67244
rect 72 67229 76 67244
rect 38 67211 80 67229
rect 16 67205 102 67211
rect 144 67205 148 67357
rect 174 67333 181 67361
rect 224 67323 226 67370
rect 300 67361 308 67374
rect 278 67350 305 67361
rect 332 67333 342 67383
rect 400 67363 404 67383
rect 497 67379 500 67395
rect 596 67379 599 67395
rect 466 67378 500 67379
rect 442 67371 500 67378
rect 565 67371 599 67379
rect 612 67362 614 67412
rect 256 67323 328 67331
rect 336 67325 342 67333
rect 400 67325 404 67333
rect 196 67293 204 67323
rect 216 67293 232 67323
rect 196 67289 232 67293
rect 196 67281 226 67289
rect 224 67265 226 67281
rect 332 67253 336 67321
rect 400 67291 408 67325
rect 434 67291 438 67325
rect 454 67309 504 67311
rect 504 67293 506 67309
rect 514 67303 530 67309
rect 532 67303 548 67309
rect 525 67293 548 67302
rect 400 67283 404 67291
rect 498 67283 506 67293
rect 504 67259 506 67283
rect 514 67273 515 67293
rect 525 67268 528 67293
rect 547 67273 548 67293
rect 557 67283 564 67293
rect 514 67259 548 67263
rect 400 67253 442 67254
rect 174 67243 246 67251
rect 400 67246 404 67253
rect 295 67212 300 67246
rect 324 67212 329 67246
rect 367 67229 438 67246
rect 367 67212 442 67229
rect 400 67211 442 67212
rect 378 67205 464 67211
rect 38 67189 80 67205
rect 400 67189 442 67205
rect -25 67175 25 67177
rect 42 67175 76 67189
rect 404 67175 438 67189
rect 455 67175 505 67177
rect 557 67175 607 67177
rect 16 67167 102 67175
rect 378 67167 464 67175
rect 8 67133 17 67167
rect 18 67165 51 67167
rect 80 67165 100 67167
rect 18 67133 100 67165
rect 380 67165 404 67167
rect 429 67165 438 67167
rect 442 67165 462 67167
rect 16 67125 102 67133
rect 42 67109 76 67125
rect 16 67089 38 67095
rect 42 67086 76 67090
rect 80 67089 102 67095
rect 42 67056 46 67086
rect 72 67056 76 67086
rect 42 66975 46 67009
rect 72 66975 76 67009
rect -25 66938 25 66940
rect -8 66930 14 66937
rect -8 66929 17 66930
rect 25 66929 27 66938
rect -12 66922 38 66929
rect -12 66921 34 66922
rect -12 66917 8 66921
rect 0 66905 8 66917
rect 14 66905 34 66921
rect 0 66904 34 66905
rect 0 66897 38 66904
rect 14 66896 17 66897
rect 25 66888 27 66897
rect 42 66868 45 66958
rect 69 66943 80 66975
rect 107 66943 143 66971
rect 144 66943 148 67163
rect 332 67095 336 67163
rect 380 67133 462 67165
rect 463 67133 472 67167
rect 480 67133 497 67167
rect 378 67125 464 67133
rect 505 67125 507 67175
rect 514 67133 548 67167
rect 565 67133 582 67167
rect 607 67125 609 67175
rect 404 67109 438 67125
rect 400 67095 442 67096
rect 378 67089 404 67095
rect 442 67089 464 67095
rect 400 67088 404 67089
rect 174 67049 246 67057
rect 295 67054 300 67088
rect 324 67054 329 67088
rect 224 67019 226 67035
rect 196 67011 226 67019
rect 332 67017 336 67085
rect 367 67054 438 67088
rect 400 67047 404 67054
rect 454 67041 504 67043
rect 494 67037 548 67041
rect 494 67032 514 67037
rect 504 67017 506 67032
rect 196 67007 232 67011
rect 196 66977 204 67007
rect 216 66977 232 67007
rect 400 67009 404 67017
rect 107 66937 119 66943
rect 109 66909 119 66937
rect 129 66909 149 66943
rect 174 66939 181 66969
rect 224 66930 226 66977
rect 256 66969 328 66977
rect 332 66975 336 67005
rect 400 66975 408 67009
rect 434 66975 438 67009
rect 498 67007 506 67017
rect 514 67007 515 67027
rect 504 66991 506 67007
rect 525 66998 528 67032
rect 547 67007 548 67027
rect 557 67007 564 67017
rect 514 66991 530 66997
rect 532 66991 548 66997
rect 278 66939 305 66950
rect 42 66817 46 66851
rect 72 66817 76 66851
rect 38 66779 80 66780
rect 42 66738 76 66772
rect 79 66738 113 66772
rect 42 66659 46 66693
rect 72 66659 76 66693
rect -25 66622 25 66624
rect -8 66614 14 66621
rect -8 66613 17 66614
rect 25 66613 27 66622
rect -12 66606 38 66613
rect -12 66605 34 66606
rect -12 66601 8 66605
rect 0 66589 8 66601
rect 14 66589 34 66605
rect 0 66588 34 66589
rect 0 66581 38 66588
rect 14 66580 17 66581
rect 25 66572 27 66581
rect 42 66552 45 66642
rect 71 66611 80 66639
rect 69 66573 80 66611
rect 144 66601 148 66909
rect 196 66896 204 66930
rect 216 66896 232 66930
rect 244 66926 257 66930
rect 300 66926 308 66939
rect 332 66937 342 66975
rect 400 66967 404 66975
rect 336 66927 342 66937
rect 244 66902 291 66926
rect 244 66896 257 66902
rect 224 66849 226 66896
rect 278 66892 291 66902
rect 300 66902 329 66926
rect 332 66917 342 66927
rect 400 66927 409 66955
rect 562 66938 612 66940
rect 466 66929 497 66937
rect 565 66929 596 66937
rect 300 66892 321 66902
rect 300 66886 308 66892
rect 289 66876 308 66886
rect 196 66819 204 66849
rect 216 66819 232 66849
rect 196 66815 232 66819
rect 196 66807 226 66815
rect 300 66807 308 66876
rect 332 66883 351 66917
rect 361 66889 381 66917
rect 361 66883 375 66889
rect 400 66883 411 66927
rect 442 66922 500 66929
rect 466 66921 500 66922
rect 565 66921 599 66929
rect 497 66905 500 66921
rect 596 66905 599 66921
rect 466 66904 500 66905
rect 442 66897 500 66904
rect 565 66897 599 66905
rect 612 66888 614 66938
rect 332 66859 342 66883
rect 336 66847 342 66859
rect 224 66791 226 66807
rect 332 66779 342 66847
rect 400 66851 404 66859
rect 400 66817 408 66851
rect 434 66817 438 66851
rect 454 66835 504 66837
rect 504 66819 506 66835
rect 514 66829 530 66835
rect 532 66829 548 66835
rect 525 66819 548 66828
rect 400 66809 404 66817
rect 498 66809 506 66819
rect 504 66785 506 66809
rect 514 66799 515 66819
rect 525 66794 528 66819
rect 547 66799 548 66819
rect 557 66809 564 66819
rect 514 66785 548 66789
rect 151 66738 156 66772
rect 174 66769 246 66777
rect 256 66769 328 66777
rect 336 66771 342 66779
rect 400 66774 404 66779
rect 180 66741 185 66769
rect 174 66733 246 66741
rect 256 66733 328 66741
rect 332 66739 336 66769
rect 400 66740 438 66774
rect 224 66703 226 66719
rect 196 66695 226 66703
rect 196 66691 232 66695
rect 196 66661 204 66691
rect 216 66661 232 66691
rect 224 66614 226 66661
rect 300 66634 308 66703
rect 332 66701 342 66739
rect 400 66731 404 66740
rect 454 66725 504 66727
rect 494 66721 548 66725
rect 494 66716 514 66721
rect 504 66701 506 66716
rect 336 66689 342 66701
rect 289 66624 308 66634
rect 300 66618 308 66624
rect 332 66655 342 66689
rect 400 66693 404 66701
rect 400 66659 408 66693
rect 434 66659 438 66693
rect 498 66691 506 66701
rect 514 66691 515 66711
rect 504 66675 506 66691
rect 525 66682 528 66716
rect 547 66691 548 66711
rect 557 66691 564 66701
rect 514 66675 530 66681
rect 532 66675 548 66681
rect 332 66627 373 66655
rect 332 66621 351 66627
rect 107 66567 119 66601
rect 129 66567 149 66601
rect 196 66580 204 66614
rect 216 66580 232 66614
rect 244 66608 257 66614
rect 278 66608 291 66618
rect 244 66584 291 66608
rect 300 66608 321 66618
rect 336 66611 351 66621
rect 300 66584 329 66608
rect 332 66593 351 66611
rect 361 66621 375 66627
rect 400 66621 411 66659
rect 562 66622 612 66624
rect 361 66593 381 66621
rect 400 66593 409 66621
rect 466 66613 497 66621
rect 565 66613 596 66621
rect 442 66606 500 66613
rect 466 66605 500 66606
rect 565 66605 599 66613
rect 244 66580 257 66584
rect 42 66501 46 66535
rect 72 66501 76 66535
rect 42 66454 76 66458
rect 42 66439 46 66454
rect 72 66439 76 66454
rect 38 66421 80 66439
rect 16 66415 102 66421
rect 144 66415 148 66567
rect 174 66543 181 66571
rect 224 66533 226 66580
rect 300 66571 308 66584
rect 278 66560 305 66571
rect 332 66543 342 66593
rect 400 66573 404 66593
rect 497 66589 500 66605
rect 596 66589 599 66605
rect 466 66588 500 66589
rect 442 66581 500 66588
rect 565 66581 599 66589
rect 612 66572 614 66622
rect 256 66533 328 66541
rect 336 66535 342 66543
rect 400 66535 404 66543
rect 196 66503 204 66533
rect 216 66503 232 66533
rect 196 66499 232 66503
rect 196 66491 226 66499
rect 224 66475 226 66491
rect 332 66463 336 66531
rect 400 66501 408 66535
rect 434 66501 438 66535
rect 454 66519 504 66521
rect 504 66503 506 66519
rect 514 66513 530 66519
rect 532 66513 548 66519
rect 525 66503 548 66512
rect 400 66493 404 66501
rect 498 66493 506 66503
rect 504 66469 506 66493
rect 514 66483 515 66503
rect 525 66478 528 66503
rect 547 66483 548 66503
rect 557 66493 564 66503
rect 514 66469 548 66473
rect 400 66463 442 66464
rect 174 66453 246 66461
rect 400 66456 404 66463
rect 295 66422 300 66456
rect 324 66422 329 66456
rect 367 66439 438 66456
rect 367 66422 442 66439
rect 400 66421 442 66422
rect 378 66415 464 66421
rect 38 66399 80 66415
rect 400 66399 442 66415
rect -25 66385 25 66387
rect 42 66385 76 66399
rect 404 66385 438 66399
rect 455 66385 505 66387
rect 557 66385 607 66387
rect 16 66377 102 66385
rect 378 66377 464 66385
rect 8 66343 17 66377
rect 18 66375 51 66377
rect 80 66375 100 66377
rect 18 66343 100 66375
rect 380 66375 404 66377
rect 429 66375 438 66377
rect 442 66375 462 66377
rect 16 66335 102 66343
rect 42 66319 76 66335
rect 16 66299 38 66305
rect 42 66296 76 66300
rect 80 66299 102 66305
rect 42 66266 46 66296
rect 72 66266 76 66296
rect 42 66185 46 66219
rect 72 66185 76 66219
rect -25 66148 25 66150
rect -8 66140 14 66147
rect -8 66139 17 66140
rect 25 66139 27 66148
rect -12 66132 38 66139
rect -12 66131 34 66132
rect -12 66127 8 66131
rect 0 66115 8 66127
rect 14 66115 34 66131
rect 0 66114 34 66115
rect 0 66107 38 66114
rect 14 66106 17 66107
rect 25 66098 27 66107
rect 42 66078 45 66168
rect 69 66153 80 66185
rect 107 66153 143 66181
rect 144 66153 148 66373
rect 332 66305 336 66373
rect 380 66343 462 66375
rect 463 66343 472 66377
rect 480 66343 497 66377
rect 378 66335 464 66343
rect 505 66335 507 66385
rect 514 66343 548 66377
rect 565 66343 582 66377
rect 607 66335 609 66385
rect 404 66319 438 66335
rect 400 66305 442 66306
rect 378 66299 404 66305
rect 442 66299 464 66305
rect 400 66298 404 66299
rect 174 66259 246 66267
rect 295 66264 300 66298
rect 324 66264 329 66298
rect 224 66229 226 66245
rect 196 66221 226 66229
rect 332 66227 336 66295
rect 367 66264 438 66298
rect 400 66257 404 66264
rect 454 66251 504 66253
rect 494 66247 548 66251
rect 494 66242 514 66247
rect 504 66227 506 66242
rect 196 66217 232 66221
rect 196 66187 204 66217
rect 216 66187 232 66217
rect 400 66219 404 66227
rect 107 66147 119 66153
rect 109 66119 119 66147
rect 129 66119 149 66153
rect 174 66149 181 66179
rect 224 66140 226 66187
rect 256 66179 328 66187
rect 332 66185 336 66215
rect 400 66185 408 66219
rect 434 66185 438 66219
rect 498 66217 506 66227
rect 514 66217 515 66237
rect 504 66201 506 66217
rect 525 66208 528 66242
rect 547 66217 548 66237
rect 557 66217 564 66227
rect 514 66201 530 66207
rect 532 66201 548 66207
rect 278 66149 305 66160
rect 42 66027 46 66061
rect 72 66027 76 66061
rect 38 65989 80 65990
rect 42 65948 76 65982
rect 79 65948 113 65982
rect 42 65869 46 65903
rect 72 65869 76 65903
rect -25 65832 25 65834
rect -8 65824 14 65831
rect -8 65823 17 65824
rect 25 65823 27 65832
rect -12 65816 38 65823
rect -12 65815 34 65816
rect -12 65811 8 65815
rect 0 65799 8 65811
rect 14 65799 34 65815
rect 0 65798 34 65799
rect 0 65791 38 65798
rect 14 65790 17 65791
rect 25 65782 27 65791
rect 42 65762 45 65852
rect 71 65821 80 65849
rect 69 65783 80 65821
rect 144 65811 148 66119
rect 196 66106 204 66140
rect 216 66106 232 66140
rect 244 66136 257 66140
rect 300 66136 308 66149
rect 332 66147 342 66185
rect 400 66177 404 66185
rect 336 66137 342 66147
rect 244 66112 291 66136
rect 244 66106 257 66112
rect 224 66059 226 66106
rect 278 66102 291 66112
rect 300 66112 329 66136
rect 332 66127 342 66137
rect 400 66137 409 66165
rect 562 66148 612 66150
rect 466 66139 497 66147
rect 565 66139 596 66147
rect 300 66102 321 66112
rect 300 66096 308 66102
rect 289 66086 308 66096
rect 196 66029 204 66059
rect 216 66029 232 66059
rect 196 66025 232 66029
rect 196 66017 226 66025
rect 300 66017 308 66086
rect 332 66093 351 66127
rect 361 66099 381 66127
rect 361 66093 375 66099
rect 400 66093 411 66137
rect 442 66132 500 66139
rect 466 66131 500 66132
rect 565 66131 599 66139
rect 497 66115 500 66131
rect 596 66115 599 66131
rect 466 66114 500 66115
rect 442 66107 500 66114
rect 565 66107 599 66115
rect 612 66098 614 66148
rect 332 66069 342 66093
rect 336 66057 342 66069
rect 224 66001 226 66017
rect 332 65989 342 66057
rect 400 66061 404 66069
rect 400 66027 408 66061
rect 434 66027 438 66061
rect 454 66045 504 66047
rect 504 66029 506 66045
rect 514 66039 530 66045
rect 532 66039 548 66045
rect 525 66029 548 66038
rect 400 66019 404 66027
rect 498 66019 506 66029
rect 504 65995 506 66019
rect 514 66009 515 66029
rect 525 66004 528 66029
rect 547 66009 548 66029
rect 557 66019 564 66029
rect 514 65995 548 65999
rect 151 65948 156 65982
rect 174 65979 246 65987
rect 256 65979 328 65987
rect 336 65981 342 65989
rect 400 65984 404 65989
rect 180 65951 185 65979
rect 174 65943 246 65951
rect 256 65943 328 65951
rect 332 65949 336 65979
rect 400 65950 438 65984
rect 224 65913 226 65929
rect 196 65905 226 65913
rect 196 65901 232 65905
rect 196 65871 204 65901
rect 216 65871 232 65901
rect 224 65824 226 65871
rect 300 65844 308 65913
rect 332 65911 342 65949
rect 400 65941 404 65950
rect 454 65935 504 65937
rect 494 65931 548 65935
rect 494 65926 514 65931
rect 504 65911 506 65926
rect 336 65899 342 65911
rect 289 65834 308 65844
rect 300 65828 308 65834
rect 332 65865 342 65899
rect 400 65903 404 65911
rect 400 65869 408 65903
rect 434 65869 438 65903
rect 498 65901 506 65911
rect 514 65901 515 65921
rect 504 65885 506 65901
rect 525 65892 528 65926
rect 547 65901 548 65921
rect 557 65901 564 65911
rect 514 65885 530 65891
rect 532 65885 548 65891
rect 332 65837 373 65865
rect 332 65831 351 65837
rect 107 65777 119 65811
rect 129 65777 149 65811
rect 196 65790 204 65824
rect 216 65790 232 65824
rect 244 65818 257 65824
rect 278 65818 291 65828
rect 244 65794 291 65818
rect 300 65818 321 65828
rect 336 65821 351 65831
rect 300 65794 329 65818
rect 332 65803 351 65821
rect 361 65831 375 65837
rect 400 65831 411 65869
rect 562 65832 612 65834
rect 361 65803 381 65831
rect 400 65803 409 65831
rect 466 65823 497 65831
rect 565 65823 596 65831
rect 442 65816 500 65823
rect 466 65815 500 65816
rect 565 65815 599 65823
rect 244 65790 257 65794
rect 42 65711 46 65745
rect 72 65711 76 65745
rect 42 65664 76 65668
rect 42 65649 46 65664
rect 72 65649 76 65664
rect 38 65631 80 65649
rect 16 65625 102 65631
rect 144 65625 148 65777
rect 174 65753 181 65781
rect 224 65743 226 65790
rect 300 65781 308 65794
rect 278 65770 305 65781
rect 332 65753 342 65803
rect 400 65783 404 65803
rect 497 65799 500 65815
rect 596 65799 599 65815
rect 466 65798 500 65799
rect 442 65791 500 65798
rect 565 65791 599 65799
rect 612 65782 614 65832
rect 256 65743 328 65751
rect 336 65745 342 65753
rect 400 65745 404 65753
rect 196 65713 204 65743
rect 216 65713 232 65743
rect 196 65709 232 65713
rect 196 65701 226 65709
rect 224 65685 226 65701
rect 332 65673 336 65741
rect 400 65711 408 65745
rect 434 65711 438 65745
rect 454 65729 504 65731
rect 504 65713 506 65729
rect 514 65723 530 65729
rect 532 65723 548 65729
rect 525 65713 548 65722
rect 400 65703 404 65711
rect 498 65703 506 65713
rect 504 65679 506 65703
rect 514 65693 515 65713
rect 525 65688 528 65713
rect 547 65693 548 65713
rect 557 65703 564 65713
rect 514 65679 548 65683
rect 400 65673 442 65674
rect 174 65663 246 65671
rect 400 65666 404 65673
rect 295 65632 300 65666
rect 324 65632 329 65666
rect 367 65649 438 65666
rect 367 65632 442 65649
rect 400 65631 442 65632
rect 378 65625 464 65631
rect 38 65609 80 65625
rect 400 65609 442 65625
rect -25 65595 25 65597
rect 42 65595 76 65609
rect 404 65595 438 65609
rect 455 65595 505 65597
rect 557 65595 607 65597
rect 16 65587 102 65595
rect 378 65587 464 65595
rect 8 65553 17 65587
rect 18 65585 51 65587
rect 80 65585 100 65587
rect 18 65553 100 65585
rect 380 65585 404 65587
rect 429 65585 438 65587
rect 442 65585 462 65587
rect 16 65545 102 65553
rect 42 65529 76 65545
rect 16 65509 38 65515
rect 42 65506 76 65510
rect 80 65509 102 65515
rect 42 65476 46 65506
rect 72 65476 76 65506
rect 42 65395 46 65429
rect 72 65395 76 65429
rect -25 65358 25 65360
rect -8 65350 14 65357
rect -8 65349 17 65350
rect 25 65349 27 65358
rect -12 65342 38 65349
rect -12 65341 34 65342
rect -12 65337 8 65341
rect 0 65325 8 65337
rect 14 65325 34 65341
rect 0 65324 34 65325
rect 0 65317 38 65324
rect 14 65316 17 65317
rect 25 65308 27 65317
rect 42 65288 45 65378
rect 69 65363 80 65395
rect 107 65363 143 65391
rect 144 65363 148 65583
rect 332 65515 336 65583
rect 380 65553 462 65585
rect 463 65553 472 65587
rect 480 65553 497 65587
rect 378 65545 464 65553
rect 505 65545 507 65595
rect 514 65553 548 65587
rect 565 65553 582 65587
rect 607 65545 609 65595
rect 404 65529 438 65545
rect 400 65515 442 65516
rect 378 65509 404 65515
rect 442 65509 464 65515
rect 400 65508 404 65509
rect 174 65469 246 65477
rect 295 65474 300 65508
rect 324 65474 329 65508
rect 224 65439 226 65455
rect 196 65431 226 65439
rect 332 65437 336 65505
rect 367 65474 438 65508
rect 400 65467 404 65474
rect 454 65461 504 65463
rect 494 65457 548 65461
rect 494 65452 514 65457
rect 504 65437 506 65452
rect 196 65427 232 65431
rect 196 65397 204 65427
rect 216 65397 232 65427
rect 400 65429 404 65437
rect 107 65357 119 65363
rect 109 65329 119 65357
rect 129 65329 149 65363
rect 174 65359 181 65389
rect 224 65350 226 65397
rect 256 65389 328 65397
rect 332 65395 336 65425
rect 400 65395 408 65429
rect 434 65395 438 65429
rect 498 65427 506 65437
rect 514 65427 515 65447
rect 504 65411 506 65427
rect 525 65418 528 65452
rect 547 65427 548 65447
rect 557 65427 564 65437
rect 514 65411 530 65417
rect 532 65411 548 65417
rect 278 65359 305 65370
rect 42 65237 46 65271
rect 72 65237 76 65271
rect 38 65199 80 65200
rect 42 65158 76 65192
rect 79 65158 113 65192
rect 42 65079 46 65113
rect 72 65079 76 65113
rect -25 65042 25 65044
rect -8 65034 14 65041
rect -8 65033 17 65034
rect 25 65033 27 65042
rect -12 65026 38 65033
rect -12 65025 34 65026
rect -12 65021 8 65025
rect 0 65009 8 65021
rect 14 65009 34 65025
rect 0 65008 34 65009
rect 0 65001 38 65008
rect 14 65000 17 65001
rect 25 64992 27 65001
rect 42 64972 45 65062
rect 71 65031 80 65059
rect 69 64993 80 65031
rect 144 65021 148 65329
rect 196 65316 204 65350
rect 216 65316 232 65350
rect 244 65346 257 65350
rect 300 65346 308 65359
rect 332 65357 342 65395
rect 400 65387 404 65395
rect 336 65347 342 65357
rect 244 65322 291 65346
rect 244 65316 257 65322
rect 224 65269 226 65316
rect 278 65312 291 65322
rect 300 65322 329 65346
rect 332 65337 342 65347
rect 400 65347 409 65375
rect 562 65358 612 65360
rect 466 65349 497 65357
rect 565 65349 596 65357
rect 300 65312 321 65322
rect 300 65306 308 65312
rect 289 65296 308 65306
rect 196 65239 204 65269
rect 216 65239 232 65269
rect 196 65235 232 65239
rect 196 65227 226 65235
rect 300 65227 308 65296
rect 332 65303 351 65337
rect 361 65309 381 65337
rect 361 65303 375 65309
rect 400 65303 411 65347
rect 442 65342 500 65349
rect 466 65341 500 65342
rect 565 65341 599 65349
rect 497 65325 500 65341
rect 596 65325 599 65341
rect 466 65324 500 65325
rect 442 65317 500 65324
rect 565 65317 599 65325
rect 612 65308 614 65358
rect 332 65279 342 65303
rect 336 65267 342 65279
rect 224 65211 226 65227
rect 332 65199 342 65267
rect 400 65271 404 65279
rect 400 65237 408 65271
rect 434 65237 438 65271
rect 454 65255 504 65257
rect 504 65239 506 65255
rect 514 65249 530 65255
rect 532 65249 548 65255
rect 525 65239 548 65248
rect 400 65229 404 65237
rect 498 65229 506 65239
rect 504 65205 506 65229
rect 514 65219 515 65239
rect 525 65214 528 65239
rect 547 65219 548 65239
rect 557 65229 564 65239
rect 514 65205 548 65209
rect 151 65158 156 65192
rect 174 65189 246 65197
rect 256 65189 328 65197
rect 336 65191 342 65199
rect 400 65194 404 65199
rect 180 65161 185 65189
rect 174 65153 246 65161
rect 256 65153 328 65161
rect 332 65159 336 65189
rect 400 65160 438 65194
rect 224 65123 226 65139
rect 196 65115 226 65123
rect 196 65111 232 65115
rect 196 65081 204 65111
rect 216 65081 232 65111
rect 224 65034 226 65081
rect 300 65054 308 65123
rect 332 65121 342 65159
rect 400 65151 404 65160
rect 454 65145 504 65147
rect 494 65141 548 65145
rect 494 65136 514 65141
rect 504 65121 506 65136
rect 336 65109 342 65121
rect 289 65044 308 65054
rect 300 65038 308 65044
rect 332 65075 342 65109
rect 400 65113 404 65121
rect 400 65079 408 65113
rect 434 65079 438 65113
rect 498 65111 506 65121
rect 514 65111 515 65131
rect 504 65095 506 65111
rect 525 65102 528 65136
rect 547 65111 548 65131
rect 557 65111 564 65121
rect 514 65095 530 65101
rect 532 65095 548 65101
rect 332 65047 373 65075
rect 332 65041 351 65047
rect 107 64987 119 65021
rect 129 64987 149 65021
rect 196 65000 204 65034
rect 216 65000 232 65034
rect 244 65028 257 65034
rect 278 65028 291 65038
rect 244 65004 291 65028
rect 300 65028 321 65038
rect 336 65031 351 65041
rect 300 65004 329 65028
rect 332 65013 351 65031
rect 361 65041 375 65047
rect 400 65041 411 65079
rect 562 65042 612 65044
rect 361 65013 381 65041
rect 400 65013 409 65041
rect 466 65033 497 65041
rect 565 65033 596 65041
rect 442 65026 500 65033
rect 466 65025 500 65026
rect 565 65025 599 65033
rect 244 65000 257 65004
rect 42 64921 46 64955
rect 72 64921 76 64955
rect 42 64874 76 64878
rect 42 64859 46 64874
rect 72 64859 76 64874
rect 38 64841 80 64859
rect 16 64835 102 64841
rect 144 64835 148 64987
rect 174 64963 181 64991
rect 224 64953 226 65000
rect 300 64991 308 65004
rect 278 64980 305 64991
rect 332 64963 342 65013
rect 400 64993 404 65013
rect 497 65009 500 65025
rect 596 65009 599 65025
rect 466 65008 500 65009
rect 442 65001 500 65008
rect 565 65001 599 65009
rect 612 64992 614 65042
rect 256 64953 328 64961
rect 336 64955 342 64963
rect 400 64955 404 64963
rect 196 64923 204 64953
rect 216 64923 232 64953
rect 196 64919 232 64923
rect 196 64911 226 64919
rect 224 64895 226 64911
rect 332 64883 336 64951
rect 400 64921 408 64955
rect 434 64921 438 64955
rect 454 64939 504 64941
rect 504 64923 506 64939
rect 514 64933 530 64939
rect 532 64933 548 64939
rect 525 64923 548 64932
rect 400 64913 404 64921
rect 498 64913 506 64923
rect 504 64889 506 64913
rect 514 64903 515 64923
rect 525 64898 528 64923
rect 547 64903 548 64923
rect 557 64913 564 64923
rect 514 64889 548 64893
rect 400 64883 442 64884
rect 174 64873 246 64881
rect 400 64876 404 64883
rect 295 64842 300 64876
rect 324 64842 329 64876
rect 367 64859 438 64876
rect 367 64842 442 64859
rect 400 64841 442 64842
rect 378 64835 464 64841
rect 38 64819 80 64835
rect 400 64819 442 64835
rect -25 64805 25 64807
rect 42 64805 76 64819
rect 404 64805 438 64819
rect 455 64805 505 64807
rect 557 64805 607 64807
rect 16 64797 102 64805
rect 378 64797 464 64805
rect 8 64763 17 64797
rect 18 64795 51 64797
rect 80 64795 100 64797
rect 18 64763 100 64795
rect 380 64795 404 64797
rect 429 64795 438 64797
rect 442 64795 462 64797
rect 16 64755 102 64763
rect 42 64739 76 64755
rect 16 64719 38 64725
rect 42 64716 76 64720
rect 80 64719 102 64725
rect 42 64686 46 64716
rect 72 64686 76 64716
rect 42 64605 46 64639
rect 72 64605 76 64639
rect -25 64568 25 64570
rect -8 64560 14 64567
rect -8 64559 17 64560
rect 25 64559 27 64568
rect -12 64552 38 64559
rect -12 64551 34 64552
rect -12 64547 8 64551
rect 0 64535 8 64547
rect 14 64535 34 64551
rect 0 64534 34 64535
rect 0 64527 38 64534
rect 14 64526 17 64527
rect 25 64518 27 64527
rect 42 64498 45 64588
rect 69 64573 80 64605
rect 107 64573 143 64601
rect 144 64573 148 64793
rect 332 64725 336 64793
rect 380 64763 462 64795
rect 463 64763 472 64797
rect 480 64763 497 64797
rect 378 64755 464 64763
rect 505 64755 507 64805
rect 514 64763 548 64797
rect 565 64763 582 64797
rect 607 64755 609 64805
rect 404 64739 438 64755
rect 400 64725 442 64726
rect 378 64719 404 64725
rect 442 64719 464 64725
rect 400 64718 404 64719
rect 174 64679 246 64687
rect 295 64684 300 64718
rect 324 64684 329 64718
rect 224 64649 226 64665
rect 196 64641 226 64649
rect 332 64647 336 64715
rect 367 64684 438 64718
rect 400 64677 404 64684
rect 454 64671 504 64673
rect 494 64667 548 64671
rect 494 64662 514 64667
rect 504 64647 506 64662
rect 196 64637 232 64641
rect 196 64607 204 64637
rect 216 64607 232 64637
rect 400 64639 404 64647
rect 107 64567 119 64573
rect 109 64539 119 64567
rect 129 64539 149 64573
rect 174 64569 181 64599
rect 224 64560 226 64607
rect 256 64599 328 64607
rect 332 64605 336 64635
rect 400 64605 408 64639
rect 434 64605 438 64639
rect 498 64637 506 64647
rect 514 64637 515 64657
rect 504 64621 506 64637
rect 525 64628 528 64662
rect 547 64637 548 64657
rect 557 64637 564 64647
rect 514 64621 530 64627
rect 532 64621 548 64627
rect 278 64569 305 64580
rect 42 64447 46 64481
rect 72 64447 76 64481
rect 38 64409 80 64410
rect 42 64368 76 64402
rect 79 64368 113 64402
rect 42 64289 46 64323
rect 72 64289 76 64323
rect -25 64252 25 64254
rect -8 64244 14 64251
rect -8 64243 17 64244
rect 25 64243 27 64252
rect -12 64236 38 64243
rect -12 64235 34 64236
rect -12 64231 8 64235
rect 0 64219 8 64231
rect 14 64219 34 64235
rect 0 64218 34 64219
rect 0 64211 38 64218
rect 14 64210 17 64211
rect 25 64202 27 64211
rect 42 64182 45 64272
rect 71 64241 80 64269
rect 69 64203 80 64241
rect 144 64231 148 64539
rect 196 64526 204 64560
rect 216 64526 232 64560
rect 244 64556 257 64560
rect 300 64556 308 64569
rect 332 64567 342 64605
rect 400 64597 404 64605
rect 336 64557 342 64567
rect 244 64532 291 64556
rect 244 64526 257 64532
rect 224 64479 226 64526
rect 278 64522 291 64532
rect 300 64532 329 64556
rect 332 64547 342 64557
rect 400 64557 409 64585
rect 562 64568 612 64570
rect 466 64559 497 64567
rect 565 64559 596 64567
rect 300 64522 321 64532
rect 300 64516 308 64522
rect 289 64506 308 64516
rect 196 64449 204 64479
rect 216 64449 232 64479
rect 196 64445 232 64449
rect 196 64437 226 64445
rect 300 64437 308 64506
rect 332 64513 351 64547
rect 361 64519 381 64547
rect 361 64513 375 64519
rect 400 64513 411 64557
rect 442 64552 500 64559
rect 466 64551 500 64552
rect 565 64551 599 64559
rect 497 64535 500 64551
rect 596 64535 599 64551
rect 466 64534 500 64535
rect 442 64527 500 64534
rect 565 64527 599 64535
rect 612 64518 614 64568
rect 332 64489 342 64513
rect 336 64477 342 64489
rect 224 64421 226 64437
rect 332 64409 342 64477
rect 400 64481 404 64489
rect 400 64447 408 64481
rect 434 64447 438 64481
rect 454 64465 504 64467
rect 504 64449 506 64465
rect 514 64459 530 64465
rect 532 64459 548 64465
rect 525 64449 548 64458
rect 400 64439 404 64447
rect 498 64439 506 64449
rect 504 64415 506 64439
rect 514 64429 515 64449
rect 525 64424 528 64449
rect 547 64429 548 64449
rect 557 64439 564 64449
rect 514 64415 548 64419
rect 151 64368 156 64402
rect 174 64399 246 64407
rect 256 64399 328 64407
rect 336 64401 342 64409
rect 400 64404 404 64409
rect 180 64371 185 64399
rect 174 64363 246 64371
rect 256 64363 328 64371
rect 332 64369 336 64399
rect 400 64370 438 64404
rect 224 64333 226 64349
rect 196 64325 226 64333
rect 196 64321 232 64325
rect 196 64291 204 64321
rect 216 64291 232 64321
rect 224 64244 226 64291
rect 300 64264 308 64333
rect 332 64331 342 64369
rect 400 64361 404 64370
rect 454 64355 504 64357
rect 494 64351 548 64355
rect 494 64346 514 64351
rect 504 64331 506 64346
rect 336 64319 342 64331
rect 289 64254 308 64264
rect 300 64248 308 64254
rect 332 64285 342 64319
rect 400 64323 404 64331
rect 400 64289 408 64323
rect 434 64289 438 64323
rect 498 64321 506 64331
rect 514 64321 515 64341
rect 504 64305 506 64321
rect 525 64312 528 64346
rect 547 64321 548 64341
rect 557 64321 564 64331
rect 514 64305 530 64311
rect 532 64305 548 64311
rect 332 64257 373 64285
rect 332 64251 351 64257
rect 107 64197 119 64231
rect 129 64197 149 64231
rect 196 64210 204 64244
rect 216 64210 232 64244
rect 244 64238 257 64244
rect 278 64238 291 64248
rect 244 64214 291 64238
rect 300 64238 321 64248
rect 336 64241 351 64251
rect 300 64214 329 64238
rect 332 64223 351 64241
rect 361 64251 375 64257
rect 400 64251 411 64289
rect 562 64252 612 64254
rect 361 64223 381 64251
rect 400 64223 409 64251
rect 466 64243 497 64251
rect 565 64243 596 64251
rect 442 64236 500 64243
rect 466 64235 500 64236
rect 565 64235 599 64243
rect 244 64210 257 64214
rect 42 64131 46 64165
rect 72 64131 76 64165
rect 42 64084 76 64088
rect 42 64069 46 64084
rect 72 64069 76 64084
rect 38 64051 80 64069
rect 16 64045 102 64051
rect 144 64045 148 64197
rect 174 64173 181 64201
rect 224 64163 226 64210
rect 300 64201 308 64214
rect 278 64190 305 64201
rect 332 64173 342 64223
rect 400 64203 404 64223
rect 497 64219 500 64235
rect 596 64219 599 64235
rect 466 64218 500 64219
rect 442 64211 500 64218
rect 565 64211 599 64219
rect 612 64202 614 64252
rect 256 64163 328 64171
rect 336 64165 342 64173
rect 400 64165 404 64173
rect 196 64133 204 64163
rect 216 64133 232 64163
rect 196 64129 232 64133
rect 196 64121 226 64129
rect 224 64105 226 64121
rect 332 64093 336 64161
rect 400 64131 408 64165
rect 434 64131 438 64165
rect 454 64149 504 64151
rect 504 64133 506 64149
rect 514 64143 530 64149
rect 532 64143 548 64149
rect 525 64133 548 64142
rect 400 64123 404 64131
rect 498 64123 506 64133
rect 504 64099 506 64123
rect 514 64113 515 64133
rect 525 64108 528 64133
rect 547 64113 548 64133
rect 557 64123 564 64133
rect 514 64099 548 64103
rect 400 64093 442 64094
rect 174 64083 246 64091
rect 400 64086 404 64093
rect 295 64052 300 64086
rect 324 64052 329 64086
rect 367 64069 438 64086
rect 367 64052 442 64069
rect 400 64051 442 64052
rect 378 64045 464 64051
rect 38 64029 80 64045
rect 400 64029 442 64045
rect -25 64015 25 64017
rect 42 64015 76 64029
rect 404 64015 438 64029
rect 455 64015 505 64017
rect 557 64015 607 64017
rect 16 64007 102 64015
rect 378 64007 464 64015
rect 8 63973 17 64007
rect 18 64005 51 64007
rect 80 64005 100 64007
rect 18 63973 100 64005
rect 380 64005 404 64007
rect 429 64005 438 64007
rect 442 64005 462 64007
rect 16 63965 102 63973
rect 42 63949 76 63965
rect 16 63929 38 63935
rect 42 63926 76 63930
rect 80 63929 102 63935
rect 42 63896 46 63926
rect 72 63896 76 63926
rect 42 63815 46 63849
rect 72 63815 76 63849
rect -25 63778 25 63780
rect -8 63770 14 63777
rect -8 63769 17 63770
rect 25 63769 27 63778
rect -12 63762 38 63769
rect -12 63761 34 63762
rect -12 63757 8 63761
rect 0 63745 8 63757
rect 14 63745 34 63761
rect 0 63744 34 63745
rect 0 63737 38 63744
rect 14 63736 17 63737
rect 25 63728 27 63737
rect 42 63708 45 63798
rect 69 63783 80 63815
rect 107 63783 143 63811
rect 144 63783 148 64003
rect 332 63935 336 64003
rect 380 63973 462 64005
rect 463 63973 472 64007
rect 480 63973 497 64007
rect 378 63965 464 63973
rect 505 63965 507 64015
rect 514 63973 548 64007
rect 565 63973 582 64007
rect 607 63965 609 64015
rect 404 63949 438 63965
rect 400 63935 442 63936
rect 378 63929 404 63935
rect 442 63929 464 63935
rect 400 63928 404 63929
rect 174 63889 246 63897
rect 295 63894 300 63928
rect 324 63894 329 63928
rect 224 63859 226 63875
rect 196 63851 226 63859
rect 332 63857 336 63925
rect 367 63894 438 63928
rect 400 63887 404 63894
rect 454 63881 504 63883
rect 494 63877 548 63881
rect 494 63872 514 63877
rect 504 63857 506 63872
rect 196 63847 232 63851
rect 196 63817 204 63847
rect 216 63817 232 63847
rect 400 63849 404 63857
rect 107 63777 119 63783
rect 109 63749 119 63777
rect 129 63749 149 63783
rect 174 63779 181 63809
rect 224 63770 226 63817
rect 256 63809 328 63817
rect 332 63815 336 63845
rect 400 63815 408 63849
rect 434 63815 438 63849
rect 498 63847 506 63857
rect 514 63847 515 63867
rect 504 63831 506 63847
rect 525 63838 528 63872
rect 547 63847 548 63867
rect 557 63847 564 63857
rect 514 63831 530 63837
rect 532 63831 548 63837
rect 278 63779 305 63790
rect 42 63657 46 63691
rect 72 63657 76 63691
rect 38 63619 80 63620
rect 42 63578 76 63612
rect 79 63578 113 63612
rect 42 63499 46 63533
rect 72 63499 76 63533
rect -25 63462 25 63464
rect -8 63454 14 63461
rect -8 63453 17 63454
rect 25 63453 27 63462
rect -12 63446 38 63453
rect -12 63445 34 63446
rect -12 63441 8 63445
rect 0 63429 8 63441
rect 14 63429 34 63445
rect 0 63428 34 63429
rect 0 63421 38 63428
rect 14 63420 17 63421
rect 25 63412 27 63421
rect 42 63392 45 63482
rect 71 63451 80 63479
rect 69 63413 80 63451
rect 144 63441 148 63749
rect 196 63736 204 63770
rect 216 63736 232 63770
rect 244 63766 257 63770
rect 300 63766 308 63779
rect 332 63777 342 63815
rect 400 63807 404 63815
rect 336 63767 342 63777
rect 244 63742 291 63766
rect 244 63736 257 63742
rect 224 63689 226 63736
rect 278 63732 291 63742
rect 300 63742 329 63766
rect 332 63757 342 63767
rect 400 63767 409 63795
rect 562 63778 612 63780
rect 466 63769 497 63777
rect 565 63769 596 63777
rect 300 63732 321 63742
rect 300 63726 308 63732
rect 289 63716 308 63726
rect 196 63659 204 63689
rect 216 63659 232 63689
rect 196 63655 232 63659
rect 196 63647 226 63655
rect 300 63647 308 63716
rect 332 63723 351 63757
rect 361 63729 381 63757
rect 361 63723 375 63729
rect 400 63723 411 63767
rect 442 63762 500 63769
rect 466 63761 500 63762
rect 565 63761 599 63769
rect 497 63745 500 63761
rect 596 63745 599 63761
rect 466 63744 500 63745
rect 442 63737 500 63744
rect 565 63737 599 63745
rect 612 63728 614 63778
rect 332 63699 342 63723
rect 336 63687 342 63699
rect 224 63631 226 63647
rect 332 63619 342 63687
rect 400 63691 404 63699
rect 400 63657 408 63691
rect 434 63657 438 63691
rect 454 63675 504 63677
rect 504 63659 506 63675
rect 514 63669 530 63675
rect 532 63669 548 63675
rect 525 63659 548 63668
rect 400 63649 404 63657
rect 498 63649 506 63659
rect 504 63625 506 63649
rect 514 63639 515 63659
rect 525 63634 528 63659
rect 547 63639 548 63659
rect 557 63649 564 63659
rect 514 63625 548 63629
rect 151 63578 156 63612
rect 174 63609 246 63617
rect 256 63609 328 63617
rect 336 63611 342 63619
rect 400 63614 404 63619
rect 180 63581 185 63609
rect 174 63573 246 63581
rect 256 63573 328 63581
rect 332 63579 336 63609
rect 400 63580 438 63614
rect 224 63543 226 63559
rect 196 63535 226 63543
rect 196 63531 232 63535
rect 196 63501 204 63531
rect 216 63501 232 63531
rect 224 63454 226 63501
rect 300 63474 308 63543
rect 332 63541 342 63579
rect 400 63571 404 63580
rect 454 63565 504 63567
rect 494 63561 548 63565
rect 494 63556 514 63561
rect 504 63541 506 63556
rect 336 63529 342 63541
rect 289 63464 308 63474
rect 300 63458 308 63464
rect 332 63495 342 63529
rect 400 63533 404 63541
rect 400 63499 408 63533
rect 434 63499 438 63533
rect 498 63531 506 63541
rect 514 63531 515 63551
rect 504 63515 506 63531
rect 525 63522 528 63556
rect 547 63531 548 63551
rect 557 63531 564 63541
rect 514 63515 530 63521
rect 532 63515 548 63521
rect 332 63467 373 63495
rect 332 63461 351 63467
rect 107 63407 119 63441
rect 129 63407 149 63441
rect 196 63420 204 63454
rect 216 63420 232 63454
rect 244 63448 257 63454
rect 278 63448 291 63458
rect 244 63424 291 63448
rect 300 63448 321 63458
rect 336 63451 351 63461
rect 300 63424 329 63448
rect 332 63433 351 63451
rect 361 63461 375 63467
rect 400 63461 411 63499
rect 562 63462 612 63464
rect 361 63433 381 63461
rect 400 63433 409 63461
rect 466 63453 497 63461
rect 565 63453 596 63461
rect 442 63446 500 63453
rect 466 63445 500 63446
rect 565 63445 599 63453
rect 244 63420 257 63424
rect 42 63341 46 63375
rect 72 63341 76 63375
rect 42 63294 76 63298
rect 42 63279 46 63294
rect 72 63279 76 63294
rect 38 63261 80 63279
rect 16 63255 102 63261
rect 144 63255 148 63407
rect 174 63383 181 63411
rect 224 63373 226 63420
rect 300 63411 308 63424
rect 278 63400 305 63411
rect 332 63383 342 63433
rect 400 63413 404 63433
rect 497 63429 500 63445
rect 596 63429 599 63445
rect 466 63428 500 63429
rect 442 63421 500 63428
rect 565 63421 599 63429
rect 612 63412 614 63462
rect 256 63373 328 63381
rect 336 63375 342 63383
rect 400 63375 404 63383
rect 196 63343 204 63373
rect 216 63343 232 63373
rect 196 63339 232 63343
rect 196 63331 226 63339
rect 224 63315 226 63331
rect 332 63303 336 63371
rect 400 63341 408 63375
rect 434 63341 438 63375
rect 454 63359 504 63361
rect 504 63343 506 63359
rect 514 63353 530 63359
rect 532 63353 548 63359
rect 525 63343 548 63352
rect 400 63333 404 63341
rect 498 63333 506 63343
rect 504 63309 506 63333
rect 514 63323 515 63343
rect 525 63318 528 63343
rect 547 63323 548 63343
rect 557 63333 564 63343
rect 514 63309 548 63313
rect 400 63303 442 63304
rect 174 63293 246 63301
rect 400 63296 404 63303
rect 295 63262 300 63296
rect 324 63262 329 63296
rect 367 63279 438 63296
rect 367 63262 442 63279
rect 400 63261 442 63262
rect 378 63255 464 63261
rect 38 63239 80 63255
rect 400 63239 442 63255
rect -25 63225 25 63227
rect 42 63225 76 63239
rect 404 63225 438 63239
rect 455 63225 505 63227
rect 557 63225 607 63227
rect 16 63217 102 63225
rect 378 63217 464 63225
rect 8 63183 17 63217
rect 18 63215 51 63217
rect 80 63215 100 63217
rect 18 63183 100 63215
rect 380 63215 404 63217
rect 429 63215 438 63217
rect 442 63215 462 63217
rect 16 63175 102 63183
rect 42 63159 76 63175
rect 16 63139 38 63145
rect 42 63136 76 63140
rect 80 63139 102 63145
rect 42 63106 46 63136
rect 72 63106 76 63136
rect 42 63025 46 63059
rect 72 63025 76 63059
rect -25 62988 25 62990
rect -8 62980 14 62987
rect -8 62979 17 62980
rect 25 62979 27 62988
rect -12 62972 38 62979
rect -12 62971 34 62972
rect -12 62967 8 62971
rect 0 62955 8 62967
rect 14 62955 34 62971
rect 0 62954 34 62955
rect 0 62947 38 62954
rect 14 62946 17 62947
rect 25 62938 27 62947
rect 42 62918 45 63008
rect 69 62993 80 63025
rect 107 62993 143 63021
rect 144 62993 148 63213
rect 332 63145 336 63213
rect 380 63183 462 63215
rect 463 63183 472 63217
rect 480 63183 497 63217
rect 378 63175 464 63183
rect 505 63175 507 63225
rect 514 63183 548 63217
rect 565 63183 582 63217
rect 607 63175 609 63225
rect 404 63159 438 63175
rect 400 63145 442 63146
rect 378 63139 404 63145
rect 442 63139 464 63145
rect 400 63138 404 63139
rect 174 63099 246 63107
rect 295 63104 300 63138
rect 324 63104 329 63138
rect 224 63069 226 63085
rect 196 63061 226 63069
rect 332 63067 336 63135
rect 367 63104 438 63138
rect 400 63097 404 63104
rect 454 63091 504 63093
rect 494 63087 548 63091
rect 494 63082 514 63087
rect 504 63067 506 63082
rect 196 63057 232 63061
rect 196 63027 204 63057
rect 216 63027 232 63057
rect 400 63059 404 63067
rect 107 62987 119 62993
rect 109 62959 119 62987
rect 129 62959 149 62993
rect 174 62989 181 63019
rect 224 62980 226 63027
rect 256 63019 328 63027
rect 332 63025 336 63055
rect 400 63025 408 63059
rect 434 63025 438 63059
rect 498 63057 506 63067
rect 514 63057 515 63077
rect 504 63041 506 63057
rect 525 63048 528 63082
rect 547 63057 548 63077
rect 557 63057 564 63067
rect 514 63041 530 63047
rect 532 63041 548 63047
rect 278 62989 305 63000
rect 42 62867 46 62901
rect 72 62867 76 62901
rect 38 62829 80 62830
rect 42 62788 76 62822
rect 79 62788 113 62822
rect 42 62709 46 62743
rect 72 62709 76 62743
rect -25 62672 25 62674
rect -8 62664 14 62671
rect -8 62663 17 62664
rect 25 62663 27 62672
rect -12 62656 38 62663
rect -12 62655 34 62656
rect -12 62651 8 62655
rect 0 62639 8 62651
rect 14 62639 34 62655
rect 0 62638 34 62639
rect 0 62631 38 62638
rect 14 62630 17 62631
rect 25 62622 27 62631
rect 42 62602 45 62692
rect 71 62661 80 62689
rect 69 62623 80 62661
rect 144 62651 148 62959
rect 196 62946 204 62980
rect 216 62946 232 62980
rect 244 62976 257 62980
rect 300 62976 308 62989
rect 332 62987 342 63025
rect 400 63017 404 63025
rect 336 62977 342 62987
rect 244 62952 291 62976
rect 244 62946 257 62952
rect 224 62899 226 62946
rect 278 62942 291 62952
rect 300 62952 329 62976
rect 332 62967 342 62977
rect 400 62977 409 63005
rect 562 62988 612 62990
rect 466 62979 497 62987
rect 565 62979 596 62987
rect 300 62942 321 62952
rect 300 62936 308 62942
rect 289 62926 308 62936
rect 196 62869 204 62899
rect 216 62869 232 62899
rect 196 62865 232 62869
rect 196 62857 226 62865
rect 300 62857 308 62926
rect 332 62933 351 62967
rect 361 62939 381 62967
rect 361 62933 375 62939
rect 400 62933 411 62977
rect 442 62972 500 62979
rect 466 62971 500 62972
rect 565 62971 599 62979
rect 497 62955 500 62971
rect 596 62955 599 62971
rect 466 62954 500 62955
rect 442 62947 500 62954
rect 565 62947 599 62955
rect 612 62938 614 62988
rect 332 62909 342 62933
rect 336 62897 342 62909
rect 224 62841 226 62857
rect 332 62829 342 62897
rect 400 62901 404 62909
rect 400 62867 408 62901
rect 434 62867 438 62901
rect 454 62885 504 62887
rect 504 62869 506 62885
rect 514 62879 530 62885
rect 532 62879 548 62885
rect 525 62869 548 62878
rect 400 62859 404 62867
rect 498 62859 506 62869
rect 504 62835 506 62859
rect 514 62849 515 62869
rect 525 62844 528 62869
rect 547 62849 548 62869
rect 557 62859 564 62869
rect 514 62835 548 62839
rect 151 62788 156 62822
rect 174 62819 246 62827
rect 256 62819 328 62827
rect 336 62821 342 62829
rect 400 62824 404 62829
rect 180 62791 185 62819
rect 174 62783 246 62791
rect 256 62783 328 62791
rect 332 62789 336 62819
rect 400 62790 438 62824
rect 224 62753 226 62769
rect 196 62745 226 62753
rect 196 62741 232 62745
rect 196 62711 204 62741
rect 216 62711 232 62741
rect 224 62664 226 62711
rect 300 62684 308 62753
rect 332 62751 342 62789
rect 400 62781 404 62790
rect 454 62775 504 62777
rect 494 62771 548 62775
rect 494 62766 514 62771
rect 504 62751 506 62766
rect 336 62739 342 62751
rect 289 62674 308 62684
rect 300 62668 308 62674
rect 332 62705 342 62739
rect 400 62743 404 62751
rect 400 62709 408 62743
rect 434 62709 438 62743
rect 498 62741 506 62751
rect 514 62741 515 62761
rect 504 62725 506 62741
rect 525 62732 528 62766
rect 547 62741 548 62761
rect 557 62741 564 62751
rect 514 62725 530 62731
rect 532 62725 548 62731
rect 332 62677 373 62705
rect 332 62671 351 62677
rect 107 62617 119 62651
rect 129 62617 149 62651
rect 196 62630 204 62664
rect 216 62630 232 62664
rect 244 62658 257 62664
rect 278 62658 291 62668
rect 244 62634 291 62658
rect 300 62658 321 62668
rect 336 62661 351 62671
rect 300 62634 329 62658
rect 332 62643 351 62661
rect 361 62671 375 62677
rect 400 62671 411 62709
rect 562 62672 612 62674
rect 361 62643 381 62671
rect 400 62643 409 62671
rect 466 62663 497 62671
rect 565 62663 596 62671
rect 442 62656 500 62663
rect 466 62655 500 62656
rect 565 62655 599 62663
rect 244 62630 257 62634
rect 42 62551 46 62585
rect 72 62551 76 62585
rect 42 62504 76 62508
rect 42 62489 46 62504
rect 72 62489 76 62504
rect 38 62471 80 62489
rect 16 62465 102 62471
rect 144 62465 148 62617
rect 174 62593 181 62621
rect 224 62583 226 62630
rect 300 62621 308 62634
rect 278 62610 305 62621
rect 332 62593 342 62643
rect 400 62623 404 62643
rect 497 62639 500 62655
rect 596 62639 599 62655
rect 466 62638 500 62639
rect 442 62631 500 62638
rect 565 62631 599 62639
rect 612 62622 614 62672
rect 256 62583 328 62591
rect 336 62585 342 62593
rect 400 62585 404 62593
rect 196 62553 204 62583
rect 216 62553 232 62583
rect 196 62549 232 62553
rect 196 62541 226 62549
rect 224 62525 226 62541
rect 332 62513 336 62581
rect 400 62551 408 62585
rect 434 62551 438 62585
rect 454 62569 504 62571
rect 504 62553 506 62569
rect 514 62563 530 62569
rect 532 62563 548 62569
rect 525 62553 548 62562
rect 400 62543 404 62551
rect 498 62543 506 62553
rect 504 62519 506 62543
rect 514 62533 515 62553
rect 525 62528 528 62553
rect 547 62533 548 62553
rect 557 62543 564 62553
rect 514 62519 548 62523
rect 400 62513 442 62514
rect 174 62503 246 62511
rect 400 62506 404 62513
rect 295 62472 300 62506
rect 324 62472 329 62506
rect 367 62489 438 62506
rect 367 62472 442 62489
rect 400 62471 442 62472
rect 378 62465 464 62471
rect 38 62449 80 62465
rect 400 62449 442 62465
rect -25 62435 25 62437
rect 42 62435 76 62449
rect 404 62435 438 62449
rect 455 62435 505 62437
rect 557 62435 607 62437
rect 16 62427 102 62435
rect 378 62427 464 62435
rect 8 62393 17 62427
rect 18 62425 51 62427
rect 80 62425 100 62427
rect 18 62393 100 62425
rect 380 62425 404 62427
rect 429 62425 438 62427
rect 442 62425 462 62427
rect 16 62385 102 62393
rect 42 62369 76 62385
rect 16 62349 38 62355
rect 42 62346 76 62350
rect 80 62349 102 62355
rect 42 62316 46 62346
rect 72 62316 76 62346
rect 42 62235 46 62269
rect 72 62235 76 62269
rect -25 62198 25 62200
rect -8 62190 14 62197
rect -8 62189 17 62190
rect 25 62189 27 62198
rect -12 62182 38 62189
rect -12 62181 34 62182
rect -12 62177 8 62181
rect 0 62165 8 62177
rect 14 62165 34 62181
rect 0 62164 34 62165
rect 0 62157 38 62164
rect 14 62156 17 62157
rect 25 62148 27 62157
rect 42 62128 45 62218
rect 69 62203 80 62235
rect 107 62203 143 62231
rect 144 62203 148 62423
rect 332 62355 336 62423
rect 380 62393 462 62425
rect 463 62393 472 62427
rect 480 62393 497 62427
rect 378 62385 464 62393
rect 505 62385 507 62435
rect 514 62393 548 62427
rect 565 62393 582 62427
rect 607 62385 609 62435
rect 404 62369 438 62385
rect 400 62355 442 62356
rect 378 62349 404 62355
rect 442 62349 464 62355
rect 400 62348 404 62349
rect 174 62309 246 62317
rect 295 62314 300 62348
rect 324 62314 329 62348
rect 224 62279 226 62295
rect 196 62271 226 62279
rect 332 62277 336 62345
rect 367 62314 438 62348
rect 400 62307 404 62314
rect 454 62301 504 62303
rect 494 62297 548 62301
rect 494 62292 514 62297
rect 504 62277 506 62292
rect 196 62267 232 62271
rect 196 62237 204 62267
rect 216 62237 232 62267
rect 400 62269 404 62277
rect 107 62197 119 62203
rect 109 62169 119 62197
rect 129 62169 149 62203
rect 174 62199 181 62229
rect 224 62190 226 62237
rect 256 62229 328 62237
rect 332 62235 336 62265
rect 400 62235 408 62269
rect 434 62235 438 62269
rect 498 62267 506 62277
rect 514 62267 515 62287
rect 504 62251 506 62267
rect 525 62258 528 62292
rect 547 62267 548 62287
rect 557 62267 564 62277
rect 514 62251 530 62257
rect 532 62251 548 62257
rect 278 62199 305 62210
rect 42 62077 46 62111
rect 72 62077 76 62111
rect 38 62039 80 62040
rect 42 61998 76 62032
rect 79 61998 113 62032
rect 42 61919 46 61953
rect 72 61919 76 61953
rect -25 61882 25 61884
rect -8 61874 14 61881
rect -8 61873 17 61874
rect 25 61873 27 61882
rect -12 61866 38 61873
rect -12 61865 34 61866
rect -12 61861 8 61865
rect 0 61849 8 61861
rect 14 61849 34 61865
rect 0 61848 34 61849
rect 0 61841 38 61848
rect 14 61840 17 61841
rect 25 61832 27 61841
rect 42 61812 45 61902
rect 71 61871 80 61899
rect 69 61833 80 61871
rect 144 61861 148 62169
rect 196 62156 204 62190
rect 216 62156 232 62190
rect 244 62186 257 62190
rect 300 62186 308 62199
rect 332 62197 342 62235
rect 400 62227 404 62235
rect 336 62187 342 62197
rect 244 62162 291 62186
rect 244 62156 257 62162
rect 224 62109 226 62156
rect 278 62152 291 62162
rect 300 62162 329 62186
rect 332 62177 342 62187
rect 400 62187 409 62215
rect 562 62198 612 62200
rect 466 62189 497 62197
rect 565 62189 596 62197
rect 300 62152 321 62162
rect 300 62146 308 62152
rect 289 62136 308 62146
rect 196 62079 204 62109
rect 216 62079 232 62109
rect 196 62075 232 62079
rect 196 62067 226 62075
rect 300 62067 308 62136
rect 332 62143 351 62177
rect 361 62149 381 62177
rect 361 62143 375 62149
rect 400 62143 411 62187
rect 442 62182 500 62189
rect 466 62181 500 62182
rect 565 62181 599 62189
rect 497 62165 500 62181
rect 596 62165 599 62181
rect 466 62164 500 62165
rect 442 62157 500 62164
rect 565 62157 599 62165
rect 612 62148 614 62198
rect 332 62119 342 62143
rect 336 62107 342 62119
rect 224 62051 226 62067
rect 332 62039 342 62107
rect 400 62111 404 62119
rect 400 62077 408 62111
rect 434 62077 438 62111
rect 454 62095 504 62097
rect 504 62079 506 62095
rect 514 62089 530 62095
rect 532 62089 548 62095
rect 525 62079 548 62088
rect 400 62069 404 62077
rect 498 62069 506 62079
rect 504 62045 506 62069
rect 514 62059 515 62079
rect 525 62054 528 62079
rect 547 62059 548 62079
rect 557 62069 564 62079
rect 514 62045 548 62049
rect 151 61998 156 62032
rect 174 62029 246 62037
rect 256 62029 328 62037
rect 336 62031 342 62039
rect 400 62034 404 62039
rect 180 62001 185 62029
rect 174 61993 246 62001
rect 256 61993 328 62001
rect 332 61999 336 62029
rect 400 62000 438 62034
rect 224 61963 226 61979
rect 196 61955 226 61963
rect 196 61951 232 61955
rect 196 61921 204 61951
rect 216 61921 232 61951
rect 224 61874 226 61921
rect 300 61894 308 61963
rect 332 61961 342 61999
rect 400 61991 404 62000
rect 454 61985 504 61987
rect 494 61981 548 61985
rect 494 61976 514 61981
rect 504 61961 506 61976
rect 336 61949 342 61961
rect 289 61884 308 61894
rect 300 61878 308 61884
rect 332 61915 342 61949
rect 400 61953 404 61961
rect 400 61919 408 61953
rect 434 61919 438 61953
rect 498 61951 506 61961
rect 514 61951 515 61971
rect 504 61935 506 61951
rect 525 61942 528 61976
rect 547 61951 548 61971
rect 557 61951 564 61961
rect 514 61935 530 61941
rect 532 61935 548 61941
rect 332 61887 373 61915
rect 332 61881 351 61887
rect 107 61827 119 61861
rect 129 61827 149 61861
rect 196 61840 204 61874
rect 216 61840 232 61874
rect 244 61868 257 61874
rect 278 61868 291 61878
rect 244 61844 291 61868
rect 300 61868 321 61878
rect 336 61871 351 61881
rect 300 61844 329 61868
rect 332 61853 351 61871
rect 361 61881 375 61887
rect 400 61881 411 61919
rect 562 61882 612 61884
rect 361 61853 381 61881
rect 400 61853 409 61881
rect 466 61873 497 61881
rect 565 61873 596 61881
rect 442 61866 500 61873
rect 466 61865 500 61866
rect 565 61865 599 61873
rect 244 61840 257 61844
rect 42 61761 46 61795
rect 72 61761 76 61795
rect 42 61714 76 61718
rect 42 61699 46 61714
rect 72 61699 76 61714
rect 38 61681 80 61699
rect 16 61675 102 61681
rect 144 61675 148 61827
rect 174 61803 181 61831
rect 224 61793 226 61840
rect 300 61831 308 61844
rect 278 61820 305 61831
rect 332 61803 342 61853
rect 400 61833 404 61853
rect 497 61849 500 61865
rect 596 61849 599 61865
rect 466 61848 500 61849
rect 442 61841 500 61848
rect 565 61841 599 61849
rect 612 61832 614 61882
rect 256 61793 328 61801
rect 336 61795 342 61803
rect 400 61795 404 61803
rect 196 61763 204 61793
rect 216 61763 232 61793
rect 196 61759 232 61763
rect 196 61751 226 61759
rect 224 61735 226 61751
rect 332 61723 336 61791
rect 400 61761 408 61795
rect 434 61761 438 61795
rect 454 61779 504 61781
rect 504 61763 506 61779
rect 514 61773 530 61779
rect 532 61773 548 61779
rect 525 61763 548 61772
rect 400 61753 404 61761
rect 498 61753 506 61763
rect 504 61729 506 61753
rect 514 61743 515 61763
rect 525 61738 528 61763
rect 547 61743 548 61763
rect 557 61753 564 61763
rect 514 61729 548 61733
rect 400 61723 442 61724
rect 174 61713 246 61721
rect 400 61716 404 61723
rect 295 61682 300 61716
rect 324 61682 329 61716
rect 367 61699 438 61716
rect 367 61682 442 61699
rect 400 61681 442 61682
rect 378 61675 464 61681
rect 38 61659 80 61675
rect 400 61659 442 61675
rect -25 61645 25 61647
rect 42 61645 76 61659
rect 404 61645 438 61659
rect 455 61645 505 61647
rect 557 61645 607 61647
rect 16 61637 102 61645
rect 378 61637 464 61645
rect 8 61603 17 61637
rect 18 61635 51 61637
rect 80 61635 100 61637
rect 18 61603 100 61635
rect 380 61635 404 61637
rect 429 61635 438 61637
rect 442 61635 462 61637
rect 16 61595 102 61603
rect 42 61579 76 61595
rect 16 61559 38 61565
rect 42 61556 76 61560
rect 80 61559 102 61565
rect 42 61526 46 61556
rect 72 61526 76 61556
rect 42 61445 46 61479
rect 72 61445 76 61479
rect -25 61408 25 61410
rect -8 61400 14 61407
rect -8 61399 17 61400
rect 25 61399 27 61408
rect -12 61392 38 61399
rect -12 61391 34 61392
rect -12 61387 8 61391
rect 0 61375 8 61387
rect 14 61375 34 61391
rect 0 61374 34 61375
rect 0 61367 38 61374
rect 14 61366 17 61367
rect 25 61358 27 61367
rect 42 61338 45 61428
rect 69 61413 80 61445
rect 107 61413 143 61441
rect 144 61413 148 61633
rect 332 61565 336 61633
rect 380 61603 462 61635
rect 463 61603 472 61637
rect 480 61603 497 61637
rect 378 61595 464 61603
rect 505 61595 507 61645
rect 514 61603 548 61637
rect 565 61603 582 61637
rect 607 61595 609 61645
rect 404 61579 438 61595
rect 400 61565 442 61566
rect 378 61559 404 61565
rect 442 61559 464 61565
rect 400 61558 404 61559
rect 174 61519 246 61527
rect 295 61524 300 61558
rect 324 61524 329 61558
rect 224 61489 226 61505
rect 196 61481 226 61489
rect 332 61487 336 61555
rect 367 61524 438 61558
rect 400 61517 404 61524
rect 454 61511 504 61513
rect 494 61507 548 61511
rect 494 61502 514 61507
rect 504 61487 506 61502
rect 196 61477 232 61481
rect 196 61447 204 61477
rect 216 61447 232 61477
rect 400 61479 404 61487
rect 107 61407 119 61413
rect 109 61379 119 61407
rect 129 61379 149 61413
rect 174 61409 181 61439
rect 224 61400 226 61447
rect 256 61439 328 61447
rect 332 61445 336 61475
rect 400 61445 408 61479
rect 434 61445 438 61479
rect 498 61477 506 61487
rect 514 61477 515 61497
rect 504 61461 506 61477
rect 525 61468 528 61502
rect 547 61477 548 61497
rect 557 61477 564 61487
rect 514 61461 530 61467
rect 532 61461 548 61467
rect 278 61409 305 61420
rect 42 61287 46 61321
rect 72 61287 76 61321
rect 38 61249 80 61250
rect 42 61208 76 61242
rect 79 61208 113 61242
rect 42 61129 46 61163
rect 72 61129 76 61163
rect -25 61092 25 61094
rect -8 61084 14 61091
rect -8 61083 17 61084
rect 25 61083 27 61092
rect -12 61076 38 61083
rect -12 61075 34 61076
rect -12 61071 8 61075
rect 0 61059 8 61071
rect 14 61059 34 61075
rect 0 61058 34 61059
rect 0 61051 38 61058
rect 14 61050 17 61051
rect 25 61042 27 61051
rect 42 61022 45 61112
rect 71 61081 80 61109
rect 69 61043 80 61081
rect 144 61071 148 61379
rect 196 61366 204 61400
rect 216 61366 232 61400
rect 244 61396 257 61400
rect 300 61396 308 61409
rect 332 61407 342 61445
rect 400 61437 404 61445
rect 336 61397 342 61407
rect 244 61372 291 61396
rect 244 61366 257 61372
rect 224 61319 226 61366
rect 278 61362 291 61372
rect 300 61372 329 61396
rect 332 61387 342 61397
rect 400 61397 409 61425
rect 562 61408 612 61410
rect 466 61399 497 61407
rect 565 61399 596 61407
rect 300 61362 321 61372
rect 300 61356 308 61362
rect 289 61346 308 61356
rect 196 61289 204 61319
rect 216 61289 232 61319
rect 196 61285 232 61289
rect 196 61277 226 61285
rect 300 61277 308 61346
rect 332 61353 351 61387
rect 361 61359 381 61387
rect 361 61353 375 61359
rect 400 61353 411 61397
rect 442 61392 500 61399
rect 466 61391 500 61392
rect 565 61391 599 61399
rect 497 61375 500 61391
rect 596 61375 599 61391
rect 466 61374 500 61375
rect 442 61367 500 61374
rect 565 61367 599 61375
rect 612 61358 614 61408
rect 332 61329 342 61353
rect 336 61317 342 61329
rect 224 61261 226 61277
rect 332 61249 342 61317
rect 400 61321 404 61329
rect 400 61287 408 61321
rect 434 61287 438 61321
rect 454 61305 504 61307
rect 504 61289 506 61305
rect 514 61299 530 61305
rect 532 61299 548 61305
rect 525 61289 548 61298
rect 400 61279 404 61287
rect 498 61279 506 61289
rect 504 61255 506 61279
rect 514 61269 515 61289
rect 525 61264 528 61289
rect 547 61269 548 61289
rect 557 61279 564 61289
rect 514 61255 548 61259
rect 151 61208 156 61242
rect 174 61239 246 61247
rect 256 61239 328 61247
rect 336 61241 342 61249
rect 400 61244 404 61249
rect 180 61211 185 61239
rect 174 61203 246 61211
rect 256 61203 328 61211
rect 332 61209 336 61239
rect 400 61210 438 61244
rect 224 61173 226 61189
rect 196 61165 226 61173
rect 196 61161 232 61165
rect 196 61131 204 61161
rect 216 61131 232 61161
rect 224 61084 226 61131
rect 300 61104 308 61173
rect 332 61171 342 61209
rect 400 61201 404 61210
rect 454 61195 504 61197
rect 494 61191 548 61195
rect 494 61186 514 61191
rect 504 61171 506 61186
rect 336 61159 342 61171
rect 289 61094 308 61104
rect 300 61088 308 61094
rect 332 61125 342 61159
rect 400 61163 404 61171
rect 400 61129 408 61163
rect 434 61129 438 61163
rect 498 61161 506 61171
rect 514 61161 515 61181
rect 504 61145 506 61161
rect 525 61152 528 61186
rect 547 61161 548 61181
rect 557 61161 564 61171
rect 514 61145 530 61151
rect 532 61145 548 61151
rect 332 61097 373 61125
rect 332 61091 351 61097
rect 107 61037 119 61071
rect 129 61037 149 61071
rect 196 61050 204 61084
rect 216 61050 232 61084
rect 244 61078 257 61084
rect 278 61078 291 61088
rect 244 61054 291 61078
rect 300 61078 321 61088
rect 336 61081 351 61091
rect 300 61054 329 61078
rect 332 61063 351 61081
rect 361 61091 375 61097
rect 400 61091 411 61129
rect 562 61092 612 61094
rect 361 61063 381 61091
rect 400 61063 409 61091
rect 466 61083 497 61091
rect 565 61083 596 61091
rect 442 61076 500 61083
rect 466 61075 500 61076
rect 565 61075 599 61083
rect 244 61050 257 61054
rect 42 60971 46 61005
rect 72 60971 76 61005
rect 42 60924 76 60928
rect 42 60909 46 60924
rect 72 60909 76 60924
rect 38 60891 80 60909
rect 16 60885 102 60891
rect 144 60885 148 61037
rect 174 61013 181 61041
rect 224 61003 226 61050
rect 300 61041 308 61054
rect 278 61030 305 61041
rect 332 61013 342 61063
rect 400 61043 404 61063
rect 497 61059 500 61075
rect 596 61059 599 61075
rect 466 61058 500 61059
rect 442 61051 500 61058
rect 565 61051 599 61059
rect 612 61042 614 61092
rect 256 61003 328 61011
rect 336 61005 342 61013
rect 400 61005 404 61013
rect 196 60973 204 61003
rect 216 60973 232 61003
rect 196 60969 232 60973
rect 196 60961 226 60969
rect 224 60945 226 60961
rect 332 60933 336 61001
rect 400 60971 408 61005
rect 434 60971 438 61005
rect 454 60989 504 60991
rect 504 60973 506 60989
rect 514 60983 530 60989
rect 532 60983 548 60989
rect 525 60973 548 60982
rect 400 60963 404 60971
rect 498 60963 506 60973
rect 504 60939 506 60963
rect 514 60953 515 60973
rect 525 60948 528 60973
rect 547 60953 548 60973
rect 557 60963 564 60973
rect 514 60939 548 60943
rect 400 60933 442 60934
rect 174 60923 246 60931
rect 400 60926 404 60933
rect 295 60892 300 60926
rect 324 60892 329 60926
rect 367 60909 438 60926
rect 367 60892 442 60909
rect 400 60891 442 60892
rect 378 60885 464 60891
rect 38 60869 80 60885
rect 400 60869 442 60885
rect -25 60855 25 60857
rect 42 60855 76 60869
rect 404 60855 438 60869
rect 455 60855 505 60857
rect 557 60855 607 60857
rect 16 60847 102 60855
rect 378 60847 464 60855
rect 8 60813 17 60847
rect 18 60845 51 60847
rect 80 60845 100 60847
rect 18 60813 100 60845
rect 380 60845 404 60847
rect 429 60845 438 60847
rect 442 60845 462 60847
rect 16 60805 102 60813
rect 42 60789 76 60805
rect 16 60769 38 60775
rect 42 60766 76 60770
rect 80 60769 102 60775
rect 42 60736 46 60766
rect 72 60736 76 60766
rect 42 60655 46 60689
rect 72 60655 76 60689
rect -25 60618 25 60620
rect -8 60610 14 60617
rect -8 60609 17 60610
rect 25 60609 27 60618
rect -12 60602 38 60609
rect -12 60601 34 60602
rect -12 60597 8 60601
rect 0 60585 8 60597
rect 14 60585 34 60601
rect 0 60584 34 60585
rect 0 60577 38 60584
rect 14 60576 17 60577
rect 25 60568 27 60577
rect 42 60548 45 60638
rect 69 60623 80 60655
rect 107 60623 143 60651
rect 144 60623 148 60843
rect 332 60775 336 60843
rect 380 60813 462 60845
rect 463 60813 472 60847
rect 480 60813 497 60847
rect 378 60805 464 60813
rect 505 60805 507 60855
rect 514 60813 548 60847
rect 565 60813 582 60847
rect 607 60805 609 60855
rect 404 60789 438 60805
rect 400 60775 442 60776
rect 378 60769 404 60775
rect 442 60769 464 60775
rect 400 60768 404 60769
rect 174 60729 246 60737
rect 295 60734 300 60768
rect 324 60734 329 60768
rect 224 60699 226 60715
rect 196 60691 226 60699
rect 332 60697 336 60765
rect 367 60734 438 60768
rect 400 60727 404 60734
rect 454 60721 504 60723
rect 494 60717 548 60721
rect 494 60712 514 60717
rect 504 60697 506 60712
rect 196 60687 232 60691
rect 196 60657 204 60687
rect 216 60657 232 60687
rect 400 60689 404 60697
rect 107 60617 119 60623
rect 109 60589 119 60617
rect 129 60589 149 60623
rect 174 60619 181 60649
rect 224 60610 226 60657
rect 256 60649 328 60657
rect 332 60655 336 60685
rect 400 60655 408 60689
rect 434 60655 438 60689
rect 498 60687 506 60697
rect 514 60687 515 60707
rect 504 60671 506 60687
rect 525 60678 528 60712
rect 547 60687 548 60707
rect 557 60687 564 60697
rect 514 60671 530 60677
rect 532 60671 548 60677
rect 278 60619 305 60630
rect 42 60497 46 60531
rect 72 60497 76 60531
rect 38 60459 80 60460
rect 42 60418 76 60452
rect 79 60418 113 60452
rect 42 60339 46 60373
rect 72 60339 76 60373
rect -25 60302 25 60304
rect -8 60294 14 60301
rect -8 60293 17 60294
rect 25 60293 27 60302
rect -12 60286 38 60293
rect -12 60285 34 60286
rect -12 60281 8 60285
rect 0 60269 8 60281
rect 14 60269 34 60285
rect 0 60268 34 60269
rect 0 60261 38 60268
rect 14 60260 17 60261
rect 25 60252 27 60261
rect 42 60232 45 60322
rect 71 60291 80 60319
rect 69 60253 80 60291
rect 144 60281 148 60589
rect 196 60576 204 60610
rect 216 60576 232 60610
rect 244 60606 257 60610
rect 300 60606 308 60619
rect 332 60617 342 60655
rect 400 60647 404 60655
rect 336 60607 342 60617
rect 244 60582 291 60606
rect 244 60576 257 60582
rect 224 60529 226 60576
rect 278 60572 291 60582
rect 300 60582 329 60606
rect 332 60597 342 60607
rect 400 60607 409 60635
rect 562 60618 612 60620
rect 466 60609 497 60617
rect 565 60609 596 60617
rect 300 60572 321 60582
rect 300 60566 308 60572
rect 289 60556 308 60566
rect 196 60499 204 60529
rect 216 60499 232 60529
rect 196 60495 232 60499
rect 196 60487 226 60495
rect 300 60487 308 60556
rect 332 60563 351 60597
rect 361 60569 381 60597
rect 361 60563 375 60569
rect 400 60563 411 60607
rect 442 60602 500 60609
rect 466 60601 500 60602
rect 565 60601 599 60609
rect 497 60585 500 60601
rect 596 60585 599 60601
rect 466 60584 500 60585
rect 442 60577 500 60584
rect 565 60577 599 60585
rect 612 60568 614 60618
rect 332 60539 342 60563
rect 336 60527 342 60539
rect 224 60471 226 60487
rect 332 60459 342 60527
rect 400 60531 404 60539
rect 400 60497 408 60531
rect 434 60497 438 60531
rect 454 60515 504 60517
rect 504 60499 506 60515
rect 514 60509 530 60515
rect 532 60509 548 60515
rect 525 60499 548 60508
rect 400 60489 404 60497
rect 498 60489 506 60499
rect 504 60465 506 60489
rect 514 60480 515 60499
rect 525 60474 528 60499
rect 547 60480 548 60499
rect 557 60489 564 60499
rect 514 60465 548 60469
rect 151 60418 156 60452
rect 174 60449 246 60457
rect 256 60449 328 60457
rect 336 60451 342 60459
rect 400 60454 404 60459
rect 180 60421 185 60449
rect 174 60413 246 60421
rect 256 60413 328 60421
rect 332 60419 336 60449
rect 400 60420 438 60454
rect 224 60383 226 60399
rect 196 60375 226 60383
rect 196 60371 232 60375
rect 196 60341 204 60371
rect 216 60341 232 60371
rect 224 60294 226 60341
rect 300 60314 308 60383
rect 332 60381 342 60419
rect 400 60411 404 60420
rect 454 60405 504 60407
rect 494 60401 548 60405
rect 494 60396 514 60401
rect 504 60381 506 60396
rect 336 60369 342 60381
rect 289 60304 308 60314
rect 300 60298 308 60304
rect 332 60335 342 60369
rect 400 60373 404 60381
rect 400 60339 408 60373
rect 434 60339 438 60373
rect 498 60371 506 60381
rect 514 60371 515 60391
rect 504 60355 506 60371
rect 525 60362 528 60396
rect 547 60371 548 60391
rect 557 60371 564 60381
rect 514 60355 530 60361
rect 532 60355 548 60361
rect 332 60307 373 60335
rect 332 60301 351 60307
rect 107 60247 119 60281
rect 129 60247 149 60281
rect 196 60260 204 60294
rect 216 60260 232 60294
rect 244 60288 257 60294
rect 278 60288 291 60298
rect 244 60264 291 60288
rect 300 60288 321 60298
rect 336 60291 351 60301
rect 300 60264 329 60288
rect 332 60273 351 60291
rect 361 60301 375 60307
rect 400 60301 411 60339
rect 562 60302 612 60304
rect 361 60273 381 60301
rect 400 60273 409 60301
rect 466 60293 497 60301
rect 565 60293 596 60301
rect 442 60286 500 60293
rect 466 60285 500 60286
rect 565 60285 599 60293
rect 244 60260 257 60264
rect 42 60181 46 60215
rect 72 60181 76 60215
rect 42 60134 76 60138
rect 42 60119 46 60134
rect 72 60119 76 60134
rect 38 60101 80 60119
rect 16 60095 102 60101
rect 144 60095 148 60247
rect 174 60223 181 60251
rect 224 60213 226 60260
rect 300 60251 308 60264
rect 278 60240 305 60251
rect 332 60223 342 60273
rect 400 60253 404 60273
rect 497 60269 500 60285
rect 596 60269 599 60285
rect 466 60268 500 60269
rect 442 60261 500 60268
rect 565 60261 599 60269
rect 612 60252 614 60302
rect 256 60213 328 60221
rect 336 60215 342 60223
rect 400 60215 404 60223
rect 196 60183 204 60213
rect 216 60183 232 60213
rect 196 60179 232 60183
rect 196 60171 226 60179
rect 224 60155 226 60171
rect 332 60143 336 60211
rect 400 60181 408 60215
rect 434 60181 438 60215
rect 454 60199 504 60201
rect 504 60183 506 60199
rect 514 60193 530 60199
rect 532 60193 548 60199
rect 525 60183 548 60192
rect 400 60173 404 60181
rect 498 60173 506 60183
rect 504 60149 506 60173
rect 514 60163 515 60183
rect 525 60158 528 60183
rect 547 60163 548 60183
rect 557 60173 564 60183
rect 514 60149 548 60153
rect 400 60143 442 60144
rect 174 60133 246 60141
rect 400 60136 404 60143
rect 295 60102 300 60136
rect 324 60102 329 60136
rect 367 60119 438 60136
rect 367 60102 442 60119
rect 400 60101 442 60102
rect 378 60095 464 60101
rect 38 60079 80 60095
rect 400 60079 442 60095
rect -25 60065 25 60067
rect 42 60065 76 60079
rect 404 60065 438 60079
rect 455 60065 505 60067
rect 557 60065 607 60067
rect 16 60057 102 60065
rect 378 60057 464 60065
rect 8 60023 17 60057
rect 18 60055 51 60057
rect 80 60055 100 60057
rect 18 60023 100 60055
rect 380 60055 404 60057
rect 429 60055 438 60057
rect 442 60055 462 60057
rect 16 60015 102 60023
rect 42 59999 76 60015
rect 16 59979 38 59985
rect 42 59976 76 59980
rect 80 59979 102 59985
rect 42 59946 46 59976
rect 72 59946 76 59976
rect 42 59865 46 59899
rect 72 59865 76 59899
rect -25 59828 25 59830
rect -8 59820 14 59827
rect -8 59819 17 59820
rect 25 59819 27 59828
rect -12 59812 38 59819
rect -12 59811 34 59812
rect -12 59807 8 59811
rect 0 59795 8 59807
rect 14 59795 34 59811
rect 0 59794 34 59795
rect 0 59787 38 59794
rect 14 59786 17 59787
rect 25 59778 27 59787
rect 42 59758 45 59848
rect 69 59833 80 59865
rect 107 59833 143 59861
rect 144 59833 148 60053
rect 332 59985 336 60053
rect 380 60023 462 60055
rect 463 60023 472 60057
rect 480 60023 497 60057
rect 378 60015 464 60023
rect 505 60015 507 60065
rect 514 60023 548 60057
rect 565 60023 582 60057
rect 607 60015 609 60065
rect 404 59999 438 60015
rect 400 59985 442 59986
rect 378 59979 404 59985
rect 442 59979 464 59985
rect 400 59978 404 59979
rect 174 59939 246 59947
rect 295 59944 300 59978
rect 324 59944 329 59978
rect 224 59909 226 59925
rect 196 59901 226 59909
rect 332 59907 336 59975
rect 367 59944 438 59978
rect 400 59937 404 59944
rect 454 59931 504 59933
rect 494 59927 548 59931
rect 494 59922 514 59927
rect 504 59907 506 59922
rect 196 59897 232 59901
rect 196 59867 204 59897
rect 216 59867 232 59897
rect 400 59899 404 59907
rect 107 59827 119 59833
rect 109 59799 119 59827
rect 129 59799 149 59833
rect 174 59829 181 59859
rect 224 59820 226 59867
rect 256 59859 328 59867
rect 332 59865 336 59895
rect 400 59865 408 59899
rect 434 59865 438 59899
rect 498 59897 506 59907
rect 514 59897 515 59917
rect 504 59881 506 59897
rect 525 59888 528 59922
rect 547 59897 548 59917
rect 557 59897 564 59907
rect 514 59881 530 59887
rect 532 59881 548 59887
rect 278 59829 305 59840
rect 42 59707 46 59741
rect 72 59707 76 59741
rect 38 59669 80 59670
rect 42 59628 76 59662
rect 79 59628 113 59662
rect 42 59549 46 59583
rect 72 59549 76 59583
rect -25 59512 25 59514
rect -8 59504 14 59511
rect -8 59503 17 59504
rect 25 59503 27 59512
rect -12 59496 38 59503
rect -12 59495 34 59496
rect -12 59491 8 59495
rect 0 59479 8 59491
rect 14 59479 34 59495
rect 0 59478 34 59479
rect 0 59471 38 59478
rect 14 59470 17 59471
rect 25 59462 27 59471
rect 42 59442 45 59532
rect 71 59501 80 59529
rect 69 59463 80 59501
rect 144 59491 148 59799
rect 196 59786 204 59820
rect 216 59786 232 59820
rect 244 59816 257 59820
rect 300 59816 308 59829
rect 332 59827 342 59865
rect 400 59857 404 59865
rect 336 59817 342 59827
rect 244 59792 291 59816
rect 244 59786 257 59792
rect 224 59739 226 59786
rect 278 59782 291 59792
rect 300 59792 329 59816
rect 332 59807 342 59817
rect 400 59817 409 59845
rect 562 59828 612 59830
rect 466 59819 497 59827
rect 565 59819 596 59827
rect 300 59782 321 59792
rect 300 59776 308 59782
rect 289 59766 308 59776
rect 196 59709 204 59739
rect 216 59709 232 59739
rect 196 59705 232 59709
rect 196 59697 226 59705
rect 300 59697 308 59766
rect 332 59773 351 59807
rect 361 59779 381 59807
rect 361 59773 375 59779
rect 400 59773 411 59817
rect 442 59812 500 59819
rect 466 59811 500 59812
rect 565 59811 599 59819
rect 497 59795 500 59811
rect 596 59795 599 59811
rect 466 59794 500 59795
rect 442 59787 500 59794
rect 565 59787 599 59795
rect 612 59778 614 59828
rect 332 59749 342 59773
rect 336 59737 342 59749
rect 224 59681 226 59697
rect 332 59669 342 59737
rect 400 59741 404 59749
rect 400 59707 408 59741
rect 434 59707 438 59741
rect 454 59725 504 59727
rect 504 59709 506 59725
rect 514 59719 530 59725
rect 532 59719 548 59725
rect 525 59709 548 59718
rect 400 59699 404 59707
rect 498 59699 506 59709
rect 504 59675 506 59699
rect 514 59689 515 59709
rect 525 59684 528 59709
rect 547 59689 548 59709
rect 557 59699 564 59709
rect 514 59675 548 59679
rect 151 59628 156 59662
rect 174 59659 246 59667
rect 256 59659 328 59667
rect 336 59661 342 59669
rect 400 59664 404 59669
rect 180 59631 185 59659
rect 174 59623 246 59631
rect 256 59623 328 59631
rect 332 59629 336 59659
rect 400 59630 438 59664
rect 224 59593 226 59609
rect 196 59585 226 59593
rect 196 59581 232 59585
rect 196 59551 204 59581
rect 216 59551 232 59581
rect 224 59504 226 59551
rect 300 59524 308 59593
rect 332 59591 342 59629
rect 400 59621 404 59630
rect 454 59615 504 59617
rect 494 59611 548 59615
rect 494 59606 514 59611
rect 504 59591 506 59606
rect 336 59579 342 59591
rect 289 59514 308 59524
rect 300 59508 308 59514
rect 332 59545 342 59579
rect 400 59583 404 59591
rect 400 59549 408 59583
rect 434 59549 438 59583
rect 498 59581 506 59591
rect 514 59581 515 59601
rect 504 59565 506 59581
rect 525 59572 528 59606
rect 547 59581 548 59601
rect 557 59581 564 59591
rect 514 59565 530 59571
rect 532 59565 548 59571
rect 332 59517 373 59545
rect 332 59511 351 59517
rect 107 59457 119 59491
rect 129 59457 149 59491
rect 196 59470 204 59504
rect 216 59470 232 59504
rect 244 59498 257 59504
rect 278 59498 291 59508
rect 244 59474 291 59498
rect 300 59498 321 59508
rect 336 59501 351 59511
rect 300 59474 329 59498
rect 332 59483 351 59501
rect 361 59511 375 59517
rect 400 59511 411 59549
rect 562 59512 612 59514
rect 361 59483 381 59511
rect 400 59483 409 59511
rect 466 59503 497 59511
rect 565 59503 596 59511
rect 442 59496 500 59503
rect 466 59495 500 59496
rect 565 59495 599 59503
rect 244 59470 257 59474
rect 42 59391 46 59425
rect 72 59391 76 59425
rect 42 59344 76 59348
rect 42 59329 46 59344
rect 72 59329 76 59344
rect 38 59311 80 59329
rect 16 59305 102 59311
rect 144 59305 148 59457
rect 174 59433 181 59461
rect 224 59423 226 59470
rect 300 59461 308 59474
rect 278 59450 305 59461
rect 332 59433 342 59483
rect 400 59463 404 59483
rect 497 59479 500 59495
rect 596 59479 599 59495
rect 466 59478 500 59479
rect 442 59471 500 59478
rect 565 59471 599 59479
rect 612 59462 614 59512
rect 256 59423 328 59431
rect 336 59425 342 59433
rect 400 59425 404 59433
rect 196 59393 204 59423
rect 216 59393 232 59423
rect 196 59389 232 59393
rect 196 59381 226 59389
rect 224 59365 226 59381
rect 332 59353 336 59421
rect 400 59391 408 59425
rect 434 59391 438 59425
rect 454 59409 504 59411
rect 504 59393 506 59409
rect 514 59403 530 59409
rect 532 59403 548 59409
rect 525 59393 548 59402
rect 400 59383 404 59391
rect 498 59383 506 59393
rect 504 59359 506 59383
rect 514 59373 515 59393
rect 525 59368 528 59393
rect 547 59373 548 59393
rect 557 59383 564 59393
rect 514 59359 548 59363
rect 400 59353 442 59354
rect 174 59343 246 59351
rect 400 59346 404 59353
rect 295 59312 300 59346
rect 324 59312 329 59346
rect 367 59329 438 59346
rect 367 59312 442 59329
rect 400 59311 442 59312
rect 378 59305 464 59311
rect 38 59289 80 59305
rect 400 59289 442 59305
rect -25 59275 25 59277
rect 42 59275 76 59289
rect 404 59275 438 59289
rect 455 59275 505 59277
rect 557 59275 607 59277
rect 16 59267 102 59275
rect 378 59267 464 59275
rect 8 59233 17 59267
rect 18 59265 51 59267
rect 80 59265 100 59267
rect 18 59233 100 59265
rect 380 59265 404 59267
rect 429 59265 438 59267
rect 442 59265 462 59267
rect 16 59225 102 59233
rect 42 59209 76 59225
rect 16 59189 38 59195
rect 42 59186 76 59190
rect 80 59189 102 59195
rect 42 59156 46 59186
rect 72 59156 76 59186
rect 42 59075 46 59109
rect 72 59075 76 59109
rect -25 59038 25 59040
rect -8 59030 14 59037
rect -8 59029 17 59030
rect 25 59029 27 59038
rect -12 59022 38 59029
rect -12 59021 34 59022
rect -12 59017 8 59021
rect 0 59005 8 59017
rect 14 59005 34 59021
rect 0 59004 34 59005
rect 0 58997 38 59004
rect 14 58996 17 58997
rect 25 58988 27 58997
rect 42 58968 45 59058
rect 69 59043 80 59075
rect 107 59043 143 59071
rect 144 59043 148 59263
rect 332 59195 336 59263
rect 380 59233 462 59265
rect 463 59233 472 59267
rect 480 59233 497 59267
rect 378 59225 464 59233
rect 505 59225 507 59275
rect 514 59233 548 59267
rect 565 59233 582 59267
rect 607 59225 609 59275
rect 404 59209 438 59225
rect 400 59195 442 59196
rect 378 59189 404 59195
rect 442 59189 464 59195
rect 400 59188 404 59189
rect 174 59149 246 59157
rect 295 59154 300 59188
rect 324 59154 329 59188
rect 224 59119 226 59135
rect 196 59111 226 59119
rect 332 59117 336 59185
rect 367 59154 438 59188
rect 400 59147 404 59154
rect 454 59141 504 59143
rect 494 59137 548 59141
rect 494 59132 514 59137
rect 504 59117 506 59132
rect 196 59107 232 59111
rect 196 59077 204 59107
rect 216 59077 232 59107
rect 400 59109 404 59117
rect 107 59037 119 59043
rect 109 59009 119 59037
rect 129 59009 149 59043
rect 174 59039 181 59069
rect 224 59030 226 59077
rect 256 59069 328 59077
rect 332 59075 336 59105
rect 400 59075 408 59109
rect 434 59075 438 59109
rect 498 59107 506 59117
rect 514 59107 515 59127
rect 504 59091 506 59107
rect 525 59098 528 59132
rect 547 59107 548 59127
rect 557 59107 564 59117
rect 514 59091 530 59097
rect 532 59091 548 59097
rect 278 59039 305 59050
rect 42 58917 46 58951
rect 72 58917 76 58951
rect 38 58879 80 58880
rect 42 58838 76 58872
rect 79 58838 113 58872
rect 42 58759 46 58793
rect 72 58759 76 58793
rect -25 58722 25 58724
rect -8 58714 14 58721
rect -8 58713 17 58714
rect 25 58713 27 58722
rect -12 58706 38 58713
rect -12 58705 34 58706
rect -12 58701 8 58705
rect 0 58689 8 58701
rect 14 58689 34 58705
rect 0 58688 34 58689
rect 0 58681 38 58688
rect 14 58680 17 58681
rect 25 58672 27 58681
rect 42 58652 45 58742
rect 71 58711 80 58739
rect 69 58673 80 58711
rect 144 58701 148 59009
rect 196 58996 204 59030
rect 216 58996 232 59030
rect 244 59026 257 59030
rect 300 59026 308 59039
rect 332 59037 342 59075
rect 400 59067 404 59075
rect 336 59027 342 59037
rect 244 59002 291 59026
rect 244 58996 257 59002
rect 224 58949 226 58996
rect 278 58992 291 59002
rect 300 59002 329 59026
rect 332 59017 342 59027
rect 400 59027 409 59055
rect 562 59038 612 59040
rect 466 59029 497 59037
rect 565 59029 596 59037
rect 300 58992 321 59002
rect 300 58986 308 58992
rect 289 58976 308 58986
rect 196 58919 204 58949
rect 216 58919 232 58949
rect 196 58915 232 58919
rect 196 58907 226 58915
rect 300 58907 308 58976
rect 332 58983 351 59017
rect 361 58989 381 59017
rect 361 58983 375 58989
rect 400 58983 411 59027
rect 442 59022 500 59029
rect 466 59021 500 59022
rect 565 59021 599 59029
rect 497 59005 500 59021
rect 596 59005 599 59021
rect 466 59004 500 59005
rect 442 58997 500 59004
rect 565 58997 599 59005
rect 612 58988 614 59038
rect 332 58959 342 58983
rect 336 58947 342 58959
rect 224 58891 226 58907
rect 332 58879 342 58947
rect 400 58951 404 58959
rect 400 58917 408 58951
rect 434 58917 438 58951
rect 454 58935 504 58937
rect 504 58919 506 58935
rect 514 58929 530 58935
rect 532 58929 548 58935
rect 525 58919 548 58928
rect 400 58909 404 58917
rect 498 58909 506 58919
rect 504 58885 506 58909
rect 514 58899 515 58919
rect 525 58894 528 58919
rect 547 58899 548 58919
rect 557 58909 564 58919
rect 514 58885 548 58889
rect 151 58838 156 58872
rect 174 58869 246 58877
rect 256 58869 328 58877
rect 336 58871 342 58879
rect 400 58874 404 58879
rect 180 58841 185 58869
rect 174 58833 246 58841
rect 256 58833 328 58841
rect 332 58839 336 58869
rect 400 58840 438 58874
rect 224 58803 226 58819
rect 196 58795 226 58803
rect 196 58791 232 58795
rect 196 58761 204 58791
rect 216 58761 232 58791
rect 224 58714 226 58761
rect 300 58734 308 58803
rect 332 58801 342 58839
rect 400 58831 404 58840
rect 454 58825 504 58827
rect 494 58821 548 58825
rect 494 58816 514 58821
rect 504 58801 506 58816
rect 336 58789 342 58801
rect 289 58724 308 58734
rect 300 58718 308 58724
rect 332 58755 342 58789
rect 400 58793 404 58801
rect 400 58759 408 58793
rect 434 58759 438 58793
rect 498 58791 506 58801
rect 514 58791 515 58811
rect 504 58775 506 58791
rect 525 58782 528 58816
rect 547 58791 548 58811
rect 557 58791 564 58801
rect 514 58775 530 58781
rect 532 58775 548 58781
rect 332 58727 373 58755
rect 332 58721 351 58727
rect 107 58667 119 58701
rect 129 58667 149 58701
rect 196 58680 204 58714
rect 216 58680 232 58714
rect 244 58708 257 58714
rect 278 58708 291 58718
rect 244 58684 291 58708
rect 300 58708 321 58718
rect 336 58711 351 58721
rect 300 58684 329 58708
rect 332 58693 351 58711
rect 361 58721 375 58727
rect 400 58721 411 58759
rect 562 58722 612 58724
rect 361 58693 381 58721
rect 400 58693 409 58721
rect 466 58713 497 58721
rect 565 58713 596 58721
rect 442 58706 500 58713
rect 466 58705 500 58706
rect 565 58705 599 58713
rect 244 58680 257 58684
rect 42 58601 46 58635
rect 72 58601 76 58635
rect 42 58554 76 58558
rect 42 58539 46 58554
rect 72 58539 76 58554
rect 38 58521 80 58539
rect 16 58515 102 58521
rect 144 58515 148 58667
rect 174 58643 181 58671
rect 224 58633 226 58680
rect 300 58671 308 58684
rect 278 58660 305 58671
rect 332 58643 342 58693
rect 400 58673 404 58693
rect 497 58689 500 58705
rect 596 58689 599 58705
rect 466 58688 500 58689
rect 442 58681 500 58688
rect 565 58681 599 58689
rect 612 58672 614 58722
rect 256 58633 328 58641
rect 336 58635 342 58643
rect 400 58635 404 58643
rect 196 58603 204 58633
rect 216 58603 232 58633
rect 196 58599 232 58603
rect 196 58591 226 58599
rect 224 58575 226 58591
rect 332 58563 336 58631
rect 400 58601 408 58635
rect 434 58601 438 58635
rect 454 58619 504 58621
rect 504 58603 506 58619
rect 514 58613 530 58619
rect 532 58613 548 58619
rect 525 58603 548 58612
rect 400 58593 404 58601
rect 498 58593 506 58603
rect 504 58569 506 58593
rect 514 58583 515 58603
rect 525 58578 528 58603
rect 547 58583 548 58603
rect 557 58593 564 58603
rect 514 58569 548 58573
rect 400 58563 442 58564
rect 174 58553 246 58561
rect 400 58556 404 58563
rect 295 58522 300 58556
rect 324 58522 329 58556
rect 367 58539 438 58556
rect 367 58522 442 58539
rect 400 58521 442 58522
rect 378 58515 464 58521
rect 38 58499 80 58515
rect 400 58499 442 58515
rect -25 58485 25 58487
rect 42 58485 76 58499
rect 404 58485 438 58499
rect 455 58485 505 58487
rect 557 58485 607 58487
rect 16 58477 102 58485
rect 378 58477 464 58485
rect 8 58443 17 58477
rect 18 58475 51 58477
rect 80 58475 100 58477
rect 18 58443 100 58475
rect 380 58475 404 58477
rect 429 58475 438 58477
rect 442 58475 462 58477
rect 16 58435 102 58443
rect 42 58419 76 58435
rect 16 58399 38 58405
rect 42 58396 76 58400
rect 80 58399 102 58405
rect 42 58366 46 58396
rect 72 58366 76 58396
rect 42 58285 46 58319
rect 72 58285 76 58319
rect -25 58248 25 58250
rect -8 58240 14 58247
rect -8 58239 17 58240
rect 25 58239 27 58248
rect -12 58232 38 58239
rect -12 58231 34 58232
rect -12 58227 8 58231
rect 0 58215 8 58227
rect 14 58215 34 58231
rect 0 58214 34 58215
rect 0 58207 38 58214
rect 14 58206 17 58207
rect 25 58198 27 58207
rect 42 58178 45 58268
rect 69 58253 80 58285
rect 107 58253 143 58281
rect 144 58253 148 58473
rect 332 58405 336 58473
rect 380 58443 462 58475
rect 463 58443 472 58477
rect 480 58443 497 58477
rect 378 58435 464 58443
rect 505 58435 507 58485
rect 514 58443 548 58477
rect 565 58443 582 58477
rect 607 58435 609 58485
rect 404 58419 438 58435
rect 400 58405 442 58406
rect 378 58399 404 58405
rect 442 58399 464 58405
rect 400 58398 404 58399
rect 174 58359 246 58367
rect 295 58364 300 58398
rect 324 58364 329 58398
rect 224 58329 226 58345
rect 196 58321 226 58329
rect 332 58327 336 58395
rect 367 58364 438 58398
rect 400 58357 404 58364
rect 454 58351 504 58353
rect 494 58347 548 58351
rect 494 58342 514 58347
rect 504 58327 506 58342
rect 196 58317 232 58321
rect 196 58287 204 58317
rect 216 58287 232 58317
rect 400 58319 404 58327
rect 107 58247 119 58253
rect 109 58219 119 58247
rect 129 58219 149 58253
rect 174 58249 181 58279
rect 224 58240 226 58287
rect 256 58279 328 58287
rect 332 58285 336 58315
rect 400 58285 408 58319
rect 434 58285 438 58319
rect 498 58317 506 58327
rect 514 58317 515 58337
rect 504 58301 506 58317
rect 525 58308 528 58342
rect 547 58317 548 58337
rect 557 58317 564 58327
rect 514 58301 530 58307
rect 532 58301 548 58307
rect 278 58249 305 58260
rect 42 58127 46 58161
rect 72 58127 76 58161
rect 38 58089 80 58090
rect 42 58048 76 58082
rect 79 58048 113 58082
rect 42 57969 46 58003
rect 72 57969 76 58003
rect -25 57932 25 57934
rect -8 57924 14 57931
rect -8 57923 17 57924
rect 25 57923 27 57932
rect -12 57916 38 57923
rect -12 57915 34 57916
rect -12 57911 8 57915
rect 0 57899 8 57911
rect 14 57899 34 57915
rect 0 57898 34 57899
rect 0 57891 38 57898
rect 14 57890 17 57891
rect 25 57882 27 57891
rect 42 57862 45 57952
rect 71 57921 80 57949
rect 69 57883 80 57921
rect 144 57911 148 58219
rect 196 58206 204 58240
rect 216 58206 232 58240
rect 244 58236 257 58240
rect 300 58236 308 58249
rect 332 58247 342 58285
rect 400 58277 404 58285
rect 336 58237 342 58247
rect 244 58212 291 58236
rect 244 58206 257 58212
rect 224 58159 226 58206
rect 278 58202 291 58212
rect 300 58212 329 58236
rect 332 58227 342 58237
rect 400 58237 409 58265
rect 562 58248 612 58250
rect 466 58239 497 58247
rect 565 58239 596 58247
rect 300 58202 321 58212
rect 300 58196 308 58202
rect 289 58186 308 58196
rect 196 58129 204 58159
rect 216 58129 232 58159
rect 196 58125 232 58129
rect 196 58117 226 58125
rect 300 58117 308 58186
rect 332 58193 351 58227
rect 361 58199 381 58227
rect 361 58193 375 58199
rect 400 58193 411 58237
rect 442 58232 500 58239
rect 466 58231 500 58232
rect 565 58231 599 58239
rect 497 58215 500 58231
rect 596 58215 599 58231
rect 466 58214 500 58215
rect 442 58207 500 58214
rect 565 58207 599 58215
rect 612 58198 614 58248
rect 332 58169 342 58193
rect 336 58157 342 58169
rect 224 58101 226 58117
rect 332 58089 342 58157
rect 400 58161 404 58169
rect 400 58127 408 58161
rect 434 58127 438 58161
rect 454 58145 504 58147
rect 504 58129 506 58145
rect 514 58139 530 58145
rect 532 58139 548 58145
rect 525 58129 548 58138
rect 400 58119 404 58127
rect 498 58119 506 58129
rect 504 58095 506 58119
rect 514 58109 515 58129
rect 525 58104 528 58129
rect 547 58109 548 58129
rect 557 58119 564 58129
rect 514 58095 548 58099
rect 151 58048 156 58082
rect 174 58079 246 58087
rect 256 58079 328 58087
rect 336 58081 342 58089
rect 400 58084 404 58089
rect 180 58051 185 58079
rect 174 58043 246 58051
rect 256 58043 328 58051
rect 332 58049 336 58079
rect 400 58050 438 58084
rect 224 58013 226 58029
rect 196 58005 226 58013
rect 196 58001 232 58005
rect 196 57971 204 58001
rect 216 57971 232 58001
rect 224 57924 226 57971
rect 300 57944 308 58013
rect 332 58011 342 58049
rect 400 58041 404 58050
rect 454 58035 504 58037
rect 494 58031 548 58035
rect 494 58026 514 58031
rect 504 58011 506 58026
rect 336 57999 342 58011
rect 289 57934 308 57944
rect 300 57928 308 57934
rect 332 57965 342 57999
rect 400 58003 404 58011
rect 400 57969 408 58003
rect 434 57969 438 58003
rect 498 58001 506 58011
rect 514 58001 515 58021
rect 504 57985 506 58001
rect 525 57992 528 58026
rect 547 58001 548 58021
rect 557 58001 564 58011
rect 514 57985 530 57991
rect 532 57985 548 57991
rect 332 57937 373 57965
rect 332 57931 351 57937
rect 107 57877 119 57911
rect 129 57877 149 57911
rect 196 57890 204 57924
rect 216 57890 232 57924
rect 244 57918 257 57924
rect 278 57918 291 57928
rect 244 57894 291 57918
rect 300 57918 321 57928
rect 336 57921 351 57931
rect 300 57894 329 57918
rect 332 57903 351 57921
rect 361 57931 375 57937
rect 400 57931 411 57969
rect 562 57932 612 57934
rect 361 57903 381 57931
rect 400 57903 409 57931
rect 466 57923 497 57931
rect 565 57923 596 57931
rect 442 57916 500 57923
rect 466 57915 500 57916
rect 565 57915 599 57923
rect 244 57890 257 57894
rect 42 57811 46 57845
rect 72 57811 76 57845
rect 42 57764 76 57768
rect 42 57749 46 57764
rect 72 57749 76 57764
rect 38 57731 80 57749
rect 16 57725 102 57731
rect 144 57725 148 57877
rect 174 57853 181 57881
rect 224 57843 226 57890
rect 300 57881 308 57894
rect 278 57870 305 57881
rect 332 57853 342 57903
rect 400 57883 404 57903
rect 497 57899 500 57915
rect 596 57899 599 57915
rect 466 57898 500 57899
rect 442 57891 500 57898
rect 565 57891 599 57899
rect 612 57882 614 57932
rect 256 57843 328 57851
rect 336 57845 342 57853
rect 400 57845 404 57853
rect 196 57813 204 57843
rect 216 57813 232 57843
rect 196 57809 232 57813
rect 196 57801 226 57809
rect 224 57785 226 57801
rect 332 57773 336 57841
rect 400 57811 408 57845
rect 434 57811 438 57845
rect 454 57829 504 57831
rect 504 57813 506 57829
rect 514 57823 530 57829
rect 532 57823 548 57829
rect 525 57813 548 57822
rect 400 57803 404 57811
rect 498 57803 506 57813
rect 504 57779 506 57803
rect 514 57793 515 57813
rect 525 57788 528 57813
rect 547 57793 548 57813
rect 557 57803 564 57813
rect 514 57779 548 57783
rect 400 57773 442 57774
rect 174 57763 246 57771
rect 400 57766 404 57773
rect 295 57732 300 57766
rect 324 57732 329 57766
rect 367 57749 438 57766
rect 367 57732 442 57749
rect 400 57731 442 57732
rect 378 57725 464 57731
rect 38 57709 80 57725
rect 400 57709 442 57725
rect -25 57695 25 57697
rect 42 57695 76 57709
rect 404 57695 438 57709
rect 455 57695 505 57697
rect 557 57695 607 57697
rect 16 57687 102 57695
rect 378 57687 464 57695
rect 8 57653 17 57687
rect 18 57685 51 57687
rect 80 57685 100 57687
rect 18 57653 100 57685
rect 380 57685 404 57687
rect 429 57685 438 57687
rect 442 57685 462 57687
rect 16 57645 102 57653
rect 42 57629 76 57645
rect 16 57609 38 57615
rect 42 57606 76 57610
rect 80 57609 102 57615
rect 42 57576 46 57606
rect 72 57576 76 57606
rect 42 57495 46 57529
rect 72 57495 76 57529
rect -25 57458 25 57460
rect -8 57450 14 57457
rect -8 57449 17 57450
rect 25 57449 27 57458
rect -12 57442 38 57449
rect -12 57441 34 57442
rect -12 57437 8 57441
rect 0 57425 8 57437
rect 14 57425 34 57441
rect 0 57424 34 57425
rect 0 57417 38 57424
rect 14 57416 17 57417
rect 25 57408 27 57417
rect 42 57388 45 57478
rect 69 57463 80 57495
rect 107 57463 143 57491
rect 144 57463 148 57683
rect 332 57615 336 57683
rect 380 57653 462 57685
rect 463 57653 472 57687
rect 480 57653 497 57687
rect 378 57645 464 57653
rect 505 57645 507 57695
rect 514 57653 548 57687
rect 565 57653 582 57687
rect 607 57645 609 57695
rect 404 57629 438 57645
rect 400 57615 442 57616
rect 378 57609 404 57615
rect 442 57609 464 57615
rect 400 57608 404 57609
rect 174 57569 246 57577
rect 295 57574 300 57608
rect 324 57574 329 57608
rect 224 57539 226 57555
rect 196 57531 226 57539
rect 332 57537 336 57605
rect 367 57574 438 57608
rect 400 57567 404 57574
rect 454 57561 504 57563
rect 494 57557 548 57561
rect 494 57552 514 57557
rect 504 57537 506 57552
rect 196 57527 232 57531
rect 196 57497 204 57527
rect 216 57497 232 57527
rect 400 57529 404 57537
rect 107 57457 119 57463
rect 109 57429 119 57457
rect 129 57429 149 57463
rect 174 57459 181 57489
rect 224 57450 226 57497
rect 256 57489 328 57497
rect 332 57495 336 57525
rect 400 57495 408 57529
rect 434 57495 438 57529
rect 498 57527 506 57537
rect 514 57527 515 57547
rect 504 57511 506 57527
rect 525 57518 528 57552
rect 547 57527 548 57547
rect 557 57527 564 57537
rect 514 57511 530 57517
rect 532 57511 548 57517
rect 278 57459 305 57470
rect 42 57337 46 57371
rect 72 57337 76 57371
rect 38 57299 80 57300
rect 42 57258 76 57292
rect 79 57258 113 57292
rect 42 57179 46 57213
rect 72 57179 76 57213
rect -25 57142 25 57144
rect -8 57134 14 57141
rect -8 57133 17 57134
rect 25 57133 27 57142
rect -12 57126 38 57133
rect -12 57125 34 57126
rect -12 57121 8 57125
rect 0 57109 8 57121
rect 14 57109 34 57125
rect 0 57108 34 57109
rect 0 57101 38 57108
rect 14 57100 17 57101
rect 25 57092 27 57101
rect 42 57072 45 57162
rect 71 57131 80 57159
rect 69 57093 80 57131
rect 144 57121 148 57429
rect 196 57416 204 57450
rect 216 57416 232 57450
rect 244 57446 257 57450
rect 300 57446 308 57459
rect 332 57457 342 57495
rect 400 57487 404 57495
rect 336 57447 342 57457
rect 244 57422 291 57446
rect 244 57416 257 57422
rect 224 57369 226 57416
rect 278 57412 291 57422
rect 300 57422 329 57446
rect 332 57437 342 57447
rect 400 57447 409 57475
rect 562 57458 612 57460
rect 466 57449 497 57457
rect 565 57449 596 57457
rect 300 57412 321 57422
rect 300 57406 308 57412
rect 289 57396 308 57406
rect 196 57339 204 57369
rect 216 57339 232 57369
rect 196 57335 232 57339
rect 196 57327 226 57335
rect 300 57327 308 57396
rect 332 57403 351 57437
rect 361 57409 381 57437
rect 361 57403 375 57409
rect 400 57403 411 57447
rect 442 57442 500 57449
rect 466 57441 500 57442
rect 565 57441 599 57449
rect 497 57425 500 57441
rect 596 57425 599 57441
rect 466 57424 500 57425
rect 442 57417 500 57424
rect 565 57417 599 57425
rect 612 57408 614 57458
rect 332 57379 342 57403
rect 336 57367 342 57379
rect 224 57311 226 57327
rect 332 57299 342 57367
rect 400 57371 404 57379
rect 400 57337 408 57371
rect 434 57337 438 57371
rect 454 57355 504 57357
rect 504 57339 506 57355
rect 514 57349 530 57355
rect 532 57349 548 57355
rect 525 57339 548 57348
rect 400 57329 404 57337
rect 498 57329 506 57339
rect 504 57305 506 57329
rect 514 57319 515 57339
rect 525 57314 528 57339
rect 547 57319 548 57339
rect 557 57329 564 57339
rect 514 57305 548 57309
rect 151 57258 156 57292
rect 174 57289 246 57297
rect 256 57289 328 57297
rect 336 57291 342 57299
rect 400 57294 404 57299
rect 180 57261 185 57289
rect 174 57253 246 57261
rect 256 57253 328 57261
rect 332 57259 336 57289
rect 400 57260 438 57294
rect 224 57223 226 57239
rect 196 57215 226 57223
rect 196 57211 232 57215
rect 196 57181 204 57211
rect 216 57181 232 57211
rect 224 57134 226 57181
rect 300 57154 308 57223
rect 332 57221 342 57259
rect 400 57251 404 57260
rect 454 57245 504 57247
rect 494 57241 548 57245
rect 494 57236 514 57241
rect 504 57221 506 57236
rect 336 57209 342 57221
rect 289 57144 308 57154
rect 300 57138 308 57144
rect 332 57175 342 57209
rect 400 57213 404 57221
rect 400 57179 408 57213
rect 434 57179 438 57213
rect 498 57211 506 57221
rect 514 57211 515 57231
rect 504 57195 506 57211
rect 525 57202 528 57236
rect 547 57211 548 57231
rect 557 57211 564 57221
rect 514 57195 530 57201
rect 532 57195 548 57201
rect 332 57147 373 57175
rect 332 57141 351 57147
rect 107 57087 119 57121
rect 129 57087 149 57121
rect 196 57100 204 57134
rect 216 57100 232 57134
rect 244 57128 257 57134
rect 278 57128 291 57138
rect 244 57104 291 57128
rect 300 57128 321 57138
rect 336 57131 351 57141
rect 300 57104 329 57128
rect 332 57113 351 57131
rect 361 57141 375 57147
rect 400 57141 411 57179
rect 562 57142 612 57144
rect 361 57113 381 57141
rect 400 57113 409 57141
rect 466 57133 497 57141
rect 565 57133 596 57141
rect 442 57126 500 57133
rect 466 57125 500 57126
rect 565 57125 599 57133
rect 244 57100 257 57104
rect 42 57021 46 57055
rect 72 57021 76 57055
rect 42 56974 76 56978
rect 42 56959 46 56974
rect 72 56959 76 56974
rect 38 56941 80 56959
rect 16 56935 102 56941
rect 144 56935 148 57087
rect 174 57063 181 57091
rect 224 57053 226 57100
rect 300 57091 308 57104
rect 278 57080 305 57091
rect 332 57063 342 57113
rect 400 57093 404 57113
rect 497 57109 500 57125
rect 596 57109 599 57125
rect 466 57108 500 57109
rect 442 57101 500 57108
rect 565 57101 599 57109
rect 612 57092 614 57142
rect 256 57053 328 57061
rect 336 57055 342 57063
rect 400 57055 404 57063
rect 196 57023 204 57053
rect 216 57023 232 57053
rect 196 57019 232 57023
rect 196 57011 226 57019
rect 224 56995 226 57011
rect 332 56983 336 57051
rect 400 57021 408 57055
rect 434 57021 438 57055
rect 454 57039 504 57041
rect 504 57023 506 57039
rect 514 57033 530 57039
rect 532 57033 548 57039
rect 525 57023 548 57032
rect 400 57013 404 57021
rect 498 57013 506 57023
rect 504 56989 506 57013
rect 514 57003 515 57023
rect 525 56998 528 57023
rect 547 57003 548 57023
rect 557 57013 564 57023
rect 514 56989 548 56993
rect 400 56983 442 56984
rect 174 56973 246 56981
rect 400 56976 404 56983
rect 295 56942 300 56976
rect 324 56942 329 56976
rect 367 56959 438 56976
rect 367 56942 442 56959
rect 400 56941 442 56942
rect 378 56935 464 56941
rect 38 56919 80 56935
rect 400 56919 442 56935
rect -25 56905 25 56907
rect 42 56905 76 56919
rect 404 56905 438 56919
rect 455 56905 505 56907
rect 557 56905 607 56907
rect 16 56897 102 56905
rect 378 56897 464 56905
rect 8 56863 17 56897
rect 18 56895 51 56897
rect 80 56895 100 56897
rect 18 56863 100 56895
rect 380 56895 404 56897
rect 429 56895 438 56897
rect 442 56895 462 56897
rect 16 56855 102 56863
rect 42 56839 76 56855
rect 16 56819 38 56825
rect 42 56816 76 56820
rect 80 56819 102 56825
rect 42 56786 46 56816
rect 72 56786 76 56816
rect 42 56705 46 56739
rect 72 56705 76 56739
rect -25 56668 25 56670
rect -8 56660 14 56667
rect -8 56659 17 56660
rect 25 56659 27 56668
rect -12 56652 38 56659
rect -12 56651 34 56652
rect -12 56647 8 56651
rect 0 56635 8 56647
rect 14 56635 34 56651
rect 0 56634 34 56635
rect 0 56627 38 56634
rect 14 56626 17 56627
rect 25 56618 27 56627
rect 42 56598 45 56688
rect 69 56673 80 56705
rect 107 56673 143 56701
rect 144 56673 148 56893
rect 332 56825 336 56893
rect 380 56863 462 56895
rect 463 56863 472 56897
rect 480 56863 497 56897
rect 378 56855 464 56863
rect 505 56855 507 56905
rect 514 56863 548 56897
rect 565 56863 582 56897
rect 607 56855 609 56905
rect 404 56839 438 56855
rect 400 56825 442 56826
rect 378 56819 404 56825
rect 442 56819 464 56825
rect 400 56818 404 56819
rect 174 56779 246 56787
rect 295 56784 300 56818
rect 324 56784 329 56818
rect 224 56749 226 56765
rect 196 56741 226 56749
rect 332 56747 336 56815
rect 367 56784 438 56818
rect 400 56777 404 56784
rect 454 56771 504 56773
rect 494 56767 548 56771
rect 494 56762 514 56767
rect 504 56747 506 56762
rect 196 56737 232 56741
rect 196 56707 204 56737
rect 216 56707 232 56737
rect 400 56739 404 56747
rect 107 56667 119 56673
rect 109 56639 119 56667
rect 129 56639 149 56673
rect 174 56669 181 56699
rect 224 56660 226 56707
rect 256 56699 328 56707
rect 332 56705 336 56735
rect 400 56705 408 56739
rect 434 56705 438 56739
rect 498 56737 506 56747
rect 514 56737 515 56757
rect 504 56721 506 56737
rect 525 56728 528 56762
rect 547 56737 548 56757
rect 557 56737 564 56747
rect 514 56721 530 56727
rect 532 56721 548 56727
rect 278 56669 305 56680
rect 42 56547 46 56581
rect 72 56547 76 56581
rect 38 56509 80 56510
rect 42 56468 76 56502
rect 79 56468 113 56502
rect 42 56389 46 56423
rect 72 56389 76 56423
rect -25 56352 25 56354
rect -8 56344 14 56351
rect -8 56343 17 56344
rect 25 56343 27 56352
rect -12 56336 38 56343
rect -12 56335 34 56336
rect -12 56331 8 56335
rect 0 56319 8 56331
rect 14 56319 34 56335
rect 0 56318 34 56319
rect 0 56311 38 56318
rect 14 56310 17 56311
rect 25 56302 27 56311
rect 42 56282 45 56372
rect 71 56341 80 56369
rect 69 56303 80 56341
rect 144 56331 148 56639
rect 196 56626 204 56660
rect 216 56626 232 56660
rect 244 56656 257 56660
rect 300 56656 308 56669
rect 332 56667 342 56705
rect 400 56697 404 56705
rect 336 56657 342 56667
rect 244 56632 291 56656
rect 244 56626 257 56632
rect 224 56579 226 56626
rect 278 56622 291 56632
rect 300 56632 329 56656
rect 332 56647 342 56657
rect 400 56657 409 56685
rect 562 56668 612 56670
rect 466 56659 497 56667
rect 565 56659 596 56667
rect 300 56622 321 56632
rect 300 56616 308 56622
rect 289 56606 308 56616
rect 196 56549 204 56579
rect 216 56549 232 56579
rect 196 56545 232 56549
rect 196 56537 226 56545
rect 300 56537 308 56606
rect 332 56613 351 56647
rect 361 56619 381 56647
rect 361 56613 375 56619
rect 400 56613 411 56657
rect 442 56652 500 56659
rect 466 56651 500 56652
rect 565 56651 599 56659
rect 497 56635 500 56651
rect 596 56635 599 56651
rect 466 56634 500 56635
rect 442 56627 500 56634
rect 565 56627 599 56635
rect 612 56618 614 56668
rect 332 56589 342 56613
rect 336 56577 342 56589
rect 224 56521 226 56537
rect 332 56509 342 56577
rect 400 56581 404 56589
rect 400 56547 408 56581
rect 434 56547 438 56581
rect 454 56565 504 56567
rect 504 56549 506 56565
rect 514 56559 530 56565
rect 532 56559 548 56565
rect 525 56549 548 56558
rect 400 56539 404 56547
rect 498 56539 506 56549
rect 504 56515 506 56539
rect 514 56529 515 56549
rect 525 56524 528 56549
rect 547 56529 548 56549
rect 557 56539 564 56549
rect 514 56515 548 56519
rect 151 56468 156 56502
rect 174 56499 246 56507
rect 256 56499 328 56507
rect 336 56501 342 56509
rect 400 56504 404 56509
rect 180 56471 185 56499
rect 174 56463 246 56471
rect 256 56463 328 56471
rect 332 56469 336 56499
rect 400 56470 438 56504
rect 224 56433 226 56449
rect 196 56425 226 56433
rect 196 56421 232 56425
rect 196 56391 204 56421
rect 216 56391 232 56421
rect 224 56344 226 56391
rect 300 56364 308 56433
rect 332 56431 342 56469
rect 400 56461 404 56470
rect 454 56455 504 56457
rect 494 56451 548 56455
rect 494 56446 514 56451
rect 504 56431 506 56446
rect 336 56419 342 56431
rect 289 56354 308 56364
rect 300 56348 308 56354
rect 332 56385 342 56419
rect 400 56423 404 56431
rect 400 56389 408 56423
rect 434 56389 438 56423
rect 498 56421 506 56431
rect 514 56421 515 56441
rect 504 56405 506 56421
rect 525 56412 528 56446
rect 547 56421 548 56441
rect 557 56421 564 56431
rect 514 56405 530 56411
rect 532 56405 548 56411
rect 332 56357 373 56385
rect 332 56351 351 56357
rect 107 56297 119 56331
rect 129 56297 149 56331
rect 196 56310 204 56344
rect 216 56310 232 56344
rect 244 56338 257 56344
rect 278 56338 291 56348
rect 244 56314 291 56338
rect 300 56338 321 56348
rect 336 56341 351 56351
rect 300 56314 329 56338
rect 332 56323 351 56341
rect 361 56351 375 56357
rect 400 56351 411 56389
rect 562 56352 612 56354
rect 361 56323 381 56351
rect 400 56323 409 56351
rect 466 56343 497 56351
rect 565 56343 596 56351
rect 442 56336 500 56343
rect 466 56335 500 56336
rect 565 56335 599 56343
rect 244 56310 257 56314
rect 42 56231 46 56265
rect 72 56231 76 56265
rect 42 56184 76 56188
rect 42 56169 46 56184
rect 72 56169 76 56184
rect 38 56151 80 56169
rect 16 56145 102 56151
rect 144 56145 148 56297
rect 174 56273 181 56301
rect 224 56263 226 56310
rect 300 56301 308 56314
rect 278 56290 305 56301
rect 332 56273 342 56323
rect 400 56303 404 56323
rect 497 56319 500 56335
rect 596 56319 599 56335
rect 466 56318 500 56319
rect 442 56311 500 56318
rect 565 56311 599 56319
rect 612 56302 614 56352
rect 256 56263 328 56271
rect 336 56265 342 56273
rect 400 56265 404 56273
rect 196 56233 204 56263
rect 216 56233 232 56263
rect 196 56229 232 56233
rect 196 56221 226 56229
rect 224 56205 226 56221
rect 332 56193 336 56261
rect 400 56231 408 56265
rect 434 56231 438 56265
rect 454 56249 504 56251
rect 504 56233 506 56249
rect 514 56243 530 56249
rect 532 56243 548 56249
rect 525 56233 548 56242
rect 400 56223 404 56231
rect 498 56223 506 56233
rect 504 56199 506 56223
rect 514 56213 515 56233
rect 525 56208 528 56233
rect 547 56213 548 56233
rect 557 56223 564 56233
rect 514 56199 548 56203
rect 400 56193 442 56194
rect 174 56183 246 56191
rect 400 56186 404 56193
rect 295 56152 300 56186
rect 324 56152 329 56186
rect 367 56169 438 56186
rect 367 56152 442 56169
rect 400 56151 442 56152
rect 378 56145 464 56151
rect 38 56129 80 56145
rect 400 56129 442 56145
rect -25 56115 25 56117
rect 42 56115 76 56129
rect 404 56115 438 56129
rect 455 56115 505 56117
rect 557 56115 607 56117
rect 16 56107 102 56115
rect 378 56107 464 56115
rect 8 56073 17 56107
rect 18 56105 51 56107
rect 80 56105 100 56107
rect 18 56073 100 56105
rect 380 56105 404 56107
rect 429 56105 438 56107
rect 442 56105 462 56107
rect 16 56065 102 56073
rect 42 56049 76 56065
rect 16 56029 38 56035
rect 42 56026 76 56030
rect 80 56029 102 56035
rect 42 55996 46 56026
rect 72 55996 76 56026
rect 42 55915 46 55949
rect 72 55915 76 55949
rect -25 55878 25 55880
rect -8 55870 14 55877
rect -8 55869 17 55870
rect 25 55869 27 55878
rect -12 55862 38 55869
rect -12 55861 34 55862
rect -12 55857 8 55861
rect 0 55845 8 55857
rect 14 55845 34 55861
rect 0 55844 34 55845
rect 0 55837 38 55844
rect 14 55836 17 55837
rect 25 55828 27 55837
rect 42 55808 45 55898
rect 69 55883 80 55915
rect 107 55883 143 55911
rect 144 55883 148 56103
rect 332 56035 336 56103
rect 380 56073 462 56105
rect 463 56073 472 56107
rect 480 56073 497 56107
rect 378 56065 464 56073
rect 505 56065 507 56115
rect 514 56073 548 56107
rect 565 56073 582 56107
rect 607 56065 609 56115
rect 404 56049 438 56065
rect 400 56035 442 56036
rect 378 56029 404 56035
rect 442 56029 464 56035
rect 400 56028 404 56029
rect 174 55989 246 55997
rect 295 55994 300 56028
rect 324 55994 329 56028
rect 224 55959 226 55975
rect 196 55951 226 55959
rect 332 55957 336 56025
rect 367 55994 438 56028
rect 400 55987 404 55994
rect 454 55981 504 55983
rect 494 55977 548 55981
rect 494 55972 514 55977
rect 504 55957 506 55972
rect 196 55947 232 55951
rect 196 55917 204 55947
rect 216 55917 232 55947
rect 400 55949 404 55957
rect 107 55877 119 55883
rect 109 55849 119 55877
rect 129 55849 149 55883
rect 174 55879 181 55909
rect 224 55870 226 55917
rect 256 55909 328 55917
rect 332 55915 336 55945
rect 400 55915 408 55949
rect 434 55915 438 55949
rect 498 55947 506 55957
rect 514 55947 515 55967
rect 504 55931 506 55947
rect 525 55938 528 55972
rect 547 55947 548 55967
rect 557 55947 564 55957
rect 514 55931 530 55937
rect 532 55931 548 55937
rect 278 55879 305 55890
rect 42 55757 46 55791
rect 72 55757 76 55791
rect 38 55719 80 55720
rect 42 55678 76 55712
rect 79 55678 113 55712
rect 42 55599 46 55633
rect 72 55599 76 55633
rect -25 55562 25 55564
rect -8 55554 14 55561
rect -8 55553 17 55554
rect 25 55553 27 55562
rect -12 55546 38 55553
rect -12 55545 34 55546
rect -12 55541 8 55545
rect 0 55529 8 55541
rect 14 55529 34 55545
rect 0 55528 34 55529
rect 0 55521 38 55528
rect 14 55520 17 55521
rect 25 55512 27 55521
rect 42 55492 45 55582
rect 71 55551 80 55579
rect 69 55513 80 55551
rect 144 55541 148 55849
rect 196 55836 204 55870
rect 216 55836 232 55870
rect 244 55866 257 55870
rect 300 55866 308 55879
rect 332 55877 342 55915
rect 400 55907 404 55915
rect 336 55867 342 55877
rect 244 55842 291 55866
rect 244 55836 257 55842
rect 224 55789 226 55836
rect 278 55832 291 55842
rect 300 55842 329 55866
rect 332 55857 342 55867
rect 400 55867 409 55895
rect 562 55878 612 55880
rect 466 55869 497 55877
rect 565 55869 596 55877
rect 300 55832 321 55842
rect 300 55826 308 55832
rect 289 55816 308 55826
rect 196 55759 204 55789
rect 216 55759 232 55789
rect 196 55755 232 55759
rect 196 55747 226 55755
rect 300 55747 308 55816
rect 332 55823 351 55857
rect 361 55829 381 55857
rect 361 55823 375 55829
rect 400 55823 411 55867
rect 442 55862 500 55869
rect 466 55861 500 55862
rect 565 55861 599 55869
rect 497 55845 500 55861
rect 596 55845 599 55861
rect 466 55844 500 55845
rect 442 55837 500 55844
rect 565 55837 599 55845
rect 612 55828 614 55878
rect 332 55799 342 55823
rect 336 55787 342 55799
rect 224 55731 226 55747
rect 332 55719 342 55787
rect 400 55791 404 55799
rect 400 55757 408 55791
rect 434 55757 438 55791
rect 454 55775 504 55777
rect 504 55759 506 55775
rect 514 55769 530 55775
rect 532 55769 548 55775
rect 525 55759 548 55768
rect 400 55749 404 55757
rect 498 55749 506 55759
rect 504 55725 506 55749
rect 514 55739 515 55759
rect 525 55734 528 55759
rect 547 55739 548 55759
rect 557 55749 564 55759
rect 514 55725 548 55729
rect 151 55678 156 55712
rect 174 55709 246 55717
rect 256 55709 328 55717
rect 336 55711 342 55719
rect 400 55714 404 55719
rect 180 55681 185 55709
rect 174 55673 246 55681
rect 256 55673 328 55681
rect 332 55679 336 55709
rect 400 55680 438 55714
rect 224 55643 226 55659
rect 196 55635 226 55643
rect 196 55631 232 55635
rect 196 55601 204 55631
rect 216 55601 232 55631
rect 224 55554 226 55601
rect 300 55574 308 55643
rect 332 55641 342 55679
rect 400 55671 404 55680
rect 454 55665 504 55667
rect 494 55661 548 55665
rect 494 55656 514 55661
rect 504 55641 506 55656
rect 336 55629 342 55641
rect 289 55564 308 55574
rect 300 55558 308 55564
rect 332 55595 342 55629
rect 400 55633 404 55641
rect 400 55599 408 55633
rect 434 55599 438 55633
rect 498 55631 506 55641
rect 514 55631 515 55651
rect 504 55615 506 55631
rect 525 55622 528 55656
rect 547 55631 548 55651
rect 557 55631 564 55641
rect 514 55615 530 55621
rect 532 55615 548 55621
rect 332 55567 373 55595
rect 332 55561 351 55567
rect 107 55507 119 55541
rect 129 55507 149 55541
rect 196 55520 204 55554
rect 216 55520 232 55554
rect 244 55548 257 55554
rect 278 55548 291 55558
rect 244 55524 291 55548
rect 300 55548 321 55558
rect 336 55551 351 55561
rect 300 55524 329 55548
rect 332 55533 351 55551
rect 361 55561 375 55567
rect 400 55561 411 55599
rect 562 55562 612 55564
rect 361 55533 381 55561
rect 400 55533 409 55561
rect 466 55553 497 55561
rect 565 55553 596 55561
rect 442 55546 500 55553
rect 466 55545 500 55546
rect 565 55545 599 55553
rect 244 55520 257 55524
rect 42 55441 46 55475
rect 72 55441 76 55475
rect 42 55394 76 55398
rect 42 55379 46 55394
rect 72 55379 76 55394
rect 38 55361 80 55379
rect 16 55355 102 55361
rect 144 55355 148 55507
rect 174 55483 181 55511
rect 224 55473 226 55520
rect 300 55511 308 55524
rect 278 55500 305 55511
rect 332 55483 342 55533
rect 400 55513 404 55533
rect 497 55529 500 55545
rect 596 55529 599 55545
rect 466 55528 500 55529
rect 442 55521 500 55528
rect 565 55521 599 55529
rect 612 55512 614 55562
rect 256 55473 328 55481
rect 336 55475 342 55483
rect 400 55475 404 55483
rect 196 55443 204 55473
rect 216 55443 232 55473
rect 196 55439 232 55443
rect 196 55431 226 55439
rect 224 55415 226 55431
rect 332 55403 336 55471
rect 400 55441 408 55475
rect 434 55441 438 55475
rect 454 55459 504 55461
rect 504 55443 506 55459
rect 514 55453 530 55459
rect 532 55453 548 55459
rect 525 55443 548 55452
rect 400 55433 404 55441
rect 498 55433 506 55443
rect 504 55409 506 55433
rect 514 55423 515 55443
rect 525 55418 528 55443
rect 547 55423 548 55443
rect 557 55433 564 55443
rect 514 55409 548 55413
rect 400 55403 442 55404
rect 174 55393 246 55401
rect 400 55396 404 55403
rect 295 55362 300 55396
rect 324 55362 329 55396
rect 367 55379 438 55396
rect 367 55362 442 55379
rect 400 55361 442 55362
rect 378 55355 464 55361
rect 38 55339 80 55355
rect 400 55339 442 55355
rect -25 55325 25 55327
rect 42 55325 76 55339
rect 404 55325 438 55339
rect 455 55325 505 55327
rect 557 55325 607 55327
rect 16 55317 102 55325
rect 378 55317 464 55325
rect 8 55283 17 55317
rect 18 55315 51 55317
rect 80 55315 100 55317
rect 18 55283 100 55315
rect 380 55315 404 55317
rect 429 55315 438 55317
rect 442 55315 462 55317
rect 16 55275 102 55283
rect 42 55259 76 55275
rect 16 55239 38 55245
rect 42 55236 76 55240
rect 80 55239 102 55245
rect 42 55206 46 55236
rect 72 55206 76 55236
rect 42 55125 46 55159
rect 72 55125 76 55159
rect -25 55088 25 55090
rect -8 55080 14 55087
rect -8 55079 17 55080
rect 25 55079 27 55088
rect -12 55072 38 55079
rect -12 55071 34 55072
rect -12 55067 8 55071
rect 0 55055 8 55067
rect 14 55055 34 55071
rect 0 55054 34 55055
rect 0 55047 38 55054
rect 14 55046 17 55047
rect 25 55038 27 55047
rect 42 55018 45 55108
rect 69 55093 80 55125
rect 107 55093 143 55121
rect 144 55093 148 55313
rect 332 55245 336 55313
rect 380 55283 462 55315
rect 463 55283 472 55317
rect 480 55283 497 55317
rect 378 55275 464 55283
rect 505 55275 507 55325
rect 514 55283 548 55317
rect 565 55283 582 55317
rect 607 55275 609 55325
rect 404 55259 438 55275
rect 400 55245 442 55246
rect 378 55239 404 55245
rect 442 55239 464 55245
rect 400 55238 404 55239
rect 174 55199 246 55207
rect 295 55204 300 55238
rect 324 55204 329 55238
rect 224 55169 226 55185
rect 196 55161 226 55169
rect 332 55167 336 55235
rect 367 55204 438 55238
rect 400 55197 404 55204
rect 454 55191 504 55193
rect 494 55187 548 55191
rect 494 55182 514 55187
rect 504 55167 506 55182
rect 196 55157 232 55161
rect 196 55127 204 55157
rect 216 55127 232 55157
rect 400 55159 404 55167
rect 107 55087 119 55093
rect 109 55059 119 55087
rect 129 55059 149 55093
rect 174 55089 181 55119
rect 224 55080 226 55127
rect 256 55119 328 55127
rect 332 55125 336 55155
rect 400 55125 408 55159
rect 434 55125 438 55159
rect 498 55157 506 55167
rect 514 55157 515 55177
rect 504 55141 506 55157
rect 525 55148 528 55182
rect 547 55157 548 55177
rect 557 55157 564 55167
rect 514 55141 530 55147
rect 532 55141 548 55147
rect 278 55089 305 55100
rect 42 54967 46 55001
rect 72 54967 76 55001
rect 38 54929 80 54930
rect 42 54888 76 54922
rect 79 54888 113 54922
rect 42 54809 46 54843
rect 72 54809 76 54843
rect -25 54772 25 54774
rect -8 54764 14 54771
rect -8 54763 17 54764
rect 25 54763 27 54772
rect -12 54756 38 54763
rect -12 54755 34 54756
rect -12 54751 8 54755
rect 0 54739 8 54751
rect 14 54739 34 54755
rect 0 54738 34 54739
rect 0 54731 38 54738
rect 14 54730 17 54731
rect 25 54722 27 54731
rect 42 54702 45 54792
rect 71 54761 80 54789
rect 69 54723 80 54761
rect 144 54751 148 55059
rect 196 55046 204 55080
rect 216 55046 232 55080
rect 244 55076 257 55080
rect 300 55076 308 55089
rect 332 55087 342 55125
rect 400 55117 404 55125
rect 336 55077 342 55087
rect 244 55052 291 55076
rect 244 55046 257 55052
rect 224 54999 226 55046
rect 278 55042 291 55052
rect 300 55052 329 55076
rect 332 55067 342 55077
rect 400 55077 409 55105
rect 562 55088 612 55090
rect 466 55079 497 55087
rect 565 55079 596 55087
rect 300 55042 321 55052
rect 300 55036 308 55042
rect 289 55026 308 55036
rect 196 54969 204 54999
rect 216 54969 232 54999
rect 196 54965 232 54969
rect 196 54957 226 54965
rect 300 54957 308 55026
rect 332 55033 351 55067
rect 361 55039 381 55067
rect 361 55033 375 55039
rect 400 55033 411 55077
rect 442 55072 500 55079
rect 466 55071 500 55072
rect 565 55071 599 55079
rect 497 55055 500 55071
rect 596 55055 599 55071
rect 466 55054 500 55055
rect 442 55047 500 55054
rect 565 55047 599 55055
rect 612 55038 614 55088
rect 332 55009 342 55033
rect 336 54997 342 55009
rect 224 54941 226 54957
rect 332 54929 342 54997
rect 400 55001 404 55009
rect 400 54967 408 55001
rect 434 54967 438 55001
rect 454 54985 504 54987
rect 504 54969 506 54985
rect 514 54979 530 54985
rect 532 54979 548 54985
rect 525 54969 548 54978
rect 400 54959 404 54967
rect 498 54959 506 54969
rect 504 54935 506 54959
rect 514 54949 515 54969
rect 525 54944 528 54969
rect 547 54949 548 54969
rect 557 54959 564 54969
rect 514 54935 548 54939
rect 151 54888 156 54922
rect 174 54919 246 54927
rect 256 54919 328 54927
rect 336 54921 342 54929
rect 400 54924 404 54929
rect 180 54891 185 54919
rect 174 54883 246 54891
rect 256 54883 328 54891
rect 332 54889 336 54919
rect 400 54890 438 54924
rect 224 54853 226 54869
rect 196 54845 226 54853
rect 196 54841 232 54845
rect 196 54811 204 54841
rect 216 54811 232 54841
rect 224 54764 226 54811
rect 300 54784 308 54853
rect 332 54851 342 54889
rect 400 54881 404 54890
rect 454 54875 504 54877
rect 494 54871 548 54875
rect 494 54866 514 54871
rect 504 54851 506 54866
rect 336 54839 342 54851
rect 289 54774 308 54784
rect 300 54768 308 54774
rect 332 54805 342 54839
rect 400 54843 404 54851
rect 400 54809 408 54843
rect 434 54809 438 54843
rect 498 54841 506 54851
rect 514 54841 515 54861
rect 504 54825 506 54841
rect 525 54832 528 54866
rect 547 54841 548 54861
rect 557 54841 564 54851
rect 514 54825 530 54831
rect 532 54825 548 54831
rect 332 54777 373 54805
rect 332 54771 351 54777
rect 107 54717 119 54751
rect 129 54717 149 54751
rect 196 54730 204 54764
rect 216 54730 232 54764
rect 244 54758 257 54764
rect 278 54758 291 54768
rect 244 54734 291 54758
rect 300 54758 321 54768
rect 336 54761 351 54771
rect 300 54734 329 54758
rect 332 54743 351 54761
rect 361 54771 375 54777
rect 400 54771 411 54809
rect 562 54772 612 54774
rect 361 54743 381 54771
rect 400 54743 409 54771
rect 466 54763 497 54771
rect 565 54763 596 54771
rect 442 54756 500 54763
rect 466 54755 500 54756
rect 565 54755 599 54763
rect 244 54730 257 54734
rect 42 54651 46 54685
rect 72 54651 76 54685
rect 42 54604 76 54608
rect 42 54589 46 54604
rect 72 54589 76 54604
rect 38 54571 80 54589
rect 16 54565 102 54571
rect 144 54565 148 54717
rect 174 54693 181 54721
rect 224 54683 226 54730
rect 300 54721 308 54734
rect 278 54710 305 54721
rect 332 54693 342 54743
rect 400 54723 404 54743
rect 497 54739 500 54755
rect 596 54739 599 54755
rect 466 54738 500 54739
rect 442 54731 500 54738
rect 565 54731 599 54739
rect 612 54722 614 54772
rect 256 54683 328 54691
rect 336 54685 342 54693
rect 400 54685 404 54693
rect 196 54653 204 54683
rect 216 54653 232 54683
rect 196 54649 232 54653
rect 196 54641 226 54649
rect 224 54625 226 54641
rect 332 54613 336 54681
rect 400 54651 408 54685
rect 434 54651 438 54685
rect 454 54669 504 54671
rect 504 54653 506 54669
rect 514 54663 530 54669
rect 532 54663 548 54669
rect 525 54653 548 54662
rect 400 54643 404 54651
rect 498 54643 506 54653
rect 504 54619 506 54643
rect 514 54633 515 54653
rect 525 54628 528 54653
rect 547 54633 548 54653
rect 557 54643 564 54653
rect 514 54619 548 54623
rect 400 54613 442 54614
rect 174 54603 246 54611
rect 400 54606 404 54613
rect 295 54572 300 54606
rect 324 54572 329 54606
rect 367 54589 438 54606
rect 367 54572 442 54589
rect 400 54571 442 54572
rect 378 54565 464 54571
rect 38 54549 80 54565
rect 400 54549 442 54565
rect -25 54535 25 54537
rect 42 54535 76 54549
rect 404 54535 438 54549
rect 455 54535 505 54537
rect 557 54535 607 54537
rect 16 54527 102 54535
rect 378 54527 464 54535
rect 8 54493 17 54527
rect 18 54525 51 54527
rect 80 54525 100 54527
rect 18 54493 100 54525
rect 380 54525 404 54527
rect 429 54525 438 54527
rect 442 54525 462 54527
rect 16 54485 102 54493
rect 42 54469 76 54485
rect 16 54449 38 54455
rect 42 54446 76 54450
rect 80 54449 102 54455
rect 42 54416 46 54446
rect 72 54416 76 54446
rect 42 54335 46 54369
rect 72 54335 76 54369
rect -25 54298 25 54300
rect -8 54290 14 54297
rect -8 54289 17 54290
rect 25 54289 27 54298
rect -12 54282 38 54289
rect -12 54281 34 54282
rect -12 54277 8 54281
rect 0 54265 8 54277
rect 14 54265 34 54281
rect 0 54264 34 54265
rect 0 54257 38 54264
rect 14 54256 17 54257
rect 25 54248 27 54257
rect 42 54228 45 54318
rect 69 54303 80 54335
rect 107 54303 143 54331
rect 144 54303 148 54523
rect 332 54455 336 54523
rect 380 54493 462 54525
rect 463 54493 472 54527
rect 480 54493 497 54527
rect 378 54485 464 54493
rect 505 54485 507 54535
rect 514 54493 548 54527
rect 565 54493 582 54527
rect 607 54485 609 54535
rect 404 54469 438 54485
rect 400 54455 442 54456
rect 378 54449 404 54455
rect 442 54449 464 54455
rect 400 54448 404 54449
rect 174 54409 246 54417
rect 295 54414 300 54448
rect 324 54414 329 54448
rect 224 54379 226 54395
rect 196 54371 226 54379
rect 332 54377 336 54445
rect 367 54414 438 54448
rect 400 54407 404 54414
rect 454 54401 504 54403
rect 494 54397 548 54401
rect 494 54392 514 54397
rect 504 54377 506 54392
rect 196 54367 232 54371
rect 196 54337 204 54367
rect 216 54337 232 54367
rect 400 54369 404 54377
rect 107 54297 119 54303
rect 109 54269 119 54297
rect 129 54269 149 54303
rect 174 54299 181 54329
rect 224 54290 226 54337
rect 256 54329 328 54337
rect 332 54335 336 54365
rect 400 54335 408 54369
rect 434 54335 438 54369
rect 498 54367 506 54377
rect 514 54367 515 54387
rect 504 54351 506 54367
rect 525 54358 528 54392
rect 547 54367 548 54387
rect 557 54367 564 54377
rect 514 54351 530 54357
rect 532 54351 548 54357
rect 278 54299 305 54310
rect 42 54177 46 54211
rect 72 54177 76 54211
rect 38 54139 80 54140
rect 42 54098 76 54132
rect 79 54098 113 54132
rect 42 54019 46 54053
rect 72 54019 76 54053
rect -25 53982 25 53984
rect -8 53974 14 53981
rect -8 53973 17 53974
rect 25 53973 27 53982
rect -12 53966 38 53973
rect -12 53965 34 53966
rect -12 53961 8 53965
rect 0 53949 8 53961
rect 14 53949 34 53965
rect 0 53948 34 53949
rect 0 53941 38 53948
rect 14 53940 17 53941
rect 25 53932 27 53941
rect 42 53912 45 54002
rect 71 53971 80 53999
rect 69 53933 80 53971
rect 144 53961 148 54269
rect 196 54256 204 54290
rect 216 54256 232 54290
rect 244 54286 257 54290
rect 300 54286 308 54299
rect 332 54297 342 54335
rect 400 54327 404 54335
rect 336 54287 342 54297
rect 244 54262 291 54286
rect 244 54256 257 54262
rect 224 54209 226 54256
rect 278 54252 291 54262
rect 300 54262 329 54286
rect 332 54277 342 54287
rect 400 54287 409 54315
rect 562 54298 612 54300
rect 466 54289 497 54297
rect 565 54289 596 54297
rect 300 54252 321 54262
rect 300 54246 308 54252
rect 289 54236 308 54246
rect 196 54179 204 54209
rect 216 54179 232 54209
rect 196 54175 232 54179
rect 196 54167 226 54175
rect 300 54167 308 54236
rect 332 54243 351 54277
rect 361 54249 381 54277
rect 361 54243 375 54249
rect 400 54243 411 54287
rect 442 54282 500 54289
rect 466 54281 500 54282
rect 565 54281 599 54289
rect 497 54265 500 54281
rect 596 54265 599 54281
rect 466 54264 500 54265
rect 442 54257 500 54264
rect 565 54257 599 54265
rect 612 54248 614 54298
rect 332 54219 342 54243
rect 336 54207 342 54219
rect 224 54151 226 54167
rect 332 54139 342 54207
rect 400 54211 404 54219
rect 400 54177 408 54211
rect 434 54177 438 54211
rect 454 54195 504 54197
rect 504 54179 506 54195
rect 514 54189 530 54195
rect 532 54189 548 54195
rect 525 54179 548 54188
rect 400 54169 404 54177
rect 498 54169 506 54179
rect 504 54145 506 54169
rect 514 54159 515 54179
rect 525 54154 528 54179
rect 547 54159 548 54179
rect 557 54169 564 54179
rect 514 54145 548 54149
rect 151 54098 156 54132
rect 174 54129 246 54137
rect 256 54129 328 54137
rect 336 54131 342 54139
rect 400 54134 404 54139
rect 180 54101 185 54129
rect 174 54093 246 54101
rect 256 54093 328 54101
rect 332 54099 336 54129
rect 400 54100 438 54134
rect 224 54063 226 54079
rect 196 54055 226 54063
rect 196 54051 232 54055
rect 196 54021 204 54051
rect 216 54021 232 54051
rect 224 53974 226 54021
rect 300 53994 308 54063
rect 332 54061 342 54099
rect 400 54091 404 54100
rect 454 54085 504 54087
rect 494 54081 548 54085
rect 494 54076 514 54081
rect 504 54061 506 54076
rect 336 54049 342 54061
rect 289 53984 308 53994
rect 300 53978 308 53984
rect 332 54015 342 54049
rect 400 54053 404 54061
rect 400 54019 408 54053
rect 434 54019 438 54053
rect 498 54051 506 54061
rect 514 54051 515 54071
rect 504 54035 506 54051
rect 525 54042 528 54076
rect 547 54051 548 54071
rect 557 54051 564 54061
rect 514 54035 530 54041
rect 532 54035 548 54041
rect 332 53987 373 54015
rect 332 53981 351 53987
rect 107 53927 119 53961
rect 129 53927 149 53961
rect 196 53940 204 53974
rect 216 53940 232 53974
rect 244 53968 257 53974
rect 278 53968 291 53978
rect 244 53944 291 53968
rect 300 53968 321 53978
rect 336 53971 351 53981
rect 300 53944 329 53968
rect 332 53953 351 53971
rect 361 53981 375 53987
rect 400 53981 411 54019
rect 562 53982 612 53984
rect 361 53953 381 53981
rect 400 53953 409 53981
rect 466 53973 497 53981
rect 565 53973 596 53981
rect 442 53966 500 53973
rect 466 53965 500 53966
rect 565 53965 599 53973
rect 244 53940 257 53944
rect 42 53861 46 53895
rect 72 53861 76 53895
rect 42 53814 76 53818
rect 42 53799 46 53814
rect 72 53799 76 53814
rect 38 53781 80 53799
rect 16 53775 102 53781
rect 144 53775 148 53927
rect 174 53903 181 53931
rect 224 53893 226 53940
rect 300 53931 308 53944
rect 278 53920 305 53931
rect 332 53903 342 53953
rect 400 53933 404 53953
rect 497 53949 500 53965
rect 596 53949 599 53965
rect 466 53948 500 53949
rect 442 53941 500 53948
rect 565 53941 599 53949
rect 612 53932 614 53982
rect 256 53893 328 53901
rect 336 53895 342 53903
rect 400 53895 404 53903
rect 196 53863 204 53893
rect 216 53863 232 53893
rect 196 53859 232 53863
rect 196 53851 226 53859
rect 224 53835 226 53851
rect 332 53823 336 53891
rect 400 53861 408 53895
rect 434 53861 438 53895
rect 454 53879 504 53881
rect 504 53863 506 53879
rect 514 53873 530 53879
rect 532 53873 548 53879
rect 525 53863 548 53872
rect 400 53853 404 53861
rect 498 53853 506 53863
rect 504 53829 506 53853
rect 514 53843 515 53863
rect 525 53838 528 53863
rect 547 53843 548 53863
rect 557 53853 564 53863
rect 514 53829 548 53833
rect 400 53823 442 53824
rect 174 53813 246 53821
rect 400 53816 404 53823
rect 295 53782 300 53816
rect 324 53782 329 53816
rect 367 53799 438 53816
rect 367 53782 442 53799
rect 400 53781 442 53782
rect 378 53775 464 53781
rect 38 53759 80 53775
rect 400 53759 442 53775
rect -25 53745 25 53747
rect 42 53745 76 53759
rect 404 53745 438 53759
rect 455 53745 505 53747
rect 557 53745 607 53747
rect 16 53737 102 53745
rect 378 53737 464 53745
rect 8 53703 17 53737
rect 18 53735 51 53737
rect 80 53735 100 53737
rect 18 53703 100 53735
rect 380 53735 404 53737
rect 429 53735 438 53737
rect 442 53735 462 53737
rect 16 53695 102 53703
rect 42 53679 76 53695
rect 16 53659 38 53665
rect 42 53656 76 53660
rect 80 53659 102 53665
rect 42 53626 46 53656
rect 72 53626 76 53656
rect 42 53545 46 53579
rect 72 53545 76 53579
rect -25 53508 25 53510
rect -8 53500 14 53507
rect -8 53499 17 53500
rect 25 53499 27 53508
rect -12 53492 38 53499
rect -12 53491 34 53492
rect -12 53487 8 53491
rect 0 53475 8 53487
rect 14 53475 34 53491
rect 0 53474 34 53475
rect 0 53467 38 53474
rect 14 53466 17 53467
rect 25 53458 27 53467
rect 42 53438 45 53528
rect 69 53513 80 53545
rect 107 53513 143 53541
rect 144 53513 148 53733
rect 332 53665 336 53733
rect 380 53703 462 53735
rect 463 53703 472 53737
rect 480 53703 497 53737
rect 378 53695 464 53703
rect 505 53695 507 53745
rect 514 53703 548 53737
rect 565 53703 582 53737
rect 607 53695 609 53745
rect 404 53679 438 53695
rect 400 53665 442 53666
rect 378 53659 404 53665
rect 442 53659 464 53665
rect 400 53658 404 53659
rect 174 53619 246 53627
rect 295 53624 300 53658
rect 324 53624 329 53658
rect 224 53589 226 53605
rect 196 53581 226 53589
rect 332 53587 336 53655
rect 367 53624 438 53658
rect 400 53617 404 53624
rect 454 53611 504 53613
rect 494 53607 548 53611
rect 494 53602 514 53607
rect 504 53587 506 53602
rect 196 53577 232 53581
rect 196 53547 204 53577
rect 216 53547 232 53577
rect 400 53579 404 53587
rect 107 53507 119 53513
rect 109 53479 119 53507
rect 129 53479 149 53513
rect 174 53509 181 53539
rect 224 53500 226 53547
rect 256 53539 328 53547
rect 332 53545 336 53575
rect 400 53545 408 53579
rect 434 53545 438 53579
rect 498 53577 506 53587
rect 514 53577 515 53597
rect 504 53561 506 53577
rect 525 53568 528 53602
rect 547 53577 548 53597
rect 557 53577 564 53587
rect 514 53561 530 53567
rect 532 53561 548 53567
rect 278 53509 305 53520
rect 42 53387 46 53421
rect 72 53387 76 53421
rect 38 53349 80 53350
rect 42 53308 76 53342
rect 79 53308 113 53342
rect 42 53229 46 53263
rect 72 53229 76 53263
rect -25 53192 25 53194
rect -8 53184 14 53191
rect -8 53183 17 53184
rect 25 53183 27 53192
rect -12 53176 38 53183
rect -12 53175 34 53176
rect -12 53171 8 53175
rect 0 53159 8 53171
rect 14 53159 34 53175
rect 0 53158 34 53159
rect 0 53151 38 53158
rect 14 53150 17 53151
rect 25 53142 27 53151
rect 42 53122 45 53212
rect 71 53181 80 53209
rect 69 53143 80 53181
rect 144 53171 148 53479
rect 196 53466 204 53500
rect 216 53466 232 53500
rect 244 53496 257 53500
rect 300 53496 308 53509
rect 332 53507 342 53545
rect 400 53537 404 53545
rect 336 53497 342 53507
rect 244 53472 291 53496
rect 244 53466 257 53472
rect 224 53419 226 53466
rect 278 53462 291 53472
rect 300 53472 329 53496
rect 332 53487 342 53497
rect 400 53497 409 53525
rect 562 53508 612 53510
rect 466 53499 497 53507
rect 565 53499 596 53507
rect 300 53462 321 53472
rect 300 53456 308 53462
rect 289 53446 308 53456
rect 196 53389 204 53419
rect 216 53389 232 53419
rect 196 53385 232 53389
rect 196 53377 226 53385
rect 300 53377 308 53446
rect 332 53453 351 53487
rect 361 53459 381 53487
rect 361 53453 375 53459
rect 400 53453 411 53497
rect 442 53492 500 53499
rect 466 53491 500 53492
rect 565 53491 599 53499
rect 497 53475 500 53491
rect 596 53475 599 53491
rect 466 53474 500 53475
rect 442 53467 500 53474
rect 565 53467 599 53475
rect 612 53458 614 53508
rect 332 53429 342 53453
rect 336 53417 342 53429
rect 224 53361 226 53377
rect 332 53349 342 53417
rect 400 53421 404 53429
rect 400 53387 408 53421
rect 434 53387 438 53421
rect 454 53405 504 53407
rect 504 53389 506 53405
rect 514 53399 530 53405
rect 532 53399 548 53405
rect 525 53389 548 53398
rect 400 53379 404 53387
rect 498 53379 506 53389
rect 504 53355 506 53379
rect 514 53369 515 53389
rect 525 53364 528 53389
rect 547 53369 548 53389
rect 557 53379 564 53389
rect 514 53355 548 53359
rect 151 53308 156 53342
rect 174 53339 246 53347
rect 256 53339 328 53347
rect 336 53341 342 53349
rect 400 53344 404 53349
rect 180 53311 185 53339
rect 174 53303 246 53311
rect 256 53303 328 53311
rect 332 53309 336 53339
rect 400 53310 438 53344
rect 224 53273 226 53289
rect 196 53265 226 53273
rect 196 53261 232 53265
rect 196 53231 204 53261
rect 216 53231 232 53261
rect 224 53184 226 53231
rect 300 53204 308 53273
rect 332 53271 342 53309
rect 400 53301 404 53310
rect 454 53295 504 53297
rect 494 53291 548 53295
rect 494 53286 514 53291
rect 504 53271 506 53286
rect 336 53259 342 53271
rect 289 53194 308 53204
rect 300 53188 308 53194
rect 332 53225 342 53259
rect 400 53263 404 53271
rect 400 53229 408 53263
rect 434 53229 438 53263
rect 498 53261 506 53271
rect 514 53261 515 53281
rect 504 53245 506 53261
rect 525 53252 528 53286
rect 547 53261 548 53281
rect 557 53261 564 53271
rect 514 53245 530 53251
rect 532 53245 548 53251
rect 332 53197 373 53225
rect 332 53191 351 53197
rect 107 53137 119 53171
rect 129 53137 149 53171
rect 196 53150 204 53184
rect 216 53150 232 53184
rect 244 53178 257 53184
rect 278 53178 291 53188
rect 244 53154 291 53178
rect 300 53178 321 53188
rect 336 53181 351 53191
rect 300 53154 329 53178
rect 332 53163 351 53181
rect 361 53191 375 53197
rect 400 53191 411 53229
rect 562 53192 612 53194
rect 361 53163 381 53191
rect 400 53163 409 53191
rect 466 53183 497 53191
rect 565 53183 596 53191
rect 442 53176 500 53183
rect 466 53175 500 53176
rect 565 53175 599 53183
rect 244 53150 257 53154
rect 42 53071 46 53105
rect 72 53071 76 53105
rect 42 53024 76 53028
rect 42 53009 46 53024
rect 72 53009 76 53024
rect 38 52991 80 53009
rect 16 52985 102 52991
rect 144 52985 148 53137
rect 174 53113 181 53141
rect 224 53103 226 53150
rect 300 53141 308 53154
rect 278 53130 305 53141
rect 332 53113 342 53163
rect 400 53143 404 53163
rect 497 53159 500 53175
rect 596 53159 599 53175
rect 466 53158 500 53159
rect 442 53151 500 53158
rect 565 53151 599 53159
rect 612 53142 614 53192
rect 256 53103 328 53111
rect 336 53105 342 53113
rect 400 53105 404 53113
rect 196 53073 204 53103
rect 216 53073 232 53103
rect 196 53069 232 53073
rect 196 53061 226 53069
rect 224 53045 226 53061
rect 332 53033 336 53101
rect 400 53071 408 53105
rect 434 53071 438 53105
rect 454 53089 504 53091
rect 504 53073 506 53089
rect 514 53083 530 53089
rect 532 53083 548 53089
rect 525 53073 548 53082
rect 400 53063 404 53071
rect 498 53063 506 53073
rect 504 53039 506 53063
rect 514 53053 515 53073
rect 525 53048 528 53073
rect 547 53053 548 53073
rect 557 53063 564 53073
rect 514 53039 548 53043
rect 400 53033 442 53034
rect 174 53023 246 53031
rect 400 53026 404 53033
rect 295 52992 300 53026
rect 324 52992 329 53026
rect 367 53009 438 53026
rect 367 52992 442 53009
rect 400 52991 442 52992
rect 378 52985 464 52991
rect 38 52969 80 52985
rect 400 52969 442 52985
rect -25 52955 25 52957
rect 42 52955 76 52969
rect 404 52955 438 52969
rect 455 52955 505 52957
rect 557 52955 607 52957
rect 16 52947 102 52955
rect 378 52947 464 52955
rect 8 52913 17 52947
rect 18 52945 51 52947
rect 80 52945 100 52947
rect 18 52913 100 52945
rect 380 52945 404 52947
rect 429 52945 438 52947
rect 442 52945 462 52947
rect 16 52905 102 52913
rect 42 52889 76 52905
rect 16 52869 38 52875
rect 42 52866 76 52870
rect 80 52869 102 52875
rect 42 52836 46 52866
rect 72 52836 76 52866
rect 42 52755 46 52789
rect 72 52755 76 52789
rect -25 52718 25 52720
rect -8 52710 14 52717
rect -8 52709 17 52710
rect 25 52709 27 52718
rect -12 52702 38 52709
rect -12 52701 34 52702
rect -12 52697 8 52701
rect 0 52685 8 52697
rect 14 52685 34 52701
rect 0 52684 34 52685
rect 0 52677 38 52684
rect 14 52676 17 52677
rect 25 52668 27 52677
rect 42 52648 45 52738
rect 69 52723 80 52755
rect 107 52723 143 52751
rect 144 52723 148 52943
rect 332 52875 336 52943
rect 380 52913 462 52945
rect 463 52913 472 52947
rect 480 52913 497 52947
rect 378 52905 464 52913
rect 505 52905 507 52955
rect 514 52913 548 52947
rect 565 52913 582 52947
rect 607 52905 609 52955
rect 404 52889 438 52905
rect 400 52875 442 52876
rect 378 52869 404 52875
rect 442 52869 464 52875
rect 400 52868 404 52869
rect 174 52829 246 52837
rect 295 52834 300 52868
rect 324 52834 329 52868
rect 224 52799 226 52815
rect 196 52791 226 52799
rect 332 52797 336 52865
rect 367 52834 438 52868
rect 400 52827 404 52834
rect 454 52821 504 52823
rect 494 52817 548 52821
rect 494 52812 514 52817
rect 504 52797 506 52812
rect 196 52787 232 52791
rect 196 52757 204 52787
rect 216 52757 232 52787
rect 400 52789 404 52797
rect 107 52717 119 52723
rect 109 52689 119 52717
rect 129 52689 149 52723
rect 174 52719 181 52749
rect 224 52710 226 52757
rect 256 52749 328 52757
rect 332 52755 336 52785
rect 400 52755 408 52789
rect 434 52755 438 52789
rect 498 52787 506 52797
rect 514 52787 515 52807
rect 504 52771 506 52787
rect 525 52778 528 52812
rect 547 52787 548 52807
rect 557 52787 564 52797
rect 514 52771 530 52777
rect 532 52771 548 52777
rect 278 52719 305 52730
rect 42 52597 46 52631
rect 72 52597 76 52631
rect 38 52559 80 52560
rect 42 52518 76 52552
rect 79 52518 113 52552
rect 42 52439 46 52473
rect 72 52439 76 52473
rect -25 52402 25 52404
rect -8 52394 14 52401
rect -8 52393 17 52394
rect 25 52393 27 52402
rect -12 52386 38 52393
rect -12 52385 34 52386
rect -12 52381 8 52385
rect 0 52369 8 52381
rect 14 52369 34 52385
rect 0 52368 34 52369
rect 0 52361 38 52368
rect 14 52360 17 52361
rect 25 52352 27 52361
rect 42 52332 45 52422
rect 71 52391 80 52419
rect 69 52353 80 52391
rect 144 52381 148 52689
rect 196 52676 204 52710
rect 216 52676 232 52710
rect 244 52706 257 52710
rect 300 52706 308 52719
rect 332 52717 342 52755
rect 400 52747 404 52755
rect 336 52707 342 52717
rect 244 52682 291 52706
rect 244 52676 257 52682
rect 224 52629 226 52676
rect 278 52672 291 52682
rect 300 52682 329 52706
rect 332 52697 342 52707
rect 400 52707 409 52735
rect 562 52718 612 52720
rect 466 52709 497 52717
rect 565 52709 596 52717
rect 300 52672 321 52682
rect 300 52666 308 52672
rect 289 52656 308 52666
rect 196 52599 204 52629
rect 216 52599 232 52629
rect 196 52595 232 52599
rect 196 52587 226 52595
rect 300 52587 308 52656
rect 332 52663 351 52697
rect 361 52669 381 52697
rect 361 52663 375 52669
rect 400 52663 411 52707
rect 442 52702 500 52709
rect 466 52701 500 52702
rect 565 52701 599 52709
rect 497 52685 500 52701
rect 596 52685 599 52701
rect 466 52684 500 52685
rect 442 52677 500 52684
rect 565 52677 599 52685
rect 612 52668 614 52718
rect 332 52639 342 52663
rect 336 52627 342 52639
rect 224 52571 226 52587
rect 332 52559 342 52627
rect 400 52631 404 52639
rect 400 52597 408 52631
rect 434 52597 438 52631
rect 454 52615 504 52617
rect 504 52599 506 52615
rect 514 52609 530 52615
rect 532 52609 548 52615
rect 525 52599 548 52608
rect 400 52589 404 52597
rect 498 52589 506 52599
rect 504 52565 506 52589
rect 514 52579 515 52599
rect 525 52574 528 52599
rect 547 52579 548 52599
rect 557 52589 564 52599
rect 514 52565 548 52569
rect 151 52518 156 52552
rect 174 52549 246 52557
rect 256 52549 328 52557
rect 336 52551 342 52559
rect 400 52554 404 52559
rect 180 52521 185 52549
rect 174 52513 246 52521
rect 256 52513 328 52521
rect 332 52519 336 52549
rect 400 52520 438 52554
rect 224 52483 226 52499
rect 196 52475 226 52483
rect 196 52471 232 52475
rect 196 52441 204 52471
rect 216 52441 232 52471
rect 224 52394 226 52441
rect 300 52414 308 52483
rect 332 52481 342 52519
rect 400 52511 404 52520
rect 454 52505 504 52507
rect 494 52501 548 52505
rect 494 52496 514 52501
rect 504 52481 506 52496
rect 336 52469 342 52481
rect 289 52404 308 52414
rect 300 52398 308 52404
rect 332 52435 342 52469
rect 400 52473 404 52481
rect 400 52439 408 52473
rect 434 52439 438 52473
rect 498 52471 506 52481
rect 514 52471 515 52491
rect 504 52455 506 52471
rect 525 52462 528 52496
rect 547 52471 548 52491
rect 557 52471 564 52481
rect 514 52455 530 52461
rect 532 52455 548 52461
rect 332 52407 373 52435
rect 332 52401 351 52407
rect 107 52347 119 52381
rect 129 52347 149 52381
rect 196 52360 204 52394
rect 216 52360 232 52394
rect 244 52388 257 52394
rect 278 52388 291 52398
rect 244 52364 291 52388
rect 300 52388 321 52398
rect 336 52391 351 52401
rect 300 52364 329 52388
rect 332 52373 351 52391
rect 361 52401 375 52407
rect 400 52401 411 52439
rect 562 52402 612 52404
rect 361 52373 381 52401
rect 400 52373 409 52401
rect 466 52393 497 52401
rect 565 52393 596 52401
rect 442 52386 500 52393
rect 466 52385 500 52386
rect 565 52385 599 52393
rect 244 52360 257 52364
rect 42 52281 46 52315
rect 72 52281 76 52315
rect 42 52234 76 52238
rect 42 52219 46 52234
rect 72 52219 76 52234
rect 38 52201 80 52219
rect 16 52195 102 52201
rect 144 52195 148 52347
rect 174 52323 181 52351
rect 224 52313 226 52360
rect 300 52351 308 52364
rect 278 52340 305 52351
rect 332 52323 342 52373
rect 400 52353 404 52373
rect 497 52369 500 52385
rect 596 52369 599 52385
rect 466 52368 500 52369
rect 442 52361 500 52368
rect 565 52361 599 52369
rect 612 52352 614 52402
rect 256 52313 328 52321
rect 336 52315 342 52323
rect 400 52315 404 52323
rect 196 52283 204 52313
rect 216 52283 232 52313
rect 196 52279 232 52283
rect 196 52271 226 52279
rect 224 52255 226 52271
rect 332 52243 336 52311
rect 400 52281 408 52315
rect 434 52281 438 52315
rect 454 52299 504 52301
rect 504 52283 506 52299
rect 514 52293 530 52299
rect 532 52293 548 52299
rect 525 52283 548 52292
rect 400 52273 404 52281
rect 498 52273 506 52283
rect 504 52249 506 52273
rect 514 52263 515 52283
rect 525 52258 528 52283
rect 547 52263 548 52283
rect 557 52273 564 52283
rect 514 52249 548 52253
rect 400 52243 442 52244
rect 174 52233 246 52241
rect 400 52236 404 52243
rect 295 52202 300 52236
rect 324 52202 329 52236
rect 367 52219 438 52236
rect 367 52202 442 52219
rect 400 52201 442 52202
rect 378 52195 464 52201
rect 38 52179 80 52195
rect 400 52179 442 52195
rect -25 52165 25 52167
rect 42 52165 76 52179
rect 404 52165 438 52179
rect 455 52165 505 52167
rect 557 52165 607 52167
rect 16 52157 102 52165
rect 378 52157 464 52165
rect 8 52123 17 52157
rect 18 52155 51 52157
rect 80 52155 100 52157
rect 18 52123 100 52155
rect 380 52155 404 52157
rect 429 52155 438 52157
rect 442 52155 462 52157
rect 16 52115 102 52123
rect 42 52099 76 52115
rect 16 52079 38 52085
rect 42 52076 76 52080
rect 80 52079 102 52085
rect 42 52046 46 52076
rect 72 52046 76 52076
rect 42 51965 46 51999
rect 72 51965 76 51999
rect -25 51928 25 51930
rect -8 51920 14 51927
rect -8 51919 17 51920
rect 25 51919 27 51928
rect -12 51912 38 51919
rect -12 51911 34 51912
rect -12 51907 8 51911
rect 0 51895 8 51907
rect 14 51895 34 51911
rect 0 51894 34 51895
rect 0 51887 38 51894
rect 14 51886 17 51887
rect 25 51878 27 51887
rect 42 51858 45 51948
rect 69 51933 80 51965
rect 107 51933 143 51961
rect 144 51933 148 52153
rect 332 52085 336 52153
rect 380 52123 462 52155
rect 463 52123 472 52157
rect 480 52123 497 52157
rect 378 52115 464 52123
rect 505 52115 507 52165
rect 514 52123 548 52157
rect 565 52123 582 52157
rect 607 52115 609 52165
rect 404 52099 438 52115
rect 400 52085 442 52086
rect 378 52079 404 52085
rect 442 52079 464 52085
rect 400 52078 404 52079
rect 174 52039 246 52047
rect 295 52044 300 52078
rect 324 52044 329 52078
rect 224 52009 226 52025
rect 196 52001 226 52009
rect 332 52007 336 52075
rect 367 52044 438 52078
rect 400 52037 404 52044
rect 454 52031 504 52033
rect 494 52027 548 52031
rect 494 52022 514 52027
rect 504 52007 506 52022
rect 196 51997 232 52001
rect 196 51967 204 51997
rect 216 51967 232 51997
rect 400 51999 404 52007
rect 107 51927 119 51933
rect 109 51899 119 51927
rect 129 51899 149 51933
rect 174 51929 181 51959
rect 224 51920 226 51967
rect 256 51959 328 51967
rect 332 51965 336 51995
rect 400 51965 408 51999
rect 434 51965 438 51999
rect 498 51997 506 52007
rect 514 51997 515 52017
rect 504 51981 506 51997
rect 525 51988 528 52022
rect 547 51997 548 52017
rect 557 51997 564 52007
rect 514 51981 530 51987
rect 532 51981 548 51987
rect 278 51929 305 51940
rect 42 51807 46 51841
rect 72 51807 76 51841
rect 38 51769 80 51770
rect 42 51728 76 51762
rect 79 51728 113 51762
rect 42 51649 46 51683
rect 72 51649 76 51683
rect -25 51612 25 51614
rect -8 51604 14 51611
rect -8 51603 17 51604
rect 25 51603 27 51612
rect -12 51596 38 51603
rect -12 51595 34 51596
rect -12 51591 8 51595
rect 0 51579 8 51591
rect 14 51579 34 51595
rect 0 51578 34 51579
rect 0 51571 38 51578
rect 14 51570 17 51571
rect 25 51562 27 51571
rect 42 51542 45 51632
rect 71 51601 80 51629
rect 69 51563 80 51601
rect 144 51591 148 51899
rect 196 51886 204 51920
rect 216 51886 232 51920
rect 244 51916 257 51920
rect 300 51916 308 51929
rect 332 51927 342 51965
rect 400 51957 404 51965
rect 336 51917 342 51927
rect 244 51892 291 51916
rect 244 51886 257 51892
rect 224 51839 226 51886
rect 278 51882 291 51892
rect 300 51892 329 51916
rect 332 51907 342 51917
rect 400 51917 409 51945
rect 562 51928 612 51930
rect 466 51919 497 51927
rect 565 51919 596 51927
rect 300 51882 321 51892
rect 300 51876 308 51882
rect 289 51866 308 51876
rect 196 51809 204 51839
rect 216 51809 232 51839
rect 196 51805 232 51809
rect 196 51797 226 51805
rect 300 51797 308 51866
rect 332 51873 351 51907
rect 361 51879 381 51907
rect 361 51873 375 51879
rect 400 51873 411 51917
rect 442 51912 500 51919
rect 466 51911 500 51912
rect 565 51911 599 51919
rect 497 51895 500 51911
rect 596 51895 599 51911
rect 466 51894 500 51895
rect 442 51887 500 51894
rect 565 51887 599 51895
rect 612 51878 614 51928
rect 332 51849 342 51873
rect 336 51837 342 51849
rect 224 51781 226 51797
rect 332 51769 342 51837
rect 400 51841 404 51849
rect 400 51807 408 51841
rect 434 51807 438 51841
rect 454 51825 504 51827
rect 504 51809 506 51825
rect 514 51819 530 51825
rect 532 51819 548 51825
rect 525 51809 548 51818
rect 400 51799 404 51807
rect 498 51799 506 51809
rect 504 51775 506 51799
rect 514 51789 515 51809
rect 525 51784 528 51809
rect 547 51789 548 51809
rect 557 51799 564 51809
rect 514 51775 548 51779
rect 151 51728 156 51762
rect 174 51759 246 51767
rect 256 51759 328 51767
rect 336 51761 342 51769
rect 400 51764 404 51769
rect 180 51731 185 51759
rect 174 51723 246 51731
rect 256 51723 328 51731
rect 332 51729 336 51759
rect 400 51730 438 51764
rect 224 51693 226 51709
rect 196 51685 226 51693
rect 196 51681 232 51685
rect 196 51651 204 51681
rect 216 51651 232 51681
rect 224 51604 226 51651
rect 300 51624 308 51693
rect 332 51691 342 51729
rect 400 51721 404 51730
rect 454 51715 504 51717
rect 494 51711 548 51715
rect 494 51706 514 51711
rect 504 51691 506 51706
rect 336 51679 342 51691
rect 289 51614 308 51624
rect 300 51608 308 51614
rect 332 51645 342 51679
rect 400 51683 404 51691
rect 400 51649 408 51683
rect 434 51649 438 51683
rect 498 51681 506 51691
rect 514 51681 515 51701
rect 504 51665 506 51681
rect 525 51672 528 51706
rect 547 51681 548 51701
rect 557 51681 564 51691
rect 514 51665 530 51671
rect 532 51665 548 51671
rect 332 51617 373 51645
rect 332 51611 351 51617
rect 107 51557 119 51591
rect 129 51557 149 51591
rect 196 51570 204 51604
rect 216 51570 232 51604
rect 244 51598 257 51604
rect 278 51598 291 51608
rect 244 51574 291 51598
rect 300 51598 321 51608
rect 336 51601 351 51611
rect 300 51574 329 51598
rect 332 51583 351 51601
rect 361 51611 375 51617
rect 400 51611 411 51649
rect 562 51612 612 51614
rect 361 51583 381 51611
rect 400 51583 409 51611
rect 466 51603 497 51611
rect 565 51603 596 51611
rect 442 51596 500 51603
rect 466 51595 500 51596
rect 565 51595 599 51603
rect 244 51570 257 51574
rect 42 51491 46 51525
rect 72 51491 76 51525
rect 42 51444 76 51448
rect 42 51429 46 51444
rect 72 51429 76 51444
rect 38 51411 80 51429
rect 16 51405 102 51411
rect 144 51405 148 51557
rect 174 51533 181 51561
rect 224 51523 226 51570
rect 300 51561 308 51574
rect 278 51550 305 51561
rect 332 51533 342 51583
rect 400 51563 404 51583
rect 497 51579 500 51595
rect 596 51579 599 51595
rect 466 51578 500 51579
rect 442 51571 500 51578
rect 565 51571 599 51579
rect 612 51562 614 51612
rect 256 51523 328 51531
rect 336 51525 342 51533
rect 400 51525 404 51533
rect 196 51493 204 51523
rect 216 51493 232 51523
rect 196 51489 232 51493
rect 196 51481 226 51489
rect 224 51465 226 51481
rect 332 51453 336 51521
rect 400 51491 408 51525
rect 434 51491 438 51525
rect 454 51509 504 51511
rect 504 51493 506 51509
rect 514 51503 530 51509
rect 532 51503 548 51509
rect 525 51493 548 51502
rect 400 51483 404 51491
rect 498 51483 506 51493
rect 504 51459 506 51483
rect 514 51473 515 51493
rect 525 51468 528 51493
rect 547 51473 548 51493
rect 557 51483 564 51493
rect 514 51459 548 51463
rect 400 51453 442 51454
rect 174 51443 246 51451
rect 400 51446 404 51453
rect 295 51412 300 51446
rect 324 51412 329 51446
rect 367 51429 438 51446
rect 367 51412 442 51429
rect 400 51411 442 51412
rect 378 51405 464 51411
rect 38 51389 80 51405
rect 400 51389 442 51405
rect -25 51375 25 51377
rect 42 51375 76 51389
rect 404 51375 438 51389
rect 455 51375 505 51377
rect 557 51375 607 51377
rect 16 51367 102 51375
rect 378 51367 464 51375
rect 8 51333 17 51367
rect 18 51365 51 51367
rect 80 51365 100 51367
rect 18 51333 100 51365
rect 380 51365 404 51367
rect 429 51365 438 51367
rect 442 51365 462 51367
rect 16 51325 102 51333
rect 42 51309 76 51325
rect 16 51289 38 51295
rect 42 51286 76 51290
rect 80 51289 102 51295
rect 42 51256 46 51286
rect 72 51256 76 51286
rect 42 51175 46 51209
rect 72 51175 76 51209
rect -25 51138 25 51140
rect -8 51130 14 51137
rect -8 51129 17 51130
rect 25 51129 27 51138
rect -12 51122 38 51129
rect -12 51121 34 51122
rect -12 51117 8 51121
rect 0 51105 8 51117
rect 14 51105 34 51121
rect 0 51104 34 51105
rect 0 51097 38 51104
rect 14 51096 17 51097
rect 25 51088 27 51097
rect 42 51068 45 51158
rect 69 51143 80 51175
rect 107 51143 143 51171
rect 144 51143 148 51363
rect 332 51295 336 51363
rect 380 51333 462 51365
rect 463 51333 472 51367
rect 480 51333 497 51367
rect 378 51325 464 51333
rect 505 51325 507 51375
rect 514 51333 548 51367
rect 565 51333 582 51367
rect 607 51325 609 51375
rect 404 51309 438 51325
rect 400 51295 442 51296
rect 378 51289 404 51295
rect 442 51289 464 51295
rect 400 51288 404 51289
rect 174 51249 246 51257
rect 295 51254 300 51288
rect 324 51254 329 51288
rect 224 51219 226 51235
rect 196 51211 226 51219
rect 332 51217 336 51285
rect 367 51254 438 51288
rect 400 51247 404 51254
rect 454 51241 504 51243
rect 494 51237 548 51241
rect 494 51232 514 51237
rect 504 51217 506 51232
rect 196 51207 232 51211
rect 196 51177 204 51207
rect 216 51177 232 51207
rect 400 51209 404 51217
rect 107 51137 119 51143
rect 109 51109 119 51137
rect 129 51109 149 51143
rect 174 51139 181 51169
rect 224 51130 226 51177
rect 256 51169 328 51177
rect 332 51175 336 51205
rect 400 51175 408 51209
rect 434 51175 438 51209
rect 498 51207 506 51217
rect 514 51207 515 51227
rect 504 51191 506 51207
rect 525 51198 528 51232
rect 547 51207 548 51227
rect 557 51207 564 51217
rect 514 51191 530 51197
rect 532 51191 548 51197
rect 278 51139 305 51150
rect 42 51017 46 51051
rect 72 51017 76 51051
rect 38 50979 80 50980
rect 42 50938 76 50972
rect 79 50938 113 50972
rect 42 50859 46 50893
rect 72 50859 76 50893
rect -25 50822 25 50824
rect -8 50814 14 50821
rect -8 50813 17 50814
rect 25 50813 27 50822
rect -12 50806 38 50813
rect -12 50805 34 50806
rect -12 50801 8 50805
rect 0 50789 8 50801
rect 14 50789 34 50805
rect 0 50788 34 50789
rect 0 50781 38 50788
rect 14 50780 17 50781
rect 25 50772 27 50781
rect 42 50752 45 50842
rect 71 50811 80 50839
rect 69 50773 80 50811
rect 144 50801 148 51109
rect 196 51096 204 51130
rect 216 51096 232 51130
rect 244 51126 257 51130
rect 300 51126 308 51139
rect 332 51137 342 51175
rect 400 51167 404 51175
rect 336 51127 342 51137
rect 244 51102 291 51126
rect 244 51096 257 51102
rect 224 51049 226 51096
rect 278 51092 291 51102
rect 300 51102 329 51126
rect 332 51117 342 51127
rect 400 51127 409 51155
rect 562 51138 612 51140
rect 466 51129 497 51137
rect 565 51129 596 51137
rect 300 51092 321 51102
rect 300 51086 308 51092
rect 289 51076 308 51086
rect 196 51019 204 51049
rect 216 51019 232 51049
rect 196 51015 232 51019
rect 196 51007 226 51015
rect 300 51007 308 51076
rect 332 51083 351 51117
rect 361 51089 381 51117
rect 361 51083 375 51089
rect 400 51083 411 51127
rect 442 51122 500 51129
rect 466 51121 500 51122
rect 565 51121 599 51129
rect 497 51105 500 51121
rect 596 51105 599 51121
rect 466 51104 500 51105
rect 442 51097 500 51104
rect 565 51097 599 51105
rect 612 51088 614 51138
rect 332 51059 342 51083
rect 336 51047 342 51059
rect 224 50991 226 51007
rect 332 50979 342 51047
rect 400 51051 404 51059
rect 400 51017 408 51051
rect 434 51017 438 51051
rect 454 51035 504 51037
rect 504 51019 506 51035
rect 514 51029 530 51035
rect 532 51029 548 51035
rect 525 51019 548 51028
rect 400 51009 404 51017
rect 498 51009 506 51019
rect 504 50985 506 51009
rect 514 50999 515 51019
rect 525 50994 528 51019
rect 547 50999 548 51019
rect 557 51009 564 51019
rect 514 50985 548 50989
rect 151 50938 156 50972
rect 174 50969 246 50977
rect 256 50969 328 50977
rect 336 50971 342 50979
rect 400 50974 404 50979
rect 180 50941 185 50969
rect 174 50933 246 50941
rect 256 50933 328 50941
rect 332 50939 336 50969
rect 400 50940 438 50974
rect 224 50903 226 50919
rect 196 50895 226 50903
rect 196 50891 232 50895
rect 196 50861 204 50891
rect 216 50861 232 50891
rect 224 50814 226 50861
rect 300 50834 308 50903
rect 332 50901 342 50939
rect 400 50931 404 50940
rect 454 50925 504 50927
rect 494 50921 548 50925
rect 494 50916 514 50921
rect 504 50901 506 50916
rect 336 50889 342 50901
rect 289 50824 308 50834
rect 300 50818 308 50824
rect 332 50855 342 50889
rect 400 50893 404 50901
rect 400 50859 408 50893
rect 434 50859 438 50893
rect 498 50891 506 50901
rect 514 50891 515 50911
rect 504 50875 506 50891
rect 525 50882 528 50916
rect 547 50891 548 50911
rect 557 50891 564 50901
rect 514 50875 530 50881
rect 532 50875 548 50881
rect 332 50827 373 50855
rect 332 50821 351 50827
rect 107 50767 119 50801
rect 129 50767 149 50801
rect 196 50780 204 50814
rect 216 50780 232 50814
rect 244 50808 257 50814
rect 278 50808 291 50818
rect 244 50784 291 50808
rect 300 50808 321 50818
rect 336 50811 351 50821
rect 300 50784 329 50808
rect 332 50793 351 50811
rect 361 50821 375 50827
rect 400 50821 411 50859
rect 562 50822 612 50824
rect 361 50793 381 50821
rect 400 50793 409 50821
rect 466 50813 497 50821
rect 565 50813 596 50821
rect 442 50806 500 50813
rect 466 50805 500 50806
rect 565 50805 599 50813
rect 244 50780 257 50784
rect 42 50701 46 50735
rect 72 50701 76 50735
rect 42 50654 76 50658
rect 42 50639 46 50654
rect 72 50639 76 50654
rect 38 50621 80 50639
rect 16 50615 102 50621
rect 144 50615 148 50767
rect 174 50743 181 50771
rect 224 50733 226 50780
rect 300 50771 308 50784
rect 278 50760 305 50771
rect 332 50743 342 50793
rect 400 50773 404 50793
rect 497 50789 500 50805
rect 596 50789 599 50805
rect 466 50788 500 50789
rect 442 50781 500 50788
rect 565 50781 599 50789
rect 612 50772 614 50822
rect 256 50733 328 50741
rect 336 50735 342 50743
rect 400 50735 404 50743
rect 196 50703 204 50733
rect 216 50703 232 50733
rect 196 50699 232 50703
rect 196 50691 226 50699
rect 224 50675 226 50691
rect 332 50663 336 50731
rect 400 50701 408 50735
rect 434 50701 438 50735
rect 454 50719 504 50721
rect 504 50703 506 50719
rect 514 50713 530 50719
rect 532 50713 548 50719
rect 525 50703 548 50712
rect 400 50693 404 50701
rect 498 50693 506 50703
rect 504 50669 506 50693
rect 514 50683 515 50703
rect 525 50678 528 50703
rect 547 50683 548 50703
rect 557 50693 564 50703
rect 514 50669 548 50673
rect 400 50663 442 50664
rect 174 50653 246 50661
rect 400 50656 404 50663
rect 295 50622 300 50656
rect 324 50622 329 50656
rect 367 50639 438 50656
rect 367 50622 442 50639
rect 400 50621 442 50622
rect 378 50615 464 50621
rect 38 50599 80 50615
rect 400 50599 442 50615
rect -25 50585 25 50587
rect 42 50585 76 50599
rect 404 50585 438 50599
rect 455 50585 505 50587
rect 557 50585 607 50587
rect 16 50577 102 50585
rect 378 50577 464 50585
rect 8 50543 17 50577
rect 18 50575 51 50577
rect 80 50575 100 50577
rect 18 50543 100 50575
rect 380 50575 404 50577
rect 429 50575 438 50577
rect 442 50575 462 50577
rect 16 50535 102 50543
rect 42 50519 76 50535
rect 16 50499 38 50505
rect 42 50496 76 50500
rect 80 50499 102 50505
rect 42 50466 46 50496
rect 72 50466 76 50496
rect 42 50385 46 50419
rect 72 50385 76 50419
rect -25 50348 25 50350
rect -8 50340 14 50347
rect -8 50339 17 50340
rect 25 50339 27 50348
rect -12 50332 38 50339
rect -12 50331 34 50332
rect -12 50327 8 50331
rect 0 50315 8 50327
rect 14 50315 34 50331
rect 0 50314 34 50315
rect 0 50307 38 50314
rect 14 50306 17 50307
rect 25 50298 27 50307
rect 42 50278 45 50368
rect 69 50353 80 50385
rect 107 50353 143 50381
rect 144 50353 148 50573
rect 332 50505 336 50573
rect 380 50543 462 50575
rect 463 50543 472 50577
rect 480 50543 497 50577
rect 378 50535 464 50543
rect 505 50535 507 50585
rect 514 50543 548 50577
rect 565 50543 582 50577
rect 607 50535 609 50585
rect 404 50519 438 50535
rect 400 50505 442 50506
rect 378 50499 404 50505
rect 442 50499 464 50505
rect 400 50498 404 50499
rect 174 50459 246 50467
rect 295 50464 300 50498
rect 324 50464 329 50498
rect 224 50429 226 50445
rect 196 50421 226 50429
rect 332 50427 336 50495
rect 367 50464 438 50498
rect 400 50457 404 50464
rect 454 50451 504 50453
rect 494 50447 548 50451
rect 494 50442 514 50447
rect 504 50427 506 50442
rect 196 50417 232 50421
rect 196 50387 204 50417
rect 216 50387 232 50417
rect 400 50419 404 50427
rect 107 50347 119 50353
rect 109 50319 119 50347
rect 129 50319 149 50353
rect 174 50349 181 50379
rect 224 50340 226 50387
rect 256 50379 328 50387
rect 332 50385 336 50415
rect 400 50385 408 50419
rect 434 50385 438 50419
rect 498 50417 506 50427
rect 514 50417 515 50437
rect 504 50401 506 50417
rect 525 50408 528 50442
rect 547 50417 548 50437
rect 557 50417 564 50427
rect 514 50401 530 50407
rect 532 50401 548 50407
rect 278 50349 305 50360
rect 42 50227 46 50261
rect 72 50227 76 50261
rect 38 50189 80 50190
rect 42 50148 76 50182
rect 79 50148 113 50182
rect 42 50069 46 50103
rect 72 50069 76 50103
rect -25 50032 25 50034
rect -8 50024 14 50031
rect -8 50023 17 50024
rect 25 50023 27 50032
rect -12 50016 38 50023
rect -12 50015 34 50016
rect -12 50011 8 50015
rect 0 49999 8 50011
rect 14 49999 34 50015
rect 0 49998 34 49999
rect 0 49991 38 49998
rect 14 49990 17 49991
rect 25 49982 27 49991
rect 42 49962 45 50052
rect 71 50021 80 50049
rect 69 49983 80 50021
rect 144 50011 148 50319
rect 196 50306 204 50340
rect 216 50306 232 50340
rect 244 50336 257 50340
rect 300 50336 308 50349
rect 332 50347 342 50385
rect 400 50377 404 50385
rect 336 50337 342 50347
rect 244 50312 291 50336
rect 244 50306 257 50312
rect 224 50259 226 50306
rect 278 50302 291 50312
rect 300 50312 329 50336
rect 332 50327 342 50337
rect 400 50337 409 50365
rect 562 50348 612 50350
rect 466 50339 497 50347
rect 565 50339 596 50347
rect 300 50302 321 50312
rect 300 50296 308 50302
rect 289 50286 308 50296
rect 196 50229 204 50259
rect 216 50229 232 50259
rect 196 50225 232 50229
rect 196 50217 226 50225
rect 300 50217 308 50286
rect 332 50293 351 50327
rect 361 50299 381 50327
rect 361 50293 375 50299
rect 400 50293 411 50337
rect 442 50332 500 50339
rect 466 50331 500 50332
rect 565 50331 599 50339
rect 497 50315 500 50331
rect 596 50315 599 50331
rect 466 50314 500 50315
rect 442 50307 500 50314
rect 565 50307 599 50315
rect 612 50298 614 50348
rect 332 50269 342 50293
rect 336 50257 342 50269
rect 224 50201 226 50217
rect 332 50189 342 50257
rect 400 50261 404 50269
rect 400 50227 408 50261
rect 434 50227 438 50261
rect 454 50245 504 50247
rect 504 50229 506 50245
rect 514 50239 530 50245
rect 532 50239 548 50245
rect 525 50229 548 50238
rect 400 50219 404 50227
rect 498 50219 506 50229
rect 504 50195 506 50219
rect 514 50209 515 50229
rect 525 50204 528 50229
rect 547 50209 548 50229
rect 557 50219 564 50229
rect 514 50195 548 50199
rect 151 50148 156 50182
rect 174 50179 246 50187
rect 256 50179 328 50187
rect 336 50181 342 50189
rect 400 50184 404 50189
rect 180 50151 185 50179
rect 174 50143 246 50151
rect 256 50143 328 50151
rect 332 50149 336 50179
rect 400 50150 438 50184
rect 224 50113 226 50129
rect 196 50105 226 50113
rect 196 50101 232 50105
rect 196 50071 204 50101
rect 216 50071 232 50101
rect 224 50024 226 50071
rect 300 50044 308 50113
rect 332 50111 342 50149
rect 400 50141 404 50150
rect 454 50135 504 50137
rect 494 50131 548 50135
rect 494 50126 514 50131
rect 504 50111 506 50126
rect 336 50099 342 50111
rect 289 50034 308 50044
rect 300 50028 308 50034
rect 332 50065 342 50099
rect 400 50103 404 50111
rect 400 50069 408 50103
rect 434 50069 438 50103
rect 498 50101 506 50111
rect 514 50101 515 50121
rect 504 50085 506 50101
rect 525 50092 528 50126
rect 547 50101 548 50121
rect 557 50101 564 50111
rect 514 50085 530 50091
rect 532 50085 548 50091
rect 332 50037 373 50065
rect 332 50031 351 50037
rect 107 49977 119 50011
rect 129 49977 149 50011
rect 196 49990 204 50024
rect 216 49990 232 50024
rect 244 50018 257 50024
rect 278 50018 291 50028
rect 244 49994 291 50018
rect 300 50018 321 50028
rect 336 50021 351 50031
rect 300 49994 329 50018
rect 332 50003 351 50021
rect 361 50031 375 50037
rect 400 50031 411 50069
rect 562 50032 612 50034
rect 361 50003 381 50031
rect 400 50003 409 50031
rect 466 50023 497 50031
rect 565 50023 596 50031
rect 442 50016 500 50023
rect 466 50015 500 50016
rect 565 50015 599 50023
rect 244 49990 257 49994
rect 42 49911 46 49945
rect 72 49911 76 49945
rect 42 49864 76 49868
rect 42 49849 46 49864
rect 72 49849 76 49864
rect 38 49831 80 49849
rect 16 49825 102 49831
rect 144 49825 148 49977
rect 174 49953 181 49981
rect 224 49943 226 49990
rect 300 49981 308 49994
rect 278 49970 305 49981
rect 332 49953 342 50003
rect 400 49983 404 50003
rect 497 49999 500 50015
rect 596 49999 599 50015
rect 466 49998 500 49999
rect 442 49991 500 49998
rect 565 49991 599 49999
rect 612 49982 614 50032
rect 256 49943 328 49951
rect 336 49945 342 49953
rect 400 49945 404 49953
rect 196 49913 204 49943
rect 216 49913 232 49943
rect 196 49909 232 49913
rect 196 49901 226 49909
rect 224 49885 226 49901
rect 332 49873 336 49941
rect 400 49911 408 49945
rect 434 49911 438 49945
rect 454 49929 504 49931
rect 504 49913 506 49929
rect 514 49923 530 49929
rect 532 49923 548 49929
rect 525 49913 548 49922
rect 400 49903 404 49911
rect 498 49903 506 49913
rect 504 49879 506 49903
rect 514 49893 515 49913
rect 525 49888 528 49913
rect 547 49893 548 49913
rect 557 49903 564 49913
rect 514 49879 548 49883
rect 400 49873 442 49874
rect 174 49863 246 49871
rect 400 49866 404 49873
rect 295 49832 300 49866
rect 324 49832 329 49866
rect 367 49849 438 49866
rect 367 49832 442 49849
rect 400 49831 442 49832
rect 378 49825 464 49831
rect 38 49809 80 49825
rect 400 49809 442 49825
rect -25 49795 25 49797
rect 42 49795 76 49809
rect 404 49795 438 49809
rect 455 49795 505 49797
rect 557 49795 607 49797
rect 16 49787 102 49795
rect 378 49787 464 49795
rect 8 49753 17 49787
rect 18 49785 51 49787
rect 80 49785 100 49787
rect 18 49753 100 49785
rect 380 49785 404 49787
rect 429 49785 438 49787
rect 442 49785 462 49787
rect 16 49745 102 49753
rect 42 49729 76 49745
rect 16 49709 38 49715
rect 42 49706 76 49710
rect 80 49709 102 49715
rect 42 49676 46 49706
rect 72 49676 76 49706
rect 42 49595 46 49629
rect 72 49595 76 49629
rect -25 49558 25 49560
rect -8 49550 14 49557
rect -8 49549 17 49550
rect 25 49549 27 49558
rect -12 49542 38 49549
rect -12 49541 34 49542
rect -12 49537 8 49541
rect 0 49525 8 49537
rect 14 49525 34 49541
rect 0 49524 34 49525
rect 0 49517 38 49524
rect 14 49516 17 49517
rect 25 49508 27 49517
rect 42 49488 45 49578
rect 69 49563 80 49595
rect 107 49563 143 49591
rect 144 49563 148 49783
rect 332 49715 336 49783
rect 380 49753 462 49785
rect 463 49753 472 49787
rect 480 49753 497 49787
rect 378 49745 464 49753
rect 505 49745 507 49795
rect 514 49753 548 49787
rect 565 49753 582 49787
rect 607 49745 609 49795
rect 404 49729 438 49745
rect 400 49715 442 49716
rect 378 49709 404 49715
rect 442 49709 464 49715
rect 400 49708 404 49709
rect 174 49669 246 49677
rect 295 49674 300 49708
rect 324 49674 329 49708
rect 224 49639 226 49655
rect 196 49631 226 49639
rect 332 49637 336 49705
rect 367 49674 438 49708
rect 400 49667 404 49674
rect 454 49661 504 49663
rect 494 49657 548 49661
rect 494 49652 514 49657
rect 504 49637 506 49652
rect 196 49627 232 49631
rect 196 49597 204 49627
rect 216 49597 232 49627
rect 400 49629 404 49637
rect 107 49557 119 49563
rect 109 49529 119 49557
rect 129 49529 149 49563
rect 174 49559 181 49589
rect 224 49550 226 49597
rect 256 49589 328 49597
rect 332 49595 336 49625
rect 400 49595 408 49629
rect 434 49595 438 49629
rect 498 49627 506 49637
rect 514 49627 515 49647
rect 504 49611 506 49627
rect 525 49618 528 49652
rect 547 49627 548 49647
rect 557 49627 564 49637
rect 514 49611 530 49617
rect 532 49611 548 49617
rect 278 49559 305 49570
rect 42 49437 46 49471
rect 72 49437 76 49471
rect 38 49399 80 49400
rect 42 49358 76 49392
rect 79 49358 113 49392
rect 42 49279 46 49313
rect 72 49279 76 49313
rect -25 49242 25 49244
rect -8 49234 14 49241
rect -8 49233 17 49234
rect 25 49233 27 49242
rect -12 49226 38 49233
rect -12 49225 34 49226
rect -12 49221 8 49225
rect 0 49209 8 49221
rect 14 49209 34 49225
rect 0 49208 34 49209
rect 0 49201 38 49208
rect 14 49200 17 49201
rect 25 49192 27 49201
rect 42 49172 45 49262
rect 71 49231 80 49259
rect 69 49193 80 49231
rect 144 49221 148 49529
rect 196 49516 204 49550
rect 216 49516 232 49550
rect 244 49546 257 49550
rect 300 49546 308 49559
rect 332 49557 342 49595
rect 400 49587 404 49595
rect 336 49547 342 49557
rect 244 49522 291 49546
rect 244 49516 257 49522
rect 224 49469 226 49516
rect 278 49512 291 49522
rect 300 49522 329 49546
rect 332 49537 342 49547
rect 400 49547 409 49575
rect 562 49558 612 49560
rect 466 49549 497 49557
rect 565 49549 596 49557
rect 300 49512 321 49522
rect 300 49506 308 49512
rect 289 49496 308 49506
rect 196 49439 204 49469
rect 216 49439 232 49469
rect 196 49435 232 49439
rect 196 49427 226 49435
rect 300 49427 308 49496
rect 332 49503 351 49537
rect 361 49509 381 49537
rect 361 49503 375 49509
rect 400 49503 411 49547
rect 442 49542 500 49549
rect 466 49541 500 49542
rect 565 49541 599 49549
rect 497 49525 500 49541
rect 596 49525 599 49541
rect 466 49524 500 49525
rect 442 49517 500 49524
rect 565 49517 599 49525
rect 612 49508 614 49558
rect 332 49479 342 49503
rect 336 49467 342 49479
rect 224 49411 226 49427
rect 332 49399 342 49467
rect 400 49471 404 49479
rect 400 49437 408 49471
rect 434 49437 438 49471
rect 454 49455 504 49457
rect 504 49439 506 49455
rect 514 49449 530 49455
rect 532 49449 548 49455
rect 525 49439 548 49448
rect 400 49429 404 49437
rect 498 49429 506 49439
rect 504 49405 506 49429
rect 514 49419 515 49439
rect 525 49414 528 49439
rect 547 49419 548 49439
rect 557 49429 564 49439
rect 514 49405 548 49409
rect 151 49358 156 49392
rect 174 49389 246 49397
rect 256 49389 328 49397
rect 336 49391 342 49399
rect 400 49394 404 49399
rect 180 49361 185 49389
rect 174 49353 246 49361
rect 256 49353 328 49361
rect 332 49359 336 49389
rect 400 49360 438 49394
rect 224 49323 226 49339
rect 196 49315 226 49323
rect 196 49311 232 49315
rect 196 49281 204 49311
rect 216 49281 232 49311
rect 224 49234 226 49281
rect 300 49254 308 49323
rect 332 49321 342 49359
rect 400 49351 404 49360
rect 454 49345 504 49347
rect 494 49341 548 49345
rect 494 49336 514 49341
rect 504 49321 506 49336
rect 336 49309 342 49321
rect 289 49244 308 49254
rect 300 49238 308 49244
rect 332 49275 342 49309
rect 400 49313 404 49321
rect 400 49279 408 49313
rect 434 49279 438 49313
rect 498 49311 506 49321
rect 514 49311 515 49331
rect 504 49295 506 49311
rect 525 49302 528 49336
rect 547 49311 548 49331
rect 557 49311 564 49321
rect 514 49295 530 49301
rect 532 49295 548 49301
rect 332 49247 373 49275
rect 332 49241 351 49247
rect 107 49187 119 49221
rect 129 49187 149 49221
rect 196 49200 204 49234
rect 216 49200 232 49234
rect 244 49228 257 49234
rect 278 49228 291 49238
rect 244 49204 291 49228
rect 300 49228 321 49238
rect 336 49231 351 49241
rect 300 49204 329 49228
rect 332 49213 351 49231
rect 361 49241 375 49247
rect 400 49241 411 49279
rect 562 49242 612 49244
rect 361 49213 381 49241
rect 400 49213 409 49241
rect 466 49233 497 49241
rect 565 49233 596 49241
rect 442 49226 500 49233
rect 466 49225 500 49226
rect 565 49225 599 49233
rect 244 49200 257 49204
rect 42 49121 46 49155
rect 72 49121 76 49155
rect 42 49074 76 49078
rect 42 49059 46 49074
rect 72 49059 76 49074
rect 38 49041 80 49059
rect 16 49035 102 49041
rect 144 49035 148 49187
rect 174 49163 181 49191
rect 224 49153 226 49200
rect 300 49191 308 49204
rect 278 49180 305 49191
rect 332 49163 342 49213
rect 400 49193 404 49213
rect 497 49209 500 49225
rect 596 49209 599 49225
rect 466 49208 500 49209
rect 442 49201 500 49208
rect 565 49201 599 49209
rect 612 49192 614 49242
rect 256 49153 328 49161
rect 336 49155 342 49163
rect 400 49155 404 49163
rect 196 49123 204 49153
rect 216 49123 232 49153
rect 196 49119 232 49123
rect 196 49111 226 49119
rect 224 49095 226 49111
rect 332 49083 336 49151
rect 400 49121 408 49155
rect 434 49121 438 49155
rect 454 49139 504 49141
rect 504 49123 506 49139
rect 514 49133 530 49139
rect 532 49133 548 49139
rect 525 49123 548 49132
rect 400 49113 404 49121
rect 498 49113 506 49123
rect 504 49089 506 49113
rect 514 49103 515 49123
rect 525 49098 528 49123
rect 547 49103 548 49123
rect 557 49113 564 49123
rect 514 49089 548 49093
rect 400 49083 442 49084
rect 174 49073 246 49081
rect 400 49076 404 49083
rect 295 49042 300 49076
rect 324 49042 329 49076
rect 367 49059 438 49076
rect 367 49042 442 49059
rect 400 49041 442 49042
rect 378 49035 464 49041
rect 38 49019 80 49035
rect 400 49019 442 49035
rect -25 49005 25 49007
rect 42 49005 76 49019
rect 404 49005 438 49019
rect 455 49005 505 49007
rect 557 49005 607 49007
rect 16 48997 102 49005
rect 378 48997 464 49005
rect 8 48963 17 48997
rect 18 48995 51 48997
rect 80 48995 100 48997
rect 18 48963 100 48995
rect 380 48995 404 48997
rect 429 48995 438 48997
rect 442 48995 462 48997
rect 16 48955 102 48963
rect 42 48939 76 48955
rect 16 48919 38 48925
rect 42 48916 76 48920
rect 80 48919 102 48925
rect 42 48886 46 48916
rect 72 48886 76 48916
rect 42 48805 46 48839
rect 72 48805 76 48839
rect -25 48768 25 48770
rect -8 48760 14 48767
rect -8 48759 17 48760
rect 25 48759 27 48768
rect -12 48752 38 48759
rect -12 48751 34 48752
rect -12 48747 8 48751
rect 0 48735 8 48747
rect 14 48735 34 48751
rect 0 48734 34 48735
rect 0 48727 38 48734
rect 14 48726 17 48727
rect 25 48718 27 48727
rect 42 48698 45 48788
rect 69 48773 80 48805
rect 107 48773 143 48801
rect 144 48773 148 48993
rect 332 48925 336 48993
rect 380 48963 462 48995
rect 463 48963 472 48997
rect 480 48963 497 48997
rect 378 48955 464 48963
rect 505 48955 507 49005
rect 514 48963 548 48997
rect 565 48963 582 48997
rect 607 48955 609 49005
rect 404 48939 438 48955
rect 400 48925 442 48926
rect 378 48919 404 48925
rect 442 48919 464 48925
rect 400 48918 404 48919
rect 174 48879 246 48887
rect 295 48884 300 48918
rect 324 48884 329 48918
rect 224 48849 226 48865
rect 196 48841 226 48849
rect 332 48847 336 48915
rect 367 48884 438 48918
rect 400 48877 404 48884
rect 454 48871 504 48873
rect 494 48867 548 48871
rect 494 48862 514 48867
rect 504 48847 506 48862
rect 196 48837 232 48841
rect 196 48807 204 48837
rect 216 48807 232 48837
rect 400 48839 404 48847
rect 107 48767 119 48773
rect 109 48739 119 48767
rect 129 48739 149 48773
rect 174 48769 181 48799
rect 224 48760 226 48807
rect 256 48799 328 48807
rect 332 48805 336 48835
rect 400 48805 408 48839
rect 434 48805 438 48839
rect 498 48837 506 48847
rect 514 48837 515 48857
rect 504 48821 506 48837
rect 525 48828 528 48862
rect 547 48837 548 48857
rect 557 48837 564 48847
rect 514 48821 530 48827
rect 532 48821 548 48827
rect 278 48769 305 48780
rect 42 48647 46 48681
rect 72 48647 76 48681
rect 38 48609 80 48610
rect 42 48568 76 48602
rect 79 48568 113 48602
rect 42 48489 46 48523
rect 72 48489 76 48523
rect -25 48452 25 48454
rect -8 48444 14 48451
rect -8 48443 17 48444
rect 25 48443 27 48452
rect -12 48436 38 48443
rect -12 48435 34 48436
rect -12 48431 8 48435
rect 0 48419 8 48431
rect 14 48419 34 48435
rect 0 48418 34 48419
rect 0 48411 38 48418
rect 14 48410 17 48411
rect 25 48402 27 48411
rect 42 48382 45 48472
rect 71 48441 80 48469
rect 69 48403 80 48441
rect 144 48431 148 48739
rect 196 48726 204 48760
rect 216 48726 232 48760
rect 244 48756 257 48760
rect 300 48756 308 48769
rect 332 48767 342 48805
rect 400 48797 404 48805
rect 336 48757 342 48767
rect 244 48732 291 48756
rect 244 48726 257 48732
rect 224 48679 226 48726
rect 278 48722 291 48732
rect 300 48732 329 48756
rect 332 48747 342 48757
rect 400 48757 409 48785
rect 562 48768 612 48770
rect 466 48759 497 48767
rect 565 48759 596 48767
rect 300 48722 321 48732
rect 300 48716 308 48722
rect 289 48706 308 48716
rect 196 48649 204 48679
rect 216 48649 232 48679
rect 196 48645 232 48649
rect 196 48637 226 48645
rect 300 48637 308 48706
rect 332 48713 351 48747
rect 361 48719 381 48747
rect 361 48713 375 48719
rect 400 48713 411 48757
rect 442 48752 500 48759
rect 466 48751 500 48752
rect 565 48751 599 48759
rect 497 48735 500 48751
rect 596 48735 599 48751
rect 466 48734 500 48735
rect 442 48727 500 48734
rect 565 48727 599 48735
rect 612 48718 614 48768
rect 332 48689 342 48713
rect 336 48677 342 48689
rect 224 48621 226 48637
rect 332 48609 342 48677
rect 400 48681 404 48689
rect 400 48647 408 48681
rect 434 48647 438 48681
rect 454 48665 504 48667
rect 504 48649 506 48665
rect 514 48659 530 48665
rect 532 48659 548 48665
rect 525 48649 548 48658
rect 400 48639 404 48647
rect 498 48639 506 48649
rect 504 48615 506 48639
rect 514 48629 515 48649
rect 525 48624 528 48649
rect 547 48629 548 48649
rect 557 48639 564 48649
rect 514 48615 548 48619
rect 151 48568 156 48602
rect 174 48599 246 48607
rect 256 48599 328 48607
rect 336 48601 342 48609
rect 400 48604 404 48609
rect 180 48571 185 48599
rect 174 48563 246 48571
rect 256 48563 328 48571
rect 332 48569 336 48599
rect 400 48570 438 48604
rect 224 48533 226 48549
rect 196 48525 226 48533
rect 196 48521 232 48525
rect 196 48491 204 48521
rect 216 48491 232 48521
rect 224 48444 226 48491
rect 300 48464 308 48533
rect 332 48531 342 48569
rect 400 48561 404 48570
rect 454 48555 504 48557
rect 494 48551 548 48555
rect 494 48546 514 48551
rect 504 48531 506 48546
rect 336 48519 342 48531
rect 289 48454 308 48464
rect 300 48448 308 48454
rect 332 48485 342 48519
rect 400 48523 404 48531
rect 400 48489 408 48523
rect 434 48489 438 48523
rect 498 48521 506 48531
rect 514 48521 515 48541
rect 504 48505 506 48521
rect 525 48512 528 48546
rect 547 48521 548 48541
rect 557 48521 564 48531
rect 514 48505 530 48511
rect 532 48505 548 48511
rect 332 48457 373 48485
rect 332 48451 351 48457
rect 107 48397 119 48431
rect 129 48397 149 48431
rect 196 48410 204 48444
rect 216 48410 232 48444
rect 244 48438 257 48444
rect 278 48438 291 48448
rect 244 48414 291 48438
rect 300 48438 321 48448
rect 336 48441 351 48451
rect 300 48414 329 48438
rect 332 48423 351 48441
rect 361 48451 375 48457
rect 400 48451 411 48489
rect 562 48452 612 48454
rect 361 48423 381 48451
rect 400 48423 409 48451
rect 466 48443 497 48451
rect 565 48443 596 48451
rect 442 48436 500 48443
rect 466 48435 500 48436
rect 565 48435 599 48443
rect 244 48410 257 48414
rect 42 48331 46 48365
rect 72 48331 76 48365
rect 42 48284 76 48288
rect 42 48269 46 48284
rect 72 48269 76 48284
rect 38 48251 80 48269
rect 16 48245 102 48251
rect 144 48245 148 48397
rect 174 48373 181 48401
rect 224 48363 226 48410
rect 300 48401 308 48414
rect 278 48390 305 48401
rect 332 48373 342 48423
rect 400 48403 404 48423
rect 497 48419 500 48435
rect 596 48419 599 48435
rect 466 48418 500 48419
rect 442 48411 500 48418
rect 565 48411 599 48419
rect 612 48402 614 48452
rect 256 48363 328 48371
rect 336 48365 342 48373
rect 400 48365 404 48373
rect 196 48333 204 48363
rect 216 48333 232 48363
rect 196 48329 232 48333
rect 196 48321 226 48329
rect 224 48305 226 48321
rect 332 48293 336 48361
rect 400 48331 408 48365
rect 434 48331 438 48365
rect 454 48349 504 48351
rect 504 48333 506 48349
rect 514 48343 530 48349
rect 532 48343 548 48349
rect 525 48333 548 48342
rect 400 48323 404 48331
rect 498 48323 506 48333
rect 504 48299 506 48323
rect 514 48313 515 48333
rect 525 48308 528 48333
rect 547 48313 548 48333
rect 557 48323 564 48333
rect 514 48299 548 48303
rect 400 48293 442 48294
rect 174 48283 246 48291
rect 400 48286 404 48293
rect 295 48252 300 48286
rect 324 48252 329 48286
rect 367 48269 438 48286
rect 367 48252 442 48269
rect 400 48251 442 48252
rect 378 48245 464 48251
rect 38 48229 80 48245
rect 400 48229 442 48245
rect -25 48215 25 48217
rect 42 48215 76 48229
rect 404 48215 438 48229
rect 455 48215 505 48217
rect 557 48215 607 48217
rect 16 48207 102 48215
rect 378 48207 464 48215
rect 8 48173 17 48207
rect 18 48205 51 48207
rect 80 48205 100 48207
rect 18 48173 100 48205
rect 380 48205 404 48207
rect 429 48205 438 48207
rect 442 48205 462 48207
rect 16 48165 102 48173
rect 42 48149 76 48165
rect 16 48129 38 48135
rect 42 48126 76 48130
rect 80 48129 102 48135
rect 42 48096 46 48126
rect 72 48096 76 48126
rect 42 48015 46 48049
rect 72 48015 76 48049
rect -25 47978 25 47980
rect -8 47970 14 47977
rect -8 47969 17 47970
rect 25 47969 27 47978
rect -12 47962 38 47969
rect -12 47961 34 47962
rect -12 47957 8 47961
rect 0 47945 8 47957
rect 14 47945 34 47961
rect 0 47944 34 47945
rect 0 47937 38 47944
rect 14 47936 17 47937
rect 25 47928 27 47937
rect 42 47908 45 47998
rect 69 47983 80 48015
rect 107 47983 143 48011
rect 144 47983 148 48203
rect 332 48135 336 48203
rect 380 48173 462 48205
rect 463 48173 472 48207
rect 480 48173 497 48207
rect 378 48165 464 48173
rect 505 48165 507 48215
rect 514 48173 548 48207
rect 565 48173 582 48207
rect 607 48165 609 48215
rect 404 48149 438 48165
rect 400 48135 442 48136
rect 378 48129 404 48135
rect 442 48129 464 48135
rect 400 48128 404 48129
rect 174 48089 246 48097
rect 295 48094 300 48128
rect 324 48094 329 48128
rect 224 48059 226 48075
rect 196 48051 226 48059
rect 332 48057 336 48125
rect 367 48094 438 48128
rect 400 48087 404 48094
rect 454 48081 504 48083
rect 494 48077 548 48081
rect 494 48072 514 48077
rect 504 48057 506 48072
rect 196 48047 232 48051
rect 196 48017 204 48047
rect 216 48017 232 48047
rect 400 48049 404 48057
rect 107 47977 119 47983
rect 109 47949 119 47977
rect 129 47949 149 47983
rect 174 47979 181 48009
rect 224 47970 226 48017
rect 256 48009 328 48017
rect 332 48015 336 48045
rect 400 48015 408 48049
rect 434 48015 438 48049
rect 498 48047 506 48057
rect 514 48047 515 48067
rect 504 48031 506 48047
rect 525 48038 528 48072
rect 547 48047 548 48067
rect 557 48047 564 48057
rect 514 48031 530 48037
rect 532 48031 548 48037
rect 278 47979 305 47990
rect 42 47857 46 47891
rect 72 47857 76 47891
rect 38 47819 80 47820
rect 42 47778 76 47812
rect 79 47778 113 47812
rect 42 47699 46 47733
rect 72 47699 76 47733
rect -25 47662 25 47664
rect -8 47654 14 47661
rect -8 47653 17 47654
rect 25 47653 27 47662
rect -12 47646 38 47653
rect -12 47645 34 47646
rect -12 47641 8 47645
rect 0 47629 8 47641
rect 14 47629 34 47645
rect 0 47628 34 47629
rect 0 47621 38 47628
rect 14 47620 17 47621
rect 25 47612 27 47621
rect 42 47592 45 47682
rect 71 47651 80 47679
rect 69 47613 80 47651
rect 144 47641 148 47949
rect 196 47936 204 47970
rect 216 47936 232 47970
rect 244 47966 257 47970
rect 300 47966 308 47979
rect 332 47977 342 48015
rect 400 48007 404 48015
rect 336 47967 342 47977
rect 244 47942 291 47966
rect 244 47936 257 47942
rect 224 47889 226 47936
rect 278 47932 291 47942
rect 300 47942 329 47966
rect 332 47957 342 47967
rect 400 47967 409 47995
rect 562 47978 612 47980
rect 466 47969 497 47977
rect 565 47969 596 47977
rect 300 47932 321 47942
rect 300 47926 308 47932
rect 289 47916 308 47926
rect 196 47859 204 47889
rect 216 47859 232 47889
rect 196 47855 232 47859
rect 196 47847 226 47855
rect 300 47847 308 47916
rect 332 47923 351 47957
rect 361 47929 381 47957
rect 361 47923 375 47929
rect 400 47923 411 47967
rect 442 47962 500 47969
rect 466 47961 500 47962
rect 565 47961 599 47969
rect 497 47945 500 47961
rect 596 47945 599 47961
rect 466 47944 500 47945
rect 442 47937 500 47944
rect 565 47937 599 47945
rect 612 47928 614 47978
rect 332 47899 342 47923
rect 336 47887 342 47899
rect 224 47831 226 47847
rect 332 47819 342 47887
rect 400 47891 404 47899
rect 400 47857 408 47891
rect 434 47857 438 47891
rect 454 47875 504 47877
rect 504 47859 506 47875
rect 514 47869 530 47875
rect 532 47869 548 47875
rect 525 47859 548 47868
rect 400 47849 404 47857
rect 498 47849 506 47859
rect 504 47825 506 47849
rect 514 47839 515 47859
rect 525 47834 528 47859
rect 547 47839 548 47859
rect 557 47849 564 47859
rect 514 47825 548 47829
rect 151 47778 156 47812
rect 174 47809 246 47817
rect 256 47809 328 47817
rect 336 47811 342 47819
rect 400 47814 404 47819
rect 180 47781 185 47809
rect 174 47773 246 47781
rect 256 47773 328 47781
rect 332 47779 336 47809
rect 400 47780 438 47814
rect 224 47743 226 47759
rect 196 47735 226 47743
rect 196 47731 232 47735
rect 196 47701 204 47731
rect 216 47701 232 47731
rect 224 47654 226 47701
rect 300 47674 308 47743
rect 332 47741 342 47779
rect 400 47771 404 47780
rect 454 47765 504 47767
rect 494 47761 548 47765
rect 494 47756 514 47761
rect 504 47741 506 47756
rect 336 47729 342 47741
rect 289 47664 308 47674
rect 300 47658 308 47664
rect 332 47695 342 47729
rect 400 47733 404 47741
rect 400 47699 408 47733
rect 434 47699 438 47733
rect 498 47731 506 47741
rect 514 47731 515 47751
rect 504 47715 506 47731
rect 525 47722 528 47756
rect 547 47731 548 47751
rect 557 47731 564 47741
rect 514 47715 530 47721
rect 532 47715 548 47721
rect 332 47667 373 47695
rect 332 47661 351 47667
rect 107 47607 119 47641
rect 129 47607 149 47641
rect 196 47620 204 47654
rect 216 47620 232 47654
rect 244 47648 257 47654
rect 278 47648 291 47658
rect 244 47624 291 47648
rect 300 47648 321 47658
rect 336 47651 351 47661
rect 300 47624 329 47648
rect 332 47633 351 47651
rect 361 47661 375 47667
rect 400 47661 411 47699
rect 562 47662 612 47664
rect 361 47633 381 47661
rect 400 47633 409 47661
rect 466 47653 497 47661
rect 565 47653 596 47661
rect 442 47646 500 47653
rect 466 47645 500 47646
rect 565 47645 599 47653
rect 244 47620 257 47624
rect 42 47541 46 47575
rect 72 47541 76 47575
rect 42 47494 76 47498
rect 42 47479 46 47494
rect 72 47479 76 47494
rect 38 47461 80 47479
rect 16 47455 102 47461
rect 144 47455 148 47607
rect 174 47583 181 47611
rect 224 47573 226 47620
rect 300 47611 308 47624
rect 278 47600 305 47611
rect 332 47583 342 47633
rect 400 47613 404 47633
rect 497 47629 500 47645
rect 596 47629 599 47645
rect 466 47628 500 47629
rect 442 47621 500 47628
rect 565 47621 599 47629
rect 612 47612 614 47662
rect 256 47573 328 47581
rect 336 47575 342 47583
rect 400 47575 404 47583
rect 196 47543 204 47573
rect 216 47543 232 47573
rect 196 47539 232 47543
rect 196 47531 226 47539
rect 224 47515 226 47531
rect 332 47503 336 47571
rect 400 47541 408 47575
rect 434 47541 438 47575
rect 454 47559 504 47561
rect 504 47543 506 47559
rect 514 47553 530 47559
rect 532 47553 548 47559
rect 525 47543 548 47552
rect 400 47533 404 47541
rect 498 47533 506 47543
rect 504 47509 506 47533
rect 514 47523 515 47543
rect 525 47518 528 47543
rect 547 47523 548 47543
rect 557 47533 564 47543
rect 514 47509 548 47513
rect 400 47503 442 47504
rect 174 47493 246 47501
rect 400 47496 404 47503
rect 295 47462 300 47496
rect 324 47462 329 47496
rect 367 47479 438 47496
rect 367 47462 442 47479
rect 400 47461 442 47462
rect 378 47455 464 47461
rect 38 47439 80 47455
rect 400 47439 442 47455
rect -25 47425 25 47427
rect 42 47425 76 47439
rect 404 47425 438 47439
rect 455 47425 505 47427
rect 557 47425 607 47427
rect 16 47417 102 47425
rect 378 47417 464 47425
rect 8 47383 17 47417
rect 18 47415 51 47417
rect 80 47415 100 47417
rect 18 47383 100 47415
rect 380 47415 404 47417
rect 429 47415 438 47417
rect 442 47415 462 47417
rect 16 47375 102 47383
rect 42 47359 76 47375
rect 16 47339 38 47345
rect 42 47336 76 47340
rect 80 47339 102 47345
rect 42 47306 46 47336
rect 72 47306 76 47336
rect 42 47225 46 47259
rect 72 47225 76 47259
rect -25 47188 25 47190
rect -8 47180 14 47187
rect -8 47179 17 47180
rect 25 47179 27 47188
rect -12 47172 38 47179
rect -12 47171 34 47172
rect -12 47167 8 47171
rect 0 47155 8 47167
rect 14 47155 34 47171
rect 0 47154 34 47155
rect 0 47147 38 47154
rect 14 47146 17 47147
rect 25 47138 27 47147
rect 42 47118 45 47208
rect 69 47193 80 47225
rect 107 47193 143 47221
rect 144 47193 148 47413
rect 332 47345 336 47413
rect 380 47383 462 47415
rect 463 47383 472 47417
rect 480 47383 497 47417
rect 378 47375 464 47383
rect 505 47375 507 47425
rect 514 47383 548 47417
rect 565 47383 582 47417
rect 607 47375 609 47425
rect 404 47359 438 47375
rect 400 47345 442 47346
rect 378 47339 404 47345
rect 442 47339 464 47345
rect 400 47338 404 47339
rect 174 47299 246 47307
rect 295 47304 300 47338
rect 324 47304 329 47338
rect 224 47269 226 47285
rect 196 47261 226 47269
rect 332 47267 336 47335
rect 367 47304 438 47338
rect 400 47297 404 47304
rect 454 47291 504 47293
rect 494 47287 548 47291
rect 494 47282 514 47287
rect 504 47267 506 47282
rect 196 47257 232 47261
rect 196 47227 204 47257
rect 216 47227 232 47257
rect 400 47259 404 47267
rect 107 47187 119 47193
rect 109 47159 119 47187
rect 129 47159 149 47193
rect 174 47189 181 47219
rect 224 47180 226 47227
rect 256 47219 328 47227
rect 332 47225 336 47255
rect 400 47225 408 47259
rect 434 47225 438 47259
rect 498 47257 506 47267
rect 514 47257 515 47277
rect 504 47241 506 47257
rect 525 47248 528 47282
rect 547 47257 548 47277
rect 557 47257 564 47267
rect 514 47241 530 47247
rect 532 47241 548 47247
rect 278 47189 305 47200
rect 42 47067 46 47101
rect 72 47067 76 47101
rect 38 47029 80 47030
rect 42 46988 76 47022
rect 79 46988 113 47022
rect 42 46909 46 46943
rect 72 46909 76 46943
rect -25 46872 25 46874
rect -8 46864 14 46871
rect -8 46863 17 46864
rect 25 46863 27 46872
rect -12 46856 38 46863
rect -12 46855 34 46856
rect -12 46851 8 46855
rect 0 46839 8 46851
rect 14 46839 34 46855
rect 0 46838 34 46839
rect 0 46831 38 46838
rect 14 46830 17 46831
rect 25 46822 27 46831
rect 42 46802 45 46892
rect 71 46861 80 46889
rect 69 46823 80 46861
rect 144 46851 148 47159
rect 196 47146 204 47180
rect 216 47146 232 47180
rect 244 47176 257 47180
rect 300 47176 308 47189
rect 332 47187 342 47225
rect 400 47217 404 47225
rect 336 47177 342 47187
rect 244 47152 291 47176
rect 244 47146 257 47152
rect 224 47099 226 47146
rect 278 47142 291 47152
rect 300 47152 329 47176
rect 332 47167 342 47177
rect 400 47177 409 47205
rect 562 47188 612 47190
rect 466 47179 497 47187
rect 565 47179 596 47187
rect 300 47142 321 47152
rect 300 47136 308 47142
rect 289 47126 308 47136
rect 196 47069 204 47099
rect 216 47069 232 47099
rect 196 47065 232 47069
rect 196 47057 226 47065
rect 300 47057 308 47126
rect 332 47133 351 47167
rect 361 47139 381 47167
rect 361 47133 375 47139
rect 400 47133 411 47177
rect 442 47172 500 47179
rect 466 47171 500 47172
rect 565 47171 599 47179
rect 497 47155 500 47171
rect 596 47155 599 47171
rect 466 47154 500 47155
rect 442 47147 500 47154
rect 565 47147 599 47155
rect 612 47138 614 47188
rect 332 47109 342 47133
rect 336 47097 342 47109
rect 224 47041 226 47057
rect 332 47029 342 47097
rect 400 47101 404 47109
rect 400 47067 408 47101
rect 434 47067 438 47101
rect 454 47085 504 47087
rect 504 47069 506 47085
rect 514 47079 530 47085
rect 532 47079 548 47085
rect 525 47069 548 47078
rect 400 47059 404 47067
rect 498 47059 506 47069
rect 504 47035 506 47059
rect 514 47049 515 47069
rect 525 47044 528 47069
rect 547 47049 548 47069
rect 557 47059 564 47069
rect 514 47035 548 47039
rect 151 46988 156 47022
rect 174 47019 246 47027
rect 256 47019 328 47027
rect 336 47021 342 47029
rect 400 47024 404 47029
rect 180 46991 185 47019
rect 174 46983 246 46991
rect 256 46983 328 46991
rect 332 46989 336 47019
rect 400 46990 438 47024
rect 224 46953 226 46969
rect 196 46945 226 46953
rect 196 46941 232 46945
rect 196 46911 204 46941
rect 216 46911 232 46941
rect 224 46864 226 46911
rect 300 46884 308 46953
rect 332 46951 342 46989
rect 400 46981 404 46990
rect 454 46975 504 46977
rect 494 46971 548 46975
rect 494 46966 514 46971
rect 504 46951 506 46966
rect 336 46939 342 46951
rect 289 46874 308 46884
rect 300 46868 308 46874
rect 332 46905 342 46939
rect 400 46943 404 46951
rect 400 46909 408 46943
rect 434 46909 438 46943
rect 498 46941 506 46951
rect 514 46941 515 46961
rect 504 46925 506 46941
rect 525 46932 528 46966
rect 547 46941 548 46961
rect 557 46941 564 46951
rect 514 46925 530 46931
rect 532 46925 548 46931
rect 332 46877 373 46905
rect 332 46871 351 46877
rect 107 46817 119 46851
rect 129 46817 149 46851
rect 196 46830 204 46864
rect 216 46830 232 46864
rect 244 46858 257 46864
rect 278 46858 291 46868
rect 244 46834 291 46858
rect 300 46858 321 46868
rect 336 46861 351 46871
rect 300 46834 329 46858
rect 332 46843 351 46861
rect 361 46871 375 46877
rect 400 46871 411 46909
rect 562 46872 612 46874
rect 361 46843 381 46871
rect 400 46843 409 46871
rect 466 46863 497 46871
rect 565 46863 596 46871
rect 442 46856 500 46863
rect 466 46855 500 46856
rect 565 46855 599 46863
rect 244 46830 257 46834
rect 42 46751 46 46785
rect 72 46751 76 46785
rect 42 46704 76 46708
rect 42 46689 46 46704
rect 72 46689 76 46704
rect 38 46671 80 46689
rect 16 46665 102 46671
rect 144 46665 148 46817
rect 174 46793 181 46821
rect 224 46783 226 46830
rect 300 46821 308 46834
rect 278 46810 305 46821
rect 332 46793 342 46843
rect 400 46823 404 46843
rect 497 46839 500 46855
rect 596 46839 599 46855
rect 466 46838 500 46839
rect 442 46831 500 46838
rect 565 46831 599 46839
rect 612 46822 614 46872
rect 256 46783 328 46791
rect 336 46785 342 46793
rect 400 46785 404 46793
rect 196 46753 204 46783
rect 216 46753 232 46783
rect 196 46749 232 46753
rect 196 46741 226 46749
rect 224 46725 226 46741
rect 332 46713 336 46781
rect 400 46751 408 46785
rect 434 46751 438 46785
rect 454 46769 504 46771
rect 504 46753 506 46769
rect 514 46763 530 46769
rect 532 46763 548 46769
rect 525 46753 548 46762
rect 400 46743 404 46751
rect 498 46743 506 46753
rect 504 46719 506 46743
rect 514 46733 515 46753
rect 525 46728 528 46753
rect 547 46733 548 46753
rect 557 46743 564 46753
rect 514 46719 548 46723
rect 400 46713 442 46714
rect 174 46703 246 46711
rect 400 46706 404 46713
rect 295 46672 300 46706
rect 324 46672 329 46706
rect 367 46689 438 46706
rect 367 46672 442 46689
rect 400 46671 442 46672
rect 378 46665 464 46671
rect 38 46649 80 46665
rect 400 46649 442 46665
rect -25 46635 25 46637
rect 42 46635 76 46649
rect 404 46635 438 46649
rect 455 46635 505 46637
rect 557 46635 607 46637
rect 16 46627 102 46635
rect 378 46627 464 46635
rect 8 46593 17 46627
rect 18 46625 51 46627
rect 80 46625 100 46627
rect 18 46593 100 46625
rect 380 46625 404 46627
rect 429 46625 438 46627
rect 442 46625 462 46627
rect 16 46585 102 46593
rect 42 46569 76 46585
rect 16 46549 38 46555
rect 42 46546 76 46550
rect 80 46549 102 46555
rect 42 46516 46 46546
rect 72 46516 76 46546
rect 42 46435 46 46469
rect 72 46435 76 46469
rect -25 46398 25 46400
rect -8 46390 14 46397
rect -8 46389 17 46390
rect 25 46389 27 46398
rect -12 46382 38 46389
rect -12 46381 34 46382
rect -12 46377 8 46381
rect 0 46365 8 46377
rect 14 46365 34 46381
rect 0 46364 34 46365
rect 0 46357 38 46364
rect 14 46356 17 46357
rect 25 46348 27 46357
rect 42 46328 45 46418
rect 69 46403 80 46435
rect 107 46403 143 46431
rect 144 46403 148 46623
rect 332 46555 336 46623
rect 380 46593 462 46625
rect 463 46593 472 46627
rect 480 46593 497 46627
rect 378 46585 464 46593
rect 505 46585 507 46635
rect 514 46593 548 46627
rect 565 46593 582 46627
rect 607 46585 609 46635
rect 404 46569 438 46585
rect 400 46555 442 46556
rect 378 46549 404 46555
rect 442 46549 464 46555
rect 400 46548 404 46549
rect 174 46509 246 46517
rect 295 46514 300 46548
rect 324 46514 329 46548
rect 224 46479 226 46495
rect 196 46471 226 46479
rect 332 46477 336 46545
rect 367 46514 438 46548
rect 400 46507 404 46514
rect 454 46501 504 46503
rect 494 46497 548 46501
rect 494 46492 514 46497
rect 504 46477 506 46492
rect 196 46467 232 46471
rect 196 46437 204 46467
rect 216 46437 232 46467
rect 400 46469 404 46477
rect 107 46397 119 46403
rect 109 46369 119 46397
rect 129 46369 149 46403
rect 174 46399 181 46429
rect 224 46390 226 46437
rect 256 46429 328 46437
rect 332 46435 336 46465
rect 400 46435 408 46469
rect 434 46435 438 46469
rect 498 46467 506 46477
rect 514 46467 515 46487
rect 504 46451 506 46467
rect 525 46458 528 46492
rect 547 46467 548 46487
rect 557 46467 564 46477
rect 514 46451 530 46457
rect 532 46451 548 46457
rect 278 46399 305 46410
rect 42 46277 46 46311
rect 72 46277 76 46311
rect 38 46239 80 46240
rect 42 46198 76 46232
rect 79 46198 113 46232
rect 42 46119 46 46153
rect 72 46119 76 46153
rect -25 46082 25 46084
rect -8 46074 14 46081
rect -8 46073 17 46074
rect 25 46073 27 46082
rect -12 46066 38 46073
rect -12 46065 34 46066
rect -12 46061 8 46065
rect 0 46049 8 46061
rect 14 46049 34 46065
rect 0 46048 34 46049
rect 0 46041 38 46048
rect 14 46040 17 46041
rect 25 46032 27 46041
rect 42 46012 45 46102
rect 71 46071 80 46099
rect 69 46033 80 46071
rect 144 46061 148 46369
rect 196 46356 204 46390
rect 216 46356 232 46390
rect 244 46386 257 46390
rect 300 46386 308 46399
rect 332 46397 342 46435
rect 400 46427 404 46435
rect 336 46387 342 46397
rect 244 46362 291 46386
rect 244 46356 257 46362
rect 224 46309 226 46356
rect 278 46352 291 46362
rect 300 46362 329 46386
rect 332 46377 342 46387
rect 400 46387 409 46415
rect 562 46398 612 46400
rect 466 46389 497 46397
rect 565 46389 596 46397
rect 300 46352 321 46362
rect 300 46346 308 46352
rect 289 46336 308 46346
rect 196 46279 204 46309
rect 216 46279 232 46309
rect 196 46275 232 46279
rect 196 46267 226 46275
rect 300 46267 308 46336
rect 332 46343 351 46377
rect 361 46349 381 46377
rect 361 46343 375 46349
rect 400 46343 411 46387
rect 442 46382 500 46389
rect 466 46381 500 46382
rect 565 46381 599 46389
rect 497 46365 500 46381
rect 596 46365 599 46381
rect 466 46364 500 46365
rect 442 46357 500 46364
rect 565 46357 599 46365
rect 612 46348 614 46398
rect 332 46319 342 46343
rect 336 46307 342 46319
rect 224 46251 226 46267
rect 332 46239 342 46307
rect 400 46311 404 46319
rect 400 46277 408 46311
rect 434 46277 438 46311
rect 454 46295 504 46297
rect 504 46279 506 46295
rect 514 46289 530 46295
rect 532 46289 548 46295
rect 525 46279 548 46288
rect 400 46269 404 46277
rect 498 46269 506 46279
rect 504 46245 506 46269
rect 514 46259 515 46279
rect 525 46254 528 46279
rect 547 46259 548 46279
rect 557 46269 564 46279
rect 514 46245 548 46249
rect 151 46198 156 46232
rect 174 46229 246 46237
rect 256 46229 328 46237
rect 336 46231 342 46239
rect 400 46234 404 46239
rect 180 46201 185 46229
rect 174 46193 246 46201
rect 256 46193 328 46201
rect 332 46199 336 46229
rect 400 46200 438 46234
rect 224 46163 226 46179
rect 196 46155 226 46163
rect 196 46151 232 46155
rect 196 46121 204 46151
rect 216 46121 232 46151
rect 224 46074 226 46121
rect 300 46094 308 46163
rect 332 46161 342 46199
rect 400 46191 404 46200
rect 454 46185 504 46187
rect 494 46181 548 46185
rect 494 46176 514 46181
rect 504 46161 506 46176
rect 336 46149 342 46161
rect 289 46084 308 46094
rect 300 46078 308 46084
rect 332 46115 342 46149
rect 400 46153 404 46161
rect 400 46119 408 46153
rect 434 46119 438 46153
rect 498 46151 506 46161
rect 514 46151 515 46171
rect 504 46135 506 46151
rect 525 46142 528 46176
rect 547 46151 548 46171
rect 557 46151 564 46161
rect 514 46135 530 46141
rect 532 46135 548 46141
rect 332 46087 373 46115
rect 332 46081 351 46087
rect 107 46027 119 46061
rect 129 46027 149 46061
rect 196 46040 204 46074
rect 216 46040 232 46074
rect 244 46068 257 46074
rect 278 46068 291 46078
rect 244 46044 291 46068
rect 300 46068 321 46078
rect 336 46071 351 46081
rect 300 46044 329 46068
rect 332 46053 351 46071
rect 361 46081 375 46087
rect 400 46081 411 46119
rect 562 46082 612 46084
rect 361 46053 381 46081
rect 400 46053 409 46081
rect 466 46073 497 46081
rect 565 46073 596 46081
rect 442 46066 500 46073
rect 466 46065 500 46066
rect 565 46065 599 46073
rect 244 46040 257 46044
rect 42 45961 46 45995
rect 72 45961 76 45995
rect 42 45914 76 45918
rect 42 45899 46 45914
rect 72 45899 76 45914
rect 38 45881 80 45899
rect 16 45875 102 45881
rect 144 45875 148 46027
rect 174 46003 181 46031
rect 224 45993 226 46040
rect 300 46031 308 46044
rect 278 46020 305 46031
rect 332 46003 342 46053
rect 400 46033 404 46053
rect 497 46049 500 46065
rect 596 46049 599 46065
rect 466 46048 500 46049
rect 442 46041 500 46048
rect 565 46041 599 46049
rect 612 46032 614 46082
rect 256 45993 328 46001
rect 336 45995 342 46003
rect 400 45995 404 46003
rect 196 45963 204 45993
rect 216 45963 232 45993
rect 196 45959 232 45963
rect 196 45951 226 45959
rect 224 45935 226 45951
rect 332 45923 336 45991
rect 400 45961 408 45995
rect 434 45961 438 45995
rect 454 45979 504 45981
rect 504 45963 506 45979
rect 514 45973 530 45979
rect 532 45973 548 45979
rect 525 45963 548 45972
rect 400 45953 404 45961
rect 498 45953 506 45963
rect 504 45929 506 45953
rect 514 45943 515 45963
rect 525 45938 528 45963
rect 547 45943 548 45963
rect 557 45953 564 45963
rect 514 45929 548 45933
rect 400 45923 442 45924
rect 174 45913 246 45921
rect 400 45916 404 45923
rect 295 45882 300 45916
rect 324 45882 329 45916
rect 367 45899 438 45916
rect 367 45882 442 45899
rect 400 45881 442 45882
rect 378 45875 464 45881
rect 38 45859 80 45875
rect 400 45859 442 45875
rect -25 45845 25 45847
rect 42 45845 76 45859
rect 404 45845 438 45859
rect 455 45845 505 45847
rect 557 45845 607 45847
rect 16 45837 102 45845
rect 378 45837 464 45845
rect 8 45803 17 45837
rect 18 45835 51 45837
rect 80 45835 100 45837
rect 18 45803 100 45835
rect 380 45835 404 45837
rect 429 45835 438 45837
rect 442 45835 462 45837
rect 16 45795 102 45803
rect 42 45779 76 45795
rect 16 45759 38 45765
rect 42 45756 76 45760
rect 80 45759 102 45765
rect 42 45726 46 45756
rect 72 45726 76 45756
rect 42 45645 46 45679
rect 72 45645 76 45679
rect -25 45608 25 45610
rect -8 45600 14 45607
rect -8 45599 17 45600
rect 25 45599 27 45608
rect -12 45592 38 45599
rect -12 45591 34 45592
rect -12 45587 8 45591
rect 0 45575 8 45587
rect 14 45575 34 45591
rect 0 45574 34 45575
rect 0 45567 38 45574
rect 14 45566 17 45567
rect 25 45558 27 45567
rect 42 45538 45 45628
rect 69 45613 80 45645
rect 107 45613 143 45641
rect 144 45613 148 45833
rect 332 45765 336 45833
rect 380 45803 462 45835
rect 463 45803 472 45837
rect 480 45803 497 45837
rect 378 45795 464 45803
rect 505 45795 507 45845
rect 514 45803 548 45837
rect 565 45803 582 45837
rect 607 45795 609 45845
rect 404 45779 438 45795
rect 400 45765 442 45766
rect 378 45759 404 45765
rect 442 45759 464 45765
rect 400 45758 404 45759
rect 174 45719 246 45727
rect 295 45724 300 45758
rect 324 45724 329 45758
rect 224 45689 226 45705
rect 196 45681 226 45689
rect 332 45687 336 45755
rect 367 45724 438 45758
rect 400 45717 404 45724
rect 454 45711 504 45713
rect 494 45707 548 45711
rect 494 45702 514 45707
rect 504 45687 506 45702
rect 196 45677 232 45681
rect 196 45647 204 45677
rect 216 45647 232 45677
rect 400 45679 404 45687
rect 107 45607 119 45613
rect 109 45579 119 45607
rect 129 45579 149 45613
rect 174 45609 181 45639
rect 224 45600 226 45647
rect 256 45639 328 45647
rect 332 45645 336 45675
rect 400 45645 408 45679
rect 434 45645 438 45679
rect 498 45677 506 45687
rect 514 45677 515 45697
rect 504 45661 506 45677
rect 525 45668 528 45702
rect 547 45677 548 45697
rect 557 45677 564 45687
rect 514 45661 530 45667
rect 532 45661 548 45667
rect 278 45609 305 45620
rect 42 45487 46 45521
rect 72 45487 76 45521
rect 38 45449 80 45450
rect 42 45408 76 45442
rect 79 45408 113 45442
rect 42 45329 46 45363
rect 72 45329 76 45363
rect -25 45292 25 45294
rect -8 45284 14 45291
rect -8 45283 17 45284
rect 25 45283 27 45292
rect -12 45276 38 45283
rect -12 45275 34 45276
rect -12 45271 8 45275
rect 0 45259 8 45271
rect 14 45259 34 45275
rect 0 45258 34 45259
rect 0 45251 38 45258
rect 14 45250 17 45251
rect 25 45242 27 45251
rect 42 45222 45 45312
rect 71 45281 80 45309
rect 69 45243 80 45281
rect 144 45271 148 45579
rect 196 45566 204 45600
rect 216 45566 232 45600
rect 244 45596 257 45600
rect 300 45596 308 45609
rect 332 45607 342 45645
rect 400 45637 404 45645
rect 336 45597 342 45607
rect 244 45572 291 45596
rect 244 45566 257 45572
rect 224 45519 226 45566
rect 278 45562 291 45572
rect 300 45572 329 45596
rect 332 45587 342 45597
rect 400 45597 409 45625
rect 562 45608 612 45610
rect 466 45599 497 45607
rect 565 45599 596 45607
rect 300 45562 321 45572
rect 300 45556 308 45562
rect 289 45546 308 45556
rect 196 45489 204 45519
rect 216 45489 232 45519
rect 196 45485 232 45489
rect 196 45477 226 45485
rect 300 45477 308 45546
rect 332 45553 351 45587
rect 361 45559 381 45587
rect 361 45553 375 45559
rect 400 45553 411 45597
rect 442 45592 500 45599
rect 466 45591 500 45592
rect 565 45591 599 45599
rect 497 45575 500 45591
rect 596 45575 599 45591
rect 466 45574 500 45575
rect 442 45567 500 45574
rect 565 45567 599 45575
rect 612 45558 614 45608
rect 332 45529 342 45553
rect 336 45517 342 45529
rect 224 45461 226 45477
rect 332 45449 342 45517
rect 400 45521 404 45529
rect 400 45487 408 45521
rect 434 45487 438 45521
rect 454 45505 504 45507
rect 504 45489 506 45505
rect 514 45499 530 45505
rect 532 45499 548 45505
rect 525 45489 548 45498
rect 400 45479 404 45487
rect 498 45479 506 45489
rect 504 45455 506 45479
rect 514 45469 515 45489
rect 525 45464 528 45489
rect 547 45469 548 45489
rect 557 45479 564 45489
rect 514 45455 548 45459
rect 151 45408 156 45442
rect 174 45439 246 45447
rect 256 45439 328 45447
rect 336 45441 342 45449
rect 400 45444 404 45449
rect 180 45411 185 45439
rect 174 45403 246 45411
rect 256 45403 328 45411
rect 332 45409 336 45439
rect 400 45410 438 45444
rect 224 45373 226 45389
rect 196 45365 226 45373
rect 196 45361 232 45365
rect 196 45331 204 45361
rect 216 45331 232 45361
rect 224 45284 226 45331
rect 300 45304 308 45373
rect 332 45371 342 45409
rect 400 45401 404 45410
rect 454 45395 504 45397
rect 494 45391 548 45395
rect 494 45386 514 45391
rect 504 45371 506 45386
rect 336 45359 342 45371
rect 289 45294 308 45304
rect 300 45288 308 45294
rect 332 45325 342 45359
rect 400 45363 404 45371
rect 400 45329 408 45363
rect 434 45329 438 45363
rect 498 45361 506 45371
rect 514 45361 515 45381
rect 504 45345 506 45361
rect 525 45352 528 45386
rect 547 45361 548 45381
rect 557 45361 564 45371
rect 514 45345 530 45351
rect 532 45345 548 45351
rect 332 45297 373 45325
rect 332 45291 351 45297
rect 107 45237 119 45271
rect 129 45237 149 45271
rect 196 45250 204 45284
rect 216 45250 232 45284
rect 244 45278 257 45284
rect 278 45278 291 45288
rect 244 45254 291 45278
rect 300 45278 321 45288
rect 336 45281 351 45291
rect 300 45254 329 45278
rect 332 45263 351 45281
rect 361 45291 375 45297
rect 400 45291 411 45329
rect 562 45292 612 45294
rect 361 45263 381 45291
rect 400 45263 409 45291
rect 466 45283 497 45291
rect 565 45283 596 45291
rect 442 45276 500 45283
rect 466 45275 500 45276
rect 565 45275 599 45283
rect 244 45250 257 45254
rect 42 45171 46 45205
rect 72 45171 76 45205
rect 42 45124 76 45128
rect 42 45109 46 45124
rect 72 45109 76 45124
rect 38 45091 80 45109
rect 16 45085 102 45091
rect 144 45085 148 45237
rect 174 45213 181 45241
rect 224 45203 226 45250
rect 300 45241 308 45254
rect 278 45230 305 45241
rect 332 45213 342 45263
rect 400 45243 404 45263
rect 497 45259 500 45275
rect 596 45259 599 45275
rect 466 45258 500 45259
rect 442 45251 500 45258
rect 565 45251 599 45259
rect 612 45242 614 45292
rect 256 45203 328 45211
rect 336 45205 342 45213
rect 400 45205 404 45213
rect 196 45173 204 45203
rect 216 45173 232 45203
rect 196 45169 232 45173
rect 196 45161 226 45169
rect 224 45145 226 45161
rect 332 45133 336 45201
rect 400 45171 408 45205
rect 434 45171 438 45205
rect 454 45189 504 45191
rect 504 45173 506 45189
rect 514 45183 530 45189
rect 532 45183 548 45189
rect 525 45173 548 45182
rect 400 45163 404 45171
rect 498 45163 506 45173
rect 504 45139 506 45163
rect 514 45153 515 45173
rect 525 45148 528 45173
rect 547 45153 548 45173
rect 557 45163 564 45173
rect 514 45139 548 45143
rect 400 45133 442 45134
rect 174 45123 246 45131
rect 400 45126 404 45133
rect 295 45092 300 45126
rect 324 45092 329 45126
rect 367 45109 438 45126
rect 367 45092 442 45109
rect 400 45091 442 45092
rect 378 45085 464 45091
rect 38 45069 80 45085
rect 400 45069 442 45085
rect -25 45055 25 45057
rect 42 45055 76 45069
rect 404 45055 438 45069
rect 455 45055 505 45057
rect 557 45055 607 45057
rect 16 45047 102 45055
rect 378 45047 464 45055
rect 8 45013 17 45047
rect 18 45045 51 45047
rect 80 45045 100 45047
rect 18 45013 100 45045
rect 380 45045 404 45047
rect 429 45045 438 45047
rect 442 45045 462 45047
rect 16 45005 102 45013
rect 42 44989 76 45005
rect 16 44969 38 44975
rect 42 44966 76 44970
rect 80 44969 102 44975
rect 42 44936 46 44966
rect 72 44936 76 44966
rect 42 44855 46 44889
rect 72 44855 76 44889
rect -25 44818 25 44820
rect -8 44810 14 44817
rect -8 44809 17 44810
rect 25 44809 27 44818
rect -12 44802 38 44809
rect -12 44801 34 44802
rect -12 44797 8 44801
rect 0 44785 8 44797
rect 14 44785 34 44801
rect 0 44784 34 44785
rect 0 44777 38 44784
rect 14 44776 17 44777
rect 25 44768 27 44777
rect 42 44748 45 44838
rect 69 44823 80 44855
rect 107 44823 143 44851
rect 144 44823 148 45043
rect 332 44975 336 45043
rect 380 45013 462 45045
rect 463 45013 472 45047
rect 480 45013 497 45047
rect 378 45005 464 45013
rect 505 45005 507 45055
rect 514 45013 548 45047
rect 565 45013 582 45047
rect 607 45005 609 45055
rect 404 44989 438 45005
rect 400 44975 442 44976
rect 378 44969 404 44975
rect 442 44969 464 44975
rect 400 44968 404 44969
rect 174 44929 246 44937
rect 295 44934 300 44968
rect 324 44934 329 44968
rect 224 44899 226 44915
rect 196 44891 226 44899
rect 332 44897 336 44965
rect 367 44934 438 44968
rect 400 44927 404 44934
rect 454 44921 504 44923
rect 494 44917 548 44921
rect 494 44912 514 44917
rect 504 44897 506 44912
rect 196 44887 232 44891
rect 196 44857 204 44887
rect 216 44857 232 44887
rect 400 44889 404 44897
rect 107 44817 119 44823
rect 109 44789 119 44817
rect 129 44789 149 44823
rect 174 44819 181 44849
rect 224 44810 226 44857
rect 256 44849 328 44857
rect 332 44855 336 44885
rect 400 44855 408 44889
rect 434 44855 438 44889
rect 498 44887 506 44897
rect 514 44887 515 44907
rect 504 44871 506 44887
rect 525 44878 528 44912
rect 547 44887 548 44907
rect 557 44887 564 44897
rect 514 44871 530 44877
rect 532 44871 548 44877
rect 278 44819 305 44830
rect 42 44697 46 44731
rect 72 44697 76 44731
rect 38 44659 80 44660
rect 42 44618 76 44652
rect 79 44618 113 44652
rect 42 44539 46 44573
rect 72 44539 76 44573
rect -25 44502 25 44504
rect -8 44494 14 44501
rect -8 44493 17 44494
rect 25 44493 27 44502
rect -12 44486 38 44493
rect -12 44485 34 44486
rect -12 44481 8 44485
rect 0 44469 8 44481
rect 14 44469 34 44485
rect 0 44468 34 44469
rect 0 44461 38 44468
rect 14 44460 17 44461
rect 25 44452 27 44461
rect 42 44432 45 44522
rect 71 44491 80 44519
rect 69 44453 80 44491
rect 144 44481 148 44789
rect 196 44776 204 44810
rect 216 44776 232 44810
rect 244 44806 257 44810
rect 300 44806 308 44819
rect 332 44817 342 44855
rect 400 44847 404 44855
rect 336 44807 342 44817
rect 244 44782 291 44806
rect 244 44776 257 44782
rect 224 44729 226 44776
rect 278 44772 291 44782
rect 300 44782 329 44806
rect 332 44797 342 44807
rect 400 44807 409 44835
rect 562 44818 612 44820
rect 466 44809 497 44817
rect 565 44809 596 44817
rect 300 44772 321 44782
rect 300 44766 308 44772
rect 289 44756 308 44766
rect 196 44699 204 44729
rect 216 44699 232 44729
rect 196 44695 232 44699
rect 196 44687 226 44695
rect 300 44687 308 44756
rect 332 44763 351 44797
rect 361 44769 381 44797
rect 361 44763 375 44769
rect 400 44763 411 44807
rect 442 44802 500 44809
rect 466 44801 500 44802
rect 565 44801 599 44809
rect 497 44785 500 44801
rect 596 44785 599 44801
rect 466 44784 500 44785
rect 442 44777 500 44784
rect 565 44777 599 44785
rect 612 44768 614 44818
rect 332 44739 342 44763
rect 336 44727 342 44739
rect 224 44671 226 44687
rect 332 44659 342 44727
rect 400 44731 404 44739
rect 400 44697 408 44731
rect 434 44697 438 44731
rect 454 44715 504 44717
rect 504 44699 506 44715
rect 514 44709 530 44715
rect 532 44709 548 44715
rect 525 44699 548 44708
rect 400 44689 404 44697
rect 498 44689 506 44699
rect 504 44665 506 44689
rect 514 44679 515 44699
rect 525 44674 528 44699
rect 547 44679 548 44699
rect 557 44689 564 44699
rect 514 44665 548 44669
rect 151 44618 156 44652
rect 174 44649 246 44657
rect 256 44649 328 44657
rect 336 44651 342 44659
rect 400 44654 404 44659
rect 180 44621 185 44649
rect 174 44613 246 44621
rect 256 44613 328 44621
rect 332 44619 336 44649
rect 400 44620 438 44654
rect 224 44583 226 44599
rect 196 44575 226 44583
rect 196 44571 232 44575
rect 196 44541 204 44571
rect 216 44541 232 44571
rect 224 44494 226 44541
rect 300 44514 308 44583
rect 332 44581 342 44619
rect 400 44611 404 44620
rect 454 44605 504 44607
rect 494 44601 548 44605
rect 494 44596 514 44601
rect 504 44581 506 44596
rect 336 44569 342 44581
rect 289 44504 308 44514
rect 300 44498 308 44504
rect 332 44535 342 44569
rect 400 44573 404 44581
rect 400 44539 408 44573
rect 434 44539 438 44573
rect 498 44571 506 44581
rect 514 44571 515 44591
rect 504 44555 506 44571
rect 525 44562 528 44596
rect 547 44571 548 44591
rect 557 44571 564 44581
rect 514 44555 530 44561
rect 532 44555 548 44561
rect 332 44507 373 44535
rect 332 44501 351 44507
rect 107 44447 119 44481
rect 129 44447 149 44481
rect 196 44460 204 44494
rect 216 44460 232 44494
rect 244 44488 257 44494
rect 278 44488 291 44498
rect 244 44464 291 44488
rect 300 44488 321 44498
rect 336 44491 351 44501
rect 300 44464 329 44488
rect 332 44473 351 44491
rect 361 44501 375 44507
rect 400 44501 411 44539
rect 562 44502 612 44504
rect 361 44473 381 44501
rect 400 44473 409 44501
rect 466 44493 497 44501
rect 565 44493 596 44501
rect 442 44486 500 44493
rect 466 44485 500 44486
rect 565 44485 599 44493
rect 244 44460 257 44464
rect 42 44381 46 44415
rect 72 44381 76 44415
rect 42 44334 76 44338
rect 42 44319 46 44334
rect 72 44319 76 44334
rect 38 44301 80 44319
rect 16 44295 102 44301
rect 144 44295 148 44447
rect 174 44423 181 44451
rect 224 44413 226 44460
rect 300 44451 308 44464
rect 278 44440 305 44451
rect 332 44423 342 44473
rect 400 44453 404 44473
rect 497 44469 500 44485
rect 596 44469 599 44485
rect 466 44468 500 44469
rect 442 44461 500 44468
rect 565 44461 599 44469
rect 612 44452 614 44502
rect 256 44413 328 44421
rect 336 44415 342 44423
rect 400 44415 404 44423
rect 196 44383 204 44413
rect 216 44383 232 44413
rect 196 44379 232 44383
rect 196 44371 226 44379
rect 224 44355 226 44371
rect 332 44343 336 44411
rect 400 44381 408 44415
rect 434 44381 438 44415
rect 454 44399 504 44401
rect 504 44383 506 44399
rect 514 44393 530 44399
rect 532 44393 548 44399
rect 525 44383 548 44392
rect 400 44373 404 44381
rect 498 44373 506 44383
rect 504 44349 506 44373
rect 514 44363 515 44383
rect 525 44358 528 44383
rect 547 44363 548 44383
rect 557 44373 564 44383
rect 514 44349 548 44353
rect 400 44343 442 44344
rect 174 44333 246 44341
rect 400 44336 404 44343
rect 295 44302 300 44336
rect 324 44302 329 44336
rect 367 44319 438 44336
rect 367 44302 442 44319
rect 400 44301 442 44302
rect 378 44295 464 44301
rect 38 44279 80 44295
rect 400 44279 442 44295
rect -25 44265 25 44267
rect 42 44265 76 44279
rect 404 44265 438 44279
rect 455 44265 505 44267
rect 557 44265 607 44267
rect 16 44257 102 44265
rect 378 44257 464 44265
rect 8 44223 17 44257
rect 18 44255 51 44257
rect 80 44255 100 44257
rect 18 44223 100 44255
rect 380 44255 404 44257
rect 429 44255 438 44257
rect 442 44255 462 44257
rect 16 44215 102 44223
rect 42 44199 76 44215
rect 16 44179 38 44185
rect 42 44176 76 44180
rect 80 44179 102 44185
rect 42 44146 46 44176
rect 72 44146 76 44176
rect 42 44065 46 44099
rect 72 44065 76 44099
rect -25 44028 25 44030
rect -8 44020 14 44027
rect -8 44019 17 44020
rect 25 44019 27 44028
rect -12 44012 38 44019
rect -12 44011 34 44012
rect -12 44007 8 44011
rect 0 43995 8 44007
rect 14 43995 34 44011
rect 0 43994 34 43995
rect 0 43987 38 43994
rect 14 43986 17 43987
rect 25 43978 27 43987
rect 42 43958 45 44048
rect 69 44033 80 44065
rect 107 44033 143 44061
rect 144 44033 148 44253
rect 332 44185 336 44253
rect 380 44223 462 44255
rect 463 44223 472 44257
rect 480 44223 497 44257
rect 378 44215 464 44223
rect 505 44215 507 44265
rect 514 44223 548 44257
rect 565 44223 582 44257
rect 607 44215 609 44265
rect 404 44199 438 44215
rect 400 44185 442 44186
rect 378 44179 404 44185
rect 442 44179 464 44185
rect 400 44178 404 44179
rect 174 44139 246 44147
rect 295 44144 300 44178
rect 324 44144 329 44178
rect 224 44109 226 44125
rect 196 44101 226 44109
rect 332 44107 336 44175
rect 367 44144 438 44178
rect 400 44137 404 44144
rect 454 44131 504 44133
rect 494 44127 548 44131
rect 494 44122 514 44127
rect 504 44107 506 44122
rect 196 44097 232 44101
rect 196 44067 204 44097
rect 216 44067 232 44097
rect 400 44099 404 44107
rect 107 44027 119 44033
rect 109 43999 119 44027
rect 129 43999 149 44033
rect 174 44029 181 44059
rect 224 44020 226 44067
rect 256 44059 328 44067
rect 332 44065 336 44095
rect 400 44065 408 44099
rect 434 44065 438 44099
rect 498 44097 506 44107
rect 514 44097 515 44117
rect 504 44081 506 44097
rect 525 44088 528 44122
rect 547 44097 548 44117
rect 557 44097 564 44107
rect 514 44081 530 44087
rect 532 44081 548 44087
rect 278 44029 305 44040
rect 42 43907 46 43941
rect 72 43907 76 43941
rect 38 43869 80 43870
rect 42 43828 76 43862
rect 79 43828 113 43862
rect 42 43749 46 43783
rect 72 43749 76 43783
rect -25 43712 25 43714
rect -8 43704 14 43711
rect -8 43703 17 43704
rect 25 43703 27 43712
rect -12 43696 38 43703
rect -12 43695 34 43696
rect -12 43691 8 43695
rect 0 43679 8 43691
rect 14 43679 34 43695
rect 0 43678 34 43679
rect 0 43671 38 43678
rect 14 43670 17 43671
rect 25 43662 27 43671
rect 42 43642 45 43732
rect 71 43701 80 43729
rect 69 43663 80 43701
rect 144 43691 148 43999
rect 196 43986 204 44020
rect 216 43986 232 44020
rect 244 44016 257 44020
rect 300 44016 308 44029
rect 332 44027 342 44065
rect 400 44057 404 44065
rect 336 44017 342 44027
rect 244 43992 291 44016
rect 244 43986 257 43992
rect 224 43939 226 43986
rect 278 43982 291 43992
rect 300 43992 329 44016
rect 332 44007 342 44017
rect 400 44017 409 44045
rect 562 44028 612 44030
rect 466 44019 497 44027
rect 565 44019 596 44027
rect 300 43982 321 43992
rect 300 43976 308 43982
rect 289 43966 308 43976
rect 196 43909 204 43939
rect 216 43909 232 43939
rect 196 43905 232 43909
rect 196 43897 226 43905
rect 300 43897 308 43966
rect 332 43973 351 44007
rect 361 43979 381 44007
rect 361 43973 375 43979
rect 400 43973 411 44017
rect 442 44012 500 44019
rect 466 44011 500 44012
rect 565 44011 599 44019
rect 497 43995 500 44011
rect 596 43995 599 44011
rect 466 43994 500 43995
rect 442 43987 500 43994
rect 565 43987 599 43995
rect 612 43978 614 44028
rect 332 43949 342 43973
rect 336 43937 342 43949
rect 224 43881 226 43897
rect 332 43869 342 43937
rect 400 43941 404 43949
rect 400 43907 408 43941
rect 434 43907 438 43941
rect 454 43925 504 43927
rect 504 43909 506 43925
rect 514 43919 530 43925
rect 532 43919 548 43925
rect 525 43909 548 43918
rect 400 43899 404 43907
rect 498 43899 506 43909
rect 504 43875 506 43899
rect 514 43889 515 43909
rect 525 43884 528 43909
rect 547 43889 548 43909
rect 557 43899 564 43909
rect 514 43875 548 43879
rect 151 43828 156 43862
rect 174 43859 246 43867
rect 256 43859 328 43867
rect 336 43861 342 43869
rect 400 43864 404 43869
rect 180 43831 185 43859
rect 174 43823 246 43831
rect 256 43823 328 43831
rect 332 43829 336 43859
rect 400 43830 438 43864
rect 224 43793 226 43809
rect 196 43785 226 43793
rect 196 43781 232 43785
rect 196 43751 204 43781
rect 216 43751 232 43781
rect 224 43704 226 43751
rect 300 43724 308 43793
rect 332 43791 342 43829
rect 400 43821 404 43830
rect 454 43815 504 43817
rect 494 43811 548 43815
rect 494 43806 514 43811
rect 504 43791 506 43806
rect 336 43779 342 43791
rect 289 43714 308 43724
rect 300 43708 308 43714
rect 332 43745 342 43779
rect 400 43783 404 43791
rect 400 43749 408 43783
rect 434 43749 438 43783
rect 498 43781 506 43791
rect 514 43781 515 43801
rect 504 43765 506 43781
rect 525 43772 528 43806
rect 547 43781 548 43801
rect 557 43781 564 43791
rect 514 43765 530 43771
rect 532 43765 548 43771
rect 332 43717 373 43745
rect 332 43711 351 43717
rect 107 43657 119 43691
rect 129 43657 149 43691
rect 196 43670 204 43704
rect 216 43670 232 43704
rect 244 43698 257 43704
rect 278 43698 291 43708
rect 244 43674 291 43698
rect 300 43698 321 43708
rect 336 43701 351 43711
rect 300 43674 329 43698
rect 332 43683 351 43701
rect 361 43711 375 43717
rect 400 43711 411 43749
rect 562 43712 612 43714
rect 361 43683 381 43711
rect 400 43683 409 43711
rect 466 43703 497 43711
rect 565 43703 596 43711
rect 442 43696 500 43703
rect 466 43695 500 43696
rect 565 43695 599 43703
rect 244 43670 257 43674
rect 42 43591 46 43625
rect 72 43591 76 43625
rect 42 43544 76 43548
rect 42 43529 46 43544
rect 72 43529 76 43544
rect 38 43511 80 43529
rect 16 43505 102 43511
rect 144 43505 148 43657
rect 174 43633 181 43661
rect 224 43623 226 43670
rect 300 43661 308 43674
rect 278 43650 305 43661
rect 332 43633 342 43683
rect 400 43663 404 43683
rect 497 43679 500 43695
rect 596 43679 599 43695
rect 466 43678 500 43679
rect 442 43671 500 43678
rect 565 43671 599 43679
rect 612 43662 614 43712
rect 256 43623 328 43631
rect 336 43625 342 43633
rect 400 43625 404 43633
rect 196 43593 204 43623
rect 216 43593 232 43623
rect 196 43589 232 43593
rect 196 43581 226 43589
rect 224 43565 226 43581
rect 332 43553 336 43621
rect 400 43591 408 43625
rect 434 43591 438 43625
rect 454 43609 504 43611
rect 504 43593 506 43609
rect 514 43603 530 43609
rect 532 43603 548 43609
rect 525 43593 548 43602
rect 400 43583 404 43591
rect 498 43583 506 43593
rect 504 43559 506 43583
rect 514 43573 515 43593
rect 525 43568 528 43593
rect 547 43573 548 43593
rect 557 43583 564 43593
rect 514 43559 548 43563
rect 400 43553 442 43554
rect 174 43543 246 43551
rect 400 43546 404 43553
rect 295 43512 300 43546
rect 324 43512 329 43546
rect 367 43529 438 43546
rect 367 43512 442 43529
rect 400 43511 442 43512
rect 378 43505 464 43511
rect 38 43489 80 43505
rect 400 43489 442 43505
rect -25 43475 25 43477
rect 42 43475 76 43489
rect 404 43475 438 43489
rect 455 43475 505 43477
rect 557 43475 607 43477
rect 16 43467 102 43475
rect 378 43467 464 43475
rect 8 43433 17 43467
rect 18 43465 51 43467
rect 80 43465 100 43467
rect 18 43433 100 43465
rect 380 43465 404 43467
rect 429 43465 438 43467
rect 442 43465 462 43467
rect 16 43425 102 43433
rect 42 43409 76 43425
rect 16 43389 38 43395
rect 42 43386 76 43390
rect 80 43389 102 43395
rect 42 43356 46 43386
rect 72 43356 76 43386
rect 42 43275 46 43309
rect 72 43275 76 43309
rect -25 43238 25 43240
rect -8 43230 14 43237
rect -8 43229 17 43230
rect 25 43229 27 43238
rect -12 43222 38 43229
rect -12 43221 34 43222
rect -12 43217 8 43221
rect 0 43205 8 43217
rect 14 43205 34 43221
rect 0 43204 34 43205
rect 0 43197 38 43204
rect 14 43196 17 43197
rect 25 43188 27 43197
rect 42 43168 45 43258
rect 69 43243 80 43275
rect 107 43243 143 43271
rect 144 43243 148 43463
rect 332 43395 336 43463
rect 380 43433 462 43465
rect 463 43433 472 43467
rect 480 43433 497 43467
rect 378 43425 464 43433
rect 505 43425 507 43475
rect 514 43433 548 43467
rect 565 43433 582 43467
rect 607 43425 609 43475
rect 404 43409 438 43425
rect 400 43395 442 43396
rect 378 43389 404 43395
rect 442 43389 464 43395
rect 400 43388 404 43389
rect 174 43349 246 43357
rect 295 43354 300 43388
rect 324 43354 329 43388
rect 224 43319 226 43335
rect 196 43311 226 43319
rect 332 43317 336 43385
rect 367 43354 438 43388
rect 400 43347 404 43354
rect 454 43341 504 43343
rect 494 43337 548 43341
rect 494 43332 514 43337
rect 504 43317 506 43332
rect 196 43307 232 43311
rect 196 43277 204 43307
rect 216 43277 232 43307
rect 400 43309 404 43317
rect 107 43237 119 43243
rect 109 43209 119 43237
rect 129 43209 149 43243
rect 174 43239 181 43269
rect 224 43230 226 43277
rect 256 43269 328 43277
rect 332 43275 336 43305
rect 400 43275 408 43309
rect 434 43275 438 43309
rect 498 43307 506 43317
rect 514 43307 515 43327
rect 504 43291 506 43307
rect 525 43298 528 43332
rect 547 43307 548 43327
rect 557 43307 564 43317
rect 514 43291 530 43297
rect 532 43291 548 43297
rect 278 43239 305 43250
rect 42 43117 46 43151
rect 72 43117 76 43151
rect 38 43079 80 43080
rect 42 43038 76 43072
rect 79 43038 113 43072
rect 42 42959 46 42993
rect 72 42959 76 42993
rect -25 42922 25 42924
rect -8 42914 14 42921
rect -8 42913 17 42914
rect 25 42913 27 42922
rect -12 42906 38 42913
rect -12 42905 34 42906
rect -12 42901 8 42905
rect 0 42889 8 42901
rect 14 42889 34 42905
rect 0 42888 34 42889
rect 0 42881 38 42888
rect 14 42880 17 42881
rect 25 42872 27 42881
rect 42 42852 45 42942
rect 71 42911 80 42939
rect 69 42873 80 42911
rect 144 42901 148 43209
rect 196 43196 204 43230
rect 216 43196 232 43230
rect 244 43226 257 43230
rect 300 43226 308 43239
rect 332 43237 342 43275
rect 400 43267 404 43275
rect 336 43227 342 43237
rect 244 43202 291 43226
rect 244 43196 257 43202
rect 224 43149 226 43196
rect 278 43192 291 43202
rect 300 43202 329 43226
rect 332 43217 342 43227
rect 400 43227 409 43255
rect 562 43238 612 43240
rect 466 43229 497 43237
rect 565 43229 596 43237
rect 300 43192 321 43202
rect 300 43186 308 43192
rect 289 43176 308 43186
rect 196 43119 204 43149
rect 216 43119 232 43149
rect 196 43115 232 43119
rect 196 43107 226 43115
rect 300 43107 308 43176
rect 332 43183 351 43217
rect 361 43189 381 43217
rect 361 43183 375 43189
rect 400 43183 411 43227
rect 442 43222 500 43229
rect 466 43221 500 43222
rect 565 43221 599 43229
rect 497 43205 500 43221
rect 596 43205 599 43221
rect 466 43204 500 43205
rect 442 43197 500 43204
rect 565 43197 599 43205
rect 612 43188 614 43238
rect 332 43159 342 43183
rect 336 43147 342 43159
rect 224 43091 226 43107
rect 332 43079 342 43147
rect 400 43151 404 43159
rect 400 43117 408 43151
rect 434 43117 438 43151
rect 454 43135 504 43137
rect 504 43119 506 43135
rect 514 43129 530 43135
rect 532 43129 548 43135
rect 525 43119 548 43128
rect 400 43109 404 43117
rect 498 43109 506 43119
rect 504 43085 506 43109
rect 514 43099 515 43119
rect 525 43094 528 43119
rect 547 43099 548 43119
rect 557 43109 564 43119
rect 514 43085 548 43089
rect 151 43038 156 43072
rect 174 43069 246 43077
rect 256 43069 328 43077
rect 336 43071 342 43079
rect 400 43074 404 43079
rect 180 43041 185 43069
rect 174 43033 246 43041
rect 256 43033 328 43041
rect 332 43039 336 43069
rect 400 43040 438 43074
rect 224 43003 226 43019
rect 196 42995 226 43003
rect 196 42991 232 42995
rect 196 42961 204 42991
rect 216 42961 232 42991
rect 224 42914 226 42961
rect 300 42934 308 43003
rect 332 43001 342 43039
rect 400 43031 404 43040
rect 454 43025 504 43027
rect 494 43021 548 43025
rect 494 43016 514 43021
rect 504 43001 506 43016
rect 336 42989 342 43001
rect 289 42924 308 42934
rect 300 42918 308 42924
rect 332 42955 342 42989
rect 400 42993 404 43001
rect 400 42959 408 42993
rect 434 42959 438 42993
rect 498 42991 506 43001
rect 514 42991 515 43011
rect 504 42975 506 42991
rect 525 42982 528 43016
rect 547 42991 548 43011
rect 557 42991 564 43001
rect 514 42975 530 42981
rect 532 42975 548 42981
rect 332 42927 373 42955
rect 332 42921 351 42927
rect 107 42867 119 42901
rect 129 42867 149 42901
rect 196 42880 204 42914
rect 216 42880 232 42914
rect 244 42908 257 42914
rect 278 42908 291 42918
rect 244 42884 291 42908
rect 300 42908 321 42918
rect 336 42911 351 42921
rect 300 42884 329 42908
rect 332 42893 351 42911
rect 361 42921 375 42927
rect 400 42921 411 42959
rect 562 42922 612 42924
rect 361 42893 381 42921
rect 400 42893 409 42921
rect 466 42913 497 42921
rect 565 42913 596 42921
rect 442 42906 500 42913
rect 466 42905 500 42906
rect 565 42905 599 42913
rect 244 42880 257 42884
rect 42 42801 46 42835
rect 72 42801 76 42835
rect 42 42754 76 42758
rect 42 42739 46 42754
rect 72 42739 76 42754
rect 38 42721 80 42739
rect 16 42715 102 42721
rect 144 42715 148 42867
rect 174 42843 181 42871
rect 224 42833 226 42880
rect 300 42871 308 42884
rect 278 42860 305 42871
rect 332 42843 342 42893
rect 400 42873 404 42893
rect 497 42889 500 42905
rect 596 42889 599 42905
rect 466 42888 500 42889
rect 442 42881 500 42888
rect 565 42881 599 42889
rect 612 42872 614 42922
rect 256 42833 328 42841
rect 336 42835 342 42843
rect 400 42835 404 42843
rect 196 42803 204 42833
rect 216 42803 232 42833
rect 196 42799 232 42803
rect 196 42791 226 42799
rect 224 42775 226 42791
rect 332 42763 336 42831
rect 400 42801 408 42835
rect 434 42801 438 42835
rect 454 42819 504 42821
rect 504 42803 506 42819
rect 514 42813 530 42819
rect 532 42813 548 42819
rect 525 42803 548 42812
rect 400 42793 404 42801
rect 498 42793 506 42803
rect 504 42769 506 42793
rect 514 42783 515 42803
rect 525 42778 528 42803
rect 547 42783 548 42803
rect 557 42793 564 42803
rect 514 42769 548 42773
rect 400 42763 442 42764
rect 174 42753 246 42761
rect 400 42756 404 42763
rect 295 42722 300 42756
rect 324 42722 329 42756
rect 367 42739 438 42756
rect 367 42722 442 42739
rect 400 42721 442 42722
rect 378 42715 464 42721
rect 38 42699 80 42715
rect 400 42699 442 42715
rect -25 42685 25 42687
rect 42 42685 76 42699
rect 404 42685 438 42699
rect 455 42685 505 42687
rect 557 42685 607 42687
rect 16 42677 102 42685
rect 378 42677 464 42685
rect 8 42643 17 42677
rect 18 42675 51 42677
rect 80 42675 100 42677
rect 18 42643 100 42675
rect 380 42675 404 42677
rect 429 42675 438 42677
rect 442 42675 462 42677
rect 16 42635 102 42643
rect 42 42619 76 42635
rect 16 42599 38 42605
rect 42 42596 76 42600
rect 80 42599 102 42605
rect 42 42566 46 42596
rect 72 42566 76 42596
rect 42 42485 46 42519
rect 72 42485 76 42519
rect -25 42448 25 42450
rect -8 42440 14 42447
rect -8 42439 17 42440
rect 25 42439 27 42448
rect -12 42432 38 42439
rect -12 42431 34 42432
rect -12 42427 8 42431
rect 0 42415 8 42427
rect 14 42415 34 42431
rect 0 42414 34 42415
rect 0 42407 38 42414
rect 14 42406 17 42407
rect 25 42398 27 42407
rect 42 42378 45 42468
rect 69 42453 80 42485
rect 107 42453 143 42481
rect 144 42453 148 42673
rect 332 42605 336 42673
rect 380 42643 462 42675
rect 463 42643 472 42677
rect 480 42643 497 42677
rect 378 42635 464 42643
rect 505 42635 507 42685
rect 514 42643 548 42677
rect 565 42643 582 42677
rect 607 42635 609 42685
rect 404 42619 438 42635
rect 400 42605 442 42606
rect 378 42599 404 42605
rect 442 42599 464 42605
rect 400 42598 404 42599
rect 174 42559 246 42567
rect 295 42564 300 42598
rect 324 42564 329 42598
rect 224 42529 226 42545
rect 196 42521 226 42529
rect 332 42527 336 42595
rect 367 42564 438 42598
rect 400 42557 404 42564
rect 454 42551 504 42553
rect 494 42547 548 42551
rect 494 42542 514 42547
rect 504 42527 506 42542
rect 196 42517 232 42521
rect 196 42487 204 42517
rect 216 42487 232 42517
rect 400 42519 404 42527
rect 107 42447 119 42453
rect 109 42419 119 42447
rect 129 42419 149 42453
rect 174 42449 181 42479
rect 224 42440 226 42487
rect 256 42479 328 42487
rect 332 42485 336 42515
rect 400 42485 408 42519
rect 434 42485 438 42519
rect 498 42517 506 42527
rect 514 42517 515 42537
rect 504 42501 506 42517
rect 525 42508 528 42542
rect 547 42517 548 42537
rect 557 42517 564 42527
rect 514 42501 530 42507
rect 532 42501 548 42507
rect 278 42449 305 42460
rect 42 42327 46 42361
rect 72 42327 76 42361
rect 38 42289 80 42290
rect 42 42248 76 42282
rect 79 42248 113 42282
rect 42 42169 46 42203
rect 72 42169 76 42203
rect -25 42132 25 42134
rect -8 42124 14 42131
rect -8 42123 17 42124
rect 25 42123 27 42132
rect -12 42116 38 42123
rect -12 42115 34 42116
rect -12 42111 8 42115
rect 0 42099 8 42111
rect 14 42099 34 42115
rect 0 42098 34 42099
rect 0 42091 38 42098
rect 14 42090 17 42091
rect 25 42082 27 42091
rect 42 42062 45 42152
rect 71 42121 80 42149
rect 69 42083 80 42121
rect 144 42111 148 42419
rect 196 42406 204 42440
rect 216 42406 232 42440
rect 244 42436 257 42440
rect 300 42436 308 42449
rect 332 42447 342 42485
rect 400 42477 404 42485
rect 336 42437 342 42447
rect 244 42412 291 42436
rect 244 42406 257 42412
rect 224 42359 226 42406
rect 278 42402 291 42412
rect 300 42412 329 42436
rect 332 42427 342 42437
rect 400 42437 409 42465
rect 562 42448 612 42450
rect 466 42439 497 42447
rect 565 42439 596 42447
rect 300 42402 321 42412
rect 300 42396 308 42402
rect 289 42386 308 42396
rect 196 42329 204 42359
rect 216 42329 232 42359
rect 196 42325 232 42329
rect 196 42317 226 42325
rect 300 42317 308 42386
rect 332 42393 351 42427
rect 361 42399 381 42427
rect 361 42393 375 42399
rect 400 42393 411 42437
rect 442 42432 500 42439
rect 466 42431 500 42432
rect 565 42431 599 42439
rect 497 42415 500 42431
rect 596 42415 599 42431
rect 466 42414 500 42415
rect 442 42407 500 42414
rect 565 42407 599 42415
rect 612 42398 614 42448
rect 332 42369 342 42393
rect 336 42357 342 42369
rect 224 42301 226 42317
rect 332 42289 342 42357
rect 400 42361 404 42369
rect 400 42327 408 42361
rect 434 42327 438 42361
rect 454 42345 504 42347
rect 504 42329 506 42345
rect 514 42339 530 42345
rect 532 42339 548 42345
rect 525 42329 548 42338
rect 400 42319 404 42327
rect 498 42319 506 42329
rect 504 42295 506 42319
rect 514 42309 515 42329
rect 525 42304 528 42329
rect 547 42309 548 42329
rect 557 42319 564 42329
rect 514 42295 548 42299
rect 151 42248 156 42282
rect 174 42279 246 42287
rect 256 42279 328 42287
rect 336 42281 342 42289
rect 400 42284 404 42289
rect 180 42251 185 42279
rect 174 42243 246 42251
rect 256 42243 328 42251
rect 332 42249 336 42279
rect 400 42250 438 42284
rect 224 42213 226 42229
rect 196 42205 226 42213
rect 196 42201 232 42205
rect 196 42171 204 42201
rect 216 42171 232 42201
rect 224 42124 226 42171
rect 300 42144 308 42213
rect 332 42211 342 42249
rect 400 42241 404 42250
rect 454 42235 504 42237
rect 494 42231 548 42235
rect 494 42226 514 42231
rect 504 42211 506 42226
rect 336 42199 342 42211
rect 289 42134 308 42144
rect 300 42128 308 42134
rect 332 42165 342 42199
rect 400 42203 404 42211
rect 400 42169 408 42203
rect 434 42169 438 42203
rect 498 42201 506 42211
rect 514 42201 515 42221
rect 504 42185 506 42201
rect 525 42192 528 42226
rect 547 42201 548 42221
rect 557 42201 564 42211
rect 514 42185 530 42191
rect 532 42185 548 42191
rect 332 42137 373 42165
rect 332 42131 351 42137
rect 107 42077 119 42111
rect 129 42077 149 42111
rect 196 42090 204 42124
rect 216 42090 232 42124
rect 244 42118 257 42124
rect 278 42118 291 42128
rect 244 42094 291 42118
rect 300 42118 321 42128
rect 336 42121 351 42131
rect 300 42094 329 42118
rect 332 42103 351 42121
rect 361 42131 375 42137
rect 400 42131 411 42169
rect 562 42132 612 42134
rect 361 42103 381 42131
rect 400 42103 409 42131
rect 466 42123 497 42131
rect 565 42123 596 42131
rect 442 42116 500 42123
rect 466 42115 500 42116
rect 565 42115 599 42123
rect 244 42090 257 42094
rect 42 42011 46 42045
rect 72 42011 76 42045
rect 42 41964 76 41968
rect 42 41949 46 41964
rect 72 41949 76 41964
rect 38 41931 80 41949
rect 16 41925 102 41931
rect 144 41925 148 42077
rect 174 42053 181 42081
rect 224 42043 226 42090
rect 300 42081 308 42094
rect 278 42070 305 42081
rect 332 42053 342 42103
rect 400 42083 404 42103
rect 497 42099 500 42115
rect 596 42099 599 42115
rect 466 42098 500 42099
rect 442 42091 500 42098
rect 565 42091 599 42099
rect 612 42082 614 42132
rect 256 42043 328 42051
rect 336 42045 342 42053
rect 400 42045 404 42053
rect 196 42013 204 42043
rect 216 42013 232 42043
rect 196 42009 232 42013
rect 196 42001 226 42009
rect 224 41985 226 42001
rect 332 41973 336 42041
rect 400 42011 408 42045
rect 434 42011 438 42045
rect 454 42029 504 42031
rect 504 42013 506 42029
rect 514 42023 530 42029
rect 532 42023 548 42029
rect 525 42013 548 42022
rect 400 42003 404 42011
rect 498 42003 506 42013
rect 504 41979 506 42003
rect 514 41993 515 42013
rect 525 41988 528 42013
rect 547 41993 548 42013
rect 557 42003 564 42013
rect 514 41979 548 41983
rect 400 41973 442 41974
rect 174 41963 246 41971
rect 400 41966 404 41973
rect 295 41932 300 41966
rect 324 41932 329 41966
rect 367 41949 438 41966
rect 367 41932 442 41949
rect 400 41931 442 41932
rect 378 41925 464 41931
rect 38 41909 80 41925
rect 400 41909 442 41925
rect -25 41895 25 41897
rect 42 41895 76 41909
rect 404 41895 438 41909
rect 455 41895 505 41897
rect 557 41895 607 41897
rect 16 41887 102 41895
rect 378 41887 464 41895
rect 8 41853 17 41887
rect 18 41885 51 41887
rect 80 41885 100 41887
rect 18 41853 100 41885
rect 380 41885 404 41887
rect 429 41885 438 41887
rect 442 41885 462 41887
rect 16 41845 102 41853
rect 42 41829 76 41845
rect 16 41809 38 41815
rect 42 41806 76 41810
rect 80 41809 102 41815
rect 42 41776 46 41806
rect 72 41776 76 41806
rect 42 41695 46 41729
rect 72 41695 76 41729
rect -25 41658 25 41660
rect -8 41650 14 41657
rect -8 41649 17 41650
rect 25 41649 27 41658
rect -12 41642 38 41649
rect -12 41641 34 41642
rect -12 41637 8 41641
rect 0 41625 8 41637
rect 14 41625 34 41641
rect 0 41624 34 41625
rect 0 41617 38 41624
rect 14 41616 17 41617
rect 25 41608 27 41617
rect 42 41588 45 41678
rect 69 41663 80 41695
rect 107 41663 143 41691
rect 144 41663 148 41883
rect 332 41815 336 41883
rect 380 41853 462 41885
rect 463 41853 472 41887
rect 480 41853 497 41887
rect 378 41845 464 41853
rect 505 41845 507 41895
rect 514 41853 548 41887
rect 565 41853 582 41887
rect 607 41845 609 41895
rect 404 41829 438 41845
rect 400 41815 442 41816
rect 378 41809 404 41815
rect 442 41809 464 41815
rect 400 41808 404 41809
rect 174 41769 246 41777
rect 295 41774 300 41808
rect 324 41774 329 41808
rect 224 41739 226 41755
rect 196 41731 226 41739
rect 332 41737 336 41805
rect 367 41774 438 41808
rect 400 41767 404 41774
rect 454 41761 504 41763
rect 494 41757 548 41761
rect 494 41752 514 41757
rect 504 41737 506 41752
rect 196 41727 232 41731
rect 196 41697 204 41727
rect 216 41697 232 41727
rect 400 41729 404 41737
rect 107 41657 119 41663
rect 109 41629 119 41657
rect 129 41629 149 41663
rect 174 41659 181 41689
rect 224 41650 226 41697
rect 256 41689 328 41697
rect 332 41695 336 41725
rect 400 41695 408 41729
rect 434 41695 438 41729
rect 498 41727 506 41737
rect 514 41727 515 41747
rect 504 41711 506 41727
rect 525 41718 528 41752
rect 547 41727 548 41747
rect 557 41727 564 41737
rect 514 41711 530 41717
rect 532 41711 548 41717
rect 278 41659 305 41670
rect 42 41537 46 41571
rect 72 41537 76 41571
rect 38 41499 80 41500
rect 42 41458 76 41492
rect 79 41458 113 41492
rect 42 41379 46 41413
rect 72 41379 76 41413
rect -25 41342 25 41344
rect -8 41334 14 41341
rect -8 41333 17 41334
rect 25 41333 27 41342
rect -12 41326 38 41333
rect -12 41325 34 41326
rect -12 41321 8 41325
rect 0 41309 8 41321
rect 14 41309 34 41325
rect 0 41308 34 41309
rect 0 41301 38 41308
rect 14 41300 17 41301
rect 25 41292 27 41301
rect 42 41272 45 41362
rect 71 41331 80 41359
rect 69 41293 80 41331
rect 144 41321 148 41629
rect 196 41616 204 41650
rect 216 41616 232 41650
rect 244 41646 257 41650
rect 300 41646 308 41659
rect 332 41657 342 41695
rect 400 41687 404 41695
rect 336 41647 342 41657
rect 244 41622 291 41646
rect 244 41616 257 41622
rect 224 41569 226 41616
rect 278 41612 291 41622
rect 300 41622 329 41646
rect 332 41637 342 41647
rect 400 41647 409 41675
rect 562 41658 612 41660
rect 466 41649 497 41657
rect 565 41649 596 41657
rect 300 41612 321 41622
rect 300 41606 308 41612
rect 289 41596 308 41606
rect 196 41539 204 41569
rect 216 41539 232 41569
rect 196 41535 232 41539
rect 196 41527 226 41535
rect 300 41527 308 41596
rect 332 41603 351 41637
rect 361 41609 381 41637
rect 361 41603 375 41609
rect 400 41603 411 41647
rect 442 41642 500 41649
rect 466 41641 500 41642
rect 565 41641 599 41649
rect 497 41625 500 41641
rect 596 41625 599 41641
rect 466 41624 500 41625
rect 442 41617 500 41624
rect 565 41617 599 41625
rect 612 41608 614 41658
rect 332 41579 342 41603
rect 336 41567 342 41579
rect 224 41511 226 41527
rect 332 41499 342 41567
rect 400 41571 404 41579
rect 400 41537 408 41571
rect 434 41537 438 41571
rect 454 41555 504 41557
rect 504 41539 506 41555
rect 514 41549 530 41555
rect 532 41549 548 41555
rect 525 41539 548 41548
rect 400 41529 404 41537
rect 498 41529 506 41539
rect 504 41505 506 41529
rect 514 41519 515 41539
rect 525 41514 528 41539
rect 547 41519 548 41539
rect 557 41529 564 41539
rect 514 41505 548 41509
rect 151 41458 156 41492
rect 174 41489 246 41497
rect 256 41489 328 41497
rect 336 41491 342 41499
rect 400 41494 404 41499
rect 180 41461 185 41489
rect 174 41453 246 41461
rect 256 41453 328 41461
rect 332 41459 336 41489
rect 400 41460 438 41494
rect 224 41423 226 41439
rect 196 41415 226 41423
rect 196 41411 232 41415
rect 196 41381 204 41411
rect 216 41381 232 41411
rect 224 41334 226 41381
rect 300 41354 308 41423
rect 332 41421 342 41459
rect 400 41451 404 41460
rect 454 41445 504 41447
rect 494 41441 548 41445
rect 494 41436 514 41441
rect 504 41421 506 41436
rect 336 41409 342 41421
rect 289 41344 308 41354
rect 300 41338 308 41344
rect 332 41375 342 41409
rect 400 41413 404 41421
rect 400 41379 408 41413
rect 434 41379 438 41413
rect 498 41411 506 41421
rect 514 41411 515 41431
rect 504 41395 506 41411
rect 525 41402 528 41436
rect 547 41411 548 41431
rect 557 41411 564 41421
rect 514 41395 530 41401
rect 532 41395 548 41401
rect 332 41347 373 41375
rect 332 41341 351 41347
rect 107 41287 119 41321
rect 129 41287 149 41321
rect 196 41300 204 41334
rect 216 41300 232 41334
rect 244 41328 257 41334
rect 278 41328 291 41338
rect 244 41304 291 41328
rect 300 41328 321 41338
rect 336 41331 351 41341
rect 300 41304 329 41328
rect 332 41313 351 41331
rect 361 41341 375 41347
rect 400 41341 411 41379
rect 562 41342 612 41344
rect 361 41313 381 41341
rect 400 41313 409 41341
rect 466 41333 497 41341
rect 565 41333 596 41341
rect 442 41326 500 41333
rect 466 41325 500 41326
rect 565 41325 599 41333
rect 244 41300 257 41304
rect 42 41221 46 41255
rect 72 41221 76 41255
rect 42 41174 76 41178
rect 42 41159 46 41174
rect 72 41159 76 41174
rect 38 41141 80 41159
rect 16 41135 102 41141
rect 144 41135 148 41287
rect 174 41263 181 41291
rect 224 41253 226 41300
rect 300 41291 308 41304
rect 278 41280 305 41291
rect 332 41263 342 41313
rect 400 41293 404 41313
rect 497 41309 500 41325
rect 596 41309 599 41325
rect 466 41308 500 41309
rect 442 41301 500 41308
rect 565 41301 599 41309
rect 612 41292 614 41342
rect 256 41253 328 41261
rect 336 41255 342 41263
rect 400 41255 404 41263
rect 196 41223 204 41253
rect 216 41223 232 41253
rect 196 41219 232 41223
rect 196 41211 226 41219
rect 224 41195 226 41211
rect 332 41183 336 41251
rect 400 41221 408 41255
rect 434 41221 438 41255
rect 454 41239 504 41241
rect 504 41223 506 41239
rect 514 41233 530 41239
rect 532 41233 548 41239
rect 525 41223 548 41232
rect 400 41213 404 41221
rect 498 41213 506 41223
rect 504 41189 506 41213
rect 514 41203 515 41223
rect 525 41198 528 41223
rect 547 41203 548 41223
rect 557 41213 564 41223
rect 514 41189 548 41193
rect 400 41183 442 41184
rect 174 41173 246 41181
rect 400 41176 404 41183
rect 295 41142 300 41176
rect 324 41142 329 41176
rect 367 41159 438 41176
rect 367 41142 442 41159
rect 400 41141 442 41142
rect 378 41135 464 41141
rect 38 41119 80 41135
rect 400 41119 442 41135
rect -25 41105 25 41107
rect 42 41105 76 41119
rect 404 41105 438 41119
rect 455 41105 505 41107
rect 557 41105 607 41107
rect 16 41097 102 41105
rect 378 41097 464 41105
rect 8 41063 17 41097
rect 18 41095 51 41097
rect 80 41095 100 41097
rect 18 41063 100 41095
rect 380 41095 404 41097
rect 429 41095 438 41097
rect 442 41095 462 41097
rect 16 41055 102 41063
rect 42 41039 76 41055
rect 16 41019 38 41025
rect 42 41016 76 41020
rect 80 41019 102 41025
rect 42 40986 46 41016
rect 72 40986 76 41016
rect 42 40905 46 40939
rect 72 40905 76 40939
rect -25 40868 25 40870
rect -8 40860 14 40867
rect -8 40859 17 40860
rect 25 40859 27 40868
rect -12 40852 38 40859
rect -12 40851 34 40852
rect -12 40847 8 40851
rect 0 40835 8 40847
rect 14 40835 34 40851
rect 0 40834 34 40835
rect 0 40827 38 40834
rect 14 40826 17 40827
rect 25 40818 27 40827
rect 42 40798 45 40888
rect 69 40873 80 40905
rect 107 40873 143 40901
rect 144 40873 148 41093
rect 332 41025 336 41093
rect 380 41063 462 41095
rect 463 41063 472 41097
rect 480 41063 497 41097
rect 378 41055 464 41063
rect 505 41055 507 41105
rect 514 41063 548 41097
rect 565 41063 582 41097
rect 607 41055 609 41105
rect 404 41039 438 41055
rect 400 41025 442 41026
rect 378 41019 404 41025
rect 442 41019 464 41025
rect 400 41018 404 41019
rect 174 40979 246 40987
rect 295 40984 300 41018
rect 324 40984 329 41018
rect 224 40949 226 40965
rect 196 40941 226 40949
rect 332 40947 336 41015
rect 367 40984 438 41018
rect 400 40977 404 40984
rect 454 40971 504 40973
rect 494 40967 548 40971
rect 494 40962 514 40967
rect 504 40947 506 40962
rect 196 40937 232 40941
rect 196 40907 204 40937
rect 216 40907 232 40937
rect 400 40939 404 40947
rect 107 40867 119 40873
rect 109 40839 119 40867
rect 129 40839 149 40873
rect 174 40869 181 40899
rect 224 40860 226 40907
rect 256 40899 328 40907
rect 332 40905 336 40935
rect 400 40905 408 40939
rect 434 40905 438 40939
rect 498 40937 506 40947
rect 514 40937 515 40957
rect 504 40921 506 40937
rect 525 40928 528 40962
rect 547 40937 548 40957
rect 557 40937 564 40947
rect 514 40921 530 40927
rect 532 40921 548 40927
rect 278 40869 305 40880
rect 42 40747 46 40781
rect 72 40747 76 40781
rect 38 40709 80 40710
rect 42 40668 76 40702
rect 79 40668 113 40702
rect 42 40589 46 40623
rect 72 40589 76 40623
rect -25 40552 25 40554
rect -8 40544 14 40551
rect -8 40543 17 40544
rect 25 40543 27 40552
rect -12 40536 38 40543
rect -12 40535 34 40536
rect -12 40531 8 40535
rect 0 40519 8 40531
rect 14 40519 34 40535
rect 0 40518 34 40519
rect 0 40511 38 40518
rect 14 40510 17 40511
rect 25 40502 27 40511
rect 42 40482 45 40572
rect 71 40541 80 40569
rect 69 40503 80 40541
rect 144 40531 148 40839
rect 196 40826 204 40860
rect 216 40826 232 40860
rect 244 40856 257 40860
rect 300 40856 308 40869
rect 332 40867 342 40905
rect 400 40897 404 40905
rect 336 40857 342 40867
rect 244 40832 291 40856
rect 244 40826 257 40832
rect 224 40779 226 40826
rect 278 40822 291 40832
rect 300 40832 329 40856
rect 332 40847 342 40857
rect 400 40857 409 40885
rect 562 40868 612 40870
rect 466 40859 497 40867
rect 565 40859 596 40867
rect 300 40822 321 40832
rect 300 40816 308 40822
rect 289 40806 308 40816
rect 196 40749 204 40779
rect 216 40749 232 40779
rect 196 40745 232 40749
rect 196 40737 226 40745
rect 300 40737 308 40806
rect 332 40813 351 40847
rect 361 40819 381 40847
rect 361 40813 375 40819
rect 400 40813 411 40857
rect 442 40852 500 40859
rect 466 40851 500 40852
rect 565 40851 599 40859
rect 497 40835 500 40851
rect 596 40835 599 40851
rect 466 40834 500 40835
rect 442 40827 500 40834
rect 565 40827 599 40835
rect 612 40818 614 40868
rect 332 40789 342 40813
rect 336 40777 342 40789
rect 224 40721 226 40737
rect 332 40709 342 40777
rect 400 40781 404 40789
rect 400 40747 408 40781
rect 434 40747 438 40781
rect 454 40765 504 40767
rect 504 40749 506 40765
rect 514 40759 530 40765
rect 532 40759 548 40765
rect 525 40749 548 40758
rect 400 40739 404 40747
rect 498 40739 506 40749
rect 504 40715 506 40739
rect 514 40729 515 40749
rect 525 40724 528 40749
rect 547 40729 548 40749
rect 557 40739 564 40749
rect 514 40715 548 40719
rect 151 40668 156 40702
rect 174 40699 246 40707
rect 256 40699 328 40707
rect 336 40701 342 40709
rect 400 40704 404 40709
rect 180 40671 185 40699
rect 174 40663 246 40671
rect 256 40663 328 40671
rect 332 40669 336 40699
rect 400 40670 438 40704
rect 224 40633 226 40649
rect 196 40625 226 40633
rect 196 40621 232 40625
rect 196 40591 204 40621
rect 216 40591 232 40621
rect 224 40544 226 40591
rect 300 40564 308 40633
rect 332 40631 342 40669
rect 400 40661 404 40670
rect 454 40655 504 40657
rect 494 40651 548 40655
rect 494 40646 514 40651
rect 504 40631 506 40646
rect 336 40619 342 40631
rect 289 40554 308 40564
rect 300 40548 308 40554
rect 332 40585 342 40619
rect 400 40623 404 40631
rect 400 40589 408 40623
rect 434 40589 438 40623
rect 498 40621 506 40631
rect 514 40621 515 40641
rect 504 40605 506 40621
rect 525 40612 528 40646
rect 547 40621 548 40641
rect 557 40621 564 40631
rect 514 40605 530 40611
rect 532 40605 548 40611
rect 332 40557 373 40585
rect 332 40551 351 40557
rect 107 40497 119 40531
rect 129 40497 149 40531
rect 196 40510 204 40544
rect 216 40510 232 40544
rect 244 40538 257 40544
rect 278 40538 291 40548
rect 244 40514 291 40538
rect 300 40538 321 40548
rect 336 40541 351 40551
rect 300 40514 329 40538
rect 332 40523 351 40541
rect 361 40551 375 40557
rect 400 40551 411 40589
rect 562 40552 612 40554
rect 361 40523 381 40551
rect 400 40523 409 40551
rect 466 40543 497 40551
rect 565 40543 596 40551
rect 442 40536 500 40543
rect 466 40535 500 40536
rect 565 40535 599 40543
rect 244 40510 257 40514
rect 42 40431 46 40465
rect 72 40431 76 40465
rect 42 40384 76 40388
rect 42 40369 46 40384
rect 72 40369 76 40384
rect 38 40351 80 40369
rect 16 40345 102 40351
rect 144 40345 148 40497
rect 174 40473 181 40501
rect 224 40463 226 40510
rect 300 40501 308 40514
rect 278 40490 305 40501
rect 332 40473 342 40523
rect 400 40503 404 40523
rect 497 40519 500 40535
rect 596 40519 599 40535
rect 466 40518 500 40519
rect 442 40511 500 40518
rect 565 40511 599 40519
rect 612 40502 614 40552
rect 256 40463 328 40471
rect 336 40465 342 40473
rect 400 40465 404 40473
rect 196 40433 204 40463
rect 216 40433 232 40463
rect 196 40429 232 40433
rect 196 40421 226 40429
rect 224 40405 226 40421
rect 332 40393 336 40461
rect 400 40431 408 40465
rect 434 40431 438 40465
rect 454 40449 504 40451
rect 504 40433 506 40449
rect 514 40443 530 40449
rect 532 40443 548 40449
rect 525 40433 548 40442
rect 400 40423 404 40431
rect 498 40423 506 40433
rect 504 40399 506 40423
rect 514 40413 515 40433
rect 525 40408 528 40433
rect 547 40413 548 40433
rect 557 40423 564 40433
rect 514 40399 548 40403
rect 400 40393 442 40394
rect 174 40383 246 40391
rect 400 40386 404 40393
rect 295 40352 300 40386
rect 324 40352 329 40386
rect 367 40369 438 40386
rect 367 40352 442 40369
rect 400 40351 442 40352
rect 378 40345 464 40351
rect 38 40329 80 40345
rect 400 40329 442 40345
rect -25 40315 25 40317
rect 42 40315 76 40329
rect 404 40315 438 40329
rect 455 40315 505 40317
rect 557 40315 607 40317
rect 16 40307 102 40315
rect 378 40307 464 40315
rect 8 40273 17 40307
rect 18 40305 51 40307
rect 80 40305 100 40307
rect 18 40273 100 40305
rect 380 40305 404 40307
rect 429 40305 438 40307
rect 442 40305 462 40307
rect 16 40265 102 40273
rect 42 40249 76 40265
rect 16 40229 38 40235
rect 42 40226 76 40230
rect 80 40229 102 40235
rect 42 40196 46 40226
rect 72 40196 76 40226
rect 42 40115 46 40149
rect 72 40115 76 40149
rect -25 40078 25 40080
rect -8 40070 14 40077
rect -8 40069 17 40070
rect 25 40069 27 40078
rect -12 40062 38 40069
rect -12 40061 34 40062
rect -12 40057 8 40061
rect 0 40045 8 40057
rect 14 40045 34 40061
rect 0 40044 34 40045
rect 0 40037 38 40044
rect 14 40036 17 40037
rect 25 40028 27 40037
rect 42 40008 45 40098
rect 69 40083 80 40115
rect 107 40083 143 40111
rect 144 40083 148 40303
rect 332 40235 336 40303
rect 380 40273 462 40305
rect 463 40273 472 40307
rect 480 40273 497 40307
rect 378 40265 464 40273
rect 505 40265 507 40315
rect 514 40273 548 40307
rect 565 40273 582 40307
rect 607 40265 609 40315
rect 404 40249 438 40265
rect 400 40235 442 40236
rect 378 40229 404 40235
rect 442 40229 464 40235
rect 400 40228 404 40229
rect 174 40189 246 40197
rect 295 40194 300 40228
rect 324 40194 329 40228
rect 224 40159 226 40175
rect 196 40151 226 40159
rect 332 40157 336 40225
rect 367 40194 438 40228
rect 400 40187 404 40194
rect 454 40181 504 40183
rect 494 40177 548 40181
rect 494 40172 514 40177
rect 504 40157 506 40172
rect 196 40147 232 40151
rect 196 40117 204 40147
rect 216 40117 232 40147
rect 400 40149 404 40157
rect 107 40077 119 40083
rect 109 40049 119 40077
rect 129 40049 149 40083
rect 174 40079 181 40109
rect 224 40070 226 40117
rect 256 40109 328 40117
rect 332 40115 336 40145
rect 400 40115 408 40149
rect 434 40115 438 40149
rect 498 40147 506 40157
rect 514 40147 515 40167
rect 504 40131 506 40147
rect 525 40138 528 40172
rect 547 40147 548 40167
rect 557 40147 564 40157
rect 514 40131 530 40137
rect 532 40131 548 40137
rect 278 40079 305 40090
rect 42 39957 46 39991
rect 72 39957 76 39991
rect 38 39919 80 39920
rect 42 39878 76 39912
rect 79 39878 113 39912
rect 42 39799 46 39833
rect 72 39799 76 39833
rect -25 39762 25 39764
rect -8 39754 14 39761
rect -8 39753 17 39754
rect 25 39753 27 39762
rect -12 39746 38 39753
rect -12 39745 34 39746
rect -12 39741 8 39745
rect 0 39729 8 39741
rect 14 39729 34 39745
rect 0 39728 34 39729
rect 0 39721 38 39728
rect 14 39720 17 39721
rect 25 39712 27 39721
rect 42 39692 45 39782
rect 71 39751 80 39779
rect 69 39713 80 39751
rect 144 39741 148 40049
rect 196 40036 204 40070
rect 216 40036 232 40070
rect 244 40066 257 40070
rect 300 40066 308 40079
rect 332 40077 342 40115
rect 400 40107 404 40115
rect 336 40067 342 40077
rect 244 40042 291 40066
rect 244 40036 257 40042
rect 224 39989 226 40036
rect 278 40032 291 40042
rect 300 40042 329 40066
rect 332 40057 342 40067
rect 400 40067 409 40095
rect 562 40078 612 40080
rect 466 40069 497 40077
rect 565 40069 596 40077
rect 300 40032 321 40042
rect 300 40026 308 40032
rect 289 40016 308 40026
rect 196 39959 204 39989
rect 216 39959 232 39989
rect 196 39955 232 39959
rect 196 39947 226 39955
rect 300 39947 308 40016
rect 332 40023 351 40057
rect 361 40029 381 40057
rect 361 40023 375 40029
rect 400 40023 411 40067
rect 442 40062 500 40069
rect 466 40061 500 40062
rect 565 40061 599 40069
rect 497 40045 500 40061
rect 596 40045 599 40061
rect 466 40044 500 40045
rect 442 40037 500 40044
rect 565 40037 599 40045
rect 612 40028 614 40078
rect 332 39999 342 40023
rect 336 39987 342 39999
rect 224 39931 226 39947
rect 332 39919 342 39987
rect 400 39991 404 39999
rect 400 39957 408 39991
rect 434 39957 438 39991
rect 454 39975 504 39977
rect 504 39959 506 39975
rect 514 39969 530 39975
rect 532 39969 548 39975
rect 525 39959 548 39968
rect 400 39949 404 39957
rect 498 39949 506 39959
rect 504 39925 506 39949
rect 514 39939 515 39959
rect 525 39934 528 39959
rect 547 39939 548 39959
rect 557 39949 564 39959
rect 514 39925 548 39929
rect 151 39878 156 39912
rect 174 39909 246 39917
rect 256 39909 328 39917
rect 336 39911 342 39919
rect 400 39914 404 39919
rect 180 39881 185 39909
rect 174 39873 246 39881
rect 256 39873 328 39881
rect 332 39879 336 39909
rect 400 39880 438 39914
rect 224 39843 226 39859
rect 196 39835 226 39843
rect 196 39831 232 39835
rect 196 39801 204 39831
rect 216 39801 232 39831
rect 224 39754 226 39801
rect 300 39774 308 39843
rect 332 39841 342 39879
rect 400 39871 404 39880
rect 454 39865 504 39867
rect 494 39861 548 39865
rect 494 39856 514 39861
rect 504 39841 506 39856
rect 336 39829 342 39841
rect 289 39764 308 39774
rect 300 39758 308 39764
rect 332 39795 342 39829
rect 400 39833 404 39841
rect 400 39799 408 39833
rect 434 39799 438 39833
rect 498 39831 506 39841
rect 514 39831 515 39851
rect 504 39815 506 39831
rect 525 39822 528 39856
rect 547 39831 548 39851
rect 557 39831 564 39841
rect 514 39815 530 39821
rect 532 39815 548 39821
rect 332 39767 373 39795
rect 332 39761 351 39767
rect 107 39707 119 39741
rect 129 39707 149 39741
rect 196 39720 204 39754
rect 216 39720 232 39754
rect 244 39748 257 39754
rect 278 39748 291 39758
rect 244 39724 291 39748
rect 300 39748 321 39758
rect 336 39751 351 39761
rect 300 39724 329 39748
rect 332 39733 351 39751
rect 361 39761 375 39767
rect 400 39761 411 39799
rect 562 39762 612 39764
rect 361 39733 381 39761
rect 400 39733 409 39761
rect 466 39753 497 39761
rect 565 39753 596 39761
rect 442 39746 500 39753
rect 466 39745 500 39746
rect 565 39745 599 39753
rect 244 39720 257 39724
rect 42 39641 46 39675
rect 72 39641 76 39675
rect 42 39594 76 39598
rect 42 39579 46 39594
rect 72 39579 76 39594
rect 38 39561 80 39579
rect 16 39555 102 39561
rect 144 39555 148 39707
rect 174 39683 181 39711
rect 224 39673 226 39720
rect 300 39711 308 39724
rect 278 39700 305 39711
rect 332 39683 342 39733
rect 400 39713 404 39733
rect 497 39729 500 39745
rect 596 39729 599 39745
rect 466 39728 500 39729
rect 442 39721 500 39728
rect 565 39721 599 39729
rect 612 39712 614 39762
rect 256 39673 328 39681
rect 336 39675 342 39683
rect 400 39675 404 39683
rect 196 39643 204 39673
rect 216 39643 232 39673
rect 196 39639 232 39643
rect 196 39631 226 39639
rect 224 39615 226 39631
rect 332 39603 336 39671
rect 400 39641 408 39675
rect 434 39641 438 39675
rect 454 39659 504 39661
rect 504 39643 506 39659
rect 514 39653 530 39659
rect 532 39653 548 39659
rect 525 39643 548 39652
rect 400 39633 404 39641
rect 498 39633 506 39643
rect 504 39609 506 39633
rect 514 39623 515 39643
rect 525 39618 528 39643
rect 547 39623 548 39643
rect 557 39633 564 39643
rect 514 39609 548 39613
rect 400 39603 442 39604
rect 174 39593 246 39601
rect 400 39596 404 39603
rect 295 39562 300 39596
rect 324 39562 329 39596
rect 367 39579 438 39596
rect 367 39562 442 39579
rect 400 39561 442 39562
rect 378 39555 464 39561
rect 38 39539 80 39555
rect 400 39539 442 39555
rect -25 39525 25 39527
rect 42 39525 76 39539
rect 404 39525 438 39539
rect 455 39525 505 39527
rect 557 39525 607 39527
rect 16 39517 102 39525
rect 378 39517 464 39525
rect 8 39483 17 39517
rect 18 39515 51 39517
rect 80 39515 100 39517
rect 18 39483 100 39515
rect 380 39515 404 39517
rect 429 39515 438 39517
rect 442 39515 462 39517
rect 16 39475 102 39483
rect 42 39459 76 39475
rect 16 39439 38 39445
rect 42 39436 76 39440
rect 80 39439 102 39445
rect 42 39406 46 39436
rect 72 39406 76 39436
rect 42 39325 46 39359
rect 72 39325 76 39359
rect -25 39288 25 39290
rect -8 39280 14 39287
rect -8 39279 17 39280
rect 25 39279 27 39288
rect -12 39272 38 39279
rect -12 39271 34 39272
rect -12 39267 8 39271
rect 0 39255 8 39267
rect 14 39255 34 39271
rect 0 39254 34 39255
rect 0 39247 38 39254
rect 14 39246 17 39247
rect 25 39238 27 39247
rect 42 39218 45 39308
rect 69 39293 80 39325
rect 107 39293 143 39321
rect 144 39293 148 39513
rect 332 39445 336 39513
rect 380 39483 462 39515
rect 463 39483 472 39517
rect 480 39483 497 39517
rect 378 39475 464 39483
rect 505 39475 507 39525
rect 514 39483 548 39517
rect 565 39483 582 39517
rect 607 39475 609 39525
rect 404 39459 438 39475
rect 400 39445 442 39446
rect 378 39439 404 39445
rect 442 39439 464 39445
rect 400 39438 404 39439
rect 174 39399 246 39407
rect 295 39404 300 39438
rect 324 39404 329 39438
rect 224 39369 226 39385
rect 196 39361 226 39369
rect 332 39367 336 39435
rect 367 39404 438 39438
rect 400 39397 404 39404
rect 454 39391 504 39393
rect 494 39387 548 39391
rect 494 39382 514 39387
rect 504 39367 506 39382
rect 196 39357 232 39361
rect 196 39327 204 39357
rect 216 39327 232 39357
rect 400 39359 404 39367
rect 107 39287 119 39293
rect 109 39259 119 39287
rect 129 39259 149 39293
rect 174 39289 181 39319
rect 224 39280 226 39327
rect 256 39319 328 39327
rect 332 39325 336 39355
rect 400 39325 408 39359
rect 434 39325 438 39359
rect 498 39357 506 39367
rect 514 39357 515 39377
rect 504 39341 506 39357
rect 525 39348 528 39382
rect 547 39357 548 39377
rect 557 39357 564 39367
rect 514 39341 530 39347
rect 532 39341 548 39347
rect 278 39289 305 39300
rect 42 39167 46 39201
rect 72 39167 76 39201
rect 38 39129 80 39130
rect 42 39088 76 39122
rect 79 39088 113 39122
rect 42 39009 46 39043
rect 72 39009 76 39043
rect -25 38972 25 38974
rect -8 38964 14 38971
rect -8 38963 17 38964
rect 25 38963 27 38972
rect -12 38956 38 38963
rect -12 38955 34 38956
rect -12 38951 8 38955
rect 0 38939 8 38951
rect 14 38939 34 38955
rect 0 38938 34 38939
rect 0 38931 38 38938
rect 14 38930 17 38931
rect 25 38922 27 38931
rect 42 38902 45 38992
rect 71 38961 80 38989
rect 69 38923 80 38961
rect 144 38951 148 39259
rect 196 39246 204 39280
rect 216 39246 232 39280
rect 244 39276 257 39280
rect 300 39276 308 39289
rect 332 39287 342 39325
rect 400 39317 404 39325
rect 336 39277 342 39287
rect 244 39252 291 39276
rect 244 39246 257 39252
rect 224 39199 226 39246
rect 278 39242 291 39252
rect 300 39252 329 39276
rect 332 39267 342 39277
rect 400 39277 409 39305
rect 562 39288 612 39290
rect 466 39279 497 39287
rect 565 39279 596 39287
rect 300 39242 321 39252
rect 300 39236 308 39242
rect 289 39226 308 39236
rect 196 39169 204 39199
rect 216 39169 232 39199
rect 196 39165 232 39169
rect 196 39157 226 39165
rect 300 39157 308 39226
rect 332 39233 351 39267
rect 361 39239 381 39267
rect 361 39233 375 39239
rect 400 39233 411 39277
rect 442 39272 500 39279
rect 466 39271 500 39272
rect 565 39271 599 39279
rect 497 39255 500 39271
rect 596 39255 599 39271
rect 466 39254 500 39255
rect 442 39247 500 39254
rect 565 39247 599 39255
rect 612 39238 614 39288
rect 332 39209 342 39233
rect 336 39197 342 39209
rect 224 39141 226 39157
rect 332 39129 342 39197
rect 400 39201 404 39209
rect 400 39167 408 39201
rect 434 39167 438 39201
rect 454 39185 504 39187
rect 504 39169 506 39185
rect 514 39179 530 39185
rect 532 39179 548 39185
rect 525 39169 548 39178
rect 400 39159 404 39167
rect 498 39159 506 39169
rect 504 39135 506 39159
rect 514 39149 515 39169
rect 525 39144 528 39169
rect 547 39149 548 39169
rect 557 39159 564 39169
rect 514 39135 548 39139
rect 151 39088 156 39122
rect 174 39119 246 39127
rect 256 39119 328 39127
rect 336 39121 342 39129
rect 400 39124 404 39129
rect 180 39091 185 39119
rect 174 39083 246 39091
rect 256 39083 328 39091
rect 332 39089 336 39119
rect 400 39090 438 39124
rect 224 39053 226 39069
rect 196 39045 226 39053
rect 196 39041 232 39045
rect 196 39011 204 39041
rect 216 39011 232 39041
rect 224 38964 226 39011
rect 300 38984 308 39053
rect 332 39051 342 39089
rect 400 39081 404 39090
rect 454 39075 504 39077
rect 494 39071 548 39075
rect 494 39066 514 39071
rect 504 39051 506 39066
rect 336 39039 342 39051
rect 289 38974 308 38984
rect 300 38968 308 38974
rect 332 39005 342 39039
rect 400 39043 404 39051
rect 400 39009 408 39043
rect 434 39009 438 39043
rect 498 39041 506 39051
rect 514 39041 515 39061
rect 504 39025 506 39041
rect 525 39032 528 39066
rect 547 39041 548 39061
rect 557 39041 564 39051
rect 514 39025 530 39031
rect 532 39025 548 39031
rect 332 38977 373 39005
rect 332 38971 351 38977
rect 107 38917 119 38951
rect 129 38917 149 38951
rect 196 38930 204 38964
rect 216 38930 232 38964
rect 244 38958 257 38964
rect 278 38958 291 38968
rect 244 38934 291 38958
rect 300 38958 321 38968
rect 336 38961 351 38971
rect 300 38934 329 38958
rect 332 38943 351 38961
rect 361 38971 375 38977
rect 400 38971 411 39009
rect 562 38972 612 38974
rect 361 38943 381 38971
rect 400 38943 409 38971
rect 466 38963 497 38971
rect 565 38963 596 38971
rect 442 38956 500 38963
rect 466 38955 500 38956
rect 565 38955 599 38963
rect 244 38930 257 38934
rect 42 38851 46 38885
rect 72 38851 76 38885
rect 42 38804 76 38808
rect 42 38789 46 38804
rect 72 38789 76 38804
rect 38 38771 80 38789
rect 16 38765 102 38771
rect 144 38765 148 38917
rect 174 38893 181 38921
rect 224 38883 226 38930
rect 300 38921 308 38934
rect 278 38910 305 38921
rect 332 38893 342 38943
rect 400 38923 404 38943
rect 497 38939 500 38955
rect 596 38939 599 38955
rect 466 38938 500 38939
rect 442 38931 500 38938
rect 565 38931 599 38939
rect 612 38922 614 38972
rect 256 38883 328 38891
rect 336 38885 342 38893
rect 400 38885 404 38893
rect 196 38853 204 38883
rect 216 38853 232 38883
rect 196 38849 232 38853
rect 196 38841 226 38849
rect 224 38825 226 38841
rect 332 38813 336 38881
rect 400 38851 408 38885
rect 434 38851 438 38885
rect 454 38869 504 38871
rect 504 38853 506 38869
rect 514 38863 530 38869
rect 532 38863 548 38869
rect 525 38853 548 38862
rect 400 38843 404 38851
rect 498 38843 506 38853
rect 504 38819 506 38843
rect 514 38833 515 38853
rect 525 38828 528 38853
rect 547 38833 548 38853
rect 557 38843 564 38853
rect 514 38819 548 38823
rect 400 38813 442 38814
rect 174 38803 246 38811
rect 400 38806 404 38813
rect 295 38772 300 38806
rect 324 38772 329 38806
rect 367 38789 438 38806
rect 367 38772 442 38789
rect 400 38771 442 38772
rect 378 38765 464 38771
rect 38 38749 80 38765
rect 400 38749 442 38765
rect -25 38735 25 38737
rect 42 38735 76 38749
rect 404 38735 438 38749
rect 455 38735 505 38737
rect 557 38735 607 38737
rect 16 38727 102 38735
rect 378 38727 464 38735
rect 8 38693 17 38727
rect 18 38725 51 38727
rect 80 38725 100 38727
rect 18 38693 100 38725
rect 380 38725 404 38727
rect 429 38725 438 38727
rect 442 38725 462 38727
rect 16 38685 102 38693
rect 42 38669 76 38685
rect 16 38649 38 38655
rect 42 38646 76 38650
rect 80 38649 102 38655
rect 42 38616 46 38646
rect 72 38616 76 38646
rect 42 38535 46 38569
rect 72 38535 76 38569
rect -25 38498 25 38500
rect -8 38490 14 38497
rect -8 38489 17 38490
rect 25 38489 27 38498
rect -12 38482 38 38489
rect -12 38481 34 38482
rect -12 38477 8 38481
rect 0 38465 8 38477
rect 14 38465 34 38481
rect 0 38464 34 38465
rect 0 38457 38 38464
rect 14 38456 17 38457
rect 25 38448 27 38457
rect 42 38428 45 38518
rect 69 38503 80 38535
rect 107 38503 143 38531
rect 144 38503 148 38723
rect 332 38655 336 38723
rect 380 38693 462 38725
rect 463 38693 472 38727
rect 480 38693 497 38727
rect 378 38685 464 38693
rect 505 38685 507 38735
rect 514 38693 548 38727
rect 565 38693 582 38727
rect 607 38685 609 38735
rect 404 38669 438 38685
rect 400 38655 442 38656
rect 378 38649 404 38655
rect 442 38649 464 38655
rect 400 38648 404 38649
rect 174 38609 246 38617
rect 295 38614 300 38648
rect 324 38614 329 38648
rect 224 38579 226 38595
rect 196 38571 226 38579
rect 332 38577 336 38645
rect 367 38614 438 38648
rect 400 38607 404 38614
rect 454 38601 504 38603
rect 494 38597 548 38601
rect 494 38592 514 38597
rect 504 38577 506 38592
rect 196 38567 232 38571
rect 196 38537 204 38567
rect 216 38537 232 38567
rect 400 38569 404 38577
rect 107 38497 119 38503
rect 109 38469 119 38497
rect 129 38469 149 38503
rect 174 38499 181 38529
rect 224 38490 226 38537
rect 256 38529 328 38537
rect 332 38535 336 38565
rect 400 38535 408 38569
rect 434 38535 438 38569
rect 498 38567 506 38577
rect 514 38567 515 38587
rect 504 38551 506 38567
rect 525 38558 528 38592
rect 547 38567 548 38587
rect 557 38567 564 38577
rect 514 38551 530 38557
rect 532 38551 548 38557
rect 278 38499 305 38510
rect 42 38377 46 38411
rect 72 38377 76 38411
rect 38 38339 80 38340
rect 42 38298 76 38332
rect 79 38298 113 38332
rect 42 38219 46 38253
rect 72 38219 76 38253
rect -25 38182 25 38184
rect -8 38174 14 38181
rect -8 38173 17 38174
rect 25 38173 27 38182
rect -12 38166 38 38173
rect -12 38165 34 38166
rect -12 38161 8 38165
rect 0 38149 8 38161
rect 14 38149 34 38165
rect 0 38148 34 38149
rect 0 38141 38 38148
rect 14 38140 17 38141
rect 25 38132 27 38141
rect 42 38112 45 38202
rect 71 38171 80 38199
rect 69 38133 80 38171
rect 144 38161 148 38469
rect 196 38456 204 38490
rect 216 38456 232 38490
rect 244 38486 257 38490
rect 300 38486 308 38499
rect 332 38497 342 38535
rect 400 38527 404 38535
rect 336 38487 342 38497
rect 244 38462 291 38486
rect 244 38456 257 38462
rect 224 38409 226 38456
rect 278 38452 291 38462
rect 300 38462 329 38486
rect 332 38477 342 38487
rect 400 38487 409 38515
rect 562 38498 612 38500
rect 466 38489 497 38497
rect 565 38489 596 38497
rect 300 38452 321 38462
rect 300 38446 308 38452
rect 289 38436 308 38446
rect 196 38379 204 38409
rect 216 38379 232 38409
rect 196 38375 232 38379
rect 196 38367 226 38375
rect 300 38367 308 38436
rect 332 38443 351 38477
rect 361 38449 381 38477
rect 361 38443 375 38449
rect 400 38443 411 38487
rect 442 38482 500 38489
rect 466 38481 500 38482
rect 565 38481 599 38489
rect 497 38465 500 38481
rect 596 38465 599 38481
rect 466 38464 500 38465
rect 442 38457 500 38464
rect 565 38457 599 38465
rect 612 38448 614 38498
rect 332 38419 342 38443
rect 336 38407 342 38419
rect 224 38351 226 38367
rect 332 38339 342 38407
rect 400 38411 404 38419
rect 400 38377 408 38411
rect 434 38377 438 38411
rect 454 38395 504 38397
rect 504 38379 506 38395
rect 514 38389 530 38395
rect 532 38389 548 38395
rect 525 38379 548 38388
rect 400 38369 404 38377
rect 498 38369 506 38379
rect 504 38345 506 38369
rect 514 38359 515 38379
rect 525 38354 528 38379
rect 547 38359 548 38379
rect 557 38369 564 38379
rect 514 38345 548 38349
rect 151 38298 156 38332
rect 174 38329 246 38337
rect 256 38329 328 38337
rect 336 38331 342 38339
rect 400 38334 404 38339
rect 180 38301 185 38329
rect 174 38293 246 38301
rect 256 38293 328 38301
rect 332 38299 336 38329
rect 400 38300 438 38334
rect 224 38263 226 38279
rect 196 38255 226 38263
rect 196 38251 232 38255
rect 196 38221 204 38251
rect 216 38221 232 38251
rect 224 38174 226 38221
rect 300 38194 308 38263
rect 332 38261 342 38299
rect 400 38291 404 38300
rect 454 38285 504 38287
rect 494 38281 548 38285
rect 494 38276 514 38281
rect 504 38261 506 38276
rect 336 38249 342 38261
rect 289 38184 308 38194
rect 300 38178 308 38184
rect 332 38215 342 38249
rect 400 38253 404 38261
rect 400 38219 408 38253
rect 434 38219 438 38253
rect 498 38251 506 38261
rect 514 38251 515 38271
rect 504 38235 506 38251
rect 525 38242 528 38276
rect 547 38251 548 38271
rect 557 38251 564 38261
rect 514 38235 530 38241
rect 532 38235 548 38241
rect 332 38187 373 38215
rect 332 38181 351 38187
rect 107 38127 119 38161
rect 129 38127 149 38161
rect 196 38140 204 38174
rect 216 38140 232 38174
rect 244 38168 257 38174
rect 278 38168 291 38178
rect 244 38144 291 38168
rect 300 38168 321 38178
rect 336 38171 351 38181
rect 300 38144 329 38168
rect 332 38153 351 38171
rect 361 38181 375 38187
rect 400 38181 411 38219
rect 562 38182 612 38184
rect 361 38153 381 38181
rect 400 38153 409 38181
rect 466 38173 497 38181
rect 565 38173 596 38181
rect 442 38166 500 38173
rect 466 38165 500 38166
rect 565 38165 599 38173
rect 244 38140 257 38144
rect 42 38061 46 38095
rect 72 38061 76 38095
rect 42 38014 76 38018
rect 42 37999 46 38014
rect 72 37999 76 38014
rect 38 37981 80 37999
rect 16 37975 102 37981
rect 144 37975 148 38127
rect 174 38103 181 38131
rect 224 38093 226 38140
rect 300 38131 308 38144
rect 278 38120 305 38131
rect 332 38103 342 38153
rect 400 38133 404 38153
rect 497 38149 500 38165
rect 596 38149 599 38165
rect 466 38148 500 38149
rect 442 38141 500 38148
rect 565 38141 599 38149
rect 612 38132 614 38182
rect 256 38093 328 38101
rect 336 38095 342 38103
rect 400 38095 404 38103
rect 196 38063 204 38093
rect 216 38063 232 38093
rect 196 38059 232 38063
rect 196 38051 226 38059
rect 224 38035 226 38051
rect 332 38023 336 38091
rect 400 38061 408 38095
rect 434 38061 438 38095
rect 454 38079 504 38081
rect 504 38063 506 38079
rect 514 38073 530 38079
rect 532 38073 548 38079
rect 525 38063 548 38072
rect 400 38053 404 38061
rect 498 38053 506 38063
rect 504 38029 506 38053
rect 514 38043 515 38063
rect 525 38038 528 38063
rect 547 38043 548 38063
rect 557 38053 564 38063
rect 514 38029 548 38033
rect 400 38023 442 38024
rect 174 38013 246 38021
rect 400 38016 404 38023
rect 295 37982 300 38016
rect 324 37982 329 38016
rect 367 37999 438 38016
rect 367 37982 442 37999
rect 400 37981 442 37982
rect 378 37975 464 37981
rect 38 37959 80 37975
rect 400 37959 442 37975
rect -25 37945 25 37947
rect 42 37945 76 37959
rect 404 37945 438 37959
rect 455 37945 505 37947
rect 557 37945 607 37947
rect 16 37937 102 37945
rect 378 37937 464 37945
rect 8 37903 17 37937
rect 18 37935 51 37937
rect 80 37935 100 37937
rect 18 37903 100 37935
rect 380 37935 404 37937
rect 429 37935 438 37937
rect 442 37935 462 37937
rect 16 37895 102 37903
rect 42 37879 76 37895
rect 16 37859 38 37865
rect 42 37856 76 37860
rect 80 37859 102 37865
rect 42 37826 46 37856
rect 72 37826 76 37856
rect 42 37745 46 37779
rect 72 37745 76 37779
rect -25 37708 25 37710
rect -8 37700 14 37707
rect -8 37699 17 37700
rect 25 37699 27 37708
rect -12 37692 38 37699
rect -12 37691 34 37692
rect -12 37687 8 37691
rect 0 37675 8 37687
rect 14 37675 34 37691
rect 0 37674 34 37675
rect 0 37667 38 37674
rect 14 37666 17 37667
rect 25 37658 27 37667
rect 42 37638 45 37728
rect 69 37713 80 37745
rect 107 37713 143 37741
rect 144 37713 148 37933
rect 332 37865 336 37933
rect 380 37903 462 37935
rect 463 37903 472 37937
rect 480 37903 497 37937
rect 378 37895 464 37903
rect 505 37895 507 37945
rect 514 37903 548 37937
rect 565 37903 582 37937
rect 607 37895 609 37945
rect 404 37879 438 37895
rect 400 37865 442 37866
rect 378 37859 404 37865
rect 442 37859 464 37865
rect 400 37858 404 37859
rect 174 37819 246 37827
rect 295 37824 300 37858
rect 324 37824 329 37858
rect 224 37789 226 37805
rect 196 37781 226 37789
rect 332 37787 336 37855
rect 367 37824 438 37858
rect 400 37817 404 37824
rect 454 37811 504 37813
rect 494 37807 548 37811
rect 494 37802 514 37807
rect 504 37787 506 37802
rect 196 37777 232 37781
rect 196 37747 204 37777
rect 216 37747 232 37777
rect 400 37779 404 37787
rect 107 37707 119 37713
rect 109 37679 119 37707
rect 129 37679 149 37713
rect 174 37709 181 37739
rect 224 37700 226 37747
rect 256 37739 328 37747
rect 332 37745 336 37775
rect 400 37745 408 37779
rect 434 37745 438 37779
rect 498 37777 506 37787
rect 514 37777 515 37797
rect 504 37761 506 37777
rect 525 37768 528 37802
rect 547 37777 548 37797
rect 557 37777 564 37787
rect 514 37761 530 37767
rect 532 37761 548 37767
rect 278 37709 305 37720
rect 42 37587 46 37621
rect 72 37587 76 37621
rect 38 37549 80 37550
rect 42 37508 76 37542
rect 79 37508 113 37542
rect 42 37429 46 37463
rect 72 37429 76 37463
rect -25 37392 25 37394
rect -8 37384 14 37391
rect -8 37383 17 37384
rect 25 37383 27 37392
rect -12 37376 38 37383
rect -12 37375 34 37376
rect -12 37371 8 37375
rect 0 37359 8 37371
rect 14 37359 34 37375
rect 0 37358 34 37359
rect 0 37351 38 37358
rect 14 37350 17 37351
rect 25 37342 27 37351
rect 42 37322 45 37412
rect 71 37381 80 37409
rect 69 37343 80 37381
rect 144 37371 148 37679
rect 196 37666 204 37700
rect 216 37666 232 37700
rect 244 37696 257 37700
rect 300 37696 308 37709
rect 332 37707 342 37745
rect 400 37737 404 37745
rect 336 37697 342 37707
rect 244 37672 291 37696
rect 244 37666 257 37672
rect 224 37619 226 37666
rect 278 37662 291 37672
rect 300 37672 329 37696
rect 332 37687 342 37697
rect 400 37697 409 37725
rect 562 37708 612 37710
rect 466 37699 497 37707
rect 565 37699 596 37707
rect 300 37662 321 37672
rect 300 37656 308 37662
rect 289 37646 308 37656
rect 196 37589 204 37619
rect 216 37589 232 37619
rect 196 37585 232 37589
rect 196 37577 226 37585
rect 300 37577 308 37646
rect 332 37653 351 37687
rect 361 37659 381 37687
rect 361 37653 375 37659
rect 400 37653 411 37697
rect 442 37692 500 37699
rect 466 37691 500 37692
rect 565 37691 599 37699
rect 497 37675 500 37691
rect 596 37675 599 37691
rect 466 37674 500 37675
rect 442 37667 500 37674
rect 565 37667 599 37675
rect 612 37658 614 37708
rect 332 37629 342 37653
rect 336 37617 342 37629
rect 224 37561 226 37577
rect 332 37549 342 37617
rect 400 37621 404 37629
rect 400 37587 408 37621
rect 434 37587 438 37621
rect 454 37605 504 37607
rect 504 37589 506 37605
rect 514 37599 530 37605
rect 532 37599 548 37605
rect 525 37589 548 37598
rect 400 37579 404 37587
rect 498 37579 506 37589
rect 504 37555 506 37579
rect 514 37569 515 37589
rect 525 37564 528 37589
rect 547 37569 548 37589
rect 557 37579 564 37589
rect 514 37555 548 37559
rect 151 37508 156 37542
rect 174 37539 246 37547
rect 256 37539 328 37547
rect 336 37541 342 37549
rect 400 37544 404 37549
rect 180 37511 185 37539
rect 174 37503 246 37511
rect 256 37503 328 37511
rect 332 37509 336 37539
rect 400 37510 438 37544
rect 224 37473 226 37489
rect 196 37465 226 37473
rect 196 37461 232 37465
rect 196 37431 204 37461
rect 216 37431 232 37461
rect 224 37384 226 37431
rect 300 37404 308 37473
rect 332 37471 342 37509
rect 400 37501 404 37510
rect 454 37495 504 37497
rect 494 37491 548 37495
rect 494 37486 514 37491
rect 504 37471 506 37486
rect 336 37459 342 37471
rect 289 37394 308 37404
rect 300 37388 308 37394
rect 332 37425 342 37459
rect 400 37463 404 37471
rect 400 37429 408 37463
rect 434 37429 438 37463
rect 498 37461 506 37471
rect 514 37461 515 37481
rect 504 37445 506 37461
rect 525 37452 528 37486
rect 547 37461 548 37481
rect 557 37461 564 37471
rect 514 37445 530 37451
rect 532 37445 548 37451
rect 332 37397 373 37425
rect 332 37391 351 37397
rect 107 37337 119 37371
rect 129 37337 149 37371
rect 196 37350 204 37384
rect 216 37350 232 37384
rect 244 37378 257 37384
rect 278 37378 291 37388
rect 244 37354 291 37378
rect 300 37378 321 37388
rect 336 37381 351 37391
rect 300 37354 329 37378
rect 332 37363 351 37381
rect 361 37391 375 37397
rect 400 37391 411 37429
rect 562 37392 612 37394
rect 361 37363 381 37391
rect 400 37363 409 37391
rect 466 37383 497 37391
rect 565 37383 596 37391
rect 442 37376 500 37383
rect 466 37375 500 37376
rect 565 37375 599 37383
rect 244 37350 257 37354
rect 42 37271 46 37305
rect 72 37271 76 37305
rect 42 37224 76 37228
rect 42 37209 46 37224
rect 72 37209 76 37224
rect 38 37191 80 37209
rect 16 37185 102 37191
rect 144 37185 148 37337
rect 174 37313 181 37341
rect 224 37303 226 37350
rect 300 37341 308 37354
rect 278 37330 305 37341
rect 332 37313 342 37363
rect 400 37343 404 37363
rect 497 37359 500 37375
rect 596 37359 599 37375
rect 466 37358 500 37359
rect 442 37351 500 37358
rect 565 37351 599 37359
rect 612 37342 614 37392
rect 256 37303 328 37311
rect 336 37305 342 37313
rect 400 37305 404 37313
rect 196 37273 204 37303
rect 216 37273 232 37303
rect 196 37269 232 37273
rect 196 37261 226 37269
rect 224 37245 226 37261
rect 332 37233 336 37301
rect 400 37271 408 37305
rect 434 37271 438 37305
rect 454 37289 504 37291
rect 504 37273 506 37289
rect 514 37283 530 37289
rect 532 37283 548 37289
rect 525 37273 548 37282
rect 400 37263 404 37271
rect 498 37263 506 37273
rect 504 37239 506 37263
rect 514 37253 515 37273
rect 525 37248 528 37273
rect 547 37253 548 37273
rect 557 37263 564 37273
rect 514 37239 548 37243
rect 400 37233 442 37234
rect 174 37223 246 37231
rect 400 37226 404 37233
rect 295 37192 300 37226
rect 324 37192 329 37226
rect 367 37209 438 37226
rect 367 37192 442 37209
rect 400 37191 442 37192
rect 378 37185 464 37191
rect 38 37169 80 37185
rect 400 37169 442 37185
rect -25 37155 25 37157
rect 42 37155 76 37169
rect 404 37155 438 37169
rect 455 37155 505 37157
rect 557 37155 607 37157
rect 16 37147 102 37155
rect 378 37147 464 37155
rect 8 37113 17 37147
rect 18 37145 51 37147
rect 80 37145 100 37147
rect 18 37113 100 37145
rect 380 37145 404 37147
rect 429 37145 438 37147
rect 442 37145 462 37147
rect 16 37105 102 37113
rect 42 37089 76 37105
rect 16 37069 38 37075
rect 42 37066 76 37070
rect 80 37069 102 37075
rect 42 37036 46 37066
rect 72 37036 76 37066
rect 42 36955 46 36989
rect 72 36955 76 36989
rect -25 36918 25 36920
rect -8 36910 14 36917
rect -8 36909 17 36910
rect 25 36909 27 36918
rect -12 36902 38 36909
rect -12 36901 34 36902
rect -12 36897 8 36901
rect 0 36885 8 36897
rect 14 36885 34 36901
rect 0 36884 34 36885
rect 0 36877 38 36884
rect 14 36876 17 36877
rect 25 36868 27 36877
rect 42 36848 45 36938
rect 69 36923 80 36955
rect 107 36923 143 36951
rect 144 36923 148 37143
rect 332 37075 336 37143
rect 380 37113 462 37145
rect 463 37113 472 37147
rect 480 37113 497 37147
rect 378 37105 464 37113
rect 505 37105 507 37155
rect 514 37113 548 37147
rect 565 37113 582 37147
rect 607 37105 609 37155
rect 404 37089 438 37105
rect 400 37075 442 37076
rect 378 37069 404 37075
rect 442 37069 464 37075
rect 400 37068 404 37069
rect 174 37029 246 37037
rect 295 37034 300 37068
rect 324 37034 329 37068
rect 224 36999 226 37015
rect 196 36991 226 36999
rect 332 36997 336 37065
rect 367 37034 438 37068
rect 400 37027 404 37034
rect 454 37021 504 37023
rect 494 37017 548 37021
rect 494 37012 514 37017
rect 504 36997 506 37012
rect 196 36987 232 36991
rect 196 36957 204 36987
rect 216 36957 232 36987
rect 400 36989 404 36997
rect 107 36917 119 36923
rect 109 36889 119 36917
rect 129 36889 149 36923
rect 174 36919 181 36949
rect 224 36910 226 36957
rect 256 36949 328 36957
rect 332 36955 336 36985
rect 400 36955 408 36989
rect 434 36955 438 36989
rect 498 36987 506 36997
rect 514 36987 515 37007
rect 504 36971 506 36987
rect 525 36978 528 37012
rect 547 36987 548 37007
rect 557 36987 564 36997
rect 514 36971 530 36977
rect 532 36971 548 36977
rect 278 36919 305 36930
rect 42 36797 46 36831
rect 72 36797 76 36831
rect 38 36759 80 36760
rect 42 36718 76 36752
rect 79 36718 113 36752
rect 42 36639 46 36673
rect 72 36639 76 36673
rect -25 36602 25 36604
rect -8 36594 14 36601
rect -8 36593 17 36594
rect 25 36593 27 36602
rect -12 36586 38 36593
rect -12 36585 34 36586
rect -12 36581 8 36585
rect 0 36569 8 36581
rect 14 36569 34 36585
rect 0 36568 34 36569
rect 0 36561 38 36568
rect 14 36560 17 36561
rect 25 36552 27 36561
rect 42 36532 45 36622
rect 71 36591 80 36619
rect 69 36553 80 36591
rect 144 36581 148 36889
rect 196 36876 204 36910
rect 216 36876 232 36910
rect 244 36906 257 36910
rect 300 36906 308 36919
rect 332 36917 342 36955
rect 400 36947 404 36955
rect 336 36907 342 36917
rect 244 36882 291 36906
rect 244 36876 257 36882
rect 224 36829 226 36876
rect 278 36872 291 36882
rect 300 36882 329 36906
rect 332 36897 342 36907
rect 400 36907 409 36935
rect 562 36918 612 36920
rect 466 36909 497 36917
rect 565 36909 596 36917
rect 300 36872 321 36882
rect 300 36866 308 36872
rect 289 36856 308 36866
rect 196 36799 204 36829
rect 216 36799 232 36829
rect 196 36795 232 36799
rect 196 36787 226 36795
rect 300 36787 308 36856
rect 332 36863 351 36897
rect 361 36869 381 36897
rect 361 36863 375 36869
rect 400 36863 411 36907
rect 442 36902 500 36909
rect 466 36901 500 36902
rect 565 36901 599 36909
rect 497 36885 500 36901
rect 596 36885 599 36901
rect 466 36884 500 36885
rect 442 36877 500 36884
rect 565 36877 599 36885
rect 612 36868 614 36918
rect 332 36839 342 36863
rect 336 36827 342 36839
rect 224 36771 226 36787
rect 332 36759 342 36827
rect 400 36831 404 36839
rect 400 36797 408 36831
rect 434 36797 438 36831
rect 454 36815 504 36817
rect 504 36799 506 36815
rect 514 36809 530 36815
rect 532 36809 548 36815
rect 525 36799 548 36808
rect 400 36789 404 36797
rect 498 36789 506 36799
rect 504 36765 506 36789
rect 514 36779 515 36799
rect 525 36774 528 36799
rect 547 36779 548 36799
rect 557 36789 564 36799
rect 514 36765 548 36769
rect 151 36718 156 36752
rect 174 36749 246 36757
rect 256 36749 328 36757
rect 336 36751 342 36759
rect 400 36754 404 36759
rect 180 36721 185 36749
rect 174 36713 246 36721
rect 256 36713 328 36721
rect 332 36719 336 36749
rect 400 36720 438 36754
rect 224 36683 226 36699
rect 196 36675 226 36683
rect 196 36671 232 36675
rect 196 36641 204 36671
rect 216 36641 232 36671
rect 224 36594 226 36641
rect 300 36614 308 36683
rect 332 36681 342 36719
rect 400 36711 404 36720
rect 454 36705 504 36707
rect 494 36701 548 36705
rect 494 36696 514 36701
rect 504 36681 506 36696
rect 336 36669 342 36681
rect 289 36604 308 36614
rect 300 36598 308 36604
rect 332 36635 342 36669
rect 400 36673 404 36681
rect 400 36639 408 36673
rect 434 36639 438 36673
rect 498 36671 506 36681
rect 514 36671 515 36691
rect 504 36655 506 36671
rect 525 36662 528 36696
rect 547 36671 548 36691
rect 557 36671 564 36681
rect 514 36655 530 36661
rect 532 36655 548 36661
rect 332 36607 373 36635
rect 332 36601 351 36607
rect 107 36547 119 36581
rect 129 36547 149 36581
rect 196 36560 204 36594
rect 216 36560 232 36594
rect 244 36588 257 36594
rect 278 36588 291 36598
rect 244 36564 291 36588
rect 300 36588 321 36598
rect 336 36591 351 36601
rect 300 36564 329 36588
rect 332 36573 351 36591
rect 361 36601 375 36607
rect 400 36601 411 36639
rect 562 36602 612 36604
rect 361 36573 381 36601
rect 400 36573 409 36601
rect 466 36593 497 36601
rect 565 36593 596 36601
rect 442 36586 500 36593
rect 466 36585 500 36586
rect 565 36585 599 36593
rect 244 36560 257 36564
rect 42 36481 46 36515
rect 72 36481 76 36515
rect 42 36434 76 36438
rect 42 36419 46 36434
rect 72 36419 76 36434
rect 38 36401 80 36419
rect 16 36395 102 36401
rect 144 36395 148 36547
rect 174 36523 181 36551
rect 224 36513 226 36560
rect 300 36551 308 36564
rect 278 36540 305 36551
rect 332 36523 342 36573
rect 400 36553 404 36573
rect 497 36569 500 36585
rect 596 36569 599 36585
rect 466 36568 500 36569
rect 442 36561 500 36568
rect 565 36561 599 36569
rect 612 36552 614 36602
rect 256 36513 328 36521
rect 336 36515 342 36523
rect 400 36515 404 36523
rect 196 36483 204 36513
rect 216 36483 232 36513
rect 196 36479 232 36483
rect 196 36471 226 36479
rect 224 36455 226 36471
rect 332 36443 336 36511
rect 400 36481 408 36515
rect 434 36481 438 36515
rect 454 36499 504 36501
rect 504 36483 506 36499
rect 514 36493 530 36499
rect 532 36493 548 36499
rect 525 36483 548 36492
rect 400 36473 404 36481
rect 498 36473 506 36483
rect 504 36449 506 36473
rect 514 36463 515 36483
rect 525 36458 528 36483
rect 547 36463 548 36483
rect 557 36473 564 36483
rect 514 36449 548 36453
rect 400 36443 442 36444
rect 174 36433 246 36441
rect 400 36436 404 36443
rect 295 36402 300 36436
rect 324 36402 329 36436
rect 367 36419 438 36436
rect 367 36402 442 36419
rect 400 36401 442 36402
rect 378 36395 464 36401
rect 38 36379 80 36395
rect 400 36379 442 36395
rect -25 36365 25 36367
rect 42 36365 76 36379
rect 404 36365 438 36379
rect 455 36365 505 36367
rect 557 36365 607 36367
rect 16 36357 102 36365
rect 378 36357 464 36365
rect 8 36323 17 36357
rect 18 36355 51 36357
rect 80 36355 100 36357
rect 18 36323 100 36355
rect 380 36355 404 36357
rect 429 36355 438 36357
rect 442 36355 462 36357
rect 16 36315 102 36323
rect 42 36299 76 36315
rect 16 36279 38 36285
rect 42 36276 76 36280
rect 80 36279 102 36285
rect 42 36246 46 36276
rect 72 36246 76 36276
rect 42 36165 46 36199
rect 72 36165 76 36199
rect -25 36128 25 36130
rect -8 36120 14 36127
rect -8 36119 17 36120
rect 25 36119 27 36128
rect -12 36112 38 36119
rect -12 36111 34 36112
rect -12 36107 8 36111
rect 0 36095 8 36107
rect 14 36095 34 36111
rect 0 36094 34 36095
rect 0 36087 38 36094
rect 14 36086 17 36087
rect 25 36078 27 36087
rect 42 36058 45 36148
rect 69 36133 80 36165
rect 107 36133 143 36161
rect 144 36133 148 36353
rect 332 36285 336 36353
rect 380 36323 462 36355
rect 463 36323 472 36357
rect 480 36323 497 36357
rect 378 36315 464 36323
rect 505 36315 507 36365
rect 514 36323 548 36357
rect 565 36323 582 36357
rect 607 36315 609 36365
rect 404 36299 438 36315
rect 400 36285 442 36286
rect 378 36279 404 36285
rect 442 36279 464 36285
rect 400 36278 404 36279
rect 174 36239 246 36247
rect 295 36244 300 36278
rect 324 36244 329 36278
rect 224 36209 226 36225
rect 196 36201 226 36209
rect 332 36207 336 36275
rect 367 36244 438 36278
rect 400 36237 404 36244
rect 454 36231 504 36233
rect 494 36227 548 36231
rect 494 36222 514 36227
rect 504 36207 506 36222
rect 196 36197 232 36201
rect 196 36167 204 36197
rect 216 36167 232 36197
rect 400 36199 404 36207
rect 107 36127 119 36133
rect 109 36099 119 36127
rect 129 36099 149 36133
rect 174 36129 181 36159
rect 224 36120 226 36167
rect 256 36159 328 36167
rect 332 36165 336 36195
rect 400 36165 408 36199
rect 434 36165 438 36199
rect 498 36197 506 36207
rect 514 36197 515 36217
rect 504 36181 506 36197
rect 525 36188 528 36222
rect 547 36197 548 36217
rect 557 36197 564 36207
rect 514 36181 530 36187
rect 532 36181 548 36187
rect 278 36129 305 36140
rect 42 36007 46 36041
rect 72 36007 76 36041
rect 38 35969 80 35970
rect 42 35928 76 35962
rect 79 35928 113 35962
rect 42 35849 46 35883
rect 72 35849 76 35883
rect -25 35812 25 35814
rect -8 35804 14 35811
rect -8 35803 17 35804
rect 25 35803 27 35812
rect -12 35796 38 35803
rect -12 35795 34 35796
rect -12 35791 8 35795
rect 0 35779 8 35791
rect 14 35779 34 35795
rect 0 35778 34 35779
rect 0 35771 38 35778
rect 14 35770 17 35771
rect 25 35762 27 35771
rect 42 35742 45 35832
rect 71 35801 80 35829
rect 69 35763 80 35801
rect 144 35791 148 36099
rect 196 36086 204 36120
rect 216 36086 232 36120
rect 244 36116 257 36120
rect 300 36116 308 36129
rect 332 36127 342 36165
rect 400 36157 404 36165
rect 336 36117 342 36127
rect 244 36092 291 36116
rect 244 36086 257 36092
rect 224 36039 226 36086
rect 278 36082 291 36092
rect 300 36092 329 36116
rect 332 36107 342 36117
rect 400 36117 409 36145
rect 562 36128 612 36130
rect 466 36119 497 36127
rect 565 36119 596 36127
rect 300 36082 321 36092
rect 300 36076 308 36082
rect 289 36066 308 36076
rect 196 36009 204 36039
rect 216 36009 232 36039
rect 196 36005 232 36009
rect 196 35997 226 36005
rect 300 35997 308 36066
rect 332 36073 351 36107
rect 361 36079 381 36107
rect 361 36073 375 36079
rect 400 36073 411 36117
rect 442 36112 500 36119
rect 466 36111 500 36112
rect 565 36111 599 36119
rect 497 36095 500 36111
rect 596 36095 599 36111
rect 466 36094 500 36095
rect 442 36087 500 36094
rect 565 36087 599 36095
rect 612 36078 614 36128
rect 332 36049 342 36073
rect 336 36037 342 36049
rect 224 35981 226 35997
rect 332 35969 342 36037
rect 400 36041 404 36049
rect 400 36007 408 36041
rect 434 36007 438 36041
rect 454 36025 504 36027
rect 504 36009 506 36025
rect 514 36019 530 36025
rect 532 36019 548 36025
rect 525 36009 548 36018
rect 400 35999 404 36007
rect 498 35999 506 36009
rect 504 35975 506 35999
rect 514 35989 515 36009
rect 525 35984 528 36009
rect 547 35989 548 36009
rect 557 35999 564 36009
rect 514 35975 548 35979
rect 151 35928 156 35962
rect 174 35959 246 35967
rect 256 35959 328 35967
rect 336 35961 342 35969
rect 400 35964 404 35969
rect 180 35931 185 35959
rect 174 35923 246 35931
rect 256 35923 328 35931
rect 332 35929 336 35959
rect 400 35930 438 35964
rect 224 35893 226 35909
rect 196 35885 226 35893
rect 196 35881 232 35885
rect 196 35851 204 35881
rect 216 35851 232 35881
rect 224 35804 226 35851
rect 300 35824 308 35893
rect 332 35891 342 35929
rect 400 35921 404 35930
rect 454 35915 504 35917
rect 494 35911 548 35915
rect 494 35906 514 35911
rect 504 35891 506 35906
rect 336 35879 342 35891
rect 289 35814 308 35824
rect 300 35808 308 35814
rect 332 35845 342 35879
rect 400 35883 404 35891
rect 400 35849 408 35883
rect 434 35849 438 35883
rect 498 35881 506 35891
rect 514 35881 515 35901
rect 504 35865 506 35881
rect 525 35872 528 35906
rect 547 35881 548 35901
rect 557 35881 564 35891
rect 514 35865 530 35871
rect 532 35865 548 35871
rect 332 35817 373 35845
rect 332 35811 351 35817
rect 107 35757 119 35791
rect 129 35757 149 35791
rect 196 35770 204 35804
rect 216 35770 232 35804
rect 244 35798 257 35804
rect 278 35798 291 35808
rect 244 35774 291 35798
rect 300 35798 321 35808
rect 336 35801 351 35811
rect 300 35774 329 35798
rect 332 35783 351 35801
rect 361 35811 375 35817
rect 400 35811 411 35849
rect 562 35812 612 35814
rect 361 35783 381 35811
rect 400 35783 409 35811
rect 466 35803 497 35811
rect 565 35803 596 35811
rect 442 35796 500 35803
rect 466 35795 500 35796
rect 565 35795 599 35803
rect 244 35770 257 35774
rect 42 35691 46 35725
rect 72 35691 76 35725
rect 42 35644 76 35648
rect 42 35629 46 35644
rect 72 35629 76 35644
rect 38 35611 80 35629
rect 16 35605 102 35611
rect 144 35605 148 35757
rect 174 35733 181 35761
rect 224 35723 226 35770
rect 300 35761 308 35774
rect 278 35750 305 35761
rect 332 35733 342 35783
rect 400 35763 404 35783
rect 497 35779 500 35795
rect 596 35779 599 35795
rect 466 35778 500 35779
rect 442 35771 500 35778
rect 565 35771 599 35779
rect 612 35762 614 35812
rect 256 35723 328 35731
rect 336 35725 342 35733
rect 400 35725 404 35733
rect 196 35693 204 35723
rect 216 35693 232 35723
rect 196 35689 232 35693
rect 196 35681 226 35689
rect 224 35665 226 35681
rect 332 35653 336 35721
rect 400 35691 408 35725
rect 434 35691 438 35725
rect 454 35709 504 35711
rect 504 35693 506 35709
rect 514 35703 530 35709
rect 532 35703 548 35709
rect 525 35693 548 35702
rect 400 35683 404 35691
rect 498 35683 506 35693
rect 504 35659 506 35683
rect 514 35673 515 35693
rect 525 35668 528 35693
rect 547 35673 548 35693
rect 557 35683 564 35693
rect 514 35659 548 35663
rect 400 35653 442 35654
rect 174 35643 246 35651
rect 400 35646 404 35653
rect 295 35612 300 35646
rect 324 35612 329 35646
rect 367 35629 438 35646
rect 367 35612 442 35629
rect 400 35611 442 35612
rect 378 35605 464 35611
rect 38 35589 80 35605
rect 400 35589 442 35605
rect -25 35575 25 35577
rect 42 35575 76 35589
rect 404 35575 438 35589
rect 455 35575 505 35577
rect 557 35575 607 35577
rect 16 35567 102 35575
rect 378 35567 464 35575
rect 8 35533 17 35567
rect 18 35565 51 35567
rect 80 35565 100 35567
rect 18 35533 100 35565
rect 380 35565 404 35567
rect 429 35565 438 35567
rect 442 35565 462 35567
rect 16 35525 102 35533
rect 42 35509 76 35525
rect 16 35489 38 35495
rect 42 35486 76 35490
rect 80 35489 102 35495
rect 42 35456 46 35486
rect 72 35456 76 35486
rect 42 35375 46 35409
rect 72 35375 76 35409
rect -25 35338 25 35340
rect -8 35330 14 35337
rect -8 35329 17 35330
rect 25 35329 27 35338
rect -12 35322 38 35329
rect -12 35321 34 35322
rect -12 35317 8 35321
rect 0 35305 8 35317
rect 14 35305 34 35321
rect 0 35304 34 35305
rect 0 35297 38 35304
rect 14 35296 17 35297
rect 25 35288 27 35297
rect 42 35268 45 35358
rect 69 35343 80 35375
rect 107 35343 143 35371
rect 144 35343 148 35563
rect 332 35495 336 35563
rect 380 35533 462 35565
rect 463 35533 472 35567
rect 480 35533 497 35567
rect 378 35525 464 35533
rect 505 35525 507 35575
rect 514 35533 548 35567
rect 565 35533 582 35567
rect 607 35525 609 35575
rect 404 35509 438 35525
rect 400 35495 442 35496
rect 378 35489 404 35495
rect 442 35489 464 35495
rect 400 35488 404 35489
rect 174 35449 246 35457
rect 295 35454 300 35488
rect 324 35454 329 35488
rect 224 35419 226 35435
rect 196 35411 226 35419
rect 332 35417 336 35485
rect 367 35454 438 35488
rect 400 35447 404 35454
rect 454 35441 504 35443
rect 494 35437 548 35441
rect 494 35432 514 35437
rect 504 35417 506 35432
rect 196 35407 232 35411
rect 196 35377 204 35407
rect 216 35377 232 35407
rect 400 35409 404 35417
rect 107 35337 119 35343
rect 109 35309 119 35337
rect 129 35309 149 35343
rect 174 35339 181 35369
rect 224 35330 226 35377
rect 256 35369 328 35377
rect 332 35375 336 35405
rect 400 35375 408 35409
rect 434 35375 438 35409
rect 498 35407 506 35417
rect 514 35407 515 35427
rect 504 35391 506 35407
rect 525 35398 528 35432
rect 547 35407 548 35427
rect 557 35407 564 35417
rect 514 35391 530 35397
rect 532 35391 548 35397
rect 278 35339 305 35350
rect 42 35217 46 35251
rect 72 35217 76 35251
rect 38 35179 80 35180
rect 42 35138 76 35172
rect 79 35138 113 35172
rect 42 35059 46 35093
rect 72 35059 76 35093
rect -25 35022 25 35024
rect -8 35014 14 35021
rect -8 35013 17 35014
rect 25 35013 27 35022
rect -12 35006 38 35013
rect -12 35005 34 35006
rect -12 35001 8 35005
rect 0 34989 8 35001
rect 14 34989 34 35005
rect 0 34988 34 34989
rect 0 34981 38 34988
rect 14 34980 17 34981
rect 25 34972 27 34981
rect 42 34952 45 35042
rect 71 35011 80 35039
rect 69 34973 80 35011
rect 144 35001 148 35309
rect 196 35296 204 35330
rect 216 35296 232 35330
rect 244 35326 257 35330
rect 300 35326 308 35339
rect 332 35337 342 35375
rect 400 35367 404 35375
rect 336 35327 342 35337
rect 244 35302 291 35326
rect 244 35296 257 35302
rect 224 35249 226 35296
rect 278 35292 291 35302
rect 300 35302 329 35326
rect 332 35317 342 35327
rect 400 35327 409 35355
rect 562 35338 612 35340
rect 466 35329 497 35337
rect 565 35329 596 35337
rect 300 35292 321 35302
rect 300 35286 308 35292
rect 289 35276 308 35286
rect 196 35219 204 35249
rect 216 35219 232 35249
rect 196 35215 232 35219
rect 196 35207 226 35215
rect 300 35207 308 35276
rect 332 35283 351 35317
rect 361 35289 381 35317
rect 361 35283 375 35289
rect 400 35283 411 35327
rect 442 35322 500 35329
rect 466 35321 500 35322
rect 565 35321 599 35329
rect 497 35305 500 35321
rect 596 35305 599 35321
rect 466 35304 500 35305
rect 442 35297 500 35304
rect 565 35297 599 35305
rect 612 35288 614 35338
rect 332 35259 342 35283
rect 336 35247 342 35259
rect 224 35191 226 35207
rect 332 35179 342 35247
rect 400 35251 404 35259
rect 400 35217 408 35251
rect 434 35217 438 35251
rect 454 35235 504 35237
rect 504 35219 506 35235
rect 514 35229 530 35235
rect 532 35229 548 35235
rect 525 35219 548 35228
rect 400 35209 404 35217
rect 498 35209 506 35219
rect 504 35185 506 35209
rect 514 35199 515 35219
rect 525 35194 528 35219
rect 547 35199 548 35219
rect 557 35209 564 35219
rect 514 35185 548 35189
rect 151 35138 156 35172
rect 174 35169 246 35177
rect 256 35169 328 35177
rect 336 35171 342 35179
rect 400 35174 404 35179
rect 180 35141 185 35169
rect 174 35133 246 35141
rect 256 35133 328 35141
rect 332 35139 336 35169
rect 400 35140 438 35174
rect 224 35103 226 35119
rect 196 35095 226 35103
rect 196 35091 232 35095
rect 196 35061 204 35091
rect 216 35061 232 35091
rect 224 35014 226 35061
rect 300 35034 308 35103
rect 332 35101 342 35139
rect 400 35131 404 35140
rect 454 35125 504 35127
rect 494 35121 548 35125
rect 494 35116 514 35121
rect 504 35101 506 35116
rect 336 35089 342 35101
rect 289 35024 308 35034
rect 300 35018 308 35024
rect 332 35055 342 35089
rect 400 35093 404 35101
rect 400 35059 408 35093
rect 434 35059 438 35093
rect 498 35091 506 35101
rect 514 35091 515 35111
rect 504 35075 506 35091
rect 525 35082 528 35116
rect 547 35091 548 35111
rect 557 35091 564 35101
rect 514 35075 530 35081
rect 532 35075 548 35081
rect 332 35027 373 35055
rect 332 35021 351 35027
rect 107 34967 119 35001
rect 129 34967 149 35001
rect 196 34980 204 35014
rect 216 34980 232 35014
rect 244 35008 257 35014
rect 278 35008 291 35018
rect 244 34984 291 35008
rect 300 35008 321 35018
rect 336 35011 351 35021
rect 300 34984 329 35008
rect 332 34993 351 35011
rect 361 35021 375 35027
rect 400 35021 411 35059
rect 562 35022 612 35024
rect 361 34993 381 35021
rect 400 34993 409 35021
rect 466 35013 497 35021
rect 565 35013 596 35021
rect 442 35006 500 35013
rect 466 35005 500 35006
rect 565 35005 599 35013
rect 244 34980 257 34984
rect 42 34901 46 34935
rect 72 34901 76 34935
rect 42 34854 76 34858
rect 42 34839 46 34854
rect 72 34839 76 34854
rect 38 34821 80 34839
rect 16 34815 102 34821
rect 144 34815 148 34967
rect 174 34943 181 34971
rect 224 34933 226 34980
rect 300 34971 308 34984
rect 278 34960 305 34971
rect 332 34943 342 34993
rect 400 34973 404 34993
rect 497 34989 500 35005
rect 596 34989 599 35005
rect 466 34988 500 34989
rect 442 34981 500 34988
rect 565 34981 599 34989
rect 612 34972 614 35022
rect 256 34933 328 34941
rect 336 34935 342 34943
rect 400 34935 404 34943
rect 196 34903 204 34933
rect 216 34903 232 34933
rect 196 34899 232 34903
rect 196 34891 226 34899
rect 224 34875 226 34891
rect 332 34863 336 34931
rect 400 34901 408 34935
rect 434 34901 438 34935
rect 454 34919 504 34921
rect 504 34903 506 34919
rect 514 34913 530 34919
rect 532 34913 548 34919
rect 525 34903 548 34912
rect 400 34893 404 34901
rect 498 34893 506 34903
rect 504 34869 506 34893
rect 514 34883 515 34903
rect 525 34878 528 34903
rect 547 34883 548 34903
rect 557 34893 564 34903
rect 514 34869 548 34873
rect 400 34863 442 34864
rect 174 34853 246 34861
rect 400 34856 404 34863
rect 295 34822 300 34856
rect 324 34822 329 34856
rect 367 34839 438 34856
rect 367 34822 442 34839
rect 400 34821 442 34822
rect 378 34815 464 34821
rect 38 34799 80 34815
rect 400 34799 442 34815
rect -25 34785 25 34787
rect 42 34785 76 34799
rect 404 34785 438 34799
rect 455 34785 505 34787
rect 557 34785 607 34787
rect 16 34777 102 34785
rect 378 34777 464 34785
rect 8 34743 17 34777
rect 18 34775 51 34777
rect 80 34775 100 34777
rect 18 34743 100 34775
rect 380 34775 404 34777
rect 429 34775 438 34777
rect 442 34775 462 34777
rect 16 34735 102 34743
rect 42 34719 76 34735
rect 16 34699 38 34705
rect 42 34696 76 34700
rect 80 34699 102 34705
rect 42 34666 46 34696
rect 72 34666 76 34696
rect 42 34585 46 34619
rect 72 34585 76 34619
rect -25 34548 25 34550
rect -8 34540 14 34547
rect -8 34539 17 34540
rect 25 34539 27 34548
rect -12 34532 38 34539
rect -12 34531 34 34532
rect -12 34527 8 34531
rect 0 34515 8 34527
rect 14 34515 34 34531
rect 0 34514 34 34515
rect 0 34507 38 34514
rect 14 34506 17 34507
rect 25 34498 27 34507
rect 42 34478 45 34568
rect 69 34553 80 34585
rect 107 34553 143 34581
rect 144 34553 148 34773
rect 332 34705 336 34773
rect 380 34743 462 34775
rect 463 34743 472 34777
rect 480 34743 497 34777
rect 378 34735 464 34743
rect 505 34735 507 34785
rect 514 34743 548 34777
rect 565 34743 582 34777
rect 607 34735 609 34785
rect 404 34719 438 34735
rect 400 34705 442 34706
rect 378 34699 404 34705
rect 442 34699 464 34705
rect 400 34698 404 34699
rect 174 34659 246 34667
rect 295 34664 300 34698
rect 324 34664 329 34698
rect 224 34629 226 34645
rect 196 34621 226 34629
rect 332 34627 336 34695
rect 367 34664 438 34698
rect 400 34657 404 34664
rect 454 34651 504 34653
rect 494 34647 548 34651
rect 494 34642 514 34647
rect 504 34627 506 34642
rect 196 34617 232 34621
rect 196 34587 204 34617
rect 216 34587 232 34617
rect 400 34619 404 34627
rect 107 34547 119 34553
rect 109 34519 119 34547
rect 129 34519 149 34553
rect 174 34549 181 34579
rect 224 34540 226 34587
rect 256 34579 328 34587
rect 332 34585 336 34615
rect 400 34585 408 34619
rect 434 34585 438 34619
rect 498 34617 506 34627
rect 514 34617 515 34637
rect 504 34601 506 34617
rect 525 34608 528 34642
rect 547 34617 548 34637
rect 557 34617 564 34627
rect 514 34601 530 34607
rect 532 34601 548 34607
rect 278 34549 305 34560
rect 42 34427 46 34461
rect 72 34427 76 34461
rect 38 34389 80 34390
rect 42 34348 76 34382
rect 79 34348 113 34382
rect 42 34269 46 34303
rect 72 34269 76 34303
rect -25 34232 25 34234
rect -8 34224 14 34231
rect -8 34223 17 34224
rect 25 34223 27 34232
rect -12 34216 38 34223
rect -12 34215 34 34216
rect -12 34211 8 34215
rect 0 34199 8 34211
rect 14 34199 34 34215
rect 0 34198 34 34199
rect 0 34191 38 34198
rect 14 34190 17 34191
rect 25 34182 27 34191
rect 42 34162 45 34252
rect 71 34221 80 34249
rect 69 34183 80 34221
rect 144 34211 148 34519
rect 196 34506 204 34540
rect 216 34506 232 34540
rect 244 34536 257 34540
rect 300 34536 308 34549
rect 332 34547 342 34585
rect 400 34577 404 34585
rect 336 34537 342 34547
rect 244 34512 291 34536
rect 244 34506 257 34512
rect 224 34459 226 34506
rect 278 34502 291 34512
rect 300 34512 329 34536
rect 332 34527 342 34537
rect 400 34537 409 34565
rect 562 34548 612 34550
rect 466 34539 497 34547
rect 565 34539 596 34547
rect 300 34502 321 34512
rect 300 34496 308 34502
rect 289 34486 308 34496
rect 196 34429 204 34459
rect 216 34429 232 34459
rect 196 34425 232 34429
rect 196 34417 226 34425
rect 300 34417 308 34486
rect 332 34493 351 34527
rect 361 34499 381 34527
rect 361 34493 375 34499
rect 400 34493 411 34537
rect 442 34532 500 34539
rect 466 34531 500 34532
rect 565 34531 599 34539
rect 497 34515 500 34531
rect 596 34515 599 34531
rect 466 34514 500 34515
rect 442 34507 500 34514
rect 565 34507 599 34515
rect 612 34498 614 34548
rect 332 34469 342 34493
rect 336 34457 342 34469
rect 224 34401 226 34417
rect 332 34389 342 34457
rect 400 34461 404 34469
rect 400 34427 408 34461
rect 434 34427 438 34461
rect 454 34445 504 34447
rect 504 34429 506 34445
rect 514 34439 530 34445
rect 532 34439 548 34445
rect 525 34429 548 34438
rect 400 34419 404 34427
rect 498 34419 506 34429
rect 504 34395 506 34419
rect 514 34409 515 34429
rect 525 34404 528 34429
rect 547 34409 548 34429
rect 557 34419 564 34429
rect 514 34395 548 34399
rect 151 34348 156 34382
rect 174 34379 246 34387
rect 256 34379 328 34387
rect 336 34381 342 34389
rect 400 34384 404 34389
rect 180 34351 185 34379
rect 174 34343 246 34351
rect 256 34343 328 34351
rect 332 34349 336 34379
rect 400 34350 438 34384
rect 224 34313 226 34329
rect 196 34305 226 34313
rect 196 34301 232 34305
rect 196 34271 204 34301
rect 216 34271 232 34301
rect 224 34224 226 34271
rect 300 34244 308 34313
rect 332 34311 342 34349
rect 400 34341 404 34350
rect 454 34335 504 34337
rect 494 34331 548 34335
rect 494 34326 514 34331
rect 504 34311 506 34326
rect 336 34299 342 34311
rect 289 34234 308 34244
rect 300 34228 308 34234
rect 332 34265 342 34299
rect 400 34303 404 34311
rect 400 34269 408 34303
rect 434 34269 438 34303
rect 498 34301 506 34311
rect 514 34301 515 34321
rect 504 34285 506 34301
rect 525 34292 528 34326
rect 547 34301 548 34321
rect 557 34301 564 34311
rect 514 34285 530 34291
rect 532 34285 548 34291
rect 332 34237 373 34265
rect 332 34231 351 34237
rect 107 34177 119 34211
rect 129 34177 149 34211
rect 196 34190 204 34224
rect 216 34190 232 34224
rect 244 34218 257 34224
rect 278 34218 291 34228
rect 244 34194 291 34218
rect 300 34218 321 34228
rect 336 34221 351 34231
rect 300 34194 329 34218
rect 332 34203 351 34221
rect 361 34231 375 34237
rect 400 34231 411 34269
rect 562 34232 612 34234
rect 361 34203 381 34231
rect 400 34203 409 34231
rect 466 34223 497 34231
rect 565 34223 596 34231
rect 442 34216 500 34223
rect 466 34215 500 34216
rect 565 34215 599 34223
rect 244 34190 257 34194
rect 42 34111 46 34145
rect 72 34111 76 34145
rect 42 34064 76 34068
rect 42 34049 46 34064
rect 72 34049 76 34064
rect 38 34031 80 34049
rect 16 34025 102 34031
rect 144 34025 148 34177
rect 174 34153 181 34181
rect 224 34143 226 34190
rect 300 34181 308 34194
rect 278 34170 305 34181
rect 332 34153 342 34203
rect 400 34183 404 34203
rect 497 34199 500 34215
rect 596 34199 599 34215
rect 466 34198 500 34199
rect 442 34191 500 34198
rect 565 34191 599 34199
rect 612 34182 614 34232
rect 256 34143 328 34151
rect 336 34145 342 34153
rect 400 34145 404 34153
rect 196 34113 204 34143
rect 216 34113 232 34143
rect 196 34109 232 34113
rect 196 34101 226 34109
rect 224 34085 226 34101
rect 332 34073 336 34141
rect 400 34111 408 34145
rect 434 34111 438 34145
rect 454 34129 504 34131
rect 504 34113 506 34129
rect 514 34123 530 34129
rect 532 34123 548 34129
rect 525 34113 548 34122
rect 400 34103 404 34111
rect 498 34103 506 34113
rect 504 34079 506 34103
rect 514 34093 515 34113
rect 525 34088 528 34113
rect 547 34093 548 34113
rect 557 34103 564 34113
rect 514 34079 548 34083
rect 400 34073 442 34074
rect 174 34063 246 34071
rect 400 34066 404 34073
rect 295 34032 300 34066
rect 324 34032 329 34066
rect 367 34049 438 34066
rect 367 34032 442 34049
rect 400 34031 442 34032
rect 378 34025 464 34031
rect 38 34009 80 34025
rect 400 34009 442 34025
rect -25 33995 25 33997
rect 42 33995 76 34009
rect 404 33995 438 34009
rect 455 33995 505 33997
rect 557 33995 607 33997
rect 16 33987 102 33995
rect 378 33987 464 33995
rect 8 33953 17 33987
rect 18 33985 51 33987
rect 80 33985 100 33987
rect 18 33953 100 33985
rect 380 33985 404 33987
rect 429 33985 438 33987
rect 442 33985 462 33987
rect 16 33945 102 33953
rect 42 33929 76 33945
rect 16 33909 38 33915
rect 42 33906 76 33910
rect 80 33909 102 33915
rect 42 33876 46 33906
rect 72 33876 76 33906
rect 42 33795 46 33829
rect 72 33795 76 33829
rect -25 33758 25 33760
rect -8 33750 14 33757
rect -8 33749 17 33750
rect 25 33749 27 33758
rect -12 33742 38 33749
rect -12 33741 34 33742
rect -12 33737 8 33741
rect 0 33725 8 33737
rect 14 33725 34 33741
rect 0 33724 34 33725
rect 0 33717 38 33724
rect 14 33716 17 33717
rect 25 33708 27 33717
rect 42 33688 45 33778
rect 69 33763 80 33795
rect 107 33763 143 33791
rect 144 33763 148 33983
rect 332 33915 336 33983
rect 380 33953 462 33985
rect 463 33953 472 33987
rect 480 33953 497 33987
rect 378 33945 464 33953
rect 505 33945 507 33995
rect 514 33953 548 33987
rect 565 33953 582 33987
rect 607 33945 609 33995
rect 404 33929 438 33945
rect 400 33915 442 33916
rect 378 33909 404 33915
rect 442 33909 464 33915
rect 400 33908 404 33909
rect 174 33869 246 33877
rect 295 33874 300 33908
rect 324 33874 329 33908
rect 224 33839 226 33855
rect 196 33831 226 33839
rect 332 33837 336 33905
rect 367 33874 438 33908
rect 400 33867 404 33874
rect 454 33861 504 33863
rect 494 33857 548 33861
rect 494 33852 514 33857
rect 504 33837 506 33852
rect 196 33827 232 33831
rect 196 33797 204 33827
rect 216 33797 232 33827
rect 400 33829 404 33837
rect 107 33757 119 33763
rect 109 33729 119 33757
rect 129 33729 149 33763
rect 174 33759 181 33789
rect 224 33750 226 33797
rect 256 33789 328 33797
rect 332 33795 336 33825
rect 400 33795 408 33829
rect 434 33795 438 33829
rect 498 33827 506 33837
rect 514 33827 515 33847
rect 504 33811 506 33827
rect 525 33818 528 33852
rect 547 33827 548 33847
rect 557 33827 564 33837
rect 514 33811 530 33817
rect 532 33811 548 33817
rect 278 33759 305 33770
rect 42 33637 46 33671
rect 72 33637 76 33671
rect 38 33599 80 33600
rect 42 33558 76 33592
rect 79 33558 113 33592
rect 42 33479 46 33513
rect 72 33479 76 33513
rect -25 33442 25 33444
rect -8 33434 14 33441
rect -8 33433 17 33434
rect 25 33433 27 33442
rect -12 33426 38 33433
rect -12 33425 34 33426
rect -12 33421 8 33425
rect 0 33409 8 33421
rect 14 33409 34 33425
rect 0 33408 34 33409
rect 0 33401 38 33408
rect 14 33400 17 33401
rect 25 33392 27 33401
rect 42 33372 45 33462
rect 71 33431 80 33459
rect 69 33393 80 33431
rect 144 33421 148 33729
rect 196 33716 204 33750
rect 216 33716 232 33750
rect 244 33746 257 33750
rect 300 33746 308 33759
rect 332 33757 342 33795
rect 400 33787 404 33795
rect 336 33747 342 33757
rect 244 33722 291 33746
rect 244 33716 257 33722
rect 224 33669 226 33716
rect 278 33712 291 33722
rect 300 33722 329 33746
rect 332 33737 342 33747
rect 400 33747 409 33775
rect 562 33758 612 33760
rect 466 33749 497 33757
rect 565 33749 596 33757
rect 300 33712 321 33722
rect 300 33706 308 33712
rect 289 33696 308 33706
rect 196 33639 204 33669
rect 216 33639 232 33669
rect 196 33635 232 33639
rect 196 33627 226 33635
rect 300 33627 308 33696
rect 332 33703 351 33737
rect 361 33709 381 33737
rect 361 33703 375 33709
rect 400 33703 411 33747
rect 442 33742 500 33749
rect 466 33741 500 33742
rect 565 33741 599 33749
rect 497 33725 500 33741
rect 596 33725 599 33741
rect 466 33724 500 33725
rect 442 33717 500 33724
rect 565 33717 599 33725
rect 612 33708 614 33758
rect 332 33679 342 33703
rect 336 33667 342 33679
rect 224 33611 226 33627
rect 332 33599 342 33667
rect 400 33671 404 33679
rect 400 33637 408 33671
rect 434 33637 438 33671
rect 454 33655 504 33657
rect 504 33639 506 33655
rect 514 33649 530 33655
rect 532 33649 548 33655
rect 525 33639 548 33648
rect 400 33629 404 33637
rect 498 33629 506 33639
rect 504 33605 506 33629
rect 514 33619 515 33639
rect 525 33614 528 33639
rect 547 33619 548 33639
rect 557 33629 564 33639
rect 514 33605 548 33609
rect 151 33558 156 33592
rect 174 33589 246 33597
rect 256 33589 328 33597
rect 336 33591 342 33599
rect 400 33594 404 33599
rect 180 33561 185 33589
rect 174 33553 246 33561
rect 256 33553 328 33561
rect 332 33559 336 33589
rect 400 33560 438 33594
rect 224 33523 226 33539
rect 196 33515 226 33523
rect 196 33511 232 33515
rect 196 33481 204 33511
rect 216 33481 232 33511
rect 224 33434 226 33481
rect 300 33454 308 33523
rect 332 33521 342 33559
rect 400 33551 404 33560
rect 454 33545 504 33547
rect 494 33541 548 33545
rect 494 33536 514 33541
rect 504 33521 506 33536
rect 336 33509 342 33521
rect 289 33444 308 33454
rect 300 33438 308 33444
rect 332 33475 342 33509
rect 400 33513 404 33521
rect 400 33479 408 33513
rect 434 33479 438 33513
rect 498 33511 506 33521
rect 514 33511 515 33531
rect 504 33495 506 33511
rect 525 33502 528 33536
rect 547 33511 548 33531
rect 557 33511 564 33521
rect 514 33495 530 33501
rect 532 33495 548 33501
rect 332 33447 373 33475
rect 332 33441 351 33447
rect 107 33387 119 33421
rect 129 33387 149 33421
rect 196 33400 204 33434
rect 216 33400 232 33434
rect 244 33428 257 33434
rect 278 33428 291 33438
rect 244 33404 291 33428
rect 300 33428 321 33438
rect 336 33431 351 33441
rect 300 33404 329 33428
rect 332 33413 351 33431
rect 361 33441 375 33447
rect 400 33441 411 33479
rect 562 33442 612 33444
rect 361 33413 381 33441
rect 400 33413 409 33441
rect 466 33433 497 33441
rect 565 33433 596 33441
rect 442 33426 500 33433
rect 466 33425 500 33426
rect 565 33425 599 33433
rect 244 33400 257 33404
rect 42 33321 46 33355
rect 72 33321 76 33355
rect 42 33274 76 33278
rect 42 33259 46 33274
rect 72 33259 76 33274
rect 38 33241 80 33259
rect 16 33235 102 33241
rect 144 33235 148 33387
rect 174 33363 181 33391
rect 224 33353 226 33400
rect 300 33391 308 33404
rect 278 33380 305 33391
rect 332 33363 342 33413
rect 400 33393 404 33413
rect 497 33409 500 33425
rect 596 33409 599 33425
rect 466 33408 500 33409
rect 442 33401 500 33408
rect 565 33401 599 33409
rect 612 33392 614 33442
rect 256 33353 328 33361
rect 336 33355 342 33363
rect 400 33355 404 33363
rect 196 33323 204 33353
rect 216 33323 232 33353
rect 196 33319 232 33323
rect 196 33311 226 33319
rect 224 33295 226 33311
rect 332 33283 336 33351
rect 400 33321 408 33355
rect 434 33321 438 33355
rect 454 33339 504 33341
rect 504 33323 506 33339
rect 514 33333 530 33339
rect 532 33333 548 33339
rect 525 33323 548 33332
rect 400 33313 404 33321
rect 498 33313 506 33323
rect 504 33289 506 33313
rect 514 33303 515 33323
rect 525 33298 528 33323
rect 547 33303 548 33323
rect 557 33313 564 33323
rect 514 33289 548 33293
rect 400 33283 442 33284
rect 174 33273 246 33281
rect 400 33276 404 33283
rect 295 33242 300 33276
rect 324 33242 329 33276
rect 367 33259 438 33276
rect 367 33242 442 33259
rect 400 33241 442 33242
rect 378 33235 464 33241
rect 38 33219 80 33235
rect 400 33219 442 33235
rect -25 33205 25 33207
rect 42 33205 76 33219
rect 404 33205 438 33219
rect 455 33205 505 33207
rect 557 33205 607 33207
rect 16 33197 102 33205
rect 378 33197 464 33205
rect 8 33163 17 33197
rect 18 33195 51 33197
rect 80 33195 100 33197
rect 18 33163 100 33195
rect 380 33195 404 33197
rect 429 33195 438 33197
rect 442 33195 462 33197
rect 16 33155 102 33163
rect 42 33139 76 33155
rect 16 33119 38 33125
rect 42 33116 76 33120
rect 80 33119 102 33125
rect 42 33086 46 33116
rect 72 33086 76 33116
rect 42 33005 46 33039
rect 72 33005 76 33039
rect -25 32968 25 32970
rect -8 32960 14 32967
rect -8 32959 17 32960
rect 25 32959 27 32968
rect -12 32952 38 32959
rect -12 32951 34 32952
rect -12 32947 8 32951
rect 0 32935 8 32947
rect 14 32935 34 32951
rect 0 32934 34 32935
rect 0 32927 38 32934
rect 14 32926 17 32927
rect 25 32918 27 32927
rect 42 32898 45 32988
rect 69 32973 80 33005
rect 107 32973 143 33001
rect 144 32973 148 33193
rect 332 33125 336 33193
rect 380 33163 462 33195
rect 463 33163 472 33197
rect 480 33163 497 33197
rect 378 33155 464 33163
rect 505 33155 507 33205
rect 514 33163 548 33197
rect 565 33163 582 33197
rect 607 33155 609 33205
rect 404 33139 438 33155
rect 400 33125 442 33126
rect 378 33119 404 33125
rect 442 33119 464 33125
rect 400 33118 404 33119
rect 174 33079 246 33087
rect 295 33084 300 33118
rect 324 33084 329 33118
rect 224 33049 226 33065
rect 196 33041 226 33049
rect 332 33047 336 33115
rect 367 33084 438 33118
rect 400 33077 404 33084
rect 454 33071 504 33073
rect 494 33067 548 33071
rect 494 33062 514 33067
rect 504 33047 506 33062
rect 196 33037 232 33041
rect 196 33007 204 33037
rect 216 33007 232 33037
rect 400 33039 404 33047
rect 107 32967 119 32973
rect 109 32939 119 32967
rect 129 32939 149 32973
rect 174 32969 181 32999
rect 224 32960 226 33007
rect 256 32999 328 33007
rect 332 33005 336 33035
rect 400 33005 408 33039
rect 434 33005 438 33039
rect 498 33037 506 33047
rect 514 33037 515 33057
rect 504 33021 506 33037
rect 525 33028 528 33062
rect 547 33037 548 33057
rect 557 33037 564 33047
rect 514 33021 530 33027
rect 532 33021 548 33027
rect 278 32969 305 32980
rect 42 32847 46 32881
rect 72 32847 76 32881
rect 38 32809 80 32810
rect 42 32768 76 32802
rect 79 32768 113 32802
rect 42 32689 46 32723
rect 72 32689 76 32723
rect -25 32652 25 32654
rect -8 32644 14 32651
rect -8 32643 17 32644
rect 25 32643 27 32652
rect -12 32636 38 32643
rect -12 32635 34 32636
rect -12 32631 8 32635
rect 0 32619 8 32631
rect 14 32619 34 32635
rect 0 32618 34 32619
rect 0 32611 38 32618
rect 14 32610 17 32611
rect 25 32602 27 32611
rect 42 32582 45 32672
rect 71 32641 80 32669
rect 69 32603 80 32641
rect 144 32631 148 32939
rect 196 32926 204 32960
rect 216 32926 232 32960
rect 244 32956 257 32960
rect 300 32956 308 32969
rect 332 32967 342 33005
rect 400 32997 404 33005
rect 336 32957 342 32967
rect 244 32932 291 32956
rect 244 32926 257 32932
rect 224 32879 226 32926
rect 278 32922 291 32932
rect 300 32932 329 32956
rect 332 32947 342 32957
rect 400 32957 409 32985
rect 562 32968 612 32970
rect 466 32959 497 32967
rect 565 32959 596 32967
rect 300 32922 321 32932
rect 300 32916 308 32922
rect 289 32906 308 32916
rect 196 32849 204 32879
rect 216 32849 232 32879
rect 196 32845 232 32849
rect 196 32837 226 32845
rect 300 32837 308 32906
rect 332 32913 351 32947
rect 361 32919 381 32947
rect 361 32913 375 32919
rect 400 32913 411 32957
rect 442 32952 500 32959
rect 466 32951 500 32952
rect 565 32951 599 32959
rect 497 32935 500 32951
rect 596 32935 599 32951
rect 466 32934 500 32935
rect 442 32927 500 32934
rect 565 32927 599 32935
rect 612 32918 614 32968
rect 332 32889 342 32913
rect 336 32877 342 32889
rect 224 32821 226 32837
rect 332 32809 342 32877
rect 400 32881 404 32889
rect 400 32847 408 32881
rect 434 32847 438 32881
rect 454 32865 504 32867
rect 504 32849 506 32865
rect 514 32859 530 32865
rect 532 32859 548 32865
rect 525 32849 548 32858
rect 400 32839 404 32847
rect 498 32839 506 32849
rect 504 32815 506 32839
rect 514 32829 515 32849
rect 525 32824 528 32849
rect 547 32829 548 32849
rect 557 32839 564 32849
rect 514 32815 548 32819
rect 151 32768 156 32802
rect 174 32799 246 32807
rect 256 32799 328 32807
rect 336 32801 342 32809
rect 400 32804 404 32809
rect 180 32771 185 32799
rect 174 32763 246 32771
rect 256 32763 328 32771
rect 332 32769 336 32799
rect 400 32770 438 32804
rect 224 32733 226 32749
rect 196 32725 226 32733
rect 196 32721 232 32725
rect 196 32691 204 32721
rect 216 32691 232 32721
rect 224 32644 226 32691
rect 300 32664 308 32733
rect 332 32731 342 32769
rect 400 32761 404 32770
rect 454 32755 504 32757
rect 494 32751 548 32755
rect 494 32746 514 32751
rect 504 32731 506 32746
rect 336 32719 342 32731
rect 289 32654 308 32664
rect 300 32648 308 32654
rect 332 32685 342 32719
rect 400 32723 404 32731
rect 400 32689 408 32723
rect 434 32689 438 32723
rect 498 32721 506 32731
rect 514 32721 515 32741
rect 504 32705 506 32721
rect 525 32712 528 32746
rect 547 32721 548 32741
rect 557 32721 564 32731
rect 514 32705 530 32711
rect 532 32705 548 32711
rect 332 32657 373 32685
rect 332 32651 351 32657
rect 107 32597 119 32631
rect 129 32597 149 32631
rect 196 32610 204 32644
rect 216 32610 232 32644
rect 244 32638 257 32644
rect 278 32638 291 32648
rect 244 32614 291 32638
rect 300 32638 321 32648
rect 336 32641 351 32651
rect 300 32614 329 32638
rect 332 32623 351 32641
rect 361 32651 375 32657
rect 400 32651 411 32689
rect 562 32652 612 32654
rect 361 32623 381 32651
rect 400 32623 409 32651
rect 466 32643 497 32651
rect 565 32643 596 32651
rect 442 32636 500 32643
rect 466 32635 500 32636
rect 565 32635 599 32643
rect 244 32610 257 32614
rect 42 32531 46 32565
rect 72 32531 76 32565
rect 42 32484 76 32488
rect 42 32469 46 32484
rect 72 32469 76 32484
rect 38 32451 80 32469
rect 16 32445 102 32451
rect 144 32445 148 32597
rect 174 32573 181 32601
rect 224 32563 226 32610
rect 300 32601 308 32614
rect 278 32590 305 32601
rect 332 32573 342 32623
rect 400 32603 404 32623
rect 497 32619 500 32635
rect 596 32619 599 32635
rect 466 32618 500 32619
rect 442 32611 500 32618
rect 565 32611 599 32619
rect 612 32602 614 32652
rect 256 32563 328 32571
rect 336 32565 342 32573
rect 400 32565 404 32573
rect 196 32533 204 32563
rect 216 32533 232 32563
rect 196 32529 232 32533
rect 196 32521 226 32529
rect 224 32505 226 32521
rect 332 32493 336 32561
rect 400 32531 408 32565
rect 434 32531 438 32565
rect 454 32549 504 32551
rect 504 32533 506 32549
rect 514 32543 530 32549
rect 532 32543 548 32549
rect 525 32533 548 32542
rect 400 32523 404 32531
rect 498 32523 506 32533
rect 504 32499 506 32523
rect 514 32513 515 32533
rect 525 32508 528 32533
rect 547 32513 548 32533
rect 557 32523 564 32533
rect 514 32499 548 32503
rect 400 32493 442 32494
rect 174 32483 246 32491
rect 400 32486 404 32493
rect 295 32452 300 32486
rect 324 32452 329 32486
rect 367 32469 438 32486
rect 367 32452 442 32469
rect 400 32451 442 32452
rect 378 32445 464 32451
rect 38 32429 80 32445
rect 400 32429 442 32445
rect -25 32415 25 32417
rect 42 32415 76 32429
rect 404 32415 438 32429
rect 455 32415 505 32417
rect 557 32415 607 32417
rect 16 32407 102 32415
rect 378 32407 464 32415
rect 8 32373 17 32407
rect 18 32405 51 32407
rect 80 32405 100 32407
rect 18 32373 100 32405
rect 380 32405 404 32407
rect 429 32405 438 32407
rect 442 32405 462 32407
rect 16 32365 102 32373
rect 42 32349 76 32365
rect 16 32329 38 32335
rect 42 32326 76 32330
rect 80 32329 102 32335
rect 42 32296 46 32326
rect 72 32296 76 32326
rect 42 32215 46 32249
rect 72 32215 76 32249
rect -25 32178 25 32180
rect -8 32170 14 32177
rect -8 32169 17 32170
rect 25 32169 27 32178
rect -12 32162 38 32169
rect -12 32161 34 32162
rect -12 32157 8 32161
rect 0 32145 8 32157
rect 14 32145 34 32161
rect 0 32144 34 32145
rect 0 32137 38 32144
rect 14 32136 17 32137
rect 25 32128 27 32137
rect 42 32108 45 32198
rect 69 32183 80 32215
rect 107 32183 143 32211
rect 144 32183 148 32403
rect 332 32335 336 32403
rect 380 32373 462 32405
rect 463 32373 472 32407
rect 480 32373 497 32407
rect 378 32365 464 32373
rect 505 32365 507 32415
rect 514 32373 548 32407
rect 565 32373 582 32407
rect 607 32365 609 32415
rect 404 32349 438 32365
rect 400 32335 442 32336
rect 378 32329 404 32335
rect 442 32329 464 32335
rect 400 32328 404 32329
rect 174 32289 246 32297
rect 295 32294 300 32328
rect 324 32294 329 32328
rect 224 32259 226 32275
rect 196 32251 226 32259
rect 332 32257 336 32325
rect 367 32294 438 32328
rect 400 32287 404 32294
rect 454 32281 504 32283
rect 494 32277 548 32281
rect 494 32272 514 32277
rect 504 32257 506 32272
rect 196 32247 232 32251
rect 196 32217 204 32247
rect 216 32217 232 32247
rect 400 32249 404 32257
rect 107 32177 119 32183
rect 109 32149 119 32177
rect 129 32149 149 32183
rect 174 32179 181 32209
rect 224 32170 226 32217
rect 256 32209 328 32217
rect 332 32215 336 32245
rect 400 32215 408 32249
rect 434 32215 438 32249
rect 498 32247 506 32257
rect 514 32247 515 32267
rect 504 32231 506 32247
rect 525 32238 528 32272
rect 547 32247 548 32267
rect 557 32247 564 32257
rect 514 32231 530 32237
rect 532 32231 548 32237
rect 278 32179 305 32190
rect 42 32057 46 32091
rect 72 32057 76 32091
rect 38 32019 80 32020
rect 42 31978 76 32012
rect 79 31978 113 32012
rect 42 31899 46 31933
rect 72 31899 76 31933
rect -25 31862 25 31864
rect -8 31854 14 31861
rect -8 31853 17 31854
rect 25 31853 27 31862
rect -12 31846 38 31853
rect -12 31845 34 31846
rect -12 31841 8 31845
rect 0 31829 8 31841
rect 14 31829 34 31845
rect 0 31828 34 31829
rect 0 31821 38 31828
rect 14 31820 17 31821
rect 25 31812 27 31821
rect 42 31792 45 31882
rect 71 31851 80 31879
rect 69 31813 80 31851
rect 144 31841 148 32149
rect 196 32136 204 32170
rect 216 32136 232 32170
rect 244 32166 257 32170
rect 300 32166 308 32179
rect 332 32177 342 32215
rect 400 32207 404 32215
rect 336 32167 342 32177
rect 244 32142 291 32166
rect 244 32136 257 32142
rect 224 32089 226 32136
rect 278 32132 291 32142
rect 300 32142 329 32166
rect 332 32157 342 32167
rect 400 32167 409 32195
rect 562 32178 612 32180
rect 466 32169 497 32177
rect 565 32169 596 32177
rect 300 32132 321 32142
rect 300 32126 308 32132
rect 289 32116 308 32126
rect 196 32059 204 32089
rect 216 32059 232 32089
rect 196 32055 232 32059
rect 196 32047 226 32055
rect 300 32047 308 32116
rect 332 32123 351 32157
rect 361 32129 381 32157
rect 361 32123 375 32129
rect 400 32123 411 32167
rect 442 32162 500 32169
rect 466 32161 500 32162
rect 565 32161 599 32169
rect 497 32145 500 32161
rect 596 32145 599 32161
rect 466 32144 500 32145
rect 442 32137 500 32144
rect 565 32137 599 32145
rect 612 32128 614 32178
rect 332 32099 342 32123
rect 336 32087 342 32099
rect 224 32031 226 32047
rect 332 32019 342 32087
rect 400 32091 404 32099
rect 400 32057 408 32091
rect 434 32057 438 32091
rect 454 32075 504 32077
rect 504 32059 506 32075
rect 514 32069 530 32075
rect 532 32069 548 32075
rect 525 32059 548 32068
rect 400 32049 404 32057
rect 498 32049 506 32059
rect 504 32025 506 32049
rect 514 32039 515 32059
rect 525 32034 528 32059
rect 547 32039 548 32059
rect 557 32049 564 32059
rect 514 32025 548 32029
rect 151 31978 156 32012
rect 174 32009 246 32017
rect 256 32009 328 32017
rect 336 32011 342 32019
rect 400 32014 404 32019
rect 180 31981 185 32009
rect 174 31973 246 31981
rect 256 31973 328 31981
rect 332 31979 336 32009
rect 400 31980 438 32014
rect 224 31943 226 31959
rect 196 31935 226 31943
rect 196 31931 232 31935
rect 196 31901 204 31931
rect 216 31901 232 31931
rect 224 31854 226 31901
rect 300 31874 308 31943
rect 332 31941 342 31979
rect 400 31971 404 31980
rect 454 31965 504 31967
rect 494 31961 548 31965
rect 494 31956 514 31961
rect 504 31941 506 31956
rect 336 31929 342 31941
rect 289 31864 308 31874
rect 300 31858 308 31864
rect 332 31895 342 31929
rect 400 31933 404 31941
rect 400 31899 408 31933
rect 434 31899 438 31933
rect 498 31931 506 31941
rect 514 31931 515 31951
rect 504 31915 506 31931
rect 525 31922 528 31956
rect 547 31931 548 31951
rect 557 31931 564 31941
rect 514 31915 530 31921
rect 532 31915 548 31921
rect 332 31867 373 31895
rect 332 31861 351 31867
rect 107 31807 119 31841
rect 129 31807 149 31841
rect 196 31820 204 31854
rect 216 31820 232 31854
rect 244 31848 257 31854
rect 278 31848 291 31858
rect 244 31824 291 31848
rect 300 31848 321 31858
rect 336 31851 351 31861
rect 300 31824 329 31848
rect 332 31833 351 31851
rect 361 31861 375 31867
rect 400 31861 411 31899
rect 562 31862 612 31864
rect 361 31833 381 31861
rect 400 31833 409 31861
rect 466 31853 497 31861
rect 565 31853 596 31861
rect 442 31846 500 31853
rect 466 31845 500 31846
rect 565 31845 599 31853
rect 244 31820 257 31824
rect 42 31741 46 31775
rect 72 31741 76 31775
rect 42 31694 76 31698
rect 42 31679 46 31694
rect 72 31679 76 31694
rect 38 31661 80 31679
rect 16 31655 102 31661
rect 144 31655 148 31807
rect 174 31783 181 31811
rect 224 31773 226 31820
rect 300 31811 308 31824
rect 278 31800 305 31811
rect 332 31783 342 31833
rect 400 31813 404 31833
rect 497 31829 500 31845
rect 596 31829 599 31845
rect 466 31828 500 31829
rect 442 31821 500 31828
rect 565 31821 599 31829
rect 612 31812 614 31862
rect 256 31773 328 31781
rect 336 31775 342 31783
rect 400 31775 404 31783
rect 196 31743 204 31773
rect 216 31743 232 31773
rect 196 31739 232 31743
rect 196 31731 226 31739
rect 224 31715 226 31731
rect 332 31703 336 31771
rect 400 31741 408 31775
rect 434 31741 438 31775
rect 454 31759 504 31761
rect 504 31743 506 31759
rect 514 31753 530 31759
rect 532 31753 548 31759
rect 525 31743 548 31752
rect 400 31733 404 31741
rect 498 31733 506 31743
rect 504 31709 506 31733
rect 514 31723 515 31743
rect 525 31718 528 31743
rect 547 31723 548 31743
rect 557 31733 564 31743
rect 514 31709 548 31713
rect 400 31703 442 31704
rect 174 31693 246 31701
rect 400 31696 404 31703
rect 295 31662 300 31696
rect 324 31662 329 31696
rect 367 31679 438 31696
rect 367 31662 442 31679
rect 400 31661 442 31662
rect 378 31655 464 31661
rect 38 31639 80 31655
rect 400 31639 442 31655
rect -25 31625 25 31627
rect 42 31625 76 31639
rect 404 31625 438 31639
rect 455 31625 505 31627
rect 557 31625 607 31627
rect 16 31617 102 31625
rect 378 31617 464 31625
rect 8 31583 17 31617
rect 18 31615 51 31617
rect 80 31615 100 31617
rect 18 31583 100 31615
rect 380 31615 404 31617
rect 429 31615 438 31617
rect 442 31615 462 31617
rect 16 31575 102 31583
rect 42 31559 76 31575
rect 16 31539 38 31545
rect 42 31536 76 31540
rect 80 31539 102 31545
rect 42 31506 46 31536
rect 72 31506 76 31536
rect 42 31425 46 31459
rect 72 31425 76 31459
rect -25 31388 25 31390
rect -8 31380 14 31387
rect -8 31379 17 31380
rect 25 31379 27 31388
rect -12 31372 38 31379
rect -12 31371 34 31372
rect -12 31367 8 31371
rect 0 31355 8 31367
rect 14 31355 34 31371
rect 0 31354 34 31355
rect 0 31347 38 31354
rect 14 31346 17 31347
rect 25 31338 27 31347
rect 42 31318 45 31408
rect 69 31393 80 31425
rect 107 31393 143 31421
rect 144 31393 148 31613
rect 332 31545 336 31613
rect 380 31583 462 31615
rect 463 31583 472 31617
rect 480 31583 497 31617
rect 378 31575 464 31583
rect 505 31575 507 31625
rect 514 31583 548 31617
rect 565 31583 582 31617
rect 607 31575 609 31625
rect 404 31559 438 31575
rect 400 31545 442 31546
rect 378 31539 404 31545
rect 442 31539 464 31545
rect 400 31538 404 31539
rect 174 31499 246 31507
rect 295 31504 300 31538
rect 324 31504 329 31538
rect 224 31469 226 31485
rect 196 31461 226 31469
rect 332 31467 336 31535
rect 367 31504 438 31538
rect 400 31497 404 31504
rect 454 31491 504 31493
rect 494 31487 548 31491
rect 494 31482 514 31487
rect 504 31467 506 31482
rect 196 31457 232 31461
rect 196 31427 204 31457
rect 216 31427 232 31457
rect 400 31459 404 31467
rect 107 31387 119 31393
rect 109 31359 119 31387
rect 129 31359 149 31393
rect 174 31389 181 31419
rect 224 31380 226 31427
rect 256 31419 328 31427
rect 332 31425 336 31455
rect 400 31425 408 31459
rect 434 31425 438 31459
rect 498 31457 506 31467
rect 514 31457 515 31477
rect 504 31441 506 31457
rect 525 31448 528 31482
rect 547 31457 548 31477
rect 557 31457 564 31467
rect 514 31441 530 31447
rect 532 31441 548 31447
rect 278 31389 305 31400
rect 42 31267 46 31301
rect 72 31267 76 31301
rect 38 31229 80 31230
rect 42 31188 76 31222
rect 79 31188 113 31222
rect 42 31109 46 31143
rect 72 31109 76 31143
rect -25 31072 25 31074
rect -8 31064 14 31071
rect -8 31063 17 31064
rect 25 31063 27 31072
rect -12 31056 38 31063
rect -12 31055 34 31056
rect -12 31051 8 31055
rect 0 31039 8 31051
rect 14 31039 34 31055
rect 0 31038 34 31039
rect 0 31031 38 31038
rect 14 31030 17 31031
rect 25 31022 27 31031
rect 42 31002 45 31092
rect 71 31061 80 31089
rect 69 31023 80 31061
rect 144 31051 148 31359
rect 196 31346 204 31380
rect 216 31346 232 31380
rect 244 31376 257 31380
rect 300 31376 308 31389
rect 332 31387 342 31425
rect 400 31417 404 31425
rect 336 31377 342 31387
rect 244 31352 291 31376
rect 244 31346 257 31352
rect 224 31299 226 31346
rect 278 31342 291 31352
rect 300 31352 329 31376
rect 332 31367 342 31377
rect 400 31377 409 31405
rect 562 31388 612 31390
rect 466 31379 497 31387
rect 565 31379 596 31387
rect 300 31342 321 31352
rect 300 31336 308 31342
rect 289 31326 308 31336
rect 196 31269 204 31299
rect 216 31269 232 31299
rect 196 31265 232 31269
rect 196 31257 226 31265
rect 300 31257 308 31326
rect 332 31333 351 31367
rect 361 31339 381 31367
rect 361 31333 375 31339
rect 400 31333 411 31377
rect 442 31372 500 31379
rect 466 31371 500 31372
rect 565 31371 599 31379
rect 497 31355 500 31371
rect 596 31355 599 31371
rect 466 31354 500 31355
rect 442 31347 500 31354
rect 565 31347 599 31355
rect 612 31338 614 31388
rect 332 31309 342 31333
rect 336 31297 342 31309
rect 224 31241 226 31257
rect 332 31229 342 31297
rect 400 31301 404 31309
rect 400 31267 408 31301
rect 434 31267 438 31301
rect 454 31285 504 31287
rect 504 31269 506 31285
rect 514 31279 530 31285
rect 532 31279 548 31285
rect 525 31269 548 31278
rect 400 31259 404 31267
rect 498 31259 506 31269
rect 504 31235 506 31259
rect 514 31249 515 31269
rect 525 31244 528 31269
rect 547 31249 548 31269
rect 557 31259 564 31269
rect 514 31235 548 31239
rect 151 31188 156 31222
rect 174 31219 246 31227
rect 256 31219 328 31227
rect 336 31221 342 31229
rect 400 31224 404 31229
rect 180 31191 185 31219
rect 174 31183 246 31191
rect 256 31183 328 31191
rect 332 31189 336 31219
rect 400 31190 438 31224
rect 224 31153 226 31169
rect 196 31145 226 31153
rect 196 31141 232 31145
rect 196 31111 204 31141
rect 216 31111 232 31141
rect 224 31064 226 31111
rect 300 31084 308 31153
rect 332 31151 342 31189
rect 400 31181 404 31190
rect 454 31175 504 31177
rect 494 31171 548 31175
rect 494 31166 514 31171
rect 504 31151 506 31166
rect 336 31139 342 31151
rect 289 31074 308 31084
rect 300 31068 308 31074
rect 332 31105 342 31139
rect 400 31143 404 31151
rect 400 31109 408 31143
rect 434 31109 438 31143
rect 498 31141 506 31151
rect 514 31141 515 31161
rect 504 31125 506 31141
rect 525 31132 528 31166
rect 547 31141 548 31161
rect 557 31141 564 31151
rect 514 31125 530 31131
rect 532 31125 548 31131
rect 332 31077 373 31105
rect 332 31071 351 31077
rect 107 31017 119 31051
rect 129 31017 149 31051
rect 196 31030 204 31064
rect 216 31030 232 31064
rect 244 31058 257 31064
rect 278 31058 291 31068
rect 244 31034 291 31058
rect 300 31058 321 31068
rect 336 31061 351 31071
rect 300 31034 329 31058
rect 332 31043 351 31061
rect 361 31071 375 31077
rect 400 31071 411 31109
rect 562 31072 612 31074
rect 361 31043 381 31071
rect 400 31043 409 31071
rect 466 31063 497 31071
rect 565 31063 596 31071
rect 442 31056 500 31063
rect 466 31055 500 31056
rect 565 31055 599 31063
rect 244 31030 257 31034
rect 42 30951 46 30985
rect 72 30951 76 30985
rect 42 30904 76 30908
rect 42 30889 46 30904
rect 72 30889 76 30904
rect 38 30871 80 30889
rect 16 30865 102 30871
rect 144 30865 148 31017
rect 174 30993 181 31021
rect 224 30983 226 31030
rect 300 31021 308 31034
rect 278 31010 305 31021
rect 332 30993 342 31043
rect 400 31023 404 31043
rect 497 31039 500 31055
rect 596 31039 599 31055
rect 466 31038 500 31039
rect 442 31031 500 31038
rect 565 31031 599 31039
rect 612 31022 614 31072
rect 256 30983 328 30991
rect 336 30985 342 30993
rect 400 30985 404 30993
rect 196 30953 204 30983
rect 216 30953 232 30983
rect 196 30949 232 30953
rect 196 30941 226 30949
rect 224 30925 226 30941
rect 332 30913 336 30981
rect 400 30951 408 30985
rect 434 30951 438 30985
rect 454 30969 504 30971
rect 504 30953 506 30969
rect 514 30963 530 30969
rect 532 30963 548 30969
rect 525 30953 548 30962
rect 400 30943 404 30951
rect 498 30943 506 30953
rect 504 30919 506 30943
rect 514 30933 515 30953
rect 525 30928 528 30953
rect 547 30933 548 30953
rect 557 30943 564 30953
rect 514 30919 548 30923
rect 400 30913 442 30914
rect 174 30903 246 30911
rect 400 30906 404 30913
rect 295 30872 300 30906
rect 324 30872 329 30906
rect 367 30889 438 30906
rect 367 30872 442 30889
rect 400 30871 442 30872
rect 378 30865 464 30871
rect 38 30849 80 30865
rect 400 30849 442 30865
rect -25 30835 25 30837
rect 42 30835 76 30849
rect 404 30835 438 30849
rect 455 30835 505 30837
rect 557 30835 607 30837
rect 16 30827 102 30835
rect 378 30827 464 30835
rect 8 30793 17 30827
rect 18 30825 51 30827
rect 80 30825 100 30827
rect 18 30793 100 30825
rect 380 30825 404 30827
rect 429 30825 438 30827
rect 442 30825 462 30827
rect 16 30785 102 30793
rect 42 30769 76 30785
rect 16 30749 38 30755
rect 42 30746 76 30750
rect 80 30749 102 30755
rect 42 30716 46 30746
rect 72 30716 76 30746
rect 42 30635 46 30669
rect 72 30635 76 30669
rect -25 30598 25 30600
rect -8 30590 14 30597
rect -8 30589 17 30590
rect 25 30589 27 30598
rect -12 30582 38 30589
rect -12 30581 34 30582
rect -12 30577 8 30581
rect 0 30565 8 30577
rect 14 30565 34 30581
rect 0 30564 34 30565
rect 0 30557 38 30564
rect 14 30556 17 30557
rect 25 30548 27 30557
rect 42 30528 45 30618
rect 69 30603 80 30635
rect 107 30603 143 30631
rect 144 30603 148 30823
rect 332 30755 336 30823
rect 380 30793 462 30825
rect 463 30793 472 30827
rect 480 30793 497 30827
rect 378 30785 464 30793
rect 505 30785 507 30835
rect 514 30793 548 30827
rect 565 30793 582 30827
rect 607 30785 609 30835
rect 404 30769 438 30785
rect 400 30755 442 30756
rect 378 30749 404 30755
rect 442 30749 464 30755
rect 400 30748 404 30749
rect 174 30709 246 30717
rect 295 30714 300 30748
rect 324 30714 329 30748
rect 224 30679 226 30695
rect 196 30671 226 30679
rect 332 30677 336 30745
rect 367 30714 438 30748
rect 400 30707 404 30714
rect 454 30701 504 30703
rect 494 30697 548 30701
rect 494 30692 514 30697
rect 504 30677 506 30692
rect 196 30667 232 30671
rect 196 30637 204 30667
rect 216 30637 232 30667
rect 400 30669 404 30677
rect 107 30597 119 30603
rect 109 30569 119 30597
rect 129 30569 149 30603
rect 174 30599 181 30629
rect 224 30590 226 30637
rect 256 30629 328 30637
rect 332 30635 336 30665
rect 400 30635 408 30669
rect 434 30635 438 30669
rect 498 30667 506 30677
rect 514 30667 515 30687
rect 504 30651 506 30667
rect 525 30658 528 30692
rect 547 30667 548 30687
rect 557 30667 564 30677
rect 514 30651 530 30657
rect 532 30651 548 30657
rect 278 30599 305 30610
rect 42 30477 46 30511
rect 72 30477 76 30511
rect 38 30439 80 30440
rect 42 30398 76 30432
rect 79 30398 113 30432
rect 42 30319 46 30353
rect 72 30319 76 30353
rect -25 30282 25 30284
rect -8 30274 14 30281
rect -8 30273 17 30274
rect 25 30273 27 30282
rect -12 30266 38 30273
rect -12 30265 34 30266
rect -12 30261 8 30265
rect 0 30249 8 30261
rect 14 30249 34 30265
rect 0 30248 34 30249
rect 0 30241 38 30248
rect 14 30240 17 30241
rect 25 30232 27 30241
rect 42 30212 45 30302
rect 71 30271 80 30299
rect 69 30233 80 30271
rect 144 30261 148 30569
rect 196 30556 204 30590
rect 216 30556 232 30590
rect 244 30586 257 30590
rect 300 30586 308 30599
rect 332 30597 342 30635
rect 400 30627 404 30635
rect 336 30587 342 30597
rect 244 30562 291 30586
rect 244 30556 257 30562
rect 224 30509 226 30556
rect 278 30552 291 30562
rect 300 30562 329 30586
rect 332 30577 342 30587
rect 400 30587 409 30615
rect 562 30598 612 30600
rect 466 30589 497 30597
rect 565 30589 596 30597
rect 300 30552 321 30562
rect 300 30546 308 30552
rect 289 30536 308 30546
rect 196 30479 204 30509
rect 216 30479 232 30509
rect 196 30475 232 30479
rect 196 30467 226 30475
rect 300 30467 308 30536
rect 332 30543 351 30577
rect 361 30549 381 30577
rect 361 30543 375 30549
rect 400 30543 411 30587
rect 442 30582 500 30589
rect 466 30581 500 30582
rect 565 30581 599 30589
rect 497 30565 500 30581
rect 596 30565 599 30581
rect 466 30564 500 30565
rect 442 30557 500 30564
rect 565 30557 599 30565
rect 612 30548 614 30598
rect 332 30519 342 30543
rect 336 30507 342 30519
rect 224 30451 226 30467
rect 332 30439 342 30507
rect 400 30511 404 30519
rect 400 30477 408 30511
rect 434 30477 438 30511
rect 454 30495 504 30497
rect 504 30479 506 30495
rect 514 30489 530 30495
rect 532 30489 548 30495
rect 525 30479 548 30488
rect 400 30469 404 30477
rect 498 30469 506 30479
rect 504 30445 506 30469
rect 514 30459 515 30479
rect 525 30454 528 30479
rect 547 30459 548 30479
rect 557 30469 564 30479
rect 514 30445 548 30449
rect 151 30398 156 30432
rect 174 30429 246 30437
rect 256 30429 328 30437
rect 336 30431 342 30439
rect 400 30434 404 30439
rect 180 30401 185 30429
rect 174 30393 246 30401
rect 256 30393 328 30401
rect 332 30399 336 30429
rect 400 30400 438 30434
rect 224 30363 226 30379
rect 196 30355 226 30363
rect 196 30351 232 30355
rect 196 30321 204 30351
rect 216 30321 232 30351
rect 224 30274 226 30321
rect 300 30294 308 30363
rect 332 30361 342 30399
rect 400 30391 404 30400
rect 454 30385 504 30387
rect 494 30381 548 30385
rect 494 30376 514 30381
rect 504 30361 506 30376
rect 336 30349 342 30361
rect 289 30284 308 30294
rect 300 30278 308 30284
rect 332 30315 342 30349
rect 400 30353 404 30361
rect 400 30319 408 30353
rect 434 30319 438 30353
rect 498 30351 506 30361
rect 514 30351 515 30371
rect 504 30335 506 30351
rect 525 30342 528 30376
rect 547 30351 548 30371
rect 557 30351 564 30361
rect 514 30335 530 30341
rect 532 30335 548 30341
rect 332 30287 373 30315
rect 332 30281 351 30287
rect 107 30227 119 30261
rect 129 30227 149 30261
rect 196 30240 204 30274
rect 216 30240 232 30274
rect 244 30268 257 30274
rect 278 30268 291 30278
rect 244 30244 291 30268
rect 300 30268 321 30278
rect 336 30271 351 30281
rect 300 30244 329 30268
rect 332 30253 351 30271
rect 361 30281 375 30287
rect 400 30281 411 30319
rect 562 30282 612 30284
rect 361 30253 381 30281
rect 400 30253 409 30281
rect 466 30273 497 30281
rect 565 30273 596 30281
rect 442 30266 500 30273
rect 466 30265 500 30266
rect 565 30265 599 30273
rect 244 30240 257 30244
rect 42 30161 46 30195
rect 72 30161 76 30195
rect 42 30114 76 30118
rect 42 30099 46 30114
rect 72 30099 76 30114
rect 38 30081 80 30099
rect 16 30075 102 30081
rect 144 30075 148 30227
rect 174 30203 181 30231
rect 224 30193 226 30240
rect 300 30231 308 30244
rect 278 30220 305 30231
rect 332 30203 342 30253
rect 400 30233 404 30253
rect 497 30249 500 30265
rect 596 30249 599 30265
rect 466 30248 500 30249
rect 442 30241 500 30248
rect 565 30241 599 30249
rect 612 30232 614 30282
rect 256 30193 328 30201
rect 336 30195 342 30203
rect 400 30195 404 30203
rect 196 30163 204 30193
rect 216 30163 232 30193
rect 196 30159 232 30163
rect 196 30151 226 30159
rect 224 30135 226 30151
rect 332 30123 336 30191
rect 400 30161 408 30195
rect 434 30161 438 30195
rect 454 30179 504 30181
rect 504 30163 506 30179
rect 514 30173 530 30179
rect 532 30173 548 30179
rect 525 30163 548 30172
rect 400 30153 404 30161
rect 498 30153 506 30163
rect 504 30129 506 30153
rect 514 30143 515 30163
rect 525 30138 528 30163
rect 547 30143 548 30163
rect 557 30153 564 30163
rect 514 30129 548 30133
rect 400 30123 442 30124
rect 174 30113 246 30121
rect 400 30116 404 30123
rect 295 30082 300 30116
rect 324 30082 329 30116
rect 367 30099 438 30116
rect 367 30082 442 30099
rect 400 30081 442 30082
rect 378 30075 464 30081
rect 38 30059 80 30075
rect 400 30059 442 30075
rect -25 30045 25 30047
rect 42 30045 76 30059
rect 404 30045 438 30059
rect 455 30045 505 30047
rect 557 30045 607 30047
rect 16 30037 102 30045
rect 378 30037 464 30045
rect 8 30003 17 30037
rect 18 30035 51 30037
rect 80 30035 100 30037
rect 18 30003 100 30035
rect 380 30035 404 30037
rect 429 30035 438 30037
rect 442 30035 462 30037
rect 16 29995 102 30003
rect 42 29979 76 29995
rect 16 29959 38 29965
rect 42 29956 76 29960
rect 80 29959 102 29965
rect 42 29926 46 29956
rect 72 29926 76 29956
rect 42 29845 46 29879
rect 72 29845 76 29879
rect -25 29808 25 29810
rect -8 29800 14 29807
rect -8 29799 17 29800
rect 25 29799 27 29808
rect -12 29792 38 29799
rect -12 29791 34 29792
rect -12 29787 8 29791
rect 0 29775 8 29787
rect 14 29775 34 29791
rect 0 29774 34 29775
rect 0 29767 38 29774
rect 14 29766 17 29767
rect 25 29758 27 29767
rect 42 29738 45 29828
rect 69 29813 80 29845
rect 107 29813 143 29841
rect 144 29813 148 30033
rect 332 29965 336 30033
rect 380 30003 462 30035
rect 463 30003 472 30037
rect 480 30003 497 30037
rect 378 29995 464 30003
rect 505 29995 507 30045
rect 514 30003 548 30037
rect 565 30003 582 30037
rect 607 29995 609 30045
rect 404 29979 438 29995
rect 400 29965 442 29966
rect 378 29959 404 29965
rect 442 29959 464 29965
rect 400 29958 404 29959
rect 174 29919 246 29927
rect 295 29924 300 29958
rect 324 29924 329 29958
rect 224 29889 226 29905
rect 196 29881 226 29889
rect 332 29887 336 29955
rect 367 29924 438 29958
rect 400 29917 404 29924
rect 454 29911 504 29913
rect 494 29907 548 29911
rect 494 29902 514 29907
rect 504 29887 506 29902
rect 196 29877 232 29881
rect 196 29847 204 29877
rect 216 29847 232 29877
rect 400 29879 404 29887
rect 107 29807 119 29813
rect 109 29779 119 29807
rect 129 29779 149 29813
rect 174 29809 181 29839
rect 224 29800 226 29847
rect 256 29839 328 29847
rect 332 29845 336 29875
rect 400 29845 408 29879
rect 434 29845 438 29879
rect 498 29877 506 29887
rect 514 29877 515 29897
rect 504 29861 506 29877
rect 525 29868 528 29902
rect 547 29877 548 29897
rect 557 29877 564 29887
rect 514 29861 530 29867
rect 532 29861 548 29867
rect 278 29809 305 29820
rect 42 29687 46 29721
rect 72 29687 76 29721
rect 38 29649 80 29650
rect 42 29608 76 29642
rect 79 29608 113 29642
rect 42 29529 46 29563
rect 72 29529 76 29563
rect -25 29492 25 29494
rect -8 29484 14 29491
rect -8 29483 17 29484
rect 25 29483 27 29492
rect -12 29476 38 29483
rect -12 29475 34 29476
rect -12 29471 8 29475
rect 0 29459 8 29471
rect 14 29459 34 29475
rect 0 29458 34 29459
rect 0 29451 38 29458
rect 14 29450 17 29451
rect 25 29442 27 29451
rect 42 29422 45 29512
rect 71 29481 80 29509
rect 69 29443 80 29481
rect 144 29471 148 29779
rect 196 29766 204 29800
rect 216 29766 232 29800
rect 244 29796 257 29800
rect 300 29796 308 29809
rect 332 29807 342 29845
rect 400 29837 404 29845
rect 336 29797 342 29807
rect 244 29772 291 29796
rect 244 29766 257 29772
rect 224 29719 226 29766
rect 278 29762 291 29772
rect 300 29772 329 29796
rect 332 29787 342 29797
rect 400 29797 409 29825
rect 562 29808 612 29810
rect 466 29799 497 29807
rect 565 29799 596 29807
rect 300 29762 321 29772
rect 300 29756 308 29762
rect 289 29746 308 29756
rect 196 29689 204 29719
rect 216 29689 232 29719
rect 196 29685 232 29689
rect 196 29677 226 29685
rect 300 29677 308 29746
rect 332 29753 351 29787
rect 361 29759 381 29787
rect 361 29753 375 29759
rect 400 29753 411 29797
rect 442 29792 500 29799
rect 466 29791 500 29792
rect 565 29791 599 29799
rect 497 29775 500 29791
rect 596 29775 599 29791
rect 466 29774 500 29775
rect 442 29767 500 29774
rect 565 29767 599 29775
rect 612 29758 614 29808
rect 332 29729 342 29753
rect 336 29717 342 29729
rect 224 29661 226 29677
rect 332 29649 342 29717
rect 400 29721 404 29729
rect 400 29687 408 29721
rect 434 29687 438 29721
rect 454 29705 504 29707
rect 504 29689 506 29705
rect 514 29699 530 29705
rect 532 29699 548 29705
rect 525 29689 548 29698
rect 400 29679 404 29687
rect 498 29679 506 29689
rect 504 29655 506 29679
rect 514 29669 515 29689
rect 525 29664 528 29689
rect 547 29669 548 29689
rect 557 29679 564 29689
rect 514 29655 548 29659
rect 151 29608 156 29642
rect 174 29639 246 29647
rect 256 29639 328 29647
rect 336 29641 342 29649
rect 400 29644 404 29649
rect 180 29611 185 29639
rect 174 29603 246 29611
rect 256 29603 328 29611
rect 332 29609 336 29639
rect 400 29610 438 29644
rect 224 29573 226 29589
rect 196 29565 226 29573
rect 196 29561 232 29565
rect 196 29531 204 29561
rect 216 29531 232 29561
rect 224 29484 226 29531
rect 300 29504 308 29573
rect 332 29571 342 29609
rect 400 29601 404 29610
rect 454 29595 504 29597
rect 494 29591 548 29595
rect 494 29586 514 29591
rect 504 29571 506 29586
rect 336 29559 342 29571
rect 289 29494 308 29504
rect 300 29488 308 29494
rect 332 29525 342 29559
rect 400 29563 404 29571
rect 400 29529 408 29563
rect 434 29529 438 29563
rect 498 29561 506 29571
rect 514 29561 515 29581
rect 504 29545 506 29561
rect 525 29552 528 29586
rect 547 29561 548 29581
rect 557 29561 564 29571
rect 514 29545 530 29551
rect 532 29545 548 29551
rect 332 29497 373 29525
rect 332 29491 351 29497
rect 107 29437 119 29471
rect 129 29437 149 29471
rect 196 29450 204 29484
rect 216 29450 232 29484
rect 244 29478 257 29484
rect 278 29478 291 29488
rect 244 29454 291 29478
rect 300 29478 321 29488
rect 336 29481 351 29491
rect 300 29454 329 29478
rect 332 29463 351 29481
rect 361 29491 375 29497
rect 400 29491 411 29529
rect 562 29492 612 29494
rect 361 29463 381 29491
rect 400 29463 409 29491
rect 466 29483 497 29491
rect 565 29483 596 29491
rect 442 29476 500 29483
rect 466 29475 500 29476
rect 565 29475 599 29483
rect 244 29450 257 29454
rect 42 29371 46 29405
rect 72 29371 76 29405
rect 42 29324 76 29328
rect 42 29309 46 29324
rect 72 29309 76 29324
rect 38 29291 80 29309
rect 16 29285 102 29291
rect 144 29285 148 29437
rect 174 29413 181 29441
rect 224 29403 226 29450
rect 300 29441 308 29454
rect 278 29430 305 29441
rect 332 29413 342 29463
rect 400 29443 404 29463
rect 497 29459 500 29475
rect 596 29459 599 29475
rect 466 29458 500 29459
rect 442 29451 500 29458
rect 565 29451 599 29459
rect 612 29442 614 29492
rect 256 29403 328 29411
rect 336 29405 342 29413
rect 400 29405 404 29413
rect 196 29373 204 29403
rect 216 29373 232 29403
rect 196 29369 232 29373
rect 196 29361 226 29369
rect 224 29345 226 29361
rect 332 29333 336 29401
rect 400 29371 408 29405
rect 434 29371 438 29405
rect 454 29389 504 29391
rect 504 29373 506 29389
rect 514 29383 530 29389
rect 532 29383 548 29389
rect 525 29373 548 29382
rect 400 29363 404 29371
rect 498 29363 506 29373
rect 504 29339 506 29363
rect 514 29353 515 29373
rect 525 29348 528 29373
rect 547 29353 548 29373
rect 557 29363 564 29373
rect 514 29339 548 29343
rect 400 29333 442 29334
rect 174 29323 246 29331
rect 400 29326 404 29333
rect 295 29292 300 29326
rect 324 29292 329 29326
rect 367 29309 438 29326
rect 367 29292 442 29309
rect 400 29291 442 29292
rect 378 29285 464 29291
rect 38 29269 80 29285
rect 400 29269 442 29285
rect -25 29255 25 29257
rect 42 29255 76 29269
rect 404 29255 438 29269
rect 455 29255 505 29257
rect 557 29255 607 29257
rect 16 29247 102 29255
rect 378 29247 464 29255
rect 8 29213 17 29247
rect 18 29245 51 29247
rect 80 29245 100 29247
rect 18 29213 100 29245
rect 380 29245 404 29247
rect 429 29245 438 29247
rect 442 29245 462 29247
rect 16 29205 102 29213
rect 42 29189 76 29205
rect 16 29169 38 29175
rect 42 29166 76 29170
rect 80 29169 102 29175
rect 42 29136 46 29166
rect 72 29136 76 29166
rect 42 29055 46 29089
rect 72 29055 76 29089
rect -25 29018 25 29020
rect -8 29010 14 29017
rect -8 29009 17 29010
rect 25 29009 27 29018
rect -12 29002 38 29009
rect -12 29001 34 29002
rect -12 28997 8 29001
rect 0 28985 8 28997
rect 14 28985 34 29001
rect 0 28984 34 28985
rect 0 28977 38 28984
rect 14 28976 17 28977
rect 25 28968 27 28977
rect 42 28948 45 29038
rect 69 29023 80 29055
rect 107 29023 143 29051
rect 144 29023 148 29243
rect 332 29175 336 29243
rect 380 29213 462 29245
rect 463 29213 472 29247
rect 480 29213 497 29247
rect 378 29205 464 29213
rect 505 29205 507 29255
rect 514 29213 548 29247
rect 565 29213 582 29247
rect 607 29205 609 29255
rect 404 29189 438 29205
rect 400 29175 442 29176
rect 378 29169 404 29175
rect 442 29169 464 29175
rect 400 29168 404 29169
rect 174 29129 246 29137
rect 295 29134 300 29168
rect 324 29134 329 29168
rect 224 29099 226 29115
rect 196 29091 226 29099
rect 332 29097 336 29165
rect 367 29134 438 29168
rect 400 29127 404 29134
rect 454 29121 504 29123
rect 494 29117 548 29121
rect 494 29112 514 29117
rect 504 29097 506 29112
rect 196 29087 232 29091
rect 196 29057 204 29087
rect 216 29057 232 29087
rect 400 29089 404 29097
rect 107 29017 119 29023
rect 109 28989 119 29017
rect 129 28989 149 29023
rect 174 29019 181 29049
rect 224 29010 226 29057
rect 256 29049 328 29057
rect 332 29055 336 29085
rect 400 29055 408 29089
rect 434 29055 438 29089
rect 498 29087 506 29097
rect 514 29087 515 29107
rect 504 29071 506 29087
rect 525 29078 528 29112
rect 547 29087 548 29107
rect 557 29087 564 29097
rect 514 29071 530 29077
rect 532 29071 548 29077
rect 278 29019 305 29030
rect 42 28897 46 28931
rect 72 28897 76 28931
rect 38 28859 80 28860
rect 42 28818 76 28852
rect 79 28818 113 28852
rect 42 28739 46 28773
rect 72 28739 76 28773
rect -25 28702 25 28704
rect -8 28694 14 28701
rect -8 28693 17 28694
rect 25 28693 27 28702
rect -12 28686 38 28693
rect -12 28685 34 28686
rect -12 28681 8 28685
rect 0 28669 8 28681
rect 14 28669 34 28685
rect 0 28668 34 28669
rect 0 28661 38 28668
rect 14 28660 17 28661
rect 25 28652 27 28661
rect 42 28632 45 28722
rect 71 28691 80 28719
rect 69 28653 80 28691
rect 144 28681 148 28989
rect 196 28976 204 29010
rect 216 28976 232 29010
rect 244 29006 257 29010
rect 300 29006 308 29019
rect 332 29017 342 29055
rect 400 29047 404 29055
rect 336 29007 342 29017
rect 244 28982 291 29006
rect 244 28976 257 28982
rect 224 28929 226 28976
rect 278 28972 291 28982
rect 300 28982 329 29006
rect 332 28997 342 29007
rect 400 29007 409 29035
rect 562 29018 612 29020
rect 466 29009 497 29017
rect 565 29009 596 29017
rect 300 28972 321 28982
rect 300 28966 308 28972
rect 289 28956 308 28966
rect 196 28899 204 28929
rect 216 28899 232 28929
rect 196 28895 232 28899
rect 196 28887 226 28895
rect 300 28887 308 28956
rect 332 28963 351 28997
rect 361 28969 381 28997
rect 361 28963 375 28969
rect 400 28963 411 29007
rect 442 29002 500 29009
rect 466 29001 500 29002
rect 565 29001 599 29009
rect 497 28985 500 29001
rect 596 28985 599 29001
rect 466 28984 500 28985
rect 442 28977 500 28984
rect 565 28977 599 28985
rect 612 28968 614 29018
rect 332 28939 342 28963
rect 336 28927 342 28939
rect 224 28871 226 28887
rect 332 28859 342 28927
rect 400 28931 404 28939
rect 400 28897 408 28931
rect 434 28897 438 28931
rect 454 28915 504 28917
rect 504 28899 506 28915
rect 514 28909 530 28915
rect 532 28909 548 28915
rect 525 28899 548 28908
rect 400 28889 404 28897
rect 498 28889 506 28899
rect 504 28865 506 28889
rect 514 28879 515 28899
rect 525 28874 528 28899
rect 547 28879 548 28899
rect 557 28889 564 28899
rect 514 28865 548 28869
rect 151 28818 156 28852
rect 174 28849 246 28857
rect 256 28849 328 28857
rect 336 28851 342 28859
rect 400 28854 404 28859
rect 180 28821 185 28849
rect 174 28813 246 28821
rect 256 28813 328 28821
rect 332 28819 336 28849
rect 400 28820 438 28854
rect 224 28783 226 28799
rect 196 28775 226 28783
rect 196 28771 232 28775
rect 196 28741 204 28771
rect 216 28741 232 28771
rect 224 28694 226 28741
rect 300 28714 308 28783
rect 332 28781 342 28819
rect 400 28811 404 28820
rect 454 28805 504 28807
rect 494 28801 548 28805
rect 494 28796 514 28801
rect 504 28781 506 28796
rect 336 28769 342 28781
rect 289 28704 308 28714
rect 300 28698 308 28704
rect 332 28735 342 28769
rect 400 28773 404 28781
rect 400 28739 408 28773
rect 434 28739 438 28773
rect 498 28771 506 28781
rect 514 28771 515 28791
rect 504 28755 506 28771
rect 525 28762 528 28796
rect 547 28771 548 28791
rect 557 28771 564 28781
rect 514 28755 530 28761
rect 532 28755 548 28761
rect 332 28707 373 28735
rect 332 28701 351 28707
rect 107 28647 119 28681
rect 129 28647 149 28681
rect 196 28660 204 28694
rect 216 28660 232 28694
rect 244 28688 257 28694
rect 278 28688 291 28698
rect 244 28664 291 28688
rect 300 28688 321 28698
rect 336 28691 351 28701
rect 300 28664 329 28688
rect 332 28673 351 28691
rect 361 28701 375 28707
rect 400 28701 411 28739
rect 562 28702 612 28704
rect 361 28673 381 28701
rect 400 28673 409 28701
rect 466 28693 497 28701
rect 565 28693 596 28701
rect 442 28686 500 28693
rect 466 28685 500 28686
rect 565 28685 599 28693
rect 244 28660 257 28664
rect 42 28581 46 28615
rect 72 28581 76 28615
rect 42 28534 76 28538
rect 42 28519 46 28534
rect 72 28519 76 28534
rect 38 28501 80 28519
rect 16 28495 102 28501
rect 144 28495 148 28647
rect 174 28623 181 28651
rect 224 28613 226 28660
rect 300 28651 308 28664
rect 278 28640 305 28651
rect 332 28623 342 28673
rect 400 28653 404 28673
rect 497 28669 500 28685
rect 596 28669 599 28685
rect 466 28668 500 28669
rect 442 28661 500 28668
rect 565 28661 599 28669
rect 612 28652 614 28702
rect 256 28613 328 28621
rect 336 28615 342 28623
rect 400 28615 404 28623
rect 196 28583 204 28613
rect 216 28583 232 28613
rect 196 28579 232 28583
rect 196 28571 226 28579
rect 224 28555 226 28571
rect 332 28543 336 28611
rect 400 28581 408 28615
rect 434 28581 438 28615
rect 454 28599 504 28601
rect 504 28583 506 28599
rect 514 28593 530 28599
rect 532 28593 548 28599
rect 525 28583 548 28592
rect 400 28573 404 28581
rect 498 28573 506 28583
rect 504 28549 506 28573
rect 514 28563 515 28583
rect 525 28558 528 28583
rect 547 28563 548 28583
rect 557 28573 564 28583
rect 514 28549 548 28553
rect 400 28543 442 28544
rect 174 28533 246 28541
rect 400 28536 404 28543
rect 295 28502 300 28536
rect 324 28502 329 28536
rect 367 28519 438 28536
rect 367 28502 442 28519
rect 400 28501 442 28502
rect 378 28495 464 28501
rect 38 28479 80 28495
rect 400 28479 442 28495
rect -25 28465 25 28467
rect 42 28465 76 28479
rect 404 28465 438 28479
rect 455 28465 505 28467
rect 557 28465 607 28467
rect 16 28457 102 28465
rect 378 28457 464 28465
rect 8 28423 17 28457
rect 18 28455 51 28457
rect 80 28455 100 28457
rect 18 28423 100 28455
rect 380 28455 404 28457
rect 429 28455 438 28457
rect 442 28455 462 28457
rect 16 28415 102 28423
rect 42 28399 76 28415
rect 16 28379 38 28385
rect 42 28376 76 28380
rect 80 28379 102 28385
rect 42 28346 46 28376
rect 72 28346 76 28376
rect 42 28265 46 28299
rect 72 28265 76 28299
rect -25 28228 25 28230
rect -8 28220 14 28227
rect -8 28219 17 28220
rect 25 28219 27 28228
rect -12 28212 38 28219
rect -12 28211 34 28212
rect -12 28207 8 28211
rect 0 28195 8 28207
rect 14 28195 34 28211
rect 0 28194 34 28195
rect 0 28187 38 28194
rect 14 28186 17 28187
rect 25 28178 27 28187
rect 42 28158 45 28248
rect 69 28233 80 28265
rect 107 28233 143 28261
rect 144 28233 148 28453
rect 332 28385 336 28453
rect 380 28423 462 28455
rect 463 28423 472 28457
rect 480 28423 497 28457
rect 378 28415 464 28423
rect 505 28415 507 28465
rect 514 28423 548 28457
rect 565 28423 582 28457
rect 607 28415 609 28465
rect 404 28399 438 28415
rect 400 28385 442 28386
rect 378 28379 404 28385
rect 442 28379 464 28385
rect 400 28378 404 28379
rect 174 28339 246 28347
rect 295 28344 300 28378
rect 324 28344 329 28378
rect 224 28309 226 28325
rect 196 28301 226 28309
rect 332 28307 336 28375
rect 367 28344 438 28378
rect 400 28337 404 28344
rect 454 28331 504 28333
rect 494 28327 548 28331
rect 494 28322 514 28327
rect 504 28307 506 28322
rect 196 28297 232 28301
rect 196 28267 204 28297
rect 216 28267 232 28297
rect 400 28299 404 28307
rect 107 28227 119 28233
rect 109 28199 119 28227
rect 129 28199 149 28233
rect 174 28229 181 28259
rect 224 28220 226 28267
rect 256 28259 328 28267
rect 332 28265 336 28295
rect 400 28265 408 28299
rect 434 28265 438 28299
rect 498 28297 506 28307
rect 514 28297 515 28317
rect 504 28281 506 28297
rect 525 28288 528 28322
rect 547 28297 548 28317
rect 557 28297 564 28307
rect 514 28281 530 28287
rect 532 28281 548 28287
rect 278 28229 305 28240
rect 42 28107 46 28141
rect 72 28107 76 28141
rect 38 28069 80 28070
rect 42 28028 76 28062
rect 79 28028 113 28062
rect 42 27949 46 27983
rect 72 27949 76 27983
rect -25 27912 25 27914
rect -8 27904 14 27911
rect -8 27903 17 27904
rect 25 27903 27 27912
rect -12 27896 38 27903
rect -12 27895 34 27896
rect -12 27891 8 27895
rect 0 27879 8 27891
rect 14 27879 34 27895
rect 0 27878 34 27879
rect 0 27871 38 27878
rect 14 27870 17 27871
rect 25 27862 27 27871
rect 42 27842 45 27932
rect 71 27901 80 27929
rect 69 27863 80 27901
rect 144 27891 148 28199
rect 196 28186 204 28220
rect 216 28186 232 28220
rect 244 28216 257 28220
rect 300 28216 308 28229
rect 332 28227 342 28265
rect 400 28257 404 28265
rect 336 28217 342 28227
rect 244 28192 291 28216
rect 244 28186 257 28192
rect 224 28139 226 28186
rect 278 28182 291 28192
rect 300 28192 329 28216
rect 332 28207 342 28217
rect 400 28217 409 28245
rect 562 28228 612 28230
rect 466 28219 497 28227
rect 565 28219 596 28227
rect 300 28182 321 28192
rect 300 28176 308 28182
rect 289 28166 308 28176
rect 196 28109 204 28139
rect 216 28109 232 28139
rect 196 28105 232 28109
rect 196 28097 226 28105
rect 300 28097 308 28166
rect 332 28173 351 28207
rect 361 28179 381 28207
rect 361 28173 375 28179
rect 400 28173 411 28217
rect 442 28212 500 28219
rect 466 28211 500 28212
rect 565 28211 599 28219
rect 497 28195 500 28211
rect 596 28195 599 28211
rect 466 28194 500 28195
rect 442 28187 500 28194
rect 565 28187 599 28195
rect 612 28178 614 28228
rect 332 28149 342 28173
rect 336 28137 342 28149
rect 224 28081 226 28097
rect 332 28069 342 28137
rect 400 28141 404 28149
rect 400 28107 408 28141
rect 434 28107 438 28141
rect 454 28125 504 28127
rect 504 28109 506 28125
rect 514 28119 530 28125
rect 532 28119 548 28125
rect 525 28109 548 28118
rect 400 28099 404 28107
rect 498 28099 506 28109
rect 504 28075 506 28099
rect 514 28089 515 28109
rect 525 28084 528 28109
rect 547 28089 548 28109
rect 557 28099 564 28109
rect 514 28075 548 28079
rect 151 28028 156 28062
rect 174 28059 246 28067
rect 256 28059 328 28067
rect 336 28061 342 28069
rect 400 28064 404 28069
rect 180 28031 185 28059
rect 174 28023 246 28031
rect 256 28023 328 28031
rect 332 28029 336 28059
rect 400 28030 438 28064
rect 224 27993 226 28009
rect 196 27985 226 27993
rect 196 27981 232 27985
rect 196 27951 204 27981
rect 216 27951 232 27981
rect 224 27904 226 27951
rect 300 27924 308 27993
rect 332 27991 342 28029
rect 400 28021 404 28030
rect 454 28015 504 28017
rect 494 28011 548 28015
rect 494 28006 514 28011
rect 504 27991 506 28006
rect 336 27979 342 27991
rect 289 27914 308 27924
rect 300 27908 308 27914
rect 332 27945 342 27979
rect 400 27983 404 27991
rect 400 27949 408 27983
rect 434 27949 438 27983
rect 498 27981 506 27991
rect 514 27981 515 28001
rect 504 27965 506 27981
rect 525 27972 528 28006
rect 547 27981 548 28001
rect 557 27981 564 27991
rect 514 27965 530 27971
rect 532 27965 548 27971
rect 332 27917 373 27945
rect 332 27911 351 27917
rect 107 27857 119 27891
rect 129 27857 149 27891
rect 196 27870 204 27904
rect 216 27870 232 27904
rect 244 27898 257 27904
rect 278 27898 291 27908
rect 244 27874 291 27898
rect 300 27898 321 27908
rect 336 27901 351 27911
rect 300 27874 329 27898
rect 332 27883 351 27901
rect 361 27911 375 27917
rect 400 27911 411 27949
rect 562 27912 612 27914
rect 361 27883 381 27911
rect 400 27883 409 27911
rect 466 27903 497 27911
rect 565 27903 596 27911
rect 442 27896 500 27903
rect 466 27895 500 27896
rect 565 27895 599 27903
rect 244 27870 257 27874
rect 42 27791 46 27825
rect 72 27791 76 27825
rect 42 27744 76 27748
rect 42 27729 46 27744
rect 72 27729 76 27744
rect 38 27711 80 27729
rect 16 27705 102 27711
rect 144 27705 148 27857
rect 174 27833 181 27861
rect 224 27823 226 27870
rect 300 27861 308 27874
rect 278 27850 305 27861
rect 332 27833 342 27883
rect 400 27863 404 27883
rect 497 27879 500 27895
rect 596 27879 599 27895
rect 466 27878 500 27879
rect 442 27871 500 27878
rect 565 27871 599 27879
rect 612 27862 614 27912
rect 256 27823 328 27831
rect 336 27825 342 27833
rect 400 27825 404 27833
rect 196 27793 204 27823
rect 216 27793 232 27823
rect 196 27789 232 27793
rect 196 27781 226 27789
rect 224 27765 226 27781
rect 332 27753 336 27821
rect 400 27791 408 27825
rect 434 27791 438 27825
rect 454 27809 504 27811
rect 504 27793 506 27809
rect 514 27803 530 27809
rect 532 27803 548 27809
rect 525 27793 548 27802
rect 400 27783 404 27791
rect 498 27783 506 27793
rect 504 27759 506 27783
rect 514 27773 515 27793
rect 525 27768 528 27793
rect 547 27773 548 27793
rect 557 27783 564 27793
rect 514 27759 548 27763
rect 400 27753 442 27754
rect 174 27743 246 27751
rect 400 27746 404 27753
rect 295 27712 300 27746
rect 324 27712 329 27746
rect 367 27729 438 27746
rect 367 27712 442 27729
rect 400 27711 442 27712
rect 378 27705 464 27711
rect 38 27689 80 27705
rect 400 27689 442 27705
rect -25 27675 25 27677
rect 42 27675 76 27689
rect 404 27675 438 27689
rect 455 27675 505 27677
rect 557 27675 607 27677
rect 16 27667 102 27675
rect 378 27667 464 27675
rect 8 27633 17 27667
rect 18 27665 51 27667
rect 80 27665 100 27667
rect 18 27633 100 27665
rect 380 27665 404 27667
rect 429 27665 438 27667
rect 442 27665 462 27667
rect 16 27625 102 27633
rect 42 27609 76 27625
rect 16 27589 38 27595
rect 42 27586 76 27590
rect 80 27589 102 27595
rect 42 27556 46 27586
rect 72 27556 76 27586
rect 42 27475 46 27509
rect 72 27475 76 27509
rect -25 27438 25 27440
rect -8 27430 14 27437
rect -8 27429 17 27430
rect 25 27429 27 27438
rect -12 27422 38 27429
rect -12 27421 34 27422
rect -12 27417 8 27421
rect 0 27405 8 27417
rect 14 27405 34 27421
rect 0 27404 34 27405
rect 0 27397 38 27404
rect 14 27396 17 27397
rect 25 27388 27 27397
rect 42 27368 45 27458
rect 69 27443 80 27475
rect 107 27443 143 27471
rect 144 27443 148 27663
rect 332 27595 336 27663
rect 380 27633 462 27665
rect 463 27633 472 27667
rect 480 27633 497 27667
rect 378 27625 464 27633
rect 505 27625 507 27675
rect 514 27633 548 27667
rect 565 27633 582 27667
rect 607 27625 609 27675
rect 404 27609 438 27625
rect 400 27595 442 27596
rect 378 27589 404 27595
rect 442 27589 464 27595
rect 400 27588 404 27589
rect 174 27549 246 27557
rect 295 27554 300 27588
rect 324 27554 329 27588
rect 224 27519 226 27535
rect 196 27511 226 27519
rect 332 27517 336 27585
rect 367 27554 438 27588
rect 400 27547 404 27554
rect 454 27541 504 27543
rect 494 27537 548 27541
rect 494 27532 514 27537
rect 504 27517 506 27532
rect 196 27507 232 27511
rect 196 27477 204 27507
rect 216 27477 232 27507
rect 400 27509 404 27517
rect 107 27437 119 27443
rect 109 27409 119 27437
rect 129 27409 149 27443
rect 174 27439 181 27469
rect 224 27430 226 27477
rect 256 27469 328 27477
rect 332 27475 336 27505
rect 400 27475 408 27509
rect 434 27475 438 27509
rect 498 27507 506 27517
rect 514 27507 515 27527
rect 504 27491 506 27507
rect 525 27498 528 27532
rect 547 27507 548 27527
rect 557 27507 564 27517
rect 514 27491 530 27497
rect 532 27491 548 27497
rect 278 27439 305 27450
rect 42 27317 46 27351
rect 72 27317 76 27351
rect 38 27279 80 27280
rect 42 27238 76 27272
rect 79 27238 113 27272
rect 42 27159 46 27193
rect 72 27159 76 27193
rect -25 27122 25 27124
rect -8 27114 14 27121
rect -8 27113 17 27114
rect 25 27113 27 27122
rect -12 27106 38 27113
rect -12 27105 34 27106
rect -12 27101 8 27105
rect 0 27089 8 27101
rect 14 27089 34 27105
rect 0 27088 34 27089
rect 0 27081 38 27088
rect 14 27080 17 27081
rect 25 27072 27 27081
rect 42 27052 45 27142
rect 71 27111 80 27139
rect 69 27073 80 27111
rect 144 27101 148 27409
rect 196 27396 204 27430
rect 216 27396 232 27430
rect 244 27426 257 27430
rect 300 27426 308 27439
rect 332 27437 342 27475
rect 400 27467 404 27475
rect 336 27427 342 27437
rect 244 27402 291 27426
rect 244 27396 257 27402
rect 224 27349 226 27396
rect 278 27392 291 27402
rect 300 27402 329 27426
rect 332 27417 342 27427
rect 400 27427 409 27455
rect 562 27438 612 27440
rect 466 27429 497 27437
rect 565 27429 596 27437
rect 300 27392 321 27402
rect 300 27386 308 27392
rect 289 27376 308 27386
rect 196 27319 204 27349
rect 216 27319 232 27349
rect 196 27315 232 27319
rect 196 27307 226 27315
rect 300 27307 308 27376
rect 332 27383 351 27417
rect 361 27389 381 27417
rect 361 27383 375 27389
rect 400 27383 411 27427
rect 442 27422 500 27429
rect 466 27421 500 27422
rect 565 27421 599 27429
rect 497 27405 500 27421
rect 596 27405 599 27421
rect 466 27404 500 27405
rect 442 27397 500 27404
rect 565 27397 599 27405
rect 612 27388 614 27438
rect 332 27359 342 27383
rect 336 27347 342 27359
rect 224 27291 226 27307
rect 332 27279 342 27347
rect 400 27351 404 27359
rect 400 27317 408 27351
rect 434 27317 438 27351
rect 454 27335 504 27337
rect 504 27319 506 27335
rect 514 27329 530 27335
rect 532 27329 548 27335
rect 525 27319 548 27328
rect 400 27309 404 27317
rect 498 27309 506 27319
rect 504 27285 506 27309
rect 514 27299 515 27319
rect 525 27294 528 27319
rect 547 27299 548 27319
rect 557 27309 564 27319
rect 514 27285 548 27289
rect 151 27238 156 27272
rect 174 27269 246 27277
rect 256 27269 328 27277
rect 336 27271 342 27279
rect 400 27274 404 27279
rect 180 27241 185 27269
rect 174 27233 246 27241
rect 256 27233 328 27241
rect 332 27239 336 27269
rect 400 27240 438 27274
rect 224 27203 226 27219
rect 196 27195 226 27203
rect 196 27191 232 27195
rect 196 27161 204 27191
rect 216 27161 232 27191
rect 224 27114 226 27161
rect 300 27134 308 27203
rect 332 27201 342 27239
rect 400 27231 404 27240
rect 454 27225 504 27227
rect 494 27221 548 27225
rect 494 27216 514 27221
rect 504 27201 506 27216
rect 336 27189 342 27201
rect 289 27124 308 27134
rect 300 27118 308 27124
rect 332 27155 342 27189
rect 400 27193 404 27201
rect 400 27159 408 27193
rect 434 27159 438 27193
rect 498 27191 506 27201
rect 514 27191 515 27211
rect 504 27175 506 27191
rect 525 27182 528 27216
rect 547 27191 548 27211
rect 557 27191 564 27201
rect 514 27175 530 27181
rect 532 27175 548 27181
rect 332 27127 373 27155
rect 332 27121 351 27127
rect 107 27067 119 27101
rect 129 27067 149 27101
rect 196 27080 204 27114
rect 216 27080 232 27114
rect 244 27108 257 27114
rect 278 27108 291 27118
rect 244 27084 291 27108
rect 300 27108 321 27118
rect 336 27111 351 27121
rect 300 27084 329 27108
rect 332 27093 351 27111
rect 361 27121 375 27127
rect 400 27121 411 27159
rect 562 27122 612 27124
rect 361 27093 381 27121
rect 400 27093 409 27121
rect 466 27113 497 27121
rect 565 27113 596 27121
rect 442 27106 500 27113
rect 466 27105 500 27106
rect 565 27105 599 27113
rect 244 27080 257 27084
rect 42 27001 46 27035
rect 72 27001 76 27035
rect 42 26954 76 26958
rect 42 26939 46 26954
rect 72 26939 76 26954
rect 38 26921 80 26939
rect 16 26915 102 26921
rect 144 26915 148 27067
rect 174 27043 181 27071
rect 224 27033 226 27080
rect 300 27071 308 27084
rect 278 27060 305 27071
rect 332 27043 342 27093
rect 400 27073 404 27093
rect 497 27089 500 27105
rect 596 27089 599 27105
rect 466 27088 500 27089
rect 442 27081 500 27088
rect 565 27081 599 27089
rect 612 27072 614 27122
rect 256 27033 328 27041
rect 336 27035 342 27043
rect 400 27035 404 27043
rect 196 27003 204 27033
rect 216 27003 232 27033
rect 196 26999 232 27003
rect 196 26991 226 26999
rect 224 26975 226 26991
rect 332 26963 336 27031
rect 400 27001 408 27035
rect 434 27001 438 27035
rect 454 27019 504 27021
rect 504 27003 506 27019
rect 514 27013 530 27019
rect 532 27013 548 27019
rect 525 27003 548 27012
rect 400 26993 404 27001
rect 498 26993 506 27003
rect 504 26969 506 26993
rect 514 26983 515 27003
rect 525 26978 528 27003
rect 547 26983 548 27003
rect 557 26993 564 27003
rect 514 26969 548 26973
rect 400 26963 442 26964
rect 174 26953 246 26961
rect 400 26956 404 26963
rect 295 26922 300 26956
rect 324 26922 329 26956
rect 367 26939 438 26956
rect 367 26922 442 26939
rect 400 26921 442 26922
rect 378 26915 464 26921
rect 38 26899 80 26915
rect 400 26899 442 26915
rect -25 26885 25 26887
rect 42 26885 76 26899
rect 404 26885 438 26899
rect 455 26885 505 26887
rect 557 26885 607 26887
rect 16 26877 102 26885
rect 378 26877 464 26885
rect 8 26843 17 26877
rect 18 26875 51 26877
rect 80 26875 100 26877
rect 18 26843 100 26875
rect 380 26875 404 26877
rect 429 26875 438 26877
rect 442 26875 462 26877
rect 16 26835 102 26843
rect 42 26819 76 26835
rect 16 26799 38 26805
rect 42 26796 76 26800
rect 80 26799 102 26805
rect 42 26766 46 26796
rect 72 26766 76 26796
rect 42 26685 46 26719
rect 72 26685 76 26719
rect -25 26648 25 26650
rect -8 26640 14 26647
rect -8 26639 17 26640
rect 25 26639 27 26648
rect -12 26632 38 26639
rect -12 26631 34 26632
rect -12 26627 8 26631
rect 0 26615 8 26627
rect 14 26615 34 26631
rect 0 26614 34 26615
rect 0 26607 38 26614
rect 14 26606 17 26607
rect 25 26598 27 26607
rect 42 26578 45 26668
rect 69 26653 80 26685
rect 107 26653 143 26681
rect 144 26653 148 26873
rect 332 26805 336 26873
rect 380 26843 462 26875
rect 463 26843 472 26877
rect 480 26843 497 26877
rect 378 26835 464 26843
rect 505 26835 507 26885
rect 514 26843 548 26877
rect 565 26843 582 26877
rect 607 26835 609 26885
rect 404 26819 438 26835
rect 400 26805 442 26806
rect 378 26799 404 26805
rect 442 26799 464 26805
rect 400 26798 404 26799
rect 174 26759 246 26767
rect 295 26764 300 26798
rect 324 26764 329 26798
rect 224 26729 226 26745
rect 196 26721 226 26729
rect 332 26727 336 26795
rect 367 26764 438 26798
rect 400 26757 404 26764
rect 454 26751 504 26753
rect 494 26747 548 26751
rect 494 26742 514 26747
rect 504 26727 506 26742
rect 196 26717 232 26721
rect 196 26687 204 26717
rect 216 26687 232 26717
rect 400 26719 404 26727
rect 107 26647 119 26653
rect 109 26619 119 26647
rect 129 26619 149 26653
rect 174 26649 181 26679
rect 224 26640 226 26687
rect 256 26679 328 26687
rect 332 26685 336 26715
rect 400 26685 408 26719
rect 434 26685 438 26719
rect 498 26717 506 26727
rect 514 26717 515 26737
rect 504 26701 506 26717
rect 525 26708 528 26742
rect 547 26717 548 26737
rect 557 26717 564 26727
rect 514 26701 530 26707
rect 532 26701 548 26707
rect 278 26649 305 26660
rect 42 26527 46 26561
rect 72 26527 76 26561
rect 38 26489 80 26490
rect 42 26448 76 26482
rect 79 26448 113 26482
rect 42 26369 46 26403
rect 72 26369 76 26403
rect -25 26332 25 26334
rect -8 26324 14 26331
rect -8 26323 17 26324
rect 25 26323 27 26332
rect -12 26316 38 26323
rect -12 26315 34 26316
rect -12 26311 8 26315
rect 0 26299 8 26311
rect 14 26299 34 26315
rect 0 26298 34 26299
rect 0 26291 38 26298
rect 14 26290 17 26291
rect 25 26282 27 26291
rect 42 26262 45 26352
rect 71 26321 80 26349
rect 69 26283 80 26321
rect 144 26311 148 26619
rect 196 26606 204 26640
rect 216 26606 232 26640
rect 244 26636 257 26640
rect 300 26636 308 26649
rect 332 26647 342 26685
rect 400 26677 404 26685
rect 336 26637 342 26647
rect 244 26612 291 26636
rect 244 26606 257 26612
rect 224 26559 226 26606
rect 278 26602 291 26612
rect 300 26612 329 26636
rect 332 26627 342 26637
rect 400 26637 409 26665
rect 562 26648 612 26650
rect 466 26639 497 26647
rect 565 26639 596 26647
rect 300 26602 321 26612
rect 300 26596 308 26602
rect 289 26586 308 26596
rect 196 26529 204 26559
rect 216 26529 232 26559
rect 196 26525 232 26529
rect 196 26517 226 26525
rect 300 26517 308 26586
rect 332 26593 351 26627
rect 361 26599 381 26627
rect 361 26593 375 26599
rect 400 26593 411 26637
rect 442 26632 500 26639
rect 466 26631 500 26632
rect 565 26631 599 26639
rect 497 26615 500 26631
rect 596 26615 599 26631
rect 466 26614 500 26615
rect 442 26607 500 26614
rect 565 26607 599 26615
rect 612 26598 614 26648
rect 332 26569 342 26593
rect 336 26557 342 26569
rect 224 26501 226 26517
rect 332 26489 342 26557
rect 400 26561 404 26569
rect 400 26527 408 26561
rect 434 26527 438 26561
rect 454 26545 504 26547
rect 504 26529 506 26545
rect 514 26539 530 26545
rect 532 26539 548 26545
rect 525 26529 548 26538
rect 400 26519 404 26527
rect 498 26519 506 26529
rect 504 26495 506 26519
rect 514 26509 515 26529
rect 525 26504 528 26529
rect 547 26509 548 26529
rect 557 26519 564 26529
rect 514 26495 548 26499
rect 151 26448 156 26482
rect 174 26479 246 26487
rect 256 26479 328 26487
rect 336 26481 342 26489
rect 400 26484 404 26489
rect 180 26451 185 26479
rect 174 26443 246 26451
rect 256 26443 328 26451
rect 332 26449 336 26479
rect 400 26450 438 26484
rect 224 26413 226 26429
rect 196 26405 226 26413
rect 196 26401 232 26405
rect 196 26371 204 26401
rect 216 26371 232 26401
rect 224 26324 226 26371
rect 300 26344 308 26413
rect 332 26411 342 26449
rect 400 26441 404 26450
rect 454 26435 504 26437
rect 494 26431 548 26435
rect 494 26426 514 26431
rect 504 26411 506 26426
rect 336 26399 342 26411
rect 289 26334 308 26344
rect 300 26328 308 26334
rect 332 26365 342 26399
rect 400 26403 404 26411
rect 400 26369 408 26403
rect 434 26369 438 26403
rect 498 26401 506 26411
rect 514 26401 515 26421
rect 504 26385 506 26401
rect 525 26392 528 26426
rect 547 26401 548 26421
rect 557 26401 564 26411
rect 514 26385 530 26391
rect 532 26385 548 26391
rect 332 26337 373 26365
rect 332 26331 351 26337
rect 107 26277 119 26311
rect 129 26277 149 26311
rect 196 26290 204 26324
rect 216 26290 232 26324
rect 244 26318 257 26324
rect 278 26318 291 26328
rect 244 26294 291 26318
rect 300 26318 321 26328
rect 336 26321 351 26331
rect 300 26294 329 26318
rect 332 26303 351 26321
rect 361 26331 375 26337
rect 400 26331 411 26369
rect 562 26332 612 26334
rect 361 26303 381 26331
rect 400 26303 409 26331
rect 466 26323 497 26331
rect 565 26323 596 26331
rect 442 26316 500 26323
rect 466 26315 500 26316
rect 565 26315 599 26323
rect 244 26290 257 26294
rect 42 26211 46 26245
rect 72 26211 76 26245
rect 42 26164 76 26168
rect 42 26149 46 26164
rect 72 26149 76 26164
rect 38 26131 80 26149
rect 16 26125 102 26131
rect 144 26125 148 26277
rect 174 26253 181 26281
rect 224 26243 226 26290
rect 300 26281 308 26294
rect 278 26270 305 26281
rect 332 26253 342 26303
rect 400 26283 404 26303
rect 497 26299 500 26315
rect 596 26299 599 26315
rect 466 26298 500 26299
rect 442 26291 500 26298
rect 565 26291 599 26299
rect 612 26282 614 26332
rect 256 26243 328 26251
rect 336 26245 342 26253
rect 400 26245 404 26253
rect 196 26213 204 26243
rect 216 26213 232 26243
rect 196 26209 232 26213
rect 196 26201 226 26209
rect 224 26185 226 26201
rect 332 26173 336 26241
rect 400 26211 408 26245
rect 434 26211 438 26245
rect 454 26229 504 26231
rect 504 26213 506 26229
rect 514 26223 530 26229
rect 532 26223 548 26229
rect 525 26213 548 26222
rect 400 26203 404 26211
rect 498 26203 506 26213
rect 504 26179 506 26203
rect 514 26193 515 26213
rect 525 26188 528 26213
rect 547 26193 548 26213
rect 557 26203 564 26213
rect 514 26179 548 26183
rect 400 26173 442 26174
rect 174 26163 246 26171
rect 400 26166 404 26173
rect 295 26132 300 26166
rect 324 26132 329 26166
rect 367 26149 438 26166
rect 367 26132 442 26149
rect 400 26131 442 26132
rect 378 26125 464 26131
rect 38 26109 80 26125
rect 400 26109 442 26125
rect -25 26095 25 26097
rect 42 26095 76 26109
rect 404 26095 438 26109
rect 455 26095 505 26097
rect 557 26095 607 26097
rect 16 26087 102 26095
rect 378 26087 464 26095
rect 8 26053 17 26087
rect 18 26085 51 26087
rect 80 26085 100 26087
rect 18 26053 100 26085
rect 380 26085 404 26087
rect 429 26085 438 26087
rect 442 26085 462 26087
rect 16 26045 102 26053
rect 42 26029 76 26045
rect 16 26009 38 26015
rect 42 26006 76 26010
rect 80 26009 102 26015
rect 42 25976 46 26006
rect 72 25976 76 26006
rect 42 25895 46 25929
rect 72 25895 76 25929
rect -25 25858 25 25860
rect -8 25850 14 25857
rect -8 25849 17 25850
rect 25 25849 27 25858
rect -12 25842 38 25849
rect -12 25841 34 25842
rect -12 25837 8 25841
rect 0 25825 8 25837
rect 14 25825 34 25841
rect 0 25824 34 25825
rect 0 25817 38 25824
rect 14 25816 17 25817
rect 25 25808 27 25817
rect 42 25788 45 25878
rect 69 25863 80 25895
rect 107 25863 143 25891
rect 144 25863 148 26083
rect 332 26015 336 26083
rect 380 26053 462 26085
rect 463 26053 472 26087
rect 480 26053 497 26087
rect 378 26045 464 26053
rect 505 26045 507 26095
rect 514 26053 548 26087
rect 565 26053 582 26087
rect 607 26045 609 26095
rect 404 26029 438 26045
rect 400 26015 442 26016
rect 378 26009 404 26015
rect 442 26009 464 26015
rect 400 26008 404 26009
rect 174 25969 246 25977
rect 295 25974 300 26008
rect 324 25974 329 26008
rect 224 25939 226 25955
rect 196 25931 226 25939
rect 332 25937 336 26005
rect 367 25974 438 26008
rect 400 25967 404 25974
rect 454 25961 504 25963
rect 494 25957 548 25961
rect 494 25952 514 25957
rect 504 25937 506 25952
rect 196 25927 232 25931
rect 196 25897 204 25927
rect 216 25897 232 25927
rect 400 25929 404 25937
rect 107 25857 119 25863
rect 109 25829 119 25857
rect 129 25829 149 25863
rect 174 25859 181 25889
rect 224 25850 226 25897
rect 256 25889 328 25897
rect 332 25895 336 25925
rect 400 25895 408 25929
rect 434 25895 438 25929
rect 498 25927 506 25937
rect 514 25927 515 25947
rect 504 25911 506 25927
rect 525 25918 528 25952
rect 547 25927 548 25947
rect 557 25927 564 25937
rect 514 25911 530 25917
rect 532 25911 548 25917
rect 278 25859 305 25870
rect 42 25737 46 25771
rect 72 25737 76 25771
rect 38 25699 80 25700
rect 42 25658 76 25692
rect 79 25658 113 25692
rect 42 25579 46 25613
rect 72 25579 76 25613
rect -25 25542 25 25544
rect -8 25534 14 25541
rect -8 25533 17 25534
rect 25 25533 27 25542
rect -12 25526 38 25533
rect -12 25525 34 25526
rect -12 25521 8 25525
rect 0 25509 8 25521
rect 14 25509 34 25525
rect 0 25508 34 25509
rect 0 25501 38 25508
rect 14 25500 17 25501
rect 25 25492 27 25501
rect 42 25472 45 25562
rect 71 25531 80 25559
rect 69 25493 80 25531
rect 144 25521 148 25829
rect 196 25816 204 25850
rect 216 25816 232 25850
rect 244 25846 257 25850
rect 300 25846 308 25859
rect 332 25857 342 25895
rect 400 25887 404 25895
rect 336 25847 342 25857
rect 244 25822 291 25846
rect 244 25816 257 25822
rect 224 25769 226 25816
rect 278 25812 291 25822
rect 300 25822 329 25846
rect 332 25837 342 25847
rect 400 25847 409 25875
rect 562 25858 612 25860
rect 466 25849 497 25857
rect 565 25849 596 25857
rect 300 25812 321 25822
rect 300 25806 308 25812
rect 289 25796 308 25806
rect 196 25739 204 25769
rect 216 25739 232 25769
rect 196 25735 232 25739
rect 196 25727 226 25735
rect 300 25727 308 25796
rect 332 25803 351 25837
rect 361 25809 381 25837
rect 361 25803 375 25809
rect 400 25803 411 25847
rect 442 25842 500 25849
rect 466 25841 500 25842
rect 565 25841 599 25849
rect 497 25825 500 25841
rect 596 25825 599 25841
rect 466 25824 500 25825
rect 442 25817 500 25824
rect 565 25817 599 25825
rect 612 25808 614 25858
rect 332 25779 342 25803
rect 336 25767 342 25779
rect 224 25711 226 25727
rect 332 25699 342 25767
rect 400 25771 404 25779
rect 400 25737 408 25771
rect 434 25737 438 25771
rect 454 25755 504 25757
rect 504 25739 506 25755
rect 514 25749 530 25755
rect 532 25749 548 25755
rect 525 25739 548 25748
rect 400 25729 404 25737
rect 498 25729 506 25739
rect 504 25705 506 25729
rect 514 25719 515 25739
rect 525 25714 528 25739
rect 547 25719 548 25739
rect 557 25729 564 25739
rect 514 25705 548 25709
rect 151 25658 156 25692
rect 174 25689 246 25697
rect 256 25689 328 25697
rect 336 25691 342 25699
rect 400 25694 404 25699
rect 180 25661 185 25689
rect 174 25653 246 25661
rect 256 25653 328 25661
rect 332 25659 336 25689
rect 400 25660 438 25694
rect 224 25623 226 25639
rect 196 25615 226 25623
rect 196 25611 232 25615
rect 196 25581 204 25611
rect 216 25581 232 25611
rect 224 25534 226 25581
rect 300 25554 308 25623
rect 332 25621 342 25659
rect 400 25651 404 25660
rect 454 25645 504 25647
rect 494 25641 548 25645
rect 494 25636 514 25641
rect 504 25621 506 25636
rect 336 25609 342 25621
rect 289 25544 308 25554
rect 300 25538 308 25544
rect 332 25575 342 25609
rect 400 25613 404 25621
rect 400 25579 408 25613
rect 434 25579 438 25613
rect 498 25611 506 25621
rect 514 25611 515 25631
rect 504 25595 506 25611
rect 525 25602 528 25636
rect 547 25611 548 25631
rect 557 25611 564 25621
rect 514 25595 530 25601
rect 532 25595 548 25601
rect 332 25547 373 25575
rect 332 25541 351 25547
rect 107 25487 119 25521
rect 129 25487 149 25521
rect 196 25500 204 25534
rect 216 25500 232 25534
rect 244 25528 257 25534
rect 278 25528 291 25538
rect 244 25504 291 25528
rect 300 25528 321 25538
rect 336 25531 351 25541
rect 300 25504 329 25528
rect 332 25513 351 25531
rect 361 25541 375 25547
rect 400 25541 411 25579
rect 562 25542 612 25544
rect 361 25513 381 25541
rect 400 25513 409 25541
rect 466 25533 497 25541
rect 565 25533 596 25541
rect 442 25526 500 25533
rect 466 25525 500 25526
rect 565 25525 599 25533
rect 244 25500 257 25504
rect 42 25421 46 25455
rect 72 25421 76 25455
rect 42 25374 76 25378
rect 42 25359 46 25374
rect 72 25359 76 25374
rect 38 25341 80 25359
rect 16 25335 102 25341
rect 144 25335 148 25487
rect 174 25463 181 25491
rect 224 25453 226 25500
rect 300 25491 308 25504
rect 278 25480 305 25491
rect 332 25463 342 25513
rect 400 25493 404 25513
rect 497 25509 500 25525
rect 596 25509 599 25525
rect 466 25508 500 25509
rect 442 25501 500 25508
rect 565 25501 599 25509
rect 612 25492 614 25542
rect 256 25453 328 25461
rect 336 25455 342 25463
rect 400 25455 404 25463
rect 196 25423 204 25453
rect 216 25423 232 25453
rect 196 25419 232 25423
rect 196 25411 226 25419
rect 224 25395 226 25411
rect 332 25383 336 25451
rect 400 25421 408 25455
rect 434 25421 438 25455
rect 454 25439 504 25441
rect 504 25423 506 25439
rect 514 25433 530 25439
rect 532 25433 548 25439
rect 525 25423 548 25432
rect 400 25413 404 25421
rect 498 25413 506 25423
rect 504 25389 506 25413
rect 514 25403 515 25423
rect 525 25398 528 25423
rect 547 25403 548 25423
rect 557 25413 564 25423
rect 514 25389 548 25393
rect 400 25383 442 25384
rect 174 25373 246 25381
rect 400 25376 404 25383
rect 295 25342 300 25376
rect 324 25342 329 25376
rect 367 25359 438 25376
rect 367 25342 442 25359
rect 400 25341 442 25342
rect 378 25335 464 25341
rect 38 25319 80 25335
rect 400 25319 442 25335
rect -25 25305 25 25307
rect 42 25305 76 25319
rect 404 25305 438 25319
rect 455 25305 505 25307
rect 557 25305 607 25307
rect 16 25297 102 25305
rect 378 25297 464 25305
rect 8 25263 17 25297
rect 18 25295 51 25297
rect 80 25295 100 25297
rect 18 25263 100 25295
rect 380 25295 404 25297
rect 429 25295 438 25297
rect 442 25295 462 25297
rect 16 25255 102 25263
rect 42 25239 76 25255
rect 16 25219 38 25225
rect 42 25216 76 25220
rect 80 25219 102 25225
rect 42 25186 46 25216
rect 72 25186 76 25216
rect 42 25105 46 25139
rect 72 25105 76 25139
rect -25 25068 25 25070
rect -8 25060 14 25067
rect -8 25059 17 25060
rect 25 25059 27 25068
rect -12 25052 38 25059
rect -12 25051 34 25052
rect -12 25047 8 25051
rect 0 25035 8 25047
rect 14 25035 34 25051
rect 0 25034 34 25035
rect 0 25027 38 25034
rect 14 25026 17 25027
rect 25 25018 27 25027
rect 42 24998 45 25088
rect 69 25073 80 25105
rect 107 25073 143 25101
rect 144 25073 148 25293
rect 332 25225 336 25293
rect 380 25263 462 25295
rect 463 25263 472 25297
rect 480 25263 497 25297
rect 378 25255 464 25263
rect 505 25255 507 25305
rect 514 25263 548 25297
rect 565 25263 582 25297
rect 607 25255 609 25305
rect 404 25239 438 25255
rect 400 25225 442 25226
rect 378 25219 404 25225
rect 442 25219 464 25225
rect 400 25218 404 25219
rect 174 25179 246 25187
rect 295 25184 300 25218
rect 324 25184 329 25218
rect 224 25149 226 25165
rect 196 25141 226 25149
rect 332 25147 336 25215
rect 367 25184 438 25218
rect 400 25177 404 25184
rect 454 25171 504 25173
rect 494 25167 548 25171
rect 494 25162 514 25167
rect 504 25147 506 25162
rect 196 25137 232 25141
rect 196 25107 204 25137
rect 216 25107 232 25137
rect 400 25139 404 25147
rect 107 25067 119 25073
rect 109 25039 119 25067
rect 129 25039 149 25073
rect 174 25069 181 25099
rect 224 25060 226 25107
rect 256 25099 328 25107
rect 332 25105 336 25135
rect 400 25105 408 25139
rect 434 25105 438 25139
rect 498 25137 506 25147
rect 514 25137 515 25157
rect 504 25121 506 25137
rect 525 25128 528 25162
rect 547 25137 548 25157
rect 557 25137 564 25147
rect 514 25121 530 25127
rect 532 25121 548 25127
rect 278 25069 305 25080
rect 42 24947 46 24981
rect 72 24947 76 24981
rect 38 24909 80 24910
rect 42 24868 76 24902
rect 79 24868 113 24902
rect 42 24789 46 24823
rect 72 24789 76 24823
rect -25 24752 25 24754
rect -8 24744 14 24751
rect -8 24743 17 24744
rect 25 24743 27 24752
rect -12 24736 38 24743
rect -12 24735 34 24736
rect -12 24731 8 24735
rect 0 24719 8 24731
rect 14 24719 34 24735
rect 0 24718 34 24719
rect 0 24711 38 24718
rect 14 24710 17 24711
rect 25 24702 27 24711
rect 42 24682 45 24772
rect 71 24741 80 24769
rect 69 24703 80 24741
rect 144 24731 148 25039
rect 196 25026 204 25060
rect 216 25026 232 25060
rect 244 25056 257 25060
rect 300 25056 308 25069
rect 332 25067 342 25105
rect 400 25097 404 25105
rect 336 25057 342 25067
rect 244 25032 291 25056
rect 244 25026 257 25032
rect 224 24979 226 25026
rect 278 25022 291 25032
rect 300 25032 329 25056
rect 332 25047 342 25057
rect 400 25057 409 25085
rect 562 25068 612 25070
rect 466 25059 497 25067
rect 565 25059 596 25067
rect 300 25022 321 25032
rect 300 25016 308 25022
rect 289 25006 308 25016
rect 196 24949 204 24979
rect 216 24949 232 24979
rect 196 24945 232 24949
rect 196 24937 226 24945
rect 300 24937 308 25006
rect 332 25013 351 25047
rect 361 25019 381 25047
rect 361 25013 375 25019
rect 400 25013 411 25057
rect 442 25052 500 25059
rect 466 25051 500 25052
rect 565 25051 599 25059
rect 497 25035 500 25051
rect 596 25035 599 25051
rect 466 25034 500 25035
rect 442 25027 500 25034
rect 565 25027 599 25035
rect 612 25018 614 25068
rect 332 24989 342 25013
rect 336 24977 342 24989
rect 224 24921 226 24937
rect 332 24909 342 24977
rect 400 24981 404 24989
rect 400 24947 408 24981
rect 434 24947 438 24981
rect 454 24965 504 24967
rect 504 24949 506 24965
rect 514 24959 530 24965
rect 532 24959 548 24965
rect 525 24949 548 24958
rect 400 24939 404 24947
rect 498 24939 506 24949
rect 504 24915 506 24939
rect 514 24929 515 24949
rect 525 24924 528 24949
rect 547 24929 548 24949
rect 557 24939 564 24949
rect 514 24915 548 24919
rect 151 24868 156 24902
rect 174 24899 246 24907
rect 256 24899 328 24907
rect 336 24901 342 24909
rect 400 24904 404 24909
rect 180 24871 185 24899
rect 174 24863 246 24871
rect 256 24863 328 24871
rect 332 24869 336 24899
rect 400 24870 438 24904
rect 224 24833 226 24849
rect 196 24825 226 24833
rect 196 24821 232 24825
rect 196 24791 204 24821
rect 216 24791 232 24821
rect 224 24744 226 24791
rect 300 24764 308 24833
rect 332 24831 342 24869
rect 400 24861 404 24870
rect 454 24855 504 24857
rect 494 24851 548 24855
rect 494 24846 514 24851
rect 504 24831 506 24846
rect 336 24819 342 24831
rect 289 24754 308 24764
rect 300 24748 308 24754
rect 332 24785 342 24819
rect 400 24823 404 24831
rect 400 24789 408 24823
rect 434 24789 438 24823
rect 498 24821 506 24831
rect 514 24821 515 24841
rect 504 24805 506 24821
rect 525 24812 528 24846
rect 547 24821 548 24841
rect 557 24821 564 24831
rect 514 24805 530 24811
rect 532 24805 548 24811
rect 332 24757 373 24785
rect 332 24751 351 24757
rect 107 24697 119 24731
rect 129 24697 149 24731
rect 196 24710 204 24744
rect 216 24710 232 24744
rect 244 24738 257 24744
rect 278 24738 291 24748
rect 244 24714 291 24738
rect 300 24738 321 24748
rect 336 24741 351 24751
rect 300 24714 329 24738
rect 332 24723 351 24741
rect 361 24751 375 24757
rect 400 24751 411 24789
rect 562 24752 612 24754
rect 361 24723 381 24751
rect 400 24723 409 24751
rect 466 24743 497 24751
rect 565 24743 596 24751
rect 442 24736 500 24743
rect 466 24735 500 24736
rect 565 24735 599 24743
rect 244 24710 257 24714
rect 42 24631 46 24665
rect 72 24631 76 24665
rect 42 24584 76 24588
rect 42 24569 46 24584
rect 72 24569 76 24584
rect 38 24551 80 24569
rect 16 24545 102 24551
rect 144 24545 148 24697
rect 174 24673 181 24701
rect 224 24663 226 24710
rect 300 24701 308 24714
rect 278 24690 305 24701
rect 332 24673 342 24723
rect 400 24703 404 24723
rect 497 24719 500 24735
rect 596 24719 599 24735
rect 466 24718 500 24719
rect 442 24711 500 24718
rect 565 24711 599 24719
rect 612 24702 614 24752
rect 256 24663 328 24671
rect 336 24665 342 24673
rect 400 24665 404 24673
rect 196 24633 204 24663
rect 216 24633 232 24663
rect 196 24629 232 24633
rect 196 24621 226 24629
rect 224 24605 226 24621
rect 332 24593 336 24661
rect 400 24631 408 24665
rect 434 24631 438 24665
rect 454 24649 504 24651
rect 504 24633 506 24649
rect 514 24643 530 24649
rect 532 24643 548 24649
rect 525 24633 548 24642
rect 400 24623 404 24631
rect 498 24623 506 24633
rect 504 24599 506 24623
rect 514 24613 515 24633
rect 525 24608 528 24633
rect 547 24613 548 24633
rect 557 24623 564 24633
rect 514 24599 548 24603
rect 400 24593 442 24594
rect 174 24583 246 24591
rect 400 24586 404 24593
rect 295 24552 300 24586
rect 324 24552 329 24586
rect 367 24569 438 24586
rect 367 24552 442 24569
rect 400 24551 442 24552
rect 378 24545 464 24551
rect 38 24529 80 24545
rect 400 24529 442 24545
rect -25 24515 25 24517
rect 42 24515 76 24529
rect 404 24515 438 24529
rect 455 24515 505 24517
rect 557 24515 607 24517
rect 16 24507 102 24515
rect 378 24507 464 24515
rect 8 24473 17 24507
rect 18 24505 51 24507
rect 80 24505 100 24507
rect 18 24473 100 24505
rect 380 24505 404 24507
rect 429 24505 438 24507
rect 442 24505 462 24507
rect 16 24465 102 24473
rect 42 24449 76 24465
rect 16 24429 38 24435
rect 42 24426 76 24430
rect 80 24429 102 24435
rect 42 24396 46 24426
rect 72 24396 76 24426
rect 42 24315 46 24349
rect 72 24315 76 24349
rect -25 24278 25 24280
rect -8 24270 14 24277
rect -8 24269 17 24270
rect 25 24269 27 24278
rect -12 24262 38 24269
rect -12 24261 34 24262
rect -12 24257 8 24261
rect 0 24245 8 24257
rect 14 24245 34 24261
rect 0 24244 34 24245
rect 0 24237 38 24244
rect 14 24236 17 24237
rect 25 24228 27 24237
rect 42 24208 45 24298
rect 69 24283 80 24315
rect 107 24283 143 24311
rect 144 24283 148 24503
rect 332 24435 336 24503
rect 380 24473 462 24505
rect 463 24473 472 24507
rect 480 24473 497 24507
rect 378 24465 464 24473
rect 505 24465 507 24515
rect 514 24473 548 24507
rect 565 24473 582 24507
rect 607 24465 609 24515
rect 404 24449 438 24465
rect 400 24435 442 24436
rect 378 24429 404 24435
rect 442 24429 464 24435
rect 400 24428 404 24429
rect 174 24389 246 24397
rect 295 24394 300 24428
rect 324 24394 329 24428
rect 224 24359 226 24375
rect 196 24351 226 24359
rect 332 24357 336 24425
rect 367 24394 438 24428
rect 400 24387 404 24394
rect 454 24381 504 24383
rect 494 24377 548 24381
rect 494 24372 514 24377
rect 504 24357 506 24372
rect 196 24347 232 24351
rect 196 24317 204 24347
rect 216 24317 232 24347
rect 400 24349 404 24357
rect 107 24277 119 24283
rect 109 24249 119 24277
rect 129 24249 149 24283
rect 174 24279 181 24309
rect 224 24270 226 24317
rect 256 24309 328 24317
rect 332 24315 336 24345
rect 400 24315 408 24349
rect 434 24315 438 24349
rect 498 24347 506 24357
rect 514 24347 515 24367
rect 504 24331 506 24347
rect 525 24338 528 24372
rect 547 24347 548 24367
rect 557 24347 564 24357
rect 514 24331 530 24337
rect 532 24331 548 24337
rect 278 24279 305 24290
rect 42 24157 46 24191
rect 72 24157 76 24191
rect 38 24119 80 24120
rect 42 24078 76 24112
rect 79 24078 113 24112
rect 42 23999 46 24033
rect 72 23999 76 24033
rect -25 23962 25 23964
rect -8 23954 14 23961
rect -8 23953 17 23954
rect 25 23953 27 23962
rect -12 23946 38 23953
rect -12 23945 34 23946
rect -12 23941 8 23945
rect 0 23929 8 23941
rect 14 23929 34 23945
rect 0 23928 34 23929
rect 0 23921 38 23928
rect 14 23920 17 23921
rect 25 23912 27 23921
rect 42 23892 45 23982
rect 71 23951 80 23979
rect 69 23913 80 23951
rect 144 23941 148 24249
rect 196 24236 204 24270
rect 216 24236 232 24270
rect 244 24266 257 24270
rect 300 24266 308 24279
rect 332 24277 342 24315
rect 400 24307 404 24315
rect 336 24267 342 24277
rect 244 24242 291 24266
rect 244 24236 257 24242
rect 224 24189 226 24236
rect 278 24232 291 24242
rect 300 24242 329 24266
rect 332 24257 342 24267
rect 400 24267 409 24295
rect 562 24278 612 24280
rect 466 24269 497 24277
rect 565 24269 596 24277
rect 300 24232 321 24242
rect 300 24226 308 24232
rect 289 24216 308 24226
rect 196 24159 204 24189
rect 216 24159 232 24189
rect 196 24155 232 24159
rect 196 24147 226 24155
rect 300 24147 308 24216
rect 332 24223 351 24257
rect 361 24229 381 24257
rect 361 24223 375 24229
rect 400 24223 411 24267
rect 442 24262 500 24269
rect 466 24261 500 24262
rect 565 24261 599 24269
rect 497 24245 500 24261
rect 596 24245 599 24261
rect 466 24244 500 24245
rect 442 24237 500 24244
rect 565 24237 599 24245
rect 612 24228 614 24278
rect 332 24199 342 24223
rect 336 24187 342 24199
rect 224 24131 226 24147
rect 332 24119 342 24187
rect 400 24191 404 24199
rect 400 24157 408 24191
rect 434 24157 438 24191
rect 454 24175 504 24177
rect 504 24159 506 24175
rect 514 24169 530 24175
rect 532 24169 548 24175
rect 525 24159 548 24168
rect 400 24149 404 24157
rect 498 24149 506 24159
rect 504 24125 506 24149
rect 514 24139 515 24159
rect 525 24134 528 24159
rect 547 24139 548 24159
rect 557 24149 564 24159
rect 514 24125 548 24129
rect 151 24078 156 24112
rect 174 24109 246 24117
rect 256 24109 328 24117
rect 336 24111 342 24119
rect 400 24114 404 24119
rect 180 24081 185 24109
rect 174 24073 246 24081
rect 256 24073 328 24081
rect 332 24079 336 24109
rect 400 24080 438 24114
rect 224 24043 226 24059
rect 196 24035 226 24043
rect 196 24031 232 24035
rect 196 24001 204 24031
rect 216 24001 232 24031
rect 224 23954 226 24001
rect 300 23974 308 24043
rect 332 24041 342 24079
rect 400 24071 404 24080
rect 454 24065 504 24067
rect 494 24061 548 24065
rect 494 24056 514 24061
rect 504 24041 506 24056
rect 336 24029 342 24041
rect 289 23964 308 23974
rect 300 23958 308 23964
rect 332 23995 342 24029
rect 400 24033 404 24041
rect 400 23999 408 24033
rect 434 23999 438 24033
rect 498 24031 506 24041
rect 514 24031 515 24051
rect 504 24015 506 24031
rect 525 24022 528 24056
rect 547 24031 548 24051
rect 557 24031 564 24041
rect 514 24015 530 24021
rect 532 24015 548 24021
rect 332 23967 373 23995
rect 332 23961 351 23967
rect 107 23907 119 23941
rect 129 23907 149 23941
rect 196 23920 204 23954
rect 216 23920 232 23954
rect 244 23948 257 23954
rect 278 23948 291 23958
rect 244 23924 291 23948
rect 300 23948 321 23958
rect 336 23951 351 23961
rect 300 23924 329 23948
rect 332 23933 351 23951
rect 361 23961 375 23967
rect 400 23961 411 23999
rect 562 23962 612 23964
rect 361 23933 381 23961
rect 400 23933 409 23961
rect 466 23953 497 23961
rect 565 23953 596 23961
rect 442 23946 500 23953
rect 466 23945 500 23946
rect 565 23945 599 23953
rect 244 23920 257 23924
rect 42 23841 46 23875
rect 72 23841 76 23875
rect 42 23794 76 23798
rect 42 23779 46 23794
rect 72 23779 76 23794
rect 38 23761 80 23779
rect 16 23755 102 23761
rect 144 23755 148 23907
rect 174 23883 181 23911
rect 224 23873 226 23920
rect 300 23911 308 23924
rect 278 23900 305 23911
rect 332 23883 342 23933
rect 400 23913 404 23933
rect 497 23929 500 23945
rect 596 23929 599 23945
rect 466 23928 500 23929
rect 442 23921 500 23928
rect 565 23921 599 23929
rect 612 23912 614 23962
rect 256 23873 328 23881
rect 336 23875 342 23883
rect 400 23875 404 23883
rect 196 23843 204 23873
rect 216 23843 232 23873
rect 196 23839 232 23843
rect 196 23831 226 23839
rect 224 23815 226 23831
rect 332 23803 336 23871
rect 400 23841 408 23875
rect 434 23841 438 23875
rect 454 23859 504 23861
rect 504 23843 506 23859
rect 514 23853 530 23859
rect 532 23853 548 23859
rect 525 23843 548 23852
rect 400 23833 404 23841
rect 498 23833 506 23843
rect 504 23809 506 23833
rect 514 23823 515 23843
rect 525 23818 528 23843
rect 547 23823 548 23843
rect 557 23833 564 23843
rect 514 23809 548 23813
rect 400 23803 442 23804
rect 174 23793 246 23801
rect 400 23796 404 23803
rect 295 23762 300 23796
rect 324 23762 329 23796
rect 367 23779 438 23796
rect 367 23762 442 23779
rect 400 23761 442 23762
rect 378 23755 464 23761
rect 38 23739 80 23755
rect 400 23739 442 23755
rect -25 23725 25 23727
rect 42 23725 76 23739
rect 404 23725 438 23739
rect 455 23725 505 23727
rect 557 23725 607 23727
rect 16 23717 102 23725
rect 378 23717 464 23725
rect 8 23683 17 23717
rect 18 23715 51 23717
rect 80 23715 100 23717
rect 18 23683 100 23715
rect 380 23715 404 23717
rect 429 23715 438 23717
rect 442 23715 462 23717
rect 16 23675 102 23683
rect 42 23659 76 23675
rect 16 23639 38 23645
rect 42 23636 76 23640
rect 80 23639 102 23645
rect 42 23606 46 23636
rect 72 23606 76 23636
rect 42 23525 46 23559
rect 72 23525 76 23559
rect -25 23488 25 23490
rect -8 23480 14 23487
rect -8 23479 17 23480
rect 25 23479 27 23488
rect -12 23472 38 23479
rect -12 23471 34 23472
rect -12 23467 8 23471
rect 0 23455 8 23467
rect 14 23455 34 23471
rect 0 23454 34 23455
rect 0 23447 38 23454
rect 14 23446 17 23447
rect 25 23438 27 23447
rect 42 23418 45 23508
rect 69 23493 80 23525
rect 107 23493 143 23521
rect 144 23493 148 23713
rect 332 23645 336 23713
rect 380 23683 462 23715
rect 463 23683 472 23717
rect 480 23683 497 23717
rect 378 23675 464 23683
rect 505 23675 507 23725
rect 514 23683 548 23717
rect 565 23683 582 23717
rect 607 23675 609 23725
rect 404 23659 438 23675
rect 400 23645 442 23646
rect 378 23639 404 23645
rect 442 23639 464 23645
rect 400 23638 404 23639
rect 174 23599 246 23607
rect 295 23604 300 23638
rect 324 23604 329 23638
rect 224 23569 226 23585
rect 196 23561 226 23569
rect 332 23567 336 23635
rect 367 23604 438 23638
rect 400 23597 404 23604
rect 454 23591 504 23593
rect 494 23587 548 23591
rect 494 23582 514 23587
rect 504 23567 506 23582
rect 196 23557 232 23561
rect 196 23527 204 23557
rect 216 23527 232 23557
rect 400 23559 404 23567
rect 107 23487 119 23493
rect 109 23459 119 23487
rect 129 23459 149 23493
rect 174 23489 181 23519
rect 224 23480 226 23527
rect 256 23519 328 23527
rect 332 23525 336 23555
rect 400 23525 408 23559
rect 434 23525 438 23559
rect 498 23557 506 23567
rect 514 23557 515 23577
rect 504 23541 506 23557
rect 525 23548 528 23582
rect 547 23557 548 23577
rect 557 23557 564 23567
rect 514 23541 530 23547
rect 532 23541 548 23547
rect 278 23489 305 23500
rect 42 23367 46 23401
rect 72 23367 76 23401
rect 38 23329 80 23330
rect 42 23288 76 23322
rect 79 23288 113 23322
rect 42 23209 46 23243
rect 72 23209 76 23243
rect -25 23172 25 23174
rect -8 23164 14 23171
rect -8 23163 17 23164
rect 25 23163 27 23172
rect -12 23156 38 23163
rect -12 23155 34 23156
rect -12 23151 8 23155
rect 0 23139 8 23151
rect 14 23139 34 23155
rect 0 23138 34 23139
rect 0 23131 38 23138
rect 14 23130 17 23131
rect 25 23122 27 23131
rect 42 23102 45 23192
rect 71 23161 80 23189
rect 69 23123 80 23161
rect 144 23151 148 23459
rect 196 23446 204 23480
rect 216 23446 232 23480
rect 244 23476 257 23480
rect 300 23476 308 23489
rect 332 23487 342 23525
rect 400 23517 404 23525
rect 336 23477 342 23487
rect 244 23452 291 23476
rect 244 23446 257 23452
rect 224 23399 226 23446
rect 278 23442 291 23452
rect 300 23452 329 23476
rect 332 23467 342 23477
rect 400 23477 409 23505
rect 562 23488 612 23490
rect 466 23479 497 23487
rect 565 23479 596 23487
rect 300 23442 321 23452
rect 300 23436 308 23442
rect 289 23426 308 23436
rect 196 23369 204 23399
rect 216 23369 232 23399
rect 196 23365 232 23369
rect 196 23357 226 23365
rect 300 23357 308 23426
rect 332 23433 351 23467
rect 361 23439 381 23467
rect 361 23433 375 23439
rect 400 23433 411 23477
rect 442 23472 500 23479
rect 466 23471 500 23472
rect 565 23471 599 23479
rect 497 23455 500 23471
rect 596 23455 599 23471
rect 466 23454 500 23455
rect 442 23447 500 23454
rect 565 23447 599 23455
rect 612 23438 614 23488
rect 332 23409 342 23433
rect 336 23397 342 23409
rect 224 23341 226 23357
rect 332 23329 342 23397
rect 400 23401 404 23409
rect 400 23367 408 23401
rect 434 23367 438 23401
rect 454 23385 504 23387
rect 504 23369 506 23385
rect 514 23379 530 23385
rect 532 23379 548 23385
rect 525 23369 548 23378
rect 400 23359 404 23367
rect 498 23359 506 23369
rect 504 23335 506 23359
rect 514 23349 515 23369
rect 525 23344 528 23369
rect 547 23349 548 23369
rect 557 23359 564 23369
rect 514 23335 548 23339
rect 151 23288 156 23322
rect 174 23319 246 23327
rect 256 23319 328 23327
rect 336 23321 342 23329
rect 400 23324 404 23329
rect 180 23291 185 23319
rect 174 23283 246 23291
rect 256 23283 328 23291
rect 332 23289 336 23319
rect 400 23290 438 23324
rect 224 23253 226 23269
rect 196 23245 226 23253
rect 196 23241 232 23245
rect 196 23211 204 23241
rect 216 23211 232 23241
rect 224 23164 226 23211
rect 300 23184 308 23253
rect 332 23251 342 23289
rect 400 23281 404 23290
rect 454 23275 504 23277
rect 494 23271 548 23275
rect 494 23266 514 23271
rect 504 23251 506 23266
rect 336 23239 342 23251
rect 289 23174 308 23184
rect 300 23168 308 23174
rect 332 23205 342 23239
rect 400 23243 404 23251
rect 400 23209 408 23243
rect 434 23209 438 23243
rect 498 23241 506 23251
rect 514 23241 515 23261
rect 504 23225 506 23241
rect 525 23232 528 23266
rect 547 23241 548 23261
rect 557 23241 564 23251
rect 514 23225 530 23231
rect 532 23225 548 23231
rect 332 23177 373 23205
rect 332 23171 351 23177
rect 107 23117 119 23151
rect 129 23117 149 23151
rect 196 23130 204 23164
rect 216 23130 232 23164
rect 244 23158 257 23164
rect 278 23158 291 23168
rect 244 23134 291 23158
rect 300 23158 321 23168
rect 336 23161 351 23171
rect 300 23134 329 23158
rect 332 23143 351 23161
rect 361 23171 375 23177
rect 400 23171 411 23209
rect 562 23172 612 23174
rect 361 23143 381 23171
rect 400 23143 409 23171
rect 466 23163 497 23171
rect 565 23163 596 23171
rect 442 23156 500 23163
rect 466 23155 500 23156
rect 565 23155 599 23163
rect 244 23130 257 23134
rect 42 23051 46 23085
rect 72 23051 76 23085
rect 42 23004 76 23008
rect 42 22989 46 23004
rect 72 22989 76 23004
rect 38 22971 80 22989
rect 16 22965 102 22971
rect 144 22965 148 23117
rect 174 23093 181 23121
rect 224 23083 226 23130
rect 300 23121 308 23134
rect 278 23110 305 23121
rect 332 23093 342 23143
rect 400 23123 404 23143
rect 497 23139 500 23155
rect 596 23139 599 23155
rect 466 23138 500 23139
rect 442 23131 500 23138
rect 565 23131 599 23139
rect 612 23122 614 23172
rect 256 23083 328 23091
rect 336 23085 342 23093
rect 400 23085 404 23093
rect 196 23053 204 23083
rect 216 23053 232 23083
rect 196 23049 232 23053
rect 196 23041 226 23049
rect 224 23025 226 23041
rect 332 23013 336 23081
rect 400 23051 408 23085
rect 434 23051 438 23085
rect 454 23069 504 23071
rect 504 23053 506 23069
rect 514 23063 530 23069
rect 532 23063 548 23069
rect 525 23053 548 23062
rect 400 23043 404 23051
rect 498 23043 506 23053
rect 504 23019 506 23043
rect 514 23033 515 23053
rect 525 23028 528 23053
rect 547 23033 548 23053
rect 557 23043 564 23053
rect 514 23019 548 23023
rect 400 23013 442 23014
rect 174 23003 246 23011
rect 400 23006 404 23013
rect 295 22972 300 23006
rect 324 22972 329 23006
rect 367 22989 438 23006
rect 367 22972 442 22989
rect 400 22971 442 22972
rect 378 22965 464 22971
rect 38 22949 80 22965
rect 400 22949 442 22965
rect -25 22935 25 22937
rect 42 22935 76 22949
rect 404 22935 438 22949
rect 455 22935 505 22937
rect 557 22935 607 22937
rect 16 22927 102 22935
rect 378 22927 464 22935
rect 8 22893 17 22927
rect 18 22925 51 22927
rect 80 22925 100 22927
rect 18 22893 100 22925
rect 380 22925 404 22927
rect 429 22925 438 22927
rect 442 22925 462 22927
rect 16 22885 102 22893
rect 42 22869 76 22885
rect 16 22849 38 22855
rect 42 22846 76 22850
rect 80 22849 102 22855
rect 42 22816 46 22846
rect 72 22816 76 22846
rect 42 22735 46 22769
rect 72 22735 76 22769
rect -25 22698 25 22700
rect -8 22690 14 22697
rect -8 22689 17 22690
rect 25 22689 27 22698
rect -12 22682 38 22689
rect -12 22681 34 22682
rect -12 22677 8 22681
rect 0 22665 8 22677
rect 14 22665 34 22681
rect 0 22664 34 22665
rect 0 22657 38 22664
rect 14 22656 17 22657
rect 25 22648 27 22657
rect 42 22628 45 22718
rect 69 22703 80 22735
rect 107 22703 143 22731
rect 144 22703 148 22923
rect 332 22855 336 22923
rect 380 22893 462 22925
rect 463 22893 472 22927
rect 480 22893 497 22927
rect 378 22885 464 22893
rect 505 22885 507 22935
rect 514 22893 548 22927
rect 565 22893 582 22927
rect 607 22885 609 22935
rect 404 22869 438 22885
rect 400 22855 442 22856
rect 378 22849 404 22855
rect 442 22849 464 22855
rect 400 22848 404 22849
rect 174 22809 246 22817
rect 295 22814 300 22848
rect 324 22814 329 22848
rect 224 22779 226 22795
rect 196 22771 226 22779
rect 332 22777 336 22845
rect 367 22814 438 22848
rect 400 22807 404 22814
rect 454 22801 504 22803
rect 494 22797 548 22801
rect 494 22792 514 22797
rect 504 22777 506 22792
rect 196 22767 232 22771
rect 196 22737 204 22767
rect 216 22737 232 22767
rect 400 22769 404 22777
rect 107 22697 119 22703
rect 109 22669 119 22697
rect 129 22669 149 22703
rect 174 22699 181 22729
rect 224 22690 226 22737
rect 256 22729 328 22737
rect 332 22735 336 22765
rect 400 22735 408 22769
rect 434 22735 438 22769
rect 498 22767 506 22777
rect 514 22767 515 22787
rect 504 22751 506 22767
rect 525 22758 528 22792
rect 547 22767 548 22787
rect 557 22767 564 22777
rect 514 22751 530 22757
rect 532 22751 548 22757
rect 278 22699 305 22710
rect 42 22577 46 22611
rect 72 22577 76 22611
rect 38 22539 80 22540
rect 42 22498 76 22532
rect 79 22498 113 22532
rect 42 22419 46 22453
rect 72 22419 76 22453
rect -25 22382 25 22384
rect -8 22374 14 22381
rect -8 22373 17 22374
rect 25 22373 27 22382
rect -12 22366 38 22373
rect -12 22365 34 22366
rect -12 22361 8 22365
rect 0 22349 8 22361
rect 14 22349 34 22365
rect 0 22348 34 22349
rect 0 22341 38 22348
rect 14 22340 17 22341
rect 25 22332 27 22341
rect 42 22312 45 22402
rect 71 22371 80 22399
rect 69 22333 80 22371
rect 144 22361 148 22669
rect 196 22656 204 22690
rect 216 22656 232 22690
rect 244 22686 257 22690
rect 300 22686 308 22699
rect 332 22697 342 22735
rect 400 22727 404 22735
rect 336 22687 342 22697
rect 244 22662 291 22686
rect 244 22656 257 22662
rect 224 22609 226 22656
rect 278 22652 291 22662
rect 300 22662 329 22686
rect 332 22677 342 22687
rect 400 22687 409 22715
rect 562 22698 612 22700
rect 466 22689 497 22697
rect 565 22689 596 22697
rect 300 22652 321 22662
rect 300 22646 308 22652
rect 289 22636 308 22646
rect 196 22579 204 22609
rect 216 22579 232 22609
rect 196 22575 232 22579
rect 196 22567 226 22575
rect 300 22567 308 22636
rect 332 22643 351 22677
rect 361 22649 381 22677
rect 361 22643 375 22649
rect 400 22643 411 22687
rect 442 22682 500 22689
rect 466 22681 500 22682
rect 565 22681 599 22689
rect 497 22665 500 22681
rect 596 22665 599 22681
rect 466 22664 500 22665
rect 442 22657 500 22664
rect 565 22657 599 22665
rect 612 22648 614 22698
rect 332 22619 342 22643
rect 336 22607 342 22619
rect 224 22551 226 22567
rect 332 22539 342 22607
rect 400 22611 404 22619
rect 400 22577 408 22611
rect 434 22577 438 22611
rect 454 22595 504 22597
rect 504 22579 506 22595
rect 514 22589 530 22595
rect 532 22589 548 22595
rect 525 22579 548 22588
rect 400 22569 404 22577
rect 498 22569 506 22579
rect 504 22545 506 22569
rect 514 22559 515 22579
rect 525 22554 528 22579
rect 547 22559 548 22579
rect 557 22569 564 22579
rect 514 22545 548 22549
rect 151 22498 156 22532
rect 174 22529 246 22537
rect 256 22529 328 22537
rect 336 22531 342 22539
rect 400 22534 404 22539
rect 180 22501 185 22529
rect 174 22493 246 22501
rect 256 22493 328 22501
rect 332 22499 336 22529
rect 400 22500 438 22534
rect 224 22463 226 22479
rect 196 22455 226 22463
rect 196 22451 232 22455
rect 196 22421 204 22451
rect 216 22421 232 22451
rect 224 22374 226 22421
rect 300 22394 308 22463
rect 332 22461 342 22499
rect 400 22491 404 22500
rect 454 22485 504 22487
rect 494 22481 548 22485
rect 494 22476 514 22481
rect 504 22461 506 22476
rect 336 22449 342 22461
rect 289 22384 308 22394
rect 300 22378 308 22384
rect 332 22415 342 22449
rect 400 22453 404 22461
rect 400 22419 408 22453
rect 434 22419 438 22453
rect 498 22451 506 22461
rect 514 22451 515 22471
rect 504 22435 506 22451
rect 525 22442 528 22476
rect 547 22451 548 22471
rect 557 22451 564 22461
rect 514 22435 530 22441
rect 532 22435 548 22441
rect 332 22387 373 22415
rect 332 22381 351 22387
rect 107 22327 119 22361
rect 129 22327 149 22361
rect 196 22340 204 22374
rect 216 22340 232 22374
rect 244 22368 257 22374
rect 278 22368 291 22378
rect 244 22344 291 22368
rect 300 22368 321 22378
rect 336 22371 351 22381
rect 300 22344 329 22368
rect 332 22353 351 22371
rect 361 22381 375 22387
rect 400 22381 411 22419
rect 562 22382 612 22384
rect 361 22353 381 22381
rect 400 22353 409 22381
rect 466 22373 497 22381
rect 565 22373 596 22381
rect 442 22366 500 22373
rect 466 22365 500 22366
rect 565 22365 599 22373
rect 244 22340 257 22344
rect 42 22261 46 22295
rect 72 22261 76 22295
rect 42 22214 76 22218
rect 42 22199 46 22214
rect 72 22199 76 22214
rect 38 22181 80 22199
rect 16 22175 102 22181
rect 144 22175 148 22327
rect 174 22303 181 22331
rect 224 22293 226 22340
rect 300 22331 308 22344
rect 278 22320 305 22331
rect 332 22303 342 22353
rect 400 22333 404 22353
rect 497 22349 500 22365
rect 596 22349 599 22365
rect 466 22348 500 22349
rect 442 22341 500 22348
rect 565 22341 599 22349
rect 612 22332 614 22382
rect 256 22293 328 22301
rect 336 22295 342 22303
rect 400 22295 404 22303
rect 196 22263 204 22293
rect 216 22263 232 22293
rect 196 22259 232 22263
rect 196 22251 226 22259
rect 224 22235 226 22251
rect 332 22223 336 22291
rect 400 22261 408 22295
rect 434 22261 438 22295
rect 454 22279 504 22281
rect 504 22263 506 22279
rect 514 22273 530 22279
rect 532 22273 548 22279
rect 525 22263 548 22272
rect 400 22253 404 22261
rect 498 22253 506 22263
rect 504 22229 506 22253
rect 514 22243 515 22263
rect 525 22238 528 22263
rect 547 22243 548 22263
rect 557 22253 564 22263
rect 514 22229 548 22233
rect 400 22223 442 22224
rect 174 22213 246 22221
rect 400 22216 404 22223
rect 295 22182 300 22216
rect 324 22182 329 22216
rect 367 22199 438 22216
rect 367 22182 442 22199
rect 400 22181 442 22182
rect 378 22175 464 22181
rect 38 22159 80 22175
rect 400 22159 442 22175
rect -25 22145 25 22147
rect 42 22145 76 22159
rect 404 22145 438 22159
rect 455 22145 505 22147
rect 557 22145 607 22147
rect 16 22137 102 22145
rect 378 22137 464 22145
rect 8 22103 17 22137
rect 18 22135 51 22137
rect 80 22135 100 22137
rect 18 22103 100 22135
rect 380 22135 404 22137
rect 429 22135 438 22137
rect 442 22135 462 22137
rect 16 22095 102 22103
rect 42 22079 76 22095
rect 16 22059 38 22065
rect 42 22056 76 22060
rect 80 22059 102 22065
rect 42 22026 46 22056
rect 72 22026 76 22056
rect 42 21945 46 21979
rect 72 21945 76 21979
rect -25 21908 25 21910
rect -8 21900 14 21907
rect -8 21899 17 21900
rect 25 21899 27 21908
rect -12 21892 38 21899
rect -12 21891 34 21892
rect -12 21887 8 21891
rect 0 21875 8 21887
rect 14 21875 34 21891
rect 0 21874 34 21875
rect 0 21867 38 21874
rect 14 21866 17 21867
rect 25 21858 27 21867
rect 42 21838 45 21928
rect 69 21913 80 21945
rect 107 21913 143 21941
rect 144 21913 148 22133
rect 332 22065 336 22133
rect 380 22103 462 22135
rect 463 22103 472 22137
rect 480 22103 497 22137
rect 378 22095 464 22103
rect 505 22095 507 22145
rect 514 22103 548 22137
rect 565 22103 582 22137
rect 607 22095 609 22145
rect 404 22079 438 22095
rect 400 22065 442 22066
rect 378 22059 404 22065
rect 442 22059 464 22065
rect 400 22058 404 22059
rect 174 22019 246 22027
rect 295 22024 300 22058
rect 324 22024 329 22058
rect 224 21989 226 22005
rect 196 21981 226 21989
rect 332 21987 336 22055
rect 367 22024 438 22058
rect 400 22017 404 22024
rect 454 22011 504 22013
rect 494 22007 548 22011
rect 494 22002 514 22007
rect 504 21987 506 22002
rect 196 21977 232 21981
rect 196 21947 204 21977
rect 216 21947 232 21977
rect 400 21979 404 21987
rect 107 21907 119 21913
rect 109 21879 119 21907
rect 129 21879 149 21913
rect 174 21909 181 21939
rect 224 21900 226 21947
rect 256 21939 328 21947
rect 332 21945 336 21975
rect 400 21945 408 21979
rect 434 21945 438 21979
rect 498 21977 506 21987
rect 514 21977 515 21997
rect 504 21961 506 21977
rect 525 21968 528 22002
rect 547 21977 548 21997
rect 557 21977 564 21987
rect 514 21961 530 21967
rect 532 21961 548 21967
rect 278 21909 305 21920
rect 42 21787 46 21821
rect 72 21787 76 21821
rect 38 21749 80 21750
rect 42 21708 76 21742
rect 79 21708 113 21742
rect 42 21629 46 21663
rect 72 21629 76 21663
rect -25 21592 25 21594
rect -8 21584 14 21591
rect -8 21583 17 21584
rect 25 21583 27 21592
rect -12 21576 38 21583
rect -12 21575 34 21576
rect -12 21571 8 21575
rect 0 21559 8 21571
rect 14 21559 34 21575
rect 0 21558 34 21559
rect 0 21551 38 21558
rect 14 21550 17 21551
rect 25 21542 27 21551
rect 42 21522 45 21612
rect 71 21581 80 21609
rect 69 21543 80 21581
rect 144 21571 148 21879
rect 196 21866 204 21900
rect 216 21866 232 21900
rect 244 21896 257 21900
rect 300 21896 308 21909
rect 332 21907 342 21945
rect 400 21937 404 21945
rect 336 21897 342 21907
rect 244 21872 291 21896
rect 244 21866 257 21872
rect 224 21819 226 21866
rect 278 21862 291 21872
rect 300 21872 329 21896
rect 332 21887 342 21897
rect 400 21897 409 21925
rect 562 21908 612 21910
rect 466 21899 497 21907
rect 565 21899 596 21907
rect 300 21862 321 21872
rect 300 21856 308 21862
rect 289 21846 308 21856
rect 196 21789 204 21819
rect 216 21789 232 21819
rect 196 21785 232 21789
rect 196 21777 226 21785
rect 300 21777 308 21846
rect 332 21853 351 21887
rect 361 21859 381 21887
rect 361 21853 375 21859
rect 400 21853 411 21897
rect 442 21892 500 21899
rect 466 21891 500 21892
rect 565 21891 599 21899
rect 497 21875 500 21891
rect 596 21875 599 21891
rect 466 21874 500 21875
rect 442 21867 500 21874
rect 565 21867 599 21875
rect 612 21858 614 21908
rect 332 21829 342 21853
rect 336 21817 342 21829
rect 224 21761 226 21777
rect 332 21749 342 21817
rect 400 21821 404 21829
rect 400 21787 408 21821
rect 434 21787 438 21821
rect 454 21805 504 21807
rect 504 21789 506 21805
rect 514 21799 530 21805
rect 532 21799 548 21805
rect 525 21789 548 21798
rect 400 21779 404 21787
rect 498 21779 506 21789
rect 504 21755 506 21779
rect 514 21769 515 21789
rect 525 21764 528 21789
rect 547 21769 548 21789
rect 557 21779 564 21789
rect 514 21755 548 21759
rect 151 21708 156 21742
rect 174 21739 246 21747
rect 256 21739 328 21747
rect 336 21741 342 21749
rect 400 21744 404 21749
rect 180 21711 185 21739
rect 174 21703 246 21711
rect 256 21703 328 21711
rect 332 21709 336 21739
rect 400 21710 438 21744
rect 224 21673 226 21689
rect 196 21665 226 21673
rect 196 21661 232 21665
rect 196 21631 204 21661
rect 216 21631 232 21661
rect 224 21584 226 21631
rect 300 21604 308 21673
rect 332 21671 342 21709
rect 400 21701 404 21710
rect 454 21695 504 21697
rect 494 21691 548 21695
rect 494 21686 514 21691
rect 504 21671 506 21686
rect 336 21659 342 21671
rect 289 21594 308 21604
rect 300 21588 308 21594
rect 332 21625 342 21659
rect 400 21663 404 21671
rect 400 21629 408 21663
rect 434 21629 438 21663
rect 498 21661 506 21671
rect 514 21661 515 21681
rect 504 21645 506 21661
rect 525 21652 528 21686
rect 547 21661 548 21681
rect 557 21661 564 21671
rect 514 21645 530 21651
rect 532 21645 548 21651
rect 332 21597 373 21625
rect 332 21591 351 21597
rect 107 21537 119 21571
rect 129 21537 149 21571
rect 196 21550 204 21584
rect 216 21550 232 21584
rect 244 21578 257 21584
rect 278 21578 291 21588
rect 244 21554 291 21578
rect 300 21578 321 21588
rect 336 21581 351 21591
rect 300 21554 329 21578
rect 332 21563 351 21581
rect 361 21591 375 21597
rect 400 21591 411 21629
rect 562 21592 612 21594
rect 361 21563 381 21591
rect 400 21563 409 21591
rect 466 21583 497 21591
rect 565 21583 596 21591
rect 442 21576 500 21583
rect 466 21575 500 21576
rect 565 21575 599 21583
rect 244 21550 257 21554
rect 42 21471 46 21505
rect 72 21471 76 21505
rect 42 21424 76 21428
rect 42 21409 46 21424
rect 72 21409 76 21424
rect 38 21391 80 21409
rect 16 21385 102 21391
rect 144 21385 148 21537
rect 174 21513 181 21541
rect 224 21503 226 21550
rect 300 21541 308 21554
rect 278 21530 305 21541
rect 332 21513 342 21563
rect 400 21543 404 21563
rect 497 21559 500 21575
rect 596 21559 599 21575
rect 466 21558 500 21559
rect 442 21551 500 21558
rect 565 21551 599 21559
rect 612 21542 614 21592
rect 256 21503 328 21511
rect 336 21505 342 21513
rect 400 21505 404 21513
rect 196 21473 204 21503
rect 216 21473 232 21503
rect 196 21469 232 21473
rect 196 21461 226 21469
rect 224 21445 226 21461
rect 332 21433 336 21501
rect 400 21471 408 21505
rect 434 21471 438 21505
rect 454 21489 504 21491
rect 504 21473 506 21489
rect 514 21483 530 21489
rect 532 21483 548 21489
rect 525 21473 548 21482
rect 400 21463 404 21471
rect 498 21463 506 21473
rect 504 21439 506 21463
rect 514 21453 515 21473
rect 525 21448 528 21473
rect 547 21453 548 21473
rect 557 21463 564 21473
rect 514 21439 548 21443
rect 400 21433 442 21434
rect 174 21423 246 21431
rect 400 21426 404 21433
rect 295 21392 300 21426
rect 324 21392 329 21426
rect 367 21409 438 21426
rect 367 21392 442 21409
rect 400 21391 442 21392
rect 378 21385 464 21391
rect 38 21369 80 21385
rect 400 21369 442 21385
rect -25 21355 25 21357
rect 42 21355 76 21369
rect 404 21355 438 21369
rect 455 21355 505 21357
rect 557 21355 607 21357
rect 16 21347 102 21355
rect 378 21347 464 21355
rect 8 21313 17 21347
rect 18 21345 51 21347
rect 80 21345 100 21347
rect 18 21313 100 21345
rect 380 21345 404 21347
rect 429 21345 438 21347
rect 442 21345 462 21347
rect 16 21305 102 21313
rect 42 21289 76 21305
rect 16 21269 38 21275
rect 42 21266 76 21270
rect 80 21269 102 21275
rect 42 21236 46 21266
rect 72 21236 76 21266
rect 42 21155 46 21189
rect 72 21155 76 21189
rect -25 21118 25 21120
rect -8 21110 14 21117
rect -8 21109 17 21110
rect 25 21109 27 21118
rect -12 21102 38 21109
rect -12 21101 34 21102
rect -12 21097 8 21101
rect 0 21085 8 21097
rect 14 21085 34 21101
rect 0 21084 34 21085
rect 0 21077 38 21084
rect 14 21076 17 21077
rect 25 21068 27 21077
rect 42 21048 45 21138
rect 69 21123 80 21155
rect 107 21123 143 21151
rect 144 21123 148 21343
rect 332 21275 336 21343
rect 380 21313 462 21345
rect 463 21313 472 21347
rect 480 21313 497 21347
rect 378 21305 464 21313
rect 505 21305 507 21355
rect 514 21313 548 21347
rect 565 21313 582 21347
rect 607 21305 609 21355
rect 404 21289 438 21305
rect 400 21275 442 21276
rect 378 21269 404 21275
rect 442 21269 464 21275
rect 400 21268 404 21269
rect 174 21229 246 21237
rect 295 21234 300 21268
rect 324 21234 329 21268
rect 224 21199 226 21215
rect 196 21191 226 21199
rect 332 21197 336 21265
rect 367 21234 438 21268
rect 400 21227 404 21234
rect 454 21221 504 21223
rect 494 21217 548 21221
rect 494 21212 514 21217
rect 504 21197 506 21212
rect 196 21187 232 21191
rect 196 21157 204 21187
rect 216 21157 232 21187
rect 400 21189 404 21197
rect 107 21117 119 21123
rect 109 21089 119 21117
rect 129 21089 149 21123
rect 174 21119 181 21149
rect 224 21110 226 21157
rect 256 21149 328 21157
rect 332 21155 336 21185
rect 400 21155 408 21189
rect 434 21155 438 21189
rect 498 21187 506 21197
rect 514 21187 515 21207
rect 504 21171 506 21187
rect 525 21178 528 21212
rect 547 21187 548 21207
rect 557 21187 564 21197
rect 514 21171 530 21177
rect 532 21171 548 21177
rect 278 21119 305 21130
rect 42 20997 46 21031
rect 72 20997 76 21031
rect 38 20959 80 20960
rect 42 20918 76 20952
rect 79 20918 113 20952
rect 42 20839 46 20873
rect 72 20839 76 20873
rect -25 20802 25 20804
rect -8 20794 14 20801
rect -8 20793 17 20794
rect 25 20793 27 20802
rect -12 20786 38 20793
rect -12 20785 34 20786
rect -12 20781 8 20785
rect 0 20769 8 20781
rect 14 20769 34 20785
rect 0 20768 34 20769
rect 0 20761 38 20768
rect 14 20760 17 20761
rect 25 20752 27 20761
rect 42 20732 45 20822
rect 71 20791 80 20819
rect 69 20753 80 20791
rect 144 20781 148 21089
rect 196 21076 204 21110
rect 216 21076 232 21110
rect 244 21106 257 21110
rect 300 21106 308 21119
rect 332 21117 342 21155
rect 400 21147 404 21155
rect 336 21107 342 21117
rect 244 21082 291 21106
rect 244 21076 257 21082
rect 224 21029 226 21076
rect 278 21072 291 21082
rect 300 21082 329 21106
rect 332 21097 342 21107
rect 400 21107 409 21135
rect 562 21118 612 21120
rect 466 21109 497 21117
rect 565 21109 596 21117
rect 300 21072 321 21082
rect 300 21066 308 21072
rect 289 21056 308 21066
rect 196 20999 204 21029
rect 216 20999 232 21029
rect 196 20995 232 20999
rect 196 20987 226 20995
rect 300 20987 308 21056
rect 332 21063 351 21097
rect 361 21069 381 21097
rect 361 21063 375 21069
rect 400 21063 411 21107
rect 442 21102 500 21109
rect 466 21101 500 21102
rect 565 21101 599 21109
rect 497 21085 500 21101
rect 596 21085 599 21101
rect 466 21084 500 21085
rect 442 21077 500 21084
rect 565 21077 599 21085
rect 612 21068 614 21118
rect 332 21039 342 21063
rect 336 21027 342 21039
rect 224 20971 226 20987
rect 332 20959 342 21027
rect 400 21031 404 21039
rect 400 20997 408 21031
rect 434 20997 438 21031
rect 454 21015 504 21017
rect 504 20999 506 21015
rect 514 21009 530 21015
rect 532 21009 548 21015
rect 525 20999 548 21008
rect 400 20989 404 20997
rect 498 20989 506 20999
rect 504 20965 506 20989
rect 514 20979 515 20999
rect 525 20974 528 20999
rect 547 20979 548 20999
rect 557 20989 564 20999
rect 514 20965 548 20969
rect 151 20918 156 20952
rect 174 20949 246 20957
rect 256 20949 328 20957
rect 336 20951 342 20959
rect 400 20954 404 20959
rect 180 20921 185 20949
rect 174 20913 246 20921
rect 256 20913 328 20921
rect 332 20919 336 20949
rect 400 20920 438 20954
rect 224 20883 226 20899
rect 196 20875 226 20883
rect 196 20871 232 20875
rect 196 20841 204 20871
rect 216 20841 232 20871
rect 224 20794 226 20841
rect 300 20814 308 20883
rect 332 20881 342 20919
rect 400 20911 404 20920
rect 454 20905 504 20907
rect 494 20901 548 20905
rect 494 20896 514 20901
rect 504 20881 506 20896
rect 336 20869 342 20881
rect 289 20804 308 20814
rect 300 20798 308 20804
rect 332 20835 342 20869
rect 400 20873 404 20881
rect 400 20839 408 20873
rect 434 20839 438 20873
rect 498 20871 506 20881
rect 514 20871 515 20891
rect 504 20855 506 20871
rect 525 20862 528 20896
rect 547 20871 548 20891
rect 557 20871 564 20881
rect 514 20855 530 20861
rect 532 20855 548 20861
rect 332 20807 373 20835
rect 332 20801 351 20807
rect 107 20747 119 20781
rect 129 20747 149 20781
rect 196 20760 204 20794
rect 216 20760 232 20794
rect 244 20788 257 20794
rect 278 20788 291 20798
rect 244 20764 291 20788
rect 300 20788 321 20798
rect 336 20791 351 20801
rect 300 20764 329 20788
rect 332 20773 351 20791
rect 361 20801 375 20807
rect 400 20801 411 20839
rect 562 20802 612 20804
rect 361 20773 381 20801
rect 400 20773 409 20801
rect 466 20793 497 20801
rect 565 20793 596 20801
rect 442 20786 500 20793
rect 466 20785 500 20786
rect 565 20785 599 20793
rect 244 20760 257 20764
rect 42 20681 46 20715
rect 72 20681 76 20715
rect 42 20634 76 20638
rect 42 20619 46 20634
rect 72 20619 76 20634
rect 38 20601 80 20619
rect 16 20595 102 20601
rect 144 20595 148 20747
rect 174 20723 181 20751
rect 224 20713 226 20760
rect 300 20751 308 20764
rect 278 20740 305 20751
rect 332 20723 342 20773
rect 400 20753 404 20773
rect 497 20769 500 20785
rect 596 20769 599 20785
rect 466 20768 500 20769
rect 442 20761 500 20768
rect 565 20761 599 20769
rect 612 20752 614 20802
rect 256 20713 328 20721
rect 336 20715 342 20723
rect 400 20715 404 20723
rect 196 20683 204 20713
rect 216 20683 232 20713
rect 196 20679 232 20683
rect 196 20671 226 20679
rect 224 20655 226 20671
rect 332 20643 336 20711
rect 400 20681 408 20715
rect 434 20681 438 20715
rect 454 20699 504 20701
rect 504 20683 506 20699
rect 514 20693 530 20699
rect 532 20693 548 20699
rect 525 20683 548 20692
rect 400 20673 404 20681
rect 498 20673 506 20683
rect 504 20649 506 20673
rect 514 20663 515 20683
rect 525 20658 528 20683
rect 547 20663 548 20683
rect 557 20673 564 20683
rect 514 20649 548 20653
rect 400 20643 442 20644
rect 174 20633 246 20641
rect 400 20636 404 20643
rect 295 20602 300 20636
rect 324 20602 329 20636
rect 367 20619 438 20636
rect 367 20602 442 20619
rect 400 20601 442 20602
rect 378 20595 464 20601
rect 38 20579 80 20595
rect 400 20579 442 20595
rect -25 20565 25 20567
rect 42 20565 76 20579
rect 404 20565 438 20579
rect 455 20565 505 20567
rect 557 20565 607 20567
rect 16 20557 102 20565
rect 378 20557 464 20565
rect 8 20523 17 20557
rect 18 20555 51 20557
rect 80 20555 100 20557
rect 18 20523 100 20555
rect 380 20555 404 20557
rect 429 20555 438 20557
rect 442 20555 462 20557
rect 16 20515 102 20523
rect 42 20499 76 20515
rect 16 20479 38 20485
rect 42 20476 76 20480
rect 80 20479 102 20485
rect 42 20446 46 20476
rect 72 20446 76 20476
rect 42 20365 46 20399
rect 72 20365 76 20399
rect -25 20328 25 20330
rect -8 20320 14 20327
rect -8 20319 17 20320
rect 25 20319 27 20328
rect -12 20312 38 20319
rect -12 20311 34 20312
rect -12 20307 8 20311
rect 0 20295 8 20307
rect 14 20295 34 20311
rect 0 20294 34 20295
rect 0 20287 38 20294
rect 14 20286 17 20287
rect 25 20278 27 20287
rect 42 20258 45 20348
rect 69 20333 80 20365
rect 107 20333 143 20361
rect 144 20333 148 20553
rect 332 20485 336 20553
rect 380 20523 462 20555
rect 463 20523 472 20557
rect 480 20523 497 20557
rect 378 20515 464 20523
rect 505 20515 507 20565
rect 514 20523 548 20557
rect 565 20523 582 20557
rect 607 20515 609 20565
rect 404 20499 438 20515
rect 400 20485 442 20486
rect 378 20479 404 20485
rect 442 20479 464 20485
rect 400 20478 404 20479
rect 174 20439 246 20447
rect 295 20444 300 20478
rect 324 20444 329 20478
rect 224 20409 226 20425
rect 196 20401 226 20409
rect 332 20407 336 20475
rect 367 20444 438 20478
rect 400 20437 404 20444
rect 454 20431 504 20433
rect 494 20427 548 20431
rect 494 20422 514 20427
rect 504 20407 506 20422
rect 196 20397 232 20401
rect 196 20367 204 20397
rect 216 20367 232 20397
rect 400 20399 404 20407
rect 107 20327 119 20333
rect 109 20299 119 20327
rect 129 20299 149 20333
rect 174 20329 181 20359
rect 224 20320 226 20367
rect 256 20359 328 20367
rect 332 20365 336 20395
rect 400 20365 408 20399
rect 434 20365 438 20399
rect 498 20397 506 20407
rect 514 20397 515 20417
rect 504 20381 506 20397
rect 525 20388 528 20422
rect 547 20397 548 20417
rect 557 20397 564 20407
rect 514 20381 530 20387
rect 532 20381 548 20387
rect 278 20329 305 20340
rect 42 20207 46 20241
rect 72 20207 76 20241
rect 38 20169 80 20170
rect 42 20128 76 20162
rect 79 20128 113 20162
rect 42 20049 46 20083
rect 72 20049 76 20083
rect -25 20012 25 20014
rect -8 20004 14 20011
rect -8 20003 17 20004
rect 25 20003 27 20012
rect -12 19996 38 20003
rect -12 19995 34 19996
rect -12 19991 8 19995
rect 0 19979 8 19991
rect 14 19979 34 19995
rect 0 19978 34 19979
rect 0 19971 38 19978
rect 14 19970 17 19971
rect 25 19962 27 19971
rect 42 19942 45 20032
rect 71 20001 80 20029
rect 69 19963 80 20001
rect 144 19991 148 20299
rect 196 20286 204 20320
rect 216 20286 232 20320
rect 244 20316 257 20320
rect 300 20316 308 20329
rect 332 20327 342 20365
rect 400 20357 404 20365
rect 336 20317 342 20327
rect 244 20292 291 20316
rect 244 20286 257 20292
rect 224 20239 226 20286
rect 278 20282 291 20292
rect 300 20292 329 20316
rect 332 20307 342 20317
rect 400 20317 409 20345
rect 562 20328 612 20330
rect 466 20319 497 20327
rect 565 20319 596 20327
rect 300 20282 321 20292
rect 300 20276 308 20282
rect 289 20266 308 20276
rect 196 20209 204 20239
rect 216 20209 232 20239
rect 196 20205 232 20209
rect 196 20197 226 20205
rect 300 20197 308 20266
rect 332 20273 351 20307
rect 361 20279 381 20307
rect 361 20273 375 20279
rect 400 20273 411 20317
rect 442 20312 500 20319
rect 466 20311 500 20312
rect 565 20311 599 20319
rect 497 20295 500 20311
rect 596 20295 599 20311
rect 466 20294 500 20295
rect 442 20287 500 20294
rect 565 20287 599 20295
rect 612 20278 614 20328
rect 332 20249 342 20273
rect 336 20237 342 20249
rect 224 20181 226 20197
rect 332 20169 342 20237
rect 400 20241 404 20249
rect 400 20207 408 20241
rect 434 20207 438 20241
rect 454 20225 504 20227
rect 504 20209 506 20225
rect 514 20219 530 20225
rect 532 20219 548 20225
rect 525 20209 548 20218
rect 400 20199 404 20207
rect 498 20199 506 20209
rect 504 20175 506 20199
rect 514 20189 515 20209
rect 525 20184 528 20209
rect 547 20189 548 20209
rect 557 20199 564 20209
rect 514 20175 548 20179
rect 151 20128 156 20162
rect 174 20159 246 20167
rect 256 20159 328 20167
rect 336 20161 342 20169
rect 400 20164 404 20169
rect 180 20131 185 20159
rect 174 20123 246 20131
rect 256 20123 328 20131
rect 332 20129 336 20159
rect 400 20130 438 20164
rect 224 20093 226 20109
rect 196 20085 226 20093
rect 196 20081 232 20085
rect 196 20051 204 20081
rect 216 20051 232 20081
rect 224 20004 226 20051
rect 300 20024 308 20093
rect 332 20091 342 20129
rect 400 20121 404 20130
rect 454 20115 504 20117
rect 494 20111 548 20115
rect 494 20106 514 20111
rect 504 20091 506 20106
rect 336 20079 342 20091
rect 289 20014 308 20024
rect 300 20008 308 20014
rect 332 20045 342 20079
rect 400 20083 404 20091
rect 400 20049 408 20083
rect 434 20049 438 20083
rect 498 20081 506 20091
rect 514 20081 515 20101
rect 504 20065 506 20081
rect 525 20072 528 20106
rect 547 20081 548 20101
rect 557 20081 564 20091
rect 514 20065 530 20071
rect 532 20065 548 20071
rect 332 20017 373 20045
rect 332 20011 351 20017
rect 107 19957 119 19991
rect 129 19957 149 19991
rect 196 19970 204 20004
rect 216 19970 232 20004
rect 244 19998 257 20004
rect 278 19998 291 20008
rect 244 19974 291 19998
rect 300 19998 321 20008
rect 336 20001 351 20011
rect 300 19974 329 19998
rect 332 19983 351 20001
rect 361 20011 375 20017
rect 400 20011 411 20049
rect 562 20012 612 20014
rect 361 19983 381 20011
rect 400 19983 409 20011
rect 466 20003 497 20011
rect 565 20003 596 20011
rect 442 19996 500 20003
rect 466 19995 500 19996
rect 565 19995 599 20003
rect 244 19970 257 19974
rect 42 19891 46 19925
rect 72 19891 76 19925
rect 42 19844 76 19848
rect 42 19829 46 19844
rect 72 19829 76 19844
rect 38 19811 80 19829
rect 16 19805 102 19811
rect 144 19805 148 19957
rect 174 19933 181 19961
rect 224 19923 226 19970
rect 300 19961 308 19974
rect 278 19950 305 19961
rect 332 19933 342 19983
rect 400 19963 404 19983
rect 497 19979 500 19995
rect 596 19979 599 19995
rect 466 19978 500 19979
rect 442 19971 500 19978
rect 565 19971 599 19979
rect 612 19962 614 20012
rect 256 19923 328 19931
rect 336 19925 342 19933
rect 400 19925 404 19933
rect 196 19893 204 19923
rect 216 19893 232 19923
rect 196 19889 232 19893
rect 196 19881 226 19889
rect 224 19865 226 19881
rect 332 19853 336 19921
rect 400 19891 408 19925
rect 434 19891 438 19925
rect 454 19909 504 19911
rect 504 19893 506 19909
rect 514 19903 530 19909
rect 532 19903 548 19909
rect 525 19893 548 19902
rect 400 19883 404 19891
rect 498 19883 506 19893
rect 504 19859 506 19883
rect 514 19873 515 19893
rect 525 19868 528 19893
rect 547 19873 548 19893
rect 557 19883 564 19893
rect 514 19859 548 19863
rect 400 19853 442 19854
rect 174 19843 246 19851
rect 400 19846 404 19853
rect 295 19812 300 19846
rect 324 19812 329 19846
rect 367 19829 438 19846
rect 367 19812 442 19829
rect 400 19811 442 19812
rect 378 19805 464 19811
rect 38 19789 80 19805
rect 400 19789 442 19805
rect -25 19775 25 19777
rect 42 19775 76 19789
rect 404 19775 438 19789
rect 455 19775 505 19777
rect 557 19775 607 19777
rect 16 19767 102 19775
rect 378 19767 464 19775
rect 8 19733 17 19767
rect 18 19765 51 19767
rect 80 19765 100 19767
rect 18 19733 100 19765
rect 380 19765 404 19767
rect 429 19765 438 19767
rect 442 19765 462 19767
rect 16 19725 102 19733
rect 42 19709 76 19725
rect 16 19689 38 19695
rect 42 19686 76 19690
rect 80 19689 102 19695
rect 42 19656 46 19686
rect 72 19656 76 19686
rect 42 19575 46 19609
rect 72 19575 76 19609
rect -25 19538 25 19540
rect -8 19530 14 19537
rect -8 19529 17 19530
rect 25 19529 27 19538
rect -12 19522 38 19529
rect -12 19521 34 19522
rect -12 19517 8 19521
rect 0 19505 8 19517
rect 14 19505 34 19521
rect 0 19504 34 19505
rect 0 19497 38 19504
rect 14 19496 17 19497
rect 25 19488 27 19497
rect 42 19468 45 19558
rect 69 19543 80 19575
rect 107 19543 143 19571
rect 144 19543 148 19763
rect 332 19695 336 19763
rect 380 19733 462 19765
rect 463 19733 472 19767
rect 480 19733 497 19767
rect 378 19725 464 19733
rect 505 19725 507 19775
rect 514 19733 548 19767
rect 565 19733 582 19767
rect 607 19725 609 19775
rect 404 19709 438 19725
rect 400 19695 442 19696
rect 378 19689 404 19695
rect 442 19689 464 19695
rect 400 19688 404 19689
rect 174 19649 246 19657
rect 295 19654 300 19688
rect 324 19654 329 19688
rect 224 19619 226 19635
rect 196 19611 226 19619
rect 332 19617 336 19685
rect 367 19654 438 19688
rect 400 19647 404 19654
rect 454 19641 504 19643
rect 494 19637 548 19641
rect 494 19632 514 19637
rect 504 19617 506 19632
rect 196 19607 232 19611
rect 196 19577 204 19607
rect 216 19577 232 19607
rect 400 19609 404 19617
rect 107 19537 119 19543
rect 109 19509 119 19537
rect 129 19509 149 19543
rect 174 19539 181 19569
rect 224 19530 226 19577
rect 256 19569 328 19577
rect 332 19575 336 19605
rect 400 19575 408 19609
rect 434 19575 438 19609
rect 498 19607 506 19617
rect 514 19607 515 19627
rect 504 19591 506 19607
rect 525 19598 528 19632
rect 547 19607 548 19627
rect 557 19607 564 19617
rect 514 19591 530 19597
rect 532 19591 548 19597
rect 278 19539 305 19550
rect 42 19417 46 19451
rect 72 19417 76 19451
rect 38 19379 80 19380
rect 42 19338 76 19372
rect 79 19338 113 19372
rect 42 19259 46 19293
rect 72 19259 76 19293
rect -25 19222 25 19224
rect -8 19214 14 19221
rect -8 19213 17 19214
rect 25 19213 27 19222
rect -12 19206 38 19213
rect -12 19205 34 19206
rect -12 19201 8 19205
rect 0 19189 8 19201
rect 14 19189 34 19205
rect 0 19188 34 19189
rect 0 19181 38 19188
rect 14 19180 17 19181
rect 25 19172 27 19181
rect 42 19152 45 19242
rect 71 19211 80 19239
rect 69 19173 80 19211
rect 144 19201 148 19509
rect 196 19496 204 19530
rect 216 19496 232 19530
rect 244 19526 257 19530
rect 300 19526 308 19539
rect 332 19537 342 19575
rect 400 19567 404 19575
rect 336 19527 342 19537
rect 244 19502 291 19526
rect 244 19496 257 19502
rect 224 19449 226 19496
rect 278 19492 291 19502
rect 300 19502 329 19526
rect 332 19517 342 19527
rect 400 19527 409 19555
rect 562 19538 612 19540
rect 466 19529 497 19537
rect 565 19529 596 19537
rect 300 19492 321 19502
rect 300 19486 308 19492
rect 289 19476 308 19486
rect 196 19419 204 19449
rect 216 19419 232 19449
rect 196 19415 232 19419
rect 196 19407 226 19415
rect 300 19407 308 19476
rect 332 19483 351 19517
rect 361 19489 381 19517
rect 361 19483 375 19489
rect 400 19483 411 19527
rect 442 19522 500 19529
rect 466 19521 500 19522
rect 565 19521 599 19529
rect 497 19505 500 19521
rect 596 19505 599 19521
rect 466 19504 500 19505
rect 442 19497 500 19504
rect 565 19497 599 19505
rect 612 19488 614 19538
rect 332 19459 342 19483
rect 336 19447 342 19459
rect 224 19391 226 19407
rect 332 19379 342 19447
rect 400 19451 404 19459
rect 400 19417 408 19451
rect 434 19417 438 19451
rect 454 19435 504 19437
rect 504 19419 506 19435
rect 514 19429 530 19435
rect 532 19429 548 19435
rect 525 19419 548 19428
rect 400 19409 404 19417
rect 498 19409 506 19419
rect 504 19385 506 19409
rect 514 19399 515 19419
rect 525 19394 528 19419
rect 547 19399 548 19419
rect 557 19409 564 19419
rect 514 19385 548 19389
rect 151 19338 156 19372
rect 174 19369 246 19377
rect 256 19369 328 19377
rect 336 19371 342 19379
rect 400 19374 404 19379
rect 180 19341 185 19369
rect 174 19333 246 19341
rect 256 19333 328 19341
rect 332 19339 336 19369
rect 400 19340 438 19374
rect 224 19303 226 19319
rect 196 19295 226 19303
rect 196 19291 232 19295
rect 196 19261 204 19291
rect 216 19261 232 19291
rect 224 19214 226 19261
rect 300 19234 308 19303
rect 332 19301 342 19339
rect 400 19331 404 19340
rect 454 19325 504 19327
rect 494 19321 548 19325
rect 494 19316 514 19321
rect 504 19301 506 19316
rect 336 19289 342 19301
rect 289 19224 308 19234
rect 300 19218 308 19224
rect 332 19255 342 19289
rect 400 19293 404 19301
rect 400 19259 408 19293
rect 434 19259 438 19293
rect 498 19291 506 19301
rect 514 19291 515 19311
rect 504 19275 506 19291
rect 525 19282 528 19316
rect 547 19291 548 19311
rect 557 19291 564 19301
rect 514 19275 530 19281
rect 532 19275 548 19281
rect 332 19227 373 19255
rect 332 19221 351 19227
rect 107 19167 119 19201
rect 129 19167 149 19201
rect 196 19180 204 19214
rect 216 19180 232 19214
rect 244 19208 257 19214
rect 278 19208 291 19218
rect 244 19184 291 19208
rect 300 19208 321 19218
rect 336 19211 351 19221
rect 300 19184 329 19208
rect 332 19193 351 19211
rect 361 19221 375 19227
rect 400 19221 411 19259
rect 562 19222 612 19224
rect 361 19193 381 19221
rect 400 19193 409 19221
rect 466 19213 497 19221
rect 565 19213 596 19221
rect 442 19206 500 19213
rect 466 19205 500 19206
rect 565 19205 599 19213
rect 244 19180 257 19184
rect 42 19101 46 19135
rect 72 19101 76 19135
rect 42 19054 76 19058
rect 42 19039 46 19054
rect 72 19039 76 19054
rect 38 19021 80 19039
rect 16 19015 102 19021
rect 144 19015 148 19167
rect 174 19143 181 19171
rect 224 19133 226 19180
rect 300 19171 308 19184
rect 278 19160 305 19171
rect 332 19143 342 19193
rect 400 19173 404 19193
rect 497 19189 500 19205
rect 596 19189 599 19205
rect 466 19188 500 19189
rect 442 19181 500 19188
rect 565 19181 599 19189
rect 612 19172 614 19222
rect 256 19133 328 19141
rect 336 19135 342 19143
rect 400 19135 404 19143
rect 196 19103 204 19133
rect 216 19103 232 19133
rect 196 19099 232 19103
rect 196 19091 226 19099
rect 224 19075 226 19091
rect 332 19063 336 19131
rect 400 19101 408 19135
rect 434 19101 438 19135
rect 454 19119 504 19121
rect 504 19103 506 19119
rect 514 19113 530 19119
rect 532 19113 548 19119
rect 525 19103 548 19112
rect 400 19093 404 19101
rect 498 19093 506 19103
rect 504 19069 506 19093
rect 514 19083 515 19103
rect 525 19078 528 19103
rect 547 19083 548 19103
rect 557 19093 564 19103
rect 514 19069 548 19073
rect 400 19063 442 19064
rect 174 19053 246 19061
rect 400 19056 404 19063
rect 295 19022 300 19056
rect 324 19022 329 19056
rect 367 19039 438 19056
rect 367 19022 442 19039
rect 400 19021 442 19022
rect 378 19015 464 19021
rect 38 18999 80 19015
rect 400 18999 442 19015
rect -25 18985 25 18987
rect 42 18985 76 18999
rect 404 18985 438 18999
rect 455 18985 505 18987
rect 557 18985 607 18987
rect 16 18977 102 18985
rect 378 18977 464 18985
rect 8 18943 17 18977
rect 18 18975 51 18977
rect 80 18975 100 18977
rect 18 18943 100 18975
rect 380 18975 404 18977
rect 429 18975 438 18977
rect 442 18975 462 18977
rect 16 18935 102 18943
rect 42 18919 76 18935
rect 16 18899 38 18905
rect 42 18896 76 18900
rect 80 18899 102 18905
rect 42 18866 46 18896
rect 72 18866 76 18896
rect 42 18785 46 18819
rect 72 18785 76 18819
rect -25 18748 25 18750
rect -8 18740 14 18747
rect -8 18739 17 18740
rect 25 18739 27 18748
rect -12 18732 38 18739
rect -12 18731 34 18732
rect -12 18727 8 18731
rect 0 18715 8 18727
rect 14 18715 34 18731
rect 0 18714 34 18715
rect 0 18707 38 18714
rect 14 18706 17 18707
rect 25 18698 27 18707
rect 42 18678 45 18768
rect 69 18753 80 18785
rect 107 18753 143 18781
rect 144 18753 148 18973
rect 332 18905 336 18973
rect 380 18943 462 18975
rect 463 18943 472 18977
rect 480 18943 497 18977
rect 378 18935 464 18943
rect 505 18935 507 18985
rect 514 18943 548 18977
rect 565 18943 582 18977
rect 607 18935 609 18985
rect 404 18919 438 18935
rect 400 18905 442 18906
rect 378 18899 404 18905
rect 442 18899 464 18905
rect 400 18898 404 18899
rect 174 18859 246 18867
rect 295 18864 300 18898
rect 324 18864 329 18898
rect 224 18829 226 18845
rect 196 18821 226 18829
rect 332 18827 336 18895
rect 367 18864 438 18898
rect 400 18857 404 18864
rect 454 18851 504 18853
rect 494 18847 548 18851
rect 494 18842 514 18847
rect 504 18827 506 18842
rect 196 18817 232 18821
rect 196 18787 204 18817
rect 216 18787 232 18817
rect 400 18819 404 18827
rect 107 18747 119 18753
rect 109 18719 119 18747
rect 129 18719 149 18753
rect 174 18749 181 18779
rect 224 18740 226 18787
rect 256 18779 328 18787
rect 332 18785 336 18815
rect 400 18785 408 18819
rect 434 18785 438 18819
rect 498 18817 506 18827
rect 514 18817 515 18837
rect 504 18801 506 18817
rect 525 18808 528 18842
rect 547 18817 548 18837
rect 557 18817 564 18827
rect 514 18801 530 18807
rect 532 18801 548 18807
rect 278 18749 305 18760
rect 42 18627 46 18661
rect 72 18627 76 18661
rect 38 18589 80 18590
rect 42 18548 76 18582
rect 79 18548 113 18582
rect 42 18469 46 18503
rect 72 18469 76 18503
rect -25 18432 25 18434
rect -8 18424 14 18431
rect -8 18423 17 18424
rect 25 18423 27 18432
rect -12 18416 38 18423
rect -12 18415 34 18416
rect -12 18411 8 18415
rect 0 18399 8 18411
rect 14 18399 34 18415
rect 0 18398 34 18399
rect 0 18391 38 18398
rect 14 18390 17 18391
rect 25 18382 27 18391
rect 42 18362 45 18452
rect 71 18421 80 18449
rect 69 18383 80 18421
rect 144 18411 148 18719
rect 196 18706 204 18740
rect 216 18706 232 18740
rect 244 18736 257 18740
rect 300 18736 308 18749
rect 332 18747 342 18785
rect 400 18777 404 18785
rect 336 18737 342 18747
rect 244 18712 291 18736
rect 244 18706 257 18712
rect 224 18659 226 18706
rect 278 18702 291 18712
rect 300 18712 329 18736
rect 332 18727 342 18737
rect 400 18737 409 18765
rect 562 18748 612 18750
rect 466 18739 497 18747
rect 565 18739 596 18747
rect 300 18702 321 18712
rect 300 18696 308 18702
rect 289 18686 308 18696
rect 196 18629 204 18659
rect 216 18629 232 18659
rect 196 18625 232 18629
rect 196 18617 226 18625
rect 300 18617 308 18686
rect 332 18693 351 18727
rect 361 18699 381 18727
rect 361 18693 375 18699
rect 400 18693 411 18737
rect 442 18732 500 18739
rect 466 18731 500 18732
rect 565 18731 599 18739
rect 497 18715 500 18731
rect 596 18715 599 18731
rect 466 18714 500 18715
rect 442 18707 500 18714
rect 565 18707 599 18715
rect 612 18698 614 18748
rect 332 18669 342 18693
rect 336 18657 342 18669
rect 224 18601 226 18617
rect 332 18589 342 18657
rect 400 18661 404 18669
rect 400 18627 408 18661
rect 434 18627 438 18661
rect 454 18645 504 18647
rect 504 18629 506 18645
rect 514 18639 530 18645
rect 532 18639 548 18645
rect 525 18629 548 18638
rect 400 18619 404 18627
rect 498 18619 506 18629
rect 504 18595 506 18619
rect 514 18609 515 18629
rect 525 18604 528 18629
rect 547 18609 548 18629
rect 557 18619 564 18629
rect 514 18595 548 18599
rect 151 18548 156 18582
rect 174 18579 246 18587
rect 256 18579 328 18587
rect 336 18581 342 18589
rect 400 18584 404 18589
rect 180 18551 185 18579
rect 174 18543 246 18551
rect 256 18543 328 18551
rect 332 18549 336 18579
rect 400 18550 438 18584
rect 224 18513 226 18529
rect 196 18505 226 18513
rect 196 18501 232 18505
rect 196 18471 204 18501
rect 216 18471 232 18501
rect 224 18424 226 18471
rect 300 18444 308 18513
rect 332 18511 342 18549
rect 400 18541 404 18550
rect 454 18535 504 18537
rect 494 18531 548 18535
rect 494 18526 514 18531
rect 504 18511 506 18526
rect 336 18499 342 18511
rect 289 18434 308 18444
rect 300 18428 308 18434
rect 332 18465 342 18499
rect 400 18503 404 18511
rect 400 18469 408 18503
rect 434 18469 438 18503
rect 498 18501 506 18511
rect 514 18501 515 18521
rect 504 18485 506 18501
rect 525 18492 528 18526
rect 547 18501 548 18521
rect 557 18501 564 18511
rect 514 18485 530 18491
rect 532 18485 548 18491
rect 332 18437 373 18465
rect 332 18431 351 18437
rect 107 18377 119 18411
rect 129 18377 149 18411
rect 196 18390 204 18424
rect 216 18390 232 18424
rect 244 18418 257 18424
rect 278 18418 291 18428
rect 244 18394 291 18418
rect 300 18418 321 18428
rect 336 18421 351 18431
rect 300 18394 329 18418
rect 332 18403 351 18421
rect 361 18431 375 18437
rect 400 18431 411 18469
rect 562 18432 612 18434
rect 361 18403 381 18431
rect 400 18403 409 18431
rect 466 18423 497 18431
rect 565 18423 596 18431
rect 442 18416 500 18423
rect 466 18415 500 18416
rect 565 18415 599 18423
rect 244 18390 257 18394
rect 42 18311 46 18345
rect 72 18311 76 18345
rect 42 18264 76 18268
rect 42 18249 46 18264
rect 72 18249 76 18264
rect 38 18231 80 18249
rect 16 18225 102 18231
rect 144 18225 148 18377
rect 174 18353 181 18381
rect 224 18343 226 18390
rect 300 18381 308 18394
rect 278 18370 305 18381
rect 332 18353 342 18403
rect 400 18383 404 18403
rect 497 18399 500 18415
rect 596 18399 599 18415
rect 466 18398 500 18399
rect 442 18391 500 18398
rect 565 18391 599 18399
rect 612 18382 614 18432
rect 256 18343 328 18351
rect 336 18345 342 18353
rect 400 18345 404 18353
rect 196 18313 204 18343
rect 216 18313 232 18343
rect 196 18309 232 18313
rect 196 18301 226 18309
rect 224 18285 226 18301
rect 332 18273 336 18341
rect 400 18311 408 18345
rect 434 18311 438 18345
rect 454 18329 504 18331
rect 504 18313 506 18329
rect 514 18323 530 18329
rect 532 18323 548 18329
rect 525 18313 548 18322
rect 400 18303 404 18311
rect 498 18303 506 18313
rect 504 18279 506 18303
rect 514 18293 515 18313
rect 525 18288 528 18313
rect 547 18293 548 18313
rect 557 18303 564 18313
rect 514 18279 548 18283
rect 400 18273 442 18274
rect 174 18263 246 18271
rect 400 18266 404 18273
rect 295 18232 300 18266
rect 324 18232 329 18266
rect 367 18249 438 18266
rect 367 18232 442 18249
rect 400 18231 442 18232
rect 378 18225 464 18231
rect 38 18209 80 18225
rect 400 18209 442 18225
rect -25 18195 25 18197
rect 42 18195 76 18209
rect 404 18195 438 18209
rect 455 18195 505 18197
rect 557 18195 607 18197
rect 16 18187 102 18195
rect 378 18187 464 18195
rect 8 18153 17 18187
rect 18 18185 51 18187
rect 80 18185 100 18187
rect 18 18153 100 18185
rect 380 18185 404 18187
rect 429 18185 438 18187
rect 442 18185 462 18187
rect 16 18145 102 18153
rect 42 18129 76 18145
rect 16 18109 38 18115
rect 42 18106 76 18110
rect 80 18109 102 18115
rect 42 18076 46 18106
rect 72 18076 76 18106
rect 42 17995 46 18029
rect 72 17995 76 18029
rect -25 17958 25 17960
rect -8 17950 14 17957
rect -8 17949 17 17950
rect 25 17949 27 17958
rect -12 17942 38 17949
rect -12 17941 34 17942
rect -12 17937 8 17941
rect 0 17925 8 17937
rect 14 17925 34 17941
rect 0 17924 34 17925
rect 0 17917 38 17924
rect 14 17916 17 17917
rect 25 17908 27 17917
rect 42 17888 45 17978
rect 69 17963 80 17995
rect 107 17963 143 17991
rect 144 17963 148 18183
rect 332 18115 336 18183
rect 380 18153 462 18185
rect 463 18153 472 18187
rect 480 18153 497 18187
rect 378 18145 464 18153
rect 505 18145 507 18195
rect 514 18153 548 18187
rect 565 18153 582 18187
rect 607 18145 609 18195
rect 404 18129 438 18145
rect 400 18115 442 18116
rect 378 18109 404 18115
rect 442 18109 464 18115
rect 400 18108 404 18109
rect 174 18069 246 18077
rect 295 18074 300 18108
rect 324 18074 329 18108
rect 224 18039 226 18055
rect 196 18031 226 18039
rect 332 18037 336 18105
rect 367 18074 438 18108
rect 400 18067 404 18074
rect 454 18061 504 18063
rect 494 18057 548 18061
rect 494 18052 514 18057
rect 504 18037 506 18052
rect 196 18027 232 18031
rect 196 17997 204 18027
rect 216 17997 232 18027
rect 400 18029 404 18037
rect 107 17957 119 17963
rect 109 17929 119 17957
rect 129 17929 149 17963
rect 174 17959 181 17989
rect 224 17950 226 17997
rect 256 17989 328 17997
rect 332 17995 336 18025
rect 400 17995 408 18029
rect 434 17995 438 18029
rect 498 18027 506 18037
rect 514 18027 515 18047
rect 504 18011 506 18027
rect 525 18018 528 18052
rect 547 18027 548 18047
rect 557 18027 564 18037
rect 514 18011 530 18017
rect 532 18011 548 18017
rect 278 17959 305 17970
rect 42 17837 46 17871
rect 72 17837 76 17871
rect 38 17799 80 17800
rect 42 17758 76 17792
rect 79 17758 113 17792
rect 42 17679 46 17713
rect 72 17679 76 17713
rect -25 17642 25 17644
rect -8 17634 14 17641
rect -8 17633 17 17634
rect 25 17633 27 17642
rect -12 17626 38 17633
rect -12 17625 34 17626
rect -12 17621 8 17625
rect 0 17609 8 17621
rect 14 17609 34 17625
rect 0 17608 34 17609
rect 0 17601 38 17608
rect 14 17600 17 17601
rect 25 17592 27 17601
rect 42 17572 45 17662
rect 71 17631 80 17659
rect 69 17593 80 17631
rect 144 17621 148 17929
rect 196 17916 204 17950
rect 216 17916 232 17950
rect 244 17946 257 17950
rect 300 17946 308 17959
rect 332 17957 342 17995
rect 400 17987 404 17995
rect 336 17947 342 17957
rect 244 17922 291 17946
rect 244 17916 257 17922
rect 224 17869 226 17916
rect 278 17912 291 17922
rect 300 17922 329 17946
rect 332 17937 342 17947
rect 400 17947 409 17975
rect 562 17958 612 17960
rect 466 17949 497 17957
rect 565 17949 596 17957
rect 300 17912 321 17922
rect 300 17906 308 17912
rect 289 17896 308 17906
rect 196 17839 204 17869
rect 216 17839 232 17869
rect 196 17835 232 17839
rect 196 17827 226 17835
rect 300 17827 308 17896
rect 332 17903 351 17937
rect 361 17909 381 17937
rect 361 17903 375 17909
rect 400 17903 411 17947
rect 442 17942 500 17949
rect 466 17941 500 17942
rect 565 17941 599 17949
rect 497 17925 500 17941
rect 596 17925 599 17941
rect 466 17924 500 17925
rect 442 17917 500 17924
rect 565 17917 599 17925
rect 612 17908 614 17958
rect 332 17879 342 17903
rect 336 17867 342 17879
rect 224 17811 226 17827
rect 332 17799 342 17867
rect 400 17871 404 17879
rect 400 17837 408 17871
rect 434 17837 438 17871
rect 454 17855 504 17857
rect 504 17839 506 17855
rect 514 17849 530 17855
rect 532 17849 548 17855
rect 525 17839 548 17848
rect 400 17829 404 17837
rect 498 17829 506 17839
rect 504 17805 506 17829
rect 514 17819 515 17839
rect 525 17814 528 17839
rect 547 17819 548 17839
rect 557 17829 564 17839
rect 514 17805 548 17809
rect 151 17758 156 17792
rect 174 17789 246 17797
rect 256 17789 328 17797
rect 336 17791 342 17799
rect 400 17794 404 17799
rect 180 17761 185 17789
rect 174 17753 246 17761
rect 256 17753 328 17761
rect 332 17759 336 17789
rect 400 17760 438 17794
rect 224 17723 226 17739
rect 196 17715 226 17723
rect 196 17711 232 17715
rect 196 17681 204 17711
rect 216 17681 232 17711
rect 224 17634 226 17681
rect 300 17654 308 17723
rect 332 17721 342 17759
rect 400 17751 404 17760
rect 454 17745 504 17747
rect 494 17741 548 17745
rect 494 17736 514 17741
rect 504 17721 506 17736
rect 336 17709 342 17721
rect 289 17644 308 17654
rect 300 17638 308 17644
rect 332 17675 342 17709
rect 400 17713 404 17721
rect 400 17679 408 17713
rect 434 17679 438 17713
rect 498 17711 506 17721
rect 514 17711 515 17731
rect 504 17695 506 17711
rect 525 17702 528 17736
rect 547 17711 548 17731
rect 557 17711 564 17721
rect 514 17695 530 17701
rect 532 17695 548 17701
rect 332 17647 373 17675
rect 332 17641 351 17647
rect 107 17587 119 17621
rect 129 17587 149 17621
rect 196 17600 204 17634
rect 216 17600 232 17634
rect 244 17628 257 17634
rect 278 17628 291 17638
rect 244 17604 291 17628
rect 300 17628 321 17638
rect 336 17631 351 17641
rect 300 17604 329 17628
rect 332 17613 351 17631
rect 361 17641 375 17647
rect 400 17641 411 17679
rect 562 17642 612 17644
rect 361 17613 381 17641
rect 400 17613 409 17641
rect 466 17633 497 17641
rect 565 17633 596 17641
rect 442 17626 500 17633
rect 466 17625 500 17626
rect 565 17625 599 17633
rect 244 17600 257 17604
rect 42 17521 46 17555
rect 72 17521 76 17555
rect 42 17474 76 17478
rect 42 17459 46 17474
rect 72 17459 76 17474
rect 38 17441 80 17459
rect 16 17435 102 17441
rect 144 17435 148 17587
rect 174 17563 181 17591
rect 224 17553 226 17600
rect 300 17591 308 17604
rect 278 17580 305 17591
rect 332 17563 342 17613
rect 400 17593 404 17613
rect 497 17609 500 17625
rect 596 17609 599 17625
rect 466 17608 500 17609
rect 442 17601 500 17608
rect 565 17601 599 17609
rect 612 17592 614 17642
rect 256 17553 328 17561
rect 336 17555 342 17563
rect 400 17555 404 17563
rect 196 17523 204 17553
rect 216 17523 232 17553
rect 196 17519 232 17523
rect 196 17511 226 17519
rect 224 17495 226 17511
rect 332 17483 336 17551
rect 400 17521 408 17555
rect 434 17521 438 17555
rect 454 17539 504 17541
rect 504 17523 506 17539
rect 514 17533 530 17539
rect 532 17533 548 17539
rect 525 17523 548 17532
rect 400 17513 404 17521
rect 498 17513 506 17523
rect 504 17489 506 17513
rect 514 17503 515 17523
rect 525 17498 528 17523
rect 547 17503 548 17523
rect 557 17513 564 17523
rect 514 17489 548 17493
rect 400 17483 442 17484
rect 174 17473 246 17481
rect 400 17476 404 17483
rect 295 17442 300 17476
rect 324 17442 329 17476
rect 367 17459 438 17476
rect 367 17442 442 17459
rect 400 17441 442 17442
rect 378 17435 464 17441
rect 38 17419 80 17435
rect 400 17419 442 17435
rect -25 17405 25 17407
rect 42 17405 76 17419
rect 404 17405 438 17419
rect 455 17405 505 17407
rect 557 17405 607 17407
rect 16 17397 102 17405
rect 378 17397 464 17405
rect 8 17363 17 17397
rect 18 17395 51 17397
rect 80 17395 100 17397
rect 18 17363 100 17395
rect 380 17395 404 17397
rect 429 17395 438 17397
rect 442 17395 462 17397
rect 16 17355 102 17363
rect 42 17339 76 17355
rect 16 17319 38 17325
rect 42 17316 76 17320
rect 80 17319 102 17325
rect 42 17286 46 17316
rect 72 17286 76 17316
rect 42 17205 46 17239
rect 72 17205 76 17239
rect -25 17168 25 17170
rect -8 17160 14 17167
rect -8 17159 17 17160
rect 25 17159 27 17168
rect -12 17152 38 17159
rect -12 17151 34 17152
rect -12 17147 8 17151
rect 0 17135 8 17147
rect 14 17135 34 17151
rect 0 17134 34 17135
rect 0 17127 38 17134
rect 14 17126 17 17127
rect 25 17118 27 17127
rect 42 17098 45 17188
rect 69 17173 80 17205
rect 107 17173 143 17201
rect 144 17173 148 17393
rect 332 17325 336 17393
rect 380 17363 462 17395
rect 463 17363 472 17397
rect 480 17363 497 17397
rect 378 17355 464 17363
rect 505 17355 507 17405
rect 514 17363 548 17397
rect 565 17363 582 17397
rect 607 17355 609 17405
rect 404 17339 438 17355
rect 400 17325 442 17326
rect 378 17319 404 17325
rect 442 17319 464 17325
rect 400 17318 404 17319
rect 174 17279 246 17287
rect 295 17284 300 17318
rect 324 17284 329 17318
rect 224 17249 226 17265
rect 196 17241 226 17249
rect 332 17247 336 17315
rect 367 17284 438 17318
rect 400 17277 404 17284
rect 454 17271 504 17273
rect 494 17267 548 17271
rect 494 17262 514 17267
rect 504 17247 506 17262
rect 196 17237 232 17241
rect 196 17207 204 17237
rect 216 17207 232 17237
rect 400 17239 404 17247
rect 107 17167 119 17173
rect 109 17139 119 17167
rect 129 17139 149 17173
rect 174 17169 181 17199
rect 224 17160 226 17207
rect 256 17199 328 17207
rect 332 17205 336 17235
rect 400 17205 408 17239
rect 434 17205 438 17239
rect 498 17237 506 17247
rect 514 17237 515 17257
rect 504 17221 506 17237
rect 525 17228 528 17262
rect 547 17237 548 17257
rect 557 17237 564 17247
rect 514 17221 530 17227
rect 532 17221 548 17227
rect 278 17169 305 17180
rect 42 17047 46 17081
rect 72 17047 76 17081
rect 38 17009 80 17010
rect 42 16968 76 17002
rect 79 16968 113 17002
rect 42 16889 46 16923
rect 72 16889 76 16923
rect -25 16852 25 16854
rect -8 16844 14 16851
rect -8 16843 17 16844
rect 25 16843 27 16852
rect -12 16836 38 16843
rect -12 16835 34 16836
rect -12 16831 8 16835
rect 0 16819 8 16831
rect 14 16819 34 16835
rect 0 16818 34 16819
rect 0 16811 38 16818
rect 14 16810 17 16811
rect 25 16802 27 16811
rect 42 16782 45 16872
rect 71 16841 80 16869
rect 69 16803 80 16841
rect 144 16831 148 17139
rect 196 17126 204 17160
rect 216 17126 232 17160
rect 244 17156 257 17160
rect 300 17156 308 17169
rect 332 17167 342 17205
rect 400 17197 404 17205
rect 336 17157 342 17167
rect 244 17132 291 17156
rect 244 17126 257 17132
rect 224 17079 226 17126
rect 278 17122 291 17132
rect 300 17132 329 17156
rect 332 17147 342 17157
rect 400 17157 409 17185
rect 562 17168 612 17170
rect 466 17159 497 17167
rect 565 17159 596 17167
rect 300 17122 321 17132
rect 300 17116 308 17122
rect 289 17106 308 17116
rect 196 17049 204 17079
rect 216 17049 232 17079
rect 196 17045 232 17049
rect 196 17037 226 17045
rect 300 17037 308 17106
rect 332 17113 351 17147
rect 361 17119 381 17147
rect 361 17113 375 17119
rect 400 17113 411 17157
rect 442 17152 500 17159
rect 466 17151 500 17152
rect 565 17151 599 17159
rect 497 17135 500 17151
rect 596 17135 599 17151
rect 466 17134 500 17135
rect 442 17127 500 17134
rect 565 17127 599 17135
rect 612 17118 614 17168
rect 332 17089 342 17113
rect 336 17077 342 17089
rect 224 17021 226 17037
rect 332 17009 342 17077
rect 400 17081 404 17089
rect 400 17047 408 17081
rect 434 17047 438 17081
rect 454 17065 504 17067
rect 504 17049 506 17065
rect 514 17059 530 17065
rect 532 17059 548 17065
rect 525 17049 548 17058
rect 400 17039 404 17047
rect 498 17039 506 17049
rect 504 17015 506 17039
rect 514 17029 515 17049
rect 525 17024 528 17049
rect 547 17029 548 17049
rect 557 17039 564 17049
rect 514 17015 548 17019
rect 151 16968 156 17002
rect 174 16999 246 17007
rect 256 16999 328 17007
rect 336 17001 342 17009
rect 400 17004 404 17009
rect 180 16971 185 16999
rect 174 16963 246 16971
rect 256 16963 328 16971
rect 332 16969 336 16999
rect 400 16970 438 17004
rect 224 16933 226 16949
rect 196 16925 226 16933
rect 196 16921 232 16925
rect 196 16891 204 16921
rect 216 16891 232 16921
rect 224 16844 226 16891
rect 300 16864 308 16933
rect 332 16931 342 16969
rect 400 16961 404 16970
rect 454 16955 504 16957
rect 494 16951 548 16955
rect 494 16946 514 16951
rect 504 16931 506 16946
rect 336 16919 342 16931
rect 289 16854 308 16864
rect 300 16848 308 16854
rect 332 16885 342 16919
rect 400 16923 404 16931
rect 400 16889 408 16923
rect 434 16889 438 16923
rect 498 16921 506 16931
rect 514 16921 515 16941
rect 504 16905 506 16921
rect 525 16912 528 16946
rect 547 16921 548 16941
rect 557 16921 564 16931
rect 514 16905 530 16911
rect 532 16905 548 16911
rect 332 16857 373 16885
rect 332 16851 351 16857
rect 107 16797 119 16831
rect 129 16797 149 16831
rect 196 16810 204 16844
rect 216 16810 232 16844
rect 244 16838 257 16844
rect 278 16838 291 16848
rect 244 16814 291 16838
rect 300 16838 321 16848
rect 336 16841 351 16851
rect 300 16814 329 16838
rect 332 16823 351 16841
rect 361 16851 375 16857
rect 400 16851 411 16889
rect 562 16852 612 16854
rect 361 16823 381 16851
rect 400 16823 409 16851
rect 466 16843 497 16851
rect 565 16843 596 16851
rect 442 16836 500 16843
rect 466 16835 500 16836
rect 565 16835 599 16843
rect 244 16810 257 16814
rect 42 16731 46 16765
rect 72 16731 76 16765
rect 42 16684 76 16688
rect 42 16669 46 16684
rect 72 16669 76 16684
rect 38 16651 80 16669
rect 16 16645 102 16651
rect 144 16645 148 16797
rect 174 16773 181 16801
rect 224 16763 226 16810
rect 300 16801 308 16814
rect 278 16790 305 16801
rect 332 16773 342 16823
rect 400 16803 404 16823
rect 497 16819 500 16835
rect 596 16819 599 16835
rect 466 16818 500 16819
rect 442 16811 500 16818
rect 565 16811 599 16819
rect 612 16802 614 16852
rect 256 16763 328 16771
rect 336 16765 342 16773
rect 400 16765 404 16773
rect 196 16733 204 16763
rect 216 16733 232 16763
rect 196 16729 232 16733
rect 196 16721 226 16729
rect 224 16705 226 16721
rect 332 16693 336 16761
rect 400 16731 408 16765
rect 434 16731 438 16765
rect 454 16749 504 16751
rect 504 16733 506 16749
rect 514 16743 530 16749
rect 532 16743 548 16749
rect 525 16733 548 16742
rect 400 16723 404 16731
rect 498 16723 506 16733
rect 504 16699 506 16723
rect 514 16713 515 16733
rect 525 16708 528 16733
rect 547 16713 548 16733
rect 557 16723 564 16733
rect 514 16699 548 16703
rect 400 16693 442 16694
rect 174 16683 246 16691
rect 400 16686 404 16693
rect 295 16652 300 16686
rect 324 16652 329 16686
rect 367 16669 438 16686
rect 367 16652 442 16669
rect 400 16651 442 16652
rect 378 16645 464 16651
rect 38 16629 80 16645
rect 400 16629 442 16645
rect -25 16615 25 16617
rect 42 16615 76 16629
rect 404 16615 438 16629
rect 455 16615 505 16617
rect 557 16615 607 16617
rect 16 16607 102 16615
rect 378 16607 464 16615
rect 8 16573 17 16607
rect 18 16605 51 16607
rect 80 16605 100 16607
rect 18 16573 100 16605
rect 380 16605 404 16607
rect 429 16605 438 16607
rect 442 16605 462 16607
rect 16 16565 102 16573
rect 42 16549 76 16565
rect 16 16529 38 16535
rect 42 16526 76 16530
rect 80 16529 102 16535
rect 42 16496 46 16526
rect 72 16496 76 16526
rect 42 16415 46 16449
rect 72 16415 76 16449
rect -25 16378 25 16380
rect -8 16370 14 16377
rect -8 16369 17 16370
rect 25 16369 27 16378
rect -12 16362 38 16369
rect -12 16361 34 16362
rect -12 16357 8 16361
rect 0 16345 8 16357
rect 14 16345 34 16361
rect 0 16344 34 16345
rect 0 16337 38 16344
rect 14 16336 17 16337
rect 25 16328 27 16337
rect 42 16308 45 16398
rect 69 16383 80 16415
rect 107 16383 143 16411
rect 144 16383 148 16603
rect 332 16535 336 16603
rect 380 16573 462 16605
rect 463 16573 472 16607
rect 480 16573 497 16607
rect 378 16565 464 16573
rect 505 16565 507 16615
rect 514 16573 548 16607
rect 565 16573 582 16607
rect 607 16565 609 16615
rect 404 16549 438 16565
rect 400 16535 442 16536
rect 378 16529 404 16535
rect 442 16529 464 16535
rect 400 16528 404 16529
rect 174 16489 246 16497
rect 295 16494 300 16528
rect 324 16494 329 16528
rect 224 16459 226 16475
rect 196 16451 226 16459
rect 332 16457 336 16525
rect 367 16494 438 16528
rect 400 16487 404 16494
rect 454 16481 504 16483
rect 494 16477 548 16481
rect 494 16472 514 16477
rect 504 16457 506 16472
rect 196 16447 232 16451
rect 196 16417 204 16447
rect 216 16417 232 16447
rect 400 16449 404 16457
rect 107 16377 119 16383
rect 109 16349 119 16377
rect 129 16349 149 16383
rect 174 16379 181 16409
rect 224 16370 226 16417
rect 256 16409 328 16417
rect 332 16415 336 16445
rect 400 16415 408 16449
rect 434 16415 438 16449
rect 498 16447 506 16457
rect 514 16447 515 16467
rect 504 16431 506 16447
rect 525 16438 528 16472
rect 547 16447 548 16467
rect 557 16447 564 16457
rect 514 16431 530 16437
rect 532 16431 548 16437
rect 278 16379 305 16390
rect 42 16257 46 16291
rect 72 16257 76 16291
rect 38 16219 80 16220
rect 42 16178 76 16212
rect 79 16178 113 16212
rect 42 16099 46 16133
rect 72 16099 76 16133
rect -25 16062 25 16064
rect -8 16054 14 16061
rect -8 16053 17 16054
rect 25 16053 27 16062
rect -12 16046 38 16053
rect -12 16045 34 16046
rect -12 16041 8 16045
rect 0 16029 8 16041
rect 14 16029 34 16045
rect 0 16028 34 16029
rect 0 16021 38 16028
rect 14 16020 17 16021
rect 25 16012 27 16021
rect 42 15992 45 16082
rect 71 16051 80 16079
rect 69 16013 80 16051
rect 144 16041 148 16349
rect 196 16336 204 16370
rect 216 16336 232 16370
rect 244 16366 257 16370
rect 300 16366 308 16379
rect 332 16377 342 16415
rect 400 16407 404 16415
rect 336 16367 342 16377
rect 244 16342 291 16366
rect 244 16336 257 16342
rect 224 16289 226 16336
rect 278 16332 291 16342
rect 300 16342 329 16366
rect 332 16357 342 16367
rect 400 16367 409 16395
rect 562 16378 612 16380
rect 466 16369 497 16377
rect 565 16369 596 16377
rect 300 16332 321 16342
rect 300 16326 308 16332
rect 289 16316 308 16326
rect 196 16259 204 16289
rect 216 16259 232 16289
rect 196 16255 232 16259
rect 196 16247 226 16255
rect 300 16247 308 16316
rect 332 16323 351 16357
rect 361 16329 381 16357
rect 361 16323 375 16329
rect 400 16323 411 16367
rect 442 16362 500 16369
rect 466 16361 500 16362
rect 565 16361 599 16369
rect 497 16345 500 16361
rect 596 16345 599 16361
rect 466 16344 500 16345
rect 442 16337 500 16344
rect 565 16337 599 16345
rect 612 16328 614 16378
rect 332 16299 342 16323
rect 336 16287 342 16299
rect 224 16231 226 16247
rect 332 16219 342 16287
rect 400 16291 404 16299
rect 400 16257 408 16291
rect 434 16257 438 16291
rect 454 16275 504 16277
rect 504 16259 506 16275
rect 514 16269 530 16275
rect 532 16269 548 16275
rect 525 16259 548 16268
rect 400 16249 404 16257
rect 498 16249 506 16259
rect 504 16225 506 16249
rect 514 16239 515 16259
rect 525 16234 528 16259
rect 547 16239 548 16259
rect 557 16249 564 16259
rect 514 16225 548 16229
rect 151 16178 156 16212
rect 174 16209 246 16217
rect 256 16209 328 16217
rect 336 16211 342 16219
rect 400 16214 404 16219
rect 180 16181 185 16209
rect 174 16173 246 16181
rect 256 16173 328 16181
rect 332 16179 336 16209
rect 400 16180 438 16214
rect 224 16143 226 16159
rect 196 16135 226 16143
rect 196 16131 232 16135
rect 196 16101 204 16131
rect 216 16101 232 16131
rect 224 16054 226 16101
rect 300 16074 308 16143
rect 332 16141 342 16179
rect 400 16171 404 16180
rect 454 16165 504 16167
rect 494 16161 548 16165
rect 494 16156 514 16161
rect 504 16141 506 16156
rect 336 16129 342 16141
rect 289 16064 308 16074
rect 300 16058 308 16064
rect 332 16095 342 16129
rect 400 16133 404 16141
rect 400 16099 408 16133
rect 434 16099 438 16133
rect 498 16131 506 16141
rect 514 16131 515 16151
rect 504 16115 506 16131
rect 525 16122 528 16156
rect 547 16131 548 16151
rect 557 16131 564 16141
rect 514 16115 530 16121
rect 532 16115 548 16121
rect 332 16067 373 16095
rect 332 16061 351 16067
rect 107 16007 119 16041
rect 129 16007 149 16041
rect 196 16020 204 16054
rect 216 16020 232 16054
rect 244 16048 257 16054
rect 278 16048 291 16058
rect 244 16024 291 16048
rect 300 16048 321 16058
rect 336 16051 351 16061
rect 300 16024 329 16048
rect 332 16033 351 16051
rect 361 16061 375 16067
rect 400 16061 411 16099
rect 562 16062 612 16064
rect 361 16033 381 16061
rect 400 16033 409 16061
rect 466 16053 497 16061
rect 565 16053 596 16061
rect 442 16046 500 16053
rect 466 16045 500 16046
rect 565 16045 599 16053
rect 244 16020 257 16024
rect 42 15941 46 15975
rect 72 15941 76 15975
rect 42 15894 76 15898
rect 42 15879 46 15894
rect 72 15879 76 15894
rect 38 15861 80 15879
rect 16 15855 102 15861
rect 144 15855 148 16007
rect 174 15983 181 16011
rect 224 15973 226 16020
rect 300 16011 308 16024
rect 278 16000 305 16011
rect 332 15983 342 16033
rect 400 16013 404 16033
rect 497 16029 500 16045
rect 596 16029 599 16045
rect 466 16028 500 16029
rect 442 16021 500 16028
rect 565 16021 599 16029
rect 612 16012 614 16062
rect 256 15973 328 15981
rect 336 15975 342 15983
rect 400 15975 404 15983
rect 196 15943 204 15973
rect 216 15943 232 15973
rect 196 15939 232 15943
rect 196 15931 226 15939
rect 224 15915 226 15931
rect 332 15903 336 15971
rect 400 15941 408 15975
rect 434 15941 438 15975
rect 454 15959 504 15961
rect 504 15943 506 15959
rect 514 15953 530 15959
rect 532 15953 548 15959
rect 525 15943 548 15952
rect 400 15933 404 15941
rect 498 15933 506 15943
rect 504 15909 506 15933
rect 514 15923 515 15943
rect 525 15918 528 15943
rect 547 15923 548 15943
rect 557 15933 564 15943
rect 514 15909 548 15913
rect 400 15903 442 15904
rect 174 15893 246 15901
rect 400 15896 404 15903
rect 295 15862 300 15896
rect 324 15862 329 15896
rect 367 15879 438 15896
rect 367 15862 442 15879
rect 400 15861 442 15862
rect 378 15855 464 15861
rect 38 15839 80 15855
rect 400 15839 442 15855
rect -25 15825 25 15827
rect 42 15825 76 15839
rect 404 15825 438 15839
rect 455 15825 505 15827
rect 557 15825 607 15827
rect 16 15817 102 15825
rect 378 15817 464 15825
rect 8 15783 17 15817
rect 18 15815 51 15817
rect 80 15815 100 15817
rect 18 15783 100 15815
rect 380 15815 404 15817
rect 429 15815 438 15817
rect 442 15815 462 15817
rect 16 15775 102 15783
rect 42 15759 76 15775
rect 16 15739 38 15745
rect 42 15736 76 15740
rect 80 15739 102 15745
rect 42 15706 46 15736
rect 72 15706 76 15736
rect 42 15625 46 15659
rect 72 15625 76 15659
rect -25 15588 25 15590
rect -8 15580 14 15587
rect -8 15579 17 15580
rect 25 15579 27 15588
rect -12 15572 38 15579
rect -12 15571 34 15572
rect -12 15567 8 15571
rect 0 15555 8 15567
rect 14 15555 34 15571
rect 0 15554 34 15555
rect 0 15547 38 15554
rect 14 15546 17 15547
rect 25 15538 27 15547
rect 42 15518 45 15608
rect 69 15593 80 15625
rect 107 15593 143 15621
rect 144 15593 148 15813
rect 332 15745 336 15813
rect 380 15783 462 15815
rect 463 15783 472 15817
rect 480 15783 497 15817
rect 378 15775 464 15783
rect 505 15775 507 15825
rect 514 15783 548 15817
rect 565 15783 582 15817
rect 607 15775 609 15825
rect 404 15759 438 15775
rect 400 15745 442 15746
rect 378 15739 404 15745
rect 442 15739 464 15745
rect 400 15738 404 15739
rect 174 15699 246 15707
rect 295 15704 300 15738
rect 324 15704 329 15738
rect 224 15669 226 15685
rect 196 15661 226 15669
rect 332 15667 336 15735
rect 367 15704 438 15738
rect 400 15697 404 15704
rect 454 15691 504 15693
rect 494 15687 548 15691
rect 494 15682 514 15687
rect 504 15667 506 15682
rect 196 15657 232 15661
rect 196 15627 204 15657
rect 216 15627 232 15657
rect 400 15659 404 15667
rect 107 15587 119 15593
rect 109 15559 119 15587
rect 129 15559 149 15593
rect 174 15589 181 15619
rect 224 15580 226 15627
rect 256 15619 328 15627
rect 332 15625 336 15655
rect 400 15625 408 15659
rect 434 15625 438 15659
rect 498 15657 506 15667
rect 514 15657 515 15677
rect 504 15641 506 15657
rect 525 15648 528 15682
rect 547 15657 548 15677
rect 557 15657 564 15667
rect 514 15641 530 15647
rect 532 15641 548 15647
rect 278 15589 305 15600
rect 42 15467 46 15501
rect 72 15467 76 15501
rect 38 15429 80 15430
rect 42 15388 76 15422
rect 79 15388 113 15422
rect 42 15309 46 15343
rect 72 15309 76 15343
rect -25 15272 25 15274
rect -8 15264 14 15271
rect -8 15263 17 15264
rect 25 15263 27 15272
rect -12 15256 38 15263
rect -12 15255 34 15256
rect -12 15251 8 15255
rect 0 15239 8 15251
rect 14 15239 34 15255
rect 0 15238 34 15239
rect 0 15231 38 15238
rect 14 15230 17 15231
rect 25 15222 27 15231
rect 42 15202 45 15292
rect 71 15261 80 15289
rect 69 15223 80 15261
rect 144 15251 148 15559
rect 196 15546 204 15580
rect 216 15546 232 15580
rect 244 15576 257 15580
rect 300 15576 308 15589
rect 332 15587 342 15625
rect 400 15617 404 15625
rect 336 15577 342 15587
rect 244 15552 291 15576
rect 244 15546 257 15552
rect 224 15499 226 15546
rect 278 15542 291 15552
rect 300 15552 329 15576
rect 332 15567 342 15577
rect 400 15577 409 15605
rect 562 15588 612 15590
rect 466 15579 497 15587
rect 565 15579 596 15587
rect 300 15542 321 15552
rect 300 15536 308 15542
rect 289 15526 308 15536
rect 196 15469 204 15499
rect 216 15469 232 15499
rect 196 15465 232 15469
rect 196 15457 226 15465
rect 300 15457 308 15526
rect 332 15533 351 15567
rect 361 15539 381 15567
rect 361 15533 375 15539
rect 400 15533 411 15577
rect 442 15572 500 15579
rect 466 15571 500 15572
rect 565 15571 599 15579
rect 497 15555 500 15571
rect 596 15555 599 15571
rect 466 15554 500 15555
rect 442 15547 500 15554
rect 565 15547 599 15555
rect 612 15538 614 15588
rect 332 15509 342 15533
rect 336 15497 342 15509
rect 224 15441 226 15457
rect 332 15429 342 15497
rect 400 15501 404 15509
rect 400 15467 408 15501
rect 434 15467 438 15501
rect 454 15485 504 15487
rect 504 15469 506 15485
rect 514 15479 530 15485
rect 532 15479 548 15485
rect 525 15469 548 15478
rect 400 15459 404 15467
rect 498 15459 506 15469
rect 504 15435 506 15459
rect 514 15449 515 15469
rect 525 15444 528 15469
rect 547 15449 548 15469
rect 557 15459 564 15469
rect 514 15435 548 15439
rect 151 15388 156 15422
rect 174 15419 246 15427
rect 256 15419 328 15427
rect 336 15421 342 15429
rect 400 15424 404 15429
rect 180 15391 185 15419
rect 174 15383 246 15391
rect 256 15383 328 15391
rect 332 15389 336 15419
rect 400 15390 438 15424
rect 224 15353 226 15369
rect 196 15345 226 15353
rect 196 15341 232 15345
rect 196 15311 204 15341
rect 216 15311 232 15341
rect 224 15264 226 15311
rect 300 15284 308 15353
rect 332 15351 342 15389
rect 400 15381 404 15390
rect 454 15375 504 15377
rect 494 15371 548 15375
rect 494 15366 514 15371
rect 504 15351 506 15366
rect 336 15339 342 15351
rect 289 15274 308 15284
rect 300 15268 308 15274
rect 332 15305 342 15339
rect 400 15343 404 15351
rect 400 15309 408 15343
rect 434 15309 438 15343
rect 498 15341 506 15351
rect 514 15341 515 15361
rect 504 15325 506 15341
rect 525 15332 528 15366
rect 547 15341 548 15361
rect 557 15341 564 15351
rect 514 15325 530 15331
rect 532 15325 548 15331
rect 332 15277 373 15305
rect 332 15271 351 15277
rect 107 15217 119 15251
rect 129 15217 149 15251
rect 196 15230 204 15264
rect 216 15230 232 15264
rect 244 15258 257 15264
rect 278 15258 291 15268
rect 244 15234 291 15258
rect 300 15258 321 15268
rect 336 15261 351 15271
rect 300 15234 329 15258
rect 332 15243 351 15261
rect 361 15271 375 15277
rect 400 15271 411 15309
rect 562 15272 612 15274
rect 361 15243 381 15271
rect 400 15243 409 15271
rect 466 15263 497 15271
rect 565 15263 596 15271
rect 442 15256 500 15263
rect 466 15255 500 15256
rect 565 15255 599 15263
rect 244 15230 257 15234
rect 42 15151 46 15185
rect 72 15151 76 15185
rect 42 15104 76 15108
rect 42 15089 46 15104
rect 72 15089 76 15104
rect 38 15071 80 15089
rect 16 15065 102 15071
rect 144 15065 148 15217
rect 174 15193 181 15221
rect 224 15183 226 15230
rect 300 15221 308 15234
rect 278 15210 305 15221
rect 332 15193 342 15243
rect 400 15223 404 15243
rect 497 15239 500 15255
rect 596 15239 599 15255
rect 466 15238 500 15239
rect 442 15231 500 15238
rect 565 15231 599 15239
rect 612 15222 614 15272
rect 256 15183 328 15191
rect 336 15185 342 15193
rect 400 15185 404 15193
rect 196 15153 204 15183
rect 216 15153 232 15183
rect 196 15149 232 15153
rect 196 15141 226 15149
rect 224 15125 226 15141
rect 332 15113 336 15181
rect 400 15151 408 15185
rect 434 15151 438 15185
rect 454 15169 504 15171
rect 504 15153 506 15169
rect 514 15163 530 15169
rect 532 15163 548 15169
rect 525 15153 548 15162
rect 400 15143 404 15151
rect 498 15143 506 15153
rect 504 15119 506 15143
rect 514 15133 515 15153
rect 525 15128 528 15153
rect 547 15133 548 15153
rect 557 15143 564 15153
rect 514 15119 548 15123
rect 400 15113 442 15114
rect 174 15103 246 15111
rect 400 15106 404 15113
rect 295 15072 300 15106
rect 324 15072 329 15106
rect 367 15089 438 15106
rect 367 15072 442 15089
rect 400 15071 442 15072
rect 378 15065 464 15071
rect 38 15049 80 15065
rect 400 15049 442 15065
rect -25 15035 25 15037
rect 42 15035 76 15049
rect 404 15035 438 15049
rect 455 15035 505 15037
rect 557 15035 607 15037
rect 16 15027 102 15035
rect 378 15027 464 15035
rect 8 14993 17 15027
rect 18 15025 51 15027
rect 80 15025 100 15027
rect 18 14993 100 15025
rect 380 15025 404 15027
rect 429 15025 438 15027
rect 442 15025 462 15027
rect 16 14985 102 14993
rect 42 14969 76 14985
rect 16 14949 38 14955
rect 42 14946 76 14950
rect 80 14949 102 14955
rect 42 14916 46 14946
rect 72 14916 76 14946
rect 42 14835 46 14869
rect 72 14835 76 14869
rect -25 14798 25 14800
rect -8 14790 14 14797
rect -8 14789 17 14790
rect 25 14789 27 14798
rect -12 14782 38 14789
rect -12 14781 34 14782
rect -12 14777 8 14781
rect 0 14765 8 14777
rect 14 14765 34 14781
rect 0 14764 34 14765
rect 0 14757 38 14764
rect 14 14756 17 14757
rect 25 14748 27 14757
rect 42 14728 45 14818
rect 69 14803 80 14835
rect 107 14803 143 14831
rect 144 14803 148 15023
rect 332 14955 336 15023
rect 380 14993 462 15025
rect 463 14993 472 15027
rect 480 14993 497 15027
rect 378 14985 464 14993
rect 505 14985 507 15035
rect 514 14993 548 15027
rect 565 14993 582 15027
rect 607 14985 609 15035
rect 404 14969 438 14985
rect 400 14955 442 14956
rect 378 14949 404 14955
rect 442 14949 464 14955
rect 400 14948 404 14949
rect 174 14909 246 14917
rect 295 14914 300 14948
rect 324 14914 329 14948
rect 224 14879 226 14895
rect 196 14871 226 14879
rect 332 14877 336 14945
rect 367 14914 438 14948
rect 400 14907 404 14914
rect 454 14901 504 14903
rect 494 14897 548 14901
rect 494 14892 514 14897
rect 504 14877 506 14892
rect 196 14867 232 14871
rect 196 14837 204 14867
rect 216 14837 232 14867
rect 400 14869 404 14877
rect 107 14797 119 14803
rect 109 14769 119 14797
rect 129 14769 149 14803
rect 174 14799 181 14829
rect 224 14790 226 14837
rect 256 14829 328 14837
rect 332 14835 336 14865
rect 400 14835 408 14869
rect 434 14835 438 14869
rect 498 14867 506 14877
rect 514 14867 515 14887
rect 504 14851 506 14867
rect 525 14858 528 14892
rect 547 14867 548 14887
rect 557 14867 564 14877
rect 514 14851 530 14857
rect 532 14851 548 14857
rect 278 14799 305 14810
rect 42 14677 46 14711
rect 72 14677 76 14711
rect 38 14639 80 14640
rect 42 14598 76 14632
rect 79 14598 113 14632
rect 42 14519 46 14553
rect 72 14519 76 14553
rect -25 14482 25 14484
rect -8 14474 14 14481
rect -8 14473 17 14474
rect 25 14473 27 14482
rect -12 14466 38 14473
rect -12 14465 34 14466
rect -12 14461 8 14465
rect 0 14449 8 14461
rect 14 14449 34 14465
rect 0 14448 34 14449
rect 0 14441 38 14448
rect 14 14440 17 14441
rect 25 14432 27 14441
rect 42 14412 45 14502
rect 71 14471 80 14499
rect 69 14433 80 14471
rect 144 14461 148 14769
rect 196 14756 204 14790
rect 216 14756 232 14790
rect 244 14786 257 14790
rect 300 14786 308 14799
rect 332 14797 342 14835
rect 400 14827 404 14835
rect 336 14787 342 14797
rect 244 14762 291 14786
rect 244 14756 257 14762
rect 224 14709 226 14756
rect 278 14752 291 14762
rect 300 14762 329 14786
rect 332 14777 342 14787
rect 400 14787 409 14815
rect 562 14798 612 14800
rect 466 14789 497 14797
rect 565 14789 596 14797
rect 300 14752 321 14762
rect 300 14746 308 14752
rect 289 14736 308 14746
rect 196 14679 204 14709
rect 216 14679 232 14709
rect 196 14675 232 14679
rect 196 14667 226 14675
rect 300 14667 308 14736
rect 332 14743 351 14777
rect 361 14749 381 14777
rect 361 14743 375 14749
rect 400 14743 411 14787
rect 442 14782 500 14789
rect 466 14781 500 14782
rect 565 14781 599 14789
rect 497 14765 500 14781
rect 596 14765 599 14781
rect 466 14764 500 14765
rect 442 14757 500 14764
rect 565 14757 599 14765
rect 612 14748 614 14798
rect 332 14719 342 14743
rect 336 14707 342 14719
rect 224 14651 226 14667
rect 332 14639 342 14707
rect 400 14711 404 14719
rect 400 14677 408 14711
rect 434 14677 438 14711
rect 454 14695 504 14697
rect 504 14679 506 14695
rect 514 14689 530 14695
rect 532 14689 548 14695
rect 525 14679 548 14688
rect 400 14669 404 14677
rect 498 14669 506 14679
rect 504 14645 506 14669
rect 514 14659 515 14679
rect 525 14654 528 14679
rect 547 14659 548 14679
rect 557 14669 564 14679
rect 514 14645 548 14649
rect 151 14598 156 14632
rect 174 14629 246 14637
rect 256 14629 328 14637
rect 336 14631 342 14639
rect 400 14634 404 14639
rect 180 14601 185 14629
rect 174 14593 246 14601
rect 256 14593 328 14601
rect 332 14599 336 14629
rect 400 14600 438 14634
rect 224 14563 226 14579
rect 196 14555 226 14563
rect 196 14551 232 14555
rect 196 14521 204 14551
rect 216 14521 232 14551
rect 224 14474 226 14521
rect 300 14494 308 14563
rect 332 14561 342 14599
rect 400 14591 404 14600
rect 454 14585 504 14587
rect 494 14581 548 14585
rect 494 14576 514 14581
rect 504 14561 506 14576
rect 336 14549 342 14561
rect 289 14484 308 14494
rect 300 14478 308 14484
rect 332 14515 342 14549
rect 400 14553 404 14561
rect 400 14519 408 14553
rect 434 14519 438 14553
rect 498 14551 506 14561
rect 514 14551 515 14571
rect 504 14535 506 14551
rect 525 14542 528 14576
rect 547 14551 548 14571
rect 557 14551 564 14561
rect 514 14535 530 14541
rect 532 14535 548 14541
rect 332 14487 373 14515
rect 332 14481 351 14487
rect 107 14427 119 14461
rect 129 14427 149 14461
rect 196 14440 204 14474
rect 216 14440 232 14474
rect 244 14468 257 14474
rect 278 14468 291 14478
rect 244 14444 291 14468
rect 300 14468 321 14478
rect 336 14471 351 14481
rect 300 14444 329 14468
rect 332 14453 351 14471
rect 361 14481 375 14487
rect 400 14481 411 14519
rect 562 14482 612 14484
rect 361 14453 381 14481
rect 400 14453 409 14481
rect 466 14473 497 14481
rect 565 14473 596 14481
rect 442 14466 500 14473
rect 466 14465 500 14466
rect 565 14465 599 14473
rect 244 14440 257 14444
rect 42 14361 46 14395
rect 72 14361 76 14395
rect 42 14314 76 14318
rect 42 14299 46 14314
rect 72 14299 76 14314
rect 38 14281 80 14299
rect 16 14275 102 14281
rect 144 14275 148 14427
rect 174 14403 181 14431
rect 224 14393 226 14440
rect 300 14431 308 14444
rect 278 14420 305 14431
rect 332 14403 342 14453
rect 400 14433 404 14453
rect 497 14449 500 14465
rect 596 14449 599 14465
rect 466 14448 500 14449
rect 442 14441 500 14448
rect 565 14441 599 14449
rect 612 14432 614 14482
rect 256 14393 328 14401
rect 336 14395 342 14403
rect 400 14395 404 14403
rect 196 14363 204 14393
rect 216 14363 232 14393
rect 196 14359 232 14363
rect 196 14351 226 14359
rect 224 14335 226 14351
rect 332 14323 336 14391
rect 400 14361 408 14395
rect 434 14361 438 14395
rect 454 14379 504 14381
rect 504 14363 506 14379
rect 514 14373 530 14379
rect 532 14373 548 14379
rect 525 14363 548 14372
rect 400 14353 404 14361
rect 498 14353 506 14363
rect 504 14329 506 14353
rect 514 14343 515 14363
rect 525 14338 528 14363
rect 547 14343 548 14363
rect 557 14353 564 14363
rect 514 14329 548 14333
rect 400 14323 442 14324
rect 174 14313 246 14321
rect 400 14316 404 14323
rect 295 14282 300 14316
rect 324 14282 329 14316
rect 367 14299 438 14316
rect 367 14282 442 14299
rect 400 14281 442 14282
rect 378 14275 464 14281
rect 38 14259 80 14275
rect 400 14259 442 14275
rect -25 14245 25 14247
rect 42 14245 76 14259
rect 404 14245 438 14259
rect 455 14245 505 14247
rect 557 14245 607 14247
rect 16 14237 102 14245
rect 378 14237 464 14245
rect 8 14203 17 14237
rect 18 14235 51 14237
rect 80 14235 100 14237
rect 18 14203 100 14235
rect 380 14235 404 14237
rect 429 14235 438 14237
rect 442 14235 462 14237
rect 16 14195 102 14203
rect 42 14179 76 14195
rect 16 14159 38 14165
rect 42 14156 76 14160
rect 80 14159 102 14165
rect 42 14126 46 14156
rect 72 14126 76 14156
rect 42 14045 46 14079
rect 72 14045 76 14079
rect -25 14008 25 14010
rect -8 14000 14 14007
rect -8 13999 17 14000
rect 25 13999 27 14008
rect -12 13992 38 13999
rect -12 13991 34 13992
rect -12 13987 8 13991
rect 0 13975 8 13987
rect 14 13975 34 13991
rect 0 13974 34 13975
rect 0 13967 38 13974
rect 14 13966 17 13967
rect 25 13958 27 13967
rect 42 13938 45 14028
rect 69 14013 80 14045
rect 107 14013 143 14041
rect 144 14013 148 14233
rect 332 14165 336 14233
rect 380 14203 462 14235
rect 463 14203 472 14237
rect 480 14203 497 14237
rect 378 14195 464 14203
rect 505 14195 507 14245
rect 514 14203 548 14237
rect 565 14203 582 14237
rect 607 14195 609 14245
rect 404 14179 438 14195
rect 400 14165 442 14166
rect 378 14159 404 14165
rect 442 14159 464 14165
rect 400 14158 404 14159
rect 174 14119 246 14127
rect 295 14124 300 14158
rect 324 14124 329 14158
rect 224 14089 226 14105
rect 196 14081 226 14089
rect 332 14087 336 14155
rect 367 14124 438 14158
rect 400 14117 404 14124
rect 454 14111 504 14113
rect 494 14107 548 14111
rect 494 14102 514 14107
rect 504 14087 506 14102
rect 196 14077 232 14081
rect 196 14047 204 14077
rect 216 14047 232 14077
rect 400 14079 404 14087
rect 107 14007 119 14013
rect 109 13979 119 14007
rect 129 13979 149 14013
rect 174 14009 181 14039
rect 224 14000 226 14047
rect 256 14039 328 14047
rect 332 14045 336 14075
rect 400 14045 408 14079
rect 434 14045 438 14079
rect 498 14077 506 14087
rect 514 14077 515 14097
rect 504 14061 506 14077
rect 525 14068 528 14102
rect 547 14077 548 14097
rect 557 14077 564 14087
rect 514 14061 530 14067
rect 532 14061 548 14067
rect 278 14009 305 14020
rect 42 13887 46 13921
rect 72 13887 76 13921
rect 38 13849 80 13850
rect 42 13808 76 13842
rect 79 13808 113 13842
rect 42 13729 46 13763
rect 72 13729 76 13763
rect -25 13692 25 13694
rect -8 13684 14 13691
rect -8 13683 17 13684
rect 25 13683 27 13692
rect -12 13676 38 13683
rect -12 13675 34 13676
rect -12 13671 8 13675
rect 0 13659 8 13671
rect 14 13659 34 13675
rect 0 13658 34 13659
rect 0 13651 38 13658
rect 14 13650 17 13651
rect 25 13642 27 13651
rect 42 13622 45 13712
rect 71 13681 80 13709
rect 69 13643 80 13681
rect 144 13671 148 13979
rect 196 13966 204 14000
rect 216 13966 232 14000
rect 244 13996 257 14000
rect 300 13996 308 14009
rect 332 14007 342 14045
rect 400 14037 404 14045
rect 336 13997 342 14007
rect 244 13972 291 13996
rect 244 13966 257 13972
rect 224 13919 226 13966
rect 278 13962 291 13972
rect 300 13972 329 13996
rect 332 13987 342 13997
rect 400 13997 409 14025
rect 562 14008 612 14010
rect 466 13999 497 14007
rect 565 13999 596 14007
rect 300 13962 321 13972
rect 300 13956 308 13962
rect 289 13946 308 13956
rect 196 13889 204 13919
rect 216 13889 232 13919
rect 196 13885 232 13889
rect 196 13877 226 13885
rect 300 13877 308 13946
rect 332 13953 351 13987
rect 361 13959 381 13987
rect 361 13953 375 13959
rect 400 13953 411 13997
rect 442 13992 500 13999
rect 466 13991 500 13992
rect 565 13991 599 13999
rect 497 13975 500 13991
rect 596 13975 599 13991
rect 466 13974 500 13975
rect 442 13967 500 13974
rect 565 13967 599 13975
rect 612 13958 614 14008
rect 332 13929 342 13953
rect 336 13917 342 13929
rect 224 13861 226 13877
rect 332 13849 342 13917
rect 400 13921 404 13929
rect 400 13887 408 13921
rect 434 13887 438 13921
rect 454 13905 504 13907
rect 504 13889 506 13905
rect 514 13899 530 13905
rect 532 13899 548 13905
rect 525 13889 548 13898
rect 400 13879 404 13887
rect 498 13879 506 13889
rect 504 13855 506 13879
rect 514 13869 515 13889
rect 525 13864 528 13889
rect 547 13869 548 13889
rect 557 13879 564 13889
rect 514 13855 548 13859
rect 151 13808 156 13842
rect 174 13839 246 13847
rect 256 13839 328 13847
rect 336 13841 342 13849
rect 400 13844 404 13849
rect 180 13811 185 13839
rect 174 13803 246 13811
rect 256 13803 328 13811
rect 332 13809 336 13839
rect 400 13810 438 13844
rect 224 13773 226 13789
rect 196 13765 226 13773
rect 196 13761 232 13765
rect 196 13731 204 13761
rect 216 13731 232 13761
rect 224 13684 226 13731
rect 300 13704 308 13773
rect 332 13771 342 13809
rect 400 13801 404 13810
rect 454 13795 504 13797
rect 494 13791 548 13795
rect 494 13786 514 13791
rect 504 13771 506 13786
rect 336 13759 342 13771
rect 289 13694 308 13704
rect 300 13688 308 13694
rect 332 13725 342 13759
rect 400 13763 404 13771
rect 400 13729 408 13763
rect 434 13729 438 13763
rect 498 13761 506 13771
rect 514 13761 515 13781
rect 504 13745 506 13761
rect 525 13752 528 13786
rect 547 13761 548 13781
rect 557 13761 564 13771
rect 514 13745 530 13751
rect 532 13745 548 13751
rect 332 13697 373 13725
rect 332 13691 351 13697
rect 107 13637 119 13671
rect 129 13637 149 13671
rect 196 13650 204 13684
rect 216 13650 232 13684
rect 244 13678 257 13684
rect 278 13678 291 13688
rect 244 13654 291 13678
rect 300 13678 321 13688
rect 336 13681 351 13691
rect 300 13654 329 13678
rect 332 13663 351 13681
rect 361 13691 375 13697
rect 400 13691 411 13729
rect 562 13692 612 13694
rect 361 13663 381 13691
rect 400 13663 409 13691
rect 466 13683 497 13691
rect 565 13683 596 13691
rect 442 13676 500 13683
rect 466 13675 500 13676
rect 565 13675 599 13683
rect 244 13650 257 13654
rect 42 13571 46 13605
rect 72 13571 76 13605
rect 42 13524 76 13528
rect 42 13509 46 13524
rect 72 13509 76 13524
rect 38 13491 80 13509
rect 16 13485 102 13491
rect 144 13485 148 13637
rect 174 13613 181 13641
rect 224 13603 226 13650
rect 300 13641 308 13654
rect 278 13630 305 13641
rect 332 13613 342 13663
rect 400 13643 404 13663
rect 497 13659 500 13675
rect 596 13659 599 13675
rect 466 13658 500 13659
rect 442 13651 500 13658
rect 565 13651 599 13659
rect 612 13642 614 13692
rect 256 13603 328 13611
rect 336 13605 342 13613
rect 400 13605 404 13613
rect 196 13573 204 13603
rect 216 13573 232 13603
rect 196 13569 232 13573
rect 196 13561 226 13569
rect 224 13545 226 13561
rect 332 13533 336 13601
rect 400 13571 408 13605
rect 434 13571 438 13605
rect 454 13589 504 13591
rect 504 13573 506 13589
rect 514 13583 530 13589
rect 532 13583 548 13589
rect 525 13573 548 13582
rect 400 13563 404 13571
rect 498 13563 506 13573
rect 504 13539 506 13563
rect 514 13553 515 13573
rect 525 13548 528 13573
rect 547 13553 548 13573
rect 557 13563 564 13573
rect 514 13539 548 13543
rect 400 13533 442 13534
rect 174 13523 246 13531
rect 400 13526 404 13533
rect 295 13492 300 13526
rect 324 13492 329 13526
rect 367 13509 438 13526
rect 367 13492 442 13509
rect 400 13491 442 13492
rect 378 13485 464 13491
rect 38 13469 80 13485
rect 400 13469 442 13485
rect -25 13455 25 13457
rect 42 13455 76 13469
rect 404 13455 438 13469
rect 455 13455 505 13457
rect 557 13455 607 13457
rect 16 13447 102 13455
rect 378 13447 464 13455
rect 8 13413 17 13447
rect 18 13445 51 13447
rect 80 13445 100 13447
rect 18 13413 100 13445
rect 380 13445 404 13447
rect 429 13445 438 13447
rect 442 13445 462 13447
rect 16 13405 102 13413
rect 42 13389 76 13405
rect 16 13369 38 13375
rect 42 13366 76 13370
rect 80 13369 102 13375
rect 42 13336 46 13366
rect 72 13336 76 13366
rect 42 13255 46 13289
rect 72 13255 76 13289
rect -25 13218 25 13220
rect -8 13210 14 13217
rect -8 13209 17 13210
rect 25 13209 27 13218
rect -12 13202 38 13209
rect -12 13201 34 13202
rect -12 13197 8 13201
rect 0 13185 8 13197
rect 14 13185 34 13201
rect 0 13184 34 13185
rect 0 13177 38 13184
rect 14 13176 17 13177
rect 25 13168 27 13177
rect 42 13148 45 13238
rect 69 13223 80 13255
rect 107 13223 143 13251
rect 144 13223 148 13443
rect 332 13375 336 13443
rect 380 13413 462 13445
rect 463 13413 472 13447
rect 480 13413 497 13447
rect 378 13405 464 13413
rect 505 13405 507 13455
rect 514 13413 548 13447
rect 565 13413 582 13447
rect 607 13405 609 13455
rect 404 13389 438 13405
rect 400 13375 442 13376
rect 378 13369 404 13375
rect 442 13369 464 13375
rect 400 13368 404 13369
rect 174 13329 246 13337
rect 295 13334 300 13368
rect 324 13334 329 13368
rect 224 13299 226 13315
rect 196 13291 226 13299
rect 332 13297 336 13365
rect 367 13334 438 13368
rect 400 13327 404 13334
rect 454 13321 504 13323
rect 494 13317 548 13321
rect 494 13312 514 13317
rect 504 13297 506 13312
rect 196 13287 232 13291
rect 196 13257 204 13287
rect 216 13257 232 13287
rect 400 13289 404 13297
rect 107 13217 119 13223
rect 109 13189 119 13217
rect 129 13189 149 13223
rect 174 13219 181 13249
rect 224 13210 226 13257
rect 256 13249 328 13257
rect 332 13255 336 13285
rect 400 13255 408 13289
rect 434 13255 438 13289
rect 498 13287 506 13297
rect 514 13287 515 13307
rect 504 13271 506 13287
rect 525 13278 528 13312
rect 547 13287 548 13307
rect 557 13287 564 13297
rect 514 13271 530 13277
rect 532 13271 548 13277
rect 278 13219 305 13230
rect 42 13097 46 13131
rect 72 13097 76 13131
rect 38 13059 80 13060
rect 42 13018 76 13052
rect 79 13018 113 13052
rect 42 12939 46 12973
rect 72 12939 76 12973
rect -25 12902 25 12904
rect -8 12894 14 12901
rect -8 12893 17 12894
rect 25 12893 27 12902
rect -12 12886 38 12893
rect -12 12885 34 12886
rect -12 12881 8 12885
rect 0 12869 8 12881
rect 14 12869 34 12885
rect 0 12868 34 12869
rect 0 12861 38 12868
rect 14 12860 17 12861
rect 25 12852 27 12861
rect 42 12832 45 12922
rect 71 12891 80 12919
rect 69 12853 80 12891
rect 144 12881 148 13189
rect 196 13176 204 13210
rect 216 13176 232 13210
rect 244 13206 257 13210
rect 300 13206 308 13219
rect 332 13217 342 13255
rect 400 13247 404 13255
rect 336 13207 342 13217
rect 244 13182 291 13206
rect 244 13176 257 13182
rect 224 13129 226 13176
rect 278 13172 291 13182
rect 300 13182 329 13206
rect 332 13197 342 13207
rect 400 13207 409 13235
rect 562 13218 612 13220
rect 466 13209 497 13217
rect 565 13209 596 13217
rect 300 13172 321 13182
rect 300 13166 308 13172
rect 289 13156 308 13166
rect 196 13099 204 13129
rect 216 13099 232 13129
rect 196 13095 232 13099
rect 196 13087 226 13095
rect 300 13087 308 13156
rect 332 13163 351 13197
rect 361 13169 381 13197
rect 361 13163 375 13169
rect 400 13163 411 13207
rect 442 13202 500 13209
rect 466 13201 500 13202
rect 565 13201 599 13209
rect 497 13185 500 13201
rect 596 13185 599 13201
rect 466 13184 500 13185
rect 442 13177 500 13184
rect 565 13177 599 13185
rect 612 13168 614 13218
rect 332 13139 342 13163
rect 336 13127 342 13139
rect 224 13071 226 13087
rect 332 13059 342 13127
rect 400 13131 404 13139
rect 400 13097 408 13131
rect 434 13097 438 13131
rect 454 13115 504 13117
rect 504 13099 506 13115
rect 514 13109 530 13115
rect 532 13109 548 13115
rect 525 13099 548 13108
rect 400 13089 404 13097
rect 498 13089 506 13099
rect 504 13065 506 13089
rect 514 13079 515 13099
rect 525 13074 528 13099
rect 547 13079 548 13099
rect 557 13089 564 13099
rect 514 13065 548 13069
rect 151 13018 156 13052
rect 174 13049 246 13057
rect 256 13049 328 13057
rect 336 13051 342 13059
rect 400 13054 404 13059
rect 180 13021 185 13049
rect 174 13013 246 13021
rect 256 13013 328 13021
rect 332 13019 336 13049
rect 400 13020 438 13054
rect 224 12983 226 12999
rect 196 12975 226 12983
rect 196 12971 232 12975
rect 196 12941 204 12971
rect 216 12941 232 12971
rect 224 12894 226 12941
rect 300 12914 308 12983
rect 332 12981 342 13019
rect 400 13011 404 13020
rect 454 13005 504 13007
rect 494 13001 548 13005
rect 494 12996 514 13001
rect 504 12981 506 12996
rect 336 12969 342 12981
rect 289 12904 308 12914
rect 300 12898 308 12904
rect 332 12935 342 12969
rect 400 12973 404 12981
rect 400 12939 408 12973
rect 434 12939 438 12973
rect 498 12971 506 12981
rect 514 12971 515 12991
rect 504 12955 506 12971
rect 525 12962 528 12996
rect 547 12971 548 12991
rect 557 12971 564 12981
rect 514 12955 530 12961
rect 532 12955 548 12961
rect 332 12907 373 12935
rect 332 12901 351 12907
rect 107 12847 119 12881
rect 129 12847 149 12881
rect 196 12860 204 12894
rect 216 12860 232 12894
rect 244 12888 257 12894
rect 278 12888 291 12898
rect 244 12864 291 12888
rect 300 12888 321 12898
rect 336 12891 351 12901
rect 300 12864 329 12888
rect 332 12873 351 12891
rect 361 12901 375 12907
rect 400 12901 411 12939
rect 562 12902 612 12904
rect 361 12873 381 12901
rect 400 12873 409 12901
rect 466 12893 497 12901
rect 565 12893 596 12901
rect 442 12886 500 12893
rect 466 12885 500 12886
rect 565 12885 599 12893
rect 244 12860 257 12864
rect 42 12781 46 12815
rect 72 12781 76 12815
rect 42 12734 76 12738
rect 42 12719 46 12734
rect 72 12719 76 12734
rect 38 12701 80 12719
rect 16 12695 102 12701
rect 144 12695 148 12847
rect 174 12823 181 12851
rect 224 12813 226 12860
rect 300 12851 308 12864
rect 278 12840 305 12851
rect 332 12823 342 12873
rect 400 12853 404 12873
rect 497 12869 500 12885
rect 596 12869 599 12885
rect 466 12868 500 12869
rect 442 12861 500 12868
rect 565 12861 599 12869
rect 612 12852 614 12902
rect 256 12813 328 12821
rect 336 12815 342 12823
rect 400 12815 404 12823
rect 196 12783 204 12813
rect 216 12783 232 12813
rect 196 12779 232 12783
rect 196 12771 226 12779
rect 224 12755 226 12771
rect 332 12743 336 12811
rect 400 12781 408 12815
rect 434 12781 438 12815
rect 454 12799 504 12801
rect 504 12783 506 12799
rect 514 12793 530 12799
rect 532 12793 548 12799
rect 525 12783 548 12792
rect 400 12773 404 12781
rect 498 12773 506 12783
rect 504 12749 506 12773
rect 514 12763 515 12783
rect 525 12758 528 12783
rect 547 12763 548 12783
rect 557 12773 564 12783
rect 514 12749 548 12753
rect 400 12743 442 12744
rect 174 12733 246 12741
rect 400 12736 404 12743
rect 295 12702 300 12736
rect 324 12702 329 12736
rect 367 12719 438 12736
rect 367 12702 442 12719
rect 400 12701 442 12702
rect 378 12695 464 12701
rect 38 12679 80 12695
rect 400 12679 442 12695
rect -25 12665 25 12667
rect 42 12665 76 12679
rect 404 12665 438 12679
rect 455 12665 505 12667
rect 557 12665 607 12667
rect 16 12657 102 12665
rect 378 12657 464 12665
rect 8 12623 17 12657
rect 18 12655 51 12657
rect 80 12655 100 12657
rect 18 12623 100 12655
rect 380 12655 404 12657
rect 429 12655 438 12657
rect 442 12655 462 12657
rect 16 12615 102 12623
rect 42 12599 76 12615
rect 16 12579 38 12585
rect 42 12576 76 12580
rect 80 12579 102 12585
rect 42 12546 46 12576
rect 72 12546 76 12576
rect 42 12465 46 12499
rect 72 12465 76 12499
rect -25 12428 25 12430
rect -8 12420 14 12427
rect -8 12419 17 12420
rect 25 12419 27 12428
rect -12 12412 38 12419
rect -12 12411 34 12412
rect -12 12407 8 12411
rect 0 12395 8 12407
rect 14 12395 34 12411
rect 0 12394 34 12395
rect 0 12387 38 12394
rect 14 12386 17 12387
rect 25 12378 27 12387
rect 42 12358 45 12448
rect 69 12433 80 12465
rect 107 12433 143 12461
rect 144 12433 148 12653
rect 332 12585 336 12653
rect 380 12623 462 12655
rect 463 12623 472 12657
rect 480 12623 497 12657
rect 378 12615 464 12623
rect 505 12615 507 12665
rect 514 12623 548 12657
rect 565 12623 582 12657
rect 607 12615 609 12665
rect 404 12599 438 12615
rect 400 12585 442 12586
rect 378 12579 404 12585
rect 442 12579 464 12585
rect 400 12578 404 12579
rect 174 12539 246 12547
rect 295 12544 300 12578
rect 324 12544 329 12578
rect 224 12509 226 12525
rect 196 12501 226 12509
rect 332 12507 336 12575
rect 367 12544 438 12578
rect 400 12537 404 12544
rect 454 12531 504 12533
rect 494 12527 548 12531
rect 494 12522 514 12527
rect 504 12507 506 12522
rect 196 12497 232 12501
rect 196 12467 204 12497
rect 216 12467 232 12497
rect 400 12499 404 12507
rect 107 12427 119 12433
rect 109 12399 119 12427
rect 129 12399 149 12433
rect 174 12429 181 12459
rect 224 12420 226 12467
rect 256 12459 328 12467
rect 332 12465 336 12495
rect 400 12465 408 12499
rect 434 12465 438 12499
rect 498 12497 506 12507
rect 514 12497 515 12517
rect 504 12481 506 12497
rect 525 12488 528 12522
rect 547 12497 548 12517
rect 557 12497 564 12507
rect 514 12481 530 12487
rect 532 12481 548 12487
rect 278 12429 305 12440
rect 42 12307 46 12341
rect 72 12307 76 12341
rect 38 12269 80 12270
rect 42 12228 76 12262
rect 79 12228 113 12262
rect 42 12149 46 12183
rect 72 12149 76 12183
rect -25 12112 25 12114
rect -8 12104 14 12111
rect -8 12103 17 12104
rect 25 12103 27 12112
rect -12 12096 38 12103
rect -12 12095 34 12096
rect -12 12091 8 12095
rect 0 12079 8 12091
rect 14 12079 34 12095
rect 0 12078 34 12079
rect 0 12071 38 12078
rect 14 12070 17 12071
rect 25 12062 27 12071
rect 42 12042 45 12132
rect 71 12101 80 12129
rect 69 12063 80 12101
rect 144 12091 148 12399
rect 196 12386 204 12420
rect 216 12386 232 12420
rect 244 12416 257 12420
rect 300 12416 308 12429
rect 332 12427 342 12465
rect 400 12457 404 12465
rect 336 12417 342 12427
rect 244 12392 291 12416
rect 244 12386 257 12392
rect 224 12339 226 12386
rect 278 12382 291 12392
rect 300 12392 329 12416
rect 332 12407 342 12417
rect 400 12417 409 12445
rect 562 12428 612 12430
rect 466 12419 497 12427
rect 565 12419 596 12427
rect 300 12382 321 12392
rect 300 12376 308 12382
rect 289 12366 308 12376
rect 196 12309 204 12339
rect 216 12309 232 12339
rect 196 12305 232 12309
rect 196 12297 226 12305
rect 300 12297 308 12366
rect 332 12373 351 12407
rect 361 12379 381 12407
rect 361 12373 375 12379
rect 400 12373 411 12417
rect 442 12412 500 12419
rect 466 12411 500 12412
rect 565 12411 599 12419
rect 497 12395 500 12411
rect 596 12395 599 12411
rect 466 12394 500 12395
rect 442 12387 500 12394
rect 565 12387 599 12395
rect 612 12378 614 12428
rect 332 12349 342 12373
rect 336 12337 342 12349
rect 224 12281 226 12297
rect 332 12269 342 12337
rect 400 12341 404 12349
rect 400 12307 408 12341
rect 434 12307 438 12341
rect 454 12325 504 12327
rect 504 12309 506 12325
rect 514 12319 530 12325
rect 532 12319 548 12325
rect 525 12309 548 12318
rect 400 12299 404 12307
rect 498 12299 506 12309
rect 504 12275 506 12299
rect 514 12289 515 12309
rect 525 12284 528 12309
rect 547 12289 548 12309
rect 557 12299 564 12309
rect 514 12275 548 12279
rect 151 12228 156 12262
rect 174 12259 246 12267
rect 256 12259 328 12267
rect 336 12261 342 12269
rect 400 12264 404 12269
rect 180 12231 185 12259
rect 174 12223 246 12231
rect 256 12223 328 12231
rect 332 12229 336 12259
rect 400 12230 438 12264
rect 224 12193 226 12209
rect 196 12185 226 12193
rect 196 12181 232 12185
rect 196 12151 204 12181
rect 216 12151 232 12181
rect 224 12104 226 12151
rect 300 12124 308 12193
rect 332 12191 342 12229
rect 400 12221 404 12230
rect 454 12215 504 12217
rect 494 12211 548 12215
rect 494 12206 514 12211
rect 504 12191 506 12206
rect 336 12179 342 12191
rect 289 12114 308 12124
rect 300 12108 308 12114
rect 332 12145 342 12179
rect 400 12183 404 12191
rect 400 12149 408 12183
rect 434 12149 438 12183
rect 498 12181 506 12191
rect 514 12181 515 12201
rect 504 12165 506 12181
rect 525 12172 528 12206
rect 547 12181 548 12201
rect 557 12181 564 12191
rect 514 12165 530 12171
rect 532 12165 548 12171
rect 332 12117 373 12145
rect 332 12111 351 12117
rect 107 12057 119 12091
rect 129 12057 149 12091
rect 196 12070 204 12104
rect 216 12070 232 12104
rect 244 12098 257 12104
rect 278 12098 291 12108
rect 244 12074 291 12098
rect 300 12098 321 12108
rect 336 12101 351 12111
rect 300 12074 329 12098
rect 332 12083 351 12101
rect 361 12111 375 12117
rect 400 12111 411 12149
rect 562 12112 612 12114
rect 361 12083 381 12111
rect 400 12083 409 12111
rect 466 12103 497 12111
rect 565 12103 596 12111
rect 442 12096 500 12103
rect 466 12095 500 12096
rect 565 12095 599 12103
rect 244 12070 257 12074
rect 42 11991 46 12025
rect 72 11991 76 12025
rect 42 11944 76 11948
rect 42 11929 46 11944
rect 72 11929 76 11944
rect 38 11911 80 11929
rect 16 11905 102 11911
rect 144 11905 148 12057
rect 174 12033 181 12061
rect 224 12023 226 12070
rect 300 12061 308 12074
rect 278 12050 305 12061
rect 332 12033 342 12083
rect 400 12063 404 12083
rect 497 12079 500 12095
rect 596 12079 599 12095
rect 466 12078 500 12079
rect 442 12071 500 12078
rect 565 12071 599 12079
rect 612 12062 614 12112
rect 256 12023 328 12031
rect 336 12025 342 12033
rect 400 12025 404 12033
rect 196 11993 204 12023
rect 216 11993 232 12023
rect 196 11989 232 11993
rect 196 11981 226 11989
rect 224 11965 226 11981
rect 332 11953 336 12021
rect 400 11991 408 12025
rect 434 11991 438 12025
rect 454 12009 504 12011
rect 504 11993 506 12009
rect 514 12003 530 12009
rect 532 12003 548 12009
rect 525 11993 548 12002
rect 400 11983 404 11991
rect 498 11983 506 11993
rect 504 11959 506 11983
rect 514 11973 515 11993
rect 525 11968 528 11993
rect 547 11973 548 11993
rect 557 11983 564 11993
rect 514 11959 548 11963
rect 400 11953 442 11954
rect 174 11943 246 11951
rect 400 11946 404 11953
rect 295 11912 300 11946
rect 324 11912 329 11946
rect 367 11929 438 11946
rect 367 11912 442 11929
rect 400 11911 442 11912
rect 378 11905 464 11911
rect 38 11889 80 11905
rect 400 11889 442 11905
rect -25 11875 25 11877
rect 42 11875 76 11889
rect 404 11875 438 11889
rect 455 11875 505 11877
rect 557 11875 607 11877
rect 16 11867 102 11875
rect 378 11867 464 11875
rect 8 11833 17 11867
rect 18 11865 51 11867
rect 80 11865 100 11867
rect 18 11833 100 11865
rect 380 11865 404 11867
rect 429 11865 438 11867
rect 442 11865 462 11867
rect 16 11825 102 11833
rect 42 11809 76 11825
rect 16 11789 38 11795
rect 42 11786 76 11790
rect 80 11789 102 11795
rect 42 11756 46 11786
rect 72 11756 76 11786
rect 42 11675 46 11709
rect 72 11675 76 11709
rect -25 11638 25 11640
rect -8 11630 14 11637
rect -8 11629 17 11630
rect 25 11629 27 11638
rect -12 11622 38 11629
rect -12 11621 34 11622
rect -12 11617 8 11621
rect 0 11605 8 11617
rect 14 11605 34 11621
rect 0 11604 34 11605
rect 0 11597 38 11604
rect 14 11596 17 11597
rect 25 11588 27 11597
rect 42 11568 45 11658
rect 69 11643 80 11675
rect 107 11643 143 11671
rect 144 11643 148 11863
rect 332 11795 336 11863
rect 380 11833 462 11865
rect 463 11833 472 11867
rect 480 11833 497 11867
rect 378 11825 464 11833
rect 505 11825 507 11875
rect 514 11833 548 11867
rect 565 11833 582 11867
rect 607 11825 609 11875
rect 404 11809 438 11825
rect 400 11795 442 11796
rect 378 11789 404 11795
rect 442 11789 464 11795
rect 400 11788 404 11789
rect 174 11749 246 11757
rect 295 11754 300 11788
rect 324 11754 329 11788
rect 224 11719 226 11735
rect 196 11711 226 11719
rect 332 11717 336 11785
rect 367 11754 438 11788
rect 400 11747 404 11754
rect 454 11741 504 11743
rect 494 11737 548 11741
rect 494 11732 514 11737
rect 504 11717 506 11732
rect 196 11707 232 11711
rect 196 11677 204 11707
rect 216 11677 232 11707
rect 400 11709 404 11717
rect 107 11637 119 11643
rect 109 11609 119 11637
rect 129 11609 149 11643
rect 174 11639 181 11669
rect 224 11630 226 11677
rect 256 11669 328 11677
rect 332 11675 336 11705
rect 400 11675 408 11709
rect 434 11675 438 11709
rect 498 11707 506 11717
rect 514 11707 515 11727
rect 504 11691 506 11707
rect 525 11698 528 11732
rect 547 11707 548 11727
rect 557 11707 564 11717
rect 514 11691 530 11697
rect 532 11691 548 11697
rect 278 11639 305 11650
rect 42 11517 46 11551
rect 72 11517 76 11551
rect 38 11479 80 11480
rect 42 11438 76 11472
rect 79 11438 113 11472
rect 42 11359 46 11393
rect 72 11359 76 11393
rect -25 11322 25 11324
rect -8 11314 14 11321
rect -8 11313 17 11314
rect 25 11313 27 11322
rect -12 11306 38 11313
rect -12 11305 34 11306
rect -12 11301 8 11305
rect 0 11289 8 11301
rect 14 11289 34 11305
rect 0 11288 34 11289
rect 0 11281 38 11288
rect 14 11280 17 11281
rect 25 11272 27 11281
rect 42 11252 45 11342
rect 71 11311 80 11339
rect 69 11273 80 11311
rect 144 11301 148 11609
rect 196 11596 204 11630
rect 216 11596 232 11630
rect 244 11626 257 11630
rect 300 11626 308 11639
rect 332 11637 342 11675
rect 400 11667 404 11675
rect 336 11627 342 11637
rect 244 11602 291 11626
rect 244 11596 257 11602
rect 224 11549 226 11596
rect 278 11592 291 11602
rect 300 11602 329 11626
rect 332 11617 342 11627
rect 400 11627 409 11655
rect 562 11638 612 11640
rect 466 11629 497 11637
rect 565 11629 596 11637
rect 300 11592 321 11602
rect 300 11586 308 11592
rect 289 11576 308 11586
rect 196 11519 204 11549
rect 216 11519 232 11549
rect 196 11515 232 11519
rect 196 11507 226 11515
rect 300 11507 308 11576
rect 332 11583 351 11617
rect 361 11589 381 11617
rect 361 11583 375 11589
rect 400 11583 411 11627
rect 442 11622 500 11629
rect 466 11621 500 11622
rect 565 11621 599 11629
rect 497 11605 500 11621
rect 596 11605 599 11621
rect 466 11604 500 11605
rect 442 11597 500 11604
rect 565 11597 599 11605
rect 612 11588 614 11638
rect 332 11559 342 11583
rect 336 11547 342 11559
rect 224 11491 226 11507
rect 332 11479 342 11547
rect 400 11551 404 11559
rect 400 11517 408 11551
rect 434 11517 438 11551
rect 454 11535 504 11537
rect 504 11519 506 11535
rect 514 11529 530 11535
rect 532 11529 548 11535
rect 525 11519 548 11528
rect 400 11509 404 11517
rect 498 11509 506 11519
rect 504 11485 506 11509
rect 514 11499 515 11519
rect 525 11494 528 11519
rect 547 11499 548 11519
rect 557 11509 564 11519
rect 514 11485 548 11489
rect 151 11438 156 11472
rect 174 11469 246 11477
rect 256 11469 328 11477
rect 336 11471 342 11479
rect 400 11474 404 11479
rect 180 11441 185 11469
rect 174 11433 246 11441
rect 256 11433 328 11441
rect 332 11439 336 11469
rect 400 11440 438 11474
rect 224 11403 226 11419
rect 196 11395 226 11403
rect 196 11391 232 11395
rect 196 11361 204 11391
rect 216 11361 232 11391
rect 224 11314 226 11361
rect 300 11334 308 11403
rect 332 11401 342 11439
rect 400 11431 404 11440
rect 454 11425 504 11427
rect 494 11421 548 11425
rect 494 11416 514 11421
rect 504 11401 506 11416
rect 336 11389 342 11401
rect 289 11324 308 11334
rect 300 11318 308 11324
rect 332 11355 342 11389
rect 400 11393 404 11401
rect 400 11359 408 11393
rect 434 11359 438 11393
rect 498 11391 506 11401
rect 514 11391 515 11411
rect 504 11375 506 11391
rect 525 11382 528 11416
rect 547 11391 548 11411
rect 557 11391 564 11401
rect 514 11375 530 11381
rect 532 11375 548 11381
rect 332 11327 373 11355
rect 332 11321 351 11327
rect 107 11267 119 11301
rect 129 11267 149 11301
rect 196 11280 204 11314
rect 216 11280 232 11314
rect 244 11308 257 11314
rect 278 11308 291 11318
rect 244 11284 291 11308
rect 300 11308 321 11318
rect 336 11311 351 11321
rect 300 11284 329 11308
rect 332 11293 351 11311
rect 361 11321 375 11327
rect 400 11321 411 11359
rect 562 11322 612 11324
rect 361 11293 381 11321
rect 400 11293 409 11321
rect 466 11313 497 11321
rect 565 11313 596 11321
rect 442 11306 500 11313
rect 466 11305 500 11306
rect 565 11305 599 11313
rect 244 11280 257 11284
rect 42 11201 46 11235
rect 72 11201 76 11235
rect 42 11154 76 11158
rect 42 11139 46 11154
rect 72 11139 76 11154
rect 38 11121 80 11139
rect 16 11115 102 11121
rect 144 11115 148 11267
rect 174 11243 181 11271
rect 224 11233 226 11280
rect 300 11271 308 11284
rect 278 11260 305 11271
rect 332 11243 342 11293
rect 400 11273 404 11293
rect 497 11289 500 11305
rect 596 11289 599 11305
rect 466 11288 500 11289
rect 442 11281 500 11288
rect 565 11281 599 11289
rect 612 11272 614 11322
rect 256 11233 328 11241
rect 336 11235 342 11243
rect 400 11235 404 11243
rect 196 11203 204 11233
rect 216 11203 232 11233
rect 196 11199 232 11203
rect 196 11191 226 11199
rect 224 11175 226 11191
rect 332 11163 336 11231
rect 400 11201 408 11235
rect 434 11201 438 11235
rect 454 11219 504 11221
rect 504 11203 506 11219
rect 514 11213 530 11219
rect 532 11213 548 11219
rect 525 11203 548 11212
rect 400 11193 404 11201
rect 498 11193 506 11203
rect 504 11169 506 11193
rect 514 11183 515 11203
rect 525 11178 528 11203
rect 547 11183 548 11203
rect 557 11193 564 11203
rect 514 11169 548 11173
rect 400 11163 442 11164
rect 174 11153 246 11161
rect 400 11156 404 11163
rect 295 11122 300 11156
rect 324 11122 329 11156
rect 367 11139 438 11156
rect 367 11122 442 11139
rect 400 11121 442 11122
rect 378 11115 464 11121
rect 38 11099 80 11115
rect 400 11099 442 11115
rect -25 11085 25 11087
rect 42 11085 76 11099
rect 404 11085 438 11099
rect 455 11085 505 11087
rect 557 11085 607 11087
rect 16 11077 102 11085
rect 378 11077 464 11085
rect 8 11043 17 11077
rect 18 11075 51 11077
rect 80 11075 100 11077
rect 18 11043 100 11075
rect 380 11075 404 11077
rect 429 11075 438 11077
rect 442 11075 462 11077
rect 16 11035 102 11043
rect 42 11019 76 11035
rect 16 10999 38 11005
rect 42 10996 76 11000
rect 80 10999 102 11005
rect 42 10966 46 10996
rect 72 10966 76 10996
rect 42 10885 46 10919
rect 72 10885 76 10919
rect -25 10848 25 10850
rect -8 10840 14 10847
rect -8 10839 17 10840
rect 25 10839 27 10848
rect -12 10832 38 10839
rect -12 10831 34 10832
rect -12 10827 8 10831
rect 0 10815 8 10827
rect 14 10815 34 10831
rect 0 10814 34 10815
rect 0 10807 38 10814
rect 14 10806 17 10807
rect 25 10798 27 10807
rect 42 10778 45 10868
rect 69 10853 80 10885
rect 107 10853 143 10881
rect 144 10853 148 11073
rect 332 11005 336 11073
rect 380 11043 462 11075
rect 463 11043 472 11077
rect 480 11043 497 11077
rect 378 11035 464 11043
rect 505 11035 507 11085
rect 514 11043 548 11077
rect 565 11043 582 11077
rect 607 11035 609 11085
rect 404 11019 438 11035
rect 400 11005 442 11006
rect 378 10999 404 11005
rect 442 10999 464 11005
rect 400 10998 404 10999
rect 174 10959 246 10967
rect 295 10964 300 10998
rect 324 10964 329 10998
rect 224 10929 226 10945
rect 196 10921 226 10929
rect 332 10927 336 10995
rect 367 10964 438 10998
rect 400 10957 404 10964
rect 454 10951 504 10953
rect 494 10947 548 10951
rect 494 10942 514 10947
rect 504 10927 506 10942
rect 196 10917 232 10921
rect 196 10887 204 10917
rect 216 10887 232 10917
rect 400 10919 404 10927
rect 107 10847 119 10853
rect 109 10819 119 10847
rect 129 10819 149 10853
rect 174 10849 181 10879
rect 224 10840 226 10887
rect 256 10879 328 10887
rect 332 10885 336 10915
rect 400 10885 408 10919
rect 434 10885 438 10919
rect 498 10917 506 10927
rect 514 10917 515 10937
rect 504 10901 506 10917
rect 525 10908 528 10942
rect 547 10917 548 10937
rect 557 10917 564 10927
rect 514 10901 530 10907
rect 532 10901 548 10907
rect 278 10849 305 10860
rect 42 10727 46 10761
rect 72 10727 76 10761
rect 38 10689 80 10690
rect 42 10648 76 10682
rect 79 10648 113 10682
rect 42 10569 46 10603
rect 72 10569 76 10603
rect -25 10532 25 10534
rect -8 10524 14 10531
rect -8 10523 17 10524
rect 25 10523 27 10532
rect -12 10516 38 10523
rect -12 10515 34 10516
rect -12 10511 8 10515
rect 0 10499 8 10511
rect 14 10499 34 10515
rect 0 10498 34 10499
rect 0 10491 38 10498
rect 14 10490 17 10491
rect 25 10482 27 10491
rect 42 10462 45 10552
rect 71 10521 80 10549
rect 69 10483 80 10521
rect 144 10511 148 10819
rect 196 10806 204 10840
rect 216 10806 232 10840
rect 244 10836 257 10840
rect 300 10836 308 10849
rect 332 10847 342 10885
rect 400 10877 404 10885
rect 336 10837 342 10847
rect 244 10812 291 10836
rect 244 10806 257 10812
rect 224 10759 226 10806
rect 278 10802 291 10812
rect 300 10812 329 10836
rect 332 10827 342 10837
rect 400 10837 409 10865
rect 562 10848 612 10850
rect 466 10839 497 10847
rect 565 10839 596 10847
rect 300 10802 321 10812
rect 300 10796 308 10802
rect 289 10786 308 10796
rect 196 10729 204 10759
rect 216 10729 232 10759
rect 196 10725 232 10729
rect 196 10717 226 10725
rect 300 10717 308 10786
rect 332 10793 351 10827
rect 361 10799 381 10827
rect 361 10793 375 10799
rect 400 10793 411 10837
rect 442 10832 500 10839
rect 466 10831 500 10832
rect 565 10831 599 10839
rect 497 10815 500 10831
rect 596 10815 599 10831
rect 466 10814 500 10815
rect 442 10807 500 10814
rect 565 10807 599 10815
rect 612 10798 614 10848
rect 332 10769 342 10793
rect 336 10757 342 10769
rect 224 10701 226 10717
rect 332 10689 342 10757
rect 400 10761 404 10769
rect 400 10727 408 10761
rect 434 10727 438 10761
rect 454 10745 504 10747
rect 504 10729 506 10745
rect 514 10739 530 10745
rect 532 10739 548 10745
rect 525 10729 548 10738
rect 400 10719 404 10727
rect 498 10719 506 10729
rect 504 10695 506 10719
rect 514 10709 515 10729
rect 525 10704 528 10729
rect 547 10709 548 10729
rect 557 10719 564 10729
rect 514 10695 548 10699
rect 151 10648 156 10682
rect 174 10679 246 10687
rect 256 10679 328 10687
rect 336 10681 342 10689
rect 400 10684 404 10689
rect 180 10651 185 10679
rect 174 10643 246 10651
rect 256 10643 328 10651
rect 332 10649 336 10679
rect 400 10650 438 10684
rect 224 10613 226 10629
rect 196 10605 226 10613
rect 196 10601 232 10605
rect 196 10571 204 10601
rect 216 10571 232 10601
rect 224 10524 226 10571
rect 300 10544 308 10613
rect 332 10611 342 10649
rect 400 10641 404 10650
rect 454 10635 504 10637
rect 494 10631 548 10635
rect 494 10626 514 10631
rect 504 10611 506 10626
rect 336 10599 342 10611
rect 289 10534 308 10544
rect 300 10528 308 10534
rect 332 10565 342 10599
rect 400 10603 404 10611
rect 400 10569 408 10603
rect 434 10569 438 10603
rect 498 10601 506 10611
rect 514 10601 515 10621
rect 504 10585 506 10601
rect 525 10592 528 10626
rect 547 10601 548 10621
rect 557 10601 564 10611
rect 514 10585 530 10591
rect 532 10585 548 10591
rect 332 10537 373 10565
rect 332 10531 351 10537
rect 107 10477 119 10511
rect 129 10477 149 10511
rect 196 10490 204 10524
rect 216 10490 232 10524
rect 244 10518 257 10524
rect 278 10518 291 10528
rect 244 10494 291 10518
rect 300 10518 321 10528
rect 336 10521 351 10531
rect 300 10494 329 10518
rect 332 10503 351 10521
rect 361 10531 375 10537
rect 400 10531 411 10569
rect 562 10532 612 10534
rect 361 10503 381 10531
rect 400 10503 409 10531
rect 466 10523 497 10531
rect 565 10523 596 10531
rect 442 10516 500 10523
rect 466 10515 500 10516
rect 565 10515 599 10523
rect 244 10490 257 10494
rect 42 10411 46 10445
rect 72 10411 76 10445
rect 42 10364 76 10368
rect 42 10349 46 10364
rect 72 10349 76 10364
rect 38 10331 80 10349
rect 16 10325 102 10331
rect 144 10325 148 10477
rect 174 10453 181 10481
rect 224 10443 226 10490
rect 300 10481 308 10494
rect 278 10470 305 10481
rect 332 10453 342 10503
rect 400 10483 404 10503
rect 497 10499 500 10515
rect 596 10499 599 10515
rect 466 10498 500 10499
rect 442 10491 500 10498
rect 565 10491 599 10499
rect 612 10482 614 10532
rect 256 10443 328 10451
rect 336 10445 342 10453
rect 400 10445 404 10453
rect 196 10413 204 10443
rect 216 10413 232 10443
rect 196 10409 232 10413
rect 196 10401 226 10409
rect 224 10385 226 10401
rect 332 10373 336 10441
rect 400 10411 408 10445
rect 434 10411 438 10445
rect 454 10429 504 10431
rect 504 10413 506 10429
rect 514 10423 530 10429
rect 532 10423 548 10429
rect 525 10413 548 10422
rect 400 10403 404 10411
rect 498 10403 506 10413
rect 504 10379 506 10403
rect 514 10393 515 10413
rect 525 10388 528 10413
rect 547 10393 548 10413
rect 557 10403 564 10413
rect 514 10379 548 10383
rect 400 10373 442 10374
rect 174 10363 246 10371
rect 400 10366 404 10373
rect 295 10332 300 10366
rect 324 10332 329 10366
rect 367 10349 438 10366
rect 367 10332 442 10349
rect 400 10331 442 10332
rect 378 10325 464 10331
rect 38 10309 80 10325
rect 400 10309 442 10325
rect -25 10295 25 10297
rect 42 10295 76 10309
rect 404 10295 438 10309
rect 455 10295 505 10297
rect 557 10295 607 10297
rect 16 10287 102 10295
rect 378 10287 464 10295
rect 8 10253 17 10287
rect 18 10285 51 10287
rect 80 10285 100 10287
rect 18 10253 100 10285
rect 380 10285 404 10287
rect 429 10285 438 10287
rect 442 10285 462 10287
rect 16 10245 102 10253
rect 42 10229 76 10245
rect 16 10209 38 10215
rect 42 10206 76 10210
rect 80 10209 102 10215
rect 42 10176 46 10206
rect 72 10176 76 10206
rect 42 10095 46 10129
rect 72 10095 76 10129
rect -25 10058 25 10060
rect -8 10050 14 10057
rect -8 10049 17 10050
rect 25 10049 27 10058
rect -12 10042 38 10049
rect -12 10041 34 10042
rect -12 10037 8 10041
rect 0 10025 8 10037
rect 14 10025 34 10041
rect 0 10024 34 10025
rect 0 10017 38 10024
rect 14 10016 17 10017
rect 25 10008 27 10017
rect 42 9988 45 10078
rect 69 10063 80 10095
rect 107 10063 143 10091
rect 144 10063 148 10283
rect 332 10215 336 10283
rect 380 10253 462 10285
rect 463 10253 472 10287
rect 480 10253 497 10287
rect 378 10245 464 10253
rect 505 10245 507 10295
rect 514 10253 548 10287
rect 565 10253 582 10287
rect 607 10245 609 10295
rect 404 10229 438 10245
rect 400 10215 442 10216
rect 378 10209 404 10215
rect 442 10209 464 10215
rect 400 10208 404 10209
rect 174 10169 246 10177
rect 295 10174 300 10208
rect 324 10174 329 10208
rect 224 10139 226 10155
rect 196 10131 226 10139
rect 332 10137 336 10205
rect 367 10174 438 10208
rect 400 10167 404 10174
rect 454 10161 504 10163
rect 494 10157 548 10161
rect 494 10152 514 10157
rect 504 10137 506 10152
rect 196 10127 232 10131
rect 196 10097 204 10127
rect 216 10097 232 10127
rect 400 10129 404 10137
rect 107 10057 119 10063
rect 109 10029 119 10057
rect 129 10029 149 10063
rect 174 10059 181 10089
rect 224 10050 226 10097
rect 256 10089 328 10097
rect 332 10095 336 10125
rect 400 10095 408 10129
rect 434 10095 438 10129
rect 498 10127 506 10137
rect 514 10127 515 10147
rect 504 10111 506 10127
rect 525 10118 528 10152
rect 547 10127 548 10147
rect 557 10127 564 10137
rect 514 10111 530 10117
rect 532 10111 548 10117
rect 278 10059 305 10070
rect 42 9937 46 9971
rect 72 9937 76 9971
rect 38 9899 80 9900
rect 42 9858 76 9892
rect 79 9858 113 9892
rect 42 9779 46 9813
rect 72 9779 76 9813
rect -25 9742 25 9744
rect -8 9734 14 9741
rect -8 9733 17 9734
rect 25 9733 27 9742
rect -12 9726 38 9733
rect -12 9725 34 9726
rect -12 9721 8 9725
rect 0 9709 8 9721
rect 14 9709 34 9725
rect 0 9708 34 9709
rect 0 9701 38 9708
rect 14 9700 17 9701
rect 25 9692 27 9701
rect 42 9672 45 9762
rect 71 9731 80 9759
rect 69 9693 80 9731
rect 144 9721 148 10029
rect 196 10016 204 10050
rect 216 10016 232 10050
rect 244 10046 257 10050
rect 300 10046 308 10059
rect 332 10057 342 10095
rect 400 10087 404 10095
rect 336 10047 342 10057
rect 244 10022 291 10046
rect 244 10016 257 10022
rect 224 9969 226 10016
rect 278 10012 291 10022
rect 300 10022 329 10046
rect 332 10037 342 10047
rect 400 10047 409 10075
rect 562 10058 612 10060
rect 466 10049 497 10057
rect 565 10049 596 10057
rect 300 10012 321 10022
rect 300 10006 308 10012
rect 289 9996 308 10006
rect 196 9939 204 9969
rect 216 9939 232 9969
rect 196 9935 232 9939
rect 196 9927 226 9935
rect 300 9927 308 9996
rect 332 10003 351 10037
rect 361 10009 381 10037
rect 361 10003 375 10009
rect 400 10003 411 10047
rect 442 10042 500 10049
rect 466 10041 500 10042
rect 565 10041 599 10049
rect 497 10025 500 10041
rect 596 10025 599 10041
rect 466 10024 500 10025
rect 442 10017 500 10024
rect 565 10017 599 10025
rect 612 10008 614 10058
rect 332 9979 342 10003
rect 336 9967 342 9979
rect 224 9911 226 9927
rect 332 9899 342 9967
rect 400 9971 404 9979
rect 400 9937 408 9971
rect 434 9937 438 9971
rect 454 9955 504 9957
rect 504 9939 506 9955
rect 514 9949 530 9955
rect 532 9949 548 9955
rect 525 9939 548 9948
rect 400 9929 404 9937
rect 498 9929 506 9939
rect 504 9905 506 9929
rect 514 9919 515 9939
rect 525 9914 528 9939
rect 547 9919 548 9939
rect 557 9929 564 9939
rect 514 9905 548 9909
rect 151 9858 156 9892
rect 174 9889 246 9897
rect 256 9889 328 9897
rect 336 9891 342 9899
rect 400 9894 404 9899
rect 180 9861 185 9889
rect 174 9853 246 9861
rect 256 9853 328 9861
rect 332 9859 336 9889
rect 400 9860 438 9894
rect 224 9823 226 9839
rect 196 9815 226 9823
rect 196 9811 232 9815
rect 196 9781 204 9811
rect 216 9781 232 9811
rect 224 9734 226 9781
rect 300 9754 308 9823
rect 332 9821 342 9859
rect 400 9851 404 9860
rect 454 9845 504 9847
rect 494 9841 548 9845
rect 494 9836 514 9841
rect 504 9821 506 9836
rect 336 9809 342 9821
rect 289 9744 308 9754
rect 300 9738 308 9744
rect 332 9775 342 9809
rect 400 9813 404 9821
rect 400 9779 408 9813
rect 434 9779 438 9813
rect 498 9811 506 9821
rect 514 9811 515 9831
rect 504 9795 506 9811
rect 525 9802 528 9836
rect 547 9811 548 9831
rect 557 9811 564 9821
rect 514 9795 530 9801
rect 532 9795 548 9801
rect 332 9747 373 9775
rect 332 9741 351 9747
rect 107 9687 119 9721
rect 129 9687 149 9721
rect 196 9700 204 9734
rect 216 9700 232 9734
rect 244 9728 257 9734
rect 278 9728 291 9738
rect 244 9704 291 9728
rect 300 9728 321 9738
rect 336 9731 351 9741
rect 300 9704 329 9728
rect 332 9713 351 9731
rect 361 9741 375 9747
rect 400 9741 411 9779
rect 562 9742 612 9744
rect 361 9713 381 9741
rect 400 9713 409 9741
rect 466 9733 497 9741
rect 565 9733 596 9741
rect 442 9726 500 9733
rect 466 9725 500 9726
rect 565 9725 599 9733
rect 244 9700 257 9704
rect 42 9621 46 9655
rect 72 9621 76 9655
rect 42 9574 76 9578
rect 42 9559 46 9574
rect 72 9559 76 9574
rect 38 9541 80 9559
rect 16 9535 102 9541
rect 144 9535 148 9687
rect 174 9663 181 9691
rect 224 9653 226 9700
rect 300 9691 308 9704
rect 278 9680 305 9691
rect 332 9663 342 9713
rect 400 9693 404 9713
rect 497 9709 500 9725
rect 596 9709 599 9725
rect 466 9708 500 9709
rect 442 9701 500 9708
rect 565 9701 599 9709
rect 612 9692 614 9742
rect 256 9653 328 9661
rect 336 9655 342 9663
rect 400 9655 404 9663
rect 196 9623 204 9653
rect 216 9623 232 9653
rect 196 9619 232 9623
rect 196 9611 226 9619
rect 224 9595 226 9611
rect 332 9583 336 9651
rect 400 9621 408 9655
rect 434 9621 438 9655
rect 454 9639 504 9641
rect 504 9623 506 9639
rect 514 9633 530 9639
rect 532 9633 548 9639
rect 525 9623 548 9632
rect 400 9613 404 9621
rect 498 9613 506 9623
rect 504 9589 506 9613
rect 514 9603 515 9623
rect 525 9598 528 9623
rect 547 9603 548 9623
rect 557 9613 564 9623
rect 514 9589 548 9593
rect 400 9583 442 9584
rect 174 9573 246 9581
rect 400 9576 404 9583
rect 295 9542 300 9576
rect 324 9542 329 9576
rect 367 9559 438 9576
rect 367 9542 442 9559
rect 400 9541 442 9542
rect 378 9535 464 9541
rect 38 9519 80 9535
rect 400 9519 442 9535
rect -25 9505 25 9507
rect 42 9505 76 9519
rect 404 9505 438 9519
rect 455 9505 505 9507
rect 557 9505 607 9507
rect 16 9497 102 9505
rect 378 9497 464 9505
rect 8 9463 17 9497
rect 18 9495 51 9497
rect 80 9495 100 9497
rect 18 9463 100 9495
rect 380 9495 404 9497
rect 429 9495 438 9497
rect 442 9495 462 9497
rect 16 9455 102 9463
rect 42 9439 76 9455
rect 16 9419 38 9425
rect 42 9416 76 9420
rect 80 9419 102 9425
rect 42 9386 46 9416
rect 72 9386 76 9416
rect 42 9305 46 9339
rect 72 9305 76 9339
rect -25 9268 25 9270
rect -8 9260 14 9267
rect -8 9259 17 9260
rect 25 9259 27 9268
rect -12 9252 38 9259
rect -12 9251 34 9252
rect -12 9247 8 9251
rect 0 9235 8 9247
rect 14 9235 34 9251
rect 0 9234 34 9235
rect 0 9227 38 9234
rect 14 9226 17 9227
rect 25 9218 27 9227
rect 42 9198 45 9288
rect 69 9273 80 9305
rect 107 9273 143 9301
rect 144 9273 148 9493
rect 332 9425 336 9493
rect 380 9463 462 9495
rect 463 9463 472 9497
rect 480 9463 497 9497
rect 378 9455 464 9463
rect 505 9455 507 9505
rect 514 9463 548 9497
rect 565 9463 582 9497
rect 607 9455 609 9505
rect 404 9439 438 9455
rect 400 9425 442 9426
rect 378 9419 404 9425
rect 442 9419 464 9425
rect 400 9418 404 9419
rect 174 9379 246 9387
rect 295 9384 300 9418
rect 324 9384 329 9418
rect 224 9349 226 9365
rect 196 9341 226 9349
rect 332 9347 336 9415
rect 367 9384 438 9418
rect 400 9377 404 9384
rect 454 9371 504 9373
rect 494 9367 548 9371
rect 494 9362 514 9367
rect 504 9347 506 9362
rect 196 9337 232 9341
rect 196 9307 204 9337
rect 216 9307 232 9337
rect 400 9339 404 9347
rect 107 9267 119 9273
rect 109 9239 119 9267
rect 129 9239 149 9273
rect 174 9269 181 9299
rect 224 9260 226 9307
rect 256 9299 328 9307
rect 332 9305 336 9335
rect 400 9305 408 9339
rect 434 9305 438 9339
rect 498 9337 506 9347
rect 514 9337 515 9357
rect 504 9321 506 9337
rect 525 9328 528 9362
rect 547 9337 548 9357
rect 557 9337 564 9347
rect 514 9321 530 9327
rect 532 9321 548 9327
rect 278 9269 305 9280
rect 42 9147 46 9181
rect 72 9147 76 9181
rect 38 9109 80 9110
rect 42 9068 76 9102
rect 79 9068 113 9102
rect 42 8989 46 9023
rect 72 8989 76 9023
rect -25 8952 25 8954
rect -8 8944 14 8951
rect -8 8943 17 8944
rect 25 8943 27 8952
rect -12 8936 38 8943
rect -12 8935 34 8936
rect -12 8931 8 8935
rect 0 8919 8 8931
rect 14 8919 34 8935
rect 0 8918 34 8919
rect 0 8911 38 8918
rect 14 8910 17 8911
rect 25 8902 27 8911
rect 42 8882 45 8972
rect 71 8941 80 8969
rect 69 8903 80 8941
rect 144 8931 148 9239
rect 196 9226 204 9260
rect 216 9226 232 9260
rect 244 9256 257 9260
rect 300 9256 308 9269
rect 332 9267 342 9305
rect 400 9297 404 9305
rect 336 9257 342 9267
rect 244 9232 291 9256
rect 244 9226 257 9232
rect 224 9179 226 9226
rect 278 9222 291 9232
rect 300 9232 329 9256
rect 332 9247 342 9257
rect 400 9257 409 9285
rect 562 9268 612 9270
rect 466 9259 497 9267
rect 565 9259 596 9267
rect 300 9222 321 9232
rect 300 9216 308 9222
rect 289 9206 308 9216
rect 196 9149 204 9179
rect 216 9149 232 9179
rect 196 9145 232 9149
rect 196 9137 226 9145
rect 300 9137 308 9206
rect 332 9213 351 9247
rect 361 9219 381 9247
rect 361 9213 375 9219
rect 400 9213 411 9257
rect 442 9252 500 9259
rect 466 9251 500 9252
rect 565 9251 599 9259
rect 497 9235 500 9251
rect 596 9235 599 9251
rect 466 9234 500 9235
rect 442 9227 500 9234
rect 565 9227 599 9235
rect 612 9218 614 9268
rect 332 9189 342 9213
rect 336 9177 342 9189
rect 224 9121 226 9137
rect 332 9109 342 9177
rect 400 9181 404 9189
rect 400 9147 408 9181
rect 434 9147 438 9181
rect 454 9165 504 9167
rect 504 9149 506 9165
rect 514 9159 530 9165
rect 532 9159 548 9165
rect 525 9149 548 9158
rect 400 9139 404 9147
rect 498 9139 506 9149
rect 504 9115 506 9139
rect 514 9129 515 9149
rect 525 9124 528 9149
rect 547 9129 548 9149
rect 557 9139 564 9149
rect 514 9115 548 9119
rect 151 9068 156 9102
rect 174 9099 246 9107
rect 256 9099 328 9107
rect 336 9101 342 9109
rect 400 9104 404 9109
rect 180 9071 185 9099
rect 174 9063 246 9071
rect 256 9063 328 9071
rect 332 9069 336 9099
rect 400 9070 438 9104
rect 224 9033 226 9049
rect 196 9025 226 9033
rect 196 9021 232 9025
rect 196 8991 204 9021
rect 216 8991 232 9021
rect 224 8944 226 8991
rect 300 8964 308 9033
rect 332 9031 342 9069
rect 400 9061 404 9070
rect 454 9055 504 9057
rect 494 9051 548 9055
rect 494 9046 514 9051
rect 504 9031 506 9046
rect 336 9019 342 9031
rect 289 8954 308 8964
rect 300 8948 308 8954
rect 332 8985 342 9019
rect 400 9023 404 9031
rect 400 8989 408 9023
rect 434 8989 438 9023
rect 498 9021 506 9031
rect 514 9021 515 9041
rect 504 9005 506 9021
rect 525 9012 528 9046
rect 547 9021 548 9041
rect 557 9021 564 9031
rect 514 9005 530 9011
rect 532 9005 548 9011
rect 332 8957 373 8985
rect 332 8951 351 8957
rect 107 8897 119 8931
rect 129 8897 149 8931
rect 196 8910 204 8944
rect 216 8910 232 8944
rect 244 8938 257 8944
rect 278 8938 291 8948
rect 244 8914 291 8938
rect 300 8938 321 8948
rect 336 8941 351 8951
rect 300 8914 329 8938
rect 332 8923 351 8941
rect 361 8951 375 8957
rect 400 8951 411 8989
rect 562 8952 612 8954
rect 361 8923 381 8951
rect 400 8923 409 8951
rect 466 8943 497 8951
rect 565 8943 596 8951
rect 442 8936 500 8943
rect 466 8935 500 8936
rect 565 8935 599 8943
rect 244 8910 257 8914
rect 42 8831 46 8865
rect 72 8831 76 8865
rect 42 8784 76 8788
rect 42 8769 46 8784
rect 72 8769 76 8784
rect 38 8751 80 8769
rect 16 8745 102 8751
rect 144 8745 148 8897
rect 174 8873 181 8901
rect 224 8863 226 8910
rect 300 8901 308 8914
rect 278 8890 305 8901
rect 332 8873 342 8923
rect 400 8903 404 8923
rect 497 8919 500 8935
rect 596 8919 599 8935
rect 466 8918 500 8919
rect 442 8911 500 8918
rect 565 8911 599 8919
rect 612 8902 614 8952
rect 256 8863 328 8871
rect 336 8865 342 8873
rect 400 8865 404 8873
rect 196 8833 204 8863
rect 216 8833 232 8863
rect 196 8829 232 8833
rect 196 8821 226 8829
rect 224 8805 226 8821
rect 332 8793 336 8861
rect 400 8831 408 8865
rect 434 8831 438 8865
rect 454 8849 504 8851
rect 504 8833 506 8849
rect 514 8843 530 8849
rect 532 8843 548 8849
rect 525 8833 548 8842
rect 400 8823 404 8831
rect 498 8823 506 8833
rect 504 8799 506 8823
rect 514 8813 515 8833
rect 525 8808 528 8833
rect 547 8813 548 8833
rect 557 8823 564 8833
rect 514 8799 548 8803
rect 400 8793 442 8794
rect 174 8783 246 8791
rect 400 8786 404 8793
rect 295 8752 300 8786
rect 324 8752 329 8786
rect 367 8769 438 8786
rect 367 8752 442 8769
rect 400 8751 442 8752
rect 378 8745 464 8751
rect 38 8729 80 8745
rect 400 8729 442 8745
rect -25 8715 25 8717
rect 42 8715 76 8729
rect 404 8715 438 8729
rect 455 8715 505 8717
rect 557 8715 607 8717
rect 16 8707 102 8715
rect 378 8707 464 8715
rect 8 8673 17 8707
rect 18 8705 51 8707
rect 80 8705 100 8707
rect 18 8673 100 8705
rect 380 8705 404 8707
rect 429 8705 438 8707
rect 442 8705 462 8707
rect 16 8665 102 8673
rect 42 8649 76 8665
rect 16 8629 38 8635
rect 42 8626 76 8630
rect 80 8629 102 8635
rect 42 8596 46 8626
rect 72 8596 76 8626
rect 42 8515 46 8549
rect 72 8515 76 8549
rect -25 8478 25 8480
rect -8 8470 14 8477
rect -8 8469 17 8470
rect 25 8469 27 8478
rect -12 8462 38 8469
rect -12 8461 34 8462
rect -12 8457 8 8461
rect 0 8445 8 8457
rect 14 8445 34 8461
rect 0 8444 34 8445
rect 0 8437 38 8444
rect 14 8436 17 8437
rect 25 8428 27 8437
rect 42 8408 45 8498
rect 69 8483 80 8515
rect 107 8483 143 8511
rect 144 8483 148 8703
rect 332 8635 336 8703
rect 380 8673 462 8705
rect 463 8673 472 8707
rect 480 8673 497 8707
rect 378 8665 464 8673
rect 505 8665 507 8715
rect 514 8673 548 8707
rect 565 8673 582 8707
rect 607 8665 609 8715
rect 404 8649 438 8665
rect 400 8635 442 8636
rect 378 8629 404 8635
rect 442 8629 464 8635
rect 400 8628 404 8629
rect 174 8589 246 8597
rect 295 8594 300 8628
rect 324 8594 329 8628
rect 224 8559 226 8575
rect 196 8551 226 8559
rect 332 8557 336 8625
rect 367 8594 438 8628
rect 400 8587 404 8594
rect 454 8581 504 8583
rect 494 8577 548 8581
rect 494 8572 514 8577
rect 504 8557 506 8572
rect 196 8547 232 8551
rect 196 8517 204 8547
rect 216 8517 232 8547
rect 400 8549 404 8557
rect 107 8477 119 8483
rect 109 8449 119 8477
rect 129 8449 149 8483
rect 174 8479 181 8509
rect 224 8470 226 8517
rect 256 8509 328 8517
rect 332 8515 336 8545
rect 400 8515 408 8549
rect 434 8515 438 8549
rect 498 8547 506 8557
rect 514 8547 515 8567
rect 504 8531 506 8547
rect 525 8538 528 8572
rect 547 8547 548 8567
rect 557 8547 564 8557
rect 514 8531 530 8537
rect 532 8531 548 8537
rect 278 8479 305 8490
rect 42 8357 46 8391
rect 72 8357 76 8391
rect 38 8319 80 8320
rect 42 8278 76 8312
rect 79 8278 113 8312
rect 42 8199 46 8233
rect 72 8199 76 8233
rect -25 8162 25 8164
rect -8 8154 14 8161
rect -8 8153 17 8154
rect 25 8153 27 8162
rect -12 8146 38 8153
rect -12 8145 34 8146
rect -12 8141 8 8145
rect 0 8129 8 8141
rect 14 8129 34 8145
rect 0 8128 34 8129
rect 0 8121 38 8128
rect 14 8120 17 8121
rect 25 8112 27 8121
rect 42 8092 45 8182
rect 71 8151 80 8179
rect 69 8113 80 8151
rect 144 8141 148 8449
rect 196 8436 204 8470
rect 216 8436 232 8470
rect 244 8466 257 8470
rect 300 8466 308 8479
rect 332 8477 342 8515
rect 400 8507 404 8515
rect 336 8467 342 8477
rect 244 8442 291 8466
rect 244 8436 257 8442
rect 224 8389 226 8436
rect 278 8432 291 8442
rect 300 8442 329 8466
rect 332 8457 342 8467
rect 400 8467 409 8495
rect 562 8478 612 8480
rect 466 8469 497 8477
rect 565 8469 596 8477
rect 300 8432 321 8442
rect 300 8426 308 8432
rect 289 8416 308 8426
rect 196 8359 204 8389
rect 216 8359 232 8389
rect 196 8355 232 8359
rect 196 8347 226 8355
rect 300 8347 308 8416
rect 332 8423 351 8457
rect 361 8429 381 8457
rect 361 8423 375 8429
rect 400 8423 411 8467
rect 442 8462 500 8469
rect 466 8461 500 8462
rect 565 8461 599 8469
rect 497 8445 500 8461
rect 596 8445 599 8461
rect 466 8444 500 8445
rect 442 8437 500 8444
rect 565 8437 599 8445
rect 612 8428 614 8478
rect 332 8399 342 8423
rect 336 8387 342 8399
rect 224 8331 226 8347
rect 332 8319 342 8387
rect 400 8391 404 8399
rect 400 8357 408 8391
rect 434 8357 438 8391
rect 454 8375 504 8377
rect 504 8359 506 8375
rect 514 8369 530 8375
rect 532 8369 548 8375
rect 525 8359 548 8368
rect 400 8349 404 8357
rect 498 8349 506 8359
rect 504 8325 506 8349
rect 514 8339 515 8359
rect 525 8334 528 8359
rect 547 8339 548 8359
rect 557 8349 564 8359
rect 514 8325 548 8329
rect 151 8278 156 8312
rect 174 8309 246 8317
rect 256 8309 328 8317
rect 336 8311 342 8319
rect 400 8314 404 8319
rect 180 8281 185 8309
rect 174 8273 246 8281
rect 256 8273 328 8281
rect 332 8279 336 8309
rect 400 8280 438 8314
rect 224 8243 226 8259
rect 196 8235 226 8243
rect 196 8231 232 8235
rect 196 8201 204 8231
rect 216 8201 232 8231
rect 224 8154 226 8201
rect 300 8174 308 8243
rect 332 8241 342 8279
rect 400 8271 404 8280
rect 454 8265 504 8267
rect 494 8261 548 8265
rect 494 8256 514 8261
rect 504 8241 506 8256
rect 336 8229 342 8241
rect 289 8164 308 8174
rect 300 8158 308 8164
rect 332 8195 342 8229
rect 400 8233 404 8241
rect 400 8199 408 8233
rect 434 8199 438 8233
rect 498 8231 506 8241
rect 514 8231 515 8251
rect 504 8215 506 8231
rect 525 8222 528 8256
rect 547 8231 548 8251
rect 557 8231 564 8241
rect 514 8215 530 8221
rect 532 8215 548 8221
rect 332 8167 373 8195
rect 332 8161 351 8167
rect 107 8107 119 8141
rect 129 8107 149 8141
rect 196 8120 204 8154
rect 216 8120 232 8154
rect 244 8148 257 8154
rect 278 8148 291 8158
rect 244 8124 291 8148
rect 300 8148 321 8158
rect 336 8151 351 8161
rect 300 8124 329 8148
rect 332 8133 351 8151
rect 361 8161 375 8167
rect 400 8161 411 8199
rect 562 8162 612 8164
rect 361 8133 381 8161
rect 400 8133 409 8161
rect 466 8153 497 8161
rect 565 8153 596 8161
rect 442 8146 500 8153
rect 466 8145 500 8146
rect 565 8145 599 8153
rect 244 8120 257 8124
rect 42 8041 46 8075
rect 72 8041 76 8075
rect 42 7994 76 7998
rect 42 7979 46 7994
rect 72 7979 76 7994
rect 38 7961 80 7979
rect 16 7955 102 7961
rect 144 7955 148 8107
rect 174 8083 181 8111
rect 224 8073 226 8120
rect 300 8111 308 8124
rect 278 8100 305 8111
rect 332 8083 342 8133
rect 400 8113 404 8133
rect 497 8129 500 8145
rect 596 8129 599 8145
rect 466 8128 500 8129
rect 442 8121 500 8128
rect 565 8121 599 8129
rect 612 8112 614 8162
rect 256 8073 328 8081
rect 336 8075 342 8083
rect 400 8075 404 8083
rect 196 8043 204 8073
rect 216 8043 232 8073
rect 196 8039 232 8043
rect 196 8031 226 8039
rect 224 8015 226 8031
rect 332 8003 336 8071
rect 400 8041 408 8075
rect 434 8041 438 8075
rect 454 8059 504 8061
rect 504 8043 506 8059
rect 514 8053 530 8059
rect 532 8053 548 8059
rect 525 8043 548 8052
rect 400 8033 404 8041
rect 498 8033 506 8043
rect 504 8009 506 8033
rect 514 8023 515 8043
rect 525 8018 528 8043
rect 547 8023 548 8043
rect 557 8033 564 8043
rect 514 8009 548 8013
rect 400 8003 442 8004
rect 174 7993 246 8001
rect 400 7996 404 8003
rect 295 7962 300 7996
rect 324 7962 329 7996
rect 367 7979 438 7996
rect 367 7962 442 7979
rect 400 7961 442 7962
rect 378 7955 464 7961
rect 38 7939 80 7955
rect 400 7939 442 7955
rect -25 7925 25 7927
rect 42 7925 76 7939
rect 404 7925 438 7939
rect 455 7925 505 7927
rect 557 7925 607 7927
rect 16 7917 102 7925
rect 378 7917 464 7925
rect 8 7883 17 7917
rect 18 7915 51 7917
rect 80 7915 100 7917
rect 18 7883 100 7915
rect 380 7915 404 7917
rect 429 7915 438 7917
rect 442 7915 462 7917
rect 16 7875 102 7883
rect 42 7859 76 7875
rect 16 7839 38 7845
rect 42 7836 76 7840
rect 80 7839 102 7845
rect 42 7806 46 7836
rect 72 7806 76 7836
rect 42 7725 46 7759
rect 72 7725 76 7759
rect -25 7688 25 7690
rect -8 7680 14 7687
rect -8 7679 17 7680
rect 25 7679 27 7688
rect -12 7672 38 7679
rect -12 7671 34 7672
rect -12 7667 8 7671
rect 0 7655 8 7667
rect 14 7655 34 7671
rect 0 7654 34 7655
rect 0 7647 38 7654
rect 14 7646 17 7647
rect 25 7638 27 7647
rect 42 7618 45 7708
rect 69 7693 80 7725
rect 107 7693 143 7721
rect 144 7693 148 7913
rect 332 7845 336 7913
rect 380 7883 462 7915
rect 463 7883 472 7917
rect 480 7883 497 7917
rect 378 7875 464 7883
rect 505 7875 507 7925
rect 514 7883 548 7917
rect 565 7883 582 7917
rect 607 7875 609 7925
rect 404 7859 438 7875
rect 400 7845 442 7846
rect 378 7839 404 7845
rect 442 7839 464 7845
rect 400 7838 404 7839
rect 174 7799 246 7807
rect 295 7804 300 7838
rect 324 7804 329 7838
rect 224 7769 226 7785
rect 196 7761 226 7769
rect 332 7767 336 7835
rect 367 7804 438 7838
rect 400 7797 404 7804
rect 454 7791 504 7793
rect 494 7787 548 7791
rect 494 7782 514 7787
rect 504 7767 506 7782
rect 196 7757 232 7761
rect 196 7727 204 7757
rect 216 7727 232 7757
rect 400 7759 404 7767
rect 107 7687 119 7693
rect 109 7659 119 7687
rect 129 7659 149 7693
rect 174 7689 181 7719
rect 224 7680 226 7727
rect 256 7719 328 7727
rect 332 7725 336 7755
rect 400 7725 408 7759
rect 434 7725 438 7759
rect 498 7757 506 7767
rect 514 7757 515 7777
rect 504 7741 506 7757
rect 525 7748 528 7782
rect 547 7757 548 7777
rect 557 7757 564 7767
rect 514 7741 530 7747
rect 532 7741 548 7747
rect 278 7689 305 7700
rect 42 7567 46 7601
rect 72 7567 76 7601
rect 38 7529 80 7530
rect 42 7488 76 7522
rect 79 7488 113 7522
rect 42 7409 46 7443
rect 72 7409 76 7443
rect -25 7372 25 7374
rect -8 7364 14 7371
rect -8 7363 17 7364
rect 25 7363 27 7372
rect -12 7356 38 7363
rect -12 7355 34 7356
rect -12 7351 8 7355
rect 0 7339 8 7351
rect 14 7339 34 7355
rect 0 7338 34 7339
rect 0 7331 38 7338
rect 14 7330 17 7331
rect 25 7322 27 7331
rect 42 7302 45 7392
rect 71 7361 80 7389
rect 69 7323 80 7361
rect 144 7351 148 7659
rect 196 7646 204 7680
rect 216 7646 232 7680
rect 244 7676 257 7680
rect 300 7676 308 7689
rect 332 7687 342 7725
rect 400 7717 404 7725
rect 336 7677 342 7687
rect 244 7652 291 7676
rect 244 7646 257 7652
rect 224 7599 226 7646
rect 278 7642 291 7652
rect 300 7652 329 7676
rect 332 7667 342 7677
rect 400 7677 409 7705
rect 562 7688 612 7690
rect 466 7679 497 7687
rect 565 7679 596 7687
rect 300 7642 321 7652
rect 300 7636 308 7642
rect 289 7626 308 7636
rect 196 7569 204 7599
rect 216 7569 232 7599
rect 196 7565 232 7569
rect 196 7557 226 7565
rect 300 7557 308 7626
rect 332 7633 351 7667
rect 361 7639 381 7667
rect 361 7633 375 7639
rect 400 7633 411 7677
rect 442 7672 500 7679
rect 466 7671 500 7672
rect 565 7671 599 7679
rect 497 7655 500 7671
rect 596 7655 599 7671
rect 466 7654 500 7655
rect 442 7647 500 7654
rect 565 7647 599 7655
rect 612 7638 614 7688
rect 332 7609 342 7633
rect 336 7597 342 7609
rect 224 7541 226 7557
rect 332 7529 342 7597
rect 400 7601 404 7609
rect 400 7567 408 7601
rect 434 7567 438 7601
rect 454 7585 504 7587
rect 504 7569 506 7585
rect 514 7579 530 7585
rect 532 7579 548 7585
rect 525 7569 548 7578
rect 400 7559 404 7567
rect 498 7559 506 7569
rect 504 7535 506 7559
rect 514 7549 515 7569
rect 525 7544 528 7569
rect 547 7549 548 7569
rect 557 7559 564 7569
rect 514 7535 548 7539
rect 151 7488 156 7522
rect 174 7519 246 7527
rect 256 7519 328 7527
rect 336 7521 342 7529
rect 400 7524 404 7529
rect 180 7491 185 7519
rect 174 7483 246 7491
rect 256 7483 328 7491
rect 332 7489 336 7519
rect 400 7490 438 7524
rect 224 7453 226 7469
rect 196 7445 226 7453
rect 196 7441 232 7445
rect 196 7411 204 7441
rect 216 7411 232 7441
rect 224 7364 226 7411
rect 300 7384 308 7453
rect 332 7451 342 7489
rect 400 7481 404 7490
rect 454 7475 504 7477
rect 494 7471 548 7475
rect 494 7466 514 7471
rect 504 7451 506 7466
rect 336 7439 342 7451
rect 289 7374 308 7384
rect 300 7368 308 7374
rect 332 7405 342 7439
rect 400 7443 404 7451
rect 400 7409 408 7443
rect 434 7409 438 7443
rect 498 7441 506 7451
rect 514 7441 515 7461
rect 504 7425 506 7441
rect 525 7432 528 7466
rect 547 7441 548 7461
rect 557 7441 564 7451
rect 514 7425 530 7431
rect 532 7425 548 7431
rect 332 7377 373 7405
rect 332 7371 351 7377
rect 107 7317 119 7351
rect 129 7317 149 7351
rect 196 7330 204 7364
rect 216 7330 232 7364
rect 244 7358 257 7364
rect 278 7358 291 7368
rect 244 7334 291 7358
rect 300 7358 321 7368
rect 336 7361 351 7371
rect 300 7334 329 7358
rect 332 7343 351 7361
rect 361 7371 375 7377
rect 400 7371 411 7409
rect 562 7372 612 7374
rect 361 7343 381 7371
rect 400 7343 409 7371
rect 466 7363 497 7371
rect 565 7363 596 7371
rect 442 7356 500 7363
rect 466 7355 500 7356
rect 565 7355 599 7363
rect 244 7330 257 7334
rect 42 7251 46 7285
rect 72 7251 76 7285
rect 42 7204 76 7208
rect 42 7189 46 7204
rect 72 7189 76 7204
rect 38 7171 80 7189
rect 16 7165 102 7171
rect 144 7165 148 7317
rect 174 7293 181 7321
rect 224 7283 226 7330
rect 300 7321 308 7334
rect 278 7310 305 7321
rect 332 7293 342 7343
rect 400 7323 404 7343
rect 497 7339 500 7355
rect 596 7339 599 7355
rect 466 7338 500 7339
rect 442 7331 500 7338
rect 565 7331 599 7339
rect 612 7322 614 7372
rect 256 7283 328 7291
rect 336 7285 342 7293
rect 400 7285 404 7293
rect 196 7253 204 7283
rect 216 7253 232 7283
rect 196 7249 232 7253
rect 196 7241 226 7249
rect 224 7225 226 7241
rect 332 7213 336 7281
rect 400 7251 408 7285
rect 434 7251 438 7285
rect 454 7269 504 7271
rect 504 7253 506 7269
rect 514 7263 530 7269
rect 532 7263 548 7269
rect 525 7253 548 7262
rect 400 7243 404 7251
rect 498 7243 506 7253
rect 504 7219 506 7243
rect 514 7233 515 7253
rect 525 7228 528 7253
rect 547 7233 548 7253
rect 557 7243 564 7253
rect 514 7219 548 7223
rect 400 7213 442 7214
rect 174 7203 246 7211
rect 400 7206 404 7213
rect 295 7172 300 7206
rect 324 7172 329 7206
rect 367 7189 438 7206
rect 367 7172 442 7189
rect 400 7171 442 7172
rect 378 7165 464 7171
rect 38 7149 80 7165
rect 400 7149 442 7165
rect -25 7135 25 7137
rect 42 7135 76 7149
rect 404 7135 438 7149
rect 455 7135 505 7137
rect 557 7135 607 7137
rect 16 7127 102 7135
rect 378 7127 464 7135
rect 8 7093 17 7127
rect 18 7125 51 7127
rect 80 7125 100 7127
rect 18 7093 100 7125
rect 380 7125 404 7127
rect 429 7125 438 7127
rect 442 7125 462 7127
rect 16 7085 102 7093
rect 42 7069 76 7085
rect 16 7049 38 7055
rect 42 7046 76 7050
rect 80 7049 102 7055
rect 42 7016 46 7046
rect 72 7016 76 7046
rect 42 6935 46 6969
rect 72 6935 76 6969
rect -25 6898 25 6900
rect -8 6890 14 6897
rect -8 6889 17 6890
rect 25 6889 27 6898
rect -12 6882 38 6889
rect -12 6881 34 6882
rect -12 6877 8 6881
rect 0 6865 8 6877
rect 14 6865 34 6881
rect 0 6864 34 6865
rect 0 6857 38 6864
rect 14 6856 17 6857
rect 25 6848 27 6857
rect 42 6828 45 6918
rect 69 6903 80 6935
rect 107 6903 143 6931
rect 144 6903 148 7123
rect 332 7055 336 7123
rect 380 7093 462 7125
rect 463 7093 472 7127
rect 480 7093 497 7127
rect 378 7085 464 7093
rect 505 7085 507 7135
rect 514 7093 548 7127
rect 565 7093 582 7127
rect 607 7085 609 7135
rect 404 7069 438 7085
rect 400 7055 442 7056
rect 378 7049 404 7055
rect 442 7049 464 7055
rect 400 7048 404 7049
rect 174 7009 246 7017
rect 295 7014 300 7048
rect 324 7014 329 7048
rect 224 6979 226 6995
rect 196 6971 226 6979
rect 332 6977 336 7045
rect 367 7014 438 7048
rect 400 7007 404 7014
rect 454 7001 504 7003
rect 494 6997 548 7001
rect 494 6992 514 6997
rect 504 6977 506 6992
rect 196 6967 232 6971
rect 196 6937 204 6967
rect 216 6937 232 6967
rect 400 6969 404 6977
rect 107 6897 119 6903
rect 109 6869 119 6897
rect 129 6869 149 6903
rect 174 6899 181 6929
rect 224 6890 226 6937
rect 256 6929 328 6937
rect 332 6935 336 6965
rect 400 6935 408 6969
rect 434 6935 438 6969
rect 498 6967 506 6977
rect 514 6967 515 6987
rect 504 6951 506 6967
rect 525 6958 528 6992
rect 547 6967 548 6987
rect 557 6967 564 6977
rect 514 6951 530 6957
rect 532 6951 548 6957
rect 278 6899 305 6910
rect 42 6777 46 6811
rect 72 6777 76 6811
rect 38 6739 80 6740
rect 42 6698 76 6732
rect 79 6698 113 6732
rect 42 6619 46 6653
rect 72 6619 76 6653
rect -25 6582 25 6584
rect -8 6574 14 6581
rect -8 6573 17 6574
rect 25 6573 27 6582
rect -12 6566 38 6573
rect -12 6565 34 6566
rect -12 6561 8 6565
rect 0 6549 8 6561
rect 14 6549 34 6565
rect 0 6548 34 6549
rect 0 6541 38 6548
rect 14 6540 17 6541
rect 25 6532 27 6541
rect 42 6512 45 6602
rect 71 6571 80 6599
rect 69 6533 80 6571
rect 144 6561 148 6869
rect 196 6856 204 6890
rect 216 6856 232 6890
rect 244 6886 257 6890
rect 300 6886 308 6899
rect 332 6897 342 6935
rect 400 6927 404 6935
rect 336 6887 342 6897
rect 244 6862 291 6886
rect 244 6856 257 6862
rect 224 6809 226 6856
rect 278 6852 291 6862
rect 300 6862 329 6886
rect 332 6877 342 6887
rect 400 6887 409 6915
rect 562 6898 612 6900
rect 466 6889 497 6897
rect 565 6889 596 6897
rect 300 6852 321 6862
rect 300 6846 308 6852
rect 289 6836 308 6846
rect 196 6779 204 6809
rect 216 6779 232 6809
rect 196 6775 232 6779
rect 196 6767 226 6775
rect 300 6767 308 6836
rect 332 6843 351 6877
rect 361 6849 381 6877
rect 361 6843 375 6849
rect 400 6843 411 6887
rect 442 6882 500 6889
rect 466 6881 500 6882
rect 565 6881 599 6889
rect 497 6865 500 6881
rect 596 6865 599 6881
rect 466 6864 500 6865
rect 442 6857 500 6864
rect 565 6857 599 6865
rect 612 6848 614 6898
rect 332 6819 342 6843
rect 336 6807 342 6819
rect 224 6751 226 6767
rect 332 6739 342 6807
rect 400 6811 404 6819
rect 400 6777 408 6811
rect 434 6777 438 6811
rect 454 6795 504 6797
rect 504 6779 506 6795
rect 514 6789 530 6795
rect 532 6789 548 6795
rect 525 6779 548 6788
rect 400 6769 404 6777
rect 498 6769 506 6779
rect 504 6745 506 6769
rect 514 6759 515 6779
rect 525 6754 528 6779
rect 547 6759 548 6779
rect 557 6769 564 6779
rect 514 6745 548 6749
rect 151 6698 156 6732
rect 174 6729 246 6737
rect 256 6729 328 6737
rect 336 6731 342 6739
rect 400 6734 404 6739
rect 180 6701 185 6729
rect 174 6693 246 6701
rect 256 6693 328 6701
rect 332 6699 336 6729
rect 400 6700 438 6734
rect 224 6663 226 6679
rect 196 6655 226 6663
rect 196 6651 232 6655
rect 196 6621 204 6651
rect 216 6621 232 6651
rect 224 6574 226 6621
rect 300 6594 308 6663
rect 332 6661 342 6699
rect 400 6691 404 6700
rect 454 6685 504 6687
rect 494 6681 548 6685
rect 494 6676 514 6681
rect 504 6661 506 6676
rect 336 6649 342 6661
rect 289 6584 308 6594
rect 300 6578 308 6584
rect 332 6615 342 6649
rect 400 6653 404 6661
rect 400 6619 408 6653
rect 434 6619 438 6653
rect 498 6651 506 6661
rect 514 6651 515 6671
rect 504 6635 506 6651
rect 525 6642 528 6676
rect 547 6651 548 6671
rect 557 6651 564 6661
rect 514 6635 530 6641
rect 532 6635 548 6641
rect 332 6587 373 6615
rect 332 6581 351 6587
rect 107 6527 119 6561
rect 129 6527 149 6561
rect 196 6540 204 6574
rect 216 6540 232 6574
rect 244 6568 257 6574
rect 278 6568 291 6578
rect 244 6544 291 6568
rect 300 6568 321 6578
rect 336 6571 351 6581
rect 300 6544 329 6568
rect 332 6553 351 6571
rect 361 6581 375 6587
rect 400 6581 411 6619
rect 562 6582 612 6584
rect 361 6553 381 6581
rect 400 6553 409 6581
rect 466 6573 497 6581
rect 565 6573 596 6581
rect 442 6566 500 6573
rect 466 6565 500 6566
rect 565 6565 599 6573
rect 244 6540 257 6544
rect 42 6461 46 6495
rect 72 6461 76 6495
rect 42 6414 76 6418
rect 42 6399 46 6414
rect 72 6399 76 6414
rect 38 6381 80 6399
rect 16 6375 102 6381
rect 144 6375 148 6527
rect 174 6503 181 6531
rect 224 6493 226 6540
rect 300 6531 308 6544
rect 278 6520 305 6531
rect 332 6503 342 6553
rect 400 6533 404 6553
rect 497 6549 500 6565
rect 596 6549 599 6565
rect 466 6548 500 6549
rect 442 6541 500 6548
rect 565 6541 599 6549
rect 612 6532 614 6582
rect 256 6493 328 6501
rect 336 6495 342 6503
rect 400 6495 404 6503
rect 196 6463 204 6493
rect 216 6463 232 6493
rect 196 6459 232 6463
rect 196 6451 226 6459
rect 224 6435 226 6451
rect 332 6423 336 6491
rect 400 6461 408 6495
rect 434 6461 438 6495
rect 454 6479 504 6481
rect 504 6463 506 6479
rect 514 6473 530 6479
rect 532 6473 548 6479
rect 525 6463 548 6472
rect 400 6453 404 6461
rect 498 6453 506 6463
rect 504 6429 506 6453
rect 514 6443 515 6463
rect 525 6438 528 6463
rect 547 6443 548 6463
rect 557 6453 564 6463
rect 514 6429 548 6433
rect 400 6423 442 6424
rect 174 6413 246 6421
rect 400 6416 404 6423
rect 295 6382 300 6416
rect 324 6382 329 6416
rect 367 6399 438 6416
rect 367 6382 442 6399
rect 400 6381 442 6382
rect 378 6375 464 6381
rect 38 6359 80 6375
rect 400 6359 442 6375
rect -25 6345 25 6347
rect 42 6345 76 6359
rect 404 6345 438 6359
rect 455 6345 505 6347
rect 557 6345 607 6347
rect 16 6337 102 6345
rect 378 6337 464 6345
rect 8 6303 17 6337
rect 18 6335 51 6337
rect 80 6335 100 6337
rect 18 6303 100 6335
rect 380 6335 404 6337
rect 429 6335 438 6337
rect 442 6335 462 6337
rect 16 6295 102 6303
rect 42 6279 76 6295
rect 16 6259 38 6265
rect 42 6256 76 6260
rect 80 6259 102 6265
rect 42 6226 46 6256
rect 72 6226 76 6256
rect 42 6145 46 6179
rect 72 6145 76 6179
rect -25 6108 25 6110
rect -8 6100 14 6107
rect -8 6099 17 6100
rect 25 6099 27 6108
rect -12 6092 38 6099
rect -12 6091 34 6092
rect -12 6087 8 6091
rect 0 6075 8 6087
rect 14 6075 34 6091
rect 0 6074 34 6075
rect 0 6067 38 6074
rect 14 6066 17 6067
rect 25 6058 27 6067
rect 42 6038 45 6128
rect 69 6113 80 6145
rect 107 6113 143 6141
rect 144 6113 148 6333
rect 332 6265 336 6333
rect 380 6303 462 6335
rect 463 6303 472 6337
rect 480 6303 497 6337
rect 378 6295 464 6303
rect 505 6295 507 6345
rect 514 6303 548 6337
rect 565 6303 582 6337
rect 607 6295 609 6345
rect 404 6279 438 6295
rect 400 6265 442 6266
rect 378 6259 404 6265
rect 442 6259 464 6265
rect 400 6258 404 6259
rect 174 6219 246 6227
rect 295 6224 300 6258
rect 324 6224 329 6258
rect 224 6189 226 6205
rect 196 6181 226 6189
rect 332 6187 336 6255
rect 367 6224 438 6258
rect 400 6217 404 6224
rect 454 6211 504 6213
rect 494 6207 548 6211
rect 494 6202 514 6207
rect 504 6187 506 6202
rect 196 6177 232 6181
rect 196 6147 204 6177
rect 216 6147 232 6177
rect 400 6179 404 6187
rect 107 6107 119 6113
rect 109 6079 119 6107
rect 129 6079 149 6113
rect 174 6109 181 6139
rect 224 6100 226 6147
rect 256 6139 328 6147
rect 332 6145 336 6175
rect 400 6145 408 6179
rect 434 6145 438 6179
rect 498 6177 506 6187
rect 514 6177 515 6197
rect 504 6161 506 6177
rect 525 6168 528 6202
rect 547 6177 548 6197
rect 557 6177 564 6187
rect 514 6161 530 6167
rect 532 6161 548 6167
rect 278 6109 305 6120
rect 42 5987 46 6021
rect 72 5987 76 6021
rect 38 5949 80 5950
rect 42 5908 76 5942
rect 79 5908 113 5942
rect 42 5829 46 5863
rect 72 5829 76 5863
rect -25 5792 25 5794
rect -8 5784 14 5791
rect -8 5783 17 5784
rect 25 5783 27 5792
rect -12 5776 38 5783
rect -12 5775 34 5776
rect -12 5771 8 5775
rect 0 5759 8 5771
rect 14 5759 34 5775
rect 0 5758 34 5759
rect 0 5751 38 5758
rect 14 5750 17 5751
rect 25 5742 27 5751
rect 42 5722 45 5812
rect 71 5781 80 5809
rect 69 5743 80 5781
rect 144 5771 148 6079
rect 196 6066 204 6100
rect 216 6066 232 6100
rect 244 6096 257 6100
rect 300 6096 308 6109
rect 332 6107 342 6145
rect 400 6137 404 6145
rect 336 6097 342 6107
rect 244 6072 291 6096
rect 244 6066 257 6072
rect 224 6019 226 6066
rect 278 6062 291 6072
rect 300 6072 329 6096
rect 332 6087 342 6097
rect 400 6097 409 6125
rect 562 6108 612 6110
rect 466 6099 497 6107
rect 565 6099 596 6107
rect 300 6062 321 6072
rect 300 6056 308 6062
rect 289 6046 308 6056
rect 196 5989 204 6019
rect 216 5989 232 6019
rect 196 5985 232 5989
rect 196 5977 226 5985
rect 300 5977 308 6046
rect 332 6053 351 6087
rect 361 6059 381 6087
rect 361 6053 375 6059
rect 400 6053 411 6097
rect 442 6092 500 6099
rect 466 6091 500 6092
rect 565 6091 599 6099
rect 497 6075 500 6091
rect 596 6075 599 6091
rect 466 6074 500 6075
rect 442 6067 500 6074
rect 565 6067 599 6075
rect 612 6058 614 6108
rect 332 6029 342 6053
rect 336 6017 342 6029
rect 224 5961 226 5977
rect 332 5949 342 6017
rect 400 6021 404 6029
rect 400 5987 408 6021
rect 434 5987 438 6021
rect 454 6005 504 6007
rect 504 5989 506 6005
rect 514 5999 530 6005
rect 532 5999 548 6005
rect 525 5989 548 5998
rect 400 5979 404 5987
rect 498 5979 506 5989
rect 504 5955 506 5979
rect 514 5969 515 5989
rect 525 5964 528 5989
rect 547 5969 548 5989
rect 557 5979 564 5989
rect 514 5955 548 5959
rect 151 5908 156 5942
rect 174 5939 246 5947
rect 256 5939 328 5947
rect 336 5941 342 5949
rect 400 5944 404 5949
rect 180 5911 185 5939
rect 174 5903 246 5911
rect 256 5903 328 5911
rect 332 5909 336 5939
rect 400 5910 438 5944
rect 224 5873 226 5889
rect 196 5865 226 5873
rect 196 5861 232 5865
rect 196 5831 204 5861
rect 216 5831 232 5861
rect 224 5784 226 5831
rect 300 5804 308 5873
rect 332 5871 342 5909
rect 400 5901 404 5910
rect 454 5895 504 5897
rect 494 5891 548 5895
rect 494 5886 514 5891
rect 504 5871 506 5886
rect 336 5859 342 5871
rect 289 5794 308 5804
rect 300 5788 308 5794
rect 332 5825 342 5859
rect 400 5863 404 5871
rect 400 5829 408 5863
rect 434 5829 438 5863
rect 498 5861 506 5871
rect 514 5861 515 5881
rect 504 5845 506 5861
rect 525 5852 528 5886
rect 547 5861 548 5881
rect 557 5861 564 5871
rect 514 5845 530 5851
rect 532 5845 548 5851
rect 332 5797 373 5825
rect 332 5791 351 5797
rect 107 5737 119 5771
rect 129 5737 149 5771
rect 196 5750 204 5784
rect 216 5750 232 5784
rect 244 5778 257 5784
rect 278 5778 291 5788
rect 244 5754 291 5778
rect 300 5778 321 5788
rect 336 5781 351 5791
rect 300 5754 329 5778
rect 332 5763 351 5781
rect 361 5791 375 5797
rect 400 5791 411 5829
rect 562 5792 612 5794
rect 361 5763 381 5791
rect 400 5763 409 5791
rect 466 5783 497 5791
rect 565 5783 596 5791
rect 442 5776 500 5783
rect 466 5775 500 5776
rect 565 5775 599 5783
rect 244 5750 257 5754
rect 42 5671 46 5705
rect 72 5671 76 5705
rect 42 5624 76 5628
rect 42 5609 46 5624
rect 72 5609 76 5624
rect 38 5591 80 5609
rect 16 5585 102 5591
rect 144 5585 148 5737
rect 174 5713 181 5741
rect 224 5703 226 5750
rect 300 5741 308 5754
rect 278 5730 305 5741
rect 332 5713 342 5763
rect 400 5743 404 5763
rect 497 5759 500 5775
rect 596 5759 599 5775
rect 466 5758 500 5759
rect 442 5751 500 5758
rect 565 5751 599 5759
rect 612 5742 614 5792
rect 256 5703 328 5711
rect 336 5705 342 5713
rect 400 5705 404 5713
rect 196 5673 204 5703
rect 216 5673 232 5703
rect 196 5669 232 5673
rect 196 5661 226 5669
rect 224 5645 226 5661
rect 332 5633 336 5701
rect 400 5671 408 5705
rect 434 5671 438 5705
rect 454 5689 504 5691
rect 504 5673 506 5689
rect 514 5683 530 5689
rect 532 5683 548 5689
rect 525 5673 548 5682
rect 400 5663 404 5671
rect 498 5663 506 5673
rect 504 5639 506 5663
rect 514 5653 515 5673
rect 525 5648 528 5673
rect 547 5653 548 5673
rect 557 5663 564 5673
rect 514 5639 548 5643
rect 400 5633 442 5634
rect 174 5623 246 5631
rect 400 5626 404 5633
rect 295 5592 300 5626
rect 324 5592 329 5626
rect 367 5609 438 5626
rect 367 5592 442 5609
rect 400 5591 442 5592
rect 378 5585 464 5591
rect 38 5569 80 5585
rect 400 5569 442 5585
rect -25 5555 25 5557
rect 42 5555 76 5569
rect 404 5555 438 5569
rect 455 5555 505 5557
rect 557 5555 607 5557
rect 16 5547 102 5555
rect 378 5547 464 5555
rect 8 5513 17 5547
rect 18 5545 51 5547
rect 80 5545 100 5547
rect 18 5513 100 5545
rect 380 5545 404 5547
rect 429 5545 438 5547
rect 442 5545 462 5547
rect 16 5505 102 5513
rect 42 5489 76 5505
rect 16 5469 38 5475
rect 42 5466 76 5470
rect 80 5469 102 5475
rect 42 5436 46 5466
rect 72 5436 76 5466
rect 42 5355 46 5389
rect 72 5355 76 5389
rect -25 5318 25 5320
rect -8 5310 14 5317
rect -8 5309 17 5310
rect 25 5309 27 5318
rect -12 5302 38 5309
rect -12 5301 34 5302
rect -12 5297 8 5301
rect 0 5285 8 5297
rect 14 5285 34 5301
rect 0 5284 34 5285
rect 0 5277 38 5284
rect 14 5276 17 5277
rect 25 5268 27 5277
rect 42 5248 45 5338
rect 69 5323 80 5355
rect 107 5323 143 5351
rect 144 5323 148 5543
rect 332 5475 336 5543
rect 380 5513 462 5545
rect 463 5513 472 5547
rect 480 5513 497 5547
rect 378 5505 464 5513
rect 505 5505 507 5555
rect 514 5513 548 5547
rect 565 5513 582 5547
rect 607 5505 609 5555
rect 404 5489 438 5505
rect 400 5475 442 5476
rect 378 5469 404 5475
rect 442 5469 464 5475
rect 400 5468 404 5469
rect 174 5429 246 5437
rect 295 5434 300 5468
rect 324 5434 329 5468
rect 224 5399 226 5415
rect 196 5391 226 5399
rect 332 5397 336 5465
rect 367 5434 438 5468
rect 400 5427 404 5434
rect 454 5421 504 5423
rect 494 5417 548 5421
rect 494 5412 514 5417
rect 504 5397 506 5412
rect 196 5387 232 5391
rect 196 5357 204 5387
rect 216 5357 232 5387
rect 400 5389 404 5397
rect 107 5317 119 5323
rect 109 5289 119 5317
rect 129 5289 149 5323
rect 174 5319 181 5349
rect 224 5310 226 5357
rect 256 5349 328 5357
rect 332 5355 336 5385
rect 400 5355 408 5389
rect 434 5355 438 5389
rect 498 5387 506 5397
rect 514 5387 515 5407
rect 504 5371 506 5387
rect 525 5378 528 5412
rect 547 5387 548 5407
rect 557 5387 564 5397
rect 514 5371 530 5377
rect 532 5371 548 5377
rect 278 5319 305 5330
rect 42 5197 46 5231
rect 72 5197 76 5231
rect 38 5159 80 5160
rect 42 5118 76 5152
rect 79 5118 113 5152
rect 42 5039 46 5073
rect 72 5039 76 5073
rect -25 5002 25 5004
rect -8 4994 14 5001
rect -8 4993 17 4994
rect 25 4993 27 5002
rect -12 4986 38 4993
rect -12 4985 34 4986
rect -12 4981 8 4985
rect 0 4969 8 4981
rect 14 4969 34 4985
rect 0 4968 34 4969
rect 0 4961 38 4968
rect 14 4960 17 4961
rect 25 4952 27 4961
rect 42 4932 45 5022
rect 71 4991 80 5019
rect 69 4953 80 4991
rect 144 4981 148 5289
rect 196 5276 204 5310
rect 216 5276 232 5310
rect 244 5306 257 5310
rect 300 5306 308 5319
rect 332 5317 342 5355
rect 400 5347 404 5355
rect 336 5307 342 5317
rect 244 5282 291 5306
rect 244 5276 257 5282
rect 224 5229 226 5276
rect 278 5272 291 5282
rect 300 5282 329 5306
rect 332 5297 342 5307
rect 400 5307 409 5335
rect 562 5318 612 5320
rect 466 5309 497 5317
rect 565 5309 596 5317
rect 300 5272 321 5282
rect 300 5266 308 5272
rect 289 5256 308 5266
rect 196 5199 204 5229
rect 216 5199 232 5229
rect 196 5195 232 5199
rect 196 5187 226 5195
rect 300 5187 308 5256
rect 332 5263 351 5297
rect 361 5269 381 5297
rect 361 5263 375 5269
rect 400 5263 411 5307
rect 442 5302 500 5309
rect 466 5301 500 5302
rect 565 5301 599 5309
rect 497 5285 500 5301
rect 596 5285 599 5301
rect 466 5284 500 5285
rect 442 5277 500 5284
rect 565 5277 599 5285
rect 612 5268 614 5318
rect 332 5239 342 5263
rect 336 5227 342 5239
rect 224 5171 226 5187
rect 332 5159 342 5227
rect 400 5231 404 5239
rect 400 5197 408 5231
rect 434 5197 438 5231
rect 454 5215 504 5217
rect 504 5199 506 5215
rect 514 5209 530 5215
rect 532 5209 548 5215
rect 525 5199 548 5208
rect 400 5189 404 5197
rect 498 5189 506 5199
rect 504 5165 506 5189
rect 514 5179 515 5199
rect 525 5174 528 5199
rect 547 5179 548 5199
rect 557 5189 564 5199
rect 514 5165 548 5169
rect 151 5118 156 5152
rect 174 5149 246 5157
rect 256 5149 328 5157
rect 336 5151 342 5159
rect 400 5154 404 5159
rect 180 5121 185 5149
rect 174 5113 246 5121
rect 256 5113 328 5121
rect 332 5119 336 5149
rect 400 5120 438 5154
rect 224 5083 226 5099
rect 196 5075 226 5083
rect 196 5071 232 5075
rect 196 5041 204 5071
rect 216 5041 232 5071
rect 224 4994 226 5041
rect 300 5014 308 5083
rect 332 5081 342 5119
rect 400 5111 404 5120
rect 454 5105 504 5107
rect 494 5101 548 5105
rect 494 5096 514 5101
rect 504 5081 506 5096
rect 336 5069 342 5081
rect 289 5004 308 5014
rect 300 4998 308 5004
rect 332 5035 342 5069
rect 400 5073 404 5081
rect 400 5039 408 5073
rect 434 5039 438 5073
rect 498 5071 506 5081
rect 514 5071 515 5091
rect 504 5055 506 5071
rect 525 5062 528 5096
rect 547 5071 548 5091
rect 557 5071 564 5081
rect 514 5055 530 5061
rect 532 5055 548 5061
rect 332 5007 373 5035
rect 332 5001 351 5007
rect 107 4947 119 4981
rect 129 4947 149 4981
rect 196 4960 204 4994
rect 216 4960 232 4994
rect 244 4988 257 4994
rect 278 4988 291 4998
rect 244 4964 291 4988
rect 300 4988 321 4998
rect 336 4991 351 5001
rect 300 4964 329 4988
rect 332 4973 351 4991
rect 361 5001 375 5007
rect 400 5001 411 5039
rect 562 5002 612 5004
rect 361 4973 381 5001
rect 400 4973 409 5001
rect 466 4993 497 5001
rect 565 4993 596 5001
rect 442 4986 500 4993
rect 466 4985 500 4986
rect 565 4985 599 4993
rect 244 4960 257 4964
rect 42 4881 46 4915
rect 72 4881 76 4915
rect 42 4834 76 4838
rect 42 4819 46 4834
rect 72 4819 76 4834
rect 38 4801 80 4819
rect 16 4795 102 4801
rect 144 4795 148 4947
rect 174 4923 181 4951
rect 224 4913 226 4960
rect 300 4951 308 4964
rect 278 4940 305 4951
rect 332 4923 342 4973
rect 400 4953 404 4973
rect 497 4969 500 4985
rect 596 4969 599 4985
rect 466 4968 500 4969
rect 442 4961 500 4968
rect 565 4961 599 4969
rect 612 4952 614 5002
rect 256 4913 328 4921
rect 336 4915 342 4923
rect 400 4915 404 4923
rect 196 4883 204 4913
rect 216 4883 232 4913
rect 196 4879 232 4883
rect 196 4871 226 4879
rect 224 4855 226 4871
rect 332 4843 336 4911
rect 400 4881 408 4915
rect 434 4881 438 4915
rect 454 4899 504 4901
rect 504 4883 506 4899
rect 514 4893 530 4899
rect 532 4893 548 4899
rect 525 4883 548 4892
rect 400 4873 404 4881
rect 498 4873 506 4883
rect 504 4849 506 4873
rect 514 4863 515 4883
rect 525 4858 528 4883
rect 547 4863 548 4883
rect 557 4873 564 4883
rect 514 4849 548 4853
rect 400 4843 442 4844
rect 174 4833 246 4841
rect 400 4836 404 4843
rect 295 4802 300 4836
rect 324 4802 329 4836
rect 367 4819 438 4836
rect 367 4802 442 4819
rect 400 4801 442 4802
rect 378 4795 464 4801
rect 38 4779 80 4795
rect 400 4779 442 4795
rect -25 4765 25 4767
rect 42 4765 76 4779
rect 404 4765 438 4779
rect 455 4765 505 4767
rect 557 4765 607 4767
rect 16 4757 102 4765
rect 378 4757 464 4765
rect 8 4723 17 4757
rect 18 4755 51 4757
rect 80 4755 100 4757
rect 18 4723 100 4755
rect 380 4755 404 4757
rect 429 4755 438 4757
rect 442 4755 462 4757
rect 16 4715 102 4723
rect 42 4699 76 4715
rect 16 4679 38 4685
rect 42 4676 76 4680
rect 80 4679 102 4685
rect 42 4646 46 4676
rect 72 4646 76 4676
rect 42 4565 46 4599
rect 72 4565 76 4599
rect -25 4528 25 4530
rect -8 4520 14 4527
rect -8 4519 17 4520
rect 25 4519 27 4528
rect -12 4512 38 4519
rect -12 4511 34 4512
rect -12 4507 8 4511
rect 0 4495 8 4507
rect 14 4495 34 4511
rect 0 4494 34 4495
rect 0 4487 38 4494
rect 14 4486 17 4487
rect 25 4478 27 4487
rect 42 4458 45 4548
rect 69 4533 80 4565
rect 107 4533 143 4561
rect 144 4533 148 4753
rect 332 4685 336 4753
rect 380 4723 462 4755
rect 463 4723 472 4757
rect 480 4723 497 4757
rect 378 4715 464 4723
rect 505 4715 507 4765
rect 514 4723 548 4757
rect 565 4723 582 4757
rect 607 4715 609 4765
rect 404 4699 438 4715
rect 400 4685 442 4686
rect 378 4679 404 4685
rect 442 4679 464 4685
rect 400 4678 404 4679
rect 174 4639 246 4647
rect 295 4644 300 4678
rect 324 4644 329 4678
rect 224 4609 226 4625
rect 196 4601 226 4609
rect 332 4607 336 4675
rect 367 4644 438 4678
rect 400 4637 404 4644
rect 454 4631 504 4633
rect 494 4627 548 4631
rect 494 4622 514 4627
rect 504 4607 506 4622
rect 196 4597 232 4601
rect 196 4567 204 4597
rect 216 4567 232 4597
rect 400 4599 404 4607
rect 107 4527 119 4533
rect 109 4499 119 4527
rect 129 4499 149 4533
rect 174 4529 181 4559
rect 224 4520 226 4567
rect 256 4559 328 4567
rect 332 4565 336 4595
rect 400 4565 408 4599
rect 434 4565 438 4599
rect 498 4597 506 4607
rect 514 4597 515 4617
rect 504 4581 506 4597
rect 525 4588 528 4622
rect 547 4597 548 4617
rect 557 4597 564 4607
rect 514 4581 530 4587
rect 532 4581 548 4587
rect 278 4529 305 4540
rect 42 4407 46 4441
rect 72 4407 76 4441
rect 38 4369 80 4370
rect 42 4328 76 4362
rect 79 4328 113 4362
rect 42 4249 46 4283
rect 72 4249 76 4283
rect -25 4212 25 4214
rect -8 4204 14 4211
rect -8 4203 17 4204
rect 25 4203 27 4212
rect -12 4196 38 4203
rect -12 4195 34 4196
rect -12 4191 8 4195
rect 0 4179 8 4191
rect 14 4179 34 4195
rect 0 4178 34 4179
rect 0 4171 38 4178
rect 14 4170 17 4171
rect 25 4162 27 4171
rect 42 4142 45 4232
rect 71 4201 80 4229
rect 69 4163 80 4201
rect 144 4191 148 4499
rect 196 4486 204 4520
rect 216 4486 232 4520
rect 244 4516 257 4520
rect 300 4516 308 4529
rect 332 4527 342 4565
rect 400 4557 404 4565
rect 336 4517 342 4527
rect 244 4492 291 4516
rect 244 4486 257 4492
rect 224 4439 226 4486
rect 278 4482 291 4492
rect 300 4492 329 4516
rect 332 4507 342 4517
rect 400 4517 409 4545
rect 562 4528 612 4530
rect 466 4519 497 4527
rect 565 4519 596 4527
rect 300 4482 321 4492
rect 300 4476 308 4482
rect 289 4466 308 4476
rect 196 4409 204 4439
rect 216 4409 232 4439
rect 196 4405 232 4409
rect 196 4397 226 4405
rect 300 4397 308 4466
rect 332 4473 351 4507
rect 361 4479 381 4507
rect 361 4473 375 4479
rect 400 4473 411 4517
rect 442 4512 500 4519
rect 466 4511 500 4512
rect 565 4511 599 4519
rect 497 4495 500 4511
rect 596 4495 599 4511
rect 466 4494 500 4495
rect 442 4487 500 4494
rect 565 4487 599 4495
rect 612 4478 614 4528
rect 332 4449 342 4473
rect 336 4437 342 4449
rect 224 4381 226 4397
rect 332 4369 342 4437
rect 400 4441 404 4449
rect 400 4407 408 4441
rect 434 4407 438 4441
rect 454 4425 504 4427
rect 504 4409 506 4425
rect 514 4419 530 4425
rect 532 4419 548 4425
rect 525 4409 548 4418
rect 400 4399 404 4407
rect 498 4399 506 4409
rect 504 4375 506 4399
rect 514 4389 515 4409
rect 525 4384 528 4409
rect 547 4389 548 4409
rect 557 4399 564 4409
rect 514 4375 548 4379
rect 151 4328 156 4362
rect 174 4359 246 4367
rect 256 4359 328 4367
rect 336 4361 342 4369
rect 400 4364 404 4369
rect 180 4331 185 4359
rect 174 4323 246 4331
rect 256 4323 328 4331
rect 332 4329 336 4359
rect 400 4330 438 4364
rect 224 4293 226 4309
rect 196 4285 226 4293
rect 196 4281 232 4285
rect 196 4251 204 4281
rect 216 4251 232 4281
rect 224 4204 226 4251
rect 300 4224 308 4293
rect 332 4291 342 4329
rect 400 4321 404 4330
rect 454 4315 504 4317
rect 494 4311 548 4315
rect 494 4306 514 4311
rect 504 4291 506 4306
rect 336 4279 342 4291
rect 289 4214 308 4224
rect 300 4208 308 4214
rect 332 4245 342 4279
rect 400 4283 404 4291
rect 400 4249 408 4283
rect 434 4249 438 4283
rect 498 4281 506 4291
rect 514 4281 515 4301
rect 504 4265 506 4281
rect 525 4272 528 4306
rect 547 4281 548 4301
rect 557 4281 564 4291
rect 514 4265 530 4271
rect 532 4265 548 4271
rect 332 4217 373 4245
rect 332 4211 351 4217
rect 107 4157 119 4191
rect 129 4157 149 4191
rect 196 4170 204 4204
rect 216 4170 232 4204
rect 244 4198 257 4204
rect 278 4198 291 4208
rect 244 4174 291 4198
rect 300 4198 321 4208
rect 336 4201 351 4211
rect 300 4174 329 4198
rect 332 4183 351 4201
rect 361 4211 375 4217
rect 400 4211 411 4249
rect 562 4212 612 4214
rect 361 4183 381 4211
rect 400 4183 409 4211
rect 466 4203 497 4211
rect 565 4203 596 4211
rect 442 4196 500 4203
rect 466 4195 500 4196
rect 565 4195 599 4203
rect 244 4170 257 4174
rect 42 4091 46 4125
rect 72 4091 76 4125
rect 42 4044 76 4048
rect 42 4029 46 4044
rect 72 4029 76 4044
rect 38 4011 80 4029
rect 16 4005 102 4011
rect 144 4005 148 4157
rect 174 4133 181 4161
rect 224 4123 226 4170
rect 300 4161 308 4174
rect 278 4150 305 4161
rect 332 4133 342 4183
rect 400 4163 404 4183
rect 497 4179 500 4195
rect 596 4179 599 4195
rect 466 4178 500 4179
rect 442 4171 500 4178
rect 565 4171 599 4179
rect 612 4162 614 4212
rect 256 4123 328 4131
rect 336 4125 342 4133
rect 400 4125 404 4133
rect 196 4093 204 4123
rect 216 4093 232 4123
rect 196 4089 232 4093
rect 196 4081 226 4089
rect 224 4065 226 4081
rect 332 4053 336 4121
rect 400 4091 408 4125
rect 434 4091 438 4125
rect 454 4109 504 4111
rect 504 4093 506 4109
rect 514 4103 530 4109
rect 532 4103 548 4109
rect 525 4093 548 4102
rect 400 4083 404 4091
rect 498 4083 506 4093
rect 504 4059 506 4083
rect 514 4073 515 4093
rect 525 4068 528 4093
rect 547 4073 548 4093
rect 557 4083 564 4093
rect 514 4059 548 4063
rect 400 4053 442 4054
rect 174 4043 246 4051
rect 400 4046 404 4053
rect 295 4012 300 4046
rect 324 4012 329 4046
rect 367 4029 438 4046
rect 367 4012 442 4029
rect 400 4011 442 4012
rect 378 4005 464 4011
rect 38 3989 80 4005
rect 400 3989 442 4005
rect -25 3975 25 3977
rect 42 3975 76 3989
rect 404 3975 438 3989
rect 455 3975 505 3977
rect 557 3975 607 3977
rect 16 3967 102 3975
rect 378 3967 464 3975
rect 8 3933 17 3967
rect 18 3965 51 3967
rect 80 3965 100 3967
rect 18 3933 100 3965
rect 380 3965 404 3967
rect 429 3965 438 3967
rect 442 3965 462 3967
rect 16 3925 102 3933
rect 42 3909 76 3925
rect 16 3889 38 3895
rect 42 3886 76 3890
rect 80 3889 102 3895
rect 42 3856 46 3886
rect 72 3856 76 3886
rect 42 3775 46 3809
rect 72 3775 76 3809
rect -25 3738 25 3740
rect -8 3730 14 3737
rect -8 3729 17 3730
rect 25 3729 27 3738
rect -12 3722 38 3729
rect -12 3721 34 3722
rect -12 3717 8 3721
rect 0 3705 8 3717
rect 14 3705 34 3721
rect 0 3704 34 3705
rect 0 3697 38 3704
rect 14 3696 17 3697
rect 25 3688 27 3697
rect 42 3668 45 3758
rect 69 3743 80 3775
rect 107 3743 143 3771
rect 144 3743 148 3963
rect 332 3895 336 3963
rect 380 3933 462 3965
rect 463 3933 472 3967
rect 480 3933 497 3967
rect 378 3925 464 3933
rect 505 3925 507 3975
rect 514 3933 548 3967
rect 565 3933 582 3967
rect 607 3925 609 3975
rect 404 3909 438 3925
rect 400 3895 442 3896
rect 378 3889 404 3895
rect 442 3889 464 3895
rect 400 3888 404 3889
rect 174 3849 246 3857
rect 295 3854 300 3888
rect 324 3854 329 3888
rect 224 3819 226 3835
rect 196 3811 226 3819
rect 332 3817 336 3885
rect 367 3854 438 3888
rect 400 3847 404 3854
rect 454 3841 504 3843
rect 494 3837 548 3841
rect 494 3832 514 3837
rect 504 3817 506 3832
rect 196 3807 232 3811
rect 196 3777 204 3807
rect 216 3777 232 3807
rect 400 3809 404 3817
rect 107 3737 119 3743
rect 109 3709 119 3737
rect 129 3709 149 3743
rect 174 3739 181 3769
rect 224 3730 226 3777
rect 256 3769 328 3777
rect 332 3775 336 3805
rect 400 3775 408 3809
rect 434 3775 438 3809
rect 498 3807 506 3817
rect 514 3807 515 3827
rect 504 3791 506 3807
rect 525 3798 528 3832
rect 547 3807 548 3827
rect 557 3807 564 3817
rect 514 3791 530 3797
rect 532 3791 548 3797
rect 278 3739 305 3750
rect 42 3617 46 3651
rect 72 3617 76 3651
rect 38 3579 80 3580
rect 42 3538 76 3572
rect 79 3538 113 3572
rect 42 3459 46 3493
rect 72 3459 76 3493
rect -25 3422 25 3424
rect -8 3414 14 3421
rect -8 3413 17 3414
rect 25 3413 27 3422
rect -12 3406 38 3413
rect -12 3405 34 3406
rect -12 3401 8 3405
rect 0 3389 8 3401
rect 14 3389 34 3405
rect 0 3388 34 3389
rect 0 3381 38 3388
rect 14 3380 17 3381
rect 25 3372 27 3381
rect 42 3352 45 3442
rect 71 3411 80 3439
rect 69 3373 80 3411
rect 144 3401 148 3709
rect 196 3696 204 3730
rect 216 3696 232 3730
rect 244 3726 257 3730
rect 300 3726 308 3739
rect 332 3737 342 3775
rect 400 3767 404 3775
rect 336 3727 342 3737
rect 244 3702 291 3726
rect 244 3696 257 3702
rect 224 3649 226 3696
rect 278 3692 291 3702
rect 300 3702 329 3726
rect 332 3717 342 3727
rect 400 3727 409 3755
rect 562 3738 612 3740
rect 466 3729 497 3737
rect 565 3729 596 3737
rect 300 3692 321 3702
rect 300 3686 308 3692
rect 289 3676 308 3686
rect 196 3619 204 3649
rect 216 3619 232 3649
rect 196 3615 232 3619
rect 196 3607 226 3615
rect 300 3607 308 3676
rect 332 3683 351 3717
rect 361 3689 381 3717
rect 361 3683 375 3689
rect 400 3683 411 3727
rect 442 3722 500 3729
rect 466 3721 500 3722
rect 565 3721 599 3729
rect 497 3705 500 3721
rect 596 3705 599 3721
rect 466 3704 500 3705
rect 442 3697 500 3704
rect 565 3697 599 3705
rect 612 3688 614 3738
rect 332 3659 342 3683
rect 336 3647 342 3659
rect 224 3591 226 3607
rect 332 3579 342 3647
rect 400 3651 404 3659
rect 400 3617 408 3651
rect 434 3617 438 3651
rect 454 3635 504 3637
rect 504 3619 506 3635
rect 514 3629 530 3635
rect 532 3629 548 3635
rect 525 3619 548 3628
rect 400 3609 404 3617
rect 498 3609 506 3619
rect 504 3585 506 3609
rect 514 3599 515 3619
rect 525 3594 528 3619
rect 547 3599 548 3619
rect 557 3609 564 3619
rect 514 3585 548 3589
rect 151 3538 156 3572
rect 174 3569 246 3577
rect 256 3569 328 3577
rect 336 3571 342 3579
rect 400 3574 404 3579
rect 180 3541 185 3569
rect 174 3533 246 3541
rect 256 3533 328 3541
rect 332 3539 336 3569
rect 400 3540 438 3574
rect 224 3503 226 3519
rect 196 3495 226 3503
rect 196 3491 232 3495
rect 196 3461 204 3491
rect 216 3461 232 3491
rect 224 3414 226 3461
rect 300 3434 308 3503
rect 332 3501 342 3539
rect 400 3531 404 3540
rect 454 3525 504 3527
rect 494 3521 548 3525
rect 494 3516 514 3521
rect 504 3501 506 3516
rect 336 3489 342 3501
rect 289 3424 308 3434
rect 300 3418 308 3424
rect 332 3455 342 3489
rect 400 3493 404 3501
rect 400 3459 408 3493
rect 434 3459 438 3493
rect 498 3491 506 3501
rect 514 3491 515 3511
rect 504 3475 506 3491
rect 525 3482 528 3516
rect 547 3491 548 3511
rect 557 3491 564 3501
rect 514 3475 530 3481
rect 532 3475 548 3481
rect 332 3427 373 3455
rect 332 3421 351 3427
rect 107 3367 119 3401
rect 129 3367 149 3401
rect 196 3380 204 3414
rect 216 3380 232 3414
rect 244 3408 257 3414
rect 278 3408 291 3418
rect 244 3384 291 3408
rect 300 3408 321 3418
rect 336 3411 351 3421
rect 300 3384 329 3408
rect 332 3393 351 3411
rect 361 3421 375 3427
rect 400 3421 411 3459
rect 562 3422 612 3424
rect 361 3393 381 3421
rect 400 3393 409 3421
rect 466 3413 497 3421
rect 565 3413 596 3421
rect 442 3406 500 3413
rect 466 3405 500 3406
rect 565 3405 599 3413
rect 244 3380 257 3384
rect 42 3301 46 3335
rect 72 3301 76 3335
rect 42 3254 76 3258
rect 42 3239 46 3254
rect 72 3239 76 3254
rect 38 3221 80 3239
rect 16 3215 102 3221
rect 144 3215 148 3367
rect 174 3343 181 3371
rect 224 3333 226 3380
rect 300 3371 308 3384
rect 278 3360 305 3371
rect 332 3343 342 3393
rect 400 3373 404 3393
rect 497 3389 500 3405
rect 596 3389 599 3405
rect 466 3388 500 3389
rect 442 3381 500 3388
rect 565 3381 599 3389
rect 612 3372 614 3422
rect 256 3333 328 3341
rect 336 3335 342 3343
rect 400 3335 404 3343
rect 196 3303 204 3333
rect 216 3303 232 3333
rect 196 3299 232 3303
rect 196 3291 226 3299
rect 224 3275 226 3291
rect 332 3263 336 3331
rect 400 3301 408 3335
rect 434 3301 438 3335
rect 454 3319 504 3321
rect 504 3303 506 3319
rect 514 3313 530 3319
rect 532 3313 548 3319
rect 525 3303 548 3312
rect 400 3293 404 3301
rect 498 3293 506 3303
rect 504 3269 506 3293
rect 514 3283 515 3303
rect 525 3278 528 3303
rect 547 3283 548 3303
rect 557 3293 564 3303
rect 514 3269 548 3273
rect 400 3263 442 3264
rect 174 3253 246 3261
rect 400 3256 404 3263
rect 295 3222 300 3256
rect 324 3222 329 3256
rect 367 3239 438 3256
rect 367 3222 442 3239
rect 400 3221 442 3222
rect 378 3215 464 3221
rect 38 3199 80 3215
rect 400 3199 442 3215
rect -25 3185 25 3187
rect 42 3185 76 3199
rect 404 3185 438 3199
rect 455 3185 505 3187
rect 557 3185 607 3187
rect 16 3177 102 3185
rect 378 3177 464 3185
rect 8 3143 17 3177
rect 18 3175 51 3177
rect 80 3175 100 3177
rect 18 3143 100 3175
rect 380 3175 404 3177
rect 429 3175 438 3177
rect 442 3175 462 3177
rect 16 3135 102 3143
rect 42 3119 76 3135
rect 16 3099 38 3105
rect 42 3096 76 3100
rect 80 3099 102 3105
rect 42 3066 46 3096
rect 72 3066 76 3096
rect 42 2985 46 3019
rect 72 2985 76 3019
rect -25 2948 25 2950
rect -8 2940 14 2947
rect -8 2939 17 2940
rect 25 2939 27 2948
rect -12 2932 38 2939
rect -12 2931 34 2932
rect -12 2927 8 2931
rect 0 2915 8 2927
rect 14 2915 34 2931
rect 0 2914 34 2915
rect 0 2907 38 2914
rect 14 2906 17 2907
rect 25 2898 27 2907
rect 42 2878 45 2968
rect 69 2953 80 2985
rect 107 2953 143 2981
rect 144 2953 148 3173
rect 332 3105 336 3173
rect 380 3143 462 3175
rect 463 3143 472 3177
rect 480 3143 497 3177
rect 378 3135 464 3143
rect 505 3135 507 3185
rect 514 3143 548 3177
rect 565 3143 582 3177
rect 607 3135 609 3185
rect 404 3119 438 3135
rect 400 3105 442 3106
rect 378 3099 404 3105
rect 442 3099 464 3105
rect 400 3098 404 3099
rect 174 3059 246 3067
rect 295 3064 300 3098
rect 324 3064 329 3098
rect 224 3029 226 3045
rect 196 3021 226 3029
rect 332 3027 336 3095
rect 367 3064 438 3098
rect 400 3057 404 3064
rect 454 3051 504 3053
rect 494 3047 548 3051
rect 494 3042 514 3047
rect 504 3027 506 3042
rect 196 3017 232 3021
rect 196 2987 204 3017
rect 216 2987 232 3017
rect 400 3019 404 3027
rect 107 2947 119 2953
rect 109 2919 119 2947
rect 129 2919 149 2953
rect 174 2949 181 2979
rect 224 2940 226 2987
rect 256 2979 328 2987
rect 332 2985 336 3015
rect 400 2985 408 3019
rect 434 2985 438 3019
rect 498 3017 506 3027
rect 514 3017 515 3037
rect 504 3001 506 3017
rect 525 3008 528 3042
rect 547 3017 548 3037
rect 557 3017 564 3027
rect 514 3001 530 3007
rect 532 3001 548 3007
rect 278 2949 305 2960
rect 42 2827 46 2861
rect 72 2827 76 2861
rect 38 2789 80 2790
rect 42 2748 76 2782
rect 79 2748 113 2782
rect 42 2669 46 2703
rect 72 2669 76 2703
rect -25 2632 25 2634
rect -8 2624 14 2631
rect -8 2623 17 2624
rect 25 2623 27 2632
rect -12 2616 38 2623
rect -12 2615 34 2616
rect -12 2611 8 2615
rect 0 2599 8 2611
rect 14 2599 34 2615
rect 0 2598 34 2599
rect 0 2591 38 2598
rect 14 2590 17 2591
rect 25 2582 27 2591
rect 42 2562 45 2652
rect 71 2621 80 2649
rect 69 2583 80 2621
rect 144 2611 148 2919
rect 196 2906 204 2940
rect 216 2906 232 2940
rect 244 2936 257 2940
rect 300 2936 308 2949
rect 332 2947 342 2985
rect 400 2977 404 2985
rect 336 2937 342 2947
rect 244 2912 291 2936
rect 244 2906 257 2912
rect 224 2859 226 2906
rect 278 2902 291 2912
rect 300 2912 329 2936
rect 332 2927 342 2937
rect 400 2937 409 2965
rect 562 2948 612 2950
rect 466 2939 497 2947
rect 565 2939 596 2947
rect 300 2902 321 2912
rect 300 2896 308 2902
rect 289 2886 308 2896
rect 196 2829 204 2859
rect 216 2829 232 2859
rect 196 2825 232 2829
rect 196 2817 226 2825
rect 300 2817 308 2886
rect 332 2893 351 2927
rect 361 2899 381 2927
rect 361 2893 375 2899
rect 400 2893 411 2937
rect 442 2932 500 2939
rect 466 2931 500 2932
rect 565 2931 599 2939
rect 497 2915 500 2931
rect 596 2915 599 2931
rect 466 2914 500 2915
rect 442 2907 500 2914
rect 565 2907 599 2915
rect 612 2898 614 2948
rect 332 2869 342 2893
rect 336 2857 342 2869
rect 224 2801 226 2817
rect 332 2789 342 2857
rect 400 2861 404 2869
rect 400 2827 408 2861
rect 434 2827 438 2861
rect 454 2845 504 2847
rect 504 2829 506 2845
rect 514 2839 530 2845
rect 532 2839 548 2845
rect 525 2829 548 2838
rect 400 2819 404 2827
rect 498 2819 506 2829
rect 504 2795 506 2819
rect 514 2809 515 2829
rect 525 2804 528 2829
rect 547 2809 548 2829
rect 557 2819 564 2829
rect 514 2795 548 2799
rect 151 2748 156 2782
rect 174 2779 246 2787
rect 256 2779 328 2787
rect 336 2781 342 2789
rect 400 2784 404 2789
rect 180 2751 185 2779
rect 174 2743 246 2751
rect 256 2743 328 2751
rect 332 2749 336 2779
rect 400 2750 438 2784
rect 224 2713 226 2729
rect 196 2705 226 2713
rect 196 2701 232 2705
rect 196 2671 204 2701
rect 216 2671 232 2701
rect 224 2624 226 2671
rect 300 2644 308 2713
rect 332 2711 342 2749
rect 400 2741 404 2750
rect 454 2735 504 2737
rect 494 2731 548 2735
rect 494 2726 514 2731
rect 504 2711 506 2726
rect 336 2699 342 2711
rect 289 2634 308 2644
rect 300 2628 308 2634
rect 332 2665 342 2699
rect 400 2703 404 2711
rect 400 2669 408 2703
rect 434 2669 438 2703
rect 498 2701 506 2711
rect 514 2701 515 2721
rect 504 2685 506 2701
rect 525 2692 528 2726
rect 547 2701 548 2721
rect 557 2701 564 2711
rect 514 2685 530 2691
rect 532 2685 548 2691
rect 332 2637 373 2665
rect 332 2631 351 2637
rect 107 2577 119 2611
rect 129 2577 149 2611
rect 196 2590 204 2624
rect 216 2590 232 2624
rect 244 2618 257 2624
rect 278 2618 291 2628
rect 244 2594 291 2618
rect 300 2618 321 2628
rect 336 2621 351 2631
rect 300 2594 329 2618
rect 332 2603 351 2621
rect 361 2631 375 2637
rect 400 2631 411 2669
rect 562 2632 612 2634
rect 361 2603 381 2631
rect 400 2603 409 2631
rect 466 2623 497 2631
rect 565 2623 596 2631
rect 442 2616 500 2623
rect 466 2615 500 2616
rect 565 2615 599 2623
rect 244 2590 257 2594
rect 42 2511 46 2545
rect 72 2511 76 2545
rect 42 2464 76 2468
rect 42 2449 46 2464
rect 72 2449 76 2464
rect 38 2431 80 2449
rect 16 2425 102 2431
rect 144 2425 148 2577
rect 174 2553 181 2581
rect 224 2543 226 2590
rect 300 2581 308 2594
rect 278 2570 305 2581
rect 332 2553 342 2603
rect 400 2583 404 2603
rect 497 2599 500 2615
rect 596 2599 599 2615
rect 466 2598 500 2599
rect 442 2591 500 2598
rect 565 2591 599 2599
rect 612 2582 614 2632
rect 256 2543 328 2551
rect 336 2545 342 2553
rect 400 2545 404 2553
rect 196 2513 204 2543
rect 216 2513 232 2543
rect 196 2509 232 2513
rect 196 2501 226 2509
rect 224 2485 226 2501
rect 332 2473 336 2541
rect 400 2511 408 2545
rect 434 2511 438 2545
rect 454 2529 504 2531
rect 504 2513 506 2529
rect 514 2523 530 2529
rect 532 2523 548 2529
rect 525 2513 548 2522
rect 400 2503 404 2511
rect 498 2503 506 2513
rect 504 2479 506 2503
rect 514 2493 515 2513
rect 525 2488 528 2513
rect 547 2493 548 2513
rect 557 2503 564 2513
rect 514 2479 548 2483
rect 400 2473 442 2474
rect 174 2463 246 2471
rect 400 2466 404 2473
rect 295 2432 300 2466
rect 324 2432 329 2466
rect 367 2449 438 2466
rect 367 2432 442 2449
rect 400 2431 442 2432
rect 378 2425 464 2431
rect 38 2409 80 2425
rect 400 2409 442 2425
rect -25 2395 25 2397
rect 42 2395 76 2409
rect 404 2395 438 2409
rect 455 2395 505 2397
rect 557 2395 607 2397
rect 16 2387 102 2395
rect 378 2387 464 2395
rect 8 2353 17 2387
rect 18 2385 51 2387
rect 80 2385 100 2387
rect 18 2353 100 2385
rect 380 2385 404 2387
rect 429 2385 438 2387
rect 442 2385 462 2387
rect 16 2345 102 2353
rect 42 2329 76 2345
rect 16 2309 38 2315
rect 42 2306 76 2310
rect 80 2309 102 2315
rect 42 2276 46 2306
rect 72 2276 76 2306
rect 42 2195 46 2229
rect 72 2195 76 2229
rect -25 2158 25 2160
rect -8 2150 14 2157
rect -8 2149 17 2150
rect 25 2149 27 2158
rect -12 2142 38 2149
rect -12 2141 34 2142
rect -12 2137 8 2141
rect 0 2125 8 2137
rect 14 2125 34 2141
rect 0 2124 34 2125
rect 0 2117 38 2124
rect 14 2116 17 2117
rect 25 2108 27 2117
rect 42 2088 45 2178
rect 69 2163 80 2195
rect 107 2163 143 2191
rect 144 2163 148 2383
rect 332 2315 336 2383
rect 380 2353 462 2385
rect 463 2353 472 2387
rect 480 2353 497 2387
rect 378 2345 464 2353
rect 505 2345 507 2395
rect 514 2353 548 2387
rect 565 2353 582 2387
rect 607 2345 609 2395
rect 404 2329 438 2345
rect 400 2315 442 2316
rect 378 2309 404 2315
rect 442 2309 464 2315
rect 400 2308 404 2309
rect 174 2269 246 2277
rect 295 2274 300 2308
rect 324 2274 329 2308
rect 224 2239 226 2255
rect 196 2231 226 2239
rect 332 2237 336 2305
rect 367 2274 438 2308
rect 400 2267 404 2274
rect 454 2261 504 2263
rect 494 2257 548 2261
rect 494 2252 514 2257
rect 504 2237 506 2252
rect 196 2227 232 2231
rect 196 2197 204 2227
rect 216 2197 232 2227
rect 400 2229 404 2237
rect 107 2157 119 2163
rect 109 2129 119 2157
rect 129 2129 149 2163
rect 174 2159 181 2189
rect 224 2150 226 2197
rect 256 2189 328 2197
rect 332 2195 336 2225
rect 400 2195 408 2229
rect 434 2195 438 2229
rect 498 2227 506 2237
rect 514 2227 515 2247
rect 504 2211 506 2227
rect 525 2218 528 2252
rect 547 2227 548 2247
rect 557 2227 564 2237
rect 514 2211 530 2217
rect 532 2211 548 2217
rect 278 2159 305 2170
rect 42 2037 46 2071
rect 72 2037 76 2071
rect 38 1999 80 2000
rect 42 1958 76 1992
rect 79 1958 113 1992
rect 42 1879 46 1913
rect 72 1879 76 1913
rect -25 1842 25 1844
rect -8 1834 14 1841
rect -8 1833 17 1834
rect 25 1833 27 1842
rect -12 1826 38 1833
rect -12 1825 34 1826
rect -12 1821 8 1825
rect 0 1809 8 1821
rect 14 1809 34 1825
rect 0 1808 34 1809
rect 0 1801 38 1808
rect 14 1800 17 1801
rect 25 1792 27 1801
rect 42 1772 45 1862
rect 71 1831 80 1859
rect 69 1793 80 1831
rect 144 1821 148 2129
rect 196 2116 204 2150
rect 216 2116 232 2150
rect 244 2146 257 2150
rect 300 2146 308 2159
rect 332 2157 342 2195
rect 400 2187 404 2195
rect 336 2147 342 2157
rect 244 2122 291 2146
rect 244 2116 257 2122
rect 224 2069 226 2116
rect 278 2112 291 2122
rect 300 2122 329 2146
rect 332 2137 342 2147
rect 400 2147 409 2175
rect 562 2158 612 2160
rect 466 2149 497 2157
rect 565 2149 596 2157
rect 300 2112 321 2122
rect 300 2106 308 2112
rect 289 2096 308 2106
rect 196 2039 204 2069
rect 216 2039 232 2069
rect 196 2035 232 2039
rect 196 2027 226 2035
rect 300 2027 308 2096
rect 332 2103 351 2137
rect 361 2109 381 2137
rect 361 2103 375 2109
rect 400 2103 411 2147
rect 442 2142 500 2149
rect 466 2141 500 2142
rect 565 2141 599 2149
rect 497 2125 500 2141
rect 596 2125 599 2141
rect 466 2124 500 2125
rect 442 2117 500 2124
rect 565 2117 599 2125
rect 612 2108 614 2158
rect 332 2079 342 2103
rect 336 2067 342 2079
rect 224 2011 226 2027
rect 332 1999 342 2067
rect 400 2071 404 2079
rect 400 2037 408 2071
rect 434 2037 438 2071
rect 454 2055 504 2057
rect 504 2039 506 2055
rect 514 2049 530 2055
rect 532 2049 548 2055
rect 525 2039 548 2048
rect 400 2029 404 2037
rect 498 2029 506 2039
rect 504 2005 506 2029
rect 514 2019 515 2039
rect 525 2014 528 2039
rect 547 2019 548 2039
rect 557 2029 564 2039
rect 514 2005 548 2009
rect 151 1958 156 1992
rect 174 1989 246 1997
rect 256 1989 328 1997
rect 336 1991 342 1999
rect 400 1994 404 1999
rect 180 1961 185 1989
rect 174 1953 246 1961
rect 256 1953 328 1961
rect 332 1959 336 1989
rect 400 1960 438 1994
rect 224 1923 226 1939
rect 196 1915 226 1923
rect 196 1911 232 1915
rect 196 1881 204 1911
rect 216 1881 232 1911
rect 224 1834 226 1881
rect 300 1854 308 1923
rect 332 1921 342 1959
rect 400 1951 404 1960
rect 454 1945 504 1947
rect 494 1941 548 1945
rect 494 1936 514 1941
rect 504 1921 506 1936
rect 336 1909 342 1921
rect 289 1844 308 1854
rect 300 1838 308 1844
rect 332 1875 342 1909
rect 400 1913 404 1921
rect 400 1879 408 1913
rect 434 1879 438 1913
rect 498 1911 506 1921
rect 514 1911 515 1931
rect 504 1895 506 1911
rect 525 1902 528 1936
rect 547 1911 548 1931
rect 557 1911 564 1921
rect 514 1895 530 1901
rect 532 1895 548 1901
rect 332 1847 373 1875
rect 332 1841 351 1847
rect 107 1787 119 1821
rect 129 1787 149 1821
rect 196 1800 204 1834
rect 216 1800 232 1834
rect 244 1828 257 1834
rect 278 1828 291 1838
rect 244 1804 291 1828
rect 300 1828 321 1838
rect 336 1831 351 1841
rect 300 1804 329 1828
rect 332 1813 351 1831
rect 361 1841 375 1847
rect 400 1841 411 1879
rect 562 1842 612 1844
rect 361 1813 381 1841
rect 400 1813 409 1841
rect 466 1833 497 1841
rect 565 1833 596 1841
rect 442 1826 500 1833
rect 466 1825 500 1826
rect 565 1825 599 1833
rect 244 1800 257 1804
rect 42 1721 46 1755
rect 72 1721 76 1755
rect 42 1674 76 1678
rect 42 1659 46 1674
rect 72 1659 76 1674
rect 38 1641 80 1659
rect 16 1635 102 1641
rect 144 1635 148 1787
rect 174 1763 181 1791
rect 224 1753 226 1800
rect 300 1791 308 1804
rect 278 1780 305 1791
rect 332 1763 342 1813
rect 400 1793 404 1813
rect 497 1809 500 1825
rect 596 1809 599 1825
rect 466 1808 500 1809
rect 442 1801 500 1808
rect 565 1801 599 1809
rect 612 1792 614 1842
rect 256 1753 328 1761
rect 336 1755 342 1763
rect 400 1755 404 1763
rect 196 1723 204 1753
rect 216 1723 232 1753
rect 196 1719 232 1723
rect 196 1711 226 1719
rect 224 1695 226 1711
rect 332 1683 336 1751
rect 400 1721 408 1755
rect 434 1721 438 1755
rect 454 1739 504 1741
rect 504 1723 506 1739
rect 514 1733 530 1739
rect 532 1733 548 1739
rect 525 1723 548 1732
rect 400 1713 404 1721
rect 498 1713 506 1723
rect 504 1689 506 1713
rect 514 1703 515 1723
rect 525 1698 528 1723
rect 547 1703 548 1723
rect 557 1713 564 1723
rect 514 1689 548 1693
rect 400 1683 442 1684
rect 174 1673 246 1681
rect 400 1676 404 1683
rect 295 1642 300 1676
rect 324 1642 329 1676
rect 367 1659 438 1676
rect 367 1642 442 1659
rect 400 1641 442 1642
rect 378 1635 464 1641
rect 38 1619 80 1635
rect 400 1619 442 1635
rect -25 1605 25 1607
rect 42 1605 76 1619
rect 404 1605 438 1619
rect 455 1605 505 1607
rect 557 1605 607 1607
rect 16 1597 102 1605
rect 378 1597 464 1605
rect 8 1563 17 1597
rect 18 1595 51 1597
rect 80 1595 100 1597
rect 18 1563 100 1595
rect 380 1595 404 1597
rect 429 1595 438 1597
rect 442 1595 462 1597
rect 16 1555 102 1563
rect 42 1539 76 1555
rect 16 1519 38 1525
rect 42 1516 76 1520
rect 80 1519 102 1525
rect 42 1486 46 1516
rect 72 1486 76 1516
rect 42 1405 46 1439
rect 72 1405 76 1439
rect -25 1368 25 1370
rect -8 1360 14 1367
rect -8 1359 17 1360
rect 25 1359 27 1368
rect -12 1352 38 1359
rect -12 1351 34 1352
rect -12 1347 8 1351
rect 0 1335 8 1347
rect 14 1335 34 1351
rect 0 1334 34 1335
rect 0 1327 38 1334
rect 14 1326 17 1327
rect 25 1318 27 1327
rect 42 1298 45 1388
rect 69 1373 80 1405
rect 107 1373 143 1401
rect 144 1373 148 1593
rect 332 1525 336 1593
rect 380 1563 462 1595
rect 463 1563 472 1597
rect 480 1563 497 1597
rect 378 1555 464 1563
rect 505 1555 507 1605
rect 514 1563 548 1597
rect 565 1563 582 1597
rect 607 1555 609 1605
rect 404 1539 438 1555
rect 400 1525 442 1526
rect 378 1519 404 1525
rect 442 1519 464 1525
rect 400 1518 404 1519
rect 174 1479 246 1487
rect 295 1484 300 1518
rect 324 1484 329 1518
rect 224 1449 226 1465
rect 196 1441 226 1449
rect 332 1447 336 1515
rect 367 1484 438 1518
rect 400 1477 404 1484
rect 454 1471 504 1473
rect 494 1467 548 1471
rect 494 1462 514 1467
rect 504 1447 506 1462
rect 196 1437 232 1441
rect 196 1407 204 1437
rect 216 1407 232 1437
rect 400 1439 404 1447
rect 107 1367 119 1373
rect 109 1339 119 1367
rect 129 1339 149 1373
rect 174 1369 181 1399
rect 224 1360 226 1407
rect 256 1399 328 1407
rect 332 1405 336 1435
rect 400 1405 408 1439
rect 434 1405 438 1439
rect 498 1437 506 1447
rect 514 1437 515 1457
rect 504 1421 506 1437
rect 525 1428 528 1462
rect 547 1437 548 1457
rect 557 1437 564 1447
rect 514 1421 530 1427
rect 532 1421 548 1427
rect 278 1369 305 1380
rect 42 1247 46 1281
rect 72 1247 76 1281
rect 38 1209 80 1210
rect 42 1168 76 1202
rect 79 1168 113 1202
rect 42 1089 46 1123
rect 72 1089 76 1123
rect -25 1052 25 1054
rect -8 1044 14 1051
rect -8 1043 17 1044
rect 25 1043 27 1052
rect -12 1036 38 1043
rect -12 1035 34 1036
rect -12 1031 8 1035
rect 0 1019 8 1031
rect 14 1019 34 1035
rect 0 1018 34 1019
rect 0 1011 38 1018
rect 14 1010 17 1011
rect 25 1002 27 1011
rect 42 982 45 1072
rect 71 1041 80 1069
rect 69 1003 80 1041
rect 144 1031 148 1339
rect 196 1326 204 1360
rect 216 1326 232 1360
rect 244 1356 257 1360
rect 300 1356 308 1369
rect 332 1367 342 1405
rect 400 1397 404 1405
rect 336 1357 342 1367
rect 244 1332 291 1356
rect 244 1326 257 1332
rect 224 1279 226 1326
rect 278 1322 291 1332
rect 300 1332 329 1356
rect 332 1347 342 1357
rect 400 1357 409 1385
rect 562 1368 612 1370
rect 466 1359 497 1367
rect 565 1359 596 1367
rect 300 1322 321 1332
rect 300 1316 308 1322
rect 289 1306 308 1316
rect 196 1249 204 1279
rect 216 1249 232 1279
rect 196 1245 232 1249
rect 196 1237 226 1245
rect 300 1237 308 1306
rect 332 1313 351 1347
rect 361 1319 381 1347
rect 361 1313 375 1319
rect 400 1313 411 1357
rect 442 1352 500 1359
rect 466 1351 500 1352
rect 565 1351 599 1359
rect 497 1335 500 1351
rect 596 1335 599 1351
rect 466 1334 500 1335
rect 442 1327 500 1334
rect 565 1327 599 1335
rect 612 1318 614 1368
rect 332 1289 342 1313
rect 336 1277 342 1289
rect 224 1221 226 1237
rect 332 1209 342 1277
rect 400 1281 404 1289
rect 400 1247 408 1281
rect 434 1247 438 1281
rect 454 1265 504 1267
rect 504 1249 506 1265
rect 514 1259 530 1265
rect 532 1259 548 1265
rect 525 1249 548 1258
rect 400 1239 404 1247
rect 498 1239 506 1249
rect 504 1215 506 1239
rect 514 1229 515 1249
rect 525 1224 528 1249
rect 547 1229 548 1249
rect 557 1239 564 1249
rect 514 1215 548 1219
rect 151 1168 156 1202
rect 174 1199 246 1207
rect 256 1199 328 1207
rect 336 1201 342 1209
rect 400 1204 404 1209
rect 180 1171 185 1199
rect 174 1163 246 1171
rect 256 1163 328 1171
rect 332 1169 336 1199
rect 400 1170 438 1204
rect 224 1133 226 1149
rect 196 1125 226 1133
rect 196 1121 232 1125
rect 196 1091 204 1121
rect 216 1091 232 1121
rect 224 1044 226 1091
rect 300 1064 308 1133
rect 332 1131 342 1169
rect 400 1161 404 1170
rect 454 1155 504 1157
rect 494 1151 548 1155
rect 494 1146 514 1151
rect 504 1131 506 1146
rect 336 1119 342 1131
rect 289 1054 308 1064
rect 300 1048 308 1054
rect 332 1085 342 1119
rect 400 1123 404 1131
rect 400 1089 408 1123
rect 434 1089 438 1123
rect 498 1121 506 1131
rect 514 1121 515 1141
rect 504 1105 506 1121
rect 525 1112 528 1146
rect 547 1121 548 1141
rect 557 1121 564 1131
rect 514 1105 530 1111
rect 532 1105 548 1111
rect 332 1057 373 1085
rect 332 1051 351 1057
rect 107 997 119 1031
rect 129 997 149 1031
rect 196 1010 204 1044
rect 216 1010 232 1044
rect 244 1038 257 1044
rect 278 1038 291 1048
rect 244 1014 291 1038
rect 300 1038 321 1048
rect 336 1041 351 1051
rect 300 1014 329 1038
rect 332 1023 351 1041
rect 361 1051 375 1057
rect 400 1051 411 1089
rect 562 1052 612 1054
rect 361 1023 381 1051
rect 400 1023 409 1051
rect 466 1043 497 1051
rect 565 1043 596 1051
rect 442 1036 500 1043
rect 466 1035 500 1036
rect 565 1035 599 1043
rect 244 1010 257 1014
rect 42 931 46 965
rect 72 931 76 965
rect 42 884 76 888
rect 42 869 46 884
rect 72 869 76 884
rect 38 851 80 869
rect 16 845 102 851
rect 144 845 148 997
rect 174 973 181 1001
rect 224 963 226 1010
rect 300 1001 308 1014
rect 278 990 305 1001
rect 332 973 342 1023
rect 400 1003 404 1023
rect 497 1019 500 1035
rect 596 1019 599 1035
rect 466 1018 500 1019
rect 442 1011 500 1018
rect 565 1011 599 1019
rect 612 1002 614 1052
rect 256 963 328 971
rect 336 965 342 973
rect 400 965 404 973
rect 196 933 204 963
rect 216 933 232 963
rect 196 929 232 933
rect 196 921 226 929
rect 224 905 226 921
rect 332 893 336 961
rect 400 931 408 965
rect 434 931 438 965
rect 454 949 504 951
rect 504 933 506 949
rect 514 943 530 949
rect 532 943 548 949
rect 525 933 548 942
rect 400 923 404 931
rect 498 923 506 933
rect 504 899 506 923
rect 514 913 515 933
rect 525 908 528 933
rect 547 913 548 933
rect 557 923 564 933
rect 514 899 548 903
rect 400 893 442 894
rect 174 883 246 891
rect 400 886 404 893
rect 295 852 300 886
rect 324 852 329 886
rect 367 869 438 886
rect 367 852 442 869
rect 400 851 442 852
rect 378 845 464 851
rect 38 829 80 845
rect 400 829 442 845
rect -25 815 25 817
rect 42 815 76 829
rect 404 815 438 829
rect 455 815 505 817
rect 557 815 607 817
rect 16 807 102 815
rect 378 807 464 815
rect 8 773 17 807
rect 18 805 51 807
rect 80 805 100 807
rect 18 773 100 805
rect 380 805 404 807
rect 429 805 438 807
rect 442 805 462 807
rect 16 765 102 773
rect 42 749 76 765
rect 16 729 38 735
rect 42 726 76 730
rect 80 729 102 735
rect 42 696 46 726
rect 72 696 76 726
rect 69 583 80 621
rect 107 583 143 611
rect 144 583 148 803
rect 332 735 336 803
rect 380 773 462 805
rect 463 773 472 807
rect 480 773 497 807
rect 378 765 464 773
rect 505 765 507 815
rect 514 773 548 807
rect 565 773 582 807
rect 607 765 609 815
rect 404 749 438 765
rect 400 735 442 736
rect 378 729 404 735
rect 442 729 464 735
rect 400 728 404 729
rect 295 694 300 728
rect 324 694 329 728
rect 332 657 336 725
rect 367 694 438 728
rect 400 687 404 694
rect 454 681 504 683
rect 494 677 548 681
rect 494 672 514 677
rect 504 657 506 672
rect -25 578 25 580
rect -8 569 17 577
rect 25 569 27 578
rect 107 577 119 583
rect -12 562 38 569
rect -12 561 34 562
rect -12 557 8 561
rect 0 545 8 557
rect 17 545 34 561
rect 109 549 119 577
rect 129 549 149 583
rect 174 579 181 609
rect 332 577 336 645
rect 400 607 404 657
rect 498 647 506 657
rect 514 647 515 667
rect 504 631 506 647
rect 525 638 528 672
rect 547 647 548 667
rect 557 647 564 657
rect 514 631 530 637
rect 532 631 548 637
rect 400 567 409 595
rect 562 578 612 580
rect 463 569 497 577
rect 0 544 34 545
rect 0 537 38 544
rect 25 528 27 537
rect 42 420 76 429
rect 38 419 80 420
rect 42 395 76 419
rect 79 395 113 412
rect 144 395 148 549
rect 332 499 336 567
rect 341 523 351 557
rect 361 529 381 557
rect 361 523 375 529
rect 400 523 411 567
rect 442 562 497 569
rect 463 561 497 562
rect 565 569 596 577
rect 565 561 599 569
rect 596 545 599 561
rect 463 544 497 545
rect 442 537 497 544
rect 565 537 599 545
rect 612 528 614 578
rect 332 419 336 487
rect 400 449 404 499
rect 454 475 504 477
rect 504 459 506 475
rect 514 469 530 475
rect 532 469 548 475
rect 525 459 548 468
rect 498 449 506 459
rect 404 419 438 429
rect 504 425 506 449
rect 514 439 515 459
rect 525 434 528 459
rect 547 439 548 459
rect 557 449 564 459
rect 514 425 548 429
rect 38 378 113 395
rect 151 378 156 412
rect 180 378 185 412
rect 400 411 438 419
rect 388 410 454 411
rect 400 403 408 410
rect 434 403 438 410
rect 400 395 438 403
rect 38 369 80 378
rect 400 369 442 395
<< metal1 >>
rect 78 0 114 102700
rect 150 0 186 102700
rect 222 101989 258 102330
rect 222 101199 258 101831
rect 222 100409 258 101041
rect 222 99619 258 100251
rect 222 98829 258 99461
rect 222 98039 258 98671
rect 222 97249 258 97881
rect 222 96459 258 97091
rect 222 95669 258 96301
rect 222 94879 258 95511
rect 222 94089 258 94721
rect 222 93299 258 93931
rect 222 92509 258 93141
rect 222 91719 258 92351
rect 222 90929 258 91561
rect 222 90139 258 90771
rect 222 89349 258 89981
rect 222 88559 258 89191
rect 222 87769 258 88401
rect 222 86979 258 87611
rect 222 86189 258 86821
rect 222 85399 258 86031
rect 222 84609 258 85241
rect 222 83819 258 84451
rect 222 83029 258 83661
rect 222 82239 258 82871
rect 222 81449 258 82081
rect 222 80659 258 81291
rect 222 79869 258 80501
rect 222 79079 258 79711
rect 222 78289 258 78921
rect 222 77499 258 78131
rect 222 76709 258 77341
rect 222 75919 258 76551
rect 222 75129 258 75761
rect 222 74339 258 74971
rect 222 73549 258 74181
rect 222 72759 258 73391
rect 222 71969 258 72601
rect 222 71179 258 71811
rect 222 70389 258 71021
rect 222 69599 258 70231
rect 222 68809 258 69441
rect 222 68019 258 68651
rect 222 67229 258 67861
rect 222 66439 258 67071
rect 222 65649 258 66281
rect 222 64859 258 65491
rect 222 64069 258 64701
rect 222 63279 258 63911
rect 222 62489 258 63121
rect 222 61699 258 62331
rect 222 60909 258 61541
rect 222 60119 258 60751
rect 222 59329 258 59961
rect 222 58539 258 59171
rect 222 57749 258 58381
rect 222 56959 258 57591
rect 222 56169 258 56801
rect 222 55379 258 56011
rect 222 54589 258 55221
rect 222 53799 258 54431
rect 222 53009 258 53641
rect 222 52219 258 52851
rect 222 51429 258 52061
rect 222 50639 258 51271
rect 222 49849 258 50481
rect 222 49059 258 49691
rect 222 48269 258 48901
rect 222 47479 258 48111
rect 222 46689 258 47321
rect 222 45899 258 46531
rect 222 45109 258 45741
rect 222 44319 258 44951
rect 222 43529 258 44161
rect 222 42739 258 43371
rect 222 41949 258 42581
rect 222 41159 258 41791
rect 222 40369 258 41001
rect 222 39579 258 40211
rect 222 38789 258 39421
rect 222 37999 258 38631
rect 222 37209 258 37841
rect 222 36419 258 37051
rect 222 35629 258 36261
rect 222 34839 258 35471
rect 222 34049 258 34681
rect 222 33259 258 33891
rect 222 32469 258 33101
rect 222 31679 258 32311
rect 222 30889 258 31521
rect 222 30099 258 30731
rect 222 29309 258 29941
rect 222 28519 258 29151
rect 222 27729 258 28361
rect 222 26939 258 27571
rect 222 26149 258 26781
rect 222 25359 258 25991
rect 222 24569 258 25201
rect 222 23779 258 24411
rect 222 22989 258 23621
rect 222 22199 258 22831
rect 222 21409 258 22041
rect 222 20619 258 21251
rect 222 19829 258 20461
rect 222 19039 258 19671
rect 222 18249 258 18881
rect 222 17459 258 18091
rect 222 16669 258 17301
rect 222 15879 258 16511
rect 222 15089 258 15721
rect 222 14299 258 14931
rect 222 13509 258 14141
rect 222 12719 258 13351
rect 222 11929 258 12561
rect 222 11139 258 11771
rect 222 10349 258 10981
rect 222 9559 258 10191
rect 222 8769 258 9401
rect 222 7979 258 8611
rect 222 7189 258 7821
rect 222 6399 258 7031
rect 222 5609 258 6241
rect 222 4819 258 5451
rect 222 4029 258 4661
rect 222 3239 258 3871
rect 222 2449 258 3081
rect 222 1659 258 2291
rect 222 869 258 1501
rect 222 370 258 711
rect 294 0 330 102700
rect 366 0 402 102700
<< metal2 >>
rect 0 102233 624 102281
rect 186 102109 294 102185
rect 0 102013 624 102061
rect 186 101855 294 101965
rect 0 101759 624 101807
rect 186 101635 294 101711
rect 0 101539 624 101587
rect 0 101443 624 101491
rect 186 101319 294 101395
rect 0 101223 624 101271
rect 186 101065 294 101175
rect 0 100969 624 101017
rect 186 100845 294 100921
rect 0 100749 624 100797
rect 0 100653 624 100701
rect 186 100529 294 100605
rect 0 100433 624 100481
rect 186 100275 294 100385
rect 0 100179 624 100227
rect 186 100055 294 100131
rect 0 99959 624 100007
rect 0 99863 624 99911
rect 186 99739 294 99815
rect 0 99643 624 99691
rect 186 99485 294 99595
rect 0 99389 624 99437
rect 186 99265 294 99341
rect 0 99169 624 99217
rect 0 99073 624 99121
rect 186 98949 294 99025
rect 0 98853 624 98901
rect 186 98695 294 98805
rect 0 98599 624 98647
rect 186 98475 294 98551
rect 0 98379 624 98427
rect 0 98283 624 98331
rect 186 98159 294 98235
rect 0 98063 624 98111
rect 186 97905 294 98015
rect 0 97809 624 97857
rect 186 97685 294 97761
rect 0 97589 624 97637
rect 0 97493 624 97541
rect 186 97369 294 97445
rect 0 97273 624 97321
rect 186 97115 294 97225
rect 0 97019 624 97067
rect 186 96895 294 96971
rect 0 96799 624 96847
rect 0 96703 624 96751
rect 186 96579 294 96655
rect 0 96483 624 96531
rect 186 96325 294 96435
rect 0 96229 624 96277
rect 186 96105 294 96181
rect 0 96009 624 96057
rect 0 95913 624 95961
rect 186 95789 294 95865
rect 0 95693 624 95741
rect 186 95535 294 95645
rect 0 95439 624 95487
rect 186 95315 294 95391
rect 0 95219 624 95267
rect 0 95123 624 95171
rect 186 94999 294 95075
rect 0 94903 624 94951
rect 186 94745 294 94855
rect 0 94649 624 94697
rect 186 94525 294 94601
rect 0 94429 624 94477
rect 0 94333 624 94381
rect 186 94209 294 94285
rect 0 94113 624 94161
rect 186 93955 294 94065
rect 0 93859 624 93907
rect 186 93735 294 93811
rect 0 93639 624 93687
rect 0 93543 624 93591
rect 186 93419 294 93495
rect 0 93323 624 93371
rect 186 93165 294 93275
rect 0 93069 624 93117
rect 186 92945 294 93021
rect 0 92849 624 92897
rect 0 92753 624 92801
rect 186 92629 294 92705
rect 0 92533 624 92581
rect 186 92375 294 92485
rect 0 92279 624 92327
rect 186 92155 294 92231
rect 0 92059 624 92107
rect 0 91963 624 92011
rect 186 91839 294 91915
rect 0 91743 624 91791
rect 186 91585 294 91695
rect 0 91489 624 91537
rect 186 91365 294 91441
rect 0 91269 624 91317
rect 0 91173 624 91221
rect 186 91049 294 91125
rect 0 90953 624 91001
rect 186 90795 294 90905
rect 0 90699 624 90747
rect 186 90575 294 90651
rect 0 90479 624 90527
rect 0 90383 624 90431
rect 186 90259 294 90335
rect 0 90163 624 90211
rect 186 90005 294 90115
rect 0 89909 624 89957
rect 186 89785 294 89861
rect 0 89689 624 89737
rect 0 89593 624 89641
rect 186 89469 294 89545
rect 0 89373 624 89421
rect 186 89215 294 89325
rect 0 89119 624 89167
rect 186 88995 294 89071
rect 0 88899 624 88947
rect 0 88803 624 88851
rect 186 88679 294 88755
rect 0 88583 624 88631
rect 186 88425 294 88535
rect 0 88329 624 88377
rect 186 88205 294 88281
rect 0 88109 624 88157
rect 0 88013 624 88061
rect 186 87889 294 87965
rect 0 87793 624 87841
rect 186 87635 294 87745
rect 0 87539 624 87587
rect 186 87415 294 87491
rect 0 87319 624 87367
rect 0 87223 624 87271
rect 186 87099 294 87175
rect 0 87003 624 87051
rect 186 86845 294 86955
rect 0 86749 624 86797
rect 186 86625 294 86701
rect 0 86529 624 86577
rect 0 86433 624 86481
rect 186 86309 294 86385
rect 0 86213 624 86261
rect 186 86055 294 86165
rect 0 85959 624 86007
rect 186 85835 294 85911
rect 0 85739 624 85787
rect 0 85643 624 85691
rect 186 85519 294 85595
rect 0 85423 624 85471
rect 186 85265 294 85375
rect 0 85169 624 85217
rect 186 85045 294 85121
rect 0 84949 624 84997
rect 0 84853 624 84901
rect 186 84729 294 84805
rect 0 84633 624 84681
rect 186 84475 294 84585
rect 0 84379 624 84427
rect 186 84255 294 84331
rect 0 84159 624 84207
rect 0 84063 624 84111
rect 186 83939 294 84015
rect 0 83843 624 83891
rect 186 83685 294 83795
rect 0 83589 624 83637
rect 186 83465 294 83541
rect 0 83369 624 83417
rect 0 83273 624 83321
rect 186 83149 294 83225
rect 0 83053 624 83101
rect 186 82895 294 83005
rect 0 82799 624 82847
rect 186 82675 294 82751
rect 0 82579 624 82627
rect 0 82483 624 82531
rect 186 82359 294 82435
rect 0 82263 624 82311
rect 186 82105 294 82215
rect 0 82009 624 82057
rect 186 81885 294 81961
rect 0 81789 624 81837
rect 0 81693 624 81741
rect 186 81569 294 81645
rect 0 81473 624 81521
rect 186 81315 294 81425
rect 0 81219 624 81267
rect 186 81095 294 81171
rect 0 80999 624 81047
rect 0 80903 624 80951
rect 186 80779 294 80855
rect 0 80683 624 80731
rect 186 80525 294 80635
rect 0 80429 624 80477
rect 186 80305 294 80381
rect 0 80209 624 80257
rect 0 80113 624 80161
rect 186 79989 294 80065
rect 0 79893 624 79941
rect 186 79735 294 79845
rect 0 79639 624 79687
rect 186 79515 294 79591
rect 0 79419 624 79467
rect 0 79323 624 79371
rect 186 79199 294 79275
rect 0 79103 624 79151
rect 186 78945 294 79055
rect 0 78849 624 78897
rect 186 78725 294 78801
rect 0 78629 624 78677
rect 0 78533 624 78581
rect 186 78409 294 78485
rect 0 78313 624 78361
rect 186 78155 294 78265
rect 0 78059 624 78107
rect 186 77935 294 78011
rect 0 77839 624 77887
rect 0 77743 624 77791
rect 186 77619 294 77695
rect 0 77523 624 77571
rect 186 77365 294 77475
rect 0 77269 624 77317
rect 186 77145 294 77221
rect 0 77049 624 77097
rect 0 76953 624 77001
rect 186 76829 294 76905
rect 0 76733 624 76781
rect 186 76575 294 76685
rect 0 76479 624 76527
rect 186 76355 294 76431
rect 0 76259 624 76307
rect 0 76163 624 76211
rect 186 76039 294 76115
rect 0 75943 624 75991
rect 186 75785 294 75895
rect 0 75689 624 75737
rect 186 75565 294 75641
rect 0 75469 624 75517
rect 0 75373 624 75421
rect 186 75249 294 75325
rect 0 75153 624 75201
rect 186 74995 294 75105
rect 0 74899 624 74947
rect 186 74775 294 74851
rect 0 74679 624 74727
rect 0 74583 624 74631
rect 186 74459 294 74535
rect 0 74363 624 74411
rect 186 74205 294 74315
rect 0 74109 624 74157
rect 186 73985 294 74061
rect 0 73889 624 73937
rect 0 73793 624 73841
rect 186 73669 294 73745
rect 0 73573 624 73621
rect 186 73415 294 73525
rect 0 73319 624 73367
rect 186 73195 294 73271
rect 0 73099 624 73147
rect 0 73003 624 73051
rect 186 72879 294 72955
rect 0 72783 624 72831
rect 186 72625 294 72735
rect 0 72529 624 72577
rect 186 72405 294 72481
rect 0 72309 624 72357
rect 0 72213 624 72261
rect 186 72089 294 72165
rect 0 71993 624 72041
rect 186 71835 294 71945
rect 0 71739 624 71787
rect 186 71615 294 71691
rect 0 71519 624 71567
rect 0 71423 624 71471
rect 186 71299 294 71375
rect 0 71203 624 71251
rect 186 71045 294 71155
rect 0 70949 624 70997
rect 186 70825 294 70901
rect 0 70729 624 70777
rect 0 70633 624 70681
rect 186 70509 294 70585
rect 0 70413 624 70461
rect 186 70255 294 70365
rect 0 70159 624 70207
rect 186 70035 294 70111
rect 0 69939 624 69987
rect 0 69843 624 69891
rect 186 69719 294 69795
rect 0 69623 624 69671
rect 186 69465 294 69575
rect 0 69369 624 69417
rect 186 69245 294 69321
rect 0 69149 624 69197
rect 0 69053 624 69101
rect 186 68929 294 69005
rect 0 68833 624 68881
rect 186 68675 294 68785
rect 0 68579 624 68627
rect 186 68455 294 68531
rect 0 68359 624 68407
rect 0 68263 624 68311
rect 186 68139 294 68215
rect 0 68043 624 68091
rect 186 67885 294 67995
rect 0 67789 624 67837
rect 186 67665 294 67741
rect 0 67569 624 67617
rect 0 67473 624 67521
rect 186 67349 294 67425
rect 0 67253 624 67301
rect 186 67095 294 67205
rect 0 66999 624 67047
rect 186 66875 294 66951
rect 0 66779 624 66827
rect 0 66683 624 66731
rect 186 66559 294 66635
rect 0 66463 624 66511
rect 186 66305 294 66415
rect 0 66209 624 66257
rect 186 66085 294 66161
rect 0 65989 624 66037
rect 0 65893 624 65941
rect 186 65769 294 65845
rect 0 65673 624 65721
rect 186 65515 294 65625
rect 0 65419 624 65467
rect 186 65295 294 65371
rect 0 65199 624 65247
rect 0 65103 624 65151
rect 186 64979 294 65055
rect 0 64883 624 64931
rect 186 64725 294 64835
rect 0 64629 624 64677
rect 186 64505 294 64581
rect 0 64409 624 64457
rect 0 64313 624 64361
rect 186 64189 294 64265
rect 0 64093 624 64141
rect 186 63935 294 64045
rect 0 63839 624 63887
rect 186 63715 294 63791
rect 0 63619 624 63667
rect 0 63523 624 63571
rect 186 63399 294 63475
rect 0 63303 624 63351
rect 186 63145 294 63255
rect 0 63049 624 63097
rect 186 62925 294 63001
rect 0 62829 624 62877
rect 0 62733 624 62781
rect 186 62609 294 62685
rect 0 62513 624 62561
rect 186 62355 294 62465
rect 0 62259 624 62307
rect 186 62135 294 62211
rect 0 62039 624 62087
rect 0 61943 624 61991
rect 186 61819 294 61895
rect 0 61723 624 61771
rect 186 61565 294 61675
rect 0 61469 624 61517
rect 186 61345 294 61421
rect 0 61249 624 61297
rect 0 61153 624 61201
rect 186 61029 294 61105
rect 0 60933 624 60981
rect 186 60775 294 60885
rect 0 60679 624 60727
rect 186 60555 294 60631
rect 0 60459 624 60507
rect 0 60363 624 60411
rect 186 60239 294 60315
rect 0 60143 624 60191
rect 186 59985 294 60095
rect 0 59889 624 59937
rect 186 59765 294 59841
rect 0 59669 624 59717
rect 0 59573 624 59621
rect 186 59449 294 59525
rect 0 59353 624 59401
rect 186 59195 294 59305
rect 0 59099 624 59147
rect 186 58975 294 59051
rect 0 58879 624 58927
rect 0 58783 624 58831
rect 186 58659 294 58735
rect 0 58563 624 58611
rect 186 58405 294 58515
rect 0 58309 624 58357
rect 186 58185 294 58261
rect 0 58089 624 58137
rect 0 57993 624 58041
rect 186 57869 294 57945
rect 0 57773 624 57821
rect 186 57615 294 57725
rect 0 57519 624 57567
rect 186 57395 294 57471
rect 0 57299 624 57347
rect 0 57203 624 57251
rect 186 57079 294 57155
rect 0 56983 624 57031
rect 186 56825 294 56935
rect 0 56729 624 56777
rect 186 56605 294 56681
rect 0 56509 624 56557
rect 0 56413 624 56461
rect 186 56289 294 56365
rect 0 56193 624 56241
rect 186 56035 294 56145
rect 0 55939 624 55987
rect 186 55815 294 55891
rect 0 55719 624 55767
rect 0 55623 624 55671
rect 186 55499 294 55575
rect 0 55403 624 55451
rect 186 55245 294 55355
rect 0 55149 624 55197
rect 186 55025 294 55101
rect 0 54929 624 54977
rect 0 54833 624 54881
rect 186 54709 294 54785
rect 0 54613 624 54661
rect 186 54455 294 54565
rect 0 54359 624 54407
rect 186 54235 294 54311
rect 0 54139 624 54187
rect 0 54043 624 54091
rect 186 53919 294 53995
rect 0 53823 624 53871
rect 186 53665 294 53775
rect 0 53569 624 53617
rect 186 53445 294 53521
rect 0 53349 624 53397
rect 0 53253 624 53301
rect 186 53129 294 53205
rect 0 53033 624 53081
rect 186 52875 294 52985
rect 0 52779 624 52827
rect 186 52655 294 52731
rect 0 52559 624 52607
rect 0 52463 624 52511
rect 186 52339 294 52415
rect 0 52243 624 52291
rect 186 52085 294 52195
rect 0 51989 624 52037
rect 186 51865 294 51941
rect 0 51769 624 51817
rect 0 51673 624 51721
rect 186 51549 294 51625
rect 0 51453 624 51501
rect 186 51295 294 51405
rect 0 51199 624 51247
rect 186 51075 294 51151
rect 0 50979 624 51027
rect 0 50883 624 50931
rect 186 50759 294 50835
rect 0 50663 624 50711
rect 186 50505 294 50615
rect 0 50409 624 50457
rect 186 50285 294 50361
rect 0 50189 624 50237
rect 0 50093 624 50141
rect 186 49969 294 50045
rect 0 49873 624 49921
rect 186 49715 294 49825
rect 0 49619 624 49667
rect 186 49495 294 49571
rect 0 49399 624 49447
rect 0 49303 624 49351
rect 186 49179 294 49255
rect 0 49083 624 49131
rect 186 48925 294 49035
rect 0 48829 624 48877
rect 186 48705 294 48781
rect 0 48609 624 48657
rect 0 48513 624 48561
rect 186 48389 294 48465
rect 0 48293 624 48341
rect 186 48135 294 48245
rect 0 48039 624 48087
rect 186 47915 294 47991
rect 0 47819 624 47867
rect 0 47723 624 47771
rect 186 47599 294 47675
rect 0 47503 624 47551
rect 186 47345 294 47455
rect 0 47249 624 47297
rect 186 47125 294 47201
rect 0 47029 624 47077
rect 0 46933 624 46981
rect 186 46809 294 46885
rect 0 46713 624 46761
rect 186 46555 294 46665
rect 0 46459 624 46507
rect 186 46335 294 46411
rect 0 46239 624 46287
rect 0 46143 624 46191
rect 186 46019 294 46095
rect 0 45923 624 45971
rect 186 45765 294 45875
rect 0 45669 624 45717
rect 186 45545 294 45621
rect 0 45449 624 45497
rect 0 45353 624 45401
rect 186 45229 294 45305
rect 0 45133 624 45181
rect 186 44975 294 45085
rect 0 44879 624 44927
rect 186 44755 294 44831
rect 0 44659 624 44707
rect 0 44563 624 44611
rect 186 44439 294 44515
rect 0 44343 624 44391
rect 186 44185 294 44295
rect 0 44089 624 44137
rect 186 43965 294 44041
rect 0 43869 624 43917
rect 0 43773 624 43821
rect 186 43649 294 43725
rect 0 43553 624 43601
rect 186 43395 294 43505
rect 0 43299 624 43347
rect 186 43175 294 43251
rect 0 43079 624 43127
rect 0 42983 624 43031
rect 186 42859 294 42935
rect 0 42763 624 42811
rect 186 42605 294 42715
rect 0 42509 624 42557
rect 186 42385 294 42461
rect 0 42289 624 42337
rect 0 42193 624 42241
rect 186 42069 294 42145
rect 0 41973 624 42021
rect 186 41815 294 41925
rect 0 41719 624 41767
rect 186 41595 294 41671
rect 0 41499 624 41547
rect 0 41403 624 41451
rect 186 41279 294 41355
rect 0 41183 624 41231
rect 186 41025 294 41135
rect 0 40929 624 40977
rect 186 40805 294 40881
rect 0 40709 624 40757
rect 0 40613 624 40661
rect 186 40489 294 40565
rect 0 40393 624 40441
rect 186 40235 294 40345
rect 0 40139 624 40187
rect 186 40015 294 40091
rect 0 39919 624 39967
rect 0 39823 624 39871
rect 186 39699 294 39775
rect 0 39603 624 39651
rect 186 39445 294 39555
rect 0 39349 624 39397
rect 186 39225 294 39301
rect 0 39129 624 39177
rect 0 39033 624 39081
rect 186 38909 294 38985
rect 0 38813 624 38861
rect 186 38655 294 38765
rect 0 38559 624 38607
rect 186 38435 294 38511
rect 0 38339 624 38387
rect 0 38243 624 38291
rect 186 38119 294 38195
rect 0 38023 624 38071
rect 186 37865 294 37975
rect 0 37769 624 37817
rect 186 37645 294 37721
rect 0 37549 624 37597
rect 0 37453 624 37501
rect 186 37329 294 37405
rect 0 37233 624 37281
rect 186 37075 294 37185
rect 0 36979 624 37027
rect 186 36855 294 36931
rect 0 36759 624 36807
rect 0 36663 624 36711
rect 186 36539 294 36615
rect 0 36443 624 36491
rect 186 36285 294 36395
rect 0 36189 624 36237
rect 186 36065 294 36141
rect 0 35969 624 36017
rect 0 35873 624 35921
rect 186 35749 294 35825
rect 0 35653 624 35701
rect 186 35495 294 35605
rect 0 35399 624 35447
rect 186 35275 294 35351
rect 0 35179 624 35227
rect 0 35083 624 35131
rect 186 34959 294 35035
rect 0 34863 624 34911
rect 186 34705 294 34815
rect 0 34609 624 34657
rect 186 34485 294 34561
rect 0 34389 624 34437
rect 0 34293 624 34341
rect 186 34169 294 34245
rect 0 34073 624 34121
rect 186 33915 294 34025
rect 0 33819 624 33867
rect 186 33695 294 33771
rect 0 33599 624 33647
rect 0 33503 624 33551
rect 186 33379 294 33455
rect 0 33283 624 33331
rect 186 33125 294 33235
rect 0 33029 624 33077
rect 186 32905 294 32981
rect 0 32809 624 32857
rect 0 32713 624 32761
rect 186 32589 294 32665
rect 0 32493 624 32541
rect 186 32335 294 32445
rect 0 32239 624 32287
rect 186 32115 294 32191
rect 0 32019 624 32067
rect 0 31923 624 31971
rect 186 31799 294 31875
rect 0 31703 624 31751
rect 186 31545 294 31655
rect 0 31449 624 31497
rect 186 31325 294 31401
rect 0 31229 624 31277
rect 0 31133 624 31181
rect 186 31009 294 31085
rect 0 30913 624 30961
rect 186 30755 294 30865
rect 0 30659 624 30707
rect 186 30535 294 30611
rect 0 30439 624 30487
rect 0 30343 624 30391
rect 186 30219 294 30295
rect 0 30123 624 30171
rect 186 29965 294 30075
rect 0 29869 624 29917
rect 186 29745 294 29821
rect 0 29649 624 29697
rect 0 29553 624 29601
rect 186 29429 294 29505
rect 0 29333 624 29381
rect 186 29175 294 29285
rect 0 29079 624 29127
rect 186 28955 294 29031
rect 0 28859 624 28907
rect 0 28763 624 28811
rect 186 28639 294 28715
rect 0 28543 624 28591
rect 186 28385 294 28495
rect 0 28289 624 28337
rect 186 28165 294 28241
rect 0 28069 624 28117
rect 0 27973 624 28021
rect 186 27849 294 27925
rect 0 27753 624 27801
rect 186 27595 294 27705
rect 0 27499 624 27547
rect 186 27375 294 27451
rect 0 27279 624 27327
rect 0 27183 624 27231
rect 186 27059 294 27135
rect 0 26963 624 27011
rect 186 26805 294 26915
rect 0 26709 624 26757
rect 186 26585 294 26661
rect 0 26489 624 26537
rect 0 26393 624 26441
rect 186 26269 294 26345
rect 0 26173 624 26221
rect 186 26015 294 26125
rect 0 25919 624 25967
rect 186 25795 294 25871
rect 0 25699 624 25747
rect 0 25603 624 25651
rect 186 25479 294 25555
rect 0 25383 624 25431
rect 186 25225 294 25335
rect 0 25129 624 25177
rect 186 25005 294 25081
rect 0 24909 624 24957
rect 0 24813 624 24861
rect 186 24689 294 24765
rect 0 24593 624 24641
rect 186 24435 294 24545
rect 0 24339 624 24387
rect 186 24215 294 24291
rect 0 24119 624 24167
rect 0 24023 624 24071
rect 186 23899 294 23975
rect 0 23803 624 23851
rect 186 23645 294 23755
rect 0 23549 624 23597
rect 186 23425 294 23501
rect 0 23329 624 23377
rect 0 23233 624 23281
rect 186 23109 294 23185
rect 0 23013 624 23061
rect 186 22855 294 22965
rect 0 22759 624 22807
rect 186 22635 294 22711
rect 0 22539 624 22587
rect 0 22443 624 22491
rect 186 22319 294 22395
rect 0 22223 624 22271
rect 186 22065 294 22175
rect 0 21969 624 22017
rect 186 21845 294 21921
rect 0 21749 624 21797
rect 0 21653 624 21701
rect 186 21529 294 21605
rect 0 21433 624 21481
rect 186 21275 294 21385
rect 0 21179 624 21227
rect 186 21055 294 21131
rect 0 20959 624 21007
rect 0 20863 624 20911
rect 186 20739 294 20815
rect 0 20643 624 20691
rect 186 20485 294 20595
rect 0 20389 624 20437
rect 186 20265 294 20341
rect 0 20169 624 20217
rect 0 20073 624 20121
rect 186 19949 294 20025
rect 0 19853 624 19901
rect 186 19695 294 19805
rect 0 19599 624 19647
rect 186 19475 294 19551
rect 0 19379 624 19427
rect 0 19283 624 19331
rect 186 19159 294 19235
rect 0 19063 624 19111
rect 186 18905 294 19015
rect 0 18809 624 18857
rect 186 18685 294 18761
rect 0 18589 624 18637
rect 0 18493 624 18541
rect 186 18369 294 18445
rect 0 18273 624 18321
rect 186 18115 294 18225
rect 0 18019 624 18067
rect 186 17895 294 17971
rect 0 17799 624 17847
rect 0 17703 624 17751
rect 186 17579 294 17655
rect 0 17483 624 17531
rect 186 17325 294 17435
rect 0 17229 624 17277
rect 186 17105 294 17181
rect 0 17009 624 17057
rect 0 16913 624 16961
rect 186 16789 294 16865
rect 0 16693 624 16741
rect 186 16535 294 16645
rect 0 16439 624 16487
rect 186 16315 294 16391
rect 0 16219 624 16267
rect 0 16123 624 16171
rect 186 15999 294 16075
rect 0 15903 624 15951
rect 186 15745 294 15855
rect 0 15649 624 15697
rect 186 15525 294 15601
rect 0 15429 624 15477
rect 0 15333 624 15381
rect 186 15209 294 15285
rect 0 15113 624 15161
rect 186 14955 294 15065
rect 0 14859 624 14907
rect 186 14735 294 14811
rect 0 14639 624 14687
rect 0 14543 624 14591
rect 186 14419 294 14495
rect 0 14323 624 14371
rect 186 14165 294 14275
rect 0 14069 624 14117
rect 186 13945 294 14021
rect 0 13849 624 13897
rect 0 13753 624 13801
rect 186 13629 294 13705
rect 0 13533 624 13581
rect 186 13375 294 13485
rect 0 13279 624 13327
rect 186 13155 294 13231
rect 0 13059 624 13107
rect 0 12963 624 13011
rect 186 12839 294 12915
rect 0 12743 624 12791
rect 186 12585 294 12695
rect 0 12489 624 12537
rect 186 12365 294 12441
rect 0 12269 624 12317
rect 0 12173 624 12221
rect 186 12049 294 12125
rect 0 11953 624 12001
rect 186 11795 294 11905
rect 0 11699 624 11747
rect 186 11575 294 11651
rect 0 11479 624 11527
rect 0 11383 624 11431
rect 186 11259 294 11335
rect 0 11163 624 11211
rect 186 11005 294 11115
rect 0 10909 624 10957
rect 186 10785 294 10861
rect 0 10689 624 10737
rect 0 10593 624 10641
rect 186 10469 294 10545
rect 0 10373 624 10421
rect 186 10215 294 10325
rect 0 10119 624 10167
rect 186 9995 294 10071
rect 0 9899 624 9947
rect 0 9803 624 9851
rect 186 9679 294 9755
rect 0 9583 624 9631
rect 186 9425 294 9535
rect 0 9329 624 9377
rect 186 9205 294 9281
rect 0 9109 624 9157
rect 0 9013 624 9061
rect 186 8889 294 8965
rect 0 8793 624 8841
rect 186 8635 294 8745
rect 0 8539 624 8587
rect 186 8415 294 8491
rect 0 8319 624 8367
rect 0 8223 624 8271
rect 186 8099 294 8175
rect 0 8003 624 8051
rect 186 7845 294 7955
rect 0 7749 624 7797
rect 186 7625 294 7701
rect 0 7529 624 7577
rect 0 7433 624 7481
rect 186 7309 294 7385
rect 0 7213 624 7261
rect 186 7055 294 7165
rect 0 6959 624 7007
rect 186 6835 294 6911
rect 0 6739 624 6787
rect 0 6643 624 6691
rect 186 6519 294 6595
rect 0 6423 624 6471
rect 186 6265 294 6375
rect 0 6169 624 6217
rect 186 6045 294 6121
rect 0 5949 624 5997
rect 0 5853 624 5901
rect 186 5729 294 5805
rect 0 5633 624 5681
rect 186 5475 294 5585
rect 0 5379 624 5427
rect 186 5255 294 5331
rect 0 5159 624 5207
rect 0 5063 624 5111
rect 186 4939 294 5015
rect 0 4843 624 4891
rect 186 4685 294 4795
rect 0 4589 624 4637
rect 186 4465 294 4541
rect 0 4369 624 4417
rect 0 4273 624 4321
rect 186 4149 294 4225
rect 0 4053 624 4101
rect 186 3895 294 4005
rect 0 3799 624 3847
rect 186 3675 294 3751
rect 0 3579 624 3627
rect 0 3483 624 3531
rect 186 3359 294 3435
rect 0 3263 624 3311
rect 186 3105 294 3215
rect 0 3009 624 3057
rect 186 2885 294 2961
rect 0 2789 624 2837
rect 0 2693 624 2741
rect 186 2569 294 2645
rect 0 2473 624 2521
rect 186 2315 294 2425
rect 0 2219 624 2267
rect 186 2095 294 2171
rect 0 1999 624 2047
rect 0 1903 624 1951
rect 186 1779 294 1855
rect 0 1683 624 1731
rect 186 1525 294 1635
rect 0 1429 624 1477
rect 186 1305 294 1381
rect 0 1209 624 1257
rect 0 1113 624 1161
rect 186 989 294 1065
rect 0 893 624 941
rect 186 735 294 845
rect 0 639 624 687
rect 186 515 294 591
rect 0 419 624 467
<< metal3 >>
rect 263 102422 361 102520
rect 263 180 361 278
use contact_9  contact_9_1
timestamp 1624494425
transform 1 0 279 0 1 192
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_1
timestamp 1624494425
transform 1 0 0 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_0
timestamp 1624494425
transform 1 0 0 0 -1 102700
box 0 0 624 474
use contact_9  contact_9_0
timestamp 1624494425
transform 1 0 279 0 1 102434
box 0 0 66 74
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_0
timestamp 1624494425
transform 1 0 0 0 -1 790
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_256
timestamp 1624494425
transform 1 0 0 0 1 790
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_255
timestamp 1624494425
transform 1 0 0 0 -1 1580
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_254
timestamp 1624494425
transform 1 0 0 0 1 1580
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_253
timestamp 1624494425
transform 1 0 0 0 -1 2370
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_252
timestamp 1624494425
transform 1 0 0 0 1 2370
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_251
timestamp 1624494425
transform 1 0 0 0 -1 3160
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_250
timestamp 1624494425
transform 1 0 0 0 1 3160
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_249
timestamp 1624494425
transform 1 0 0 0 -1 3950
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_248
timestamp 1624494425
transform 1 0 0 0 1 3950
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_247
timestamp 1624494425
transform 1 0 0 0 -1 4740
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_246
timestamp 1624494425
transform 1 0 0 0 1 4740
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_245
timestamp 1624494425
transform 1 0 0 0 -1 5530
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_244
timestamp 1624494425
transform 1 0 0 0 1 5530
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_243
timestamp 1624494425
transform 1 0 0 0 -1 6320
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_242
timestamp 1624494425
transform 1 0 0 0 1 6320
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_241
timestamp 1624494425
transform 1 0 0 0 -1 7110
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_240
timestamp 1624494425
transform 1 0 0 0 1 7110
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_239
timestamp 1624494425
transform 1 0 0 0 -1 7900
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_238
timestamp 1624494425
transform 1 0 0 0 1 7900
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_237
timestamp 1624494425
transform 1 0 0 0 -1 8690
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_236
timestamp 1624494425
transform 1 0 0 0 1 8690
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_235
timestamp 1624494425
transform 1 0 0 0 -1 9480
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_234
timestamp 1624494425
transform 1 0 0 0 1 9480
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_233
timestamp 1624494425
transform 1 0 0 0 -1 10270
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_232
timestamp 1624494425
transform 1 0 0 0 1 10270
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_231
timestamp 1624494425
transform 1 0 0 0 -1 11060
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_230
timestamp 1624494425
transform 1 0 0 0 1 11060
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_229
timestamp 1624494425
transform 1 0 0 0 -1 11850
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_228
timestamp 1624494425
transform 1 0 0 0 1 11850
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_227
timestamp 1624494425
transform 1 0 0 0 -1 12640
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_226
timestamp 1624494425
transform 1 0 0 0 1 12640
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_225
timestamp 1624494425
transform 1 0 0 0 -1 13430
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_224
timestamp 1624494425
transform 1 0 0 0 1 13430
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_223
timestamp 1624494425
transform 1 0 0 0 -1 14220
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_222
timestamp 1624494425
transform 1 0 0 0 1 14220
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_221
timestamp 1624494425
transform 1 0 0 0 -1 15010
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_220
timestamp 1624494425
transform 1 0 0 0 1 15010
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_219
timestamp 1624494425
transform 1 0 0 0 -1 15800
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_218
timestamp 1624494425
transform 1 0 0 0 1 15800
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_217
timestamp 1624494425
transform 1 0 0 0 -1 16590
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_216
timestamp 1624494425
transform 1 0 0 0 1 16590
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_215
timestamp 1624494425
transform 1 0 0 0 -1 17380
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_214
timestamp 1624494425
transform 1 0 0 0 1 17380
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_213
timestamp 1624494425
transform 1 0 0 0 -1 18170
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_212
timestamp 1624494425
transform 1 0 0 0 1 18170
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_211
timestamp 1624494425
transform 1 0 0 0 -1 18960
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_210
timestamp 1624494425
transform 1 0 0 0 1 18960
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_209
timestamp 1624494425
transform 1 0 0 0 -1 19750
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_208
timestamp 1624494425
transform 1 0 0 0 1 19750
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_207
timestamp 1624494425
transform 1 0 0 0 -1 20540
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_206
timestamp 1624494425
transform 1 0 0 0 1 20540
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_205
timestamp 1624494425
transform 1 0 0 0 -1 21330
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_204
timestamp 1624494425
transform 1 0 0 0 1 21330
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_203
timestamp 1624494425
transform 1 0 0 0 -1 22120
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_202
timestamp 1624494425
transform 1 0 0 0 1 22120
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_201
timestamp 1624494425
transform 1 0 0 0 -1 22910
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_200
timestamp 1624494425
transform 1 0 0 0 1 22910
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_199
timestamp 1624494425
transform 1 0 0 0 -1 23700
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_198
timestamp 1624494425
transform 1 0 0 0 1 23700
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_197
timestamp 1624494425
transform 1 0 0 0 -1 24490
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_196
timestamp 1624494425
transform 1 0 0 0 1 24490
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_195
timestamp 1624494425
transform 1 0 0 0 -1 25280
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_194
timestamp 1624494425
transform 1 0 0 0 1 25280
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_193
timestamp 1624494425
transform 1 0 0 0 -1 26070
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_192
timestamp 1624494425
transform 1 0 0 0 1 26070
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_191
timestamp 1624494425
transform 1 0 0 0 -1 26860
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_190
timestamp 1624494425
transform 1 0 0 0 1 26860
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_189
timestamp 1624494425
transform 1 0 0 0 -1 27650
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_188
timestamp 1624494425
transform 1 0 0 0 1 27650
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_187
timestamp 1624494425
transform 1 0 0 0 -1 28440
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_186
timestamp 1624494425
transform 1 0 0 0 1 28440
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_185
timestamp 1624494425
transform 1 0 0 0 -1 29230
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_184
timestamp 1624494425
transform 1 0 0 0 1 29230
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_183
timestamp 1624494425
transform 1 0 0 0 -1 30020
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_182
timestamp 1624494425
transform 1 0 0 0 1 30020
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_181
timestamp 1624494425
transform 1 0 0 0 -1 30810
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_180
timestamp 1624494425
transform 1 0 0 0 1 30810
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_179
timestamp 1624494425
transform 1 0 0 0 -1 31600
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_178
timestamp 1624494425
transform 1 0 0 0 1 31600
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_177
timestamp 1624494425
transform 1 0 0 0 -1 32390
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_176
timestamp 1624494425
transform 1 0 0 0 1 32390
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_175
timestamp 1624494425
transform 1 0 0 0 -1 33180
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_174
timestamp 1624494425
transform 1 0 0 0 1 33180
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_173
timestamp 1624494425
transform 1 0 0 0 -1 33970
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_172
timestamp 1624494425
transform 1 0 0 0 1 33970
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_171
timestamp 1624494425
transform 1 0 0 0 -1 34760
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_170
timestamp 1624494425
transform 1 0 0 0 1 34760
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_169
timestamp 1624494425
transform 1 0 0 0 -1 35550
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_168
timestamp 1624494425
transform 1 0 0 0 1 35550
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_167
timestamp 1624494425
transform 1 0 0 0 -1 36340
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_166
timestamp 1624494425
transform 1 0 0 0 1 36340
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_165
timestamp 1624494425
transform 1 0 0 0 -1 37130
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_164
timestamp 1624494425
transform 1 0 0 0 1 37130
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_163
timestamp 1624494425
transform 1 0 0 0 -1 37920
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_162
timestamp 1624494425
transform 1 0 0 0 1 37920
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_161
timestamp 1624494425
transform 1 0 0 0 -1 38710
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_160
timestamp 1624494425
transform 1 0 0 0 1 38710
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_159
timestamp 1624494425
transform 1 0 0 0 -1 39500
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_158
timestamp 1624494425
transform 1 0 0 0 1 39500
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_157
timestamp 1624494425
transform 1 0 0 0 -1 40290
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_156
timestamp 1624494425
transform 1 0 0 0 1 40290
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_155
timestamp 1624494425
transform 1 0 0 0 -1 41080
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_154
timestamp 1624494425
transform 1 0 0 0 1 41080
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_153
timestamp 1624494425
transform 1 0 0 0 -1 41870
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_152
timestamp 1624494425
transform 1 0 0 0 1 41870
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_151
timestamp 1624494425
transform 1 0 0 0 -1 42660
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_150
timestamp 1624494425
transform 1 0 0 0 1 42660
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_149
timestamp 1624494425
transform 1 0 0 0 -1 43450
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_148
timestamp 1624494425
transform 1 0 0 0 1 43450
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_147
timestamp 1624494425
transform 1 0 0 0 -1 44240
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_146
timestamp 1624494425
transform 1 0 0 0 1 44240
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_145
timestamp 1624494425
transform 1 0 0 0 -1 45030
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_144
timestamp 1624494425
transform 1 0 0 0 1 45030
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_143
timestamp 1624494425
transform 1 0 0 0 -1 45820
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_142
timestamp 1624494425
transform 1 0 0 0 1 45820
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_141
timestamp 1624494425
transform 1 0 0 0 -1 46610
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_140
timestamp 1624494425
transform 1 0 0 0 1 46610
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_139
timestamp 1624494425
transform 1 0 0 0 -1 47400
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_138
timestamp 1624494425
transform 1 0 0 0 1 47400
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_137
timestamp 1624494425
transform 1 0 0 0 -1 48190
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_136
timestamp 1624494425
transform 1 0 0 0 1 48190
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_135
timestamp 1624494425
transform 1 0 0 0 -1 48980
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_134
timestamp 1624494425
transform 1 0 0 0 1 48980
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_133
timestamp 1624494425
transform 1 0 0 0 -1 49770
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_132
timestamp 1624494425
transform 1 0 0 0 1 49770
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_131
timestamp 1624494425
transform 1 0 0 0 -1 50560
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_130
timestamp 1624494425
transform 1 0 0 0 1 50560
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_129
timestamp 1624494425
transform 1 0 0 0 -1 51350
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_128
timestamp 1624494425
transform 1 0 0 0 1 51350
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_127
timestamp 1624494425
transform 1 0 0 0 -1 52140
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_126
timestamp 1624494425
transform 1 0 0 0 1 52140
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_125
timestamp 1624494425
transform 1 0 0 0 -1 52930
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_124
timestamp 1624494425
transform 1 0 0 0 1 52930
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_123
timestamp 1624494425
transform 1 0 0 0 -1 53720
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_122
timestamp 1624494425
transform 1 0 0 0 1 53720
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_121
timestamp 1624494425
transform 1 0 0 0 -1 54510
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_120
timestamp 1624494425
transform 1 0 0 0 1 54510
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_119
timestamp 1624494425
transform 1 0 0 0 -1 55300
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_118
timestamp 1624494425
transform 1 0 0 0 1 55300
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_117
timestamp 1624494425
transform 1 0 0 0 -1 56090
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_116
timestamp 1624494425
transform 1 0 0 0 1 56090
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_115
timestamp 1624494425
transform 1 0 0 0 -1 56880
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_114
timestamp 1624494425
transform 1 0 0 0 1 56880
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_113
timestamp 1624494425
transform 1 0 0 0 -1 57670
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_112
timestamp 1624494425
transform 1 0 0 0 1 57670
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_111
timestamp 1624494425
transform 1 0 0 0 -1 58460
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_110
timestamp 1624494425
transform 1 0 0 0 1 58460
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_109
timestamp 1624494425
transform 1 0 0 0 -1 59250
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_108
timestamp 1624494425
transform 1 0 0 0 1 59250
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_107
timestamp 1624494425
transform 1 0 0 0 -1 60040
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_106
timestamp 1624494425
transform 1 0 0 0 1 60040
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_105
timestamp 1624494425
transform 1 0 0 0 -1 60830
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_104
timestamp 1624494425
transform 1 0 0 0 1 60830
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_103
timestamp 1624494425
transform 1 0 0 0 -1 61620
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_102
timestamp 1624494425
transform 1 0 0 0 1 61620
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_101
timestamp 1624494425
transform 1 0 0 0 -1 62410
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_100
timestamp 1624494425
transform 1 0 0 0 1 62410
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_99
timestamp 1624494425
transform 1 0 0 0 -1 63200
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_98
timestamp 1624494425
transform 1 0 0 0 1 63200
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_97
timestamp 1624494425
transform 1 0 0 0 -1 63990
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_96
timestamp 1624494425
transform 1 0 0 0 1 63990
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_95
timestamp 1624494425
transform 1 0 0 0 -1 64780
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_94
timestamp 1624494425
transform 1 0 0 0 1 64780
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_93
timestamp 1624494425
transform 1 0 0 0 -1 65570
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_92
timestamp 1624494425
transform 1 0 0 0 1 65570
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_91
timestamp 1624494425
transform 1 0 0 0 -1 66360
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_90
timestamp 1624494425
transform 1 0 0 0 1 66360
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_89
timestamp 1624494425
transform 1 0 0 0 -1 67150
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_88
timestamp 1624494425
transform 1 0 0 0 1 67150
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_87
timestamp 1624494425
transform 1 0 0 0 -1 67940
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_86
timestamp 1624494425
transform 1 0 0 0 1 67940
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_85
timestamp 1624494425
transform 1 0 0 0 -1 68730
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_84
timestamp 1624494425
transform 1 0 0 0 1 68730
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_83
timestamp 1624494425
transform 1 0 0 0 -1 69520
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_82
timestamp 1624494425
transform 1 0 0 0 1 69520
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_81
timestamp 1624494425
transform 1 0 0 0 -1 70310
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_80
timestamp 1624494425
transform 1 0 0 0 1 70310
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_79
timestamp 1624494425
transform 1 0 0 0 -1 71100
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_78
timestamp 1624494425
transform 1 0 0 0 1 71100
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_77
timestamp 1624494425
transform 1 0 0 0 -1 71890
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_76
timestamp 1624494425
transform 1 0 0 0 1 71890
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_75
timestamp 1624494425
transform 1 0 0 0 -1 72680
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_74
timestamp 1624494425
transform 1 0 0 0 1 72680
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_73
timestamp 1624494425
transform 1 0 0 0 -1 73470
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_72
timestamp 1624494425
transform 1 0 0 0 1 73470
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_71
timestamp 1624494425
transform 1 0 0 0 -1 74260
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_70
timestamp 1624494425
transform 1 0 0 0 1 74260
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_69
timestamp 1624494425
transform 1 0 0 0 -1 75050
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_68
timestamp 1624494425
transform 1 0 0 0 1 75050
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_67
timestamp 1624494425
transform 1 0 0 0 -1 75840
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_66
timestamp 1624494425
transform 1 0 0 0 1 75840
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_65
timestamp 1624494425
transform 1 0 0 0 -1 76630
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_64
timestamp 1624494425
transform 1 0 0 0 1 76630
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_63
timestamp 1624494425
transform 1 0 0 0 -1 77420
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_62
timestamp 1624494425
transform 1 0 0 0 1 77420
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_61
timestamp 1624494425
transform 1 0 0 0 -1 78210
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_60
timestamp 1624494425
transform 1 0 0 0 1 78210
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_59
timestamp 1624494425
transform 1 0 0 0 -1 79000
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_58
timestamp 1624494425
transform 1 0 0 0 1 79000
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_57
timestamp 1624494425
transform 1 0 0 0 -1 79790
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_56
timestamp 1624494425
transform 1 0 0 0 1 79790
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_55
timestamp 1624494425
transform 1 0 0 0 -1 80580
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_54
timestamp 1624494425
transform 1 0 0 0 1 80580
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_53
timestamp 1624494425
transform 1 0 0 0 -1 81370
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_52
timestamp 1624494425
transform 1 0 0 0 1 81370
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_51
timestamp 1624494425
transform 1 0 0 0 -1 82160
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_50
timestamp 1624494425
transform 1 0 0 0 1 82160
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_49
timestamp 1624494425
transform 1 0 0 0 -1 82950
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_48
timestamp 1624494425
transform 1 0 0 0 1 82950
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_47
timestamp 1624494425
transform 1 0 0 0 -1 83740
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_46
timestamp 1624494425
transform 1 0 0 0 1 83740
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_45
timestamp 1624494425
transform 1 0 0 0 -1 84530
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_44
timestamp 1624494425
transform 1 0 0 0 1 84530
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_43
timestamp 1624494425
transform 1 0 0 0 -1 85320
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_42
timestamp 1624494425
transform 1 0 0 0 1 85320
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_41
timestamp 1624494425
transform 1 0 0 0 -1 86110
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_40
timestamp 1624494425
transform 1 0 0 0 1 86110
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_39
timestamp 1624494425
transform 1 0 0 0 -1 86900
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_38
timestamp 1624494425
transform 1 0 0 0 1 86900
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_37
timestamp 1624494425
transform 1 0 0 0 -1 87690
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_36
timestamp 1624494425
transform 1 0 0 0 1 87690
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_35
timestamp 1624494425
transform 1 0 0 0 -1 88480
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_34
timestamp 1624494425
transform 1 0 0 0 1 88480
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_33
timestamp 1624494425
transform 1 0 0 0 -1 89270
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_32
timestamp 1624494425
transform 1 0 0 0 1 89270
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_31
timestamp 1624494425
transform 1 0 0 0 -1 90060
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_30
timestamp 1624494425
transform 1 0 0 0 1 90060
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_29
timestamp 1624494425
transform 1 0 0 0 -1 90850
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_28
timestamp 1624494425
transform 1 0 0 0 1 90850
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_27
timestamp 1624494425
transform 1 0 0 0 -1 91640
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_26
timestamp 1624494425
transform 1 0 0 0 1 91640
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_25
timestamp 1624494425
transform 1 0 0 0 -1 92430
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_24
timestamp 1624494425
transform 1 0 0 0 1 92430
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_23
timestamp 1624494425
transform 1 0 0 0 -1 93220
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_22
timestamp 1624494425
transform 1 0 0 0 1 93220
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_21
timestamp 1624494425
transform 1 0 0 0 -1 94010
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_20
timestamp 1624494425
transform 1 0 0 0 1 94010
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_19
timestamp 1624494425
transform 1 0 0 0 -1 94800
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_18
timestamp 1624494425
transform 1 0 0 0 1 94800
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_17
timestamp 1624494425
transform 1 0 0 0 -1 95590
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_16
timestamp 1624494425
transform 1 0 0 0 1 95590
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_15
timestamp 1624494425
transform 1 0 0 0 -1 96380
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_14
timestamp 1624494425
transform 1 0 0 0 1 96380
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_13
timestamp 1624494425
transform 1 0 0 0 -1 97170
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_12
timestamp 1624494425
transform 1 0 0 0 1 97170
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_11
timestamp 1624494425
transform 1 0 0 0 -1 97960
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_10
timestamp 1624494425
transform 1 0 0 0 1 97960
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_9
timestamp 1624494425
transform 1 0 0 0 -1 98750
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_8
timestamp 1624494425
transform 1 0 0 0 1 98750
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_7
timestamp 1624494425
transform 1 0 0 0 -1 99540
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_6
timestamp 1624494425
transform 1 0 0 0 1 99540
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_5
timestamp 1624494425
transform 1 0 0 0 -1 100330
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_4
timestamp 1624494425
transform 1 0 0 0 1 100330
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_3
timestamp 1624494425
transform 1 0 0 0 -1 101120
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_2
timestamp 1624494425
transform 1 0 0 0 1 101120
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_1
timestamp 1624494425
transform 1 0 0 0 -1 101910
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_0
timestamp 1624494425
transform 1 0 0 0 1 101910
box -42 -105 650 424
<< labels >>
rlabel metal1 s 78 0 114 102700 4 bl_0_0
rlabel metal1 s 150 0 186 102700 4 br_0_0
rlabel metal1 s 294 0 330 102700 4 bl_1_0
rlabel metal1 s 366 0 402 102700 4 br_1_0
rlabel metal2 s 0 419 624 467 4 wl_0_0
rlabel metal2 s 0 1113 624 1161 4 wl_0_1
rlabel metal2 s 0 1209 624 1257 4 wl_0_2
rlabel metal2 s 0 1903 624 1951 4 wl_0_3
rlabel metal2 s 0 1999 624 2047 4 wl_0_4
rlabel metal2 s 0 2693 624 2741 4 wl_0_5
rlabel metal2 s 0 2789 624 2837 4 wl_0_6
rlabel metal2 s 0 3483 624 3531 4 wl_0_7
rlabel metal2 s 0 3579 624 3627 4 wl_0_8
rlabel metal2 s 0 4273 624 4321 4 wl_0_9
rlabel metal2 s 0 4369 624 4417 4 wl_0_10
rlabel metal2 s 0 5063 624 5111 4 wl_0_11
rlabel metal2 s 0 5159 624 5207 4 wl_0_12
rlabel metal2 s 0 5853 624 5901 4 wl_0_13
rlabel metal2 s 0 5949 624 5997 4 wl_0_14
rlabel metal2 s 0 6643 624 6691 4 wl_0_15
rlabel metal2 s 0 6739 624 6787 4 wl_0_16
rlabel metal2 s 0 7433 624 7481 4 wl_0_17
rlabel metal2 s 0 7529 624 7577 4 wl_0_18
rlabel metal2 s 0 8223 624 8271 4 wl_0_19
rlabel metal2 s 0 8319 624 8367 4 wl_0_20
rlabel metal2 s 0 9013 624 9061 4 wl_0_21
rlabel metal2 s 0 9109 624 9157 4 wl_0_22
rlabel metal2 s 0 9803 624 9851 4 wl_0_23
rlabel metal2 s 0 9899 624 9947 4 wl_0_24
rlabel metal2 s 0 10593 624 10641 4 wl_0_25
rlabel metal2 s 0 10689 624 10737 4 wl_0_26
rlabel metal2 s 0 11383 624 11431 4 wl_0_27
rlabel metal2 s 0 11479 624 11527 4 wl_0_28
rlabel metal2 s 0 12173 624 12221 4 wl_0_29
rlabel metal2 s 0 12269 624 12317 4 wl_0_30
rlabel metal2 s 0 12963 624 13011 4 wl_0_31
rlabel metal2 s 0 13059 624 13107 4 wl_0_32
rlabel metal2 s 0 13753 624 13801 4 wl_0_33
rlabel metal2 s 0 13849 624 13897 4 wl_0_34
rlabel metal2 s 0 14543 624 14591 4 wl_0_35
rlabel metal2 s 0 14639 624 14687 4 wl_0_36
rlabel metal2 s 0 15333 624 15381 4 wl_0_37
rlabel metal2 s 0 15429 624 15477 4 wl_0_38
rlabel metal2 s 0 16123 624 16171 4 wl_0_39
rlabel metal2 s 0 16219 624 16267 4 wl_0_40
rlabel metal2 s 0 16913 624 16961 4 wl_0_41
rlabel metal2 s 0 17009 624 17057 4 wl_0_42
rlabel metal2 s 0 17703 624 17751 4 wl_0_43
rlabel metal2 s 0 17799 624 17847 4 wl_0_44
rlabel metal2 s 0 18493 624 18541 4 wl_0_45
rlabel metal2 s 0 18589 624 18637 4 wl_0_46
rlabel metal2 s 0 19283 624 19331 4 wl_0_47
rlabel metal2 s 0 19379 624 19427 4 wl_0_48
rlabel metal2 s 0 20073 624 20121 4 wl_0_49
rlabel metal2 s 0 20169 624 20217 4 wl_0_50
rlabel metal2 s 0 20863 624 20911 4 wl_0_51
rlabel metal2 s 0 20959 624 21007 4 wl_0_52
rlabel metal2 s 0 21653 624 21701 4 wl_0_53
rlabel metal2 s 0 21749 624 21797 4 wl_0_54
rlabel metal2 s 0 22443 624 22491 4 wl_0_55
rlabel metal2 s 0 22539 624 22587 4 wl_0_56
rlabel metal2 s 0 23233 624 23281 4 wl_0_57
rlabel metal2 s 0 23329 624 23377 4 wl_0_58
rlabel metal2 s 0 24023 624 24071 4 wl_0_59
rlabel metal2 s 0 24119 624 24167 4 wl_0_60
rlabel metal2 s 0 24813 624 24861 4 wl_0_61
rlabel metal2 s 0 24909 624 24957 4 wl_0_62
rlabel metal2 s 0 25603 624 25651 4 wl_0_63
rlabel metal2 s 0 25699 624 25747 4 wl_0_64
rlabel metal2 s 0 26393 624 26441 4 wl_0_65
rlabel metal2 s 0 26489 624 26537 4 wl_0_66
rlabel metal2 s 0 27183 624 27231 4 wl_0_67
rlabel metal2 s 0 27279 624 27327 4 wl_0_68
rlabel metal2 s 0 27973 624 28021 4 wl_0_69
rlabel metal2 s 0 28069 624 28117 4 wl_0_70
rlabel metal2 s 0 28763 624 28811 4 wl_0_71
rlabel metal2 s 0 28859 624 28907 4 wl_0_72
rlabel metal2 s 0 29553 624 29601 4 wl_0_73
rlabel metal2 s 0 29649 624 29697 4 wl_0_74
rlabel metal2 s 0 30343 624 30391 4 wl_0_75
rlabel metal2 s 0 30439 624 30487 4 wl_0_76
rlabel metal2 s 0 31133 624 31181 4 wl_0_77
rlabel metal2 s 0 31229 624 31277 4 wl_0_78
rlabel metal2 s 0 31923 624 31971 4 wl_0_79
rlabel metal2 s 0 32019 624 32067 4 wl_0_80
rlabel metal2 s 0 32713 624 32761 4 wl_0_81
rlabel metal2 s 0 32809 624 32857 4 wl_0_82
rlabel metal2 s 0 33503 624 33551 4 wl_0_83
rlabel metal2 s 0 33599 624 33647 4 wl_0_84
rlabel metal2 s 0 34293 624 34341 4 wl_0_85
rlabel metal2 s 0 34389 624 34437 4 wl_0_86
rlabel metal2 s 0 35083 624 35131 4 wl_0_87
rlabel metal2 s 0 35179 624 35227 4 wl_0_88
rlabel metal2 s 0 35873 624 35921 4 wl_0_89
rlabel metal2 s 0 35969 624 36017 4 wl_0_90
rlabel metal2 s 0 36663 624 36711 4 wl_0_91
rlabel metal2 s 0 36759 624 36807 4 wl_0_92
rlabel metal2 s 0 37453 624 37501 4 wl_0_93
rlabel metal2 s 0 37549 624 37597 4 wl_0_94
rlabel metal2 s 0 38243 624 38291 4 wl_0_95
rlabel metal2 s 0 38339 624 38387 4 wl_0_96
rlabel metal2 s 0 39033 624 39081 4 wl_0_97
rlabel metal2 s 0 39129 624 39177 4 wl_0_98
rlabel metal2 s 0 39823 624 39871 4 wl_0_99
rlabel metal2 s 0 39919 624 39967 4 wl_0_100
rlabel metal2 s 0 40613 624 40661 4 wl_0_101
rlabel metal2 s 0 40709 624 40757 4 wl_0_102
rlabel metal2 s 0 41403 624 41451 4 wl_0_103
rlabel metal2 s 0 41499 624 41547 4 wl_0_104
rlabel metal2 s 0 42193 624 42241 4 wl_0_105
rlabel metal2 s 0 42289 624 42337 4 wl_0_106
rlabel metal2 s 0 42983 624 43031 4 wl_0_107
rlabel metal2 s 0 43079 624 43127 4 wl_0_108
rlabel metal2 s 0 43773 624 43821 4 wl_0_109
rlabel metal2 s 0 43869 624 43917 4 wl_0_110
rlabel metal2 s 0 44563 624 44611 4 wl_0_111
rlabel metal2 s 0 44659 624 44707 4 wl_0_112
rlabel metal2 s 0 45353 624 45401 4 wl_0_113
rlabel metal2 s 0 45449 624 45497 4 wl_0_114
rlabel metal2 s 0 46143 624 46191 4 wl_0_115
rlabel metal2 s 0 46239 624 46287 4 wl_0_116
rlabel metal2 s 0 46933 624 46981 4 wl_0_117
rlabel metal2 s 0 47029 624 47077 4 wl_0_118
rlabel metal2 s 0 47723 624 47771 4 wl_0_119
rlabel metal2 s 0 47819 624 47867 4 wl_0_120
rlabel metal2 s 0 48513 624 48561 4 wl_0_121
rlabel metal2 s 0 48609 624 48657 4 wl_0_122
rlabel metal2 s 0 49303 624 49351 4 wl_0_123
rlabel metal2 s 0 49399 624 49447 4 wl_0_124
rlabel metal2 s 0 50093 624 50141 4 wl_0_125
rlabel metal2 s 0 50189 624 50237 4 wl_0_126
rlabel metal2 s 0 50883 624 50931 4 wl_0_127
rlabel metal2 s 0 50979 624 51027 4 wl_0_128
rlabel metal2 s 0 51673 624 51721 4 wl_0_129
rlabel metal2 s 0 51769 624 51817 4 wl_0_130
rlabel metal2 s 0 52463 624 52511 4 wl_0_131
rlabel metal2 s 0 52559 624 52607 4 wl_0_132
rlabel metal2 s 0 53253 624 53301 4 wl_0_133
rlabel metal2 s 0 53349 624 53397 4 wl_0_134
rlabel metal2 s 0 54043 624 54091 4 wl_0_135
rlabel metal2 s 0 54139 624 54187 4 wl_0_136
rlabel metal2 s 0 54833 624 54881 4 wl_0_137
rlabel metal2 s 0 54929 624 54977 4 wl_0_138
rlabel metal2 s 0 55623 624 55671 4 wl_0_139
rlabel metal2 s 0 55719 624 55767 4 wl_0_140
rlabel metal2 s 0 56413 624 56461 4 wl_0_141
rlabel metal2 s 0 56509 624 56557 4 wl_0_142
rlabel metal2 s 0 57203 624 57251 4 wl_0_143
rlabel metal2 s 0 57299 624 57347 4 wl_0_144
rlabel metal2 s 0 57993 624 58041 4 wl_0_145
rlabel metal2 s 0 58089 624 58137 4 wl_0_146
rlabel metal2 s 0 58783 624 58831 4 wl_0_147
rlabel metal2 s 0 58879 624 58927 4 wl_0_148
rlabel metal2 s 0 59573 624 59621 4 wl_0_149
rlabel metal2 s 0 59669 624 59717 4 wl_0_150
rlabel metal2 s 0 60363 624 60411 4 wl_0_151
rlabel metal2 s 0 60459 624 60507 4 wl_0_152
rlabel metal2 s 0 61153 624 61201 4 wl_0_153
rlabel metal2 s 0 61249 624 61297 4 wl_0_154
rlabel metal2 s 0 61943 624 61991 4 wl_0_155
rlabel metal2 s 0 62039 624 62087 4 wl_0_156
rlabel metal2 s 0 62733 624 62781 4 wl_0_157
rlabel metal2 s 0 62829 624 62877 4 wl_0_158
rlabel metal2 s 0 63523 624 63571 4 wl_0_159
rlabel metal2 s 0 63619 624 63667 4 wl_0_160
rlabel metal2 s 0 64313 624 64361 4 wl_0_161
rlabel metal2 s 0 64409 624 64457 4 wl_0_162
rlabel metal2 s 0 65103 624 65151 4 wl_0_163
rlabel metal2 s 0 65199 624 65247 4 wl_0_164
rlabel metal2 s 0 65893 624 65941 4 wl_0_165
rlabel metal2 s 0 65989 624 66037 4 wl_0_166
rlabel metal2 s 0 66683 624 66731 4 wl_0_167
rlabel metal2 s 0 66779 624 66827 4 wl_0_168
rlabel metal2 s 0 67473 624 67521 4 wl_0_169
rlabel metal2 s 0 67569 624 67617 4 wl_0_170
rlabel metal2 s 0 68263 624 68311 4 wl_0_171
rlabel metal2 s 0 68359 624 68407 4 wl_0_172
rlabel metal2 s 0 69053 624 69101 4 wl_0_173
rlabel metal2 s 0 69149 624 69197 4 wl_0_174
rlabel metal2 s 0 69843 624 69891 4 wl_0_175
rlabel metal2 s 0 69939 624 69987 4 wl_0_176
rlabel metal2 s 0 70633 624 70681 4 wl_0_177
rlabel metal2 s 0 70729 624 70777 4 wl_0_178
rlabel metal2 s 0 71423 624 71471 4 wl_0_179
rlabel metal2 s 0 71519 624 71567 4 wl_0_180
rlabel metal2 s 0 72213 624 72261 4 wl_0_181
rlabel metal2 s 0 72309 624 72357 4 wl_0_182
rlabel metal2 s 0 73003 624 73051 4 wl_0_183
rlabel metal2 s 0 73099 624 73147 4 wl_0_184
rlabel metal2 s 0 73793 624 73841 4 wl_0_185
rlabel metal2 s 0 73889 624 73937 4 wl_0_186
rlabel metal2 s 0 74583 624 74631 4 wl_0_187
rlabel metal2 s 0 74679 624 74727 4 wl_0_188
rlabel metal2 s 0 75373 624 75421 4 wl_0_189
rlabel metal2 s 0 75469 624 75517 4 wl_0_190
rlabel metal2 s 0 76163 624 76211 4 wl_0_191
rlabel metal2 s 0 76259 624 76307 4 wl_0_192
rlabel metal2 s 0 76953 624 77001 4 wl_0_193
rlabel metal2 s 0 77049 624 77097 4 wl_0_194
rlabel metal2 s 0 77743 624 77791 4 wl_0_195
rlabel metal2 s 0 77839 624 77887 4 wl_0_196
rlabel metal2 s 0 78533 624 78581 4 wl_0_197
rlabel metal2 s 0 78629 624 78677 4 wl_0_198
rlabel metal2 s 0 79323 624 79371 4 wl_0_199
rlabel metal2 s 0 79419 624 79467 4 wl_0_200
rlabel metal2 s 0 80113 624 80161 4 wl_0_201
rlabel metal2 s 0 80209 624 80257 4 wl_0_202
rlabel metal2 s 0 80903 624 80951 4 wl_0_203
rlabel metal2 s 0 80999 624 81047 4 wl_0_204
rlabel metal2 s 0 81693 624 81741 4 wl_0_205
rlabel metal2 s 0 81789 624 81837 4 wl_0_206
rlabel metal2 s 0 82483 624 82531 4 wl_0_207
rlabel metal2 s 0 82579 624 82627 4 wl_0_208
rlabel metal2 s 0 83273 624 83321 4 wl_0_209
rlabel metal2 s 0 83369 624 83417 4 wl_0_210
rlabel metal2 s 0 84063 624 84111 4 wl_0_211
rlabel metal2 s 0 84159 624 84207 4 wl_0_212
rlabel metal2 s 0 84853 624 84901 4 wl_0_213
rlabel metal2 s 0 84949 624 84997 4 wl_0_214
rlabel metal2 s 0 85643 624 85691 4 wl_0_215
rlabel metal2 s 0 85739 624 85787 4 wl_0_216
rlabel metal2 s 0 86433 624 86481 4 wl_0_217
rlabel metal2 s 0 86529 624 86577 4 wl_0_218
rlabel metal2 s 0 87223 624 87271 4 wl_0_219
rlabel metal2 s 0 87319 624 87367 4 wl_0_220
rlabel metal2 s 0 88013 624 88061 4 wl_0_221
rlabel metal2 s 0 88109 624 88157 4 wl_0_222
rlabel metal2 s 0 88803 624 88851 4 wl_0_223
rlabel metal2 s 0 88899 624 88947 4 wl_0_224
rlabel metal2 s 0 89593 624 89641 4 wl_0_225
rlabel metal2 s 0 89689 624 89737 4 wl_0_226
rlabel metal2 s 0 90383 624 90431 4 wl_0_227
rlabel metal2 s 0 90479 624 90527 4 wl_0_228
rlabel metal2 s 0 91173 624 91221 4 wl_0_229
rlabel metal2 s 0 91269 624 91317 4 wl_0_230
rlabel metal2 s 0 91963 624 92011 4 wl_0_231
rlabel metal2 s 0 92059 624 92107 4 wl_0_232
rlabel metal2 s 0 92753 624 92801 4 wl_0_233
rlabel metal2 s 0 92849 624 92897 4 wl_0_234
rlabel metal2 s 0 93543 624 93591 4 wl_0_235
rlabel metal2 s 0 93639 624 93687 4 wl_0_236
rlabel metal2 s 0 94333 624 94381 4 wl_0_237
rlabel metal2 s 0 94429 624 94477 4 wl_0_238
rlabel metal2 s 0 95123 624 95171 4 wl_0_239
rlabel metal2 s 0 95219 624 95267 4 wl_0_240
rlabel metal2 s 0 95913 624 95961 4 wl_0_241
rlabel metal2 s 0 96009 624 96057 4 wl_0_242
rlabel metal2 s 0 96703 624 96751 4 wl_0_243
rlabel metal2 s 0 96799 624 96847 4 wl_0_244
rlabel metal2 s 0 97493 624 97541 4 wl_0_245
rlabel metal2 s 0 97589 624 97637 4 wl_0_246
rlabel metal2 s 0 98283 624 98331 4 wl_0_247
rlabel metal2 s 0 98379 624 98427 4 wl_0_248
rlabel metal2 s 0 99073 624 99121 4 wl_0_249
rlabel metal2 s 0 99169 624 99217 4 wl_0_250
rlabel metal2 s 0 99863 624 99911 4 wl_0_251
rlabel metal2 s 0 99959 624 100007 4 wl_0_252
rlabel metal2 s 0 100653 624 100701 4 wl_0_253
rlabel metal2 s 0 100749 624 100797 4 wl_0_254
rlabel metal2 s 0 101443 624 101491 4 wl_0_255
rlabel metal2 s 0 101539 624 101587 4 wl_0_256
rlabel metal2 s 0 102233 624 102281 4 wl_0_257
rlabel metal2 s 0 639 624 687 4 wl_1_0
rlabel metal2 s 0 893 624 941 4 wl_1_1
rlabel metal2 s 0 1429 624 1477 4 wl_1_2
rlabel metal2 s 0 1683 624 1731 4 wl_1_3
rlabel metal2 s 0 2219 624 2267 4 wl_1_4
rlabel metal2 s 0 2473 624 2521 4 wl_1_5
rlabel metal2 s 0 3009 624 3057 4 wl_1_6
rlabel metal2 s 0 3263 624 3311 4 wl_1_7
rlabel metal2 s 0 3799 624 3847 4 wl_1_8
rlabel metal2 s 0 4053 624 4101 4 wl_1_9
rlabel metal2 s 0 4589 624 4637 4 wl_1_10
rlabel metal2 s 0 4843 624 4891 4 wl_1_11
rlabel metal2 s 0 5379 624 5427 4 wl_1_12
rlabel metal2 s 0 5633 624 5681 4 wl_1_13
rlabel metal2 s 0 6169 624 6217 4 wl_1_14
rlabel metal2 s 0 6423 624 6471 4 wl_1_15
rlabel metal2 s 0 6959 624 7007 4 wl_1_16
rlabel metal2 s 0 7213 624 7261 4 wl_1_17
rlabel metal2 s 0 7749 624 7797 4 wl_1_18
rlabel metal2 s 0 8003 624 8051 4 wl_1_19
rlabel metal2 s 0 8539 624 8587 4 wl_1_20
rlabel metal2 s 0 8793 624 8841 4 wl_1_21
rlabel metal2 s 0 9329 624 9377 4 wl_1_22
rlabel metal2 s 0 9583 624 9631 4 wl_1_23
rlabel metal2 s 0 10119 624 10167 4 wl_1_24
rlabel metal2 s 0 10373 624 10421 4 wl_1_25
rlabel metal2 s 0 10909 624 10957 4 wl_1_26
rlabel metal2 s 0 11163 624 11211 4 wl_1_27
rlabel metal2 s 0 11699 624 11747 4 wl_1_28
rlabel metal2 s 0 11953 624 12001 4 wl_1_29
rlabel metal2 s 0 12489 624 12537 4 wl_1_30
rlabel metal2 s 0 12743 624 12791 4 wl_1_31
rlabel metal2 s 0 13279 624 13327 4 wl_1_32
rlabel metal2 s 0 13533 624 13581 4 wl_1_33
rlabel metal2 s 0 14069 624 14117 4 wl_1_34
rlabel metal2 s 0 14323 624 14371 4 wl_1_35
rlabel metal2 s 0 14859 624 14907 4 wl_1_36
rlabel metal2 s 0 15113 624 15161 4 wl_1_37
rlabel metal2 s 0 15649 624 15697 4 wl_1_38
rlabel metal2 s 0 15903 624 15951 4 wl_1_39
rlabel metal2 s 0 16439 624 16487 4 wl_1_40
rlabel metal2 s 0 16693 624 16741 4 wl_1_41
rlabel metal2 s 0 17229 624 17277 4 wl_1_42
rlabel metal2 s 0 17483 624 17531 4 wl_1_43
rlabel metal2 s 0 18019 624 18067 4 wl_1_44
rlabel metal2 s 0 18273 624 18321 4 wl_1_45
rlabel metal2 s 0 18809 624 18857 4 wl_1_46
rlabel metal2 s 0 19063 624 19111 4 wl_1_47
rlabel metal2 s 0 19599 624 19647 4 wl_1_48
rlabel metal2 s 0 19853 624 19901 4 wl_1_49
rlabel metal2 s 0 20389 624 20437 4 wl_1_50
rlabel metal2 s 0 20643 624 20691 4 wl_1_51
rlabel metal2 s 0 21179 624 21227 4 wl_1_52
rlabel metal2 s 0 21433 624 21481 4 wl_1_53
rlabel metal2 s 0 21969 624 22017 4 wl_1_54
rlabel metal2 s 0 22223 624 22271 4 wl_1_55
rlabel metal2 s 0 22759 624 22807 4 wl_1_56
rlabel metal2 s 0 23013 624 23061 4 wl_1_57
rlabel metal2 s 0 23549 624 23597 4 wl_1_58
rlabel metal2 s 0 23803 624 23851 4 wl_1_59
rlabel metal2 s 0 24339 624 24387 4 wl_1_60
rlabel metal2 s 0 24593 624 24641 4 wl_1_61
rlabel metal2 s 0 25129 624 25177 4 wl_1_62
rlabel metal2 s 0 25383 624 25431 4 wl_1_63
rlabel metal2 s 0 25919 624 25967 4 wl_1_64
rlabel metal2 s 0 26173 624 26221 4 wl_1_65
rlabel metal2 s 0 26709 624 26757 4 wl_1_66
rlabel metal2 s 0 26963 624 27011 4 wl_1_67
rlabel metal2 s 0 27499 624 27547 4 wl_1_68
rlabel metal2 s 0 27753 624 27801 4 wl_1_69
rlabel metal2 s 0 28289 624 28337 4 wl_1_70
rlabel metal2 s 0 28543 624 28591 4 wl_1_71
rlabel metal2 s 0 29079 624 29127 4 wl_1_72
rlabel metal2 s 0 29333 624 29381 4 wl_1_73
rlabel metal2 s 0 29869 624 29917 4 wl_1_74
rlabel metal2 s 0 30123 624 30171 4 wl_1_75
rlabel metal2 s 0 30659 624 30707 4 wl_1_76
rlabel metal2 s 0 30913 624 30961 4 wl_1_77
rlabel metal2 s 0 31449 624 31497 4 wl_1_78
rlabel metal2 s 0 31703 624 31751 4 wl_1_79
rlabel metal2 s 0 32239 624 32287 4 wl_1_80
rlabel metal2 s 0 32493 624 32541 4 wl_1_81
rlabel metal2 s 0 33029 624 33077 4 wl_1_82
rlabel metal2 s 0 33283 624 33331 4 wl_1_83
rlabel metal2 s 0 33819 624 33867 4 wl_1_84
rlabel metal2 s 0 34073 624 34121 4 wl_1_85
rlabel metal2 s 0 34609 624 34657 4 wl_1_86
rlabel metal2 s 0 34863 624 34911 4 wl_1_87
rlabel metal2 s 0 35399 624 35447 4 wl_1_88
rlabel metal2 s 0 35653 624 35701 4 wl_1_89
rlabel metal2 s 0 36189 624 36237 4 wl_1_90
rlabel metal2 s 0 36443 624 36491 4 wl_1_91
rlabel metal2 s 0 36979 624 37027 4 wl_1_92
rlabel metal2 s 0 37233 624 37281 4 wl_1_93
rlabel metal2 s 0 37769 624 37817 4 wl_1_94
rlabel metal2 s 0 38023 624 38071 4 wl_1_95
rlabel metal2 s 0 38559 624 38607 4 wl_1_96
rlabel metal2 s 0 38813 624 38861 4 wl_1_97
rlabel metal2 s 0 39349 624 39397 4 wl_1_98
rlabel metal2 s 0 39603 624 39651 4 wl_1_99
rlabel metal2 s 0 40139 624 40187 4 wl_1_100
rlabel metal2 s 0 40393 624 40441 4 wl_1_101
rlabel metal2 s 0 40929 624 40977 4 wl_1_102
rlabel metal2 s 0 41183 624 41231 4 wl_1_103
rlabel metal2 s 0 41719 624 41767 4 wl_1_104
rlabel metal2 s 0 41973 624 42021 4 wl_1_105
rlabel metal2 s 0 42509 624 42557 4 wl_1_106
rlabel metal2 s 0 42763 624 42811 4 wl_1_107
rlabel metal2 s 0 43299 624 43347 4 wl_1_108
rlabel metal2 s 0 43553 624 43601 4 wl_1_109
rlabel metal2 s 0 44089 624 44137 4 wl_1_110
rlabel metal2 s 0 44343 624 44391 4 wl_1_111
rlabel metal2 s 0 44879 624 44927 4 wl_1_112
rlabel metal2 s 0 45133 624 45181 4 wl_1_113
rlabel metal2 s 0 45669 624 45717 4 wl_1_114
rlabel metal2 s 0 45923 624 45971 4 wl_1_115
rlabel metal2 s 0 46459 624 46507 4 wl_1_116
rlabel metal2 s 0 46713 624 46761 4 wl_1_117
rlabel metal2 s 0 47249 624 47297 4 wl_1_118
rlabel metal2 s 0 47503 624 47551 4 wl_1_119
rlabel metal2 s 0 48039 624 48087 4 wl_1_120
rlabel metal2 s 0 48293 624 48341 4 wl_1_121
rlabel metal2 s 0 48829 624 48877 4 wl_1_122
rlabel metal2 s 0 49083 624 49131 4 wl_1_123
rlabel metal2 s 0 49619 624 49667 4 wl_1_124
rlabel metal2 s 0 49873 624 49921 4 wl_1_125
rlabel metal2 s 0 50409 624 50457 4 wl_1_126
rlabel metal2 s 0 50663 624 50711 4 wl_1_127
rlabel metal2 s 0 51199 624 51247 4 wl_1_128
rlabel metal2 s 0 51453 624 51501 4 wl_1_129
rlabel metal2 s 0 51989 624 52037 4 wl_1_130
rlabel metal2 s 0 52243 624 52291 4 wl_1_131
rlabel metal2 s 0 52779 624 52827 4 wl_1_132
rlabel metal2 s 0 53033 624 53081 4 wl_1_133
rlabel metal2 s 0 53569 624 53617 4 wl_1_134
rlabel metal2 s 0 53823 624 53871 4 wl_1_135
rlabel metal2 s 0 54359 624 54407 4 wl_1_136
rlabel metal2 s 0 54613 624 54661 4 wl_1_137
rlabel metal2 s 0 55149 624 55197 4 wl_1_138
rlabel metal2 s 0 55403 624 55451 4 wl_1_139
rlabel metal2 s 0 55939 624 55987 4 wl_1_140
rlabel metal2 s 0 56193 624 56241 4 wl_1_141
rlabel metal2 s 0 56729 624 56777 4 wl_1_142
rlabel metal2 s 0 56983 624 57031 4 wl_1_143
rlabel metal2 s 0 57519 624 57567 4 wl_1_144
rlabel metal2 s 0 57773 624 57821 4 wl_1_145
rlabel metal2 s 0 58309 624 58357 4 wl_1_146
rlabel metal2 s 0 58563 624 58611 4 wl_1_147
rlabel metal2 s 0 59099 624 59147 4 wl_1_148
rlabel metal2 s 0 59353 624 59401 4 wl_1_149
rlabel metal2 s 0 59889 624 59937 4 wl_1_150
rlabel metal2 s 0 60143 624 60191 4 wl_1_151
rlabel metal2 s 0 60679 624 60727 4 wl_1_152
rlabel metal2 s 0 60933 624 60981 4 wl_1_153
rlabel metal2 s 0 61469 624 61517 4 wl_1_154
rlabel metal2 s 0 61723 624 61771 4 wl_1_155
rlabel metal2 s 0 62259 624 62307 4 wl_1_156
rlabel metal2 s 0 62513 624 62561 4 wl_1_157
rlabel metal2 s 0 63049 624 63097 4 wl_1_158
rlabel metal2 s 0 63303 624 63351 4 wl_1_159
rlabel metal2 s 0 63839 624 63887 4 wl_1_160
rlabel metal2 s 0 64093 624 64141 4 wl_1_161
rlabel metal2 s 0 64629 624 64677 4 wl_1_162
rlabel metal2 s 0 64883 624 64931 4 wl_1_163
rlabel metal2 s 0 65419 624 65467 4 wl_1_164
rlabel metal2 s 0 65673 624 65721 4 wl_1_165
rlabel metal2 s 0 66209 624 66257 4 wl_1_166
rlabel metal2 s 0 66463 624 66511 4 wl_1_167
rlabel metal2 s 0 66999 624 67047 4 wl_1_168
rlabel metal2 s 0 67253 624 67301 4 wl_1_169
rlabel metal2 s 0 67789 624 67837 4 wl_1_170
rlabel metal2 s 0 68043 624 68091 4 wl_1_171
rlabel metal2 s 0 68579 624 68627 4 wl_1_172
rlabel metal2 s 0 68833 624 68881 4 wl_1_173
rlabel metal2 s 0 69369 624 69417 4 wl_1_174
rlabel metal2 s 0 69623 624 69671 4 wl_1_175
rlabel metal2 s 0 70159 624 70207 4 wl_1_176
rlabel metal2 s 0 70413 624 70461 4 wl_1_177
rlabel metal2 s 0 70949 624 70997 4 wl_1_178
rlabel metal2 s 0 71203 624 71251 4 wl_1_179
rlabel metal2 s 0 71739 624 71787 4 wl_1_180
rlabel metal2 s 0 71993 624 72041 4 wl_1_181
rlabel metal2 s 0 72529 624 72577 4 wl_1_182
rlabel metal2 s 0 72783 624 72831 4 wl_1_183
rlabel metal2 s 0 73319 624 73367 4 wl_1_184
rlabel metal2 s 0 73573 624 73621 4 wl_1_185
rlabel metal2 s 0 74109 624 74157 4 wl_1_186
rlabel metal2 s 0 74363 624 74411 4 wl_1_187
rlabel metal2 s 0 74899 624 74947 4 wl_1_188
rlabel metal2 s 0 75153 624 75201 4 wl_1_189
rlabel metal2 s 0 75689 624 75737 4 wl_1_190
rlabel metal2 s 0 75943 624 75991 4 wl_1_191
rlabel metal2 s 0 76479 624 76527 4 wl_1_192
rlabel metal2 s 0 76733 624 76781 4 wl_1_193
rlabel metal2 s 0 77269 624 77317 4 wl_1_194
rlabel metal2 s 0 77523 624 77571 4 wl_1_195
rlabel metal2 s 0 78059 624 78107 4 wl_1_196
rlabel metal2 s 0 78313 624 78361 4 wl_1_197
rlabel metal2 s 0 78849 624 78897 4 wl_1_198
rlabel metal2 s 0 79103 624 79151 4 wl_1_199
rlabel metal2 s 0 79639 624 79687 4 wl_1_200
rlabel metal2 s 0 79893 624 79941 4 wl_1_201
rlabel metal2 s 0 80429 624 80477 4 wl_1_202
rlabel metal2 s 0 80683 624 80731 4 wl_1_203
rlabel metal2 s 0 81219 624 81267 4 wl_1_204
rlabel metal2 s 0 81473 624 81521 4 wl_1_205
rlabel metal2 s 0 82009 624 82057 4 wl_1_206
rlabel metal2 s 0 82263 624 82311 4 wl_1_207
rlabel metal2 s 0 82799 624 82847 4 wl_1_208
rlabel metal2 s 0 83053 624 83101 4 wl_1_209
rlabel metal2 s 0 83589 624 83637 4 wl_1_210
rlabel metal2 s 0 83843 624 83891 4 wl_1_211
rlabel metal2 s 0 84379 624 84427 4 wl_1_212
rlabel metal2 s 0 84633 624 84681 4 wl_1_213
rlabel metal2 s 0 85169 624 85217 4 wl_1_214
rlabel metal2 s 0 85423 624 85471 4 wl_1_215
rlabel metal2 s 0 85959 624 86007 4 wl_1_216
rlabel metal2 s 0 86213 624 86261 4 wl_1_217
rlabel metal2 s 0 86749 624 86797 4 wl_1_218
rlabel metal2 s 0 87003 624 87051 4 wl_1_219
rlabel metal2 s 0 87539 624 87587 4 wl_1_220
rlabel metal2 s 0 87793 624 87841 4 wl_1_221
rlabel metal2 s 0 88329 624 88377 4 wl_1_222
rlabel metal2 s 0 88583 624 88631 4 wl_1_223
rlabel metal2 s 0 89119 624 89167 4 wl_1_224
rlabel metal2 s 0 89373 624 89421 4 wl_1_225
rlabel metal2 s 0 89909 624 89957 4 wl_1_226
rlabel metal2 s 0 90163 624 90211 4 wl_1_227
rlabel metal2 s 0 90699 624 90747 4 wl_1_228
rlabel metal2 s 0 90953 624 91001 4 wl_1_229
rlabel metal2 s 0 91489 624 91537 4 wl_1_230
rlabel metal2 s 0 91743 624 91791 4 wl_1_231
rlabel metal2 s 0 92279 624 92327 4 wl_1_232
rlabel metal2 s 0 92533 624 92581 4 wl_1_233
rlabel metal2 s 0 93069 624 93117 4 wl_1_234
rlabel metal2 s 0 93323 624 93371 4 wl_1_235
rlabel metal2 s 0 93859 624 93907 4 wl_1_236
rlabel metal2 s 0 94113 624 94161 4 wl_1_237
rlabel metal2 s 0 94649 624 94697 4 wl_1_238
rlabel metal2 s 0 94903 624 94951 4 wl_1_239
rlabel metal2 s 0 95439 624 95487 4 wl_1_240
rlabel metal2 s 0 95693 624 95741 4 wl_1_241
rlabel metal2 s 0 96229 624 96277 4 wl_1_242
rlabel metal2 s 0 96483 624 96531 4 wl_1_243
rlabel metal2 s 0 97019 624 97067 4 wl_1_244
rlabel metal2 s 0 97273 624 97321 4 wl_1_245
rlabel metal2 s 0 97809 624 97857 4 wl_1_246
rlabel metal2 s 0 98063 624 98111 4 wl_1_247
rlabel metal2 s 0 98599 624 98647 4 wl_1_248
rlabel metal2 s 0 98853 624 98901 4 wl_1_249
rlabel metal2 s 0 99389 624 99437 4 wl_1_250
rlabel metal2 s 0 99643 624 99691 4 wl_1_251
rlabel metal2 s 0 100179 624 100227 4 wl_1_252
rlabel metal2 s 0 100433 624 100481 4 wl_1_253
rlabel metal2 s 0 100969 624 101017 4 wl_1_254
rlabel metal2 s 0 101223 624 101271 4 wl_1_255
rlabel metal2 s 0 101759 624 101807 4 wl_1_256
rlabel metal2 s 0 102013 624 102061 4 wl_1_257
rlabel metal1 s 222 61990 258 62331 4 vdd
rlabel metal1 s 222 69599 258 69940 4 vdd
rlabel metal1 s 222 51720 258 52061 4 vdd
rlabel metal1 s 222 56460 258 56801 4 vdd
rlabel metal1 s 222 45109 258 45450 4 vdd
rlabel metal1 s 222 88559 258 88900 4 vdd
rlabel metal1 s 222 24569 258 24910 4 vdd
rlabel metal1 s 222 98330 258 98671 4 vdd
rlabel metal1 s 222 43529 258 43870 4 vdd
rlabel metal1 s 222 28810 258 29151 4 vdd
rlabel metal1 s 222 13509 258 13850 4 vdd
rlabel metal1 s 222 45899 258 46240 4 vdd
rlabel metal1 s 222 80659 258 81000 4 vdd
rlabel metal1 s 222 81449 258 81790 4 vdd
rlabel metal1 s 222 83819 258 84160 4 vdd
rlabel metal1 s 222 4029 258 4370 4 vdd
rlabel metal1 s 222 46980 258 47321 4 vdd
rlabel metal1 s 222 83029 258 83370 4 vdd
rlabel metal1 s 222 95669 258 96010 4 vdd
rlabel metal1 s 222 72759 258 73100 4 vdd
rlabel metal1 s 222 19829 258 20170 4 vdd
rlabel metal1 s 222 24860 258 25201 4 vdd
rlabel metal1 s 222 17459 258 17800 4 vdd
rlabel metal1 s 222 56959 258 57300 4 vdd
rlabel metal1 s 222 101199 258 101540 4 vdd
rlabel metal1 s 222 6399 258 6740 4 vdd
rlabel metal1 s 222 57749 258 58090 4 vdd
rlabel metal1 s 222 11430 258 11771 4 vdd
rlabel metal1 s 222 26939 258 27280 4 vdd
rlabel metal1 s 222 69100 258 69441 4 vdd
rlabel metal1 s 222 8769 258 9110 4 vdd
rlabel metal1 s 222 75129 258 75470 4 vdd
rlabel metal1 s 222 30889 258 31230 4 vdd
rlabel metal1 s 222 84110 258 84451 4 vdd
rlabel metal1 s 222 53300 258 53641 4 vdd
rlabel metal1 s 222 77000 258 77341 4 vdd
rlabel metal1 s 222 31679 258 32020 4 vdd
rlabel metal1 s 222 26440 258 26781 4 vdd
rlabel metal1 s 222 20910 258 21251 4 vdd
rlabel metal1 s 222 34340 258 34681 4 vdd
rlabel metal1 s 222 91220 258 91561 4 vdd
rlabel metal1 s 222 29309 258 29650 4 vdd
rlabel metal1 s 222 37500 258 37841 4 vdd
rlabel metal1 s 222 57250 258 57591 4 vdd
rlabel metal1 s 222 20120 258 20461 4 vdd
rlabel metal1 s 222 79079 258 79420 4 vdd
rlabel metal1 s 222 18540 258 18881 4 vdd
rlabel metal1 s 222 98039 258 98380 4 vdd
rlabel metal1 s 222 22989 258 23330 4 vdd
rlabel metal1 s 222 60410 258 60751 4 vdd
rlabel metal1 s 222 869 258 1210 4 vdd
rlabel metal1 s 222 30390 258 30731 4 vdd
rlabel metal1 s 222 5110 258 5451 4 vdd
rlabel metal1 s 222 8270 258 8611 4 vdd
rlabel metal1 s 222 38290 258 38631 4 vdd
rlabel metal1 s 222 68809 258 69150 4 vdd
rlabel metal1 s 222 94380 258 94721 4 vdd
rlabel metal1 s 222 97249 258 97590 4 vdd
rlabel metal1 s 222 4819 258 5160 4 vdd
rlabel metal3 s 263 180 361 278 4 vdd
rlabel metal1 s 222 10349 258 10690 4 vdd
rlabel metal1 s 222 77790 258 78131 4 vdd
rlabel metal1 s 222 88060 258 88401 4 vdd
rlabel metal1 s 222 96750 258 97091 4 vdd
rlabel metal1 s 222 98829 258 99170 4 vdd
rlabel metal1 s 222 37209 258 37550 4 vdd
rlabel metal1 s 222 79869 258 80210 4 vdd
rlabel metal1 s 222 11139 258 11480 4 vdd
rlabel metal1 s 222 3239 258 3580 4 vdd
rlabel metal1 s 222 42240 258 42581 4 vdd
rlabel metal1 s 222 64069 258 64410 4 vdd
rlabel metal1 s 222 89640 258 89981 4 vdd
rlabel metal1 s 222 7979 258 8320 4 vdd
rlabel metal1 s 222 36419 258 36760 4 vdd
rlabel metal1 s 222 74339 258 74680 4 vdd
rlabel metal1 s 222 94089 258 94430 4 vdd
rlabel metal1 s 222 95960 258 96301 4 vdd
rlabel metal1 s 222 100409 258 100750 4 vdd
rlabel metal1 s 222 58830 258 59171 4 vdd
rlabel metal1 s 222 76709 258 77050 4 vdd
rlabel metal1 s 222 47479 258 47820 4 vdd
rlabel metal1 s 222 54880 258 55221 4 vdd
rlabel metal1 s 222 36710 258 37051 4 vdd
rlabel metal1 s 222 62489 258 62830 4 vdd
rlabel metal1 s 222 70680 258 71021 4 vdd
rlabel metal1 s 222 71470 258 71811 4 vdd
rlabel metal1 s 222 69890 258 70231 4 vdd
rlabel metal1 s 222 23779 258 24120 4 vdd
rlabel metal1 s 222 16170 258 16511 4 vdd
rlabel metal1 s 222 46190 258 46531 4 vdd
rlabel metal1 s 222 64360 258 64701 4 vdd
rlabel metal1 s 222 68019 258 68360 4 vdd
rlabel metal1 s 222 75919 258 76260 4 vdd
rlabel metal1 s 222 93590 258 93931 4 vdd
rlabel metal1 s 222 78580 258 78921 4 vdd
rlabel metal1 s 222 34839 258 35180 4 vdd
rlabel metal1 s 222 99910 258 100251 4 vdd
rlabel metal1 s 222 23280 258 23621 4 vdd
rlabel metal1 s 222 49059 258 49400 4 vdd
rlabel metal1 s 222 65940 258 66281 4 vdd
rlabel metal1 s 222 44319 258 44660 4 vdd
rlabel metal1 s 222 20619 258 20960 4 vdd
rlabel metal1 s 222 99619 258 99960 4 vdd
rlabel metal1 s 222 84900 258 85241 4 vdd
rlabel metal1 s 222 12719 258 13060 4 vdd
rlabel metal1 s 222 86480 258 86821 4 vdd
rlabel metal1 s 222 5609 258 5950 4 vdd
rlabel metal1 s 222 2740 258 3081 4 vdd
rlabel metal1 s 222 76210 258 76551 4 vdd
rlabel metal1 s 222 62780 258 63121 4 vdd
rlabel metal1 s 222 71179 258 71520 4 vdd
rlabel metal1 s 222 34049 258 34390 4 vdd
rlabel metal1 s 222 41159 258 41500 4 vdd
rlabel metal1 s 222 53799 258 54140 4 vdd
rlabel metal1 s 222 59620 258 59961 4 vdd
rlabel metal1 s 222 44610 258 44951 4 vdd
rlabel metal1 s 222 88850 258 89191 4 vdd
rlabel metal1 s 222 89349 258 89690 4 vdd
rlabel metal1 s 222 37999 258 38340 4 vdd
rlabel metal1 s 222 78289 258 78630 4 vdd
rlabel metal1 s 222 22199 258 22540 4 vdd
rlabel metal1 s 222 39870 258 40211 4 vdd
rlabel metal1 s 222 54090 258 54431 4 vdd
rlabel metal1 s 222 83320 258 83661 4 vdd
rlabel metal1 s 222 45400 258 45741 4 vdd
rlabel metal1 s 222 14299 258 14640 4 vdd
rlabel metal1 s 222 5900 258 6241 4 vdd
rlabel metal1 s 222 19039 258 19380 4 vdd
rlabel metal1 s 222 35629 258 35970 4 vdd
rlabel metal1 s 222 71969 258 72310 4 vdd
rlabel metal1 s 222 86979 258 87320 4 vdd
rlabel metal1 s 222 93299 258 93640 4 vdd
rlabel metal1 s 222 15879 258 16220 4 vdd
rlabel metal1 s 222 94879 258 95220 4 vdd
rlabel metal1 s 222 101989 258 102330 4 vdd
rlabel metal1 s 222 370 258 711 4 vdd
rlabel metal1 s 222 51429 258 51770 4 vdd
rlabel metal1 s 222 28020 258 28361 4 vdd
rlabel metal1 s 222 55670 258 56011 4 vdd
rlabel metal1 s 222 61200 258 61541 4 vdd
rlabel metal1 s 222 18249 258 18590 4 vdd
rlabel metal1 s 222 41450 258 41791 4 vdd
rlabel metal1 s 222 74630 258 74971 4 vdd
rlabel metal1 s 222 39080 258 39421 4 vdd
rlabel metal1 s 222 35130 258 35471 4 vdd
rlabel metal1 s 222 6690 258 7031 4 vdd
rlabel metal1 s 222 50639 258 50980 4 vdd
rlabel metal1 s 222 90139 258 90480 4 vdd
rlabel metal1 s 222 68310 258 68651 4 vdd
rlabel metal1 s 222 66439 258 66780 4 vdd
rlabel metal1 s 222 50930 258 51271 4 vdd
rlabel metal1 s 222 86189 258 86530 4 vdd
rlabel metal3 s 263 102422 361 102520 4 vdd
rlabel metal1 s 222 63279 258 63620 4 vdd
rlabel metal1 s 222 29600 258 29941 4 vdd
rlabel metal1 s 222 17750 258 18091 4 vdd
rlabel metal1 s 222 2449 258 2790 4 vdd
rlabel metal1 s 222 67520 258 67861 4 vdd
rlabel metal1 s 222 95170 258 95511 4 vdd
rlabel metal1 s 222 7480 258 7821 4 vdd
rlabel metal1 s 222 92010 258 92351 4 vdd
rlabel metal1 s 222 64859 258 65200 4 vdd
rlabel metal1 s 222 72260 258 72601 4 vdd
rlabel metal1 s 222 11929 258 12270 4 vdd
rlabel metal1 s 222 32760 258 33101 4 vdd
rlabel metal1 s 222 12220 258 12561 4 vdd
rlabel metal1 s 222 82530 258 82871 4 vdd
rlabel metal1 s 222 24070 258 24411 4 vdd
rlabel metal1 s 222 38789 258 39130 4 vdd
rlabel metal1 s 222 91719 258 92060 4 vdd
rlabel metal1 s 222 42739 258 43080 4 vdd
rlabel metal1 s 222 40660 258 41001 4 vdd
rlabel metal1 s 222 50140 258 50481 4 vdd
rlabel metal1 s 222 21700 258 22041 4 vdd
rlabel metal1 s 222 22490 258 22831 4 vdd
rlabel metal1 s 222 48269 258 48610 4 vdd
rlabel metal1 s 222 13800 258 14141 4 vdd
rlabel metal1 s 222 49849 258 50190 4 vdd
rlabel metal1 s 222 52219 258 52560 4 vdd
rlabel metal1 s 222 96459 258 96800 4 vdd
rlabel metal1 s 222 43030 258 43371 4 vdd
rlabel metal1 s 222 66730 258 67071 4 vdd
rlabel metal1 s 222 73840 258 74181 4 vdd
rlabel metal1 s 222 99120 258 99461 4 vdd
rlabel metal1 s 222 49350 258 49691 4 vdd
rlabel metal1 s 222 100700 258 101041 4 vdd
rlabel metal1 s 222 90929 258 91270 4 vdd
rlabel metal1 s 222 65649 258 65990 4 vdd
rlabel metal1 s 222 97540 258 97881 4 vdd
rlabel metal1 s 222 9850 258 10191 4 vdd
rlabel metal1 s 222 9559 258 9900 4 vdd
rlabel metal1 s 222 25650 258 25991 4 vdd
rlabel metal1 s 222 80950 258 81291 4 vdd
rlabel metal1 s 222 35920 258 36261 4 vdd
rlabel metal1 s 222 82239 258 82580 4 vdd
rlabel metal1 s 222 31180 258 31521 4 vdd
rlabel metal1 s 222 1160 258 1501 4 vdd
rlabel metal1 s 222 1950 258 2291 4 vdd
rlabel metal1 s 222 80160 258 80501 4 vdd
rlabel metal1 s 222 30099 258 30440 4 vdd
rlabel metal1 s 222 47770 258 48111 4 vdd
rlabel metal1 s 222 73050 258 73391 4 vdd
rlabel metal1 s 222 81740 258 82081 4 vdd
rlabel metal1 s 222 85399 258 85740 4 vdd
rlabel metal1 s 222 87769 258 88110 4 vdd
rlabel metal1 s 222 63570 258 63911 4 vdd
rlabel metal1 s 222 55379 258 55720 4 vdd
rlabel metal1 s 222 9060 258 9401 4 vdd
rlabel metal1 s 222 101490 258 101831 4 vdd
rlabel metal1 s 222 87270 258 87611 4 vdd
rlabel metal1 s 222 53009 258 53350 4 vdd
rlabel metal1 s 222 13010 258 13351 4 vdd
rlabel metal1 s 222 28519 258 28860 4 vdd
rlabel metal1 s 222 40369 258 40710 4 vdd
rlabel metal1 s 222 67229 258 67570 4 vdd
rlabel metal1 s 222 70389 258 70730 4 vdd
rlabel metal1 s 222 75420 258 75761 4 vdd
rlabel metal1 s 222 77499 258 77840 4 vdd
rlabel metal1 s 222 1659 258 2000 4 vdd
rlabel metal1 s 222 3530 258 3871 4 vdd
rlabel metal1 s 222 4320 258 4661 4 vdd
rlabel metal1 s 222 65150 258 65491 4 vdd
rlabel metal1 s 222 33259 258 33600 4 vdd
rlabel metal1 s 222 41949 258 42290 4 vdd
rlabel metal1 s 222 59329 258 59670 4 vdd
rlabel metal1 s 222 26149 258 26490 4 vdd
rlabel metal1 s 222 48560 258 48901 4 vdd
rlabel metal1 s 222 21409 258 21750 4 vdd
rlabel metal1 s 222 58539 258 58880 4 vdd
rlabel metal1 s 222 10640 258 10981 4 vdd
rlabel metal1 s 222 46689 258 47030 4 vdd
rlabel metal1 s 222 31970 258 32311 4 vdd
rlabel metal1 s 222 60119 258 60460 4 vdd
rlabel metal1 s 222 73549 258 73890 4 vdd
rlabel metal1 s 222 92800 258 93141 4 vdd
rlabel metal1 s 222 79370 258 79711 4 vdd
rlabel metal1 s 222 85690 258 86031 4 vdd
rlabel metal1 s 222 25359 258 25700 4 vdd
rlabel metal1 s 222 15380 258 15721 4 vdd
rlabel metal1 s 222 92509 258 92850 4 vdd
rlabel metal1 s 222 52510 258 52851 4 vdd
rlabel metal1 s 222 58040 258 58381 4 vdd
rlabel metal1 s 222 60909 258 61250 4 vdd
rlabel metal1 s 222 27230 258 27571 4 vdd
rlabel metal1 s 222 39579 258 39920 4 vdd
rlabel metal1 s 222 19330 258 19671 4 vdd
rlabel metal1 s 222 90430 258 90771 4 vdd
rlabel metal1 s 222 33550 258 33891 4 vdd
rlabel metal1 s 222 7189 258 7530 4 vdd
rlabel metal1 s 222 32469 258 32810 4 vdd
rlabel metal1 s 222 61699 258 62040 4 vdd
rlabel metal1 s 222 14590 258 14931 4 vdd
rlabel metal1 s 222 15089 258 15430 4 vdd
rlabel metal1 s 222 54589 258 54930 4 vdd
rlabel metal1 s 222 56169 258 56510 4 vdd
rlabel metal1 s 222 84609 258 84950 4 vdd
rlabel metal1 s 222 43820 258 44161 4 vdd
rlabel metal1 s 222 27729 258 28070 4 vdd
rlabel metal1 s 222 16669 258 17010 4 vdd
rlabel metal1 s 222 16960 258 17301 4 vdd
rlabel metal2 s 186 62609 294 62685 4 gnd
rlabel metal2 s 186 76355 294 76431 4 gnd
rlabel metal2 s 186 19695 294 19805 4 gnd
rlabel metal2 s 186 56035 294 56145 4 gnd
rlabel metal2 s 186 73195 294 73271 4 gnd
rlabel metal2 s 186 4149 294 4225 4 gnd
rlabel metal2 s 186 67665 294 67741 4 gnd
rlabel metal2 s 186 10215 294 10325 4 gnd
rlabel metal2 s 186 56289 294 56365 4 gnd
rlabel metal2 s 186 44439 294 44515 4 gnd
rlabel metal2 s 186 15745 294 15855 4 gnd
rlabel metal2 s 186 40235 294 40345 4 gnd
rlabel metal2 s 186 1305 294 1381 4 gnd
rlabel metal2 s 186 57079 294 57155 4 gnd
rlabel metal2 s 186 99485 294 99595 4 gnd
rlabel metal2 s 186 13945 294 14021 4 gnd
rlabel metal2 s 186 39699 294 39775 4 gnd
rlabel metal2 s 186 19949 294 20025 4 gnd
rlabel metal2 s 186 87415 294 87491 4 gnd
rlabel metal2 s 186 48135 294 48245 4 gnd
rlabel metal2 s 186 71299 294 71375 4 gnd
rlabel metal2 s 186 33379 294 33455 4 gnd
rlabel metal2 s 186 32589 294 32665 4 gnd
rlabel metal2 s 186 78409 294 78485 4 gnd
rlabel metal2 s 186 49495 294 49571 4 gnd
rlabel metal2 s 186 92155 294 92231 4 gnd
rlabel metal2 s 186 86309 294 86385 4 gnd
rlabel metal2 s 186 94999 294 95075 4 gnd
rlabel metal2 s 186 29745 294 29821 4 gnd
rlabel metal2 s 186 44975 294 45085 4 gnd
rlabel metal2 s 186 64189 294 64265 4 gnd
rlabel metal2 s 186 2095 294 2171 4 gnd
rlabel metal2 s 186 7309 294 7385 4 gnd
rlabel metal2 s 186 27595 294 27705 4 gnd
rlabel metal2 s 186 11005 294 11115 4 gnd
rlabel metal2 s 186 45545 294 45621 4 gnd
rlabel metal2 s 186 62135 294 62211 4 gnd
rlabel metal2 s 186 91365 294 91441 4 gnd
rlabel metal2 s 186 16535 294 16645 4 gnd
rlabel metal2 s 186 87889 294 87965 4 gnd
rlabel metal2 s 186 515 294 591 4 gnd
rlabel metal2 s 186 67095 294 67205 4 gnd
rlabel metal2 s 186 79199 294 79275 4 gnd
rlabel metal2 s 186 90575 294 90651 4 gnd
rlabel metal2 s 186 17105 294 17181 4 gnd
rlabel metal2 s 186 76039 294 76115 4 gnd
rlabel metal2 s 186 37075 294 37185 4 gnd
rlabel metal2 s 186 43395 294 43505 4 gnd
rlabel metal2 s 186 39225 294 39301 4 gnd
rlabel metal2 s 186 13155 294 13231 4 gnd
rlabel metal2 s 186 82105 294 82215 4 gnd
rlabel metal2 s 186 67349 294 67425 4 gnd
rlabel metal2 s 186 75565 294 75641 4 gnd
rlabel metal2 s 186 91049 294 91125 4 gnd
rlabel metal2 s 186 50759 294 50835 4 gnd
rlabel metal2 s 186 1779 294 1855 4 gnd
rlabel metal2 s 186 57615 294 57725 4 gnd
rlabel metal2 s 186 84475 294 84585 4 gnd
rlabel metal2 s 186 81095 294 81171 4 gnd
rlabel metal2 s 186 15525 294 15601 4 gnd
rlabel metal2 s 186 3675 294 3751 4 gnd
rlabel metal2 s 186 53665 294 53775 4 gnd
rlabel metal2 s 186 93955 294 94065 4 gnd
rlabel metal2 s 186 9995 294 10071 4 gnd
rlabel metal2 s 186 26805 294 26915 4 gnd
rlabel metal2 s 186 19159 294 19235 4 gnd
rlabel metal2 s 186 88205 294 88281 4 gnd
rlabel metal2 s 186 97905 294 98015 4 gnd
rlabel metal2 s 186 100845 294 100921 4 gnd
rlabel metal2 s 186 61819 294 61895 4 gnd
rlabel metal2 s 186 69245 294 69321 4 gnd
rlabel metal2 s 186 53445 294 53521 4 gnd
rlabel metal2 s 186 43175 294 43251 4 gnd
rlabel metal2 s 186 47345 294 47455 4 gnd
rlabel metal2 s 186 87635 294 87745 4 gnd
rlabel metal2 s 186 35275 294 35351 4 gnd
rlabel metal2 s 186 65295 294 65371 4 gnd
rlabel metal2 s 186 29175 294 29285 4 gnd
rlabel metal2 s 186 39445 294 39555 4 gnd
rlabel metal2 s 186 80525 294 80635 4 gnd
rlabel metal2 s 186 65769 294 65845 4 gnd
rlabel metal2 s 186 36285 294 36395 4 gnd
rlabel metal2 s 186 72625 294 72735 4 gnd
rlabel metal2 s 186 35495 294 35605 4 gnd
rlabel metal2 s 186 4685 294 4795 4 gnd
rlabel metal2 s 186 74995 294 75105 4 gnd
rlabel metal2 s 186 989 294 1065 4 gnd
rlabel metal2 s 186 2569 294 2645 4 gnd
rlabel metal2 s 186 91839 294 91915 4 gnd
rlabel metal2 s 186 41025 294 41135 4 gnd
rlabel metal2 s 186 88995 294 89071 4 gnd
rlabel metal2 s 186 21529 294 21605 4 gnd
rlabel metal2 s 186 9205 294 9281 4 gnd
rlabel metal2 s 186 8099 294 8175 4 gnd
rlabel metal2 s 186 12365 294 12441 4 gnd
rlabel metal2 s 186 86845 294 86955 4 gnd
rlabel metal2 s 186 77145 294 77221 4 gnd
rlabel metal2 s 186 20739 294 20815 4 gnd
rlabel metal2 s 186 3895 294 4005 4 gnd
rlabel metal2 s 186 5475 294 5585 4 gnd
rlabel metal2 s 186 86055 294 86165 4 gnd
rlabel metal2 s 186 18369 294 18445 4 gnd
rlabel metal2 s 186 6265 294 6375 4 gnd
rlabel metal2 s 186 84255 294 84331 4 gnd
rlabel metal2 s 186 28639 294 28715 4 gnd
rlabel metal2 s 186 88679 294 88755 4 gnd
rlabel metal2 s 186 42069 294 42145 4 gnd
rlabel metal2 s 186 71045 294 71155 4 gnd
rlabel metal2 s 186 63715 294 63791 4 gnd
rlabel metal2 s 186 49969 294 50045 4 gnd
rlabel metal2 s 186 74205 294 74315 4 gnd
rlabel metal2 s 186 75785 294 75895 4 gnd
rlabel metal2 s 186 98475 294 98551 4 gnd
rlabel metal2 s 186 58659 294 58735 4 gnd
rlabel metal2 s 186 51549 294 51625 4 gnd
rlabel metal2 s 186 68929 294 69005 4 gnd
rlabel metal2 s 186 6835 294 6911 4 gnd
rlabel metal2 s 186 12585 294 12695 4 gnd
rlabel metal2 s 186 25005 294 25081 4 gnd
rlabel metal2 s 186 27849 294 27925 4 gnd
rlabel metal2 s 186 14419 294 14495 4 gnd
rlabel metal2 s 186 94209 294 94285 4 gnd
rlabel metal2 s 186 101855 294 101965 4 gnd
rlabel metal2 s 186 59765 294 59841 4 gnd
rlabel metal2 s 186 47599 294 47675 4 gnd
rlabel metal2 s 186 86625 294 86701 4 gnd
rlabel metal2 s 186 57395 294 57471 4 gnd
rlabel metal2 s 186 27059 294 27135 4 gnd
rlabel metal2 s 186 4465 294 4541 4 gnd
rlabel metal2 s 186 74775 294 74851 4 gnd
rlabel metal2 s 186 47915 294 47991 4 gnd
rlabel metal2 s 186 60239 294 60315 4 gnd
rlabel metal2 s 186 85265 294 85375 4 gnd
rlabel metal2 s 186 32905 294 32981 4 gnd
rlabel metal2 s 186 66559 294 66635 4 gnd
rlabel metal2 s 186 61029 294 61105 4 gnd
rlabel metal2 s 186 70255 294 70365 4 gnd
rlabel metal2 s 186 89469 294 89545 4 gnd
rlabel metal2 s 186 83685 294 83795 4 gnd
rlabel metal2 s 186 75249 294 75325 4 gnd
rlabel metal2 s 186 14165 294 14275 4 gnd
rlabel metal2 s 186 735 294 845 4 gnd
rlabel metal2 s 186 21275 294 21385 4 gnd
rlabel metal2 s 186 55815 294 55891 4 gnd
rlabel metal2 s 186 46335 294 46411 4 gnd
rlabel metal2 s 186 24215 294 24291 4 gnd
rlabel metal2 s 186 83149 294 83225 4 gnd
rlabel metal2 s 186 52655 294 52731 4 gnd
rlabel metal2 s 186 6045 294 6121 4 gnd
rlabel metal2 s 186 79515 294 79591 4 gnd
rlabel metal2 s 186 34169 294 34245 4 gnd
rlabel metal2 s 186 48389 294 48465 4 gnd
rlabel metal2 s 186 96895 294 96971 4 gnd
rlabel metal2 s 186 52085 294 52195 4 gnd
rlabel metal2 s 186 61565 294 61675 4 gnd
rlabel metal2 s 186 78945 294 79055 4 gnd
rlabel metal2 s 186 64979 294 65055 4 gnd
rlabel metal2 s 186 81315 294 81425 4 gnd
rlabel metal2 s 186 92945 294 93021 4 gnd
rlabel metal2 s 186 37645 294 37721 4 gnd
rlabel metal2 s 186 99265 294 99341 4 gnd
rlabel metal2 s 186 55499 294 55575 4 gnd
rlabel metal2 s 186 11575 294 11651 4 gnd
rlabel metal2 s 186 36539 294 36615 4 gnd
rlabel metal2 s 186 23425 294 23501 4 gnd
rlabel metal2 s 186 25225 294 25335 4 gnd
rlabel metal2 s 186 31545 294 31655 4 gnd
rlabel metal2 s 186 45765 294 45875 4 gnd
rlabel metal2 s 186 101065 294 101175 4 gnd
rlabel metal2 s 186 12839 294 12915 4 gnd
rlabel metal2 s 186 2885 294 2961 4 gnd
rlabel metal2 s 186 33695 294 33771 4 gnd
rlabel metal2 s 186 81885 294 81961 4 gnd
rlabel metal2 s 186 13375 294 13485 4 gnd
rlabel metal2 s 186 16315 294 16391 4 gnd
rlabel metal2 s 186 99739 294 99815 4 gnd
rlabel metal2 s 186 56605 294 56681 4 gnd
rlabel metal2 s 186 60775 294 60885 4 gnd
rlabel metal2 s 186 89215 294 89325 4 gnd
rlabel metal2 s 186 25795 294 25871 4 gnd
rlabel metal2 s 186 35749 294 35825 4 gnd
rlabel metal2 s 186 40489 294 40565 4 gnd
rlabel metal2 s 186 16789 294 16865 4 gnd
rlabel metal2 s 186 93735 294 93811 4 gnd
rlabel metal2 s 186 31325 294 31401 4 gnd
rlabel metal2 s 186 70509 294 70585 4 gnd
rlabel metal2 s 186 59985 294 60095 4 gnd
rlabel metal2 s 186 95315 294 95391 4 gnd
rlabel metal2 s 186 5255 294 5331 4 gnd
rlabel metal2 s 186 41815 294 41925 4 gnd
rlabel metal2 s 186 53919 294 53995 4 gnd
rlabel metal2 s 186 54455 294 54565 4 gnd
rlabel metal2 s 186 28385 294 28495 4 gnd
rlabel metal2 s 186 22855 294 22965 4 gnd
rlabel metal2 s 186 13629 294 13705 4 gnd
rlabel metal2 s 186 22635 294 22711 4 gnd
rlabel metal2 s 186 91585 294 91695 4 gnd
rlabel metal2 s 186 64725 294 64835 4 gnd
rlabel metal2 s 186 59449 294 59525 4 gnd
rlabel metal2 s 186 96105 294 96181 4 gnd
rlabel metal2 s 186 50505 294 50615 4 gnd
rlabel metal2 s 186 72405 294 72481 4 gnd
rlabel metal2 s 186 76829 294 76905 4 gnd
rlabel metal2 s 186 93165 294 93275 4 gnd
rlabel metal2 s 186 46809 294 46885 4 gnd
rlabel metal2 s 186 100055 294 100131 4 gnd
rlabel metal2 s 186 89785 294 89861 4 gnd
rlabel metal2 s 186 77619 294 77695 4 gnd
rlabel metal2 s 186 23645 294 23755 4 gnd
rlabel metal2 s 186 70825 294 70901 4 gnd
rlabel metal2 s 186 79989 294 80065 4 gnd
rlabel metal2 s 186 43965 294 44041 4 gnd
rlabel metal2 s 186 27375 294 27451 4 gnd
rlabel metal2 s 186 31009 294 31085 4 gnd
rlabel metal2 s 186 21055 294 21131 4 gnd
rlabel metal2 s 186 24435 294 24545 4 gnd
rlabel metal2 s 186 54235 294 54311 4 gnd
rlabel metal2 s 186 40015 294 40091 4 gnd
rlabel metal2 s 186 63935 294 64045 4 gnd
rlabel metal2 s 186 26269 294 26345 4 gnd
rlabel metal2 s 186 48705 294 48781 4 gnd
rlabel metal2 s 186 36065 294 36141 4 gnd
rlabel metal2 s 186 90259 294 90335 4 gnd
rlabel metal2 s 186 94745 294 94855 4 gnd
rlabel metal2 s 186 54709 294 54785 4 gnd
rlabel metal2 s 186 25479 294 25555 4 gnd
rlabel metal2 s 186 74459 294 74535 4 gnd
rlabel metal2 s 186 42385 294 42461 4 gnd
rlabel metal2 s 186 42859 294 42935 4 gnd
rlabel metal2 s 186 28165 294 28241 4 gnd
rlabel metal2 s 186 65515 294 65625 4 gnd
rlabel metal2 s 186 18685 294 18761 4 gnd
rlabel metal2 s 186 101635 294 101711 4 gnd
rlabel metal2 s 186 63399 294 63475 4 gnd
rlabel metal2 s 186 97369 294 97445 4 gnd
rlabel metal2 s 186 38435 294 38511 4 gnd
rlabel metal2 s 186 57869 294 57945 4 gnd
rlabel metal2 s 186 58185 294 58261 4 gnd
rlabel metal2 s 186 14955 294 15065 4 gnd
rlabel metal2 s 186 37329 294 37405 4 gnd
rlabel metal2 s 186 59195 294 59305 4 gnd
rlabel metal2 s 186 66305 294 66415 4 gnd
rlabel metal2 s 186 8889 294 8965 4 gnd
rlabel metal2 s 186 84729 294 84805 4 gnd
rlabel metal2 s 186 95535 294 95645 4 gnd
rlabel metal2 s 186 38909 294 38985 4 gnd
rlabel metal2 s 186 8415 294 8491 4 gnd
rlabel metal2 s 186 26585 294 26661 4 gnd
rlabel metal2 s 186 82359 294 82435 4 gnd
rlabel metal2 s 186 52339 294 52415 4 gnd
rlabel metal2 s 186 11259 294 11335 4 gnd
rlabel metal2 s 186 100275 294 100385 4 gnd
rlabel metal2 s 186 97115 294 97225 4 gnd
rlabel metal2 s 186 4939 294 5015 4 gnd
rlabel metal2 s 186 67885 294 67995 4 gnd
rlabel metal2 s 186 17895 294 17971 4 gnd
rlabel metal2 s 186 34485 294 34561 4 gnd
rlabel metal2 s 186 68139 294 68215 4 gnd
rlabel metal2 s 186 24689 294 24765 4 gnd
rlabel metal2 s 186 51865 294 51941 4 gnd
rlabel metal2 s 186 98159 294 98235 4 gnd
rlabel metal2 s 186 34705 294 34815 4 gnd
rlabel metal2 s 186 90795 294 90905 4 gnd
rlabel metal2 s 186 78155 294 78265 4 gnd
rlabel metal2 s 186 83939 294 84015 4 gnd
rlabel metal2 s 186 58405 294 58515 4 gnd
rlabel metal2 s 186 46019 294 46095 4 gnd
rlabel metal2 s 186 15209 294 15285 4 gnd
rlabel metal2 s 186 68455 294 68531 4 gnd
rlabel metal2 s 186 33125 294 33235 4 gnd
rlabel metal2 s 186 9679 294 9755 4 gnd
rlabel metal2 s 186 38655 294 38765 4 gnd
rlabel metal2 s 186 71835 294 71945 4 gnd
rlabel metal2 s 186 62925 294 63001 4 gnd
rlabel metal2 s 186 73415 294 73525 4 gnd
rlabel metal2 s 186 22319 294 22395 4 gnd
rlabel metal2 s 186 49715 294 49825 4 gnd
rlabel metal2 s 186 87099 294 87175 4 gnd
rlabel metal2 s 186 85835 294 85911 4 gnd
rlabel metal2 s 186 72089 294 72165 4 gnd
rlabel metal2 s 186 7625 294 7701 4 gnd
rlabel metal2 s 186 10469 294 10545 4 gnd
rlabel metal2 s 186 8635 294 8745 4 gnd
rlabel metal2 s 186 48925 294 49035 4 gnd
rlabel metal2 s 186 49179 294 49255 4 gnd
rlabel metal2 s 186 51075 294 51151 4 gnd
rlabel metal2 s 186 9425 294 9535 4 gnd
rlabel metal2 s 186 73669 294 73745 4 gnd
rlabel metal2 s 186 19475 294 19551 4 gnd
rlabel metal2 s 186 70035 294 70111 4 gnd
rlabel metal2 s 186 71615 294 71691 4 gnd
rlabel metal2 s 186 30219 294 30295 4 gnd
rlabel metal2 s 186 10785 294 10861 4 gnd
rlabel metal2 s 186 28955 294 29031 4 gnd
rlabel metal2 s 186 62355 294 62465 4 gnd
rlabel metal2 s 186 1525 294 1635 4 gnd
rlabel metal2 s 186 5729 294 5805 4 gnd
rlabel metal2 s 186 3105 294 3215 4 gnd
rlabel metal2 s 186 12049 294 12125 4 gnd
rlabel metal2 s 186 38119 294 38195 4 gnd
rlabel metal2 s 186 29965 294 30075 4 gnd
rlabel metal2 s 186 93419 294 93495 4 gnd
rlabel metal2 s 186 63145 294 63255 4 gnd
rlabel metal2 s 186 7055 294 7165 4 gnd
rlabel metal2 s 186 90005 294 90115 4 gnd
rlabel metal2 s 186 58975 294 59051 4 gnd
rlabel metal2 s 186 45229 294 45305 4 gnd
rlabel metal2 s 186 31799 294 31875 4 gnd
rlabel metal2 s 186 92375 294 92485 4 gnd
rlabel metal2 s 186 30535 294 30611 4 gnd
rlabel metal2 s 186 15999 294 16075 4 gnd
rlabel metal2 s 186 88425 294 88535 4 gnd
rlabel metal2 s 186 7845 294 7955 4 gnd
rlabel metal2 s 186 85519 294 85595 4 gnd
rlabel metal2 s 186 96325 294 96435 4 gnd
rlabel metal2 s 186 18115 294 18225 4 gnd
rlabel metal2 s 186 26015 294 26125 4 gnd
rlabel metal2 s 186 69465 294 69575 4 gnd
rlabel metal2 s 186 32335 294 32445 4 gnd
rlabel metal2 s 186 102109 294 102185 4 gnd
rlabel metal2 s 186 77365 294 77475 4 gnd
rlabel metal2 s 186 52875 294 52985 4 gnd
rlabel metal2 s 186 20485 294 20595 4 gnd
rlabel metal2 s 186 98949 294 99025 4 gnd
rlabel metal2 s 186 22065 294 22175 4 gnd
rlabel metal2 s 186 17325 294 17435 4 gnd
rlabel metal2 s 186 78725 294 78801 4 gnd
rlabel metal2 s 186 42605 294 42715 4 gnd
rlabel metal2 s 186 73985 294 74061 4 gnd
rlabel metal2 s 186 29429 294 29505 4 gnd
rlabel metal2 s 186 23899 294 23975 4 gnd
rlabel metal2 s 186 37865 294 37975 4 gnd
rlabel metal2 s 186 56825 294 56935 4 gnd
rlabel metal2 s 186 98695 294 98805 4 gnd
rlabel metal2 s 186 100529 294 100605 4 gnd
rlabel metal2 s 186 30755 294 30865 4 gnd
rlabel metal2 s 186 97685 294 97761 4 gnd
rlabel metal2 s 186 80305 294 80381 4 gnd
rlabel metal2 s 186 72879 294 72955 4 gnd
rlabel metal2 s 186 68675 294 68785 4 gnd
rlabel metal2 s 186 94525 294 94601 4 gnd
rlabel metal2 s 186 6519 294 6595 4 gnd
rlabel metal2 s 186 23109 294 23185 4 gnd
rlabel metal2 s 186 33915 294 34025 4 gnd
rlabel metal2 s 186 64505 294 64581 4 gnd
rlabel metal2 s 186 34959 294 35035 4 gnd
rlabel metal2 s 186 80779 294 80855 4 gnd
rlabel metal2 s 186 77935 294 78011 4 gnd
rlabel metal2 s 186 92629 294 92705 4 gnd
rlabel metal2 s 186 66875 294 66951 4 gnd
rlabel metal2 s 186 40805 294 40881 4 gnd
rlabel metal2 s 186 44755 294 44831 4 gnd
rlabel metal2 s 186 79735 294 79845 4 gnd
rlabel metal2 s 186 83465 294 83541 4 gnd
rlabel metal2 s 186 14735 294 14811 4 gnd
rlabel metal2 s 186 3359 294 3435 4 gnd
rlabel metal2 s 186 2315 294 2425 4 gnd
rlabel metal2 s 186 66085 294 66161 4 gnd
rlabel metal2 s 186 81569 294 81645 4 gnd
rlabel metal2 s 186 17579 294 17655 4 gnd
rlabel metal2 s 186 55025 294 55101 4 gnd
rlabel metal2 s 186 82675 294 82751 4 gnd
rlabel metal2 s 186 76575 294 76685 4 gnd
rlabel metal2 s 186 20265 294 20341 4 gnd
rlabel metal2 s 186 53129 294 53205 4 gnd
rlabel metal2 s 186 41279 294 41355 4 gnd
rlabel metal2 s 186 44185 294 44295 4 gnd
rlabel metal2 s 186 46555 294 46665 4 gnd
rlabel metal2 s 186 55245 294 55355 4 gnd
rlabel metal2 s 186 18905 294 19015 4 gnd
rlabel metal2 s 186 43649 294 43725 4 gnd
rlabel metal2 s 186 61345 294 61421 4 gnd
rlabel metal2 s 186 51295 294 51405 4 gnd
rlabel metal2 s 186 82895 294 83005 4 gnd
rlabel metal2 s 186 36855 294 36931 4 gnd
rlabel metal2 s 186 96579 294 96655 4 gnd
rlabel metal2 s 186 21845 294 21921 4 gnd
rlabel metal2 s 186 69719 294 69795 4 gnd
rlabel metal2 s 186 60555 294 60631 4 gnd
rlabel metal2 s 186 32115 294 32191 4 gnd
rlabel metal2 s 186 85045 294 85121 4 gnd
rlabel metal2 s 186 95789 294 95865 4 gnd
rlabel metal2 s 186 50285 294 50361 4 gnd
rlabel metal2 s 186 47125 294 47201 4 gnd
rlabel metal2 s 186 41595 294 41671 4 gnd
rlabel metal2 s 186 11795 294 11905 4 gnd
rlabel metal2 s 186 101319 294 101395 4 gnd
<< properties >>
string FIXED_BBOX 0 0 624 102700
<< end >>
