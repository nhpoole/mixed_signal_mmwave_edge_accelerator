magic
tech sky130A
magscale 1 2
timestamp 1626065694
<< checkpaint >>
rect -2191 -1560 2191 1560
<< pwell >>
rect -931 -300 931 300
<< nmos >>
rect -745 -100 -545 100
rect -487 -100 -287 100
rect -229 -100 -29 100
rect 29 -100 229 100
rect 287 -100 487 100
rect 545 -100 745 100
<< ndiff >>
rect -803 85 -745 100
rect -803 51 -791 85
rect -757 51 -745 85
rect -803 17 -745 51
rect -803 -17 -791 17
rect -757 -17 -745 17
rect -803 -51 -745 -17
rect -803 -85 -791 -51
rect -757 -85 -745 -51
rect -803 -100 -745 -85
rect -545 85 -487 100
rect -545 51 -533 85
rect -499 51 -487 85
rect -545 17 -487 51
rect -545 -17 -533 17
rect -499 -17 -487 17
rect -545 -51 -487 -17
rect -545 -85 -533 -51
rect -499 -85 -487 -51
rect -545 -100 -487 -85
rect -287 85 -229 100
rect -287 51 -275 85
rect -241 51 -229 85
rect -287 17 -229 51
rect -287 -17 -275 17
rect -241 -17 -229 17
rect -287 -51 -229 -17
rect -287 -85 -275 -51
rect -241 -85 -229 -51
rect -287 -100 -229 -85
rect -29 85 29 100
rect -29 51 -17 85
rect 17 51 29 85
rect -29 17 29 51
rect -29 -17 -17 17
rect 17 -17 29 17
rect -29 -51 29 -17
rect -29 -85 -17 -51
rect 17 -85 29 -51
rect -29 -100 29 -85
rect 229 85 287 100
rect 229 51 241 85
rect 275 51 287 85
rect 229 17 287 51
rect 229 -17 241 17
rect 275 -17 287 17
rect 229 -51 287 -17
rect 229 -85 241 -51
rect 275 -85 287 -51
rect 229 -100 287 -85
rect 487 85 545 100
rect 487 51 499 85
rect 533 51 545 85
rect 487 17 545 51
rect 487 -17 499 17
rect 533 -17 545 17
rect 487 -51 545 -17
rect 487 -85 499 -51
rect 533 -85 545 -51
rect 487 -100 545 -85
rect 745 85 803 100
rect 745 51 757 85
rect 791 51 803 85
rect 745 17 803 51
rect 745 -17 757 17
rect 791 -17 803 17
rect 745 -51 803 -17
rect 745 -85 757 -51
rect 791 -85 803 -51
rect 745 -100 803 -85
<< ndiffc >>
rect -791 51 -757 85
rect -791 -17 -757 17
rect -791 -85 -757 -51
rect -533 51 -499 85
rect -533 -17 -499 17
rect -533 -85 -499 -51
rect -275 51 -241 85
rect -275 -17 -241 17
rect -275 -85 -241 -51
rect -17 51 17 85
rect -17 -17 17 17
rect -17 -85 17 -51
rect 241 51 275 85
rect 241 -17 275 17
rect 241 -85 275 -51
rect 499 51 533 85
rect 499 -17 533 17
rect 499 -85 533 -51
rect 757 51 791 85
rect 757 -17 791 17
rect 757 -85 791 -51
<< psubdiff >>
rect -905 240 -799 274
rect -765 240 -731 274
rect -697 240 -663 274
rect -629 240 -595 274
rect -561 240 -527 274
rect -493 240 -459 274
rect -425 240 -391 274
rect -357 240 -323 274
rect -289 240 -255 274
rect -221 240 -187 274
rect -153 240 -119 274
rect -85 240 -51 274
rect -17 240 17 274
rect 51 240 85 274
rect 119 240 153 274
rect 187 240 221 274
rect 255 240 289 274
rect 323 240 357 274
rect 391 240 425 274
rect 459 240 493 274
rect 527 240 561 274
rect 595 240 629 274
rect 663 240 697 274
rect 731 240 765 274
rect 799 240 905 274
rect -905 153 -871 240
rect -905 85 -871 119
rect 871 153 905 240
rect -905 17 -871 51
rect -905 -51 -871 -17
rect -905 -119 -871 -85
rect 871 85 905 119
rect 871 17 905 51
rect 871 -51 905 -17
rect -905 -240 -871 -153
rect 871 -119 905 -85
rect 871 -240 905 -153
rect -905 -274 -799 -240
rect -765 -274 -731 -240
rect -697 -274 -663 -240
rect -629 -274 -595 -240
rect -561 -274 -527 -240
rect -493 -274 -459 -240
rect -425 -274 -391 -240
rect -357 -274 -323 -240
rect -289 -274 -255 -240
rect -221 -274 -187 -240
rect -153 -274 -119 -240
rect -85 -274 -51 -240
rect -17 -274 17 -240
rect 51 -274 85 -240
rect 119 -274 153 -240
rect 187 -274 221 -240
rect 255 -274 289 -240
rect 323 -274 357 -240
rect 391 -274 425 -240
rect 459 -274 493 -240
rect 527 -274 561 -240
rect 595 -274 629 -240
rect 663 -274 697 -240
rect 731 -274 765 -240
rect 799 -274 905 -240
<< psubdiffcont >>
rect -799 240 -765 274
rect -731 240 -697 274
rect -663 240 -629 274
rect -595 240 -561 274
rect -527 240 -493 274
rect -459 240 -425 274
rect -391 240 -357 274
rect -323 240 -289 274
rect -255 240 -221 274
rect -187 240 -153 274
rect -119 240 -85 274
rect -51 240 -17 274
rect 17 240 51 274
rect 85 240 119 274
rect 153 240 187 274
rect 221 240 255 274
rect 289 240 323 274
rect 357 240 391 274
rect 425 240 459 274
rect 493 240 527 274
rect 561 240 595 274
rect 629 240 663 274
rect 697 240 731 274
rect 765 240 799 274
rect -905 119 -871 153
rect 871 119 905 153
rect -905 51 -871 85
rect -905 -17 -871 17
rect -905 -85 -871 -51
rect 871 51 905 85
rect 871 -17 905 17
rect 871 -85 905 -51
rect -905 -153 -871 -119
rect 871 -153 905 -119
rect -799 -274 -765 -240
rect -731 -274 -697 -240
rect -663 -274 -629 -240
rect -595 -274 -561 -240
rect -527 -274 -493 -240
rect -459 -274 -425 -240
rect -391 -274 -357 -240
rect -323 -274 -289 -240
rect -255 -274 -221 -240
rect -187 -274 -153 -240
rect -119 -274 -85 -240
rect -51 -274 -17 -240
rect 17 -274 51 -240
rect 85 -274 119 -240
rect 153 -274 187 -240
rect 221 -274 255 -240
rect 289 -274 323 -240
rect 357 -274 391 -240
rect 425 -274 459 -240
rect 493 -274 527 -240
rect 561 -274 595 -240
rect 629 -274 663 -240
rect 697 -274 731 -240
rect 765 -274 799 -240
<< poly >>
rect -711 172 -579 188
rect -711 155 -662 172
rect -745 138 -662 155
rect -628 155 -579 172
rect -453 172 -321 188
rect -453 155 -404 172
rect -628 138 -545 155
rect -745 100 -545 138
rect -487 138 -404 155
rect -370 155 -321 172
rect -195 172 -63 188
rect -195 155 -146 172
rect -370 138 -287 155
rect -487 100 -287 138
rect -229 138 -146 155
rect -112 155 -63 172
rect 63 172 195 188
rect 63 155 112 172
rect -112 138 -29 155
rect -229 100 -29 138
rect 29 138 112 155
rect 146 155 195 172
rect 321 172 453 188
rect 321 155 370 172
rect 146 138 229 155
rect 29 100 229 138
rect 287 138 370 155
rect 404 155 453 172
rect 579 172 711 188
rect 579 155 628 172
rect 404 138 487 155
rect 287 100 487 138
rect 545 138 628 155
rect 662 155 711 172
rect 662 138 745 155
rect 545 100 745 138
rect -745 -138 -545 -100
rect -745 -155 -662 -138
rect -711 -172 -662 -155
rect -628 -155 -545 -138
rect -487 -138 -287 -100
rect -487 -155 -404 -138
rect -628 -172 -579 -155
rect -711 -188 -579 -172
rect -453 -172 -404 -155
rect -370 -155 -287 -138
rect -229 -138 -29 -100
rect -229 -155 -146 -138
rect -370 -172 -321 -155
rect -453 -188 -321 -172
rect -195 -172 -146 -155
rect -112 -155 -29 -138
rect 29 -138 229 -100
rect 29 -155 112 -138
rect -112 -172 -63 -155
rect -195 -188 -63 -172
rect 63 -172 112 -155
rect 146 -155 229 -138
rect 287 -138 487 -100
rect 287 -155 370 -138
rect 146 -172 195 -155
rect 63 -188 195 -172
rect 321 -172 370 -155
rect 404 -155 487 -138
rect 545 -138 745 -100
rect 545 -155 628 -138
rect 404 -172 453 -155
rect 321 -188 453 -172
rect 579 -172 628 -155
rect 662 -155 745 -138
rect 662 -172 711 -155
rect 579 -188 711 -172
<< polycont >>
rect -662 138 -628 172
rect -404 138 -370 172
rect -146 138 -112 172
rect 112 138 146 172
rect 370 138 404 172
rect 628 138 662 172
rect -662 -172 -628 -138
rect -404 -172 -370 -138
rect -146 -172 -112 -138
rect 112 -172 146 -138
rect 370 -172 404 -138
rect 628 -172 662 -138
<< locali >>
rect -905 240 -799 274
rect -765 240 -731 274
rect -697 240 -663 274
rect -629 240 -595 274
rect -561 240 -527 274
rect -493 240 -459 274
rect -425 240 -391 274
rect -357 240 -323 274
rect -289 240 -255 274
rect -221 240 -187 274
rect -153 240 -119 274
rect -85 240 -51 274
rect -17 240 17 274
rect 51 240 85 274
rect 119 240 153 274
rect 187 240 221 274
rect 255 240 289 274
rect 323 240 357 274
rect 391 240 425 274
rect 459 240 493 274
rect 527 240 561 274
rect 595 240 629 274
rect 663 240 697 274
rect 731 240 765 274
rect 799 240 905 274
rect -905 153 -871 240
rect -711 138 -662 172
rect -628 138 -579 172
rect -453 138 -404 172
rect -370 138 -321 172
rect -195 138 -146 172
rect -112 138 -63 172
rect 63 138 112 172
rect 146 138 195 172
rect 321 138 370 172
rect 404 138 453 172
rect 579 138 628 172
rect 662 138 711 172
rect 871 153 905 240
rect -905 85 -871 119
rect -905 17 -871 51
rect -905 -51 -871 -17
rect -905 -119 -871 -85
rect -791 85 -757 104
rect -791 17 -757 19
rect -791 -19 -757 -17
rect -791 -104 -757 -85
rect -533 85 -499 104
rect -533 17 -499 19
rect -533 -19 -499 -17
rect -533 -104 -499 -85
rect -275 85 -241 104
rect -275 17 -241 19
rect -275 -19 -241 -17
rect -275 -104 -241 -85
rect -17 85 17 104
rect -17 17 17 19
rect -17 -19 17 -17
rect -17 -104 17 -85
rect 241 85 275 104
rect 241 17 275 19
rect 241 -19 275 -17
rect 241 -104 275 -85
rect 499 85 533 104
rect 499 17 533 19
rect 499 -19 533 -17
rect 499 -104 533 -85
rect 757 85 791 104
rect 757 17 791 19
rect 757 -19 791 -17
rect 757 -104 791 -85
rect 871 85 905 119
rect 871 17 905 51
rect 871 -51 905 -17
rect 871 -119 905 -85
rect -905 -240 -871 -153
rect -711 -172 -662 -138
rect -628 -172 -579 -138
rect -453 -172 -404 -138
rect -370 -172 -321 -138
rect -195 -172 -146 -138
rect -112 -172 -63 -138
rect 63 -172 112 -138
rect 146 -172 195 -138
rect 321 -172 370 -138
rect 404 -172 453 -138
rect 579 -172 628 -138
rect 662 -172 711 -138
rect 871 -240 905 -153
rect -905 -274 -799 -240
rect -765 -274 -731 -240
rect -697 -274 -663 -240
rect -629 -274 -595 -240
rect -561 -274 -527 -240
rect -493 -274 -459 -240
rect -425 -274 -391 -240
rect -357 -274 -323 -240
rect -289 -274 -255 -240
rect -221 -274 -187 -240
rect -153 -274 -119 -240
rect -85 -274 -51 -240
rect -17 -274 17 -240
rect 51 -274 85 -240
rect 119 -274 153 -240
rect 187 -274 221 -240
rect 255 -274 289 -240
rect 323 -274 357 -240
rect 391 -274 425 -240
rect 459 -274 493 -240
rect 527 -274 561 -240
rect 595 -274 629 -240
rect 663 -274 697 -240
rect 731 -274 765 -240
rect 799 -274 905 -240
<< viali >>
rect -662 138 -628 172
rect -404 138 -370 172
rect -146 138 -112 172
rect 112 138 146 172
rect 370 138 404 172
rect 628 138 662 172
rect -791 51 -757 53
rect -791 19 -757 51
rect -791 -51 -757 -19
rect -791 -53 -757 -51
rect -533 51 -499 53
rect -533 19 -499 51
rect -533 -51 -499 -19
rect -533 -53 -499 -51
rect -275 51 -241 53
rect -275 19 -241 51
rect -275 -51 -241 -19
rect -275 -53 -241 -51
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect 241 51 275 53
rect 241 19 275 51
rect 241 -51 275 -19
rect 241 -53 275 -51
rect 499 51 533 53
rect 499 19 533 51
rect 499 -51 533 -19
rect 499 -53 533 -51
rect 757 51 791 53
rect 757 19 791 51
rect 757 -51 791 -19
rect 757 -53 791 -51
rect -662 -172 -628 -138
rect -404 -172 -370 -138
rect -146 -172 -112 -138
rect 112 -172 146 -138
rect 370 -172 404 -138
rect 628 -172 662 -138
<< metal1 >>
rect -699 172 -591 178
rect -699 138 -662 172
rect -628 138 -591 172
rect -699 132 -591 138
rect -441 172 -333 178
rect -441 138 -404 172
rect -370 138 -333 172
rect -441 132 -333 138
rect -183 172 -75 178
rect -183 138 -146 172
rect -112 138 -75 172
rect -183 132 -75 138
rect 75 172 183 178
rect 75 138 112 172
rect 146 138 183 172
rect 75 132 183 138
rect 333 172 441 178
rect 333 138 370 172
rect 404 138 441 172
rect 333 132 441 138
rect 591 172 699 178
rect 591 138 628 172
rect 662 138 699 172
rect 591 132 699 138
rect -797 53 -751 100
rect -797 19 -791 53
rect -757 19 -751 53
rect -797 -19 -751 19
rect -797 -53 -791 -19
rect -757 -53 -751 -19
rect -797 -100 -751 -53
rect -539 53 -493 100
rect -539 19 -533 53
rect -499 19 -493 53
rect -539 -19 -493 19
rect -539 -53 -533 -19
rect -499 -53 -493 -19
rect -539 -100 -493 -53
rect -281 53 -235 100
rect -281 19 -275 53
rect -241 19 -235 53
rect -281 -19 -235 19
rect -281 -53 -275 -19
rect -241 -53 -235 -19
rect -281 -100 -235 -53
rect -23 53 23 100
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -100 23 -53
rect 235 53 281 100
rect 235 19 241 53
rect 275 19 281 53
rect 235 -19 281 19
rect 235 -53 241 -19
rect 275 -53 281 -19
rect 235 -100 281 -53
rect 493 53 539 100
rect 493 19 499 53
rect 533 19 539 53
rect 493 -19 539 19
rect 493 -53 499 -19
rect 533 -53 539 -19
rect 493 -100 539 -53
rect 751 53 797 100
rect 751 19 757 53
rect 791 19 797 53
rect 751 -19 797 19
rect 751 -53 757 -19
rect 791 -53 797 -19
rect 751 -100 797 -53
rect -699 -138 -591 -132
rect -699 -172 -662 -138
rect -628 -172 -591 -138
rect -699 -178 -591 -172
rect -441 -138 -333 -132
rect -441 -172 -404 -138
rect -370 -172 -333 -138
rect -441 -178 -333 -172
rect -183 -138 -75 -132
rect -183 -172 -146 -138
rect -112 -172 -75 -138
rect -183 -178 -75 -172
rect 75 -138 183 -132
rect 75 -172 112 -138
rect 146 -172 183 -138
rect 75 -178 183 -172
rect 333 -138 441 -132
rect 333 -172 370 -138
rect 404 -172 441 -138
rect 333 -178 441 -172
rect 591 -138 699 -132
rect 591 -172 628 -138
rect 662 -172 699 -138
rect 591 -178 699 -172
<< properties >>
string FIXED_BBOX -888 -257 888 257
<< end >>
