magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect -1444 -1548 1444 1548
<< pwell >>
rect -184 -226 184 226
<< nmos >>
rect -100 -200 100 200
<< ndiff >>
rect -158 187 -100 200
rect -158 153 -146 187
rect -112 153 -100 187
rect -158 119 -100 153
rect -158 85 -146 119
rect -112 85 -100 119
rect -158 51 -100 85
rect -158 17 -146 51
rect -112 17 -100 51
rect -158 -17 -100 17
rect -158 -51 -146 -17
rect -112 -51 -100 -17
rect -158 -85 -100 -51
rect -158 -119 -146 -85
rect -112 -119 -100 -85
rect -158 -153 -100 -119
rect -158 -187 -146 -153
rect -112 -187 -100 -153
rect -158 -200 -100 -187
rect 100 187 158 200
rect 100 153 112 187
rect 146 153 158 187
rect 100 119 158 153
rect 100 85 112 119
rect 146 85 158 119
rect 100 51 158 85
rect 100 17 112 51
rect 146 17 158 51
rect 100 -17 158 17
rect 100 -51 112 -17
rect 146 -51 158 -17
rect 100 -85 158 -51
rect 100 -119 112 -85
rect 146 -119 158 -85
rect 100 -153 158 -119
rect 100 -187 112 -153
rect 146 -187 158 -153
rect 100 -200 158 -187
<< ndiffc >>
rect -146 153 -112 187
rect -146 85 -112 119
rect -146 17 -112 51
rect -146 -51 -112 -17
rect -146 -119 -112 -85
rect -146 -187 -112 -153
rect 112 153 146 187
rect 112 85 146 119
rect 112 17 146 51
rect 112 -51 146 -17
rect 112 -119 146 -85
rect 112 -187 146 -153
<< poly >>
rect -66 272 66 288
rect -66 255 -17 272
rect -100 238 -17 255
rect 17 255 66 272
rect 17 238 100 255
rect -100 200 100 238
rect -100 -238 100 -200
rect -100 -255 -17 -238
rect -66 -272 -17 -255
rect 17 -255 100 -238
rect 17 -272 66 -255
rect -66 -288 66 -272
<< polycont >>
rect -17 238 17 272
rect -17 -272 17 -238
<< locali >>
rect -66 238 -17 272
rect 17 238 66 272
rect -146 187 -112 204
rect -146 119 -112 127
rect -146 51 -112 55
rect -146 -55 -112 -51
rect -146 -127 -112 -119
rect -146 -204 -112 -187
rect 112 187 146 204
rect 112 119 146 127
rect 112 51 146 55
rect 112 -55 146 -51
rect 112 -127 146 -119
rect 112 -204 146 -187
rect -66 -272 -17 -238
rect 17 -272 66 -238
<< viali >>
rect -17 238 17 272
rect -146 153 -112 161
rect -146 127 -112 153
rect -146 85 -112 89
rect -146 55 -112 85
rect -146 -17 -112 17
rect -146 -85 -112 -55
rect -146 -89 -112 -85
rect -146 -153 -112 -127
rect -146 -161 -112 -153
rect 112 153 146 161
rect 112 127 146 153
rect 112 85 146 89
rect 112 55 146 85
rect 112 -17 146 17
rect 112 -85 146 -55
rect 112 -89 146 -85
rect 112 -153 146 -127
rect 112 -161 146 -153
rect -17 -272 17 -238
<< metal1 >>
rect -54 272 54 278
rect -54 238 -17 272
rect 17 238 54 272
rect -54 232 54 238
rect -152 161 -106 200
rect -152 127 -146 161
rect -112 127 -106 161
rect -152 89 -106 127
rect -152 55 -146 89
rect -112 55 -106 89
rect -152 17 -106 55
rect -152 -17 -146 17
rect -112 -17 -106 17
rect -152 -55 -106 -17
rect -152 -89 -146 -55
rect -112 -89 -106 -55
rect -152 -127 -106 -89
rect -152 -161 -146 -127
rect -112 -161 -106 -127
rect -152 -200 -106 -161
rect 106 161 152 200
rect 106 127 112 161
rect 146 127 152 161
rect 106 89 152 127
rect 106 55 112 89
rect 146 55 152 89
rect 106 17 152 55
rect 106 -17 112 17
rect 146 -17 152 17
rect 106 -55 152 -17
rect 106 -89 112 -55
rect 146 -89 152 -55
rect 106 -127 152 -89
rect 106 -161 112 -127
rect 146 -161 152 -127
rect 106 -200 152 -161
rect -54 -238 54 -232
rect -54 -272 -17 -238
rect 17 -272 54 -238
rect -54 -278 54 -272
<< end >>
