magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect 823 -7639 6557 5632
<< metal1 >>
rect 3283 -5276 5265 -5248
rect 2115 -5378 5141 -5350
<< metal2 >>
rect 2101 -6379 2129 -5364
rect 3269 -6379 3297 -5262
rect 5127 -5364 5155 2850
rect 5251 -5262 5279 4340
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_0
timestamp 1626486988
transform 1 0 3251 0 1 -5294
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_1
timestamp 1626486988
transform 1 0 5233 0 1 4308
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_2
timestamp 1626486988
transform 1 0 5233 0 1 -5294
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_3
timestamp 1626486988
transform 1 0 2083 0 1 -5396
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_4
timestamp 1626486988
transform 1 0 5109 0 1 2818
box 0 0 64 64
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_5
timestamp 1626486988
transform 1 0 5109 0 1 -5396
box 0 0 64 64
<< properties >>
string FIXED_BBOX 2083 -6379 5297 4372
<< end >>
