magic
tech sky130A
magscale 1 2
timestamp 1623661481
<< nwell >>
rect -38 261 1418 582
<< pwell >>
rect 30 -17 64 17
<< locali >>
rect 18 197 66 325
rect 289 191 357 265
rect 1028 334 1096 493
rect 1062 149 1096 334
rect 1028 83 1096 149
rect 1311 301 1363 493
rect 1325 165 1363 301
rect 1311 51 1363 165
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1380 561
rect 35 393 69 493
rect 103 427 169 527
rect 35 359 156 393
rect 122 280 156 359
rect 203 337 248 493
rect 122 214 168 280
rect 122 161 156 214
rect 35 127 156 161
rect 35 69 69 127
rect 103 17 169 93
rect 203 69 237 337
rect 296 333 362 483
rect 396 367 459 527
rect 584 426 722 455
rect 756 435 790 527
rect 584 423 723 426
rect 584 421 724 423
rect 672 418 725 421
rect 672 415 726 418
rect 675 412 726 415
rect 684 406 726 412
rect 686 403 726 406
rect 296 299 433 333
rect 399 247 433 299
rect 499 271 556 401
rect 590 283 658 382
rect 399 181 473 247
rect 590 207 624 283
rect 692 265 726 403
rect 860 373 910 487
rect 760 324 910 373
rect 944 366 994 527
rect 760 307 916 324
rect 879 265 916 307
rect 692 233 845 265
rect 399 157 433 181
rect 307 123 433 157
rect 513 141 624 207
rect 671 199 845 233
rect 879 199 1028 265
rect 307 69 341 123
rect 671 107 705 199
rect 879 168 916 199
rect 860 132 916 168
rect 375 17 446 89
rect 558 73 705 107
rect 753 17 819 122
rect 860 83 894 132
rect 928 17 994 99
rect 1132 265 1182 493
rect 1218 367 1277 527
rect 1132 199 1291 265
rect 1132 51 1182 199
rect 1218 17 1277 109
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1380 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
<< metal1 >>
rect 0 561 1380 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1380 561
rect 0 496 1380 527
rect 0 17 1380 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1380 17
rect 0 -48 1380 -17
<< obsm1 >>
rect 202 388 260 397
rect 487 388 545 397
rect 202 360 545 388
rect 202 351 260 360
rect 487 351 545 360
rect 110 320 168 329
rect 579 320 637 329
rect 110 292 637 320
rect 110 283 168 292
rect 579 283 637 292
<< labels >>
rlabel locali s 289 191 357 265 6 D
port 1 nsew signal input
rlabel locali s 1062 149 1096 334 6 Q
port 2 nsew signal output
rlabel locali s 1028 334 1096 493 6 Q
port 2 nsew signal output
rlabel locali s 1028 83 1096 149 6 Q
port 2 nsew signal output
rlabel locali s 1325 165 1363 301 6 Q_N
port 3 nsew signal output
rlabel locali s 1311 301 1363 493 6 Q_N
port 3 nsew signal output
rlabel locali s 1311 51 1363 165 6 Q_N
port 3 nsew signal output
rlabel locali s 18 197 66 325 6 GATE_N
port 4 nsew clock input
rlabel metal1 s 0 -48 1380 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 17 8 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 1418 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 1380 592 6 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1380 544
string LEFsymmetry X Y R90
string LEFview TRUE
<< end >>
