magic
tech sky130A
magscale 1 2
timestamp 1623661481
<< nwell >>
rect -38 261 498 582
<< pwell >>
rect 30 -17 64 17
<< locali >>
rect 324 425 443 493
rect 17 199 109 345
rect 324 161 359 425
rect 395 195 443 391
rect 324 51 443 161
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 17 413 69 493
rect 103 447 290 527
rect 17 379 290 413
rect 143 165 290 379
rect 17 131 290 165
rect 17 51 69 131
rect 103 17 290 97
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
<< metal1 >>
rect 0 561 460 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 496 460 527
rect 0 17 460 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
rect 0 -48 460 -17
<< labels >>
rlabel locali s 395 195 443 391 6 A
port 1 nsew signal input
rlabel locali s 17 199 109 345 6 TE
port 2 nsew signal input
rlabel locali s 324 425 443 493 6 Z
port 3 nsew signal output
rlabel locali s 324 161 359 425 6 Z
port 3 nsew signal output
rlabel locali s 324 51 443 161 6 Z
port 3 nsew signal output
rlabel metal1 s 0 -48 460 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 17 8 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 498 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 460 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 460 544
string LEFsymmetry X Y R90
string LEFview TRUE
<< end >>
