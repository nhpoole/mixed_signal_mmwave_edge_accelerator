magic
tech sky130A
magscale 1 2
timestamp 1623661481
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 29 -17 63 17
<< locali >>
rect 226 333 292 493
rect 417 333 483 493
rect 226 299 627 333
rect 85 199 155 265
rect 193 199 247 265
rect 301 153 351 265
rect 385 153 437 265
rect 585 165 627 299
rect 539 51 627 165
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 17 319 102 385
rect 17 165 51 319
rect 142 299 192 527
rect 326 367 383 527
rect 541 367 584 527
rect 17 131 267 165
rect 471 199 551 265
rect 17 89 95 131
rect 231 119 267 131
rect 471 119 505 199
rect 131 17 197 97
rect 231 85 505 119
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
rlabel locali s 85 199 155 265 6 A_N
port 1 nsew signal input
rlabel locali s 385 153 437 265 6 B
port 2 nsew signal input
rlabel locali s 301 153 351 265 6 C
port 3 nsew signal input
rlabel locali s 193 199 247 265 6 D
port 4 nsew signal input
rlabel locali s 585 165 627 299 6 Y
port 5 nsew signal output
rlabel locali s 539 51 627 165 6 Y
port 5 nsew signal output
rlabel locali s 417 333 483 493 6 Y
port 5 nsew signal output
rlabel locali s 226 333 292 493 6 Y
port 5 nsew signal output
rlabel locali s 226 299 627 333 6 Y
port 5 nsew signal output
rlabel metal1 s 0 -48 644 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 17 8 VNB
port 7 nsew ground bidirectional
rlabel nwell s -38 261 682 582 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 496 644 592 6 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 644 544
string LEFsymmetry X Y R90
string LEFview TRUE
<< end >>
