magic
tech sky130A
magscale 1 2
timestamp 1624007260
<< error_p >>
rect 9965 14229 9999 14263
rect 8677 14161 8711 14195
rect 10149 14161 10183 14195
rect 10241 14161 10275 14195
rect 8769 14025 8803 14059
rect 9321 13957 9355 13991
rect 9965 13957 9999 13991
rect 8585 13753 8619 13787
rect 10149 13753 10183 13787
rect 8769 13549 8803 13583
rect 8493 13481 8527 13515
rect 9030 13481 9064 13515
rect 9229 13209 9263 13243
rect 8769 13141 8803 13175
rect 9030 13073 9064 13107
rect 9137 13073 9171 13107
rect 9781 13073 9815 13107
rect 9965 13073 9999 13107
rect 8585 13005 8619 13039
rect 9413 13005 9447 13039
rect 9597 12937 9631 12971
rect 9781 12937 9815 12971
rect 8769 12461 8803 12495
rect 9030 12393 9064 12427
rect 9781 12121 9815 12155
rect 8478 12053 8512 12087
rect 9965 11985 9999 12019
rect 10149 11849 10183 11883
rect 9597 11781 9631 11815
rect 10057 11577 10091 11611
rect 6193 11373 6227 11407
rect 7849 11373 7883 11407
rect 8125 11373 8159 11407
rect 8493 11373 8527 11407
rect 6377 11305 6411 11339
rect 7582 11296 7616 11330
rect 8309 11305 8343 11339
rect 8749 11296 8783 11339
rect 6469 11237 6503 11271
rect 9873 11237 9907 11271
rect 6837 11033 6871 11067
rect 10149 11033 10183 11067
rect 6101 10897 6135 10931
rect 6193 10897 6227 10931
rect 6377 10897 6411 10931
rect 6653 10897 6687 10931
rect 8769 10897 8803 10931
rect 9873 10897 9907 10931
rect 6009 10829 6043 10863
rect 6469 10829 6503 10863
rect 10149 10829 10183 10863
rect 7481 10761 7515 10795
rect 8585 10761 8619 10795
rect 6193 10693 6227 10727
rect 9965 10693 9999 10727
rect 10057 10489 10091 10523
rect 6653 10353 6687 10387
rect 6193 10285 6227 10319
rect 6929 10285 6963 10319
rect 8493 10285 8527 10319
rect 7190 10217 7224 10251
rect 8738 10207 8772 10241
rect 6837 10149 6871 10183
rect 8309 10149 8343 10183
rect 9873 10149 9907 10183
rect 9965 10149 9999 10183
rect 7466 9877 7500 9920
rect 10149 9877 10183 9911
rect 6469 9809 6503 9843
rect 6837 9809 6871 9843
rect 7205 9809 7239 9843
rect 9413 9809 9447 9843
rect 9597 9809 9631 9843
rect 9965 9809 9999 9843
rect 6469 9673 6503 9707
rect 7021 9605 7055 9639
rect 9137 9605 9171 9639
rect 9413 9605 9447 9639
rect 9781 9605 9815 9639
rect 6285 9401 6319 9435
rect 6377 9401 6411 9435
rect 8217 9401 8251 9435
rect 7849 9333 7883 9367
rect 8033 9265 8067 9299
rect 6101 9197 6135 9231
rect 7496 9197 7530 9231
rect 7757 9197 7791 9231
rect 8585 9197 8619 9231
rect 8852 9119 8886 9153
rect 6009 8857 6043 8891
rect 10149 8857 10183 8891
rect 7926 8789 7960 8823
rect 6101 8721 6135 8755
rect 6469 8721 6503 8755
rect 7665 8721 7699 8755
rect 9413 8721 9447 8755
rect 9965 8721 9999 8755
rect 6745 8653 6779 8687
rect 7389 8653 7423 8687
rect 9781 8653 9815 8687
rect 7573 8585 7607 8619
rect 9597 8585 9631 8619
rect 7205 8517 7239 8551
rect 9045 8517 9079 8551
rect 7389 8313 7423 8347
rect 9965 8313 9999 8347
rect 7297 8177 7331 8211
rect 7036 8109 7070 8143
rect 7573 8109 7607 8143
rect 7849 8109 7883 8143
rect 8493 8109 8527 8143
rect 7757 8041 7791 8075
rect 8754 8041 8788 8075
rect 7941 7973 7975 8007
rect 9873 7973 9907 8007
rect 5917 7769 5951 7803
rect 6285 7769 6319 7803
rect 7021 7701 7055 7735
rect 7466 7701 7500 7744
rect 9597 7701 9631 7735
rect 6193 7633 6227 7667
rect 6837 7633 6871 7667
rect 7205 7633 7239 7667
rect 9413 7633 9447 7667
rect 9781 7633 9815 7667
rect 9965 7633 9999 7667
rect 6009 7565 6043 7599
rect 8585 7429 8619 7463
rect 9781 7429 9815 7463
rect 6101 7225 6135 7259
rect 8309 7225 8343 7259
rect 6653 7089 6687 7123
rect 9873 7089 9907 7123
rect 6101 7021 6135 7055
rect 6193 7021 6227 7055
rect 6377 7021 6411 7055
rect 6929 7021 6963 7055
rect 6837 6953 6871 6987
rect 7190 6953 7224 6987
rect 9612 6953 9646 6987
rect 6009 6681 6043 6715
rect 7450 6613 7484 6647
rect 6653 6545 6687 6579
rect 9965 6545 9999 6579
rect 9781 6409 9815 6443
rect 6653 6341 6687 6375
rect 8585 6341 8619 6375
rect 8677 6137 8711 6171
rect 9413 6137 9447 6171
rect 9781 6137 9815 6171
rect 6469 6069 6503 6103
rect 6653 6069 6687 6103
rect 7021 6069 7055 6103
rect 8217 6069 8251 6103
rect 6837 5933 6871 5967
rect 7757 5933 7791 5967
rect 8033 5933 8067 5967
rect 8861 5933 8895 5967
rect 9137 5933 9171 5967
rect 9321 5933 9355 5967
rect 9413 5933 9447 5967
rect 9597 5933 9631 5967
rect 9965 5933 9999 5967
rect 10149 5865 10183 5899
rect 6101 5797 6135 5831
rect 6561 5797 6595 5831
<< locali >>
rect 121 14195 155 17901
rect 5457 13855 5491 14297
rect 5641 14195 5675 17085
rect 5641 14161 6026 14195
rect 8878 14161 8987 14195
rect 8953 13991 8987 14161
rect 9137 14161 9246 14195
rect 9137 14059 9171 14161
rect 5365 13821 5491 13855
rect 5365 13243 5399 13821
rect 5273 13209 5399 13243
rect 1409 119 1443 12937
rect 5273 12155 5307 13209
rect 5181 12121 5307 12155
rect 5549 13073 6118 13107
rect 5181 10931 5215 12121
rect 5549 12019 5583 13073
rect 8217 12495 8251 12665
rect 7406 12461 7483 12495
rect 8142 12461 8251 12495
rect 10166 12461 10459 12495
rect 10425 12359 10459 12461
rect 10425 12325 10643 12359
rect 7481 12019 7515 12121
rect 5457 11985 5583 12019
rect 7406 11985 7515 12019
rect 5457 11203 5491 11985
rect 5641 11849 5934 11883
rect 5641 11543 5675 11849
rect 10609 11543 10643 12325
rect 5641 11509 5767 11543
rect 10425 11509 10643 11543
rect 5733 11407 5767 11509
rect 10425 11407 10459 11509
rect 5733 11373 6026 11407
rect 10166 11373 10459 11407
rect 8749 11330 8783 11339
rect 5457 11169 5583 11203
rect 5549 11067 5583 11169
rect 5549 11033 5859 11067
rect 5825 10931 5859 11033
rect 5181 10897 5675 10931
rect 5641 10319 5675 10897
rect 5825 10897 5934 10931
rect 5825 10727 5859 10897
rect 6210 10421 6486 10455
rect 5641 10285 6026 10319
rect 2697 7599 2731 10081
rect 5641 9843 5675 10285
rect 7466 9877 7500 9886
rect 9229 9843 9263 9945
rect 8602 9809 8970 9843
rect 9154 9809 9263 9843
rect 6561 9673 6670 9707
rect 6561 9639 6595 9673
rect 5641 9197 5934 9231
rect 9982 9197 10551 9231
rect 5641 9095 5675 9197
rect 5457 9061 5675 9095
rect 10517 9095 10551 9197
rect 10517 9061 10643 9095
rect 5457 8279 5491 9061
rect 9171 8857 9246 8891
rect 5457 8245 5675 8279
rect 5641 8143 5675 8245
rect 5641 8109 5934 8143
rect 8050 8109 8159 8143
rect 5641 7735 5675 8109
rect 8125 8075 8159 8109
rect 7466 7701 7500 7710
rect 9137 7735 9171 7769
rect 9137 7701 9246 7735
rect 5641 7633 5934 7667
rect 6394 7633 6503 7667
rect 5641 7259 5675 7633
rect 6469 7531 6503 7633
rect 6561 7497 6670 7531
rect 6561 7463 6595 7497
rect 5641 7225 5767 7259
rect 5733 7055 5767 7225
rect 6394 7157 6486 7191
rect 5733 7021 5934 7055
rect 8435 7021 8510 7055
rect 10425 6715 10459 6953
rect 10166 6681 10459 6715
rect 6377 6579 6411 6681
rect 10609 6647 10643 9061
rect 10425 6613 10643 6647
rect 6118 6545 6486 6579
rect 7055 6545 7207 6579
rect 7774 6069 7866 6103
rect 9062 6069 9154 6103
rect 7331 6001 7423 6035
rect 6285 5967 6319 6001
rect 7389 5967 7423 6001
rect 10425 5967 10459 6613
rect 6210 5933 6319 5967
rect 7389 5933 7590 5967
rect 10166 5933 10459 5967
<< viali >>
rect 121 17901 155 17935
rect 5641 17085 5675 17119
rect 121 14161 155 14195
rect 5457 14297 5491 14331
rect 6193 14297 6227 14331
rect 6561 14297 6595 14331
rect 8217 14297 8251 14331
rect 8125 14229 8159 14263
rect 9965 14229 9999 14263
rect 6469 14161 6503 14195
rect 6653 14161 6687 14195
rect 8033 14161 8067 14195
rect 8309 14161 8343 14195
rect 8677 14161 8711 14195
rect 7757 14093 7791 14127
rect 7573 14025 7607 14059
rect 8769 14025 8803 14059
rect 10149 14161 10183 14195
rect 10241 14161 10275 14195
rect 9137 14025 9171 14059
rect 7941 13957 7975 13991
rect 8953 13957 8987 13991
rect 9321 13957 9355 13991
rect 9965 13957 9999 13991
rect 6745 13753 6779 13787
rect 8585 13753 8619 13787
rect 10149 13753 10183 13787
rect 6929 13685 6963 13719
rect 8048 13549 8082 13583
rect 8309 13549 8343 13583
rect 8769 13549 8803 13583
rect 8493 13481 8527 13515
rect 9030 13481 9064 13515
rect 6837 13413 6871 13447
rect 6193 13209 6227 13243
rect 9229 13209 9263 13243
rect 1409 12937 1443 12971
rect 8324 13141 8358 13175
rect 8769 13141 8803 13175
rect 6745 13073 6779 13107
rect 6929 13073 6963 13107
rect 9030 13073 9064 13107
rect 9137 13073 9171 13107
rect 9781 13073 9815 13107
rect 9965 13073 9999 13107
rect 8585 13005 8619 13039
rect 9413 13005 9447 13039
rect 7205 12937 7239 12971
rect 9597 12937 9631 12971
rect 9781 12937 9815 12971
rect 6837 12869 6871 12903
rect 8217 12665 8251 12699
rect 8033 12529 8067 12563
rect 6009 12461 6043 12495
rect 7665 12461 7699 12495
rect 7941 12461 7975 12495
rect 8769 12461 8803 12495
rect 6270 12393 6304 12427
rect 7481 12393 7515 12427
rect 7849 12393 7883 12427
rect 9030 12393 9064 12427
rect 6285 12121 6319 12155
rect 7297 12121 7331 12155
rect 7481 12121 7515 12155
rect 9781 12121 9815 12155
rect 8478 12053 8512 12087
rect 6837 11985 6871 12019
rect 7021 11985 7055 12019
rect 7205 11985 7239 12019
rect 9965 11985 9999 12019
rect 6101 11917 6135 11951
rect 6561 11917 6595 11951
rect 6745 11917 6779 11951
rect 8217 11917 8251 11951
rect 6377 11849 6411 11883
rect 10149 11849 10183 11883
rect 6837 11781 6871 11815
rect 9597 11781 9631 11815
rect 10057 11577 10091 11611
rect 7941 11509 7975 11543
rect 6193 11373 6227 11407
rect 7849 11373 7883 11407
rect 8125 11373 8159 11407
rect 8493 11373 8527 11407
rect 6377 11305 6411 11339
rect 7582 11296 7616 11330
rect 8309 11305 8343 11339
rect 8749 11296 8783 11330
rect 6469 11237 6503 11271
rect 9873 11237 9907 11271
rect 6837 11033 6871 11067
rect 10149 11033 10183 11067
rect 6101 10897 6135 10931
rect 6193 10897 6227 10931
rect 6377 10897 6411 10931
rect 6653 10897 6687 10931
rect 8769 10897 8803 10931
rect 9873 10897 9907 10931
rect 6009 10829 6043 10863
rect 6469 10829 6503 10863
rect 10149 10829 10183 10863
rect 7481 10761 7515 10795
rect 8585 10761 8619 10795
rect 5825 10693 5859 10727
rect 6193 10693 6227 10727
rect 9965 10693 9999 10727
rect 10057 10489 10091 10523
rect 6653 10353 6687 10387
rect 6193 10285 6227 10319
rect 6929 10285 6963 10319
rect 8493 10285 8527 10319
rect 2697 10081 2731 10115
rect 7190 10217 7224 10251
rect 8738 10207 8772 10241
rect 6837 10149 6871 10183
rect 8309 10149 8343 10183
rect 9873 10149 9907 10183
rect 9965 10149 9999 10183
rect 9229 9945 9263 9979
rect 7466 9886 7500 9920
rect 10149 9877 10183 9911
rect 5641 9809 5675 9843
rect 6469 9809 6503 9843
rect 6837 9809 6871 9843
rect 7205 9809 7239 9843
rect 9413 9809 9447 9843
rect 9597 9809 9631 9843
rect 9965 9809 9999 9843
rect 6469 9673 6503 9707
rect 6561 9605 6595 9639
rect 7021 9605 7055 9639
rect 9137 9605 9171 9639
rect 9413 9605 9447 9639
rect 9781 9605 9815 9639
rect 6285 9401 6319 9435
rect 6377 9401 6411 9435
rect 8217 9401 8251 9435
rect 7849 9333 7883 9367
rect 8033 9265 8067 9299
rect 6101 9197 6135 9231
rect 7496 9197 7530 9231
rect 7757 9197 7791 9231
rect 8585 9197 8619 9231
rect 8852 9119 8886 9153
rect 6009 8857 6043 8891
rect 9137 8857 9171 8891
rect 10149 8857 10183 8891
rect 7926 8789 7960 8823
rect 6101 8721 6135 8755
rect 6469 8721 6503 8755
rect 7665 8721 7699 8755
rect 9413 8721 9447 8755
rect 9965 8721 9999 8755
rect 6745 8653 6779 8687
rect 7389 8653 7423 8687
rect 9781 8653 9815 8687
rect 7573 8585 7607 8619
rect 9597 8585 9631 8619
rect 7205 8517 7239 8551
rect 9045 8517 9079 8551
rect 7389 8313 7423 8347
rect 9965 8313 9999 8347
rect 7297 8177 7331 8211
rect 7036 8109 7070 8143
rect 7573 8109 7607 8143
rect 7849 8109 7883 8143
rect 8493 8109 8527 8143
rect 7757 8041 7791 8075
rect 8125 8041 8159 8075
rect 8754 8041 8788 8075
rect 7941 7973 7975 8007
rect 9873 7973 9907 8007
rect 5917 7769 5951 7803
rect 6285 7769 6319 7803
rect 9137 7769 9171 7803
rect 5641 7701 5675 7735
rect 7021 7701 7055 7735
rect 7466 7710 7500 7744
rect 9597 7701 9631 7735
rect 2697 7565 2731 7599
rect 6193 7633 6227 7667
rect 6837 7633 6871 7667
rect 7205 7633 7239 7667
rect 9413 7633 9447 7667
rect 9781 7633 9815 7667
rect 9965 7633 9999 7667
rect 6009 7565 6043 7599
rect 6469 7497 6503 7531
rect 6561 7429 6595 7463
rect 8585 7429 8619 7463
rect 9781 7429 9815 7463
rect 6101 7225 6135 7259
rect 8309 7225 8343 7259
rect 6653 7089 6687 7123
rect 9873 7089 9907 7123
rect 6101 7021 6135 7055
rect 6193 7021 6227 7055
rect 6377 7021 6411 7055
rect 6929 7021 6963 7055
rect 8401 7021 8435 7055
rect 6837 6953 6871 6987
rect 7190 6953 7224 6987
rect 9612 6953 9646 6987
rect 10425 6953 10459 6987
rect 6009 6681 6043 6715
rect 6377 6681 6411 6715
rect 7450 6613 7484 6647
rect 6653 6545 6687 6579
rect 7021 6545 7055 6579
rect 9965 6545 9999 6579
rect 9781 6409 9815 6443
rect 6653 6341 6687 6375
rect 8585 6341 8619 6375
rect 8677 6137 8711 6171
rect 9413 6137 9447 6171
rect 9781 6137 9815 6171
rect 6469 6069 6503 6103
rect 6653 6069 6687 6103
rect 7021 6069 7055 6103
rect 8217 6069 8251 6103
rect 6285 6001 6319 6035
rect 7297 6001 7331 6035
rect 6837 5933 6871 5967
rect 7757 5933 7791 5967
rect 8033 5933 8067 5967
rect 8861 5933 8895 5967
rect 9137 5933 9171 5967
rect 9321 5933 9355 5967
rect 9413 5933 9447 5967
rect 9597 5933 9631 5967
rect 9965 5933 9999 5967
rect 10149 5865 10183 5899
rect 6101 5797 6135 5831
rect 6561 5797 6595 5831
rect 1409 85 1443 119
<< metal1 >>
rect 14 17892 20 17944
rect 72 17932 78 17944
rect 109 17935 167 17941
rect 109 17932 121 17935
rect 72 17904 121 17932
rect 72 17892 78 17904
rect 109 17901 121 17904
rect 155 17901 167 17935
rect 109 17895 167 17901
rect 14 17076 20 17128
rect 72 17116 78 17128
rect 5629 17119 5687 17125
rect 5629 17116 5641 17119
rect 72 17088 5641 17116
rect 72 17076 78 17088
rect 5629 17085 5641 17088
rect 5675 17085 5687 17119
rect 5629 17079 5687 17085
rect 5796 14442 10304 14464
rect 5796 14390 8182 14442
rect 8234 14390 8246 14442
rect 8298 14390 8310 14442
rect 8362 14390 8374 14442
rect 8426 14390 8438 14442
rect 8490 14390 8502 14442
rect 8554 14390 8566 14442
rect 8618 14390 8630 14442
rect 8682 14390 8694 14442
rect 8746 14390 8758 14442
rect 8810 14390 10304 14442
rect 5796 14368 10304 14390
rect 5445 14331 5503 14337
rect 5445 14297 5457 14331
rect 5491 14328 5503 14331
rect 6181 14331 6239 14337
rect 6181 14328 6193 14331
rect 5491 14300 6193 14328
rect 5491 14297 5503 14300
rect 5445 14291 5503 14297
rect 6181 14297 6193 14300
rect 6227 14297 6239 14331
rect 6181 14291 6239 14297
rect 6549 14331 6607 14337
rect 6549 14297 6561 14331
rect 6595 14328 6607 14331
rect 8205 14331 8263 14337
rect 6595 14300 6776 14328
rect 6595 14297 6607 14300
rect 6549 14291 6607 14297
rect 6748 14294 6776 14300
rect 8205 14297 8217 14331
rect 8251 14328 8263 14331
rect 8846 14328 8852 14340
rect 8251 14300 8852 14328
rect 8251 14297 8263 14300
rect 6748 14266 7972 14294
rect 8205 14291 8263 14297
rect 8846 14288 8852 14300
rect 8904 14288 8910 14340
rect 7944 14260 7972 14266
rect 8113 14263 8171 14269
rect 7944 14232 8064 14260
rect 109 14195 167 14201
rect 109 14161 121 14195
rect 155 14192 167 14195
rect 6457 14195 6515 14201
rect 6457 14192 6469 14195
rect 155 14164 5396 14192
rect 155 14161 167 14164
rect 109 14155 167 14161
rect 5368 14124 5396 14164
rect 6288 14164 6469 14192
rect 6288 14124 6316 14164
rect 6457 14161 6469 14164
rect 6503 14161 6515 14195
rect 6638 14192 6644 14204
rect 6583 14164 6644 14192
rect 6457 14155 6515 14161
rect 6638 14152 6644 14164
rect 6696 14192 6702 14204
rect 7558 14192 7564 14204
rect 6696 14164 6868 14192
rect 6696 14152 6702 14164
rect 5368 14096 6316 14124
rect 6840 14124 6868 14164
rect 7392 14164 7564 14192
rect 7392 14124 7420 14164
rect 7558 14152 7564 14164
rect 7616 14192 7622 14204
rect 8036 14201 8064 14232
rect 8113 14229 8125 14263
rect 8159 14260 8171 14263
rect 8386 14260 8392 14272
rect 8159 14232 8392 14260
rect 8159 14229 8171 14232
rect 8113 14223 8171 14229
rect 8386 14220 8392 14232
rect 8444 14220 8450 14272
rect 9953 14263 10011 14269
rect 9953 14229 9965 14263
rect 9999 14260 10011 14263
rect 10318 14260 10324 14272
rect 9999 14232 10324 14260
rect 9999 14229 10011 14232
rect 9953 14223 10011 14229
rect 10318 14220 10324 14232
rect 10376 14220 10382 14272
rect 8021 14195 8079 14201
rect 7616 14164 7972 14192
rect 7616 14152 7622 14164
rect 6840 14096 7420 14124
rect 7745 14127 7803 14133
rect 7745 14093 7757 14127
rect 7791 14124 7803 14127
rect 7834 14124 7840 14136
rect 7791 14096 7840 14124
rect 7791 14093 7803 14096
rect 7745 14087 7803 14093
rect 7834 14084 7840 14096
rect 7892 14084 7898 14136
rect 7944 14124 7972 14164
rect 8021 14161 8033 14195
rect 8067 14161 8079 14195
rect 8021 14155 8079 14161
rect 8202 14152 8208 14204
rect 8260 14192 8266 14204
rect 8297 14195 8355 14201
rect 8297 14192 8309 14195
rect 8260 14164 8309 14192
rect 8260 14152 8266 14164
rect 8297 14161 8309 14164
rect 8343 14161 8355 14195
rect 8665 14195 8723 14201
rect 8665 14192 8677 14195
rect 8297 14155 8355 14161
rect 8404 14164 8677 14192
rect 8404 14124 8432 14164
rect 8665 14161 8677 14164
rect 8711 14192 8723 14195
rect 9858 14192 9864 14204
rect 8711 14164 9864 14192
rect 8711 14161 8723 14164
rect 8665 14155 8723 14161
rect 9858 14152 9864 14164
rect 9916 14152 9922 14204
rect 10137 14195 10195 14201
rect 10137 14161 10149 14195
rect 10183 14161 10195 14195
rect 10137 14155 10195 14161
rect 10229 14195 10287 14201
rect 10229 14161 10241 14195
rect 10275 14192 10287 14195
rect 15838 14192 15844 14204
rect 10275 14164 15844 14192
rect 10275 14161 10287 14164
rect 10229 14155 10287 14161
rect 7944 14096 8432 14124
rect 7561 14059 7619 14065
rect 7561 14025 7573 14059
rect 7607 14056 7619 14059
rect 8757 14059 8815 14065
rect 8757 14056 8769 14059
rect 7607 14028 8769 14056
rect 7607 14025 7619 14028
rect 7561 14019 7619 14025
rect 8757 14025 8769 14028
rect 8803 14056 8815 14059
rect 9125 14059 9183 14065
rect 9125 14056 9137 14059
rect 8803 14028 9137 14056
rect 8803 14025 8815 14028
rect 8757 14019 8815 14025
rect 9125 14025 9137 14028
rect 9171 14025 9183 14059
rect 10152 14056 10180 14155
rect 15838 14152 15844 14164
rect 15896 14152 15902 14204
rect 9125 14019 9183 14025
rect 9876 14028 10180 14056
rect 7929 13991 7987 13997
rect 7929 13957 7941 13991
rect 7975 13988 7987 13991
rect 8202 13988 8208 14000
rect 7975 13960 8208 13988
rect 7975 13957 7987 13960
rect 7929 13951 7987 13957
rect 8202 13948 8208 13960
rect 8260 13948 8266 14000
rect 8662 13948 8668 14000
rect 8720 13988 8726 14000
rect 8941 13991 8999 13997
rect 8941 13988 8953 13991
rect 8720 13960 8953 13988
rect 8720 13948 8726 13960
rect 8941 13957 8953 13960
rect 8987 13957 8999 13991
rect 9306 13988 9312 14000
rect 9251 13960 9312 13988
rect 8941 13951 8999 13957
rect 9306 13948 9312 13960
rect 9364 13988 9370 14000
rect 9876 13988 9904 14028
rect 9364 13960 9904 13988
rect 9953 13991 10011 13997
rect 9364 13948 9370 13960
rect 9953 13957 9965 13991
rect 9999 13988 10011 13991
rect 10134 13988 10140 14000
rect 9999 13960 10140 13988
rect 9999 13957 10011 13960
rect 9953 13951 10011 13957
rect 10134 13948 10140 13960
rect 10192 13948 10198 14000
rect 5796 13898 10304 13920
rect 5796 13846 5800 13898
rect 5852 13846 5864 13898
rect 5916 13846 5928 13898
rect 5980 13846 5992 13898
rect 6044 13846 6056 13898
rect 6108 13846 10304 13898
rect 5796 13824 10304 13846
rect 14 13744 20 13796
rect 72 13784 78 13796
rect 6733 13787 6791 13793
rect 6733 13784 6745 13787
rect 72 13756 5764 13784
rect 72 13744 78 13756
rect 5736 13648 5764 13756
rect 6564 13756 6745 13784
rect 6564 13648 6592 13756
rect 6733 13753 6745 13756
rect 6779 13753 6791 13787
rect 6733 13747 6791 13753
rect 8573 13787 8631 13793
rect 8573 13753 8585 13787
rect 8619 13784 8631 13787
rect 8662 13784 8668 13796
rect 8619 13756 8668 13784
rect 8619 13753 8631 13756
rect 8573 13747 8631 13753
rect 8662 13744 8668 13756
rect 8720 13784 8726 13796
rect 9490 13784 9496 13796
rect 8720 13756 9496 13784
rect 8720 13744 8726 13756
rect 9490 13744 9496 13756
rect 9548 13744 9554 13796
rect 10137 13787 10195 13793
rect 10137 13753 10149 13787
rect 10183 13784 10195 13787
rect 16022 13784 16028 13796
rect 10183 13756 16028 13784
rect 10183 13753 10195 13756
rect 10137 13747 10195 13753
rect 16022 13744 16028 13756
rect 16080 13744 16086 13796
rect 6822 13676 6828 13728
rect 6880 13716 6886 13728
rect 6917 13719 6975 13725
rect 6917 13716 6929 13719
rect 6880 13688 6929 13716
rect 6880 13676 6886 13688
rect 6917 13685 6929 13688
rect 6963 13716 6975 13719
rect 6963 13688 7328 13716
rect 6963 13685 6975 13688
rect 6917 13679 6975 13685
rect 5736 13620 6592 13648
rect 7300 13512 7328 13688
rect 8036 13583 8094 13589
rect 8036 13549 8048 13583
rect 8082 13580 8094 13583
rect 8202 13580 8208 13592
rect 8082 13552 8208 13580
rect 8082 13549 8094 13552
rect 8036 13543 8094 13549
rect 8202 13540 8208 13552
rect 8260 13540 8266 13592
rect 8297 13583 8355 13589
rect 8297 13549 8309 13583
rect 8343 13580 8355 13583
rect 8757 13583 8815 13589
rect 8757 13580 8769 13583
rect 8343 13552 8769 13580
rect 8343 13549 8355 13552
rect 8297 13543 8355 13549
rect 8757 13549 8769 13552
rect 8803 13580 8815 13583
rect 8846 13580 8852 13592
rect 8803 13552 8852 13580
rect 8803 13549 8815 13552
rect 8757 13543 8815 13549
rect 8846 13540 8852 13552
rect 8904 13540 8910 13592
rect 8386 13512 8392 13524
rect 7300 13484 8392 13512
rect 8386 13472 8392 13484
rect 8444 13512 8450 13524
rect 8481 13515 8539 13521
rect 8481 13512 8493 13515
rect 8444 13484 8493 13512
rect 8444 13472 8450 13484
rect 8481 13481 8493 13484
rect 8527 13481 8539 13515
rect 8481 13475 8539 13481
rect 9018 13515 9076 13521
rect 9018 13481 9030 13515
rect 9064 13512 9076 13515
rect 9214 13512 9220 13524
rect 9064 13484 9220 13512
rect 9064 13481 9076 13484
rect 9018 13475 9076 13481
rect 9214 13472 9220 13484
rect 9272 13472 9278 13524
rect 6825 13447 6883 13453
rect 6825 13413 6837 13447
rect 6871 13444 6883 13447
rect 7006 13444 7012 13456
rect 6871 13416 7012 13444
rect 6871 13413 6883 13416
rect 6825 13407 6883 13413
rect 7006 13404 7012 13416
rect 7064 13404 7070 13456
rect 5796 13354 10304 13376
rect 5796 13302 8182 13354
rect 8234 13302 8246 13354
rect 8298 13302 8310 13354
rect 8362 13302 8374 13354
rect 8426 13302 8438 13354
rect 8490 13302 8502 13354
rect 8554 13302 8566 13354
rect 8618 13302 8630 13354
rect 8682 13302 8694 13354
rect 8746 13302 8758 13354
rect 8810 13302 10304 13354
rect 5796 13280 10304 13302
rect 14 13200 20 13252
rect 72 13240 78 13252
rect 6181 13243 6239 13249
rect 6181 13240 6193 13243
rect 72 13212 6193 13240
rect 72 13200 78 13212
rect 6181 13209 6193 13212
rect 6227 13209 6239 13243
rect 9214 13240 9220 13252
rect 9159 13212 9220 13240
rect 6181 13203 6239 13209
rect 9214 13200 9220 13212
rect 9272 13200 9278 13252
rect 8312 13175 8370 13181
rect 8312 13141 8324 13175
rect 8358 13172 8370 13175
rect 8757 13175 8815 13181
rect 8757 13172 8769 13175
rect 8358 13144 8769 13172
rect 8358 13141 8370 13144
rect 8312 13135 8370 13141
rect 8757 13141 8769 13144
rect 8803 13141 8815 13175
rect 8757 13135 8815 13141
rect 6638 13064 6644 13116
rect 6696 13104 6702 13116
rect 6733 13107 6791 13113
rect 6733 13104 6745 13107
rect 6696 13076 6745 13104
rect 6696 13064 6702 13076
rect 6733 13073 6745 13076
rect 6779 13073 6791 13107
rect 6733 13067 6791 13073
rect 6822 13064 6828 13116
rect 6880 13104 6886 13116
rect 6917 13107 6975 13113
rect 6917 13104 6929 13107
rect 6880 13076 6929 13104
rect 6880 13064 6886 13076
rect 6917 13073 6929 13076
rect 6963 13073 6975 13107
rect 6917 13067 6975 13073
rect 8018 13064 8024 13116
rect 8076 13104 8082 13116
rect 9018 13107 9076 13113
rect 9018 13104 9030 13107
rect 8076 13076 9030 13104
rect 8076 13064 8082 13076
rect 9018 13073 9030 13076
rect 9064 13073 9076 13107
rect 9018 13067 9076 13073
rect 9125 13107 9183 13113
rect 9125 13073 9137 13107
rect 9171 13104 9183 13107
rect 9306 13104 9312 13116
rect 9171 13076 9312 13104
rect 9171 13073 9183 13076
rect 9125 13067 9183 13073
rect 8573 13039 8631 13045
rect 5736 13008 6500 13036
rect 1397 12971 1455 12977
rect 1397 12937 1409 12971
rect 1443 12968 1455 12971
rect 5736 12968 5764 13008
rect 6472 13002 6500 13008
rect 8573 13005 8585 13039
rect 8619 13036 8631 13039
rect 8846 13036 8852 13048
rect 8619 13008 8852 13036
rect 8619 13005 8631 13008
rect 6472 12974 7052 13002
rect 8573 12999 8631 13005
rect 8846 12996 8852 13008
rect 8904 12996 8910 13048
rect 9033 13036 9061 13067
rect 9306 13064 9312 13076
rect 9364 13064 9370 13116
rect 9490 13064 9496 13116
rect 9548 13104 9554 13116
rect 9769 13107 9827 13113
rect 9769 13104 9781 13107
rect 9548 13076 9781 13104
rect 9548 13064 9554 13076
rect 9769 13073 9781 13076
rect 9815 13073 9827 13107
rect 9769 13067 9827 13073
rect 9858 13064 9864 13116
rect 9916 13104 9922 13116
rect 9953 13107 10011 13113
rect 9953 13104 9965 13107
rect 9916 13076 9965 13104
rect 9916 13064 9922 13076
rect 9953 13073 9965 13076
rect 9999 13073 10011 13107
rect 9953 13067 10011 13073
rect 9214 13036 9220 13048
rect 9033 13008 9220 13036
rect 9214 12996 9220 13008
rect 9272 13036 9278 13048
rect 9401 13039 9459 13045
rect 9401 13036 9413 13039
rect 9272 13008 9413 13036
rect 9272 12996 9278 13008
rect 9401 13005 9413 13008
rect 9447 13005 9459 13039
rect 9401 12999 9459 13005
rect 1443 12940 5764 12968
rect 7024 12968 7052 12974
rect 7193 12971 7251 12977
rect 7193 12968 7205 12971
rect 7024 12940 7205 12968
rect 1443 12937 1455 12940
rect 1397 12931 1455 12937
rect 7193 12937 7205 12940
rect 7239 12937 7251 12971
rect 7193 12931 7251 12937
rect 9585 12971 9643 12977
rect 9585 12937 9597 12971
rect 9631 12968 9643 12971
rect 9769 12971 9827 12977
rect 9769 12968 9781 12971
rect 9631 12940 9781 12968
rect 9631 12937 9643 12940
rect 9585 12931 9643 12937
rect 9769 12937 9781 12940
rect 9815 12968 9827 12971
rect 10318 12968 10324 12980
rect 9815 12940 10324 12968
rect 9815 12937 9827 12940
rect 9769 12931 9827 12937
rect 10318 12928 10324 12940
rect 10376 12928 10382 12980
rect 6638 12860 6644 12912
rect 6696 12900 6702 12912
rect 6825 12903 6883 12909
rect 6825 12900 6837 12903
rect 6696 12872 6837 12900
rect 6696 12860 6702 12872
rect 6825 12869 6837 12872
rect 6871 12869 6883 12903
rect 6825 12863 6883 12869
rect 5796 12810 10304 12832
rect 5796 12758 5800 12810
rect 5852 12758 5864 12810
rect 5916 12758 5928 12810
rect 5980 12758 5992 12810
rect 6044 12758 6056 12810
rect 6108 12758 10304 12810
rect 5796 12736 10304 12758
rect 6914 12656 6920 12708
rect 6972 12696 6978 12708
rect 8205 12699 8263 12705
rect 8205 12696 8217 12699
rect 6972 12668 7144 12696
rect 6972 12656 6978 12668
rect 7116 12662 7144 12668
rect 8036 12668 8217 12696
rect 8036 12662 8064 12668
rect 7116 12634 8064 12662
rect 8205 12665 8217 12668
rect 8251 12665 8263 12699
rect 8205 12659 8263 12665
rect 7558 12520 7564 12572
rect 7616 12560 7622 12572
rect 7616 12532 7788 12560
rect 7616 12520 7622 12532
rect 5997 12495 6055 12501
rect 5997 12461 6009 12495
rect 6043 12492 6055 12495
rect 6730 12492 6736 12504
rect 6043 12464 6736 12492
rect 6043 12461 6055 12464
rect 5997 12455 6055 12461
rect 6730 12452 6736 12464
rect 6788 12452 6794 12504
rect 7653 12495 7711 12501
rect 7653 12492 7665 12495
rect 6840 12464 7665 12492
rect 6258 12427 6316 12433
rect 6258 12424 6270 12427
rect 5736 12396 6270 12424
rect 5736 12152 5764 12396
rect 6258 12393 6270 12396
rect 6304 12393 6316 12427
rect 6258 12387 6316 12393
rect 6638 12384 6644 12436
rect 6696 12424 6702 12436
rect 6840 12424 6868 12464
rect 7653 12461 7665 12464
rect 7699 12461 7711 12495
rect 7760 12492 7788 12532
rect 7834 12520 7840 12572
rect 7892 12560 7898 12572
rect 8021 12563 8079 12569
rect 8021 12560 8033 12563
rect 7892 12532 8033 12560
rect 7892 12520 7898 12532
rect 8021 12529 8033 12532
rect 8067 12529 8079 12563
rect 8021 12523 8079 12529
rect 7929 12495 7987 12501
rect 7929 12492 7941 12495
rect 7760 12464 7941 12492
rect 7653 12455 7711 12461
rect 7929 12461 7941 12464
rect 7975 12461 7987 12495
rect 7929 12455 7987 12461
rect 8757 12495 8815 12501
rect 8757 12461 8769 12495
rect 8803 12492 8815 12495
rect 8846 12492 8852 12504
rect 8803 12464 8852 12492
rect 8803 12461 8815 12464
rect 8757 12455 8815 12461
rect 8846 12452 8852 12464
rect 8904 12452 8910 12504
rect 7466 12424 7472 12436
rect 6696 12396 6868 12424
rect 7411 12396 7472 12424
rect 6696 12384 6702 12396
rect 7466 12384 7472 12396
rect 7524 12384 7530 12436
rect 7742 12384 7748 12436
rect 7800 12424 7806 12436
rect 7837 12427 7895 12433
rect 7837 12424 7849 12427
rect 7800 12396 7849 12424
rect 7800 12384 7806 12396
rect 7837 12393 7849 12396
rect 7883 12393 7895 12427
rect 7837 12387 7895 12393
rect 9018 12427 9076 12433
rect 9018 12393 9030 12427
rect 9064 12424 9076 12427
rect 9064 12396 10364 12424
rect 9064 12393 9076 12396
rect 9018 12387 9076 12393
rect 5796 12266 10304 12288
rect 5796 12214 8182 12266
rect 8234 12214 8246 12266
rect 8298 12214 8310 12266
rect 8362 12214 8374 12266
rect 8426 12214 8438 12266
rect 8490 12214 8502 12266
rect 8554 12214 8566 12266
rect 8618 12214 8630 12266
rect 8682 12214 8694 12266
rect 8746 12214 8758 12266
rect 8810 12214 10304 12266
rect 5796 12192 10304 12214
rect 6273 12155 6331 12161
rect 6273 12152 6285 12155
rect 5736 12124 6285 12152
rect 6273 12121 6285 12124
rect 6319 12121 6331 12155
rect 6273 12115 6331 12121
rect 7006 12112 7012 12164
rect 7064 12152 7070 12164
rect 7285 12155 7343 12161
rect 7285 12152 7297 12155
rect 7064 12124 7297 12152
rect 7064 12112 7070 12124
rect 7285 12121 7297 12124
rect 7331 12121 7343 12155
rect 7466 12152 7472 12164
rect 7411 12124 7472 12152
rect 7285 12115 7343 12121
rect 7466 12112 7472 12124
rect 7524 12112 7530 12164
rect 9769 12155 9827 12161
rect 9769 12121 9781 12155
rect 9815 12152 9827 12155
rect 10336 12152 10364 12396
rect 9815 12124 10364 12152
rect 9815 12121 9827 12124
rect 9769 12115 9827 12121
rect 6178 11976 6184 12028
rect 6236 12016 6242 12028
rect 6638 12016 6644 12028
rect 6236 11988 6644 12016
rect 6236 11976 6242 11988
rect 6638 11976 6644 11988
rect 6696 12016 6702 12028
rect 7024 12025 7052 12112
rect 8466 12087 8524 12093
rect 8466 12084 8478 12087
rect 7116 12056 8478 12084
rect 6825 12019 6883 12025
rect 6825 12016 6837 12019
rect 6696 11988 6837 12016
rect 6696 11976 6702 11988
rect 6825 11985 6837 11988
rect 6871 11985 6883 12019
rect 6825 11979 6883 11985
rect 7009 12019 7067 12025
rect 7009 11985 7021 12019
rect 7055 11985 7067 12019
rect 7009 11979 7067 11985
rect 6089 11951 6147 11957
rect 6089 11917 6101 11951
rect 6135 11948 6147 11951
rect 6546 11948 6552 11960
rect 6135 11920 6552 11948
rect 6135 11917 6147 11920
rect 6089 11911 6147 11917
rect 6546 11908 6552 11920
rect 6604 11908 6610 11960
rect 6733 11951 6791 11957
rect 6733 11917 6745 11951
rect 6779 11948 6791 11951
rect 7116 11948 7144 12056
rect 8466 12053 8478 12056
rect 8512 12053 8524 12087
rect 8466 12047 8524 12053
rect 7193 12019 7251 12025
rect 7193 11985 7205 12019
rect 7239 11985 7251 12019
rect 7193 11979 7251 11985
rect 6779 11920 7144 11948
rect 6779 11917 6791 11920
rect 6733 11911 6791 11917
rect 6365 11883 6423 11889
rect 6365 11849 6377 11883
rect 6411 11880 6423 11883
rect 6411 11852 6684 11880
rect 6411 11849 6423 11852
rect 6365 11843 6423 11849
rect 6656 11812 6684 11852
rect 6825 11815 6883 11821
rect 6825 11812 6837 11815
rect 6656 11784 6837 11812
rect 6825 11781 6837 11784
rect 6871 11781 6883 11815
rect 7208 11812 7236 11979
rect 9214 11976 9220 12028
rect 9272 12016 9278 12028
rect 9953 12019 10011 12025
rect 9953 12016 9965 12019
rect 9272 11988 9965 12016
rect 9272 11976 9278 11988
rect 9953 11985 9965 11988
rect 9999 11985 10011 12019
rect 9953 11979 10011 11985
rect 7558 11908 7564 11960
rect 7616 11948 7622 11960
rect 8205 11951 8263 11957
rect 8205 11948 8217 11951
rect 7616 11920 8217 11948
rect 7616 11908 7622 11920
rect 8205 11917 8217 11920
rect 8251 11917 8263 11951
rect 8205 11911 8263 11917
rect 10137 11883 10195 11889
rect 10137 11849 10149 11883
rect 10183 11880 10195 11883
rect 10318 11880 10324 11892
rect 10183 11852 10324 11880
rect 10183 11849 10195 11852
rect 10137 11843 10195 11849
rect 10318 11840 10324 11852
rect 10376 11840 10382 11892
rect 9585 11815 9643 11821
rect 9585 11812 9597 11815
rect 7208 11784 9597 11812
rect 6825 11775 6883 11781
rect 9585 11781 9597 11784
rect 9631 11781 9643 11815
rect 9585 11775 9643 11781
rect 5796 11722 10304 11744
rect 5796 11670 5800 11722
rect 5852 11670 5864 11722
rect 5916 11670 5928 11722
rect 5980 11670 5992 11722
rect 6044 11670 6056 11722
rect 6108 11670 10304 11722
rect 5796 11648 10304 11670
rect 7650 11568 7656 11620
rect 7708 11608 7714 11620
rect 7708 11580 7880 11608
rect 7708 11568 7714 11580
rect 7852 11540 7880 11580
rect 9858 11568 9864 11620
rect 9916 11608 9922 11620
rect 10045 11611 10103 11617
rect 10045 11608 10057 11611
rect 9916 11580 10057 11608
rect 9916 11568 9922 11580
rect 10045 11577 10057 11580
rect 10091 11577 10103 11611
rect 10045 11571 10103 11577
rect 7929 11543 7987 11549
rect 7929 11540 7941 11543
rect 7852 11512 7941 11540
rect 7929 11509 7941 11512
rect 7975 11509 7987 11543
rect 7929 11503 7987 11509
rect 6086 11364 6092 11416
rect 6144 11404 6150 11416
rect 6181 11407 6239 11413
rect 6181 11404 6193 11407
rect 6144 11376 6193 11404
rect 6144 11364 6150 11376
rect 6181 11373 6193 11376
rect 6227 11373 6239 11407
rect 6181 11367 6239 11373
rect 7558 11364 7564 11416
rect 7616 11404 7622 11416
rect 7837 11407 7895 11413
rect 7837 11404 7849 11407
rect 7616 11376 7849 11404
rect 7616 11364 7622 11376
rect 7837 11373 7849 11376
rect 7883 11373 7895 11407
rect 7837 11367 7895 11373
rect 8018 11364 8024 11416
rect 8076 11404 8082 11416
rect 8113 11407 8171 11413
rect 8113 11404 8125 11407
rect 8076 11376 8125 11404
rect 8076 11364 8082 11376
rect 8113 11373 8125 11376
rect 8159 11373 8171 11407
rect 8113 11367 8171 11373
rect 8481 11407 8539 11413
rect 8481 11373 8493 11407
rect 8527 11404 8539 11407
rect 8754 11404 8760 11416
rect 8527 11376 8760 11404
rect 8527 11373 8539 11376
rect 8481 11367 8539 11373
rect 8754 11364 8760 11376
rect 8812 11364 8818 11416
rect 6362 11336 6368 11348
rect 6307 11308 6368 11336
rect 6362 11296 6368 11308
rect 6420 11296 6426 11348
rect 8297 11339 8355 11345
rect 7570 11330 7628 11336
rect 7570 11327 7582 11330
rect 7484 11299 7582 11327
rect 6457 11271 6515 11277
rect 6457 11268 6469 11271
rect 5736 11240 6469 11268
rect 5736 11064 5764 11240
rect 6457 11237 6469 11240
rect 6503 11237 6515 11271
rect 6457 11231 6515 11237
rect 7282 11228 7288 11280
rect 7340 11268 7346 11280
rect 7484 11268 7512 11299
rect 7570 11296 7582 11299
rect 7616 11296 7628 11330
rect 8297 11305 8309 11339
rect 8343 11336 8355 11339
rect 8343 11330 8795 11336
rect 8343 11308 8749 11330
rect 8343 11305 8355 11308
rect 8297 11299 8355 11305
rect 7570 11290 7628 11296
rect 8737 11296 8749 11308
rect 8783 11296 8795 11330
rect 8737 11290 8795 11296
rect 7340 11240 7512 11268
rect 9861 11271 9919 11277
rect 7340 11228 7346 11240
rect 9861 11237 9873 11271
rect 9907 11268 9919 11271
rect 9950 11268 9956 11280
rect 9907 11240 9956 11268
rect 9907 11237 9919 11240
rect 9861 11231 9919 11237
rect 9950 11228 9956 11240
rect 10008 11228 10014 11280
rect 5796 11178 10304 11200
rect 5796 11126 8182 11178
rect 8234 11126 8246 11178
rect 8298 11126 8310 11178
rect 8362 11126 8374 11178
rect 8426 11126 8438 11178
rect 8490 11126 8502 11178
rect 8554 11126 8566 11178
rect 8618 11126 8630 11178
rect 8682 11126 8694 11178
rect 8746 11126 8758 11178
rect 8810 11126 10304 11178
rect 5796 11104 10304 11126
rect 6825 11067 6883 11073
rect 5736 11036 6224 11064
rect 6086 10928 6092 10940
rect 6031 10900 6092 10928
rect 6086 10888 6092 10900
rect 6144 10888 6150 10940
rect 6196 10937 6224 11036
rect 6825 11033 6837 11067
rect 6871 11064 6883 11067
rect 7282 11064 7288 11076
rect 6871 11036 7288 11064
rect 6871 11033 6883 11036
rect 6825 11027 6883 11033
rect 7282 11024 7288 11036
rect 7340 11024 7346 11076
rect 7834 11064 7840 11076
rect 7576 11036 7840 11064
rect 6181 10931 6239 10937
rect 6181 10897 6193 10931
rect 6227 10897 6239 10931
rect 6362 10928 6368 10940
rect 6307 10900 6368 10928
rect 6181 10891 6239 10897
rect 6362 10888 6368 10900
rect 6420 10888 6426 10940
rect 6546 10888 6552 10940
rect 6604 10928 6610 10940
rect 6641 10931 6699 10937
rect 6641 10928 6653 10931
rect 6604 10900 6653 10928
rect 6604 10888 6610 10900
rect 6641 10897 6653 10900
rect 6687 10928 6699 10931
rect 7576 10928 7604 11036
rect 7834 11024 7840 11036
rect 7892 11024 7898 11076
rect 10137 11067 10195 11073
rect 10137 11033 10149 11067
rect 10183 11064 10195 11067
rect 10318 11064 10324 11076
rect 10183 11036 10324 11064
rect 10183 11033 10195 11036
rect 10137 11027 10195 11033
rect 10318 11024 10324 11036
rect 10376 11024 10382 11076
rect 6687 10900 7604 10928
rect 6687 10897 6699 10900
rect 6641 10891 6699 10897
rect 7650 10888 7656 10940
rect 7708 10888 7714 10940
rect 8757 10931 8815 10937
rect 8757 10897 8769 10931
rect 8803 10928 8815 10931
rect 9490 10928 9496 10940
rect 8803 10900 9496 10928
rect 8803 10897 8815 10900
rect 8757 10891 8815 10897
rect 9490 10888 9496 10900
rect 9548 10888 9554 10940
rect 9582 10888 9588 10940
rect 9640 10928 9646 10940
rect 9861 10931 9919 10937
rect 9861 10928 9873 10931
rect 9640 10900 9873 10928
rect 9640 10888 9646 10900
rect 9861 10897 9873 10900
rect 9907 10897 9919 10931
rect 9861 10891 9919 10897
rect 5997 10863 6055 10869
rect 5997 10829 6009 10863
rect 6043 10860 6055 10863
rect 6457 10863 6515 10869
rect 6457 10860 6469 10863
rect 6043 10832 6469 10860
rect 6043 10829 6055 10832
rect 5997 10823 6055 10829
rect 6457 10829 6469 10832
rect 6503 10829 6515 10863
rect 10134 10860 10140 10872
rect 10079 10832 10140 10860
rect 6457 10823 6515 10829
rect 10134 10820 10140 10832
rect 10192 10820 10198 10872
rect 7466 10792 7472 10804
rect 7411 10764 7472 10792
rect 7466 10752 7472 10764
rect 7524 10752 7530 10804
rect 8573 10795 8631 10801
rect 8573 10761 8585 10795
rect 8619 10792 8631 10795
rect 9030 10792 9036 10804
rect 8619 10764 9036 10792
rect 8619 10761 8631 10764
rect 8573 10755 8631 10761
rect 9030 10752 9036 10764
rect 9088 10752 9094 10804
rect 5813 10727 5871 10733
rect 5813 10693 5825 10727
rect 5859 10724 5871 10727
rect 6181 10727 6239 10733
rect 6181 10724 6193 10727
rect 5859 10696 6193 10724
rect 5859 10693 5871 10696
rect 5813 10687 5871 10693
rect 6181 10693 6193 10696
rect 6227 10693 6239 10727
rect 6181 10687 6239 10693
rect 9953 10727 10011 10733
rect 9953 10693 9965 10727
rect 9999 10724 10011 10727
rect 9999 10696 10364 10724
rect 9999 10693 10011 10696
rect 9953 10687 10011 10693
rect 5796 10634 10304 10656
rect 5796 10582 5800 10634
rect 5852 10582 5864 10634
rect 5916 10582 5928 10634
rect 5980 10582 5992 10634
rect 6044 10582 6056 10634
rect 6108 10582 10304 10634
rect 5796 10560 10304 10582
rect 10045 10523 10103 10529
rect 10045 10489 10057 10523
rect 10091 10520 10103 10523
rect 10336 10520 10364 10696
rect 10091 10492 10364 10520
rect 10091 10489 10103 10492
rect 10045 10483 10103 10489
rect 6546 10344 6552 10396
rect 6604 10384 6610 10396
rect 6641 10387 6699 10393
rect 6641 10384 6653 10387
rect 6604 10356 6653 10384
rect 6604 10344 6610 10356
rect 6641 10353 6653 10356
rect 6687 10353 6699 10387
rect 6641 10347 6699 10353
rect 6178 10316 6184 10328
rect 6123 10288 6184 10316
rect 6178 10276 6184 10288
rect 6236 10276 6242 10328
rect 6917 10319 6975 10325
rect 6917 10285 6929 10319
rect 6963 10316 6975 10319
rect 7466 10316 7472 10328
rect 6963 10288 7472 10316
rect 6963 10285 6975 10288
rect 6917 10279 6975 10285
rect 7466 10276 7472 10288
rect 7524 10276 7530 10328
rect 8481 10319 8539 10325
rect 8481 10285 8493 10319
rect 8527 10316 8539 10319
rect 8754 10316 8760 10328
rect 8527 10288 8760 10316
rect 8527 10285 8539 10288
rect 8481 10279 8539 10285
rect 8754 10276 8760 10288
rect 8812 10276 8818 10328
rect 7190 10257 7196 10260
rect 7178 10251 7196 10257
rect 7178 10248 7190 10251
rect 7135 10220 7190 10248
rect 7178 10217 7190 10220
rect 7178 10211 7196 10217
rect 7190 10208 7196 10211
rect 7248 10208 7254 10260
rect 7926 10208 7932 10260
rect 7984 10248 7990 10260
rect 7984 10238 8432 10248
rect 8726 10241 8784 10247
rect 8726 10238 8738 10241
rect 7984 10220 8738 10238
rect 7984 10208 7990 10220
rect 8404 10210 8738 10220
rect 8726 10207 8738 10210
rect 8772 10207 8784 10241
rect 8726 10201 8784 10207
rect 6825 10183 6883 10189
rect 6825 10149 6837 10183
rect 6871 10180 6883 10183
rect 7006 10180 7012 10192
rect 6871 10152 7012 10180
rect 6871 10149 6883 10152
rect 6825 10143 6883 10149
rect 7006 10140 7012 10152
rect 7064 10140 7070 10192
rect 8294 10180 8300 10192
rect 8239 10152 8300 10180
rect 8294 10140 8300 10152
rect 8352 10140 8358 10192
rect 9858 10180 9864 10192
rect 9803 10152 9864 10180
rect 9858 10140 9864 10152
rect 9916 10140 9922 10192
rect 9950 10140 9956 10192
rect 10008 10180 10014 10192
rect 10008 10152 10364 10180
rect 10008 10140 10014 10152
rect 14 10072 20 10124
rect 72 10112 78 10124
rect 2685 10115 2743 10121
rect 2685 10112 2697 10115
rect 72 10084 2697 10112
rect 72 10072 78 10084
rect 2685 10081 2697 10084
rect 2731 10081 2743 10115
rect 2685 10075 2743 10081
rect 5796 10090 10304 10112
rect 5796 10038 8182 10090
rect 8234 10038 8246 10090
rect 8298 10038 8310 10090
rect 8362 10038 8374 10090
rect 8426 10038 8438 10090
rect 8490 10038 8502 10090
rect 8554 10038 8566 10090
rect 8618 10038 8630 10090
rect 8682 10038 8694 10090
rect 8746 10038 8758 10090
rect 8810 10038 10304 10090
rect 5796 10016 10304 10038
rect 9217 9979 9275 9985
rect 9217 9945 9229 9979
rect 9263 9976 9275 9979
rect 10336 9976 10364 10152
rect 9263 9948 10364 9976
rect 9263 9945 9275 9948
rect 9217 9939 9275 9945
rect 7454 9920 7512 9926
rect 7006 9868 7012 9920
rect 7064 9908 7070 9920
rect 7454 9908 7466 9920
rect 7064 9886 7466 9908
rect 7500 9886 7512 9920
rect 7064 9880 7512 9886
rect 7064 9868 7070 9880
rect 9858 9868 9864 9920
rect 9916 9908 9922 9920
rect 10137 9911 10195 9917
rect 10137 9908 10149 9911
rect 9916 9880 10149 9908
rect 9916 9868 9922 9880
rect 10137 9877 10149 9880
rect 10183 9877 10195 9911
rect 10137 9871 10195 9877
rect 5629 9843 5687 9849
rect 5629 9809 5641 9843
rect 5675 9840 5687 9843
rect 6454 9840 6460 9852
rect 5675 9812 5948 9840
rect 6399 9812 6460 9840
rect 5675 9809 5687 9812
rect 5629 9803 5687 9809
rect 5920 9772 5948 9812
rect 6454 9800 6460 9812
rect 6512 9800 6518 9852
rect 6546 9800 6552 9852
rect 6604 9840 6610 9852
rect 6825 9843 6883 9849
rect 6825 9840 6837 9843
rect 6604 9812 6837 9840
rect 6604 9800 6610 9812
rect 6825 9809 6837 9812
rect 6871 9809 6883 9843
rect 6825 9803 6883 9809
rect 7193 9843 7251 9849
rect 7193 9809 7205 9843
rect 7239 9840 7251 9843
rect 7466 9840 7472 9852
rect 7239 9812 7472 9840
rect 7239 9809 7251 9812
rect 7193 9803 7251 9809
rect 7466 9800 7472 9812
rect 7524 9800 7530 9852
rect 9398 9840 9404 9852
rect 9343 9812 9404 9840
rect 9398 9800 9404 9812
rect 9456 9800 9462 9852
rect 9585 9843 9643 9849
rect 9585 9809 9597 9843
rect 9631 9840 9643 9843
rect 9876 9840 9904 9868
rect 9631 9812 9904 9840
rect 9631 9809 9643 9812
rect 9585 9803 9643 9809
rect 9950 9800 9956 9852
rect 10008 9840 10014 9852
rect 10008 9812 10069 9840
rect 10008 9800 10014 9812
rect 5920 9744 7144 9772
rect 6454 9704 6460 9716
rect 6399 9676 6460 9704
rect 6454 9664 6460 9676
rect 6512 9664 6518 9716
rect 6549 9639 6607 9645
rect 6549 9636 6561 9639
rect 5736 9608 6561 9636
rect 5736 9432 5764 9608
rect 6549 9605 6561 9608
rect 6595 9605 6607 9639
rect 7006 9636 7012 9648
rect 6951 9608 7012 9636
rect 6549 9599 6607 9605
rect 7006 9596 7012 9608
rect 7064 9596 7070 9648
rect 7116 9636 7144 9744
rect 8312 9676 8984 9704
rect 8312 9636 8340 9676
rect 7116 9608 8340 9636
rect 8956 9636 8984 9676
rect 9125 9639 9183 9645
rect 9125 9636 9137 9639
rect 8956 9608 9137 9636
rect 9125 9605 9137 9608
rect 9171 9605 9183 9639
rect 9125 9599 9183 9605
rect 9306 9596 9312 9648
rect 9364 9636 9370 9648
rect 9401 9639 9459 9645
rect 9401 9636 9413 9639
rect 9364 9608 9413 9636
rect 9364 9596 9370 9608
rect 9401 9605 9413 9608
rect 9447 9605 9459 9639
rect 9766 9636 9772 9648
rect 9711 9608 9772 9636
rect 9401 9599 9459 9605
rect 9766 9596 9772 9608
rect 9824 9596 9830 9648
rect 5796 9546 10304 9568
rect 5796 9494 5800 9546
rect 5852 9494 5864 9546
rect 5916 9494 5928 9546
rect 5980 9494 5992 9546
rect 6044 9494 6056 9546
rect 6108 9494 10304 9546
rect 5796 9472 10304 9494
rect 6273 9435 6331 9441
rect 6273 9432 6285 9435
rect 5736 9404 6285 9432
rect 6273 9401 6285 9404
rect 6319 9401 6331 9435
rect 6273 9395 6331 9401
rect 6362 9392 6368 9444
rect 6420 9432 6426 9444
rect 6420 9404 6481 9432
rect 6420 9392 6426 9404
rect 7926 9392 7932 9444
rect 7984 9432 7990 9444
rect 8205 9435 8263 9441
rect 8205 9432 8217 9435
rect 7984 9404 8217 9432
rect 7984 9392 7990 9404
rect 8205 9401 8217 9404
rect 8251 9401 8263 9435
rect 8205 9395 8263 9401
rect 7742 9324 7748 9376
rect 7800 9364 7806 9376
rect 7837 9367 7895 9373
rect 7837 9364 7849 9367
rect 7800 9336 7849 9364
rect 7800 9324 7806 9336
rect 7837 9333 7849 9336
rect 7883 9333 7895 9367
rect 7837 9327 7895 9333
rect 8018 9296 8024 9308
rect 7963 9268 8024 9296
rect 8018 9256 8024 9268
rect 8076 9256 8082 9308
rect 6089 9231 6147 9237
rect 6089 9197 6101 9231
rect 6135 9228 6147 9231
rect 6178 9228 6184 9240
rect 6135 9200 6184 9228
rect 6135 9197 6147 9200
rect 6089 9191 6147 9197
rect 6178 9188 6184 9200
rect 6236 9228 6242 9240
rect 6546 9228 6552 9240
rect 6236 9200 6552 9228
rect 6236 9188 6242 9200
rect 6546 9188 6552 9200
rect 6604 9188 6610 9240
rect 7006 9188 7012 9240
rect 7064 9228 7070 9240
rect 7484 9231 7542 9237
rect 7484 9228 7496 9231
rect 7064 9200 7496 9228
rect 7064 9188 7070 9200
rect 7484 9197 7496 9200
rect 7530 9197 7542 9231
rect 7484 9191 7542 9197
rect 7745 9231 7803 9237
rect 7745 9197 7757 9231
rect 7791 9228 7803 9231
rect 8573 9231 8631 9237
rect 8573 9228 8585 9231
rect 7791 9200 8585 9228
rect 7791 9197 7803 9200
rect 7745 9191 7803 9197
rect 8573 9197 8585 9200
rect 8619 9228 8631 9231
rect 8846 9228 8852 9240
rect 8619 9200 8852 9228
rect 8619 9197 8631 9200
rect 8573 9191 8631 9197
rect 8846 9188 8852 9200
rect 8904 9188 8910 9240
rect 9030 9160 9036 9172
rect 8840 9153 8898 9159
rect 8840 9119 8852 9153
rect 8886 9150 8898 9153
rect 8956 9150 9036 9160
rect 8886 9132 9036 9150
rect 8886 9122 8984 9132
rect 8886 9119 8898 9122
rect 9030 9120 9036 9132
rect 9088 9120 9094 9172
rect 8840 9113 8898 9119
rect 5796 9002 10304 9024
rect 5796 8950 8182 9002
rect 8234 8950 8246 9002
rect 8298 8950 8310 9002
rect 8362 8950 8374 9002
rect 8426 8950 8438 9002
rect 8490 8950 8502 9002
rect 8554 8950 8566 9002
rect 8618 8950 8630 9002
rect 8682 8950 8694 9002
rect 8746 8950 8758 9002
rect 8810 8950 10304 9002
rect 5796 8928 10304 8950
rect 14 8848 20 8900
rect 72 8888 78 8900
rect 5997 8891 6055 8897
rect 5997 8888 6009 8891
rect 72 8860 6009 8888
rect 72 8848 78 8860
rect 5997 8857 6009 8860
rect 6043 8857 6055 8891
rect 5997 8851 6055 8857
rect 7929 8860 8156 8888
rect 7929 8829 7957 8860
rect 7914 8823 7972 8829
rect 7914 8789 7926 8823
rect 7960 8789 7972 8823
rect 8128 8820 8156 8860
rect 9030 8848 9036 8900
rect 9088 8888 9094 8900
rect 9125 8891 9183 8897
rect 9125 8888 9137 8891
rect 9088 8860 9137 8888
rect 9088 8848 9094 8860
rect 9125 8857 9137 8860
rect 9171 8857 9183 8891
rect 10137 8891 10195 8897
rect 10137 8888 10149 8891
rect 9125 8851 9183 8857
rect 9968 8860 10149 8888
rect 9968 8854 9996 8860
rect 9232 8826 9996 8854
rect 10137 8857 10149 8860
rect 10183 8857 10195 8891
rect 10137 8851 10195 8857
rect 9232 8820 9260 8826
rect 8128 8792 9260 8820
rect 7914 8783 7972 8789
rect 6089 8755 6147 8761
rect 6089 8721 6101 8755
rect 6135 8752 6147 8755
rect 6178 8752 6184 8764
rect 6135 8724 6184 8752
rect 6135 8721 6147 8724
rect 6089 8715 6147 8721
rect 6178 8712 6184 8724
rect 6236 8712 6242 8764
rect 6454 8752 6460 8764
rect 6399 8724 6460 8752
rect 6454 8712 6460 8724
rect 6512 8712 6518 8764
rect 7650 8752 7656 8764
rect 7595 8724 7656 8752
rect 7650 8712 7656 8724
rect 7708 8712 7714 8764
rect 9401 8755 9459 8761
rect 9401 8752 9413 8755
rect 9048 8724 9413 8752
rect 6730 8684 6736 8696
rect 6675 8656 6736 8684
rect 6730 8644 6736 8656
rect 6788 8644 6794 8696
rect 7377 8687 7435 8693
rect 7377 8653 7389 8687
rect 7423 8653 7435 8687
rect 9048 8684 9076 8724
rect 9401 8721 9413 8724
rect 9447 8752 9459 8755
rect 9953 8755 10011 8761
rect 9953 8752 9965 8755
rect 9447 8724 9965 8752
rect 9447 8721 9459 8724
rect 9401 8715 9459 8721
rect 9953 8721 9965 8724
rect 9999 8721 10011 8755
rect 9953 8715 10011 8721
rect 9766 8684 9772 8696
rect 7377 8647 7435 8653
rect 8956 8656 9076 8684
rect 9711 8656 9772 8684
rect 5626 8576 5632 8628
rect 5684 8616 5690 8628
rect 6914 8616 6920 8628
rect 5684 8588 6920 8616
rect 5684 8576 5690 8588
rect 6914 8576 6920 8588
rect 6972 8616 6978 8628
rect 7392 8616 7420 8647
rect 7558 8616 7564 8628
rect 6972 8588 7420 8616
rect 7503 8588 7564 8616
rect 6972 8576 6978 8588
rect 7006 8508 7012 8560
rect 7064 8548 7070 8560
rect 7193 8551 7251 8557
rect 7193 8548 7205 8551
rect 7064 8520 7205 8548
rect 7064 8508 7070 8520
rect 7193 8517 7205 8520
rect 7239 8517 7251 8551
rect 7392 8548 7420 8588
rect 7558 8576 7564 8588
rect 7616 8576 7622 8628
rect 8018 8548 8024 8560
rect 7392 8520 8024 8548
rect 7193 8511 7251 8517
rect 8018 8508 8024 8520
rect 8076 8548 8082 8560
rect 8956 8548 8984 8656
rect 9766 8644 9772 8656
rect 9824 8644 9830 8696
rect 9582 8616 9588 8628
rect 9527 8588 9588 8616
rect 9582 8576 9588 8588
rect 9640 8576 9646 8628
rect 8076 8520 8984 8548
rect 9033 8551 9091 8557
rect 8076 8508 8082 8520
rect 9033 8517 9045 8551
rect 9079 8548 9091 8551
rect 9122 8548 9128 8560
rect 9079 8520 9128 8548
rect 9079 8517 9091 8520
rect 9033 8511 9091 8517
rect 9122 8508 9128 8520
rect 9180 8508 9186 8560
rect 5796 8458 10304 8480
rect 5796 8406 5800 8458
rect 5852 8406 5864 8458
rect 5916 8406 5928 8458
rect 5980 8406 5992 8458
rect 6044 8406 6056 8458
rect 6108 8406 10304 8458
rect 5796 8384 10304 8406
rect 7377 8347 7435 8353
rect 7377 8313 7389 8347
rect 7423 8344 7435 8347
rect 7558 8344 7564 8356
rect 7423 8316 7564 8344
rect 7423 8313 7435 8316
rect 7377 8307 7435 8313
rect 7558 8304 7564 8316
rect 7616 8304 7622 8356
rect 9490 8304 9496 8356
rect 9548 8344 9554 8356
rect 9953 8347 10011 8353
rect 9953 8344 9965 8347
rect 9548 8316 9965 8344
rect 9548 8304 9554 8316
rect 9953 8313 9965 8316
rect 9999 8313 10011 8347
rect 9953 8307 10011 8313
rect 7285 8211 7343 8217
rect 7285 8177 7297 8211
rect 7331 8208 7343 8211
rect 7650 8208 7656 8220
rect 7331 8180 7656 8208
rect 7331 8177 7343 8180
rect 7285 8171 7343 8177
rect 7650 8168 7656 8180
rect 7708 8168 7714 8220
rect 7006 8140 7012 8152
rect 7064 8149 7070 8152
rect 7064 8143 7082 8149
rect 6963 8112 7012 8140
rect 7006 8100 7012 8112
rect 7070 8109 7082 8143
rect 7561 8143 7619 8149
rect 7561 8140 7573 8143
rect 7064 8103 7082 8109
rect 7116 8112 7573 8140
rect 7064 8100 7070 8103
rect 6362 8032 6368 8084
rect 6420 8072 6426 8084
rect 6420 8044 6500 8072
rect 6420 8032 6426 8044
rect 6472 8004 6500 8044
rect 6730 8032 6736 8084
rect 6788 8072 6794 8084
rect 7116 8072 7144 8112
rect 7561 8109 7573 8112
rect 7607 8109 7619 8143
rect 7834 8140 7840 8152
rect 7779 8112 7840 8140
rect 7561 8103 7619 8109
rect 7834 8100 7840 8112
rect 7892 8100 7898 8152
rect 8018 8100 8024 8152
rect 8076 8140 8082 8152
rect 8481 8143 8539 8149
rect 8481 8140 8493 8143
rect 8076 8112 8493 8140
rect 8076 8100 8082 8112
rect 8481 8109 8493 8112
rect 8527 8109 8539 8143
rect 8481 8103 8539 8109
rect 6788 8044 7144 8072
rect 6788 8032 6794 8044
rect 7650 8032 7656 8084
rect 7708 8072 7714 8084
rect 7745 8075 7803 8081
rect 7745 8072 7757 8075
rect 7708 8044 7757 8072
rect 7708 8032 7714 8044
rect 7745 8041 7757 8044
rect 7791 8072 7803 8075
rect 8113 8075 8171 8081
rect 8113 8072 8125 8075
rect 7791 8044 8125 8072
rect 7791 8041 7803 8044
rect 7745 8035 7803 8041
rect 8113 8041 8125 8044
rect 8159 8041 8171 8075
rect 8113 8035 8171 8041
rect 8742 8075 8800 8081
rect 8742 8041 8754 8075
rect 8788 8072 8800 8075
rect 8846 8072 8852 8084
rect 8788 8044 8852 8072
rect 8788 8041 8800 8044
rect 8742 8035 8800 8041
rect 8846 8032 8852 8044
rect 8904 8032 8910 8084
rect 7929 8007 7987 8013
rect 7929 8004 7941 8007
rect 6472 7976 7941 8004
rect 7929 7973 7941 7976
rect 7975 7973 7987 8007
rect 7929 7967 7987 7973
rect 9861 8007 9919 8013
rect 9861 7973 9873 8007
rect 9907 8004 9919 8007
rect 9907 7976 10364 8004
rect 9907 7973 9919 7976
rect 9861 7967 9919 7973
rect 5796 7914 10304 7936
rect 5796 7862 8182 7914
rect 8234 7862 8246 7914
rect 8298 7862 8310 7914
rect 8362 7862 8374 7914
rect 8426 7862 8438 7914
rect 8490 7862 8502 7914
rect 8554 7862 8566 7914
rect 8618 7862 8630 7914
rect 8682 7862 8694 7914
rect 8746 7862 8758 7914
rect 8810 7862 10304 7914
rect 5796 7840 10304 7862
rect 5905 7803 5963 7809
rect 5905 7769 5917 7803
rect 5951 7800 5963 7803
rect 6273 7803 6331 7809
rect 6273 7800 6285 7803
rect 5951 7772 6285 7800
rect 5951 7769 5963 7772
rect 5905 7763 5963 7769
rect 6273 7769 6285 7772
rect 6319 7769 6331 7803
rect 9122 7800 9128 7812
rect 9067 7772 9128 7800
rect 6273 7763 6331 7769
rect 9122 7760 9128 7772
rect 9180 7800 9186 7812
rect 10336 7800 10364 7976
rect 9180 7772 9720 7800
rect 9180 7760 9186 7772
rect 7454 7744 7512 7750
rect 5629 7735 5687 7741
rect 5629 7701 5641 7735
rect 5675 7701 5687 7735
rect 5629 7695 5687 7701
rect 7009 7735 7067 7741
rect 7009 7701 7021 7735
rect 7055 7732 7067 7735
rect 7454 7732 7466 7744
rect 7055 7710 7466 7732
rect 7500 7710 7512 7744
rect 9582 7732 9588 7744
rect 7055 7704 7512 7710
rect 9527 7704 9588 7732
rect 7055 7701 7067 7704
rect 7009 7695 7067 7701
rect 5644 7664 5672 7695
rect 9582 7692 9588 7704
rect 9640 7692 9646 7744
rect 6181 7667 6239 7673
rect 6181 7664 6193 7667
rect 5644 7636 6193 7664
rect 6181 7633 6193 7636
rect 6227 7633 6239 7667
rect 6181 7627 6239 7633
rect 6638 7624 6644 7676
rect 6696 7664 6702 7676
rect 6825 7667 6883 7673
rect 6825 7664 6837 7667
rect 6696 7636 6837 7664
rect 6696 7624 6702 7636
rect 6825 7633 6837 7636
rect 6871 7633 6883 7667
rect 6825 7627 6883 7633
rect 7193 7667 7251 7673
rect 7193 7633 7205 7667
rect 7239 7664 7251 7667
rect 7466 7664 7472 7676
rect 7239 7636 7472 7664
rect 7239 7633 7251 7636
rect 7193 7627 7251 7633
rect 7466 7624 7472 7636
rect 7524 7624 7530 7676
rect 9401 7667 9459 7673
rect 9401 7633 9413 7667
rect 9447 7664 9459 7667
rect 9490 7664 9496 7676
rect 9447 7636 9496 7664
rect 9447 7633 9459 7636
rect 9401 7627 9459 7633
rect 9490 7624 9496 7636
rect 9548 7624 9554 7676
rect 2685 7599 2743 7605
rect 2685 7565 2697 7599
rect 2731 7596 2743 7599
rect 5997 7599 6055 7605
rect 5997 7596 6009 7599
rect 2731 7568 6009 7596
rect 2731 7565 2743 7568
rect 2685 7559 2743 7565
rect 5997 7565 6009 7568
rect 6043 7565 6055 7599
rect 9692 7596 9720 7772
rect 9876 7772 10364 7800
rect 9769 7667 9827 7673
rect 9769 7633 9781 7667
rect 9815 7664 9827 7667
rect 9876 7664 9904 7772
rect 9815 7636 9904 7664
rect 9953 7667 10011 7673
rect 9815 7633 9827 7636
rect 9769 7627 9827 7633
rect 9953 7633 9965 7667
rect 9999 7633 10011 7667
rect 9953 7627 10011 7633
rect 9968 7596 9996 7627
rect 9692 7568 9996 7596
rect 5997 7559 6055 7565
rect 6457 7531 6515 7537
rect 6457 7497 6469 7531
rect 6503 7528 6515 7531
rect 6503 7500 7236 7528
rect 6503 7497 6515 7500
rect 6457 7491 6515 7497
rect 6549 7463 6607 7469
rect 6549 7460 6561 7463
rect 5736 7432 6561 7460
rect 5736 7256 5764 7432
rect 6549 7429 6561 7432
rect 6595 7429 6607 7463
rect 7208 7460 7236 7500
rect 8573 7463 8631 7469
rect 8573 7460 8585 7463
rect 7208 7432 8585 7460
rect 6549 7423 6607 7429
rect 8573 7429 8585 7432
rect 8619 7429 8631 7463
rect 8573 7423 8631 7429
rect 9030 7420 9036 7472
rect 9088 7460 9094 7472
rect 9769 7463 9827 7469
rect 9769 7460 9781 7463
rect 9088 7432 9781 7460
rect 9088 7420 9094 7432
rect 9769 7429 9781 7432
rect 9815 7429 9827 7463
rect 9769 7423 9827 7429
rect 5796 7370 10304 7392
rect 5796 7318 5800 7370
rect 5852 7318 5864 7370
rect 5916 7318 5928 7370
rect 5980 7318 5992 7370
rect 6044 7318 6056 7370
rect 6108 7318 10304 7370
rect 5796 7296 10304 7318
rect 6089 7259 6147 7265
rect 6089 7256 6101 7259
rect 5736 7228 6101 7256
rect 6089 7225 6101 7228
rect 6135 7225 6147 7259
rect 6089 7219 6147 7225
rect 7834 7216 7840 7268
rect 7892 7256 7898 7268
rect 8297 7259 8355 7265
rect 8297 7256 8309 7259
rect 7892 7228 8309 7256
rect 7892 7216 7898 7228
rect 8297 7225 8309 7228
rect 8343 7225 8355 7259
rect 8297 7219 8355 7225
rect 5442 7080 5448 7132
rect 5500 7120 5506 7132
rect 6638 7120 6644 7132
rect 5500 7092 6644 7120
rect 5500 7080 5506 7092
rect 6638 7080 6644 7092
rect 6696 7080 6702 7132
rect 9858 7120 9864 7132
rect 9803 7092 9864 7120
rect 9858 7080 9864 7092
rect 9916 7080 9922 7132
rect 6089 7055 6147 7061
rect 6089 7021 6101 7055
rect 6135 7021 6147 7055
rect 6089 7015 6147 7021
rect 6104 6984 6132 7015
rect 6178 7012 6184 7064
rect 6236 7052 6242 7064
rect 6236 7024 6297 7052
rect 6236 7012 6242 7024
rect 6362 7012 6368 7064
rect 6420 7012 6426 7064
rect 6917 7055 6975 7061
rect 6917 7021 6929 7055
rect 6963 7052 6975 7055
rect 7466 7052 7472 7064
rect 6963 7024 7472 7052
rect 6963 7021 6975 7024
rect 6917 7015 6975 7021
rect 7466 7012 7472 7024
rect 7524 7012 7530 7064
rect 7650 7012 7656 7064
rect 7708 7052 7714 7064
rect 8389 7055 8447 7061
rect 8389 7052 8401 7055
rect 7708 7024 8401 7052
rect 7708 7012 7714 7024
rect 8389 7021 8401 7024
rect 8435 7021 8447 7055
rect 8389 7015 8447 7021
rect 6380 6984 6408 7012
rect 6104 6956 6408 6984
rect 6825 6987 6883 6993
rect 6825 6953 6837 6987
rect 6871 6984 6883 6987
rect 7178 6987 7236 6993
rect 7178 6984 7190 6987
rect 6871 6956 7190 6984
rect 6871 6953 6883 6956
rect 6825 6947 6883 6953
rect 7178 6953 7190 6956
rect 7224 6953 7236 6987
rect 7178 6947 7236 6953
rect 9600 6987 9658 6993
rect 9600 6953 9612 6987
rect 9646 6984 9658 6987
rect 10413 6987 10471 6993
rect 10413 6984 10425 6987
rect 9646 6956 10425 6984
rect 9646 6953 9658 6956
rect 9600 6947 9658 6953
rect 10413 6953 10425 6956
rect 10459 6953 10471 6987
rect 10413 6947 10471 6953
rect 5796 6826 10304 6848
rect 5796 6774 8182 6826
rect 8234 6774 8246 6826
rect 8298 6774 8310 6826
rect 8362 6774 8374 6826
rect 8426 6774 8438 6826
rect 8490 6774 8502 6826
rect 8554 6774 8566 6826
rect 8618 6774 8630 6826
rect 8682 6774 8694 6826
rect 8746 6774 8758 6826
rect 8810 6774 10304 6826
rect 5796 6752 10304 6774
rect 106 6672 112 6724
rect 164 6712 170 6724
rect 5997 6715 6055 6721
rect 5997 6712 6009 6715
rect 164 6684 6009 6712
rect 164 6672 170 6684
rect 5997 6681 6009 6684
rect 6043 6681 6055 6715
rect 5997 6675 6055 6681
rect 6365 6715 6423 6721
rect 6365 6681 6377 6715
rect 6411 6712 6423 6715
rect 9122 6712 9128 6724
rect 6411 6684 7696 6712
rect 6411 6681 6423 6684
rect 6365 6675 6423 6681
rect 7098 6604 7104 6656
rect 7156 6644 7162 6656
rect 7438 6647 7496 6653
rect 7438 6644 7450 6647
rect 7156 6616 7450 6644
rect 7156 6604 7162 6616
rect 7438 6613 7450 6616
rect 7484 6613 7496 6647
rect 7668 6644 7696 6684
rect 8496 6684 9128 6712
rect 8496 6644 8524 6684
rect 9122 6672 9128 6684
rect 9180 6672 9186 6724
rect 7668 6616 8524 6644
rect 7438 6607 7496 6613
rect 6362 6536 6368 6588
rect 6420 6576 6426 6588
rect 6641 6579 6699 6585
rect 6641 6576 6653 6579
rect 6420 6548 6653 6576
rect 6420 6536 6426 6548
rect 6641 6545 6653 6548
rect 6687 6545 6699 6579
rect 6641 6539 6699 6545
rect 6914 6536 6920 6588
rect 6972 6576 6978 6588
rect 7009 6579 7067 6585
rect 7009 6576 7021 6579
rect 6972 6548 7021 6576
rect 6972 6536 6978 6548
rect 7009 6545 7021 6548
rect 7055 6545 7067 6579
rect 7009 6539 7067 6545
rect 8662 6536 8668 6588
rect 8720 6576 8726 6588
rect 9953 6579 10011 6585
rect 9953 6576 9965 6579
rect 8720 6548 9965 6576
rect 8720 6536 8726 6548
rect 9953 6545 9965 6548
rect 9999 6545 10011 6579
rect 9953 6539 10011 6545
rect 9769 6443 9827 6449
rect 8772 6412 9352 6440
rect 6638 6372 6644 6384
rect 6583 6344 6644 6372
rect 6638 6332 6644 6344
rect 6696 6332 6702 6384
rect 8573 6375 8631 6381
rect 8573 6341 8585 6375
rect 8619 6372 8631 6375
rect 8772 6372 8800 6412
rect 8619 6344 8800 6372
rect 9324 6372 9352 6412
rect 9769 6409 9781 6443
rect 9815 6440 9827 6443
rect 9815 6412 10364 6440
rect 9815 6409 9827 6412
rect 9769 6403 9827 6409
rect 9490 6372 9496 6384
rect 9324 6344 9496 6372
rect 8619 6341 8631 6344
rect 8573 6335 8631 6341
rect 9490 6332 9496 6344
rect 9548 6332 9554 6384
rect 5796 6282 10304 6304
rect 5796 6230 5800 6282
rect 5852 6230 5864 6282
rect 5916 6230 5928 6282
rect 5980 6230 5992 6282
rect 6044 6230 6056 6282
rect 6108 6230 10304 6282
rect 5796 6208 10304 6230
rect 7190 6128 7196 6180
rect 7248 6168 7254 6180
rect 8665 6171 8723 6177
rect 8665 6168 8677 6171
rect 7248 6140 7420 6168
rect 7248 6128 7254 6140
rect 7392 6134 7420 6140
rect 8036 6140 8677 6168
rect 8036 6134 8064 6140
rect 6457 6103 6515 6109
rect 6457 6100 6469 6103
rect 216 6072 6469 6100
rect 216 6044 244 6072
rect 6457 6069 6469 6072
rect 6503 6069 6515 6103
rect 6638 6100 6644 6112
rect 6583 6072 6644 6100
rect 6457 6063 6515 6069
rect 6638 6060 6644 6072
rect 6696 6060 6702 6112
rect 7009 6103 7067 6109
rect 7009 6069 7021 6103
rect 7055 6100 7067 6103
rect 7098 6100 7104 6112
rect 7055 6072 7104 6100
rect 7055 6069 7067 6072
rect 7009 6063 7067 6069
rect 7098 6060 7104 6072
rect 7156 6060 7162 6112
rect 7392 6106 8064 6134
rect 8665 6137 8677 6140
rect 8711 6137 8723 6171
rect 8665 6131 8723 6137
rect 8846 6128 8852 6180
rect 8904 6128 8910 6180
rect 9122 6128 9128 6180
rect 9180 6168 9186 6180
rect 9401 6171 9459 6177
rect 9401 6168 9413 6171
rect 9180 6140 9413 6168
rect 9180 6128 9186 6140
rect 9401 6137 9413 6140
rect 9447 6137 9459 6171
rect 9401 6131 9459 6137
rect 9769 6171 9827 6177
rect 9769 6137 9781 6171
rect 9815 6168 9827 6171
rect 10336 6168 10364 6412
rect 9815 6140 10364 6168
rect 9815 6137 9827 6140
rect 9769 6131 9827 6137
rect 8205 6103 8263 6109
rect 8205 6069 8217 6103
rect 8251 6100 8263 6103
rect 8864 6100 8892 6128
rect 8251 6072 8892 6100
rect 8251 6069 8263 6072
rect 8205 6063 8263 6069
rect 9582 6060 9588 6112
rect 9640 6060 9646 6112
rect 198 5992 204 6044
rect 256 5992 262 6044
rect 6273 6035 6331 6041
rect 6273 6001 6285 6035
rect 6319 6032 6331 6035
rect 7285 6035 7343 6041
rect 7285 6032 7297 6035
rect 6319 6004 7297 6032
rect 6319 6001 6331 6004
rect 6273 5995 6331 6001
rect 7285 6001 7297 6004
rect 7331 6032 7343 6035
rect 8938 6032 8944 6044
rect 7331 6004 8944 6032
rect 7331 6001 7343 6004
rect 7285 5995 7343 6001
rect 8938 5992 8944 6004
rect 8996 5992 9002 6044
rect 9600 6032 9628 6060
rect 9140 6004 9996 6032
rect 6362 5924 6368 5976
rect 6420 5964 6426 5976
rect 6825 5967 6883 5973
rect 6420 5936 6776 5964
rect 6420 5924 6426 5936
rect 6748 5896 6776 5936
rect 6825 5933 6837 5967
rect 6871 5964 6883 5967
rect 7006 5964 7012 5976
rect 6871 5936 7012 5964
rect 6871 5933 6883 5936
rect 6825 5927 6883 5933
rect 7006 5924 7012 5936
rect 7064 5924 7070 5976
rect 7745 5967 7803 5973
rect 7745 5964 7757 5967
rect 7392 5936 7757 5964
rect 7392 5896 7420 5936
rect 7745 5933 7757 5936
rect 7791 5964 7803 5967
rect 7791 5936 7880 5964
rect 7791 5933 7803 5936
rect 7745 5927 7803 5933
rect 6748 5868 7420 5896
rect 7852 5896 7880 5936
rect 8018 5924 8024 5976
rect 8076 5964 8082 5976
rect 8662 5964 8668 5976
rect 8076 5936 8668 5964
rect 8076 5924 8082 5936
rect 8662 5924 8668 5936
rect 8720 5964 8726 5976
rect 9140 5973 9168 6004
rect 8849 5967 8907 5973
rect 8849 5964 8861 5967
rect 8720 5936 8861 5964
rect 8720 5924 8726 5936
rect 8849 5933 8861 5936
rect 8895 5933 8907 5967
rect 9125 5967 9183 5973
rect 9125 5964 9137 5967
rect 8849 5927 8907 5933
rect 8956 5936 9137 5964
rect 8956 5896 8984 5936
rect 9125 5933 9137 5936
rect 9171 5933 9183 5967
rect 9306 5964 9312 5976
rect 9125 5927 9183 5933
rect 9232 5936 9312 5964
rect 7852 5868 8984 5896
rect 14 5788 20 5840
rect 72 5828 78 5840
rect 6089 5831 6147 5837
rect 6089 5828 6101 5831
rect 72 5800 6101 5828
rect 72 5788 78 5800
rect 6089 5797 6101 5800
rect 6135 5797 6147 5831
rect 6089 5791 6147 5797
rect 6549 5831 6607 5837
rect 6549 5797 6561 5831
rect 6595 5828 6607 5831
rect 9232 5828 9260 5936
rect 9306 5924 9312 5936
rect 9364 5924 9370 5976
rect 9401 5967 9459 5973
rect 9401 5933 9413 5967
rect 9447 5964 9459 5967
rect 9490 5964 9496 5976
rect 9447 5936 9496 5964
rect 9447 5933 9459 5936
rect 9401 5927 9459 5933
rect 9490 5924 9496 5936
rect 9548 5924 9554 5976
rect 9968 5973 9996 6004
rect 9585 5967 9643 5973
rect 9585 5933 9597 5967
rect 9631 5964 9643 5967
rect 9953 5967 10011 5973
rect 9631 5936 9904 5964
rect 9631 5933 9643 5936
rect 9585 5927 9643 5933
rect 9876 5896 9904 5936
rect 9953 5933 9965 5967
rect 9999 5933 10011 5967
rect 9953 5927 10011 5933
rect 10137 5899 10195 5905
rect 10137 5896 10149 5899
rect 9876 5868 10149 5896
rect 10137 5865 10149 5868
rect 10183 5865 10195 5899
rect 10137 5859 10195 5865
rect 6595 5800 9260 5828
rect 6595 5797 6607 5800
rect 6549 5791 6607 5797
rect 5796 5738 10304 5760
rect 5796 5686 8182 5738
rect 8234 5686 8246 5738
rect 8298 5686 8310 5738
rect 8362 5686 8374 5738
rect 8426 5686 8438 5738
rect 8490 5686 8502 5738
rect 8554 5686 8566 5738
rect 8618 5686 8630 5738
rect 8682 5686 8694 5738
rect 8746 5686 8758 5738
rect 8810 5686 10304 5738
rect 5796 5664 10304 5686
rect 14 76 20 128
rect 72 116 78 128
rect 1397 119 1455 125
rect 1397 116 1409 119
rect 72 88 1409 116
rect 72 76 78 88
rect 1397 85 1409 88
rect 1443 85 1455 119
rect 1397 79 1455 85
<< via1 >>
rect 20 17892 72 17944
rect 20 17076 72 17128
rect 8182 14390 8234 14442
rect 8246 14390 8298 14442
rect 8310 14390 8362 14442
rect 8374 14390 8426 14442
rect 8438 14390 8490 14442
rect 8502 14390 8554 14442
rect 8566 14390 8618 14442
rect 8630 14390 8682 14442
rect 8694 14390 8746 14442
rect 8758 14390 8810 14442
rect 8852 14288 8904 14340
rect 6644 14195 6696 14204
rect 6644 14161 6653 14195
rect 6653 14161 6687 14195
rect 6687 14161 6696 14195
rect 6644 14152 6696 14161
rect 7564 14152 7616 14204
rect 8392 14220 8444 14272
rect 10324 14220 10376 14272
rect 7840 14084 7892 14136
rect 8208 14152 8260 14204
rect 9864 14152 9916 14204
rect 15844 14152 15896 14204
rect 8208 13948 8260 14000
rect 8668 13948 8720 14000
rect 9312 13991 9364 14000
rect 9312 13957 9321 13991
rect 9321 13957 9355 13991
rect 9355 13957 9364 13991
rect 9312 13948 9364 13957
rect 10140 13948 10192 14000
rect 5800 13846 5852 13898
rect 5864 13846 5916 13898
rect 5928 13846 5980 13898
rect 5992 13846 6044 13898
rect 6056 13846 6108 13898
rect 20 13744 72 13796
rect 8668 13744 8720 13796
rect 9496 13744 9548 13796
rect 16028 13744 16080 13796
rect 6828 13676 6880 13728
rect 8208 13540 8260 13592
rect 8852 13540 8904 13592
rect 8392 13472 8444 13524
rect 9220 13472 9272 13524
rect 7012 13404 7064 13456
rect 8182 13302 8234 13354
rect 8246 13302 8298 13354
rect 8310 13302 8362 13354
rect 8374 13302 8426 13354
rect 8438 13302 8490 13354
rect 8502 13302 8554 13354
rect 8566 13302 8618 13354
rect 8630 13302 8682 13354
rect 8694 13302 8746 13354
rect 8758 13302 8810 13354
rect 20 13200 72 13252
rect 9220 13243 9272 13252
rect 9220 13209 9229 13243
rect 9229 13209 9263 13243
rect 9263 13209 9272 13243
rect 9220 13200 9272 13209
rect 6644 13064 6696 13116
rect 6828 13064 6880 13116
rect 8024 13064 8076 13116
rect 8852 12996 8904 13048
rect 9312 13064 9364 13116
rect 9496 13064 9548 13116
rect 9864 13064 9916 13116
rect 9220 12996 9272 13048
rect 10324 12928 10376 12980
rect 6644 12860 6696 12912
rect 5800 12758 5852 12810
rect 5864 12758 5916 12810
rect 5928 12758 5980 12810
rect 5992 12758 6044 12810
rect 6056 12758 6108 12810
rect 6920 12656 6972 12708
rect 7564 12520 7616 12572
rect 6736 12452 6788 12504
rect 6644 12384 6696 12436
rect 7840 12520 7892 12572
rect 8852 12452 8904 12504
rect 7472 12427 7524 12436
rect 7472 12393 7481 12427
rect 7481 12393 7515 12427
rect 7515 12393 7524 12427
rect 7472 12384 7524 12393
rect 7748 12384 7800 12436
rect 8182 12214 8234 12266
rect 8246 12214 8298 12266
rect 8310 12214 8362 12266
rect 8374 12214 8426 12266
rect 8438 12214 8490 12266
rect 8502 12214 8554 12266
rect 8566 12214 8618 12266
rect 8630 12214 8682 12266
rect 8694 12214 8746 12266
rect 8758 12214 8810 12266
rect 7012 12112 7064 12164
rect 7472 12155 7524 12164
rect 7472 12121 7481 12155
rect 7481 12121 7515 12155
rect 7515 12121 7524 12155
rect 7472 12112 7524 12121
rect 6184 11976 6236 12028
rect 6644 11976 6696 12028
rect 6552 11951 6604 11960
rect 6552 11917 6561 11951
rect 6561 11917 6595 11951
rect 6595 11917 6604 11951
rect 6552 11908 6604 11917
rect 9220 11976 9272 12028
rect 7564 11908 7616 11960
rect 10324 11840 10376 11892
rect 5800 11670 5852 11722
rect 5864 11670 5916 11722
rect 5928 11670 5980 11722
rect 5992 11670 6044 11722
rect 6056 11670 6108 11722
rect 7656 11568 7708 11620
rect 9864 11568 9916 11620
rect 6092 11364 6144 11416
rect 7564 11364 7616 11416
rect 8024 11364 8076 11416
rect 8760 11364 8812 11416
rect 6368 11339 6420 11348
rect 6368 11305 6377 11339
rect 6377 11305 6411 11339
rect 6411 11305 6420 11339
rect 6368 11296 6420 11305
rect 7288 11228 7340 11280
rect 9956 11228 10008 11280
rect 8182 11126 8234 11178
rect 8246 11126 8298 11178
rect 8310 11126 8362 11178
rect 8374 11126 8426 11178
rect 8438 11126 8490 11178
rect 8502 11126 8554 11178
rect 8566 11126 8618 11178
rect 8630 11126 8682 11178
rect 8694 11126 8746 11178
rect 8758 11126 8810 11178
rect 6092 10931 6144 10940
rect 6092 10897 6101 10931
rect 6101 10897 6135 10931
rect 6135 10897 6144 10931
rect 6092 10888 6144 10897
rect 7288 11024 7340 11076
rect 6368 10931 6420 10940
rect 6368 10897 6377 10931
rect 6377 10897 6411 10931
rect 6411 10897 6420 10931
rect 6368 10888 6420 10897
rect 6552 10888 6604 10940
rect 7840 11024 7892 11076
rect 10324 11024 10376 11076
rect 7656 10888 7708 10940
rect 9496 10888 9548 10940
rect 9588 10888 9640 10940
rect 10140 10863 10192 10872
rect 10140 10829 10149 10863
rect 10149 10829 10183 10863
rect 10183 10829 10192 10863
rect 10140 10820 10192 10829
rect 7472 10795 7524 10804
rect 7472 10761 7481 10795
rect 7481 10761 7515 10795
rect 7515 10761 7524 10795
rect 7472 10752 7524 10761
rect 9036 10752 9088 10804
rect 5800 10582 5852 10634
rect 5864 10582 5916 10634
rect 5928 10582 5980 10634
rect 5992 10582 6044 10634
rect 6056 10582 6108 10634
rect 6552 10344 6604 10396
rect 6184 10319 6236 10328
rect 6184 10285 6193 10319
rect 6193 10285 6227 10319
rect 6227 10285 6236 10319
rect 6184 10276 6236 10285
rect 7472 10276 7524 10328
rect 8760 10276 8812 10328
rect 7196 10251 7248 10260
rect 7196 10217 7224 10251
rect 7224 10217 7248 10251
rect 7196 10208 7248 10217
rect 7932 10208 7984 10260
rect 7012 10140 7064 10192
rect 8300 10183 8352 10192
rect 8300 10149 8309 10183
rect 8309 10149 8343 10183
rect 8343 10149 8352 10183
rect 8300 10140 8352 10149
rect 9864 10183 9916 10192
rect 9864 10149 9873 10183
rect 9873 10149 9907 10183
rect 9907 10149 9916 10183
rect 9864 10140 9916 10149
rect 9956 10183 10008 10192
rect 9956 10149 9965 10183
rect 9965 10149 9999 10183
rect 9999 10149 10008 10183
rect 9956 10140 10008 10149
rect 20 10072 72 10124
rect 8182 10038 8234 10090
rect 8246 10038 8298 10090
rect 8310 10038 8362 10090
rect 8374 10038 8426 10090
rect 8438 10038 8490 10090
rect 8502 10038 8554 10090
rect 8566 10038 8618 10090
rect 8630 10038 8682 10090
rect 8694 10038 8746 10090
rect 8758 10038 8810 10090
rect 7012 9868 7064 9920
rect 9864 9868 9916 9920
rect 6460 9843 6512 9852
rect 6460 9809 6469 9843
rect 6469 9809 6503 9843
rect 6503 9809 6512 9843
rect 6460 9800 6512 9809
rect 6552 9800 6604 9852
rect 7472 9800 7524 9852
rect 9404 9843 9456 9852
rect 9404 9809 9413 9843
rect 9413 9809 9447 9843
rect 9447 9809 9456 9843
rect 9404 9800 9456 9809
rect 9956 9843 10008 9852
rect 9956 9809 9965 9843
rect 9965 9809 9999 9843
rect 9999 9809 10008 9843
rect 9956 9800 10008 9809
rect 6460 9707 6512 9716
rect 6460 9673 6469 9707
rect 6469 9673 6503 9707
rect 6503 9673 6512 9707
rect 6460 9664 6512 9673
rect 7012 9639 7064 9648
rect 7012 9605 7021 9639
rect 7021 9605 7055 9639
rect 7055 9605 7064 9639
rect 7012 9596 7064 9605
rect 9312 9596 9364 9648
rect 9772 9639 9824 9648
rect 9772 9605 9781 9639
rect 9781 9605 9815 9639
rect 9815 9605 9824 9639
rect 9772 9596 9824 9605
rect 5800 9494 5852 9546
rect 5864 9494 5916 9546
rect 5928 9494 5980 9546
rect 5992 9494 6044 9546
rect 6056 9494 6108 9546
rect 6368 9435 6420 9444
rect 6368 9401 6377 9435
rect 6377 9401 6411 9435
rect 6411 9401 6420 9435
rect 6368 9392 6420 9401
rect 7932 9392 7984 9444
rect 7748 9324 7800 9376
rect 8024 9299 8076 9308
rect 8024 9265 8033 9299
rect 8033 9265 8067 9299
rect 8067 9265 8076 9299
rect 8024 9256 8076 9265
rect 6184 9188 6236 9240
rect 6552 9188 6604 9240
rect 7012 9188 7064 9240
rect 8852 9188 8904 9240
rect 9036 9120 9088 9172
rect 8182 8950 8234 9002
rect 8246 8950 8298 9002
rect 8310 8950 8362 9002
rect 8374 8950 8426 9002
rect 8438 8950 8490 9002
rect 8502 8950 8554 9002
rect 8566 8950 8618 9002
rect 8630 8950 8682 9002
rect 8694 8950 8746 9002
rect 8758 8950 8810 9002
rect 20 8848 72 8900
rect 9036 8848 9088 8900
rect 6184 8712 6236 8764
rect 6460 8755 6512 8764
rect 6460 8721 6469 8755
rect 6469 8721 6503 8755
rect 6503 8721 6512 8755
rect 6460 8712 6512 8721
rect 7656 8755 7708 8764
rect 7656 8721 7665 8755
rect 7665 8721 7699 8755
rect 7699 8721 7708 8755
rect 7656 8712 7708 8721
rect 6736 8687 6788 8696
rect 6736 8653 6745 8687
rect 6745 8653 6779 8687
rect 6779 8653 6788 8687
rect 6736 8644 6788 8653
rect 9772 8687 9824 8696
rect 5632 8576 5684 8628
rect 6920 8576 6972 8628
rect 7564 8619 7616 8628
rect 7012 8508 7064 8560
rect 7564 8585 7573 8619
rect 7573 8585 7607 8619
rect 7607 8585 7616 8619
rect 7564 8576 7616 8585
rect 8024 8508 8076 8560
rect 9772 8653 9781 8687
rect 9781 8653 9815 8687
rect 9815 8653 9824 8687
rect 9772 8644 9824 8653
rect 9588 8619 9640 8628
rect 9588 8585 9597 8619
rect 9597 8585 9631 8619
rect 9631 8585 9640 8619
rect 9588 8576 9640 8585
rect 9128 8508 9180 8560
rect 5800 8406 5852 8458
rect 5864 8406 5916 8458
rect 5928 8406 5980 8458
rect 5992 8406 6044 8458
rect 6056 8406 6108 8458
rect 7564 8304 7616 8356
rect 9496 8304 9548 8356
rect 7656 8168 7708 8220
rect 7012 8143 7064 8152
rect 7012 8109 7036 8143
rect 7036 8109 7064 8143
rect 7012 8100 7064 8109
rect 6368 8032 6420 8084
rect 6736 8032 6788 8084
rect 7840 8143 7892 8152
rect 7840 8109 7849 8143
rect 7849 8109 7883 8143
rect 7883 8109 7892 8143
rect 7840 8100 7892 8109
rect 8024 8100 8076 8152
rect 7656 8032 7708 8084
rect 8852 8032 8904 8084
rect 8182 7862 8234 7914
rect 8246 7862 8298 7914
rect 8310 7862 8362 7914
rect 8374 7862 8426 7914
rect 8438 7862 8490 7914
rect 8502 7862 8554 7914
rect 8566 7862 8618 7914
rect 8630 7862 8682 7914
rect 8694 7862 8746 7914
rect 8758 7862 8810 7914
rect 9128 7803 9180 7812
rect 9128 7769 9137 7803
rect 9137 7769 9171 7803
rect 9171 7769 9180 7803
rect 9128 7760 9180 7769
rect 9588 7735 9640 7744
rect 9588 7701 9597 7735
rect 9597 7701 9631 7735
rect 9631 7701 9640 7735
rect 9588 7692 9640 7701
rect 6644 7624 6696 7676
rect 7472 7624 7524 7676
rect 9496 7624 9548 7676
rect 9036 7420 9088 7472
rect 5800 7318 5852 7370
rect 5864 7318 5916 7370
rect 5928 7318 5980 7370
rect 5992 7318 6044 7370
rect 6056 7318 6108 7370
rect 7840 7216 7892 7268
rect 5448 7080 5500 7132
rect 6644 7123 6696 7132
rect 6644 7089 6653 7123
rect 6653 7089 6687 7123
rect 6687 7089 6696 7123
rect 6644 7080 6696 7089
rect 9864 7123 9916 7132
rect 9864 7089 9873 7123
rect 9873 7089 9907 7123
rect 9907 7089 9916 7123
rect 9864 7080 9916 7089
rect 6184 7055 6236 7064
rect 6184 7021 6193 7055
rect 6193 7021 6227 7055
rect 6227 7021 6236 7055
rect 6184 7012 6236 7021
rect 6368 7055 6420 7064
rect 6368 7021 6377 7055
rect 6377 7021 6411 7055
rect 6411 7021 6420 7055
rect 6368 7012 6420 7021
rect 7472 7012 7524 7064
rect 7656 7012 7708 7064
rect 8182 6774 8234 6826
rect 8246 6774 8298 6826
rect 8310 6774 8362 6826
rect 8374 6774 8426 6826
rect 8438 6774 8490 6826
rect 8502 6774 8554 6826
rect 8566 6774 8618 6826
rect 8630 6774 8682 6826
rect 8694 6774 8746 6826
rect 8758 6774 8810 6826
rect 112 6672 164 6724
rect 7104 6604 7156 6656
rect 9128 6672 9180 6724
rect 6368 6536 6420 6588
rect 6920 6536 6972 6588
rect 8668 6536 8720 6588
rect 6644 6375 6696 6384
rect 6644 6341 6653 6375
rect 6653 6341 6687 6375
rect 6687 6341 6696 6375
rect 6644 6332 6696 6341
rect 9496 6332 9548 6384
rect 5800 6230 5852 6282
rect 5864 6230 5916 6282
rect 5928 6230 5980 6282
rect 5992 6230 6044 6282
rect 6056 6230 6108 6282
rect 7196 6128 7248 6180
rect 6644 6103 6696 6112
rect 6644 6069 6653 6103
rect 6653 6069 6687 6103
rect 6687 6069 6696 6103
rect 6644 6060 6696 6069
rect 7104 6060 7156 6112
rect 8852 6128 8904 6180
rect 9128 6128 9180 6180
rect 9588 6060 9640 6112
rect 204 5992 256 6044
rect 8944 5992 8996 6044
rect 6368 5924 6420 5976
rect 7012 5924 7064 5976
rect 8024 5967 8076 5976
rect 8024 5933 8033 5967
rect 8033 5933 8067 5967
rect 8067 5933 8076 5967
rect 8024 5924 8076 5933
rect 8668 5924 8720 5976
rect 9312 5967 9364 5976
rect 20 5788 72 5840
rect 9312 5933 9321 5967
rect 9321 5933 9355 5967
rect 9355 5933 9364 5967
rect 9312 5924 9364 5933
rect 9496 5924 9548 5976
rect 8182 5686 8234 5738
rect 8246 5686 8298 5738
rect 8310 5686 8362 5738
rect 8374 5686 8426 5738
rect 8438 5686 8490 5738
rect 8502 5686 8554 5738
rect 8566 5686 8618 5738
rect 8630 5686 8682 5738
rect 8694 5686 8746 5738
rect 8758 5686 8810 5738
rect 20 76 72 128
<< metal2 >>
rect 0 20080 97 20108
rect 32 17944 60 20080
rect 14 17892 20 17944
rect 72 17892 78 17944
rect 0 17836 97 17864
rect 32 17134 60 17836
rect 20 17128 72 17134
rect 20 17070 72 17076
rect 0 15592 97 15620
rect 32 13802 60 15592
rect 216 14933 244 20128
rect 202 14924 258 14933
rect 202 14859 258 14868
rect 6458 14924 6514 14933
rect 6458 14859 6514 14868
rect 5796 13900 6112 13920
rect 5796 13898 5806 13900
rect 5862 13898 5886 13900
rect 5942 13898 5966 13900
rect 6022 13898 6046 13900
rect 6102 13898 6112 13900
rect 5796 13846 5800 13898
rect 5862 13846 5864 13898
rect 6044 13846 6046 13898
rect 6108 13846 6112 13898
rect 5796 13844 5806 13846
rect 5862 13844 5886 13846
rect 5942 13844 5966 13846
rect 6022 13844 6046 13846
rect 6102 13844 6112 13846
rect 5796 13824 6112 13844
rect 20 13796 72 13802
rect 20 13738 72 13744
rect 0 13348 97 13376
rect 32 13258 60 13348
rect 20 13252 72 13258
rect 20 13194 72 13200
rect 5796 12812 6112 12832
rect 5796 12810 5806 12812
rect 5862 12810 5886 12812
rect 5942 12810 5966 12812
rect 6022 12810 6046 12812
rect 6102 12810 6112 12812
rect 5796 12758 5800 12810
rect 5862 12758 5864 12810
rect 6044 12758 6046 12810
rect 6108 12758 6112 12810
rect 5796 12756 5806 12758
rect 5862 12756 5886 12758
rect 5942 12756 5966 12758
rect 6022 12756 6046 12758
rect 6102 12756 6112 12758
rect 5796 12736 6112 12756
rect 6184 12028 6236 12034
rect 6184 11970 6236 11976
rect 5796 11724 6112 11744
rect 5796 11722 5806 11724
rect 5862 11722 5886 11724
rect 5942 11722 5966 11724
rect 6022 11722 6046 11724
rect 6102 11722 6112 11724
rect 5796 11670 5800 11722
rect 5862 11670 5864 11722
rect 6044 11670 6046 11722
rect 6108 11670 6112 11722
rect 5796 11668 5806 11670
rect 5862 11668 5886 11670
rect 5942 11668 5966 11670
rect 6022 11668 6046 11670
rect 6102 11668 6112 11670
rect 5796 11648 6112 11668
rect 6196 11608 6224 11970
rect 6104 11580 6224 11608
rect 6104 11422 6132 11580
rect 6092 11416 6144 11422
rect 6092 11358 6144 11364
rect 0 11104 97 11132
rect 32 10130 60 11104
rect 6104 10946 6132 11358
rect 6368 11348 6420 11354
rect 6368 11290 6420 11296
rect 6380 10946 6408 11290
rect 6092 10940 6144 10946
rect 6368 10940 6420 10946
rect 6092 10882 6144 10888
rect 6288 10900 6368 10928
rect 6104 10792 6132 10882
rect 6104 10764 6224 10792
rect 5796 10636 6112 10656
rect 5796 10634 5806 10636
rect 5862 10634 5886 10636
rect 5942 10634 5966 10636
rect 6022 10634 6046 10636
rect 6102 10634 6112 10636
rect 5796 10582 5800 10634
rect 5862 10582 5864 10634
rect 6044 10582 6046 10634
rect 6108 10582 6112 10634
rect 5796 10580 5806 10582
rect 5862 10580 5886 10582
rect 5942 10580 5966 10582
rect 6022 10580 6046 10582
rect 6102 10580 6112 10582
rect 5796 10560 6112 10580
rect 6196 10334 6224 10764
rect 6184 10328 6236 10334
rect 6184 10270 6236 10276
rect 20 10124 72 10130
rect 20 10066 72 10072
rect 5796 9548 6112 9568
rect 5796 9546 5806 9548
rect 5862 9546 5886 9548
rect 5942 9546 5966 9548
rect 6022 9546 6046 9548
rect 6102 9546 6112 9548
rect 5796 9494 5800 9546
rect 5862 9494 5864 9546
rect 6044 9494 6046 9546
rect 6108 9494 6112 9546
rect 5796 9492 5806 9494
rect 5862 9492 5886 9494
rect 5942 9492 5966 9494
rect 6022 9492 6046 9494
rect 6102 9492 6112 9494
rect 5796 9472 6112 9492
rect 6196 9246 6224 10270
rect 6288 9432 6316 10900
rect 6368 10882 6420 10888
rect 6472 10785 6500 14859
rect 6644 14204 6696 14210
rect 6644 14146 6696 14152
rect 7564 14204 7616 14210
rect 8036 14192 8064 20128
rect 15856 19904 15884 20128
rect 16003 20080 16100 20108
rect 15764 19876 15884 19904
rect 8160 14444 8832 14464
rect 8160 14442 8188 14444
rect 8244 14442 8268 14444
rect 8324 14442 8348 14444
rect 8404 14442 8428 14444
rect 8484 14442 8508 14444
rect 8564 14442 8588 14444
rect 8644 14442 8668 14444
rect 8724 14442 8748 14444
rect 8804 14442 8832 14444
rect 8160 14390 8182 14442
rect 8244 14390 8246 14442
rect 8426 14390 8428 14442
rect 8490 14390 8502 14442
rect 8564 14390 8566 14442
rect 8746 14390 8748 14442
rect 8810 14390 8832 14442
rect 8160 14388 8188 14390
rect 8244 14388 8268 14390
rect 8324 14388 8348 14390
rect 8404 14388 8428 14390
rect 8484 14388 8508 14390
rect 8564 14388 8588 14390
rect 8644 14388 8668 14390
rect 8724 14388 8748 14390
rect 8804 14388 8832 14390
rect 8160 14368 8832 14388
rect 15764 14396 15792 19876
rect 15764 14368 15884 14396
rect 8852 14340 8904 14346
rect 8852 14282 8904 14288
rect 8392 14272 8444 14278
rect 8392 14214 8444 14220
rect 8208 14204 8260 14210
rect 7564 14146 7616 14152
rect 7944 14164 8208 14192
rect 6656 13122 6684 14146
rect 6828 13728 6880 13734
rect 6828 13670 6880 13676
rect 6840 13122 6868 13670
rect 7012 13456 7064 13462
rect 7012 13398 7064 13404
rect 7024 13240 7052 13398
rect 7024 13212 7144 13240
rect 6644 13116 6696 13122
rect 6644 13058 6696 13064
rect 6828 13116 6880 13122
rect 6828 13058 6880 13064
rect 6644 12912 6696 12918
rect 6644 12854 6696 12860
rect 6656 12442 6684 12854
rect 6840 12696 6868 13058
rect 6920 12708 6972 12714
rect 6840 12668 6920 12696
rect 6920 12650 6972 12656
rect 7116 12560 7144 13212
rect 7576 12578 7604 14146
rect 7840 14136 7892 14142
rect 7944 14124 7972 14164
rect 8208 14146 8260 14152
rect 7892 14096 7972 14124
rect 7840 14078 7892 14084
rect 7944 13104 7972 14096
rect 8208 14000 8260 14006
rect 8208 13942 8260 13948
rect 8220 13598 8248 13942
rect 8208 13592 8260 13598
rect 8208 13534 8260 13540
rect 8404 13530 8432 14214
rect 8668 14000 8720 14006
rect 8668 13942 8720 13948
rect 8680 13802 8708 13942
rect 8668 13796 8720 13802
rect 8864 13784 8892 14282
rect 10324 14272 10376 14278
rect 10324 14214 10376 14220
rect 9864 14204 9916 14210
rect 9864 14146 9916 14152
rect 9312 14000 9364 14006
rect 9312 13942 9364 13948
rect 8864 13756 9076 13784
rect 8668 13738 8720 13744
rect 8852 13592 8904 13598
rect 8852 13534 8904 13540
rect 8392 13524 8444 13530
rect 8392 13466 8444 13472
rect 8160 13356 8832 13376
rect 8160 13354 8188 13356
rect 8244 13354 8268 13356
rect 8324 13354 8348 13356
rect 8404 13354 8428 13356
rect 8484 13354 8508 13356
rect 8564 13354 8588 13356
rect 8644 13354 8668 13356
rect 8724 13354 8748 13356
rect 8804 13354 8832 13356
rect 8160 13302 8182 13354
rect 8244 13302 8246 13354
rect 8426 13302 8428 13354
rect 8490 13302 8502 13354
rect 8564 13302 8566 13354
rect 8746 13302 8748 13354
rect 8810 13302 8832 13354
rect 8160 13300 8188 13302
rect 8244 13300 8268 13302
rect 8324 13300 8348 13302
rect 8404 13300 8428 13302
rect 8484 13300 8508 13302
rect 8564 13300 8588 13302
rect 8644 13300 8668 13302
rect 8724 13300 8748 13302
rect 8804 13300 8832 13302
rect 8160 13280 8832 13300
rect 8024 13116 8076 13122
rect 7944 13076 8024 13104
rect 8024 13058 8076 13064
rect 7024 12532 7144 12560
rect 7564 12572 7616 12578
rect 6736 12504 6788 12510
rect 6736 12446 6788 12452
rect 6644 12436 6696 12442
rect 6644 12378 6696 12384
rect 6656 12034 6684 12378
rect 6644 12028 6696 12034
rect 6644 11970 6696 11976
rect 6552 11960 6604 11966
rect 6552 11902 6604 11908
rect 6564 10946 6592 11902
rect 6552 10940 6604 10946
rect 6552 10882 6604 10888
rect 6458 10776 6514 10785
rect 6458 10711 6514 10720
rect 6472 9858 6500 10711
rect 6564 10402 6592 10882
rect 6552 10396 6604 10402
rect 6552 10338 6604 10344
rect 6564 9858 6592 10338
rect 6460 9852 6512 9858
rect 6460 9794 6512 9800
rect 6552 9852 6604 9858
rect 6552 9794 6604 9800
rect 6460 9716 6512 9722
rect 6460 9658 6512 9664
rect 6368 9444 6420 9450
rect 6288 9404 6368 9432
rect 6368 9386 6420 9392
rect 6184 9240 6236 9246
rect 6184 9182 6236 9188
rect 0 8928 97 8956
rect 32 8900 60 8928
rect 14 8848 20 8900
rect 72 8848 78 8900
rect 6472 8770 6500 9658
rect 6552 9240 6604 9246
rect 6552 9182 6604 9188
rect 6184 8764 6236 8770
rect 6184 8706 6236 8712
rect 6460 8764 6512 8770
rect 6460 8706 6512 8712
rect 5632 8628 5684 8634
rect 5460 8588 5632 8616
rect 5460 7138 5488 8588
rect 5632 8570 5684 8576
rect 5796 8460 6112 8480
rect 5796 8458 5806 8460
rect 5862 8458 5886 8460
rect 5942 8458 5966 8460
rect 6022 8458 6046 8460
rect 6102 8458 6112 8460
rect 5796 8406 5800 8458
rect 5862 8406 5864 8458
rect 6044 8406 6046 8458
rect 6108 8406 6112 8458
rect 5796 8404 5806 8406
rect 5862 8404 5886 8406
rect 5942 8404 5966 8406
rect 6022 8404 6046 8406
rect 6102 8404 6112 8406
rect 5796 8384 6112 8404
rect 6196 8072 6224 8706
rect 6368 8084 6420 8090
rect 6196 8044 6368 8072
rect 5796 7372 6112 7392
rect 5796 7370 5806 7372
rect 5862 7370 5886 7372
rect 5942 7370 5966 7372
rect 6022 7370 6046 7372
rect 6102 7370 6112 7372
rect 5796 7318 5800 7370
rect 5862 7318 5864 7370
rect 6044 7318 6046 7370
rect 6108 7318 6112 7370
rect 5796 7316 5806 7318
rect 5862 7316 5886 7318
rect 5942 7316 5966 7318
rect 6022 7316 6046 7318
rect 6102 7316 6112 7318
rect 5796 7296 6112 7316
rect 5448 7132 5500 7138
rect 5448 7074 5500 7080
rect 6196 7070 6224 8044
rect 6368 8026 6420 8032
rect 6564 8072 6592 9182
rect 6748 8833 6776 12446
rect 7024 12170 7052 12532
rect 7564 12514 7616 12520
rect 7840 12572 7892 12578
rect 7840 12514 7892 12520
rect 7472 12436 7524 12442
rect 7472 12378 7524 12384
rect 7748 12436 7800 12442
rect 7748 12378 7800 12384
rect 7484 12170 7512 12378
rect 7012 12164 7064 12170
rect 7012 12106 7064 12112
rect 7472 12164 7524 12170
rect 7472 12106 7524 12112
rect 7564 11960 7616 11966
rect 7564 11902 7616 11908
rect 7576 11422 7604 11902
rect 7656 11620 7708 11626
rect 7760 11608 7788 12378
rect 7852 12356 7880 12514
rect 7852 12328 7926 12356
rect 7898 11608 7926 12328
rect 8036 12084 8064 13058
rect 8864 13054 8892 13534
rect 8852 13048 8904 13054
rect 8852 12990 8904 12996
rect 8864 12510 8892 12990
rect 8852 12504 8904 12510
rect 8852 12446 8904 12452
rect 8160 12268 8832 12288
rect 8160 12266 8188 12268
rect 8244 12266 8268 12268
rect 8324 12266 8348 12268
rect 8404 12266 8428 12268
rect 8484 12266 8508 12268
rect 8564 12266 8588 12268
rect 8644 12266 8668 12268
rect 8724 12266 8748 12268
rect 8804 12266 8832 12268
rect 8160 12214 8182 12266
rect 8244 12214 8246 12266
rect 8426 12214 8428 12266
rect 8490 12214 8502 12266
rect 8564 12214 8566 12266
rect 8746 12214 8748 12266
rect 8810 12214 8832 12266
rect 8160 12212 8188 12214
rect 8244 12212 8268 12214
rect 8324 12212 8348 12214
rect 8404 12212 8428 12214
rect 8484 12212 8508 12214
rect 8564 12212 8588 12214
rect 8644 12212 8668 12214
rect 8724 12212 8748 12214
rect 8804 12212 8832 12214
rect 8160 12192 8832 12212
rect 8036 12056 8156 12084
rect 8128 11608 8156 12056
rect 7708 11580 7788 11608
rect 7852 11580 7926 11608
rect 8036 11580 8156 11608
rect 7656 11562 7708 11568
rect 7852 11472 7880 11580
rect 7760 11444 7880 11472
rect 7564 11416 7616 11422
rect 7484 11376 7564 11404
rect 7288 11280 7340 11286
rect 7288 11222 7340 11228
rect 7300 11082 7328 11222
rect 7288 11076 7340 11082
rect 7288 11018 7340 11024
rect 7484 10810 7512 11376
rect 7564 11358 7616 11364
rect 7656 10940 7708 10946
rect 7656 10882 7708 10888
rect 7472 10804 7524 10810
rect 7668 10785 7696 10882
rect 7472 10746 7524 10752
rect 7654 10776 7710 10785
rect 7484 10334 7512 10746
rect 7654 10711 7710 10720
rect 7472 10328 7524 10334
rect 7472 10270 7524 10276
rect 7196 10260 7248 10266
rect 7196 10202 7248 10208
rect 7012 10192 7064 10198
rect 7012 10134 7064 10140
rect 7024 9926 7052 10134
rect 7012 9920 7064 9926
rect 7012 9862 7064 9868
rect 7012 9648 7064 9654
rect 7012 9590 7064 9596
rect 7024 9246 7052 9590
rect 7012 9240 7064 9246
rect 7012 9182 7064 9188
rect 6734 8824 6790 8833
rect 6734 8759 6790 8768
rect 6748 8702 6776 8759
rect 6736 8696 6788 8702
rect 6736 8638 6788 8644
rect 6920 8628 6972 8634
rect 6920 8570 6972 8576
rect 6736 8084 6788 8090
rect 6564 8044 6736 8072
rect 6564 7800 6592 8044
rect 6736 8026 6788 8032
rect 6380 7772 6592 7800
rect 6380 7070 6408 7772
rect 6644 7676 6696 7682
rect 6644 7618 6696 7624
rect 6656 7138 6684 7618
rect 6644 7132 6696 7138
rect 6644 7074 6696 7080
rect 6184 7064 6236 7070
rect 6184 7006 6236 7012
rect 6368 7064 6420 7070
rect 6368 7006 6420 7012
rect 112 6724 164 6730
rect 0 6684 112 6712
rect 112 6666 164 6672
rect 6380 6594 6408 7006
rect 6932 6712 6960 8570
rect 7012 8560 7064 8566
rect 7012 8502 7064 8508
rect 7024 8158 7052 8502
rect 7012 8152 7064 8158
rect 7012 8094 7064 8100
rect 6932 6684 7052 6712
rect 6918 6628 6974 6637
rect 6368 6588 6420 6594
rect 6918 6563 6920 6572
rect 6368 6530 6420 6536
rect 6972 6563 6974 6572
rect 6920 6530 6972 6536
rect 5796 6284 6112 6304
rect 5796 6282 5806 6284
rect 5862 6282 5886 6284
rect 5942 6282 5966 6284
rect 6022 6282 6046 6284
rect 6102 6282 6112 6284
rect 5796 6230 5800 6282
rect 5862 6230 5864 6282
rect 6044 6230 6046 6282
rect 6108 6230 6112 6282
rect 5796 6228 5806 6230
rect 5862 6228 5886 6230
rect 5942 6228 5966 6230
rect 6022 6228 6046 6230
rect 6102 6228 6112 6230
rect 5796 6208 6112 6228
rect 204 6044 256 6050
rect 204 5986 256 5992
rect 20 5840 72 5846
rect 216 5828 244 5986
rect 6380 5982 6408 6530
rect 6644 6384 6696 6390
rect 6644 6326 6696 6332
rect 6656 6118 6684 6326
rect 6644 6112 6696 6118
rect 6644 6054 6696 6060
rect 7024 5982 7052 6684
rect 7104 6656 7156 6662
rect 7104 6598 7156 6604
rect 7116 6118 7144 6598
rect 7208 6186 7236 10202
rect 7484 9858 7512 10270
rect 7472 9852 7524 9858
rect 7472 9794 7524 9800
rect 7484 8101 7512 9794
rect 7760 9382 7788 11444
rect 8036 11422 8064 11580
rect 8024 11416 8076 11422
rect 8024 11358 8076 11364
rect 8760 11416 8812 11422
rect 8864 11404 8892 12446
rect 9048 11812 9076 13756
rect 9220 13524 9272 13530
rect 9220 13466 9272 13472
rect 9232 13258 9260 13466
rect 9220 13252 9272 13258
rect 9220 13194 9272 13200
rect 9324 13122 9352 13942
rect 9496 13796 9548 13802
rect 9496 13738 9548 13744
rect 9508 13122 9536 13738
rect 9876 13122 9904 14146
rect 10336 14056 10364 14214
rect 15856 14210 15884 14368
rect 15844 14204 15896 14210
rect 15844 14146 15896 14152
rect 10336 14028 10456 14056
rect 10140 14000 10192 14006
rect 10140 13942 10192 13948
rect 9312 13116 9364 13122
rect 9312 13058 9364 13064
rect 9496 13116 9548 13122
rect 9496 13058 9548 13064
rect 9864 13116 9916 13122
rect 9864 13058 9916 13064
rect 9220 13048 9272 13054
rect 9220 12990 9272 12996
rect 9232 12034 9260 12990
rect 9220 12028 9272 12034
rect 9220 11970 9272 11976
rect 9048 11784 9168 11812
rect 8812 11376 8892 11404
rect 8760 11358 8812 11364
rect 7840 11076 7892 11082
rect 8036 11064 8064 11358
rect 8160 11180 8832 11200
rect 8160 11178 8188 11180
rect 8244 11178 8268 11180
rect 8324 11178 8348 11180
rect 8404 11178 8428 11180
rect 8484 11178 8508 11180
rect 8564 11178 8588 11180
rect 8644 11178 8668 11180
rect 8724 11178 8748 11180
rect 8804 11178 8832 11180
rect 8160 11126 8182 11178
rect 8244 11126 8246 11178
rect 8426 11126 8428 11178
rect 8490 11126 8502 11178
rect 8564 11126 8566 11178
rect 8746 11126 8748 11178
rect 8810 11126 8832 11178
rect 8160 11124 8188 11126
rect 8244 11124 8268 11126
rect 8324 11124 8348 11126
rect 8404 11124 8428 11126
rect 8484 11124 8508 11126
rect 8564 11124 8588 11126
rect 8644 11124 8668 11126
rect 8724 11124 8748 11126
rect 8804 11124 8832 11126
rect 8160 11104 8832 11124
rect 7892 11036 8064 11064
rect 7840 11018 7892 11024
rect 7932 10260 7984 10266
rect 7932 10202 7984 10208
rect 7944 9450 7972 10202
rect 7932 9444 7984 9450
rect 7932 9386 7984 9392
rect 7748 9376 7800 9382
rect 7748 9318 7800 9324
rect 8036 9314 8064 11036
rect 8760 10328 8812 10334
rect 8298 10288 8354 10297
rect 8864 10316 8892 11376
rect 9140 10996 9168 11784
rect 9508 11064 9536 13058
rect 9876 11626 9904 13058
rect 9864 11620 9916 11626
rect 9864 11562 9916 11568
rect 9956 11280 10008 11286
rect 9956 11222 10008 11228
rect 9508 11036 9628 11064
rect 9048 10968 9168 10996
rect 9048 10810 9076 10968
rect 9600 10946 9628 11036
rect 9496 10940 9548 10946
rect 9496 10882 9548 10888
rect 9588 10940 9640 10946
rect 9588 10882 9640 10888
rect 9036 10804 9088 10810
rect 9036 10746 9088 10752
rect 9508 10384 9536 10882
rect 9508 10356 9628 10384
rect 8812 10288 8892 10316
rect 8760 10270 8812 10276
rect 8298 10223 8354 10232
rect 8312 10192 8340 10223
rect 8294 10140 8300 10192
rect 8352 10140 8358 10192
rect 8160 10092 8832 10112
rect 8160 10090 8188 10092
rect 8244 10090 8268 10092
rect 8324 10090 8348 10092
rect 8404 10090 8428 10092
rect 8484 10090 8508 10092
rect 8564 10090 8588 10092
rect 8644 10090 8668 10092
rect 8724 10090 8748 10092
rect 8804 10090 8832 10092
rect 8160 10038 8182 10090
rect 8244 10038 8246 10090
rect 8426 10038 8428 10090
rect 8490 10038 8502 10090
rect 8564 10038 8566 10090
rect 8746 10038 8748 10090
rect 8810 10038 8832 10090
rect 8160 10036 8188 10038
rect 8244 10036 8268 10038
rect 8324 10036 8348 10038
rect 8404 10036 8428 10038
rect 8484 10036 8508 10038
rect 8564 10036 8588 10038
rect 8644 10036 8668 10038
rect 8724 10036 8748 10038
rect 8804 10036 8832 10038
rect 8160 10016 8832 10036
rect 8024 9308 8076 9314
rect 8024 9250 8076 9256
rect 7654 8824 7710 8833
rect 7654 8764 7710 8768
rect 7654 8759 7656 8764
rect 7708 8759 7710 8764
rect 7656 8706 7708 8712
rect 7564 8628 7616 8634
rect 7564 8570 7616 8576
rect 7576 8362 7604 8570
rect 7564 8356 7616 8362
rect 7564 8298 7616 8304
rect 7668 8226 7696 8706
rect 8036 8566 8064 9250
rect 8864 9246 8892 10288
rect 9402 10288 9458 10297
rect 9402 10223 9458 10232
rect 9416 9858 9444 10223
rect 9404 9852 9456 9858
rect 9600 9840 9628 10356
rect 9968 10198 9996 11222
rect 10152 10878 10180 13942
rect 10428 13172 10456 14028
rect 16040 13802 16068 20080
rect 16028 13796 16080 13802
rect 16028 13738 16080 13744
rect 10336 13144 10456 13172
rect 10336 12986 10364 13144
rect 10324 12980 10376 12986
rect 10324 12922 10376 12928
rect 10324 11892 10376 11898
rect 10324 11834 10376 11840
rect 10336 11082 10364 11834
rect 10324 11076 10376 11082
rect 10324 11018 10376 11024
rect 10140 10872 10192 10878
rect 10140 10814 10192 10820
rect 9864 10192 9916 10198
rect 9864 10134 9916 10140
rect 9956 10192 10008 10198
rect 9956 10134 10008 10140
rect 9876 9926 9904 10134
rect 9864 9920 9916 9926
rect 9864 9862 9916 9868
rect 9404 9794 9456 9800
rect 9508 9812 9628 9840
rect 9956 9852 10008 9858
rect 9312 9648 9364 9654
rect 9312 9590 9364 9596
rect 8852 9240 8904 9246
rect 8852 9182 8904 9188
rect 8160 9004 8832 9024
rect 8160 9002 8188 9004
rect 8244 9002 8268 9004
rect 8324 9002 8348 9004
rect 8404 9002 8428 9004
rect 8484 9002 8508 9004
rect 8564 9002 8588 9004
rect 8644 9002 8668 9004
rect 8724 9002 8748 9004
rect 8804 9002 8832 9004
rect 8160 8950 8182 9002
rect 8244 8950 8246 9002
rect 8426 8950 8428 9002
rect 8490 8950 8502 9002
rect 8564 8950 8566 9002
rect 8746 8950 8748 9002
rect 8810 8950 8832 9002
rect 8160 8948 8188 8950
rect 8244 8948 8268 8950
rect 8324 8948 8348 8950
rect 8404 8948 8428 8950
rect 8484 8948 8508 8950
rect 8564 8948 8588 8950
rect 8644 8948 8668 8950
rect 8724 8948 8748 8950
rect 8804 8948 8832 8950
rect 8160 8928 8832 8948
rect 8864 8833 8892 9182
rect 9036 9172 9088 9178
rect 9036 9114 9088 9120
rect 9048 8906 9076 9114
rect 9036 8900 9088 8906
rect 9036 8842 9088 8848
rect 8850 8824 8906 8833
rect 8850 8759 8906 8768
rect 8024 8560 8076 8566
rect 8024 8502 8076 8508
rect 9128 8560 9180 8566
rect 9128 8502 9180 8508
rect 7656 8220 7708 8226
rect 7656 8162 7708 8168
rect 7840 8152 7892 8158
rect 7470 8092 7526 8101
rect 8024 8152 8076 8158
rect 7840 8094 7892 8100
rect 8022 8100 8024 8101
rect 8076 8100 8078 8101
rect 7470 8027 7526 8036
rect 7656 8084 7708 8090
rect 7484 7682 7512 8027
rect 7656 8026 7708 8032
rect 7472 7676 7524 7682
rect 7472 7618 7524 7624
rect 7484 7070 7512 7618
rect 7668 7070 7696 8026
rect 7852 7274 7880 8094
rect 8022 8092 8078 8100
rect 8022 8027 8078 8036
rect 8852 8084 8904 8090
rect 8852 8026 8904 8032
rect 8160 7916 8832 7936
rect 8160 7914 8188 7916
rect 8244 7914 8268 7916
rect 8324 7914 8348 7916
rect 8404 7914 8428 7916
rect 8484 7914 8508 7916
rect 8564 7914 8588 7916
rect 8644 7914 8668 7916
rect 8724 7914 8748 7916
rect 8804 7914 8832 7916
rect 8160 7862 8182 7914
rect 8244 7862 8246 7914
rect 8426 7862 8428 7914
rect 8490 7862 8502 7914
rect 8564 7862 8566 7914
rect 8746 7862 8748 7914
rect 8810 7862 8832 7914
rect 8160 7860 8188 7862
rect 8244 7860 8268 7862
rect 8324 7860 8348 7862
rect 8404 7860 8428 7862
rect 8484 7860 8508 7862
rect 8564 7860 8588 7862
rect 8644 7860 8668 7862
rect 8724 7860 8748 7862
rect 8804 7860 8832 7862
rect 8160 7840 8832 7860
rect 8864 7596 8892 8026
rect 9140 7818 9168 8502
rect 9128 7812 9180 7818
rect 9128 7754 9180 7760
rect 8772 7568 8892 7596
rect 7840 7268 7892 7274
rect 7840 7210 7892 7216
rect 7472 7064 7524 7070
rect 7472 7006 7524 7012
rect 7656 7064 7708 7070
rect 7656 7006 7708 7012
rect 7484 6712 7512 7006
rect 8772 6984 8800 7568
rect 9036 7472 9088 7478
rect 9036 7414 9088 7420
rect 8772 6956 8892 6984
rect 8160 6828 8832 6848
rect 8160 6826 8188 6828
rect 8244 6826 8268 6828
rect 8324 6826 8348 6828
rect 8404 6826 8428 6828
rect 8484 6826 8508 6828
rect 8564 6826 8588 6828
rect 8644 6826 8668 6828
rect 8724 6826 8748 6828
rect 8804 6826 8832 6828
rect 8160 6774 8182 6826
rect 8244 6774 8246 6826
rect 8426 6774 8428 6826
rect 8490 6774 8502 6826
rect 8564 6774 8566 6826
rect 8746 6774 8748 6826
rect 8810 6774 8832 6826
rect 8160 6772 8188 6774
rect 8244 6772 8268 6774
rect 8324 6772 8348 6774
rect 8404 6772 8428 6774
rect 8484 6772 8508 6774
rect 8564 6772 8588 6774
rect 8644 6772 8668 6774
rect 8724 6772 8748 6774
rect 8804 6772 8832 6774
rect 8160 6752 8832 6772
rect 7392 6684 7512 6712
rect 7392 6637 7420 6684
rect 7378 6628 7434 6637
rect 7378 6563 7434 6572
rect 8668 6588 8720 6594
rect 8668 6530 8720 6536
rect 7196 6180 7248 6186
rect 7196 6122 7248 6128
rect 7104 6112 7156 6118
rect 7104 6054 7156 6060
rect 8680 5982 8708 6530
rect 8864 6186 8892 6956
rect 9048 6848 9076 7414
rect 9002 6820 9076 6848
rect 9002 6304 9030 6820
rect 9128 6724 9180 6730
rect 9128 6666 9180 6672
rect 8956 6276 9030 6304
rect 8852 6180 8904 6186
rect 8852 6122 8904 6128
rect 8956 6050 8984 6276
rect 9140 6186 9168 6666
rect 9128 6180 9180 6186
rect 9128 6122 9180 6128
rect 8944 6044 8996 6050
rect 8944 5986 8996 5992
rect 9324 5982 9352 9590
rect 9508 8362 9536 9812
rect 9956 9794 10008 9800
rect 9772 9648 9824 9654
rect 9772 9590 9824 9596
rect 9784 8702 9812 9590
rect 9968 9568 9996 9794
rect 9968 9540 10088 9568
rect 10060 8956 10088 9540
rect 10060 8928 10180 8956
rect 9862 8824 9918 8833
rect 9862 8759 9918 8768
rect 9772 8696 9824 8702
rect 9772 8638 9824 8644
rect 9588 8628 9640 8634
rect 9588 8570 9640 8576
rect 9496 8356 9548 8362
rect 9496 8298 9548 8304
rect 9600 7750 9628 8570
rect 9588 7744 9640 7750
rect 9588 7686 9640 7692
rect 9496 7676 9548 7682
rect 9496 7618 9548 7624
rect 9508 6984 9536 7618
rect 9876 7138 9904 8759
rect 9864 7132 9916 7138
rect 9864 7074 9916 7080
rect 10152 6984 10180 8928
rect 9508 6956 10180 6984
rect 9496 6384 9548 6390
rect 9496 6326 9548 6332
rect 9508 5982 9536 6326
rect 9600 6118 9628 6956
rect 9588 6112 9640 6118
rect 9588 6054 9640 6060
rect 6368 5976 6420 5982
rect 6368 5918 6420 5924
rect 7012 5976 7064 5982
rect 7012 5918 7064 5924
rect 8024 5976 8076 5982
rect 8024 5918 8076 5924
rect 8668 5976 8720 5982
rect 8668 5918 8720 5924
rect 9312 5976 9364 5982
rect 9312 5918 9364 5924
rect 9496 5976 9548 5982
rect 9496 5918 9548 5924
rect 216 5800 336 5828
rect 20 5782 72 5788
rect 32 4468 60 5782
rect 0 4440 97 4468
rect 308 4400 336 5800
rect 7024 5760 7052 5918
rect 8036 5760 8064 5918
rect 7024 5732 8064 5760
rect 8160 5740 8832 5760
rect 8160 5738 8188 5740
rect 8244 5738 8268 5740
rect 8324 5738 8348 5740
rect 8404 5738 8428 5740
rect 8484 5738 8508 5740
rect 8564 5738 8588 5740
rect 8644 5738 8668 5740
rect 8724 5738 8748 5740
rect 8804 5738 8832 5740
rect 8160 5686 8182 5738
rect 8244 5686 8246 5738
rect 8426 5686 8428 5738
rect 8490 5686 8502 5738
rect 8564 5686 8566 5738
rect 8746 5686 8748 5738
rect 8810 5686 8832 5738
rect 8160 5684 8188 5686
rect 8244 5684 8268 5686
rect 8324 5684 8348 5686
rect 8404 5684 8428 5686
rect 8484 5684 8508 5686
rect 8564 5684 8588 5686
rect 8644 5684 8668 5686
rect 8724 5684 8748 5686
rect 8804 5684 8832 5686
rect 8160 5664 8832 5684
rect 216 4372 336 4400
rect 216 2224 244 4372
rect 0 2196 244 2224
rect 14 76 20 128
rect 72 76 78 128
rect 32 48 60 76
rect 0 20 97 48
<< via2 >>
rect 202 14868 258 14924
rect 6458 14868 6514 14924
rect 5806 13898 5862 13900
rect 5886 13898 5942 13900
rect 5966 13898 6022 13900
rect 6046 13898 6102 13900
rect 5806 13846 5852 13898
rect 5852 13846 5862 13898
rect 5886 13846 5916 13898
rect 5916 13846 5928 13898
rect 5928 13846 5942 13898
rect 5966 13846 5980 13898
rect 5980 13846 5992 13898
rect 5992 13846 6022 13898
rect 6046 13846 6056 13898
rect 6056 13846 6102 13898
rect 5806 13844 5862 13846
rect 5886 13844 5942 13846
rect 5966 13844 6022 13846
rect 6046 13844 6102 13846
rect 5806 12810 5862 12812
rect 5886 12810 5942 12812
rect 5966 12810 6022 12812
rect 6046 12810 6102 12812
rect 5806 12758 5852 12810
rect 5852 12758 5862 12810
rect 5886 12758 5916 12810
rect 5916 12758 5928 12810
rect 5928 12758 5942 12810
rect 5966 12758 5980 12810
rect 5980 12758 5992 12810
rect 5992 12758 6022 12810
rect 6046 12758 6056 12810
rect 6056 12758 6102 12810
rect 5806 12756 5862 12758
rect 5886 12756 5942 12758
rect 5966 12756 6022 12758
rect 6046 12756 6102 12758
rect 5806 11722 5862 11724
rect 5886 11722 5942 11724
rect 5966 11722 6022 11724
rect 6046 11722 6102 11724
rect 5806 11670 5852 11722
rect 5852 11670 5862 11722
rect 5886 11670 5916 11722
rect 5916 11670 5928 11722
rect 5928 11670 5942 11722
rect 5966 11670 5980 11722
rect 5980 11670 5992 11722
rect 5992 11670 6022 11722
rect 6046 11670 6056 11722
rect 6056 11670 6102 11722
rect 5806 11668 5862 11670
rect 5886 11668 5942 11670
rect 5966 11668 6022 11670
rect 6046 11668 6102 11670
rect 5806 10634 5862 10636
rect 5886 10634 5942 10636
rect 5966 10634 6022 10636
rect 6046 10634 6102 10636
rect 5806 10582 5852 10634
rect 5852 10582 5862 10634
rect 5886 10582 5916 10634
rect 5916 10582 5928 10634
rect 5928 10582 5942 10634
rect 5966 10582 5980 10634
rect 5980 10582 5992 10634
rect 5992 10582 6022 10634
rect 6046 10582 6056 10634
rect 6056 10582 6102 10634
rect 5806 10580 5862 10582
rect 5886 10580 5942 10582
rect 5966 10580 6022 10582
rect 6046 10580 6102 10582
rect 5806 9546 5862 9548
rect 5886 9546 5942 9548
rect 5966 9546 6022 9548
rect 6046 9546 6102 9548
rect 5806 9494 5852 9546
rect 5852 9494 5862 9546
rect 5886 9494 5916 9546
rect 5916 9494 5928 9546
rect 5928 9494 5942 9546
rect 5966 9494 5980 9546
rect 5980 9494 5992 9546
rect 5992 9494 6022 9546
rect 6046 9494 6056 9546
rect 6056 9494 6102 9546
rect 5806 9492 5862 9494
rect 5886 9492 5942 9494
rect 5966 9492 6022 9494
rect 6046 9492 6102 9494
rect 8188 14442 8244 14444
rect 8268 14442 8324 14444
rect 8348 14442 8404 14444
rect 8428 14442 8484 14444
rect 8508 14442 8564 14444
rect 8588 14442 8644 14444
rect 8668 14442 8724 14444
rect 8748 14442 8804 14444
rect 8188 14390 8234 14442
rect 8234 14390 8244 14442
rect 8268 14390 8298 14442
rect 8298 14390 8310 14442
rect 8310 14390 8324 14442
rect 8348 14390 8362 14442
rect 8362 14390 8374 14442
rect 8374 14390 8404 14442
rect 8428 14390 8438 14442
rect 8438 14390 8484 14442
rect 8508 14390 8554 14442
rect 8554 14390 8564 14442
rect 8588 14390 8618 14442
rect 8618 14390 8630 14442
rect 8630 14390 8644 14442
rect 8668 14390 8682 14442
rect 8682 14390 8694 14442
rect 8694 14390 8724 14442
rect 8748 14390 8758 14442
rect 8758 14390 8804 14442
rect 8188 14388 8244 14390
rect 8268 14388 8324 14390
rect 8348 14388 8404 14390
rect 8428 14388 8484 14390
rect 8508 14388 8564 14390
rect 8588 14388 8644 14390
rect 8668 14388 8724 14390
rect 8748 14388 8804 14390
rect 8188 13354 8244 13356
rect 8268 13354 8324 13356
rect 8348 13354 8404 13356
rect 8428 13354 8484 13356
rect 8508 13354 8564 13356
rect 8588 13354 8644 13356
rect 8668 13354 8724 13356
rect 8748 13354 8804 13356
rect 8188 13302 8234 13354
rect 8234 13302 8244 13354
rect 8268 13302 8298 13354
rect 8298 13302 8310 13354
rect 8310 13302 8324 13354
rect 8348 13302 8362 13354
rect 8362 13302 8374 13354
rect 8374 13302 8404 13354
rect 8428 13302 8438 13354
rect 8438 13302 8484 13354
rect 8508 13302 8554 13354
rect 8554 13302 8564 13354
rect 8588 13302 8618 13354
rect 8618 13302 8630 13354
rect 8630 13302 8644 13354
rect 8668 13302 8682 13354
rect 8682 13302 8694 13354
rect 8694 13302 8724 13354
rect 8748 13302 8758 13354
rect 8758 13302 8804 13354
rect 8188 13300 8244 13302
rect 8268 13300 8324 13302
rect 8348 13300 8404 13302
rect 8428 13300 8484 13302
rect 8508 13300 8564 13302
rect 8588 13300 8644 13302
rect 8668 13300 8724 13302
rect 8748 13300 8804 13302
rect 6458 10720 6514 10776
rect 5806 8458 5862 8460
rect 5886 8458 5942 8460
rect 5966 8458 6022 8460
rect 6046 8458 6102 8460
rect 5806 8406 5852 8458
rect 5852 8406 5862 8458
rect 5886 8406 5916 8458
rect 5916 8406 5928 8458
rect 5928 8406 5942 8458
rect 5966 8406 5980 8458
rect 5980 8406 5992 8458
rect 5992 8406 6022 8458
rect 6046 8406 6056 8458
rect 6056 8406 6102 8458
rect 5806 8404 5862 8406
rect 5886 8404 5942 8406
rect 5966 8404 6022 8406
rect 6046 8404 6102 8406
rect 5806 7370 5862 7372
rect 5886 7370 5942 7372
rect 5966 7370 6022 7372
rect 6046 7370 6102 7372
rect 5806 7318 5852 7370
rect 5852 7318 5862 7370
rect 5886 7318 5916 7370
rect 5916 7318 5928 7370
rect 5928 7318 5942 7370
rect 5966 7318 5980 7370
rect 5980 7318 5992 7370
rect 5992 7318 6022 7370
rect 6046 7318 6056 7370
rect 6056 7318 6102 7370
rect 5806 7316 5862 7318
rect 5886 7316 5942 7318
rect 5966 7316 6022 7318
rect 6046 7316 6102 7318
rect 8188 12266 8244 12268
rect 8268 12266 8324 12268
rect 8348 12266 8404 12268
rect 8428 12266 8484 12268
rect 8508 12266 8564 12268
rect 8588 12266 8644 12268
rect 8668 12266 8724 12268
rect 8748 12266 8804 12268
rect 8188 12214 8234 12266
rect 8234 12214 8244 12266
rect 8268 12214 8298 12266
rect 8298 12214 8310 12266
rect 8310 12214 8324 12266
rect 8348 12214 8362 12266
rect 8362 12214 8374 12266
rect 8374 12214 8404 12266
rect 8428 12214 8438 12266
rect 8438 12214 8484 12266
rect 8508 12214 8554 12266
rect 8554 12214 8564 12266
rect 8588 12214 8618 12266
rect 8618 12214 8630 12266
rect 8630 12214 8644 12266
rect 8668 12214 8682 12266
rect 8682 12214 8694 12266
rect 8694 12214 8724 12266
rect 8748 12214 8758 12266
rect 8758 12214 8804 12266
rect 8188 12212 8244 12214
rect 8268 12212 8324 12214
rect 8348 12212 8404 12214
rect 8428 12212 8484 12214
rect 8508 12212 8564 12214
rect 8588 12212 8644 12214
rect 8668 12212 8724 12214
rect 8748 12212 8804 12214
rect 7654 10720 7710 10776
rect 6734 8768 6790 8824
rect 6918 6588 6974 6628
rect 6918 6572 6920 6588
rect 6920 6572 6972 6588
rect 6972 6572 6974 6588
rect 5806 6282 5862 6284
rect 5886 6282 5942 6284
rect 5966 6282 6022 6284
rect 6046 6282 6102 6284
rect 5806 6230 5852 6282
rect 5852 6230 5862 6282
rect 5886 6230 5916 6282
rect 5916 6230 5928 6282
rect 5928 6230 5942 6282
rect 5966 6230 5980 6282
rect 5980 6230 5992 6282
rect 5992 6230 6022 6282
rect 6046 6230 6056 6282
rect 6056 6230 6102 6282
rect 5806 6228 5862 6230
rect 5886 6228 5942 6230
rect 5966 6228 6022 6230
rect 6046 6228 6102 6230
rect 8188 11178 8244 11180
rect 8268 11178 8324 11180
rect 8348 11178 8404 11180
rect 8428 11178 8484 11180
rect 8508 11178 8564 11180
rect 8588 11178 8644 11180
rect 8668 11178 8724 11180
rect 8748 11178 8804 11180
rect 8188 11126 8234 11178
rect 8234 11126 8244 11178
rect 8268 11126 8298 11178
rect 8298 11126 8310 11178
rect 8310 11126 8324 11178
rect 8348 11126 8362 11178
rect 8362 11126 8374 11178
rect 8374 11126 8404 11178
rect 8428 11126 8438 11178
rect 8438 11126 8484 11178
rect 8508 11126 8554 11178
rect 8554 11126 8564 11178
rect 8588 11126 8618 11178
rect 8618 11126 8630 11178
rect 8630 11126 8644 11178
rect 8668 11126 8682 11178
rect 8682 11126 8694 11178
rect 8694 11126 8724 11178
rect 8748 11126 8758 11178
rect 8758 11126 8804 11178
rect 8188 11124 8244 11126
rect 8268 11124 8324 11126
rect 8348 11124 8404 11126
rect 8428 11124 8484 11126
rect 8508 11124 8564 11126
rect 8588 11124 8644 11126
rect 8668 11124 8724 11126
rect 8748 11124 8804 11126
rect 8298 10232 8354 10288
rect 8188 10090 8244 10092
rect 8268 10090 8324 10092
rect 8348 10090 8404 10092
rect 8428 10090 8484 10092
rect 8508 10090 8564 10092
rect 8588 10090 8644 10092
rect 8668 10090 8724 10092
rect 8748 10090 8804 10092
rect 8188 10038 8234 10090
rect 8234 10038 8244 10090
rect 8268 10038 8298 10090
rect 8298 10038 8310 10090
rect 8310 10038 8324 10090
rect 8348 10038 8362 10090
rect 8362 10038 8374 10090
rect 8374 10038 8404 10090
rect 8428 10038 8438 10090
rect 8438 10038 8484 10090
rect 8508 10038 8554 10090
rect 8554 10038 8564 10090
rect 8588 10038 8618 10090
rect 8618 10038 8630 10090
rect 8630 10038 8644 10090
rect 8668 10038 8682 10090
rect 8682 10038 8694 10090
rect 8694 10038 8724 10090
rect 8748 10038 8758 10090
rect 8758 10038 8804 10090
rect 8188 10036 8244 10038
rect 8268 10036 8324 10038
rect 8348 10036 8404 10038
rect 8428 10036 8484 10038
rect 8508 10036 8564 10038
rect 8588 10036 8644 10038
rect 8668 10036 8724 10038
rect 8748 10036 8804 10038
rect 7654 8768 7710 8824
rect 9402 10232 9458 10288
rect 8188 9002 8244 9004
rect 8268 9002 8324 9004
rect 8348 9002 8404 9004
rect 8428 9002 8484 9004
rect 8508 9002 8564 9004
rect 8588 9002 8644 9004
rect 8668 9002 8724 9004
rect 8748 9002 8804 9004
rect 8188 8950 8234 9002
rect 8234 8950 8244 9002
rect 8268 8950 8298 9002
rect 8298 8950 8310 9002
rect 8310 8950 8324 9002
rect 8348 8950 8362 9002
rect 8362 8950 8374 9002
rect 8374 8950 8404 9002
rect 8428 8950 8438 9002
rect 8438 8950 8484 9002
rect 8508 8950 8554 9002
rect 8554 8950 8564 9002
rect 8588 8950 8618 9002
rect 8618 8950 8630 9002
rect 8630 8950 8644 9002
rect 8668 8950 8682 9002
rect 8682 8950 8694 9002
rect 8694 8950 8724 9002
rect 8748 8950 8758 9002
rect 8758 8950 8804 9002
rect 8188 8948 8244 8950
rect 8268 8948 8324 8950
rect 8348 8948 8404 8950
rect 8428 8948 8484 8950
rect 8508 8948 8564 8950
rect 8588 8948 8644 8950
rect 8668 8948 8724 8950
rect 8748 8948 8804 8950
rect 8850 8768 8906 8824
rect 7470 8036 7526 8092
rect 8022 8036 8078 8092
rect 8188 7914 8244 7916
rect 8268 7914 8324 7916
rect 8348 7914 8404 7916
rect 8428 7914 8484 7916
rect 8508 7914 8564 7916
rect 8588 7914 8644 7916
rect 8668 7914 8724 7916
rect 8748 7914 8804 7916
rect 8188 7862 8234 7914
rect 8234 7862 8244 7914
rect 8268 7862 8298 7914
rect 8298 7862 8310 7914
rect 8310 7862 8324 7914
rect 8348 7862 8362 7914
rect 8362 7862 8374 7914
rect 8374 7862 8404 7914
rect 8428 7862 8438 7914
rect 8438 7862 8484 7914
rect 8508 7862 8554 7914
rect 8554 7862 8564 7914
rect 8588 7862 8618 7914
rect 8618 7862 8630 7914
rect 8630 7862 8644 7914
rect 8668 7862 8682 7914
rect 8682 7862 8694 7914
rect 8694 7862 8724 7914
rect 8748 7862 8758 7914
rect 8758 7862 8804 7914
rect 8188 7860 8244 7862
rect 8268 7860 8324 7862
rect 8348 7860 8404 7862
rect 8428 7860 8484 7862
rect 8508 7860 8564 7862
rect 8588 7860 8644 7862
rect 8668 7860 8724 7862
rect 8748 7860 8804 7862
rect 8188 6826 8244 6828
rect 8268 6826 8324 6828
rect 8348 6826 8404 6828
rect 8428 6826 8484 6828
rect 8508 6826 8564 6828
rect 8588 6826 8644 6828
rect 8668 6826 8724 6828
rect 8748 6826 8804 6828
rect 8188 6774 8234 6826
rect 8234 6774 8244 6826
rect 8268 6774 8298 6826
rect 8298 6774 8310 6826
rect 8310 6774 8324 6826
rect 8348 6774 8362 6826
rect 8362 6774 8374 6826
rect 8374 6774 8404 6826
rect 8428 6774 8438 6826
rect 8438 6774 8484 6826
rect 8508 6774 8554 6826
rect 8554 6774 8564 6826
rect 8588 6774 8618 6826
rect 8618 6774 8630 6826
rect 8630 6774 8644 6826
rect 8668 6774 8682 6826
rect 8682 6774 8694 6826
rect 8694 6774 8724 6826
rect 8748 6774 8758 6826
rect 8758 6774 8804 6826
rect 8188 6772 8244 6774
rect 8268 6772 8324 6774
rect 8348 6772 8404 6774
rect 8428 6772 8484 6774
rect 8508 6772 8564 6774
rect 8588 6772 8644 6774
rect 8668 6772 8724 6774
rect 8748 6772 8804 6774
rect 7378 6572 7434 6628
rect 9862 8768 9918 8824
rect 8188 5738 8244 5740
rect 8268 5738 8324 5740
rect 8348 5738 8404 5740
rect 8428 5738 8484 5740
rect 8508 5738 8564 5740
rect 8588 5738 8644 5740
rect 8668 5738 8724 5740
rect 8748 5738 8804 5740
rect 8188 5686 8234 5738
rect 8234 5686 8244 5738
rect 8268 5686 8298 5738
rect 8298 5686 8310 5738
rect 8310 5686 8324 5738
rect 8348 5686 8362 5738
rect 8362 5686 8374 5738
rect 8374 5686 8404 5738
rect 8428 5686 8438 5738
rect 8438 5686 8484 5738
rect 8508 5686 8554 5738
rect 8554 5686 8564 5738
rect 8588 5686 8618 5738
rect 8618 5686 8630 5738
rect 8630 5686 8644 5738
rect 8668 5686 8682 5738
rect 8682 5686 8694 5738
rect 8694 5686 8724 5738
rect 8748 5686 8758 5738
rect 8758 5686 8804 5738
rect 8188 5684 8244 5686
rect 8268 5684 8324 5686
rect 8348 5684 8404 5686
rect 8428 5684 8484 5686
rect 8508 5684 8564 5686
rect 8588 5684 8644 5686
rect 8668 5684 8724 5686
rect 8748 5684 8804 5686
<< metal3 >>
rect 197 14926 263 14929
rect 6453 14926 6519 14929
rect 197 14924 6519 14926
rect 197 14868 202 14924
rect 258 14868 6458 14924
rect 6514 14868 6519 14924
rect 197 14866 6519 14868
rect 197 14863 263 14866
rect 6453 14863 6519 14866
rect 8160 14448 8832 14464
rect 8160 14384 8184 14448
rect 8248 14384 8264 14448
rect 8328 14384 8344 14448
rect 8408 14384 8424 14448
rect 8488 14384 8504 14448
rect 8568 14384 8584 14448
rect 8648 14384 8664 14448
rect 8728 14384 8744 14448
rect 8808 14384 8832 14448
rect 8160 14368 8832 14384
rect 5796 13904 6112 13920
rect 5796 13840 5802 13904
rect 5866 13840 5882 13904
rect 5946 13840 5962 13904
rect 6026 13840 6042 13904
rect 6106 13840 6112 13904
rect 5796 13824 6112 13840
rect 8160 13360 8832 13376
rect 8160 13296 8184 13360
rect 8248 13296 8264 13360
rect 8328 13296 8344 13360
rect 8408 13296 8424 13360
rect 8488 13296 8504 13360
rect 8568 13296 8584 13360
rect 8648 13296 8664 13360
rect 8728 13296 8744 13360
rect 8808 13296 8832 13360
rect 8160 13280 8832 13296
rect 5796 12816 6112 12832
rect 5796 12752 5802 12816
rect 5866 12752 5882 12816
rect 5946 12752 5962 12816
rect 6026 12752 6042 12816
rect 6106 12752 6112 12816
rect 5796 12736 6112 12752
rect 8160 12272 8832 12288
rect 8160 12208 8184 12272
rect 8248 12208 8264 12272
rect 8328 12208 8344 12272
rect 8408 12208 8424 12272
rect 8488 12208 8504 12272
rect 8568 12208 8584 12272
rect 8648 12208 8664 12272
rect 8728 12208 8744 12272
rect 8808 12208 8832 12272
rect 8160 12192 8832 12208
rect 5796 11728 6112 11744
rect 5796 11664 5802 11728
rect 5866 11664 5882 11728
rect 5946 11664 5962 11728
rect 6026 11664 6042 11728
rect 6106 11664 6112 11728
rect 5796 11648 6112 11664
rect 8160 11184 8832 11200
rect 8160 11120 8184 11184
rect 8248 11120 8264 11184
rect 8328 11120 8344 11184
rect 8408 11120 8424 11184
rect 8488 11120 8504 11184
rect 8568 11120 8584 11184
rect 8648 11120 8664 11184
rect 8728 11120 8744 11184
rect 8808 11120 8832 11184
rect 8160 11104 8832 11120
rect 6453 10778 6519 10781
rect 7649 10778 7715 10781
rect 6453 10776 7715 10778
rect 6453 10720 6458 10776
rect 6514 10720 7654 10776
rect 7710 10720 7715 10776
rect 6453 10718 7715 10720
rect 6453 10715 6519 10718
rect 7649 10715 7715 10718
rect 5796 10640 6112 10656
rect 5796 10576 5802 10640
rect 5866 10576 5882 10640
rect 5946 10576 5962 10640
rect 6026 10576 6042 10640
rect 6106 10576 6112 10640
rect 5796 10560 6112 10576
rect 8293 10290 8359 10293
rect 9397 10290 9463 10293
rect 8293 10288 9463 10290
rect 8293 10232 8298 10288
rect 8354 10232 9402 10288
rect 9458 10232 9463 10288
rect 8293 10230 9463 10232
rect 8293 10227 8359 10230
rect 9397 10227 9463 10230
rect 8160 10096 8832 10112
rect 8160 10032 8184 10096
rect 8248 10032 8264 10096
rect 8328 10032 8344 10096
rect 8408 10032 8424 10096
rect 8488 10032 8504 10096
rect 8568 10032 8584 10096
rect 8648 10032 8664 10096
rect 8728 10032 8744 10096
rect 8808 10032 8832 10096
rect 8160 10016 8832 10032
rect 5796 9552 6112 9568
rect 5796 9488 5802 9552
rect 5866 9488 5882 9552
rect 5946 9488 5962 9552
rect 6026 9488 6042 9552
rect 6106 9488 6112 9552
rect 5796 9472 6112 9488
rect 8160 9008 8832 9024
rect 8160 8944 8184 9008
rect 8248 8944 8264 9008
rect 8328 8944 8344 9008
rect 8408 8944 8424 9008
rect 8488 8944 8504 9008
rect 8568 8944 8584 9008
rect 8648 8944 8664 9008
rect 8728 8944 8744 9008
rect 8808 8944 8832 9008
rect 8160 8928 8832 8944
rect 6729 8826 6795 8829
rect 7649 8826 7715 8829
rect 8845 8826 8911 8829
rect 9857 8826 9923 8829
rect 6729 8824 9923 8826
rect 6729 8768 6734 8824
rect 6790 8768 7654 8824
rect 7710 8768 8850 8824
rect 8906 8768 9862 8824
rect 9918 8768 9923 8824
rect 6729 8766 9923 8768
rect 6729 8763 6795 8766
rect 7649 8763 7715 8766
rect 8845 8763 8911 8766
rect 9857 8763 9923 8766
rect 5796 8464 6112 8480
rect 5796 8400 5802 8464
rect 5866 8400 5882 8464
rect 5946 8400 5962 8464
rect 6026 8400 6042 8464
rect 6106 8400 6112 8464
rect 5796 8384 6112 8400
rect 7465 8094 7531 8097
rect 8017 8094 8083 8097
rect 7465 8092 8083 8094
rect 7465 8036 7470 8092
rect 7526 8036 8022 8092
rect 8078 8036 8083 8092
rect 7465 8034 8083 8036
rect 7465 8031 7531 8034
rect 8017 8031 8083 8034
rect 8160 7920 8832 7936
rect 8160 7856 8184 7920
rect 8248 7856 8264 7920
rect 8328 7856 8344 7920
rect 8408 7856 8424 7920
rect 8488 7856 8504 7920
rect 8568 7856 8584 7920
rect 8648 7856 8664 7920
rect 8728 7856 8744 7920
rect 8808 7856 8832 7920
rect 8160 7840 8832 7856
rect 5796 7376 6112 7392
rect 5796 7312 5802 7376
rect 5866 7312 5882 7376
rect 5946 7312 5962 7376
rect 6026 7312 6042 7376
rect 6106 7312 6112 7376
rect 5796 7296 6112 7312
rect 8160 6832 8832 6848
rect 8160 6768 8184 6832
rect 8248 6768 8264 6832
rect 8328 6768 8344 6832
rect 8408 6768 8424 6832
rect 8488 6768 8504 6832
rect 8568 6768 8584 6832
rect 8648 6768 8664 6832
rect 8728 6768 8744 6832
rect 8808 6768 8832 6832
rect 8160 6752 8832 6768
rect 6913 6630 6979 6633
rect 7373 6630 7439 6633
rect 6913 6628 7439 6630
rect 6913 6572 6918 6628
rect 6974 6572 7378 6628
rect 7434 6572 7439 6628
rect 6913 6570 7439 6572
rect 6913 6567 6979 6570
rect 7373 6567 7439 6570
rect 5796 6288 6112 6304
rect 5796 6224 5802 6288
rect 5866 6224 5882 6288
rect 5946 6224 5962 6288
rect 6026 6224 6042 6288
rect 6106 6224 6112 6288
rect 5796 6208 6112 6224
rect 8160 5744 8832 5760
rect 8160 5680 8184 5744
rect 8248 5680 8264 5744
rect 8328 5680 8344 5744
rect 8408 5680 8424 5744
rect 8488 5680 8504 5744
rect 8568 5680 8584 5744
rect 8648 5680 8664 5744
rect 8728 5680 8744 5744
rect 8808 5680 8832 5744
rect 8160 5664 8832 5680
<< via3 >>
rect 8184 14444 8248 14448
rect 8184 14388 8188 14444
rect 8188 14388 8244 14444
rect 8244 14388 8248 14444
rect 8184 14384 8248 14388
rect 8264 14444 8328 14448
rect 8264 14388 8268 14444
rect 8268 14388 8324 14444
rect 8324 14388 8328 14444
rect 8264 14384 8328 14388
rect 8344 14444 8408 14448
rect 8344 14388 8348 14444
rect 8348 14388 8404 14444
rect 8404 14388 8408 14444
rect 8344 14384 8408 14388
rect 8424 14444 8488 14448
rect 8424 14388 8428 14444
rect 8428 14388 8484 14444
rect 8484 14388 8488 14444
rect 8424 14384 8488 14388
rect 8504 14444 8568 14448
rect 8504 14388 8508 14444
rect 8508 14388 8564 14444
rect 8564 14388 8568 14444
rect 8504 14384 8568 14388
rect 8584 14444 8648 14448
rect 8584 14388 8588 14444
rect 8588 14388 8644 14444
rect 8644 14388 8648 14444
rect 8584 14384 8648 14388
rect 8664 14444 8728 14448
rect 8664 14388 8668 14444
rect 8668 14388 8724 14444
rect 8724 14388 8728 14444
rect 8664 14384 8728 14388
rect 8744 14444 8808 14448
rect 8744 14388 8748 14444
rect 8748 14388 8804 14444
rect 8804 14388 8808 14444
rect 8744 14384 8808 14388
rect 5802 13900 5866 13904
rect 5802 13844 5806 13900
rect 5806 13844 5862 13900
rect 5862 13844 5866 13900
rect 5802 13840 5866 13844
rect 5882 13900 5946 13904
rect 5882 13844 5886 13900
rect 5886 13844 5942 13900
rect 5942 13844 5946 13900
rect 5882 13840 5946 13844
rect 5962 13900 6026 13904
rect 5962 13844 5966 13900
rect 5966 13844 6022 13900
rect 6022 13844 6026 13900
rect 5962 13840 6026 13844
rect 6042 13900 6106 13904
rect 6042 13844 6046 13900
rect 6046 13844 6102 13900
rect 6102 13844 6106 13900
rect 6042 13840 6106 13844
rect 8184 13356 8248 13360
rect 8184 13300 8188 13356
rect 8188 13300 8244 13356
rect 8244 13300 8248 13356
rect 8184 13296 8248 13300
rect 8264 13356 8328 13360
rect 8264 13300 8268 13356
rect 8268 13300 8324 13356
rect 8324 13300 8328 13356
rect 8264 13296 8328 13300
rect 8344 13356 8408 13360
rect 8344 13300 8348 13356
rect 8348 13300 8404 13356
rect 8404 13300 8408 13356
rect 8344 13296 8408 13300
rect 8424 13356 8488 13360
rect 8424 13300 8428 13356
rect 8428 13300 8484 13356
rect 8484 13300 8488 13356
rect 8424 13296 8488 13300
rect 8504 13356 8568 13360
rect 8504 13300 8508 13356
rect 8508 13300 8564 13356
rect 8564 13300 8568 13356
rect 8504 13296 8568 13300
rect 8584 13356 8648 13360
rect 8584 13300 8588 13356
rect 8588 13300 8644 13356
rect 8644 13300 8648 13356
rect 8584 13296 8648 13300
rect 8664 13356 8728 13360
rect 8664 13300 8668 13356
rect 8668 13300 8724 13356
rect 8724 13300 8728 13356
rect 8664 13296 8728 13300
rect 8744 13356 8808 13360
rect 8744 13300 8748 13356
rect 8748 13300 8804 13356
rect 8804 13300 8808 13356
rect 8744 13296 8808 13300
rect 5802 12812 5866 12816
rect 5802 12756 5806 12812
rect 5806 12756 5862 12812
rect 5862 12756 5866 12812
rect 5802 12752 5866 12756
rect 5882 12812 5946 12816
rect 5882 12756 5886 12812
rect 5886 12756 5942 12812
rect 5942 12756 5946 12812
rect 5882 12752 5946 12756
rect 5962 12812 6026 12816
rect 5962 12756 5966 12812
rect 5966 12756 6022 12812
rect 6022 12756 6026 12812
rect 5962 12752 6026 12756
rect 6042 12812 6106 12816
rect 6042 12756 6046 12812
rect 6046 12756 6102 12812
rect 6102 12756 6106 12812
rect 6042 12752 6106 12756
rect 8184 12268 8248 12272
rect 8184 12212 8188 12268
rect 8188 12212 8244 12268
rect 8244 12212 8248 12268
rect 8184 12208 8248 12212
rect 8264 12268 8328 12272
rect 8264 12212 8268 12268
rect 8268 12212 8324 12268
rect 8324 12212 8328 12268
rect 8264 12208 8328 12212
rect 8344 12268 8408 12272
rect 8344 12212 8348 12268
rect 8348 12212 8404 12268
rect 8404 12212 8408 12268
rect 8344 12208 8408 12212
rect 8424 12268 8488 12272
rect 8424 12212 8428 12268
rect 8428 12212 8484 12268
rect 8484 12212 8488 12268
rect 8424 12208 8488 12212
rect 8504 12268 8568 12272
rect 8504 12212 8508 12268
rect 8508 12212 8564 12268
rect 8564 12212 8568 12268
rect 8504 12208 8568 12212
rect 8584 12268 8648 12272
rect 8584 12212 8588 12268
rect 8588 12212 8644 12268
rect 8644 12212 8648 12268
rect 8584 12208 8648 12212
rect 8664 12268 8728 12272
rect 8664 12212 8668 12268
rect 8668 12212 8724 12268
rect 8724 12212 8728 12268
rect 8664 12208 8728 12212
rect 8744 12268 8808 12272
rect 8744 12212 8748 12268
rect 8748 12212 8804 12268
rect 8804 12212 8808 12268
rect 8744 12208 8808 12212
rect 5802 11724 5866 11728
rect 5802 11668 5806 11724
rect 5806 11668 5862 11724
rect 5862 11668 5866 11724
rect 5802 11664 5866 11668
rect 5882 11724 5946 11728
rect 5882 11668 5886 11724
rect 5886 11668 5942 11724
rect 5942 11668 5946 11724
rect 5882 11664 5946 11668
rect 5962 11724 6026 11728
rect 5962 11668 5966 11724
rect 5966 11668 6022 11724
rect 6022 11668 6026 11724
rect 5962 11664 6026 11668
rect 6042 11724 6106 11728
rect 6042 11668 6046 11724
rect 6046 11668 6102 11724
rect 6102 11668 6106 11724
rect 6042 11664 6106 11668
rect 8184 11180 8248 11184
rect 8184 11124 8188 11180
rect 8188 11124 8244 11180
rect 8244 11124 8248 11180
rect 8184 11120 8248 11124
rect 8264 11180 8328 11184
rect 8264 11124 8268 11180
rect 8268 11124 8324 11180
rect 8324 11124 8328 11180
rect 8264 11120 8328 11124
rect 8344 11180 8408 11184
rect 8344 11124 8348 11180
rect 8348 11124 8404 11180
rect 8404 11124 8408 11180
rect 8344 11120 8408 11124
rect 8424 11180 8488 11184
rect 8424 11124 8428 11180
rect 8428 11124 8484 11180
rect 8484 11124 8488 11180
rect 8424 11120 8488 11124
rect 8504 11180 8568 11184
rect 8504 11124 8508 11180
rect 8508 11124 8564 11180
rect 8564 11124 8568 11180
rect 8504 11120 8568 11124
rect 8584 11180 8648 11184
rect 8584 11124 8588 11180
rect 8588 11124 8644 11180
rect 8644 11124 8648 11180
rect 8584 11120 8648 11124
rect 8664 11180 8728 11184
rect 8664 11124 8668 11180
rect 8668 11124 8724 11180
rect 8724 11124 8728 11180
rect 8664 11120 8728 11124
rect 8744 11180 8808 11184
rect 8744 11124 8748 11180
rect 8748 11124 8804 11180
rect 8804 11124 8808 11180
rect 8744 11120 8808 11124
rect 5802 10636 5866 10640
rect 5802 10580 5806 10636
rect 5806 10580 5862 10636
rect 5862 10580 5866 10636
rect 5802 10576 5866 10580
rect 5882 10636 5946 10640
rect 5882 10580 5886 10636
rect 5886 10580 5942 10636
rect 5942 10580 5946 10636
rect 5882 10576 5946 10580
rect 5962 10636 6026 10640
rect 5962 10580 5966 10636
rect 5966 10580 6022 10636
rect 6022 10580 6026 10636
rect 5962 10576 6026 10580
rect 6042 10636 6106 10640
rect 6042 10580 6046 10636
rect 6046 10580 6102 10636
rect 6102 10580 6106 10636
rect 6042 10576 6106 10580
rect 8184 10092 8248 10096
rect 8184 10036 8188 10092
rect 8188 10036 8244 10092
rect 8244 10036 8248 10092
rect 8184 10032 8248 10036
rect 8264 10092 8328 10096
rect 8264 10036 8268 10092
rect 8268 10036 8324 10092
rect 8324 10036 8328 10092
rect 8264 10032 8328 10036
rect 8344 10092 8408 10096
rect 8344 10036 8348 10092
rect 8348 10036 8404 10092
rect 8404 10036 8408 10092
rect 8344 10032 8408 10036
rect 8424 10092 8488 10096
rect 8424 10036 8428 10092
rect 8428 10036 8484 10092
rect 8484 10036 8488 10092
rect 8424 10032 8488 10036
rect 8504 10092 8568 10096
rect 8504 10036 8508 10092
rect 8508 10036 8564 10092
rect 8564 10036 8568 10092
rect 8504 10032 8568 10036
rect 8584 10092 8648 10096
rect 8584 10036 8588 10092
rect 8588 10036 8644 10092
rect 8644 10036 8648 10092
rect 8584 10032 8648 10036
rect 8664 10092 8728 10096
rect 8664 10036 8668 10092
rect 8668 10036 8724 10092
rect 8724 10036 8728 10092
rect 8664 10032 8728 10036
rect 8744 10092 8808 10096
rect 8744 10036 8748 10092
rect 8748 10036 8804 10092
rect 8804 10036 8808 10092
rect 8744 10032 8808 10036
rect 5802 9548 5866 9552
rect 5802 9492 5806 9548
rect 5806 9492 5862 9548
rect 5862 9492 5866 9548
rect 5802 9488 5866 9492
rect 5882 9548 5946 9552
rect 5882 9492 5886 9548
rect 5886 9492 5942 9548
rect 5942 9492 5946 9548
rect 5882 9488 5946 9492
rect 5962 9548 6026 9552
rect 5962 9492 5966 9548
rect 5966 9492 6022 9548
rect 6022 9492 6026 9548
rect 5962 9488 6026 9492
rect 6042 9548 6106 9552
rect 6042 9492 6046 9548
rect 6046 9492 6102 9548
rect 6102 9492 6106 9548
rect 6042 9488 6106 9492
rect 8184 9004 8248 9008
rect 8184 8948 8188 9004
rect 8188 8948 8244 9004
rect 8244 8948 8248 9004
rect 8184 8944 8248 8948
rect 8264 9004 8328 9008
rect 8264 8948 8268 9004
rect 8268 8948 8324 9004
rect 8324 8948 8328 9004
rect 8264 8944 8328 8948
rect 8344 9004 8408 9008
rect 8344 8948 8348 9004
rect 8348 8948 8404 9004
rect 8404 8948 8408 9004
rect 8344 8944 8408 8948
rect 8424 9004 8488 9008
rect 8424 8948 8428 9004
rect 8428 8948 8484 9004
rect 8484 8948 8488 9004
rect 8424 8944 8488 8948
rect 8504 9004 8568 9008
rect 8504 8948 8508 9004
rect 8508 8948 8564 9004
rect 8564 8948 8568 9004
rect 8504 8944 8568 8948
rect 8584 9004 8648 9008
rect 8584 8948 8588 9004
rect 8588 8948 8644 9004
rect 8644 8948 8648 9004
rect 8584 8944 8648 8948
rect 8664 9004 8728 9008
rect 8664 8948 8668 9004
rect 8668 8948 8724 9004
rect 8724 8948 8728 9004
rect 8664 8944 8728 8948
rect 8744 9004 8808 9008
rect 8744 8948 8748 9004
rect 8748 8948 8804 9004
rect 8804 8948 8808 9004
rect 8744 8944 8808 8948
rect 5802 8460 5866 8464
rect 5802 8404 5806 8460
rect 5806 8404 5862 8460
rect 5862 8404 5866 8460
rect 5802 8400 5866 8404
rect 5882 8460 5946 8464
rect 5882 8404 5886 8460
rect 5886 8404 5942 8460
rect 5942 8404 5946 8460
rect 5882 8400 5946 8404
rect 5962 8460 6026 8464
rect 5962 8404 5966 8460
rect 5966 8404 6022 8460
rect 6022 8404 6026 8460
rect 5962 8400 6026 8404
rect 6042 8460 6106 8464
rect 6042 8404 6046 8460
rect 6046 8404 6102 8460
rect 6102 8404 6106 8460
rect 6042 8400 6106 8404
rect 8184 7916 8248 7920
rect 8184 7860 8188 7916
rect 8188 7860 8244 7916
rect 8244 7860 8248 7916
rect 8184 7856 8248 7860
rect 8264 7916 8328 7920
rect 8264 7860 8268 7916
rect 8268 7860 8324 7916
rect 8324 7860 8328 7916
rect 8264 7856 8328 7860
rect 8344 7916 8408 7920
rect 8344 7860 8348 7916
rect 8348 7860 8404 7916
rect 8404 7860 8408 7916
rect 8344 7856 8408 7860
rect 8424 7916 8488 7920
rect 8424 7860 8428 7916
rect 8428 7860 8484 7916
rect 8484 7860 8488 7916
rect 8424 7856 8488 7860
rect 8504 7916 8568 7920
rect 8504 7860 8508 7916
rect 8508 7860 8564 7916
rect 8564 7860 8568 7916
rect 8504 7856 8568 7860
rect 8584 7916 8648 7920
rect 8584 7860 8588 7916
rect 8588 7860 8644 7916
rect 8644 7860 8648 7916
rect 8584 7856 8648 7860
rect 8664 7916 8728 7920
rect 8664 7860 8668 7916
rect 8668 7860 8724 7916
rect 8724 7860 8728 7916
rect 8664 7856 8728 7860
rect 8744 7916 8808 7920
rect 8744 7860 8748 7916
rect 8748 7860 8804 7916
rect 8804 7860 8808 7916
rect 8744 7856 8808 7860
rect 5802 7372 5866 7376
rect 5802 7316 5806 7372
rect 5806 7316 5862 7372
rect 5862 7316 5866 7372
rect 5802 7312 5866 7316
rect 5882 7372 5946 7376
rect 5882 7316 5886 7372
rect 5886 7316 5942 7372
rect 5942 7316 5946 7372
rect 5882 7312 5946 7316
rect 5962 7372 6026 7376
rect 5962 7316 5966 7372
rect 5966 7316 6022 7372
rect 6022 7316 6026 7372
rect 5962 7312 6026 7316
rect 6042 7372 6106 7376
rect 6042 7316 6046 7372
rect 6046 7316 6102 7372
rect 6102 7316 6106 7372
rect 6042 7312 6106 7316
rect 8184 6828 8248 6832
rect 8184 6772 8188 6828
rect 8188 6772 8244 6828
rect 8244 6772 8248 6828
rect 8184 6768 8248 6772
rect 8264 6828 8328 6832
rect 8264 6772 8268 6828
rect 8268 6772 8324 6828
rect 8324 6772 8328 6828
rect 8264 6768 8328 6772
rect 8344 6828 8408 6832
rect 8344 6772 8348 6828
rect 8348 6772 8404 6828
rect 8404 6772 8408 6828
rect 8344 6768 8408 6772
rect 8424 6828 8488 6832
rect 8424 6772 8428 6828
rect 8428 6772 8484 6828
rect 8484 6772 8488 6828
rect 8424 6768 8488 6772
rect 8504 6828 8568 6832
rect 8504 6772 8508 6828
rect 8508 6772 8564 6828
rect 8564 6772 8568 6828
rect 8504 6768 8568 6772
rect 8584 6828 8648 6832
rect 8584 6772 8588 6828
rect 8588 6772 8644 6828
rect 8644 6772 8648 6828
rect 8584 6768 8648 6772
rect 8664 6828 8728 6832
rect 8664 6772 8668 6828
rect 8668 6772 8724 6828
rect 8724 6772 8728 6828
rect 8664 6768 8728 6772
rect 8744 6828 8808 6832
rect 8744 6772 8748 6828
rect 8748 6772 8804 6828
rect 8804 6772 8808 6828
rect 8744 6768 8808 6772
rect 5802 6284 5866 6288
rect 5802 6228 5806 6284
rect 5806 6228 5862 6284
rect 5862 6228 5866 6284
rect 5802 6224 5866 6228
rect 5882 6284 5946 6288
rect 5882 6228 5886 6284
rect 5886 6228 5942 6284
rect 5942 6228 5946 6284
rect 5882 6224 5946 6228
rect 5962 6284 6026 6288
rect 5962 6228 5966 6284
rect 5966 6228 6022 6284
rect 6022 6228 6026 6284
rect 5962 6224 6026 6228
rect 6042 6284 6106 6288
rect 6042 6228 6046 6284
rect 6046 6228 6102 6284
rect 6102 6228 6106 6284
rect 6042 6224 6106 6228
rect 8184 5740 8248 5744
rect 8184 5684 8188 5740
rect 8188 5684 8244 5740
rect 8244 5684 8248 5740
rect 8184 5680 8248 5684
rect 8264 5740 8328 5744
rect 8264 5684 8268 5740
rect 8268 5684 8324 5740
rect 8324 5684 8328 5740
rect 8264 5680 8328 5684
rect 8344 5740 8408 5744
rect 8344 5684 8348 5740
rect 8348 5684 8404 5740
rect 8404 5684 8408 5740
rect 8344 5680 8408 5684
rect 8424 5740 8488 5744
rect 8424 5684 8428 5740
rect 8428 5684 8484 5740
rect 8484 5684 8488 5740
rect 8424 5680 8488 5684
rect 8504 5740 8568 5744
rect 8504 5684 8508 5740
rect 8508 5684 8564 5740
rect 8564 5684 8568 5740
rect 8504 5680 8568 5684
rect 8584 5740 8648 5744
rect 8584 5684 8588 5740
rect 8588 5684 8644 5740
rect 8644 5684 8648 5740
rect 8584 5680 8648 5684
rect 8664 5740 8728 5744
rect 8664 5684 8668 5740
rect 8668 5684 8724 5740
rect 8724 5684 8728 5740
rect 8664 5680 8728 5684
rect 8744 5740 8808 5744
rect 8744 5684 8748 5740
rect 8748 5684 8804 5740
rect 8804 5684 8808 5740
rect 8744 5680 8808 5684
<< metal4 >>
rect 900 19254 2532 20128
rect 900 19018 958 19254
rect 1194 19018 1278 19254
rect 1514 19018 1598 19254
rect 1834 19018 1918 19254
rect 2154 19018 2238 19254
rect 2474 19018 2532 19254
rect 900 18934 2532 19018
rect 900 18698 958 18934
rect 1194 18698 1278 18934
rect 1514 18698 1598 18934
rect 1834 18698 1918 18934
rect 2154 18698 2238 18934
rect 2474 18698 2532 18934
rect 900 18614 2532 18698
rect 900 18378 958 18614
rect 1194 18378 1278 18614
rect 1514 18378 1598 18614
rect 1834 18378 1918 18614
rect 2154 18378 2238 18614
rect 2474 18378 2532 18614
rect 900 18294 2532 18378
rect 900 18058 958 18294
rect 1194 18058 1278 18294
rect 1514 18058 1598 18294
rect 1834 18058 1918 18294
rect 2154 18058 2238 18294
rect 2474 18058 2532 18294
rect 900 17974 2532 18058
rect 900 17738 958 17974
rect 1194 17738 1278 17974
rect 1514 17738 1598 17974
rect 1834 17738 1918 17974
rect 2154 17738 2238 17974
rect 2474 17738 2532 17974
rect 900 14214 2532 17738
rect 900 13978 958 14214
rect 1194 13978 1278 14214
rect 1514 13978 1598 14214
rect 1834 13978 1918 14214
rect 2154 13978 2238 14214
rect 2474 13978 2532 14214
rect 900 13894 2532 13978
rect 900 13658 958 13894
rect 1194 13658 1278 13894
rect 1514 13658 1598 13894
rect 1834 13658 1918 13894
rect 2154 13658 2238 13894
rect 2474 13658 2532 13894
rect 900 8774 2532 13658
rect 900 8538 958 8774
rect 1194 8538 1278 8774
rect 1514 8538 1598 8774
rect 1834 8538 1918 8774
rect 2154 8538 2238 8774
rect 2474 8538 2532 8774
rect 900 8454 2532 8538
rect 900 8218 958 8454
rect 1194 8218 1278 8454
rect 1514 8218 1598 8454
rect 1834 8218 1918 8454
rect 2154 8218 2238 8454
rect 2474 8218 2532 8454
rect 900 2390 2532 8218
rect 900 2154 958 2390
rect 1194 2154 1278 2390
rect 1514 2154 1598 2390
rect 1834 2154 1918 2390
rect 2154 2154 2238 2390
rect 2474 2154 2532 2390
rect 900 2070 2532 2154
rect 900 1834 958 2070
rect 1194 1834 1278 2070
rect 1514 1834 1598 2070
rect 1834 1834 1918 2070
rect 2154 1834 2238 2070
rect 2474 1834 2532 2070
rect 900 1750 2532 1834
rect 900 1514 958 1750
rect 1194 1514 1278 1750
rect 1514 1514 1598 1750
rect 1834 1514 1918 1750
rect 2154 1514 2238 1750
rect 2474 1514 2532 1750
rect 900 1430 2532 1514
rect 900 1194 958 1430
rect 1194 1194 1278 1430
rect 1514 1194 1598 1430
rect 1834 1194 1918 1430
rect 2154 1194 2238 1430
rect 2474 1194 2532 1430
rect 900 1110 2532 1194
rect 900 874 958 1110
rect 1194 874 1278 1110
rect 1514 874 1598 1110
rect 1834 874 1918 1110
rect 2154 874 2238 1110
rect 2474 874 2532 1110
rect 900 0 2532 874
rect 3348 16806 4980 20128
rect 8160 19254 8832 19312
rect 8160 19018 8218 19254
rect 8454 19018 8538 19254
rect 8774 19018 8832 19254
rect 8160 18934 8832 19018
rect 8160 18698 8218 18934
rect 8454 18698 8538 18934
rect 8774 18698 8832 18934
rect 8160 18614 8832 18698
rect 8160 18378 8218 18614
rect 8454 18378 8538 18614
rect 8774 18378 8832 18614
rect 8160 18294 8832 18378
rect 8160 18058 8218 18294
rect 8454 18058 8538 18294
rect 8774 18058 8832 18294
rect 8160 17974 8832 18058
rect 8160 17738 8218 17974
rect 8454 17738 8538 17974
rect 8774 17738 8832 17974
rect 3348 16570 3406 16806
rect 3642 16570 3726 16806
rect 3962 16570 4046 16806
rect 4282 16570 4366 16806
rect 4602 16570 4686 16806
rect 4922 16570 4980 16806
rect 3348 16486 4980 16570
rect 3348 16250 3406 16486
rect 3642 16250 3726 16486
rect 3962 16250 4046 16486
rect 4282 16250 4366 16486
rect 4602 16250 4686 16486
rect 4922 16250 4980 16486
rect 3348 16166 4980 16250
rect 3348 15930 3406 16166
rect 3642 15930 3726 16166
rect 3962 15930 4046 16166
rect 4282 15930 4366 16166
rect 4602 15930 4686 16166
rect 4922 15930 4980 16166
rect 3348 15846 4980 15930
rect 3348 15610 3406 15846
rect 3642 15610 3726 15846
rect 3962 15610 4046 15846
rect 4282 15610 4366 15846
rect 4602 15610 4686 15846
rect 4922 15610 4980 15846
rect 3348 15526 4980 15610
rect 3348 15290 3406 15526
rect 3642 15290 3726 15526
rect 3962 15290 4046 15526
rect 4282 15290 4366 15526
rect 4602 15290 4686 15526
rect 4922 15290 4980 15526
rect 3348 11494 4980 15290
rect 3348 11258 3406 11494
rect 3642 11258 3726 11494
rect 3962 11258 4046 11494
rect 4282 11258 4366 11494
rect 4602 11258 4686 11494
rect 4922 11258 4980 11494
rect 3348 11174 4980 11258
rect 3348 10938 3406 11174
rect 3642 10938 3726 11174
rect 3962 10938 4046 11174
rect 4282 10938 4366 11174
rect 4602 10938 4686 11174
rect 4922 10938 4980 11174
rect 3348 6054 4980 10938
rect 3348 5818 3406 6054
rect 3642 5818 3726 6054
rect 3962 5818 4046 6054
rect 4282 5818 4366 6054
rect 4602 5818 4686 6054
rect 4922 5818 4980 6054
rect 3348 5734 4980 5818
rect 3348 5498 3406 5734
rect 3642 5498 3726 5734
rect 3962 5498 4046 5734
rect 4282 5498 4366 5734
rect 4602 5498 4686 5734
rect 4922 5498 4980 5734
rect 3348 4838 4980 5498
rect 3348 4602 3406 4838
rect 3642 4602 3726 4838
rect 3962 4602 4046 4838
rect 4282 4602 4366 4838
rect 4602 4602 4686 4838
rect 4922 4602 4980 4838
rect 3348 4518 4980 4602
rect 3348 4282 3406 4518
rect 3642 4282 3726 4518
rect 3962 4282 4046 4518
rect 4282 4282 4366 4518
rect 4602 4282 4686 4518
rect 4922 4282 4980 4518
rect 3348 4198 4980 4282
rect 3348 3962 3406 4198
rect 3642 3962 3726 4198
rect 3962 3962 4046 4198
rect 4282 3962 4366 4198
rect 4602 3962 4686 4198
rect 4922 3962 4980 4198
rect 3348 3878 4980 3962
rect 3348 3642 3406 3878
rect 3642 3642 3726 3878
rect 3962 3642 4046 3878
rect 4282 3642 4366 3878
rect 4602 3642 4686 3878
rect 4922 3642 4980 3878
rect 3348 3558 4980 3642
rect 3348 3322 3406 3558
rect 3642 3322 3726 3558
rect 3962 3322 4046 3558
rect 4282 3322 4366 3558
rect 4602 3322 4686 3558
rect 4922 3322 4980 3558
rect 3348 0 4980 3322
rect 5440 16806 6112 16864
rect 5440 16570 5498 16806
rect 5734 16570 5818 16806
rect 6054 16570 6112 16806
rect 5440 16486 6112 16570
rect 5440 16250 5498 16486
rect 5734 16250 5818 16486
rect 6054 16250 6112 16486
rect 5440 16166 6112 16250
rect 5440 15930 5498 16166
rect 5734 15930 5818 16166
rect 6054 15930 6112 16166
rect 5440 15846 6112 15930
rect 5440 15610 5498 15846
rect 5734 15610 5818 15846
rect 6054 15610 6112 15846
rect 5440 15526 6112 15610
rect 5440 15290 5498 15526
rect 5734 15290 5818 15526
rect 6054 15290 6112 15526
rect 5440 13904 6112 15290
rect 5440 13840 5802 13904
rect 5866 13840 5882 13904
rect 5946 13840 5962 13904
rect 6026 13840 6042 13904
rect 6106 13840 6112 13904
rect 5440 12816 6112 13840
rect 5440 12752 5802 12816
rect 5866 12752 5882 12816
rect 5946 12752 5962 12816
rect 6026 12752 6042 12816
rect 6106 12752 6112 12816
rect 5440 11728 6112 12752
rect 5440 11664 5802 11728
rect 5866 11664 5882 11728
rect 5946 11664 5962 11728
rect 6026 11664 6042 11728
rect 6106 11664 6112 11728
rect 5440 11494 6112 11664
rect 5440 11258 5498 11494
rect 5734 11258 5818 11494
rect 6054 11258 6112 11494
rect 5440 11174 6112 11258
rect 5440 10938 5498 11174
rect 5734 10938 5818 11174
rect 6054 10938 6112 11174
rect 5440 10640 6112 10938
rect 5440 10576 5802 10640
rect 5866 10576 5882 10640
rect 5946 10576 5962 10640
rect 6026 10576 6042 10640
rect 6106 10576 6112 10640
rect 5440 9552 6112 10576
rect 5440 9488 5802 9552
rect 5866 9488 5882 9552
rect 5946 9488 5962 9552
rect 6026 9488 6042 9552
rect 6106 9488 6112 9552
rect 5440 8464 6112 9488
rect 5440 8400 5802 8464
rect 5866 8400 5882 8464
rect 5946 8400 5962 8464
rect 6026 8400 6042 8464
rect 6106 8400 6112 8464
rect 5440 7376 6112 8400
rect 5440 7312 5802 7376
rect 5866 7312 5882 7376
rect 5946 7312 5962 7376
rect 6026 7312 6042 7376
rect 6106 7312 6112 7376
rect 5440 6288 6112 7312
rect 5440 6224 5802 6288
rect 5866 6224 5882 6288
rect 5946 6224 5962 6288
rect 6026 6224 6042 6288
rect 6106 6224 6112 6288
rect 5440 6054 6112 6224
rect 5440 5818 5498 6054
rect 5734 5818 5818 6054
rect 6054 5818 6112 6054
rect 5440 5734 6112 5818
rect 5440 5498 5498 5734
rect 5734 5498 5818 5734
rect 6054 5498 6112 5734
rect 5440 4838 6112 5498
rect 5440 4602 5498 4838
rect 5734 4602 5818 4838
rect 6054 4602 6112 4838
rect 5440 4518 6112 4602
rect 5440 4282 5498 4518
rect 5734 4282 5818 4518
rect 6054 4282 6112 4518
rect 5440 4198 6112 4282
rect 5440 3962 5498 4198
rect 5734 3962 5818 4198
rect 6054 3962 6112 4198
rect 5440 3878 6112 3962
rect 5440 3642 5498 3878
rect 5734 3642 5818 3878
rect 6054 3642 6112 3878
rect 5440 3558 6112 3642
rect 5440 3322 5498 3558
rect 5734 3322 5818 3558
rect 6054 3322 6112 3558
rect 5440 3264 6112 3322
rect 8160 14448 8832 17738
rect 8160 14384 8184 14448
rect 8248 14384 8264 14448
rect 8328 14384 8344 14448
rect 8408 14384 8424 14448
rect 8488 14384 8504 14448
rect 8568 14384 8584 14448
rect 8648 14384 8664 14448
rect 8728 14384 8744 14448
rect 8808 14384 8832 14448
rect 8160 14214 8832 14384
rect 8160 13978 8218 14214
rect 8454 13978 8538 14214
rect 8774 13978 8832 14214
rect 8160 13894 8832 13978
rect 8160 13658 8218 13894
rect 8454 13658 8538 13894
rect 8774 13658 8832 13894
rect 8160 13360 8832 13658
rect 8160 13296 8184 13360
rect 8248 13296 8264 13360
rect 8328 13296 8344 13360
rect 8408 13296 8424 13360
rect 8488 13296 8504 13360
rect 8568 13296 8584 13360
rect 8648 13296 8664 13360
rect 8728 13296 8744 13360
rect 8808 13296 8832 13360
rect 8160 12272 8832 13296
rect 8160 12208 8184 12272
rect 8248 12208 8264 12272
rect 8328 12208 8344 12272
rect 8408 12208 8424 12272
rect 8488 12208 8504 12272
rect 8568 12208 8584 12272
rect 8648 12208 8664 12272
rect 8728 12208 8744 12272
rect 8808 12208 8832 12272
rect 8160 11184 8832 12208
rect 8160 11120 8184 11184
rect 8248 11120 8264 11184
rect 8328 11120 8344 11184
rect 8408 11120 8424 11184
rect 8488 11120 8504 11184
rect 8568 11120 8584 11184
rect 8648 11120 8664 11184
rect 8728 11120 8744 11184
rect 8808 11120 8832 11184
rect 8160 10096 8832 11120
rect 8160 10032 8184 10096
rect 8248 10032 8264 10096
rect 8328 10032 8344 10096
rect 8408 10032 8424 10096
rect 8488 10032 8504 10096
rect 8568 10032 8584 10096
rect 8648 10032 8664 10096
rect 8728 10032 8744 10096
rect 8808 10032 8832 10096
rect 8160 9008 8832 10032
rect 8160 8944 8184 9008
rect 8248 8944 8264 9008
rect 8328 8944 8344 9008
rect 8408 8944 8424 9008
rect 8488 8944 8504 9008
rect 8568 8944 8584 9008
rect 8648 8944 8664 9008
rect 8728 8944 8744 9008
rect 8808 8944 8832 9008
rect 8160 8774 8832 8944
rect 8160 8538 8218 8774
rect 8454 8538 8538 8774
rect 8774 8538 8832 8774
rect 8160 8454 8832 8538
rect 8160 8218 8218 8454
rect 8454 8218 8538 8454
rect 8774 8218 8832 8454
rect 8160 7920 8832 8218
rect 8160 7856 8184 7920
rect 8248 7856 8264 7920
rect 8328 7856 8344 7920
rect 8408 7856 8424 7920
rect 8488 7856 8504 7920
rect 8568 7856 8584 7920
rect 8648 7856 8664 7920
rect 8728 7856 8744 7920
rect 8808 7856 8832 7920
rect 8160 6832 8832 7856
rect 8160 6768 8184 6832
rect 8248 6768 8264 6832
rect 8328 6768 8344 6832
rect 8408 6768 8424 6832
rect 8488 6768 8504 6832
rect 8568 6768 8584 6832
rect 8648 6768 8664 6832
rect 8728 6768 8744 6832
rect 8808 6768 8832 6832
rect 8160 5744 8832 6768
rect 8160 5680 8184 5744
rect 8248 5680 8264 5744
rect 8328 5680 8344 5744
rect 8408 5680 8424 5744
rect 8488 5680 8504 5744
rect 8568 5680 8584 5744
rect 8648 5680 8664 5744
rect 8728 5680 8744 5744
rect 8808 5680 8832 5744
rect 8160 2390 8832 5680
rect 8160 2154 8218 2390
rect 8454 2154 8538 2390
rect 8774 2154 8832 2390
rect 8160 2070 8832 2154
rect 8160 1834 8218 2070
rect 8454 1834 8538 2070
rect 8774 1834 8832 2070
rect 8160 1750 8832 1834
rect 8160 1514 8218 1750
rect 8454 1514 8538 1750
rect 8774 1514 8832 1750
rect 8160 1430 8832 1514
rect 8160 1194 8218 1430
rect 8454 1194 8538 1430
rect 8774 1194 8832 1430
rect 8160 1110 8832 1194
rect 8160 874 8218 1110
rect 8454 874 8538 1110
rect 8774 874 8832 1110
rect 8160 816 8832 874
rect 11120 16806 12752 20128
rect 11120 16570 11178 16806
rect 11414 16570 11498 16806
rect 11734 16570 11818 16806
rect 12054 16570 12138 16806
rect 12374 16570 12458 16806
rect 12694 16570 12752 16806
rect 11120 16486 12752 16570
rect 11120 16250 11178 16486
rect 11414 16250 11498 16486
rect 11734 16250 11818 16486
rect 12054 16250 12138 16486
rect 12374 16250 12458 16486
rect 12694 16250 12752 16486
rect 11120 16166 12752 16250
rect 11120 15930 11178 16166
rect 11414 15930 11498 16166
rect 11734 15930 11818 16166
rect 12054 15930 12138 16166
rect 12374 15930 12458 16166
rect 12694 15930 12752 16166
rect 11120 15846 12752 15930
rect 11120 15610 11178 15846
rect 11414 15610 11498 15846
rect 11734 15610 11818 15846
rect 12054 15610 12138 15846
rect 12374 15610 12458 15846
rect 12694 15610 12752 15846
rect 11120 15526 12752 15610
rect 11120 15290 11178 15526
rect 11414 15290 11498 15526
rect 11734 15290 11818 15526
rect 12054 15290 12138 15526
rect 12374 15290 12458 15526
rect 12694 15290 12752 15526
rect 11120 11494 12752 15290
rect 11120 11258 11178 11494
rect 11414 11258 11498 11494
rect 11734 11258 11818 11494
rect 12054 11258 12138 11494
rect 12374 11258 12458 11494
rect 12694 11258 12752 11494
rect 11120 11174 12752 11258
rect 11120 10938 11178 11174
rect 11414 10938 11498 11174
rect 11734 10938 11818 11174
rect 12054 10938 12138 11174
rect 12374 10938 12458 11174
rect 12694 10938 12752 11174
rect 11120 6054 12752 10938
rect 11120 5818 11178 6054
rect 11414 5818 11498 6054
rect 11734 5818 11818 6054
rect 12054 5818 12138 6054
rect 12374 5818 12458 6054
rect 12694 5818 12752 6054
rect 11120 5734 12752 5818
rect 11120 5498 11178 5734
rect 11414 5498 11498 5734
rect 11734 5498 11818 5734
rect 12054 5498 12138 5734
rect 12374 5498 12458 5734
rect 12694 5498 12752 5734
rect 11120 4838 12752 5498
rect 11120 4602 11178 4838
rect 11414 4602 11498 4838
rect 11734 4602 11818 4838
rect 12054 4602 12138 4838
rect 12374 4602 12458 4838
rect 12694 4602 12752 4838
rect 11120 4518 12752 4602
rect 11120 4282 11178 4518
rect 11414 4282 11498 4518
rect 11734 4282 11818 4518
rect 12054 4282 12138 4518
rect 12374 4282 12458 4518
rect 12694 4282 12752 4518
rect 11120 4198 12752 4282
rect 11120 3962 11178 4198
rect 11414 3962 11498 4198
rect 11734 3962 11818 4198
rect 12054 3962 12138 4198
rect 12374 3962 12458 4198
rect 12694 3962 12752 4198
rect 11120 3878 12752 3962
rect 11120 3642 11178 3878
rect 11414 3642 11498 3878
rect 11734 3642 11818 3878
rect 12054 3642 12138 3878
rect 12374 3642 12458 3878
rect 12694 3642 12752 3878
rect 11120 3558 12752 3642
rect 11120 3322 11178 3558
rect 11414 3322 11498 3558
rect 11734 3322 11818 3558
rect 12054 3322 12138 3558
rect 12374 3322 12458 3558
rect 12694 3322 12752 3558
rect 11120 0 12752 3322
rect 13568 19254 15200 20128
rect 13568 19018 13626 19254
rect 13862 19018 13946 19254
rect 14182 19018 14266 19254
rect 14502 19018 14586 19254
rect 14822 19018 14906 19254
rect 15142 19018 15200 19254
rect 13568 18934 15200 19018
rect 13568 18698 13626 18934
rect 13862 18698 13946 18934
rect 14182 18698 14266 18934
rect 14502 18698 14586 18934
rect 14822 18698 14906 18934
rect 15142 18698 15200 18934
rect 13568 18614 15200 18698
rect 13568 18378 13626 18614
rect 13862 18378 13946 18614
rect 14182 18378 14266 18614
rect 14502 18378 14586 18614
rect 14822 18378 14906 18614
rect 15142 18378 15200 18614
rect 13568 18294 15200 18378
rect 13568 18058 13626 18294
rect 13862 18058 13946 18294
rect 14182 18058 14266 18294
rect 14502 18058 14586 18294
rect 14822 18058 14906 18294
rect 15142 18058 15200 18294
rect 13568 17974 15200 18058
rect 13568 17738 13626 17974
rect 13862 17738 13946 17974
rect 14182 17738 14266 17974
rect 14502 17738 14586 17974
rect 14822 17738 14906 17974
rect 15142 17738 15200 17974
rect 13568 14214 15200 17738
rect 13568 13978 13626 14214
rect 13862 13978 13946 14214
rect 14182 13978 14266 14214
rect 14502 13978 14586 14214
rect 14822 13978 14906 14214
rect 15142 13978 15200 14214
rect 13568 13894 15200 13978
rect 13568 13658 13626 13894
rect 13862 13658 13946 13894
rect 14182 13658 14266 13894
rect 14502 13658 14586 13894
rect 14822 13658 14906 13894
rect 15142 13658 15200 13894
rect 13568 8774 15200 13658
rect 13568 8538 13626 8774
rect 13862 8538 13946 8774
rect 14182 8538 14266 8774
rect 14502 8538 14586 8774
rect 14822 8538 14906 8774
rect 15142 8538 15200 8774
rect 13568 8454 15200 8538
rect 13568 8218 13626 8454
rect 13862 8218 13946 8454
rect 14182 8218 14266 8454
rect 14502 8218 14586 8454
rect 14822 8218 14906 8454
rect 15142 8218 15200 8454
rect 13568 2390 15200 8218
rect 13568 2154 13626 2390
rect 13862 2154 13946 2390
rect 14182 2154 14266 2390
rect 14502 2154 14586 2390
rect 14822 2154 14906 2390
rect 15142 2154 15200 2390
rect 13568 2070 15200 2154
rect 13568 1834 13626 2070
rect 13862 1834 13946 2070
rect 14182 1834 14266 2070
rect 14502 1834 14586 2070
rect 14822 1834 14906 2070
rect 15142 1834 15200 2070
rect 13568 1750 15200 1834
rect 13568 1514 13626 1750
rect 13862 1514 13946 1750
rect 14182 1514 14266 1750
rect 14502 1514 14586 1750
rect 14822 1514 14906 1750
rect 15142 1514 15200 1750
rect 13568 1430 15200 1514
rect 13568 1194 13626 1430
rect 13862 1194 13946 1430
rect 14182 1194 14266 1430
rect 14502 1194 14586 1430
rect 14822 1194 14906 1430
rect 15142 1194 15200 1430
rect 13568 1110 15200 1194
rect 13568 874 13626 1110
rect 13862 874 13946 1110
rect 14182 874 14266 1110
rect 14502 874 14586 1110
rect 14822 874 14906 1110
rect 15142 874 15200 1110
rect 13568 0 15200 874
<< via4 >>
rect 958 19018 1194 19254
rect 1278 19018 1514 19254
rect 1598 19018 1834 19254
rect 1918 19018 2154 19254
rect 2238 19018 2474 19254
rect 958 18698 1194 18934
rect 1278 18698 1514 18934
rect 1598 18698 1834 18934
rect 1918 18698 2154 18934
rect 2238 18698 2474 18934
rect 958 18378 1194 18614
rect 1278 18378 1514 18614
rect 1598 18378 1834 18614
rect 1918 18378 2154 18614
rect 2238 18378 2474 18614
rect 958 18058 1194 18294
rect 1278 18058 1514 18294
rect 1598 18058 1834 18294
rect 1918 18058 2154 18294
rect 2238 18058 2474 18294
rect 958 17738 1194 17974
rect 1278 17738 1514 17974
rect 1598 17738 1834 17974
rect 1918 17738 2154 17974
rect 2238 17738 2474 17974
rect 958 13978 1194 14214
rect 1278 13978 1514 14214
rect 1598 13978 1834 14214
rect 1918 13978 2154 14214
rect 2238 13978 2474 14214
rect 958 13658 1194 13894
rect 1278 13658 1514 13894
rect 1598 13658 1834 13894
rect 1918 13658 2154 13894
rect 2238 13658 2474 13894
rect 958 8538 1194 8774
rect 1278 8538 1514 8774
rect 1598 8538 1834 8774
rect 1918 8538 2154 8774
rect 2238 8538 2474 8774
rect 958 8218 1194 8454
rect 1278 8218 1514 8454
rect 1598 8218 1834 8454
rect 1918 8218 2154 8454
rect 2238 8218 2474 8454
rect 958 2154 1194 2390
rect 1278 2154 1514 2390
rect 1598 2154 1834 2390
rect 1918 2154 2154 2390
rect 2238 2154 2474 2390
rect 958 1834 1194 2070
rect 1278 1834 1514 2070
rect 1598 1834 1834 2070
rect 1918 1834 2154 2070
rect 2238 1834 2474 2070
rect 958 1514 1194 1750
rect 1278 1514 1514 1750
rect 1598 1514 1834 1750
rect 1918 1514 2154 1750
rect 2238 1514 2474 1750
rect 958 1194 1194 1430
rect 1278 1194 1514 1430
rect 1598 1194 1834 1430
rect 1918 1194 2154 1430
rect 2238 1194 2474 1430
rect 958 874 1194 1110
rect 1278 874 1514 1110
rect 1598 874 1834 1110
rect 1918 874 2154 1110
rect 2238 874 2474 1110
rect 8218 19018 8454 19254
rect 8538 19018 8774 19254
rect 8218 18698 8454 18934
rect 8538 18698 8774 18934
rect 8218 18378 8454 18614
rect 8538 18378 8774 18614
rect 8218 18058 8454 18294
rect 8538 18058 8774 18294
rect 8218 17738 8454 17974
rect 8538 17738 8774 17974
rect 3406 16570 3642 16806
rect 3726 16570 3962 16806
rect 4046 16570 4282 16806
rect 4366 16570 4602 16806
rect 4686 16570 4922 16806
rect 3406 16250 3642 16486
rect 3726 16250 3962 16486
rect 4046 16250 4282 16486
rect 4366 16250 4602 16486
rect 4686 16250 4922 16486
rect 3406 15930 3642 16166
rect 3726 15930 3962 16166
rect 4046 15930 4282 16166
rect 4366 15930 4602 16166
rect 4686 15930 4922 16166
rect 3406 15610 3642 15846
rect 3726 15610 3962 15846
rect 4046 15610 4282 15846
rect 4366 15610 4602 15846
rect 4686 15610 4922 15846
rect 3406 15290 3642 15526
rect 3726 15290 3962 15526
rect 4046 15290 4282 15526
rect 4366 15290 4602 15526
rect 4686 15290 4922 15526
rect 3406 11258 3642 11494
rect 3726 11258 3962 11494
rect 4046 11258 4282 11494
rect 4366 11258 4602 11494
rect 4686 11258 4922 11494
rect 3406 10938 3642 11174
rect 3726 10938 3962 11174
rect 4046 10938 4282 11174
rect 4366 10938 4602 11174
rect 4686 10938 4922 11174
rect 3406 5818 3642 6054
rect 3726 5818 3962 6054
rect 4046 5818 4282 6054
rect 4366 5818 4602 6054
rect 4686 5818 4922 6054
rect 3406 5498 3642 5734
rect 3726 5498 3962 5734
rect 4046 5498 4282 5734
rect 4366 5498 4602 5734
rect 4686 5498 4922 5734
rect 3406 4602 3642 4838
rect 3726 4602 3962 4838
rect 4046 4602 4282 4838
rect 4366 4602 4602 4838
rect 4686 4602 4922 4838
rect 3406 4282 3642 4518
rect 3726 4282 3962 4518
rect 4046 4282 4282 4518
rect 4366 4282 4602 4518
rect 4686 4282 4922 4518
rect 3406 3962 3642 4198
rect 3726 3962 3962 4198
rect 4046 3962 4282 4198
rect 4366 3962 4602 4198
rect 4686 3962 4922 4198
rect 3406 3642 3642 3878
rect 3726 3642 3962 3878
rect 4046 3642 4282 3878
rect 4366 3642 4602 3878
rect 4686 3642 4922 3878
rect 3406 3322 3642 3558
rect 3726 3322 3962 3558
rect 4046 3322 4282 3558
rect 4366 3322 4602 3558
rect 4686 3322 4922 3558
rect 5498 16570 5734 16806
rect 5818 16570 6054 16806
rect 5498 16250 5734 16486
rect 5818 16250 6054 16486
rect 5498 15930 5734 16166
rect 5818 15930 6054 16166
rect 5498 15610 5734 15846
rect 5818 15610 6054 15846
rect 5498 15290 5734 15526
rect 5818 15290 6054 15526
rect 5498 11258 5734 11494
rect 5818 11258 6054 11494
rect 5498 10938 5734 11174
rect 5818 10938 6054 11174
rect 5498 5818 5734 6054
rect 5818 5818 6054 6054
rect 5498 5498 5734 5734
rect 5818 5498 6054 5734
rect 5498 4602 5734 4838
rect 5818 4602 6054 4838
rect 5498 4282 5734 4518
rect 5818 4282 6054 4518
rect 5498 3962 5734 4198
rect 5818 3962 6054 4198
rect 5498 3642 5734 3878
rect 5818 3642 6054 3878
rect 5498 3322 5734 3558
rect 5818 3322 6054 3558
rect 8218 13978 8454 14214
rect 8538 13978 8774 14214
rect 8218 13658 8454 13894
rect 8538 13658 8774 13894
rect 8218 8538 8454 8774
rect 8538 8538 8774 8774
rect 8218 8218 8454 8454
rect 8538 8218 8774 8454
rect 8218 2154 8454 2390
rect 8538 2154 8774 2390
rect 8218 1834 8454 2070
rect 8538 1834 8774 2070
rect 8218 1514 8454 1750
rect 8538 1514 8774 1750
rect 8218 1194 8454 1430
rect 8538 1194 8774 1430
rect 8218 874 8454 1110
rect 8538 874 8774 1110
rect 11178 16570 11414 16806
rect 11498 16570 11734 16806
rect 11818 16570 12054 16806
rect 12138 16570 12374 16806
rect 12458 16570 12694 16806
rect 11178 16250 11414 16486
rect 11498 16250 11734 16486
rect 11818 16250 12054 16486
rect 12138 16250 12374 16486
rect 12458 16250 12694 16486
rect 11178 15930 11414 16166
rect 11498 15930 11734 16166
rect 11818 15930 12054 16166
rect 12138 15930 12374 16166
rect 12458 15930 12694 16166
rect 11178 15610 11414 15846
rect 11498 15610 11734 15846
rect 11818 15610 12054 15846
rect 12138 15610 12374 15846
rect 12458 15610 12694 15846
rect 11178 15290 11414 15526
rect 11498 15290 11734 15526
rect 11818 15290 12054 15526
rect 12138 15290 12374 15526
rect 12458 15290 12694 15526
rect 11178 11258 11414 11494
rect 11498 11258 11734 11494
rect 11818 11258 12054 11494
rect 12138 11258 12374 11494
rect 12458 11258 12694 11494
rect 11178 10938 11414 11174
rect 11498 10938 11734 11174
rect 11818 10938 12054 11174
rect 12138 10938 12374 11174
rect 12458 10938 12694 11174
rect 11178 5818 11414 6054
rect 11498 5818 11734 6054
rect 11818 5818 12054 6054
rect 12138 5818 12374 6054
rect 12458 5818 12694 6054
rect 11178 5498 11414 5734
rect 11498 5498 11734 5734
rect 11818 5498 12054 5734
rect 12138 5498 12374 5734
rect 12458 5498 12694 5734
rect 11178 4602 11414 4838
rect 11498 4602 11734 4838
rect 11818 4602 12054 4838
rect 12138 4602 12374 4838
rect 12458 4602 12694 4838
rect 11178 4282 11414 4518
rect 11498 4282 11734 4518
rect 11818 4282 12054 4518
rect 12138 4282 12374 4518
rect 12458 4282 12694 4518
rect 11178 3962 11414 4198
rect 11498 3962 11734 4198
rect 11818 3962 12054 4198
rect 12138 3962 12374 4198
rect 12458 3962 12694 4198
rect 11178 3642 11414 3878
rect 11498 3642 11734 3878
rect 11818 3642 12054 3878
rect 12138 3642 12374 3878
rect 12458 3642 12694 3878
rect 11178 3322 11414 3558
rect 11498 3322 11734 3558
rect 11818 3322 12054 3558
rect 12138 3322 12374 3558
rect 12458 3322 12694 3558
rect 13626 19018 13862 19254
rect 13946 19018 14182 19254
rect 14266 19018 14502 19254
rect 14586 19018 14822 19254
rect 14906 19018 15142 19254
rect 13626 18698 13862 18934
rect 13946 18698 14182 18934
rect 14266 18698 14502 18934
rect 14586 18698 14822 18934
rect 14906 18698 15142 18934
rect 13626 18378 13862 18614
rect 13946 18378 14182 18614
rect 14266 18378 14502 18614
rect 14586 18378 14822 18614
rect 14906 18378 15142 18614
rect 13626 18058 13862 18294
rect 13946 18058 14182 18294
rect 14266 18058 14502 18294
rect 14586 18058 14822 18294
rect 14906 18058 15142 18294
rect 13626 17738 13862 17974
rect 13946 17738 14182 17974
rect 14266 17738 14502 17974
rect 14586 17738 14822 17974
rect 14906 17738 15142 17974
rect 13626 13978 13862 14214
rect 13946 13978 14182 14214
rect 14266 13978 14502 14214
rect 14586 13978 14822 14214
rect 14906 13978 15142 14214
rect 13626 13658 13862 13894
rect 13946 13658 14182 13894
rect 14266 13658 14502 13894
rect 14586 13658 14822 13894
rect 14906 13658 15142 13894
rect 13626 8538 13862 8774
rect 13946 8538 14182 8774
rect 14266 8538 14502 8774
rect 14586 8538 14822 8774
rect 14906 8538 15142 8774
rect 13626 8218 13862 8454
rect 13946 8218 14182 8454
rect 14266 8218 14502 8454
rect 14586 8218 14822 8454
rect 14906 8218 15142 8454
rect 13626 2154 13862 2390
rect 13946 2154 14182 2390
rect 14266 2154 14502 2390
rect 14586 2154 14822 2390
rect 14906 2154 15142 2390
rect 13626 1834 13862 2070
rect 13946 1834 14182 2070
rect 14266 1834 14502 2070
rect 14586 1834 14822 2070
rect 14906 1834 15142 2070
rect 13626 1514 13862 1750
rect 13946 1514 14182 1750
rect 14266 1514 14502 1750
rect 14586 1514 14822 1750
rect 14906 1514 15142 1750
rect 13626 1194 13862 1430
rect 13946 1194 14182 1430
rect 14266 1194 14502 1430
rect 14586 1194 14822 1430
rect 14906 1194 15142 1430
rect 13626 874 13862 1110
rect 13946 874 14182 1110
rect 14266 874 14502 1110
rect 14586 874 14822 1110
rect 14906 874 15142 1110
<< metal5 >>
rect 0 19254 16100 19312
rect 0 19018 958 19254
rect 1194 19018 1278 19254
rect 1514 19018 1598 19254
rect 1834 19018 1918 19254
rect 2154 19018 2238 19254
rect 2474 19018 8218 19254
rect 8454 19018 8538 19254
rect 8774 19018 13626 19254
rect 13862 19018 13946 19254
rect 14182 19018 14266 19254
rect 14502 19018 14586 19254
rect 14822 19018 14906 19254
rect 15142 19018 16100 19254
rect 0 18934 16100 19018
rect 0 18698 958 18934
rect 1194 18698 1278 18934
rect 1514 18698 1598 18934
rect 1834 18698 1918 18934
rect 2154 18698 2238 18934
rect 2474 18698 8218 18934
rect 8454 18698 8538 18934
rect 8774 18698 13626 18934
rect 13862 18698 13946 18934
rect 14182 18698 14266 18934
rect 14502 18698 14586 18934
rect 14822 18698 14906 18934
rect 15142 18698 16100 18934
rect 0 18614 16100 18698
rect 0 18378 958 18614
rect 1194 18378 1278 18614
rect 1514 18378 1598 18614
rect 1834 18378 1918 18614
rect 2154 18378 2238 18614
rect 2474 18378 8218 18614
rect 8454 18378 8538 18614
rect 8774 18378 13626 18614
rect 13862 18378 13946 18614
rect 14182 18378 14266 18614
rect 14502 18378 14586 18614
rect 14822 18378 14906 18614
rect 15142 18378 16100 18614
rect 0 18294 16100 18378
rect 0 18058 958 18294
rect 1194 18058 1278 18294
rect 1514 18058 1598 18294
rect 1834 18058 1918 18294
rect 2154 18058 2238 18294
rect 2474 18058 8218 18294
rect 8454 18058 8538 18294
rect 8774 18058 13626 18294
rect 13862 18058 13946 18294
rect 14182 18058 14266 18294
rect 14502 18058 14586 18294
rect 14822 18058 14906 18294
rect 15142 18058 16100 18294
rect 0 17974 16100 18058
rect 0 17738 958 17974
rect 1194 17738 1278 17974
rect 1514 17738 1598 17974
rect 1834 17738 1918 17974
rect 2154 17738 2238 17974
rect 2474 17738 8218 17974
rect 8454 17738 8538 17974
rect 8774 17738 13626 17974
rect 13862 17738 13946 17974
rect 14182 17738 14266 17974
rect 14502 17738 14586 17974
rect 14822 17738 14906 17974
rect 15142 17738 16100 17974
rect 0 17680 16100 17738
rect 0 16806 16100 16864
rect 0 16570 3406 16806
rect 3642 16570 3726 16806
rect 3962 16570 4046 16806
rect 4282 16570 4366 16806
rect 4602 16570 4686 16806
rect 4922 16570 5498 16806
rect 5734 16570 5818 16806
rect 6054 16570 11178 16806
rect 11414 16570 11498 16806
rect 11734 16570 11818 16806
rect 12054 16570 12138 16806
rect 12374 16570 12458 16806
rect 12694 16570 16100 16806
rect 0 16486 16100 16570
rect 0 16250 3406 16486
rect 3642 16250 3726 16486
rect 3962 16250 4046 16486
rect 4282 16250 4366 16486
rect 4602 16250 4686 16486
rect 4922 16250 5498 16486
rect 5734 16250 5818 16486
rect 6054 16250 11178 16486
rect 11414 16250 11498 16486
rect 11734 16250 11818 16486
rect 12054 16250 12138 16486
rect 12374 16250 12458 16486
rect 12694 16250 16100 16486
rect 0 16166 16100 16250
rect 0 15930 3406 16166
rect 3642 15930 3726 16166
rect 3962 15930 4046 16166
rect 4282 15930 4366 16166
rect 4602 15930 4686 16166
rect 4922 15930 5498 16166
rect 5734 15930 5818 16166
rect 6054 15930 11178 16166
rect 11414 15930 11498 16166
rect 11734 15930 11818 16166
rect 12054 15930 12138 16166
rect 12374 15930 12458 16166
rect 12694 15930 16100 16166
rect 0 15846 16100 15930
rect 0 15610 3406 15846
rect 3642 15610 3726 15846
rect 3962 15610 4046 15846
rect 4282 15610 4366 15846
rect 4602 15610 4686 15846
rect 4922 15610 5498 15846
rect 5734 15610 5818 15846
rect 6054 15610 11178 15846
rect 11414 15610 11498 15846
rect 11734 15610 11818 15846
rect 12054 15610 12138 15846
rect 12374 15610 12458 15846
rect 12694 15610 16100 15846
rect 0 15526 16100 15610
rect 0 15290 3406 15526
rect 3642 15290 3726 15526
rect 3962 15290 4046 15526
rect 4282 15290 4366 15526
rect 4602 15290 4686 15526
rect 4922 15290 5498 15526
rect 5734 15290 5818 15526
rect 6054 15290 11178 15526
rect 11414 15290 11498 15526
rect 11734 15290 11818 15526
rect 12054 15290 12138 15526
rect 12374 15290 12458 15526
rect 12694 15290 16100 15526
rect 0 15232 16100 15290
rect 900 14214 15200 14272
rect 900 13978 958 14214
rect 1194 13978 1278 14214
rect 1514 13978 1598 14214
rect 1834 13978 1918 14214
rect 2154 13978 2238 14214
rect 2474 13978 8218 14214
rect 8454 13978 8538 14214
rect 8774 13978 13626 14214
rect 13862 13978 13946 14214
rect 14182 13978 14266 14214
rect 14502 13978 14586 14214
rect 14822 13978 14906 14214
rect 15142 13978 15200 14214
rect 900 13894 15200 13978
rect 900 13658 958 13894
rect 1194 13658 1278 13894
rect 1514 13658 1598 13894
rect 1834 13658 1918 13894
rect 2154 13658 2238 13894
rect 2474 13658 8218 13894
rect 8454 13658 8538 13894
rect 8774 13658 13626 13894
rect 13862 13658 13946 13894
rect 14182 13658 14266 13894
rect 14502 13658 14586 13894
rect 14822 13658 14906 13894
rect 15142 13658 15200 13894
rect 900 13600 15200 13658
rect 3348 11494 12752 11552
rect 3348 11258 3406 11494
rect 3642 11258 3726 11494
rect 3962 11258 4046 11494
rect 4282 11258 4366 11494
rect 4602 11258 4686 11494
rect 4922 11258 5498 11494
rect 5734 11258 5818 11494
rect 6054 11258 11178 11494
rect 11414 11258 11498 11494
rect 11734 11258 11818 11494
rect 12054 11258 12138 11494
rect 12374 11258 12458 11494
rect 12694 11258 12752 11494
rect 3348 11174 12752 11258
rect 3348 10938 3406 11174
rect 3642 10938 3726 11174
rect 3962 10938 4046 11174
rect 4282 10938 4366 11174
rect 4602 10938 4686 11174
rect 4922 10938 5498 11174
rect 5734 10938 5818 11174
rect 6054 10938 11178 11174
rect 11414 10938 11498 11174
rect 11734 10938 11818 11174
rect 12054 10938 12138 11174
rect 12374 10938 12458 11174
rect 12694 10938 12752 11174
rect 3348 10880 12752 10938
rect 900 8774 15200 8832
rect 900 8538 958 8774
rect 1194 8538 1278 8774
rect 1514 8538 1598 8774
rect 1834 8538 1918 8774
rect 2154 8538 2238 8774
rect 2474 8538 8218 8774
rect 8454 8538 8538 8774
rect 8774 8538 13626 8774
rect 13862 8538 13946 8774
rect 14182 8538 14266 8774
rect 14502 8538 14586 8774
rect 14822 8538 14906 8774
rect 15142 8538 15200 8774
rect 900 8454 15200 8538
rect 900 8218 958 8454
rect 1194 8218 1278 8454
rect 1514 8218 1598 8454
rect 1834 8218 1918 8454
rect 2154 8218 2238 8454
rect 2474 8218 8218 8454
rect 8454 8218 8538 8454
rect 8774 8218 13626 8454
rect 13862 8218 13946 8454
rect 14182 8218 14266 8454
rect 14502 8218 14586 8454
rect 14822 8218 14906 8454
rect 15142 8218 15200 8454
rect 900 8160 15200 8218
rect 3348 6054 12752 6112
rect 3348 5818 3406 6054
rect 3642 5818 3726 6054
rect 3962 5818 4046 6054
rect 4282 5818 4366 6054
rect 4602 5818 4686 6054
rect 4922 5818 5498 6054
rect 5734 5818 5818 6054
rect 6054 5818 11178 6054
rect 11414 5818 11498 6054
rect 11734 5818 11818 6054
rect 12054 5818 12138 6054
rect 12374 5818 12458 6054
rect 12694 5818 12752 6054
rect 3348 5734 12752 5818
rect 3348 5498 3406 5734
rect 3642 5498 3726 5734
rect 3962 5498 4046 5734
rect 4282 5498 4366 5734
rect 4602 5498 4686 5734
rect 4922 5498 5498 5734
rect 5734 5498 5818 5734
rect 6054 5498 11178 5734
rect 11414 5498 11498 5734
rect 11734 5498 11818 5734
rect 12054 5498 12138 5734
rect 12374 5498 12458 5734
rect 12694 5498 12752 5734
rect 3348 5440 12752 5498
rect 0 4838 16100 4896
rect 0 4602 3406 4838
rect 3642 4602 3726 4838
rect 3962 4602 4046 4838
rect 4282 4602 4366 4838
rect 4602 4602 4686 4838
rect 4922 4602 5498 4838
rect 5734 4602 5818 4838
rect 6054 4602 11178 4838
rect 11414 4602 11498 4838
rect 11734 4602 11818 4838
rect 12054 4602 12138 4838
rect 12374 4602 12458 4838
rect 12694 4602 16100 4838
rect 0 4518 16100 4602
rect 0 4282 3406 4518
rect 3642 4282 3726 4518
rect 3962 4282 4046 4518
rect 4282 4282 4366 4518
rect 4602 4282 4686 4518
rect 4922 4282 5498 4518
rect 5734 4282 5818 4518
rect 6054 4282 11178 4518
rect 11414 4282 11498 4518
rect 11734 4282 11818 4518
rect 12054 4282 12138 4518
rect 12374 4282 12458 4518
rect 12694 4282 16100 4518
rect 0 4198 16100 4282
rect 0 3962 3406 4198
rect 3642 3962 3726 4198
rect 3962 3962 4046 4198
rect 4282 3962 4366 4198
rect 4602 3962 4686 4198
rect 4922 3962 5498 4198
rect 5734 3962 5818 4198
rect 6054 3962 11178 4198
rect 11414 3962 11498 4198
rect 11734 3962 11818 4198
rect 12054 3962 12138 4198
rect 12374 3962 12458 4198
rect 12694 3962 16100 4198
rect 0 3878 16100 3962
rect 0 3642 3406 3878
rect 3642 3642 3726 3878
rect 3962 3642 4046 3878
rect 4282 3642 4366 3878
rect 4602 3642 4686 3878
rect 4922 3642 5498 3878
rect 5734 3642 5818 3878
rect 6054 3642 11178 3878
rect 11414 3642 11498 3878
rect 11734 3642 11818 3878
rect 12054 3642 12138 3878
rect 12374 3642 12458 3878
rect 12694 3642 16100 3878
rect 0 3558 16100 3642
rect 0 3322 3406 3558
rect 3642 3322 3726 3558
rect 3962 3322 4046 3558
rect 4282 3322 4366 3558
rect 4602 3322 4686 3558
rect 4922 3322 5498 3558
rect 5734 3322 5818 3558
rect 6054 3322 11178 3558
rect 11414 3322 11498 3558
rect 11734 3322 11818 3558
rect 12054 3322 12138 3558
rect 12374 3322 12458 3558
rect 12694 3322 16100 3558
rect 0 3264 16100 3322
rect 0 2390 16100 2448
rect 0 2154 958 2390
rect 1194 2154 1278 2390
rect 1514 2154 1598 2390
rect 1834 2154 1918 2390
rect 2154 2154 2238 2390
rect 2474 2154 8218 2390
rect 8454 2154 8538 2390
rect 8774 2154 13626 2390
rect 13862 2154 13946 2390
rect 14182 2154 14266 2390
rect 14502 2154 14586 2390
rect 14822 2154 14906 2390
rect 15142 2154 16100 2390
rect 0 2070 16100 2154
rect 0 1834 958 2070
rect 1194 1834 1278 2070
rect 1514 1834 1598 2070
rect 1834 1834 1918 2070
rect 2154 1834 2238 2070
rect 2474 1834 8218 2070
rect 8454 1834 8538 2070
rect 8774 1834 13626 2070
rect 13862 1834 13946 2070
rect 14182 1834 14266 2070
rect 14502 1834 14586 2070
rect 14822 1834 14906 2070
rect 15142 1834 16100 2070
rect 0 1750 16100 1834
rect 0 1514 958 1750
rect 1194 1514 1278 1750
rect 1514 1514 1598 1750
rect 1834 1514 1918 1750
rect 2154 1514 2238 1750
rect 2474 1514 8218 1750
rect 8454 1514 8538 1750
rect 8774 1514 13626 1750
rect 13862 1514 13946 1750
rect 14182 1514 14266 1750
rect 14502 1514 14586 1750
rect 14822 1514 14906 1750
rect 15142 1514 16100 1750
rect 0 1430 16100 1514
rect 0 1194 958 1430
rect 1194 1194 1278 1430
rect 1514 1194 1598 1430
rect 1834 1194 1918 1430
rect 2154 1194 2238 1430
rect 2474 1194 8218 1430
rect 8454 1194 8538 1430
rect 8774 1194 13626 1430
rect 13862 1194 13946 1430
rect 14182 1194 14266 1430
rect 14502 1194 14586 1430
rect 14822 1194 14906 1430
rect 15142 1194 16100 1430
rect 0 1110 16100 1194
rect 0 874 958 1110
rect 1194 874 1278 1110
rect 1514 874 1598 1110
rect 1834 874 1918 1110
rect 2154 874 2238 1110
rect 2474 874 8218 1110
rect 8454 874 8538 1110
rect 8774 874 13626 1110
rect 13862 874 13946 1110
rect 14182 874 14266 1110
rect 14502 874 14586 1110
rect 14822 874 14906 1110
rect 15142 874 16100 1110
rect 0 816 16100 874
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 ~/PDKS/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623995306
transform 1 0 5796 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_1
timestamp 1623995306
transform 1 0 5796 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILL_67 ~/PDKS/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623995306
transform 1 0 5796 0 -1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILL_71
timestamp 1623995306
transform 1 0 5888 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_32
timestamp 1623995306
transform 1 0 5796 0 -1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_36
timestamp 1623995306
transform 1 0 5888 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILL_33 ~/PDKS/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623995306
transform 1 0 6164 0 -1 6800
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_21
timestamp 1623995306
transform 1 0 6164 0 -1 6800
box -38 -48 222 592
use sky130_fd_sc_hd__clkinv_1  U70 ~/PDKS/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623995306
transform -1 0 6164 0 -1 6800
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  U72
timestamp 1623995306
transform -1 0 6256 0 1 5712
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_1
timestamp 1623995306
transform -1 0 6164 0 -1 6800
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_2
timestamp 1623995306
transform -1 0 6256 0 1 5712
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_13 ~/PDKS/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623995306
transform -1 0 6716 0 -1 6800
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  U96
timestamp 1623995306
transform -1 0 6716 0 -1 6800
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_35
timestamp 1623995306
transform 1 0 6256 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_31
timestamp 1623995306
transform 1 0 6348 0 -1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILL_70
timestamp 1623995306
transform 1 0 6256 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILL_66
timestamp 1623995306
transform 1 0 6348 0 -1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_6
timestamp 1623995306
transform -1 0 6624 0 1 5712
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  U80
timestamp 1623995306
transform -1 0 6624 0 1 5712
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_7 ~/PDKS/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623995306
transform 1 0 6624 0 1 5712
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  U11
timestamp 1623995306
transform 1 0 6624 0 1 5712
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_4
timestamp 1623995306
transform 1 0 7084 0 -1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1623995306
transform 1 0 7084 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_5
timestamp 1623995306
transform 1 0 7084 0 -1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_2
timestamp 1623995306
transform 1 0 7084 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILL_10 ~/PDKS/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623995306
transform 1 0 6716 0 -1 6800
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILL_11
timestamp 1623995306
transform 1 0 7176 0 1 5712
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_5
timestamp 1623995306
transform 1 0 6716 0 -1 6800
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_6
timestamp 1623995306
transform 1 0 7176 0 1 5712
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  dac_select_bits_reg_5_ ~/PDKS/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623995306
transform 1 0 7176 0 -1 6800
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_11
timestamp 1623995306
transform 1 0 7176 0 -1 6800
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILL_69
timestamp 1623995306
transform 1 0 8280 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_34
timestamp 1623995306
transform 1 0 8280 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__and2_0  U13
timestamp 1623995306
transform 1 0 7820 0 1 5712
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_10
timestamp 1623995306
transform 1 0 7820 0 1 5712
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  U97
timestamp 1623995306
transform -1 0 7820 0 1 5712
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_14
timestamp 1623995306
transform -1 0 7820 0 1 5712
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_22
timestamp 1623995306
transform 1 0 8464 0 1 5712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILL_34
timestamp 1623995306
transform 1 0 8464 0 1 5712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1623995306
transform 1 0 8372 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_3
timestamp 1623995306
transform 1 0 8372 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_15
timestamp 1623995306
transform 1 0 9108 0 1 5712
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  U98
timestamp 1623995306
transform 1 0 9108 0 1 5712
box -38 -48 314 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_3 ~/PDKS/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623995306
transform 1 0 8648 0 -1 6800
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILL_4
timestamp 1623995306
transform 1 0 8648 0 -1 6800
box -38 -48 774 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_12
timestamp 1623995306
transform -1 0 9108 0 1 5712
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  U15
timestamp 1623995306
transform -1 0 9108 0 1 5712
box -38 -48 498 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_20
timestamp 1623995306
transform 1 0 9384 0 -1 6800
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILL_32
timestamp 1623995306
transform 1 0 9384 0 -1 6800
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_30
timestamp 1623995306
transform 1 0 9568 0 -1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILL_65
timestamp 1623995306
transform 1 0 9568 0 -1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_5
timestamp 1623995306
transform 1 0 9660 0 -1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_3
timestamp 1623995306
transform 1 0 9660 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_6
timestamp 1623995306
transform 1 0 9660 0 -1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_4
timestamp 1623995306
transform 1 0 9660 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__nor2b_1  sky130_fd_sc_hd__nor2b_1_2 ~/PDKS/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623995306
transform -1 0 10212 0 1 5712
box -38 -48 498 592
use sky130_fd_sc_hd__nor2b_1  U106
timestamp 1623995306
transform -1 0 10212 0 1 5712
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_1
timestamp 1623995306
transform 1 0 9384 0 1 5712
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  U69
timestamp 1623995306
transform 1 0 9384 0 1 5712
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_6
timestamp 1623995306
transform 1 0 9752 0 -1 6800
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  U10
timestamp 1623995306
transform 1 0 9752 0 -1 6800
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILL_64
timestamp 1623995306
transform 1 0 10212 0 -1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILL_68
timestamp 1623995306
transform 1 0 10212 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_29
timestamp 1623995306
transform 1 0 10212 0 -1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_33
timestamp 1623995306
transform 1 0 10212 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_6
timestamp 1623995306
transform 1 0 5796 0 1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_7
timestamp 1623995306
transform 1 0 5796 0 1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__and2_0  U9
timestamp 1623995306
transform 1 0 6440 0 1 6800
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_5
timestamp 1623995306
transform 1 0 6440 0 1 6800
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  U94
timestamp 1623995306
transform -1 0 6164 0 1 6800
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  U95
timestamp 1623995306
transform -1 0 6440 0 1 6800
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_11
timestamp 1623995306
transform -1 0 6164 0 1 6800
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_12
timestamp 1623995306
transform -1 0 6440 0 1 6800
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  dac_select_bits_reg_4_
timestamp 1623995306
transform 1 0 6900 0 1 6800
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_13
timestamp 1623995306
transform 1 0 6900 0 1 6800
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_12
timestamp 1623995306
transform -1 0 9936 0 1 6800
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  dac_mask_reg_4_
timestamp 1623995306
transform -1 0 9936 0 1 6800
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_7
timestamp 1623995306
transform 1 0 8372 0 1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_8
timestamp 1623995306
transform 1 0 8372 0 1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_28
timestamp 1623995306
transform 1 0 10120 0 1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILL_63
timestamp 1623995306
transform 1 0 10120 0 1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_19
timestamp 1623995306
transform 1 0 9936 0 1 6800
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILL_31
timestamp 1623995306
transform 1 0 9936 0 1 6800
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_8
timestamp 1623995306
transform 1 0 10212 0 1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_9
timestamp 1623995306
transform 1 0 10212 0 1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_3
timestamp 1623995306
transform -1 0 6440 0 -1 7888
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  U73
timestamp 1623995306
transform -1 0 6440 0 -1 7888
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_27
timestamp 1623995306
transform 1 0 5796 0 -1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILL_62
timestamp 1623995306
transform 1 0 5796 0 -1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_3
timestamp 1623995306
transform 1 0 5888 0 -1 7888
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  U74
timestamp 1623995306
transform 1 0 5888 0 -1 7888
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_18
timestamp 1623995306
transform 1 0 6440 0 -1 7888
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILL_30
timestamp 1623995306
transform 1 0 6440 0 -1 7888
box -38 -48 222 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_4
timestamp 1623995306
transform 1 0 6624 0 -1 7888
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  U7
timestamp 1623995306
transform 1 0 6624 0 -1 7888
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_9
timestamp 1623995306
transform 1 0 7084 0 -1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_10
timestamp 1623995306
transform 1 0 7084 0 -1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  dac_select_bits_reg_3_
timestamp 1623995306
transform 1 0 7176 0 -1 7888
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_15
timestamp 1623995306
transform 1 0 7176 0 -1 7888
box -38 -48 1510 592
use sky130_fd_sc_hd__nor2b_1  sky130_fd_sc_hd__nor2b_1_1
timestamp 1623995306
transform 1 0 9200 0 -1 7888
box -38 -48 498 592
use sky130_fd_sc_hd__nor2b_1  U105
timestamp 1623995306
transform 1 0 9200 0 -1 7888
box -38 -48 498 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_4
timestamp 1623995306
transform 1 0 8648 0 -1 7888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILL_9
timestamp 1623995306
transform 1 0 8648 0 -1 7888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_17
timestamp 1623995306
transform 1 0 9016 0 -1 7888
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILL_29
timestamp 1623995306
transform 1 0 9016 0 -1 7888
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_2
timestamp 1623995306
transform 1 0 9752 0 -1 7888
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  U71
timestamp 1623995306
transform 1 0 9752 0 -1 7888
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_26
timestamp 1623995306
transform 1 0 10212 0 -1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILL_61
timestamp 1623995306
transform 1 0 10212 0 -1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_16
timestamp 1623995306
transform 1 0 10028 0 -1 7888
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILL_28
timestamp 1623995306
transform 1 0 10028 0 -1 7888
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_10
timestamp 1623995306
transform 1 0 9660 0 -1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_11
timestamp 1623995306
transform 1 0 9660 0 -1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__nor2b_1  sky130_fd_sc_hd__nor2b_1_3
timestamp 1623995306
transform -1 0 7820 0 1 7888
box -38 -48 498 592
use sky130_fd_sc_hd__nor2b_1  U107
timestamp 1623995306
transform -1 0 7820 0 1 7888
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_14
timestamp 1623995306
transform -1 0 7360 0 1 7888
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  dac_mask_reg_3_
timestamp 1623995306
transform -1 0 7360 0 1 7888
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_11
timestamp 1623995306
transform 1 0 5796 0 1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_12
timestamp 1623995306
transform 1 0 5796 0 1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_12
timestamp 1623995306
transform 1 0 8372 0 1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_13
timestamp 1623995306
transform 1 0 8372 0 1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILL_27
timestamp 1623995306
transform 1 0 8096 0 1 7888
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_15
timestamp 1623995306
transform 1 0 8096 0 1 7888
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILL_60
timestamp 1623995306
transform 1 0 8280 0 1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_25
timestamp 1623995306
transform 1 0 8280 0 1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  U81
timestamp 1623995306
transform 1 0 7820 0 1 7888
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_7
timestamp 1623995306
transform 1 0 7820 0 1 7888
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  dac_select_bits_reg_6_
timestamp 1623995306
transform 1 0 8464 0 1 7888
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_9
timestamp 1623995306
transform 1 0 8464 0 1 7888
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  sky130_fd_sc_hd__conb_1_0 ~/PDKS/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623995306
transform -1 0 10212 0 1 7888
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  clk_gate_dac_select_bits_reg_LTIE
timestamp 1623995306
transform -1 0 10212 0 1 7888
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_13
timestamp 1623995306
transform 1 0 10212 0 1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_14
timestamp 1623995306
transform 1 0 10212 0 1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_1  U82
timestamp 1623995306
transform -1 0 6164 0 -1 8976
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_7
timestamp 1623995306
transform -1 0 6164 0 -1 8976
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILL_59
timestamp 1623995306
transform 1 0 5796 0 -1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_24
timestamp 1623995306
transform 1 0 5796 0 -1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_4  CTS_ccl_a_inv_00003 ~/PDKS/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623995306
transform -1 0 6808 0 -1 8976
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_0
timestamp 1623995306
transform -1 0 6808 0 -1 8976
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_14
timestamp 1623995306
transform 1 0 7084 0 -1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_15
timestamp 1623995306
transform 1 0 7084 0 -1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILL_26
timestamp 1623995306
transform 1 0 6808 0 -1 8976
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_14
timestamp 1623995306
transform 1 0 6808 0 -1 8976
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILL_58
timestamp 1623995306
transform 1 0 6992 0 -1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_23
timestamp 1623995306
transform 1 0 6992 0 -1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__and2_0  U8
timestamp 1623995306
transform -1 0 7636 0 -1 8976
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_13
timestamp 1623995306
transform -1 0 7636 0 -1 8976
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_8
timestamp 1623995306
transform 1 0 7636 0 -1 8976
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  dac_mask_reg_6_
timestamp 1623995306
transform 1 0 7636 0 -1 8976
box -38 -48 1510 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_9
timestamp 1623995306
transform -1 0 9660 0 -1 8976
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  U12
timestamp 1623995306
transform -1 0 9660 0 -1 8976
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_22
timestamp 1623995306
transform 1 0 9108 0 -1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILL_57
timestamp 1623995306
transform 1 0 9108 0 -1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_11
timestamp 1623995306
transform 1 0 9752 0 -1 8976
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  U14
timestamp 1623995306
transform 1 0 9752 0 -1 8976
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_21
timestamp 1623995306
transform 1 0 10212 0 -1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILL_56
timestamp 1623995306
transform 1 0 10212 0 -1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_15
timestamp 1623995306
transform 1 0 9660 0 -1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_16
timestamp 1623995306
transform 1 0 9660 0 -1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_16
timestamp 1623995306
transform 1 0 5796 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_17
timestamp 1623995306
transform 1 0 5796 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_18
timestamp 1623995306
transform 1 0 6532 0 -1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILL_53
timestamp 1623995306
transform 1 0 6532 0 -1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  sky130_fd_sc_hd__clkinv_2_0 ~/PDKS/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623995306
transform -1 0 6532 0 -1 10064
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  CTS_ccl_a_inv_00006
timestamp 1623995306
transform -1 0 6532 0 -1 10064
box -38 -48 406 592
use sky130_fd_sc_hd__nor2b_1  sky130_fd_sc_hd__nor2b_1_4
timestamp 1623995306
transform 1 0 5888 0 1 8976
box -38 -48 498 592
use sky130_fd_sc_hd__nor2b_1  U108
timestamp 1623995306
transform 1 0 5888 0 1 8976
box -38 -48 498 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_3
timestamp 1623995306
transform 1 0 5796 0 -1 10064
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILL_8
timestamp 1623995306
transform 1 0 5796 0 -1 10064
box -38 -48 406 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_3
timestamp 1623995306
transform 1 0 6624 0 -1 10064
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  U6
timestamp 1623995306
transform 1 0 6624 0 -1 10064
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_19
timestamp 1623995306
transform 1 0 7084 0 -1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_20
timestamp 1623995306
transform 1 0 7084 0 -1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  dac_select_bits_reg_0_
timestamp 1623995306
transform 1 0 7176 0 -1 10064
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  dac_mask_reg_2_
timestamp 1623995306
transform -1 0 7820 0 1 8976
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_6
timestamp 1623995306
transform 1 0 7176 0 -1 10064
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_16
timestamp 1623995306
transform -1 0 7820 0 1 8976
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_17
timestamp 1623995306
transform 1 0 8372 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_18
timestamp 1623995306
transform 1 0 8372 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILL_55
timestamp 1623995306
transform 1 0 8280 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_20
timestamp 1623995306
transform 1 0 8280 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__and2_0  U17
timestamp 1623995306
transform 1 0 7820 0 1 8976
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_15
timestamp 1623995306
transform 1 0 7820 0 1 8976
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_19
timestamp 1623995306
transform 1 0 8464 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILL_54
timestamp 1623995306
transform 1 0 8464 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_12
timestamp 1623995306
transform 1 0 8648 0 -1 10064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILL_24
timestamp 1623995306
transform 1 0 8648 0 -1 10064
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_0
timestamp 1623995306
transform -1 0 9200 0 -1 10064
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  U67
timestamp 1623995306
transform -1 0 9200 0 -1 10064
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_17
timestamp 1623995306
transform 1 0 8832 0 -1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILL_52
timestamp 1623995306
transform 1 0 8832 0 -1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_11
timestamp 1623995306
transform 1 0 9200 0 -1 10064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILL_23
timestamp 1623995306
transform 1 0 9200 0 -1 10064
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  dac_mask_reg_5_
timestamp 1623995306
transform 1 0 8556 0 1 8976
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_10
timestamp 1623995306
transform 1 0 8556 0 1 8976
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_20
timestamp 1623995306
transform 1 0 9660 0 -1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_21
timestamp 1623995306
transform 1 0 9660 0 -1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  U79
timestamp 1623995306
transform 1 0 9384 0 -1 10064
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_6
timestamp 1623995306
transform 1 0 9384 0 -1 10064
box -38 -48 314 592
use sky130_fd_sc_hd__nor2b_1  U104
timestamp 1623995306
transform -1 0 10212 0 -1 10064
box -38 -48 498 592
use sky130_fd_sc_hd__nor2b_1  sky130_fd_sc_hd__nor2b_1_0
timestamp 1623995306
transform -1 0 10212 0 -1 10064
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_18
timestamp 1623995306
transform 1 0 10212 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_19
timestamp 1623995306
transform 1 0 10212 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILL_25
timestamp 1623995306
transform 1 0 10028 0 1 8976
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_13
timestamp 1623995306
transform 1 0 10028 0 1 8976
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILL_51
timestamp 1623995306
transform 1 0 10212 0 -1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_16
timestamp 1623995306
transform 1 0 10212 0 -1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_8
timestamp 1623995306
transform -1 0 6256 0 1 10064
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  U91
timestamp 1623995306
transform -1 0 6256 0 1 10064
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_15
timestamp 1623995306
transform 1 0 5888 0 1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILL_50
timestamp 1623995306
transform 1 0 5888 0 1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_21
timestamp 1623995306
transform 1 0 5796 0 1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_22
timestamp 1623995306
transform 1 0 5796 0 1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_10
timestamp 1623995306
transform 1 0 6256 0 1 10064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILL_22
timestamp 1623995306
transform 1 0 6256 0 1 10064
box -38 -48 222 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_14
timestamp 1623995306
transform 1 0 6440 0 1 10064
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  U16
timestamp 1623995306
transform 1 0 6440 0 1 10064
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  dac_select_bits_reg_7_
timestamp 1623995306
transform 1 0 6900 0 1 10064
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_7
timestamp 1623995306
transform 1 0 6900 0 1 10064
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_5
timestamp 1623995306
transform 1 0 8464 0 1 10064
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  dac_mask_reg_7_
timestamp 1623995306
transform 1 0 8464 0 1 10064
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_22
timestamp 1623995306
transform 1 0 8372 0 1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_23
timestamp 1623995306
transform 1 0 8372 0 1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_11
timestamp 1623995306
transform 1 0 9936 0 1 10064
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  U100
timestamp 1623995306
transform 1 0 9936 0 1 10064
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_23
timestamp 1623995306
transform 1 0 10212 0 1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_24
timestamp 1623995306
transform 1 0 10212 0 1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILL_49
timestamp 1623995306
transform 1 0 5796 0 -1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_14
timestamp 1623995306
transform 1 0 5796 0 -1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__and2_0  U5
timestamp 1623995306
transform 1 0 6440 0 -1 11152
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_8
timestamp 1623995306
transform 1 0 6440 0 -1 11152
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  U75
timestamp 1623995306
transform 1 0 6164 0 -1 11152
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  U93
timestamp 1623995306
transform -1 0 6164 0 -1 11152
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_4
timestamp 1623995306
transform 1 0 6164 0 -1 11152
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_10
timestamp 1623995306
transform -1 0 6164 0 -1 11152
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_24
timestamp 1623995306
transform 1 0 7084 0 -1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_25
timestamp 1623995306
transform 1 0 7084 0 -1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILL_21
timestamp 1623995306
transform 1 0 6900 0 -1 11152
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_9
timestamp 1623995306
transform 1 0 6900 0 -1 11152
box -38 -48 222 592
use sky130_fd_sc_hd__sdlclkp_4  clk_gate_dac_select_bits_reg_latch ~/PDKS/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624005307
transform -1 0 8832 0 -1 11152
box -38 -48 1694 592
use sky130_fd_sc_hd__sdlclkp_4  sky130_fd_sc_hd__sdlclkp_4_0
timestamp 1624005307
transform -1 0 8832 0 -1 11152
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_2
timestamp 1623995306
transform 1 0 8832 0 -1 11152
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILL_3
timestamp 1623995306
transform 1 0 8832 0 -1 11152
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_25
timestamp 1623995306
transform 1 0 9660 0 -1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_26
timestamp 1623995306
transform 1 0 9660 0 -1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILL_48
timestamp 1623995306
transform 1 0 9568 0 -1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_13
timestamp 1623995306
transform 1 0 9568 0 -1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILL_47
timestamp 1623995306
transform 1 0 9752 0 -1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_12
timestamp 1623995306
transform 1 0 9752 0 -1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  U102 ~/PDKS/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623995306
transform 1 0 9844 0 -1 11152
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  sky130_fd_sc_hd__o21ai_1_0
timestamp 1623995306
transform 1 0 9844 0 -1 11152
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILL_46
timestamp 1623995306
transform 1 0 10212 0 -1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_11
timestamp 1623995306
transform 1 0 10212 0 -1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__nor2b_1  sky130_fd_sc_hd__nor2b_1_5
timestamp 1623995306
transform -1 0 6440 0 1 11152
box -38 -48 498 592
use sky130_fd_sc_hd__nor2b_1  U109
timestamp 1623995306
transform -1 0 6440 0 1 11152
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_17
timestamp 1623995306
transform -1 0 7912 0 1 11152
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  dac_select_bits_reg_2_
timestamp 1623995306
transform -1 0 7912 0 1 11152
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_10
timestamp 1623995306
transform 1 0 5888 0 1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILL_45
timestamp 1623995306
transform 1 0 5888 0 1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_26
timestamp 1623995306
transform 1 0 5796 0 1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_27
timestamp 1623995306
transform 1 0 5796 0 1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_0
timestamp 1623995306
transform 1 0 8464 0 1 11152
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  dac_mask_reg_0_
timestamp 1623995306
transform 1 0 8464 0 1 11152
box -38 -48 1510 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_18
timestamp 1623995306
transform 1 0 7912 0 1 11152
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  U22
timestamp 1623995306
transform 1 0 7912 0 1 11152
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_27
timestamp 1623995306
transform 1 0 8372 0 1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_28
timestamp 1623995306
transform 1 0 8372 0 1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_8
timestamp 1623995306
transform -1 0 10212 0 1 11152
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  U83
timestamp 1623995306
transform -1 0 10212 0 1 11152
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_28
timestamp 1623995306
transform 1 0 10212 0 1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_29
timestamp 1623995306
transform 1 0 10212 0 1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILL_44
timestamp 1623995306
transform 1 0 5796 0 -1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_9
timestamp 1623995306
transform 1 0 5796 0 -1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__and2_0  U4
timestamp 1623995306
transform 1 0 5888 0 -1 12240
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  U3
timestamp 1623995306
transform 1 0 6348 0 -1 12240
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_1
timestamp 1623995306
transform 1 0 5888 0 -1 12240
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_2
timestamp 1623995306
transform 1 0 6348 0 -1 12240
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_29
timestamp 1623995306
transform 1 0 7084 0 -1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_30
timestamp 1623995306
transform 1 0 7084 0 -1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  U77
timestamp 1623995306
transform 1 0 7176 0 -1 12240
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  U92
timestamp 1623995306
transform 1 0 6808 0 -1 12240
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_5
timestamp 1623995306
transform 1 0 7176 0 -1 12240
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_9
timestamp 1623995306
transform 1 0 6808 0 -1 12240
box -38 -48 314 592
use sky130_fd_sc_hd__fill_8  FILL_2
timestamp 1623995306
transform 1 0 7452 0 -1 12240
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_1
timestamp 1623995306
transform 1 0 7452 0 -1 12240
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_19
timestamp 1623995306
transform 1 0 8188 0 -1 12240
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  dac_select_bits_reg_1_
timestamp 1623995306
transform 1 0 8188 0 -1 12240
box -38 -48 1510 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_0
timestamp 1623995306
transform -1 0 10212 0 -1 12240
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  U21
timestamp 1623995306
transform -1 0 10212 0 -1 12240
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_8
timestamp 1623995306
transform 1 0 10212 0 -1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILL_43
timestamp 1623995306
transform 1 0 10212 0 -1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_30
timestamp 1623995306
transform 1 0 9660 0 -1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_31
timestamp 1623995306
transform 1 0 9660 0 -1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__nor2b_1  sky130_fd_sc_hd__nor2b_1_6
timestamp 1623995306
transform 1 0 7452 0 1 12240
box -38 -48 498 592
use sky130_fd_sc_hd__nor2b_1  U110
timestamp 1623995306
transform 1 0 7452 0 1 12240
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_18
timestamp 1623995306
transform 1 0 5980 0 1 12240
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  dac_mask_reg_1_
timestamp 1623995306
transform 1 0 5980 0 1 12240
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_7
timestamp 1623995306
transform 1 0 5888 0 1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILL_42
timestamp 1623995306
transform 1 0 5888 0 1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_31
timestamp 1623995306
transform 1 0 5796 0 1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_32
timestamp 1623995306
transform 1 0 5796 0 1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_32
timestamp 1623995306
transform 1 0 8372 0 1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_33
timestamp 1623995306
transform 1 0 8372 0 1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILL_20
timestamp 1623995306
transform 1 0 8188 0 1 12240
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_8
timestamp 1623995306
transform 1 0 8188 0 1 12240
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_1  U103
timestamp 1623995306
transform 1 0 7912 0 1 12240
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_17
timestamp 1623995306
transform 1 0 7912 0 1 12240
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILL_19
timestamp 1623995306
transform 1 0 8464 0 1 12240
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_7
timestamp 1623995306
transform 1 0 8464 0 1 12240
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILL_41
timestamp 1623995306
transform 1 0 8648 0 1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_6
timestamp 1623995306
transform 1 0 8648 0 1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  state_r_reg_0_
timestamp 1623995306
transform 1 0 8740 0 1 12240
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_1
timestamp 1623995306
transform 1 0 8740 0 1 12240
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_33
timestamp 1623995306
transform 1 0 10212 0 1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_34
timestamp 1623995306
transform 1 0 10212 0 1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_5
timestamp 1623995306
transform 1 0 5980 0 -1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILL_40
timestamp 1623995306
transform 1 0 5980 0 -1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_4
timestamp 1623995306
transform 1 0 6072 0 -1 13328
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  U76
timestamp 1623995306
transform 1 0 6072 0 -1 13328
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_6
timestamp 1623995306
transform 1 0 5796 0 -1 13328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILL_18
timestamp 1623995306
transform 1 0 5796 0 -1 13328
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_36
timestamp 1623995306
transform 1 0 5796 0 1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_37
timestamp 1623995306
transform 1 0 5796 0 1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_5
timestamp 1623995306
transform -1 0 6900 0 1 13328
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  U78
timestamp 1623995306
transform -1 0 6900 0 1 13328
box -38 -48 314 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_0
timestamp 1623995306
transform 1 0 5888 0 1 13328
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILL_1
timestamp 1623995306
transform 1 0 5888 0 1 13328
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_2
timestamp 1623995306
transform 1 0 6348 0 -1 13328
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILL_7
timestamp 1623995306
transform 1 0 6348 0 -1 13328
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_2 ~/PDKS/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623995306
transform 1 0 6716 0 -1 13328
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  U90
timestamp 1623995306
transform 1 0 6716 0 -1 13328
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_34
timestamp 1623995306
transform 1 0 7084 0 -1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_35
timestamp 1623995306
transform 1 0 7084 0 -1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILL_39
timestamp 1623995306
transform 1 0 6992 0 -1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_4
timestamp 1623995306
transform 1 0 6992 0 -1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  state_r_reg_1_
timestamp 1623995306
transform -1 0 8372 0 1 13328
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  run_adc_n_reg
timestamp 1623995306
transform -1 0 8648 0 -1 13328
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_2
timestamp 1623995306
transform -1 0 8372 0 1 13328
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_4
timestamp 1623995306
transform -1 0 8648 0 -1 13328
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_37
timestamp 1623995306
transform 1 0 8372 0 1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_38
timestamp 1623995306
transform 1 0 8372 0 1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_1  U84
timestamp 1623995306
transform 1 0 8464 0 1 13328
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_9
timestamp 1623995306
transform 1 0 8464 0 1 13328
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILL_38
timestamp 1623995306
transform 1 0 8648 0 -1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_3
timestamp 1623995306
transform 1 0 8648 0 -1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__and2_0  U19
timestamp 1623995306
transform -1 0 9660 0 -1 13328
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_17
timestamp 1623995306
transform -1 0 9660 0 -1 13328
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  U18 ~/PDKS/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623995306
transform -1 0 9200 0 -1 13328
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  sky130_fd_sc_hd__nand2b_1_0
timestamp 1623995306
transform -1 0 9200 0 -1 13328
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  out_valid_reg
timestamp 1623995306
transform 1 0 8740 0 1 13328
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_3
timestamp 1623995306
transform 1 0 8740 0 1 13328
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_35
timestamp 1623995306
transform 1 0 9660 0 -1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_36
timestamp 1623995306
transform 1 0 9660 0 -1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  U99
timestamp 1623995306
transform 1 0 9752 0 -1 13328
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_16
timestamp 1623995306
transform 1 0 9752 0 -1 13328
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_38
timestamp 1623995306
transform 1 0 10212 0 1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_39
timestamp 1623995306
transform 1 0 10212 0 1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILL_17
timestamp 1623995306
transform 1 0 10028 0 -1 13328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_5
timestamp 1623995306
transform 1 0 10028 0 -1 13328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILL_37
timestamp 1623995306
transform 1 0 10212 0 -1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_2
timestamp 1623995306
transform 1 0 10212 0 -1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_39
timestamp 1623995306
transform 1 0 5796 0 -1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_40
timestamp 1623995306
transform 1 0 5796 0 -1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_1  U68
timestamp 1623995306
transform -1 0 6256 0 -1 14416
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_0
timestamp 1623995306
transform -1 0 6256 0 -1 14416
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILL_36
timestamp 1623995306
transform 1 0 5888 0 -1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_1
timestamp 1623995306
transform 1 0 5888 0 -1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_1
timestamp 1623995306
transform -1 0 6716 0 -1 14416
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  U88
timestamp 1623995306
transform -1 0 6716 0 -1 14416
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILL_16
timestamp 1623995306
transform 1 0 6256 0 -1 14416
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_4
timestamp 1623995306
transform 1 0 6256 0 -1 14416
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_40
timestamp 1623995306
transform 1 0 7084 0 -1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_41
timestamp 1623995306
transform 1 0 7084 0 -1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILL_6
timestamp 1623995306
transform 1 0 6716 0 -1 14416
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_1
timestamp 1623995306
transform 1 0 6716 0 -1 14416
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILL_5
timestamp 1623995306
transform 1 0 7176 0 -1 14416
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_0
timestamp 1623995306
transform 1 0 7176 0 -1 14416
box -38 -48 406 592
use sky130_fd_sc_hd__and2_0  U20
timestamp 1623995306
transform 1 0 7544 0 -1 14416
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_16
timestamp 1623995306
transform 1 0 7544 0 -1 14416
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  U89 ~/PDKS/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623995306
transform -1 0 8372 0 -1 14416
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  sky130_fd_sc_hd__nand3_1_0
timestamp 1623995306
transform -1 0 8372 0 -1 14416
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_41
timestamp 1623995306
transform 1 0 8372 0 -1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_42
timestamp 1623995306
transform 1 0 8372 0 -1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILL_15
timestamp 1623995306
transform 1 0 8464 0 -1 14416
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_3
timestamp 1623995306
transform 1 0 8464 0 -1 14416
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_0
timestamp 1623995306
transform -1 0 8924 0 -1 14416
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  U85
timestamp 1623995306
transform -1 0 8924 0 -1 14416
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILL_14
timestamp 1623995306
transform 1 0 8924 0 -1 14416
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_2
timestamp 1623995306
transform 1 0 8924 0 -1 14416
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILL_35
timestamp 1623995306
transform 1 0 9108 0 -1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_0
timestamp 1623995306
transform 1 0 9108 0 -1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_1  U86
timestamp 1623995306
transform 1 0 9200 0 -1 14416
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_10
timestamp 1623995306
transform 1 0 9200 0 -1 14416
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_1
timestamp 1623995306
transform 1 0 9476 0 -1 14416
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_0
timestamp 1623995306
transform 1 0 9752 0 -1 14416
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILL_13
timestamp 1623995306
transform 1 0 9476 0 -1 14416
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILL_12
timestamp 1623995306
transform 1 0 9752 0 -1 14416
box -38 -48 222 592
use sky130_fd_sc_hd__a21oi_1  sky130_fd_sc_hd__a21oi_1_0 ~/PDKS/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623995306
transform 1 0 9936 0 -1 14416
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  U101
timestamp 1623995306
transform 1 0 9936 0 -1 14416
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_42
timestamp 1623995306
transform 1 0 9660 0 -1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  WELLTAP_43
timestamp 1623995306
transform 1 0 9660 0 -1 14416
box -38 -48 130 592
<< labels >>
rlabel metal2 s 216 20031 244 20128 6 clk
port 0 nsew signal input
rlabel metal2 s 8036 20031 8064 20128 6 rst_n
port 1 nsew signal input
rlabel metal2 s 15856 20031 15884 20128 6 adc_start
port 2 nsew signal input
rlabel metal2 s 0 20080 97 20108 6 comparator_val
port 3 nsew signal input
rlabel metal2 s 0 20 97 48 6 run_adc_n
port 4 nsew signal tristate
rlabel metal2 s 0 2196 97 2224 6 adc_val[7]
port 5 nsew signal tristate
rlabel metal2 s 0 4440 97 4468 6 adc_val[6]
port 6 nsew signal tristate
rlabel metal2 s 0 6684 97 6712 6 adc_val[5]
port 7 nsew signal tristate
rlabel metal2 s 0 8928 97 8956 6 adc_val[4]
port 8 nsew signal tristate
rlabel metal2 s 0 11104 97 11132 6 adc_val[3]
port 9 nsew signal tristate
rlabel metal2 s 0 13348 97 13376 6 adc_val[2]
port 10 nsew signal tristate
rlabel metal2 s 0 15592 97 15620 6 adc_val[1]
port 11 nsew signal tristate
rlabel metal2 s 0 17836 97 17864 6 adc_val[0]
port 12 nsew signal tristate
rlabel metal2 s 16003 20080 16100 20108 6 out_valid
port 13 nsew signal tristate
rlabel metal5 s 14468 17680 16100 19312 6 VSS
port 14 nsew ground bidirectional
rlabel metal5 s 0 17680 1632 19312 6 VSS
port 15 nsew ground bidirectional
rlabel metal5 s 14468 816 16100 2448 6 VSS
port 16 nsew ground bidirectional
rlabel metal5 s 0 816 1632 2448 6 VSS
port 17 nsew ground bidirectional
rlabel metal4 s 13568 18496 15200 20128 6 VSS
port 18 nsew ground bidirectional
rlabel metal4 s 13568 0 15200 1632 6 VSS
port 19 nsew ground bidirectional
rlabel metal4 s 900 18496 2532 20128 6 VSS
port 20 nsew ground bidirectional
rlabel metal4 s 900 0 2532 1632 6 VSS
port 21 nsew ground bidirectional
rlabel metal5 s 14468 15232 16100 16864 6 VDD
port 22 nsew power bidirectional
rlabel metal5 s 0 15232 1632 16864 6 VDD
port 23 nsew power bidirectional
rlabel metal5 s 14468 3264 16100 4896 6 VDD
port 24 nsew power bidirectional
rlabel metal5 s 0 3264 1632 4896 6 VDD
port 25 nsew power bidirectional
rlabel metal4 s 11120 18496 12752 20128 6 VDD
port 26 nsew power bidirectional
rlabel metal4 s 11120 0 12752 1632 6 VDD
port 27 nsew power bidirectional
rlabel metal4 s 3348 18496 4980 20128 6 VDD
port 28 nsew power bidirectional
rlabel metal4 s 3348 0 4980 1632 6 VDD
port 29 nsew power bidirectional
rlabel metal2 s 216 20031 244 20128 1 clk
port 0 nsew signal input
rlabel metal2 s 8036 20031 8064 20128 1 rst_n
port 1 nsew signal input
rlabel metal2 s 15856 20031 15884 20128 1 adc_start
port 2 nsew signal input
rlabel metal2 s 0 20080 97 20108 1 comparator_val
port 3 nsew signal input
rlabel metal2 s 0 20 97 48 1 run_adc_n
port 4 nsew signal tristate
rlabel metal2 s 0 2196 97 2224 1 adc_val[7]
port 5 nsew signal tristate
rlabel metal2 s 0 4440 97 4468 1 adc_val[6]
port 6 nsew signal tristate
rlabel metal2 s 0 6684 97 6712 1 adc_val[5]
port 7 nsew signal tristate
rlabel metal2 s 0 8928 97 8956 1 adc_val[4]
port 8 nsew signal tristate
rlabel metal2 s 0 11104 97 11132 1 adc_val[3]
port 9 nsew signal tristate
rlabel metal2 s 0 13348 97 13376 1 adc_val[2]
port 10 nsew signal tristate
rlabel metal2 s 0 15592 97 15620 1 adc_val[1]
port 11 nsew signal tristate
rlabel metal2 s 0 17836 97 17864 1 adc_val[0]
port 12 nsew signal tristate
rlabel metal2 s 16003 20080 16100 20108 1 out_valid
port 13 nsew signal tristate
rlabel metal5 s 14468 17680 16100 19312 1 VSS
port 14 nsew ground bidirectional
rlabel metal5 s 0 17680 1632 19312 1 VSS
port 15 nsew ground bidirectional
rlabel metal5 s 14468 816 16100 2448 1 VSS
port 16 nsew ground bidirectional
rlabel metal5 s 0 816 1632 2448 1 VSS
port 17 nsew ground bidirectional
rlabel metal4 s 13568 18496 15200 20128 1 VSS
port 18 nsew ground bidirectional
rlabel metal4 s 13568 0 15200 1632 1 VSS
port 19 nsew ground bidirectional
rlabel metal4 s 900 18496 2532 20128 1 VSS
port 20 nsew ground bidirectional
rlabel metal4 s 900 0 2532 1632 1 VSS
port 21 nsew ground bidirectional
rlabel metal5 s 14468 15232 16100 16864 1 VDD
port 22 nsew power bidirectional
rlabel metal5 s 0 15232 1632 16864 1 VDD
port 23 nsew power bidirectional
rlabel metal5 s 14468 3264 16100 4896 1 VDD
port 24 nsew power bidirectional
rlabel metal5 s 0 3264 1632 4896 1 VDD
port 25 nsew power bidirectional
rlabel metal4 s 11120 18496 12752 20128 1 VDD
port 26 nsew power bidirectional
rlabel metal4 s 11120 0 12752 1632 1 VDD
port 27 nsew power bidirectional
rlabel metal4 s 3348 18496 4980 20128 1 VDD
port 28 nsew power bidirectional
rlabel metal4 s 3348 0 4980 1632 1 VDD
port 29 nsew power bidirectional
<< end >>
