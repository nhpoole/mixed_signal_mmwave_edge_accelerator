magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect -4660 -4860 4660 4460
<< nwell >>
rect -3358 582 3358 3158
<< pwell >>
rect -3348 256 3348 408
rect -3348 56 -52 256
rect -3348 -976 -2996 56
rect -204 -976 -52 56
rect -3348 -1192 -52 -976
rect 3196 -1192 3348 256
rect -3348 -1344 3348 -1192
rect -3348 -2616 -2996 -1344
rect 2996 -2616 3348 -1344
rect -3348 -2768 3348 -2616
rect -3348 -3396 -3196 -2768
rect 3196 -3396 3348 -2768
rect -3348 -3548 3348 -3396
<< psubdiff >>
rect -3322 349 3322 382
rect -3322 315 -3145 349
rect -3111 315 -3077 349
rect -3043 315 -3009 349
rect -2975 315 -2941 349
rect -2907 315 -2873 349
rect -2839 315 -2805 349
rect -2771 315 -2737 349
rect -2703 315 -2669 349
rect -2635 315 -2601 349
rect -2567 315 -2533 349
rect -2499 315 -2465 349
rect -2431 315 -2397 349
rect -2363 315 -2329 349
rect -2295 315 -2261 349
rect -2227 315 -2193 349
rect -2159 315 -2125 349
rect -2091 315 -2057 349
rect -2023 315 -1989 349
rect -1955 315 -1921 349
rect -1887 315 -1853 349
rect -1819 315 -1785 349
rect -1751 315 -1717 349
rect -1683 315 -1649 349
rect -1615 315 -1581 349
rect -1547 315 -1513 349
rect -1479 315 -1445 349
rect -1411 315 -1377 349
rect -1343 315 -1309 349
rect -1275 315 -1241 349
rect -1207 315 -1173 349
rect -1139 315 -1105 349
rect -1071 315 -1037 349
rect -1003 315 -969 349
rect -935 315 -901 349
rect -867 315 -833 349
rect -799 315 -765 349
rect -731 315 -697 349
rect -663 315 -629 349
rect -595 315 -561 349
rect -527 315 -493 349
rect -459 315 -425 349
rect -391 315 -357 349
rect -323 315 -289 349
rect -255 315 -221 349
rect -187 315 -153 349
rect -119 315 -85 349
rect -51 315 -17 349
rect 17 315 51 349
rect 85 315 119 349
rect 153 315 187 349
rect 221 315 255 349
rect 289 315 323 349
rect 357 315 391 349
rect 425 315 459 349
rect 493 315 527 349
rect 561 315 595 349
rect 629 315 663 349
rect 697 315 731 349
rect 765 315 799 349
rect 833 315 867 349
rect 901 315 935 349
rect 969 315 1003 349
rect 1037 315 1071 349
rect 1105 315 1139 349
rect 1173 315 1207 349
rect 1241 315 1275 349
rect 1309 315 1343 349
rect 1377 315 1411 349
rect 1445 315 1479 349
rect 1513 315 1547 349
rect 1581 315 1615 349
rect 1649 315 1683 349
rect 1717 315 1751 349
rect 1785 315 1819 349
rect 1853 315 1887 349
rect 1921 315 1955 349
rect 1989 315 2023 349
rect 2057 315 2091 349
rect 2125 315 2159 349
rect 2193 315 2227 349
rect 2261 315 2295 349
rect 2329 315 2363 349
rect 2397 315 2431 349
rect 2465 315 2499 349
rect 2533 315 2567 349
rect 2601 315 2635 349
rect 2669 315 2703 349
rect 2737 315 2771 349
rect 2805 315 2839 349
rect 2873 315 2907 349
rect 2941 315 2975 349
rect 3009 315 3043 349
rect 3077 315 3111 349
rect 3145 315 3322 349
rect -3322 282 3322 315
rect -3322 215 -3222 282
rect -3322 181 -3289 215
rect -3255 181 -3222 215
rect 3222 215 3322 282
rect -3322 147 -3222 181
rect -3322 113 -3289 147
rect -3255 113 -3222 147
rect -3322 79 -3222 113
rect -3322 45 -3289 79
rect -3255 45 -3222 79
rect -3322 11 -3222 45
rect -3322 -23 -3289 11
rect -3255 -23 -3222 11
rect -3322 -57 -3222 -23
rect -3322 -91 -3289 -57
rect -3255 -91 -3222 -57
rect -3322 -125 -3222 -91
rect -3322 -159 -3289 -125
rect -3255 -159 -3222 -125
rect -3322 -193 -3222 -159
rect -3322 -227 -3289 -193
rect -3255 -227 -3222 -193
rect -3322 -261 -3222 -227
rect -3322 -295 -3289 -261
rect -3255 -295 -3222 -261
rect -3322 -329 -3222 -295
rect -3322 -363 -3289 -329
rect -3255 -363 -3222 -329
rect -3322 -397 -3222 -363
rect -3322 -431 -3289 -397
rect -3255 -431 -3222 -397
rect -3322 -465 -3222 -431
rect -3322 -499 -3289 -465
rect -3255 -499 -3222 -465
rect -3322 -533 -3222 -499
rect -3322 -567 -3289 -533
rect -3255 -567 -3222 -533
rect -3322 -601 -3222 -567
rect -3322 -635 -3289 -601
rect -3255 -635 -3222 -601
rect -3322 -669 -3222 -635
rect -3322 -703 -3289 -669
rect -3255 -703 -3222 -669
rect -3322 -737 -3222 -703
rect -3322 -771 -3289 -737
rect -3255 -771 -3222 -737
rect -3322 -805 -3222 -771
rect -3322 -839 -3289 -805
rect -3255 -839 -3222 -805
rect -3322 -873 -3222 -839
rect -3322 -907 -3289 -873
rect -3255 -907 -3222 -873
rect -3322 -941 -3222 -907
rect -3322 -975 -3289 -941
rect -3255 -975 -3222 -941
rect -3322 -1009 -3222 -975
rect -3322 -1043 -3289 -1009
rect -3255 -1043 -3222 -1009
rect -3322 -1077 -3222 -1043
rect -3322 -1111 -3289 -1077
rect -3255 -1111 -3222 -1077
rect -3122 149 -78 182
rect -3122 115 -2943 149
rect -2909 115 -2875 149
rect -2841 115 -2807 149
rect -2773 115 -2739 149
rect -2705 115 -2671 149
rect -2637 115 -2603 149
rect -2569 115 -2535 149
rect -2501 115 -2467 149
rect -2433 115 -2399 149
rect -2365 115 -2331 149
rect -2297 115 -2263 149
rect -2229 115 -2195 149
rect -2161 115 -2127 149
rect -2093 115 -2059 149
rect -2025 115 -1991 149
rect -1957 115 -1923 149
rect -1889 115 -1855 149
rect -1821 115 -1787 149
rect -1753 115 -1719 149
rect -1685 115 -1651 149
rect -1617 115 -1583 149
rect -1549 115 -1515 149
rect -1481 115 -1447 149
rect -1413 115 -1379 149
rect -1345 115 -1311 149
rect -1277 115 -1243 149
rect -1209 115 -1175 149
rect -1141 115 -1107 149
rect -1073 115 -1039 149
rect -1005 115 -971 149
rect -937 115 -903 149
rect -869 115 -835 149
rect -801 115 -767 149
rect -733 115 -699 149
rect -665 115 -631 149
rect -597 115 -563 149
rect -529 115 -495 149
rect -461 115 -427 149
rect -393 115 -359 149
rect -325 115 -291 149
rect -257 115 -78 149
rect -3122 82 -78 115
rect -3122 -1 -3022 82
rect -3122 -35 -3089 -1
rect -3055 -35 -3022 -1
rect -3122 -69 -3022 -35
rect -3122 -103 -3089 -69
rect -3055 -103 -3022 -69
rect -3122 -137 -3022 -103
rect -3122 -171 -3089 -137
rect -3055 -171 -3022 -137
rect -3122 -205 -3022 -171
rect -3122 -239 -3089 -205
rect -3055 -239 -3022 -205
rect -3122 -273 -3022 -239
rect -3122 -307 -3089 -273
rect -3055 -307 -3022 -273
rect -3122 -341 -3022 -307
rect -3122 -375 -3089 -341
rect -3055 -375 -3022 -341
rect -3122 -409 -3022 -375
rect -3122 -443 -3089 -409
rect -3055 -443 -3022 -409
rect -3122 -477 -3022 -443
rect -3122 -511 -3089 -477
rect -3055 -511 -3022 -477
rect -3122 -545 -3022 -511
rect -3122 -579 -3089 -545
rect -3055 -579 -3022 -545
rect -3122 -613 -3022 -579
rect -3122 -647 -3089 -613
rect -3055 -647 -3022 -613
rect -3122 -681 -3022 -647
rect -3122 -715 -3089 -681
rect -3055 -715 -3022 -681
rect -3122 -749 -3022 -715
rect -3122 -783 -3089 -749
rect -3055 -783 -3022 -749
rect -3122 -817 -3022 -783
rect -3122 -851 -3089 -817
rect -3055 -851 -3022 -817
rect -3122 -885 -3022 -851
rect -3122 -919 -3089 -885
rect -3055 -919 -3022 -885
rect -3122 -1002 -3022 -919
rect -178 -1 -78 82
rect -178 -35 -145 -1
rect -111 -35 -78 -1
rect -178 -69 -78 -35
rect -178 -103 -145 -69
rect -111 -103 -78 -69
rect -178 -137 -78 -103
rect -178 -171 -145 -137
rect -111 -171 -78 -137
rect -178 -205 -78 -171
rect -178 -239 -145 -205
rect -111 -239 -78 -205
rect -178 -273 -78 -239
rect -178 -307 -145 -273
rect -111 -307 -78 -273
rect -178 -341 -78 -307
rect -178 -375 -145 -341
rect -111 -375 -78 -341
rect -178 -409 -78 -375
rect -178 -443 -145 -409
rect -111 -443 -78 -409
rect -178 -477 -78 -443
rect -178 -511 -145 -477
rect -111 -511 -78 -477
rect -178 -545 -78 -511
rect -178 -579 -145 -545
rect -111 -579 -78 -545
rect -178 -613 -78 -579
rect -178 -647 -145 -613
rect -111 -647 -78 -613
rect -178 -681 -78 -647
rect -178 -715 -145 -681
rect -111 -715 -78 -681
rect -178 -749 -78 -715
rect -178 -783 -145 -749
rect -111 -783 -78 -749
rect -178 -817 -78 -783
rect -178 -851 -145 -817
rect -111 -851 -78 -817
rect -178 -885 -78 -851
rect -178 -919 -145 -885
rect -111 -919 -78 -885
rect -178 -1002 -78 -919
rect -3122 -1035 -78 -1002
rect -3122 -1069 -2943 -1035
rect -2909 -1069 -2875 -1035
rect -2841 -1069 -2807 -1035
rect -2773 -1069 -2739 -1035
rect -2705 -1069 -2671 -1035
rect -2637 -1069 -2603 -1035
rect -2569 -1069 -2535 -1035
rect -2501 -1069 -2467 -1035
rect -2433 -1069 -2399 -1035
rect -2365 -1069 -2331 -1035
rect -2297 -1069 -2263 -1035
rect -2229 -1069 -2195 -1035
rect -2161 -1069 -2127 -1035
rect -2093 -1069 -2059 -1035
rect -2025 -1069 -1991 -1035
rect -1957 -1069 -1923 -1035
rect -1889 -1069 -1855 -1035
rect -1821 -1069 -1787 -1035
rect -1753 -1069 -1719 -1035
rect -1685 -1069 -1651 -1035
rect -1617 -1069 -1583 -1035
rect -1549 -1069 -1515 -1035
rect -1481 -1069 -1447 -1035
rect -1413 -1069 -1379 -1035
rect -1345 -1069 -1311 -1035
rect -1277 -1069 -1243 -1035
rect -1209 -1069 -1175 -1035
rect -1141 -1069 -1107 -1035
rect -1073 -1069 -1039 -1035
rect -1005 -1069 -971 -1035
rect -937 -1069 -903 -1035
rect -869 -1069 -835 -1035
rect -801 -1069 -767 -1035
rect -733 -1069 -699 -1035
rect -665 -1069 -631 -1035
rect -597 -1069 -563 -1035
rect -529 -1069 -495 -1035
rect -461 -1069 -427 -1035
rect -393 -1069 -359 -1035
rect -325 -1069 -291 -1035
rect -257 -1069 -78 -1035
rect -3122 -1102 -78 -1069
rect 3222 181 3255 215
rect 3289 181 3322 215
rect 3222 147 3322 181
rect 3222 113 3255 147
rect 3289 113 3322 147
rect 3222 79 3322 113
rect 3222 45 3255 79
rect 3289 45 3322 79
rect 3222 11 3322 45
rect 3222 -23 3255 11
rect 3289 -23 3322 11
rect 3222 -57 3322 -23
rect 3222 -91 3255 -57
rect 3289 -91 3322 -57
rect 3222 -125 3322 -91
rect 3222 -159 3255 -125
rect 3289 -159 3322 -125
rect 3222 -193 3322 -159
rect 3222 -227 3255 -193
rect 3289 -227 3322 -193
rect 3222 -261 3322 -227
rect 3222 -295 3255 -261
rect 3289 -295 3322 -261
rect 3222 -329 3322 -295
rect 3222 -363 3255 -329
rect 3289 -363 3322 -329
rect 3222 -397 3322 -363
rect 3222 -431 3255 -397
rect 3289 -431 3322 -397
rect 3222 -465 3322 -431
rect 3222 -499 3255 -465
rect 3289 -499 3322 -465
rect 3222 -533 3322 -499
rect 3222 -567 3255 -533
rect 3289 -567 3322 -533
rect 3222 -601 3322 -567
rect 3222 -635 3255 -601
rect 3289 -635 3322 -601
rect 3222 -669 3322 -635
rect 3222 -703 3255 -669
rect 3289 -703 3322 -669
rect 3222 -737 3322 -703
rect 3222 -771 3255 -737
rect 3289 -771 3322 -737
rect 3222 -805 3322 -771
rect 3222 -839 3255 -805
rect 3289 -839 3322 -805
rect 3222 -873 3322 -839
rect 3222 -907 3255 -873
rect 3289 -907 3322 -873
rect 3222 -941 3322 -907
rect 3222 -975 3255 -941
rect 3289 -975 3322 -941
rect 3222 -1009 3322 -975
rect 3222 -1043 3255 -1009
rect 3289 -1043 3322 -1009
rect 3222 -1077 3322 -1043
rect -3322 -1145 -3222 -1111
rect -3322 -1179 -3289 -1145
rect -3255 -1179 -3222 -1145
rect -3322 -1213 -3222 -1179
rect -3322 -1247 -3289 -1213
rect -3255 -1247 -3222 -1213
rect 3222 -1111 3255 -1077
rect 3289 -1111 3322 -1077
rect 3222 -1145 3322 -1111
rect 3222 -1179 3255 -1145
rect 3289 -1179 3322 -1145
rect 3222 -1213 3322 -1179
rect -3322 -1281 -3222 -1247
rect -3322 -1315 -3289 -1281
rect -3255 -1315 -3222 -1281
rect -3322 -1349 -3222 -1315
rect -3322 -1383 -3289 -1349
rect -3255 -1383 -3222 -1349
rect -3322 -1417 -3222 -1383
rect -3322 -1451 -3289 -1417
rect -3255 -1451 -3222 -1417
rect -3322 -1485 -3222 -1451
rect -3322 -1519 -3289 -1485
rect -3255 -1519 -3222 -1485
rect -3322 -1553 -3222 -1519
rect -3322 -1587 -3289 -1553
rect -3255 -1587 -3222 -1553
rect -3322 -1621 -3222 -1587
rect -3322 -1655 -3289 -1621
rect -3255 -1655 -3222 -1621
rect -3322 -1689 -3222 -1655
rect -3322 -1723 -3289 -1689
rect -3255 -1723 -3222 -1689
rect -3322 -1757 -3222 -1723
rect -3322 -1791 -3289 -1757
rect -3255 -1791 -3222 -1757
rect -3322 -1825 -3222 -1791
rect -3322 -1859 -3289 -1825
rect -3255 -1859 -3222 -1825
rect -3322 -1893 -3222 -1859
rect -3322 -1927 -3289 -1893
rect -3255 -1927 -3222 -1893
rect -3322 -1961 -3222 -1927
rect -3322 -1995 -3289 -1961
rect -3255 -1995 -3222 -1961
rect -3322 -2029 -3222 -1995
rect -3322 -2063 -3289 -2029
rect -3255 -2063 -3222 -2029
rect -3322 -2097 -3222 -2063
rect -3322 -2131 -3289 -2097
rect -3255 -2131 -3222 -2097
rect -3322 -2165 -3222 -2131
rect -3322 -2199 -3289 -2165
rect -3255 -2199 -3222 -2165
rect -3322 -2233 -3222 -2199
rect -3322 -2267 -3289 -2233
rect -3255 -2267 -3222 -2233
rect -3322 -2301 -3222 -2267
rect -3322 -2335 -3289 -2301
rect -3255 -2335 -3222 -2301
rect -3322 -2369 -3222 -2335
rect -3322 -2403 -3289 -2369
rect -3255 -2403 -3222 -2369
rect -3322 -2437 -3222 -2403
rect -3322 -2471 -3289 -2437
rect -3255 -2471 -3222 -2437
rect -3322 -2505 -3222 -2471
rect -3322 -2539 -3289 -2505
rect -3255 -2539 -3222 -2505
rect -3322 -2573 -3222 -2539
rect -3322 -2607 -3289 -2573
rect -3255 -2607 -3222 -2573
rect -3322 -2641 -3222 -2607
rect -3322 -2675 -3289 -2641
rect -3255 -2675 -3222 -2641
rect -3322 -2709 -3222 -2675
rect -3322 -2743 -3289 -2709
rect -3255 -2743 -3222 -2709
rect -3122 -1251 3122 -1218
rect -3122 -1285 -2941 -1251
rect -2907 -1285 -2873 -1251
rect -2839 -1285 -2805 -1251
rect -2771 -1285 -2737 -1251
rect -2703 -1285 -2669 -1251
rect -2635 -1285 -2601 -1251
rect -2567 -1285 -2533 -1251
rect -2499 -1285 -2465 -1251
rect -2431 -1285 -2397 -1251
rect -2363 -1285 -2329 -1251
rect -2295 -1285 -2261 -1251
rect -2227 -1285 -2193 -1251
rect -2159 -1285 -2125 -1251
rect -2091 -1285 -2057 -1251
rect -2023 -1285 -1989 -1251
rect -1955 -1285 -1921 -1251
rect -1887 -1285 -1853 -1251
rect -1819 -1285 -1785 -1251
rect -1751 -1285 -1717 -1251
rect -1683 -1285 -1649 -1251
rect -1615 -1285 -1581 -1251
rect -1547 -1285 -1513 -1251
rect -1479 -1285 -1445 -1251
rect -1411 -1285 -1377 -1251
rect -1343 -1285 -1309 -1251
rect -1275 -1285 -1241 -1251
rect -1207 -1285 -1173 -1251
rect -1139 -1285 -1105 -1251
rect -1071 -1285 -1037 -1251
rect -1003 -1285 -969 -1251
rect -935 -1285 -901 -1251
rect -867 -1285 -833 -1251
rect -799 -1285 -765 -1251
rect -731 -1285 -697 -1251
rect -663 -1285 -629 -1251
rect -595 -1285 -561 -1251
rect -527 -1285 -493 -1251
rect -459 -1285 -425 -1251
rect -391 -1285 -357 -1251
rect -323 -1285 -289 -1251
rect -255 -1285 -221 -1251
rect -187 -1285 -153 -1251
rect -119 -1285 -85 -1251
rect -51 -1285 -17 -1251
rect 17 -1285 51 -1251
rect 85 -1285 119 -1251
rect 153 -1285 187 -1251
rect 221 -1285 255 -1251
rect 289 -1285 323 -1251
rect 357 -1285 391 -1251
rect 425 -1285 459 -1251
rect 493 -1285 527 -1251
rect 561 -1285 595 -1251
rect 629 -1285 663 -1251
rect 697 -1285 731 -1251
rect 765 -1285 799 -1251
rect 833 -1285 867 -1251
rect 901 -1285 935 -1251
rect 969 -1285 1003 -1251
rect 1037 -1285 1071 -1251
rect 1105 -1285 1139 -1251
rect 1173 -1285 1207 -1251
rect 1241 -1285 1275 -1251
rect 1309 -1285 1343 -1251
rect 1377 -1285 1411 -1251
rect 1445 -1285 1479 -1251
rect 1513 -1285 1547 -1251
rect 1581 -1285 1615 -1251
rect 1649 -1285 1683 -1251
rect 1717 -1285 1751 -1251
rect 1785 -1285 1819 -1251
rect 1853 -1285 1887 -1251
rect 1921 -1285 1955 -1251
rect 1989 -1285 2023 -1251
rect 2057 -1285 2091 -1251
rect 2125 -1285 2159 -1251
rect 2193 -1285 2227 -1251
rect 2261 -1285 2295 -1251
rect 2329 -1285 2363 -1251
rect 2397 -1285 2431 -1251
rect 2465 -1285 2499 -1251
rect 2533 -1285 2567 -1251
rect 2601 -1285 2635 -1251
rect 2669 -1285 2703 -1251
rect 2737 -1285 2771 -1251
rect 2805 -1285 2839 -1251
rect 2873 -1285 2907 -1251
rect 2941 -1285 3122 -1251
rect -3122 -1318 3122 -1285
rect -3122 -1385 -3022 -1318
rect -3122 -1419 -3089 -1385
rect -3055 -1419 -3022 -1385
rect -3122 -1453 -3022 -1419
rect -3122 -1487 -3089 -1453
rect -3055 -1487 -3022 -1453
rect -3122 -1521 -3022 -1487
rect -3122 -1555 -3089 -1521
rect -3055 -1555 -3022 -1521
rect -3122 -1589 -3022 -1555
rect -3122 -1623 -3089 -1589
rect -3055 -1623 -3022 -1589
rect -3122 -1657 -3022 -1623
rect -3122 -1691 -3089 -1657
rect -3055 -1691 -3022 -1657
rect -3122 -1725 -3022 -1691
rect -3122 -1759 -3089 -1725
rect -3055 -1759 -3022 -1725
rect -3122 -1793 -3022 -1759
rect -3122 -1827 -3089 -1793
rect -3055 -1827 -3022 -1793
rect -3122 -1861 -3022 -1827
rect -3122 -1895 -3089 -1861
rect -3055 -1895 -3022 -1861
rect -3122 -1929 -3022 -1895
rect -3122 -1963 -3089 -1929
rect -3055 -1963 -3022 -1929
rect -3122 -1997 -3022 -1963
rect -3122 -2031 -3089 -1997
rect -3055 -2031 -3022 -1997
rect -3122 -2065 -3022 -2031
rect -3122 -2099 -3089 -2065
rect -3055 -2099 -3022 -2065
rect -3122 -2133 -3022 -2099
rect -3122 -2167 -3089 -2133
rect -3055 -2167 -3022 -2133
rect -3122 -2201 -3022 -2167
rect -3122 -2235 -3089 -2201
rect -3055 -2235 -3022 -2201
rect -3122 -2269 -3022 -2235
rect -3122 -2303 -3089 -2269
rect -3055 -2303 -3022 -2269
rect -3122 -2337 -3022 -2303
rect -3122 -2371 -3089 -2337
rect -3055 -2371 -3022 -2337
rect -3122 -2405 -3022 -2371
rect -3122 -2439 -3089 -2405
rect -3055 -2439 -3022 -2405
rect -3122 -2473 -3022 -2439
rect -3122 -2507 -3089 -2473
rect -3055 -2507 -3022 -2473
rect -3122 -2541 -3022 -2507
rect -3122 -2575 -3089 -2541
rect -3055 -2575 -3022 -2541
rect -3122 -2642 -3022 -2575
rect 3022 -1385 3122 -1318
rect 3022 -1419 3055 -1385
rect 3089 -1419 3122 -1385
rect 3022 -1453 3122 -1419
rect 3022 -1487 3055 -1453
rect 3089 -1487 3122 -1453
rect 3022 -1521 3122 -1487
rect 3022 -1555 3055 -1521
rect 3089 -1555 3122 -1521
rect 3022 -1589 3122 -1555
rect 3022 -1623 3055 -1589
rect 3089 -1623 3122 -1589
rect 3022 -1657 3122 -1623
rect 3022 -1691 3055 -1657
rect 3089 -1691 3122 -1657
rect 3022 -1725 3122 -1691
rect 3022 -1759 3055 -1725
rect 3089 -1759 3122 -1725
rect 3022 -1793 3122 -1759
rect 3022 -1827 3055 -1793
rect 3089 -1827 3122 -1793
rect 3022 -1861 3122 -1827
rect 3022 -1895 3055 -1861
rect 3089 -1895 3122 -1861
rect 3022 -1929 3122 -1895
rect 3022 -1963 3055 -1929
rect 3089 -1963 3122 -1929
rect 3022 -1997 3122 -1963
rect 3022 -2031 3055 -1997
rect 3089 -2031 3122 -1997
rect 3022 -2065 3122 -2031
rect 3022 -2099 3055 -2065
rect 3089 -2099 3122 -2065
rect 3022 -2133 3122 -2099
rect 3022 -2167 3055 -2133
rect 3089 -2167 3122 -2133
rect 3022 -2201 3122 -2167
rect 3022 -2235 3055 -2201
rect 3089 -2235 3122 -2201
rect 3022 -2269 3122 -2235
rect 3022 -2303 3055 -2269
rect 3089 -2303 3122 -2269
rect 3022 -2337 3122 -2303
rect 3022 -2371 3055 -2337
rect 3089 -2371 3122 -2337
rect 3022 -2405 3122 -2371
rect 3022 -2439 3055 -2405
rect 3089 -2439 3122 -2405
rect 3022 -2473 3122 -2439
rect 3022 -2507 3055 -2473
rect 3089 -2507 3122 -2473
rect 3022 -2541 3122 -2507
rect 3022 -2575 3055 -2541
rect 3089 -2575 3122 -2541
rect 3022 -2642 3122 -2575
rect -3122 -2675 3122 -2642
rect -3122 -2709 -2941 -2675
rect -2907 -2709 -2873 -2675
rect -2839 -2709 -2805 -2675
rect -2771 -2709 -2737 -2675
rect -2703 -2709 -2669 -2675
rect -2635 -2709 -2601 -2675
rect -2567 -2709 -2533 -2675
rect -2499 -2709 -2465 -2675
rect -2431 -2709 -2397 -2675
rect -2363 -2709 -2329 -2675
rect -2295 -2709 -2261 -2675
rect -2227 -2709 -2193 -2675
rect -2159 -2709 -2125 -2675
rect -2091 -2709 -2057 -2675
rect -2023 -2709 -1989 -2675
rect -1955 -2709 -1921 -2675
rect -1887 -2709 -1853 -2675
rect -1819 -2709 -1785 -2675
rect -1751 -2709 -1717 -2675
rect -1683 -2709 -1649 -2675
rect -1615 -2709 -1581 -2675
rect -1547 -2709 -1513 -2675
rect -1479 -2709 -1445 -2675
rect -1411 -2709 -1377 -2675
rect -1343 -2709 -1309 -2675
rect -1275 -2709 -1241 -2675
rect -1207 -2709 -1173 -2675
rect -1139 -2709 -1105 -2675
rect -1071 -2709 -1037 -2675
rect -1003 -2709 -969 -2675
rect -935 -2709 -901 -2675
rect -867 -2709 -833 -2675
rect -799 -2709 -765 -2675
rect -731 -2709 -697 -2675
rect -663 -2709 -629 -2675
rect -595 -2709 -561 -2675
rect -527 -2709 -493 -2675
rect -459 -2709 -425 -2675
rect -391 -2709 -357 -2675
rect -323 -2709 -289 -2675
rect -255 -2709 -221 -2675
rect -187 -2709 -153 -2675
rect -119 -2709 -85 -2675
rect -51 -2709 -17 -2675
rect 17 -2709 51 -2675
rect 85 -2709 119 -2675
rect 153 -2709 187 -2675
rect 221 -2709 255 -2675
rect 289 -2709 323 -2675
rect 357 -2709 391 -2675
rect 425 -2709 459 -2675
rect 493 -2709 527 -2675
rect 561 -2709 595 -2675
rect 629 -2709 663 -2675
rect 697 -2709 731 -2675
rect 765 -2709 799 -2675
rect 833 -2709 867 -2675
rect 901 -2709 935 -2675
rect 969 -2709 1003 -2675
rect 1037 -2709 1071 -2675
rect 1105 -2709 1139 -2675
rect 1173 -2709 1207 -2675
rect 1241 -2709 1275 -2675
rect 1309 -2709 1343 -2675
rect 1377 -2709 1411 -2675
rect 1445 -2709 1479 -2675
rect 1513 -2709 1547 -2675
rect 1581 -2709 1615 -2675
rect 1649 -2709 1683 -2675
rect 1717 -2709 1751 -2675
rect 1785 -2709 1819 -2675
rect 1853 -2709 1887 -2675
rect 1921 -2709 1955 -2675
rect 1989 -2709 2023 -2675
rect 2057 -2709 2091 -2675
rect 2125 -2709 2159 -2675
rect 2193 -2709 2227 -2675
rect 2261 -2709 2295 -2675
rect 2329 -2709 2363 -2675
rect 2397 -2709 2431 -2675
rect 2465 -2709 2499 -2675
rect 2533 -2709 2567 -2675
rect 2601 -2709 2635 -2675
rect 2669 -2709 2703 -2675
rect 2737 -2709 2771 -2675
rect 2805 -2709 2839 -2675
rect 2873 -2709 2907 -2675
rect 2941 -2709 3122 -2675
rect -3122 -2742 3122 -2709
rect 3222 -1247 3255 -1213
rect 3289 -1247 3322 -1213
rect 3222 -1281 3322 -1247
rect 3222 -1315 3255 -1281
rect 3289 -1315 3322 -1281
rect 3222 -1349 3322 -1315
rect 3222 -1383 3255 -1349
rect 3289 -1383 3322 -1349
rect 3222 -1417 3322 -1383
rect 3222 -1451 3255 -1417
rect 3289 -1451 3322 -1417
rect 3222 -1485 3322 -1451
rect 3222 -1519 3255 -1485
rect 3289 -1519 3322 -1485
rect 3222 -1553 3322 -1519
rect 3222 -1587 3255 -1553
rect 3289 -1587 3322 -1553
rect 3222 -1621 3322 -1587
rect 3222 -1655 3255 -1621
rect 3289 -1655 3322 -1621
rect 3222 -1689 3322 -1655
rect 3222 -1723 3255 -1689
rect 3289 -1723 3322 -1689
rect 3222 -1757 3322 -1723
rect 3222 -1791 3255 -1757
rect 3289 -1791 3322 -1757
rect 3222 -1825 3322 -1791
rect 3222 -1859 3255 -1825
rect 3289 -1859 3322 -1825
rect 3222 -1893 3322 -1859
rect 3222 -1927 3255 -1893
rect 3289 -1927 3322 -1893
rect 3222 -1961 3322 -1927
rect 3222 -1995 3255 -1961
rect 3289 -1995 3322 -1961
rect 3222 -2029 3322 -1995
rect 3222 -2063 3255 -2029
rect 3289 -2063 3322 -2029
rect 3222 -2097 3322 -2063
rect 3222 -2131 3255 -2097
rect 3289 -2131 3322 -2097
rect 3222 -2165 3322 -2131
rect 3222 -2199 3255 -2165
rect 3289 -2199 3322 -2165
rect 3222 -2233 3322 -2199
rect 3222 -2267 3255 -2233
rect 3289 -2267 3322 -2233
rect 3222 -2301 3322 -2267
rect 3222 -2335 3255 -2301
rect 3289 -2335 3322 -2301
rect 3222 -2369 3322 -2335
rect 3222 -2403 3255 -2369
rect 3289 -2403 3322 -2369
rect 3222 -2437 3322 -2403
rect 3222 -2471 3255 -2437
rect 3289 -2471 3322 -2437
rect 3222 -2505 3322 -2471
rect 3222 -2539 3255 -2505
rect 3289 -2539 3322 -2505
rect 3222 -2573 3322 -2539
rect 3222 -2607 3255 -2573
rect 3289 -2607 3322 -2573
rect 3222 -2641 3322 -2607
rect 3222 -2675 3255 -2641
rect 3289 -2675 3322 -2641
rect 3222 -2709 3322 -2675
rect -3322 -2777 -3222 -2743
rect -3322 -2811 -3289 -2777
rect -3255 -2811 -3222 -2777
rect -3322 -2845 -3222 -2811
rect -3322 -2879 -3289 -2845
rect -3255 -2879 -3222 -2845
rect -3322 -2913 -3222 -2879
rect -3322 -2947 -3289 -2913
rect -3255 -2947 -3222 -2913
rect -3322 -2981 -3222 -2947
rect -3322 -3015 -3289 -2981
rect -3255 -3015 -3222 -2981
rect -3322 -3049 -3222 -3015
rect -3322 -3083 -3289 -3049
rect -3255 -3083 -3222 -3049
rect -3322 -3117 -3222 -3083
rect -3322 -3151 -3289 -3117
rect -3255 -3151 -3222 -3117
rect -3322 -3185 -3222 -3151
rect -3322 -3219 -3289 -3185
rect -3255 -3219 -3222 -3185
rect -3322 -3253 -3222 -3219
rect -3322 -3287 -3289 -3253
rect -3255 -3287 -3222 -3253
rect -3322 -3321 -3222 -3287
rect -3322 -3355 -3289 -3321
rect -3255 -3355 -3222 -3321
rect -3322 -3422 -3222 -3355
rect 3222 -2743 3255 -2709
rect 3289 -2743 3322 -2709
rect 3222 -2777 3322 -2743
rect 3222 -2811 3255 -2777
rect 3289 -2811 3322 -2777
rect 3222 -2845 3322 -2811
rect 3222 -2879 3255 -2845
rect 3289 -2879 3322 -2845
rect 3222 -2913 3322 -2879
rect 3222 -2947 3255 -2913
rect 3289 -2947 3322 -2913
rect 3222 -2981 3322 -2947
rect 3222 -3015 3255 -2981
rect 3289 -3015 3322 -2981
rect 3222 -3049 3322 -3015
rect 3222 -3083 3255 -3049
rect 3289 -3083 3322 -3049
rect 3222 -3117 3322 -3083
rect 3222 -3151 3255 -3117
rect 3289 -3151 3322 -3117
rect 3222 -3185 3322 -3151
rect 3222 -3219 3255 -3185
rect 3289 -3219 3322 -3185
rect 3222 -3253 3322 -3219
rect 3222 -3287 3255 -3253
rect 3289 -3287 3322 -3253
rect 3222 -3321 3322 -3287
rect 3222 -3355 3255 -3321
rect 3289 -3355 3322 -3321
rect 3222 -3422 3322 -3355
rect -3322 -3455 3322 -3422
rect -3322 -3489 -3145 -3455
rect -3111 -3489 -3077 -3455
rect -3043 -3489 -3009 -3455
rect -2975 -3489 -2941 -3455
rect -2907 -3489 -2873 -3455
rect -2839 -3489 -2805 -3455
rect -2771 -3489 -2737 -3455
rect -2703 -3489 -2669 -3455
rect -2635 -3489 -2601 -3455
rect -2567 -3489 -2533 -3455
rect -2499 -3489 -2465 -3455
rect -2431 -3489 -2397 -3455
rect -2363 -3489 -2329 -3455
rect -2295 -3489 -2261 -3455
rect -2227 -3489 -2193 -3455
rect -2159 -3489 -2125 -3455
rect -2091 -3489 -2057 -3455
rect -2023 -3489 -1989 -3455
rect -1955 -3489 -1921 -3455
rect -1887 -3489 -1853 -3455
rect -1819 -3489 -1785 -3455
rect -1751 -3489 -1717 -3455
rect -1683 -3489 -1649 -3455
rect -1615 -3489 -1581 -3455
rect -1547 -3489 -1513 -3455
rect -1479 -3489 -1445 -3455
rect -1411 -3489 -1377 -3455
rect -1343 -3489 -1309 -3455
rect -1275 -3489 -1241 -3455
rect -1207 -3489 -1173 -3455
rect -1139 -3489 -1105 -3455
rect -1071 -3489 -1037 -3455
rect -1003 -3489 -969 -3455
rect -935 -3489 -901 -3455
rect -867 -3489 -833 -3455
rect -799 -3489 -765 -3455
rect -731 -3489 -697 -3455
rect -663 -3489 -629 -3455
rect -595 -3489 -561 -3455
rect -527 -3489 -493 -3455
rect -459 -3489 -425 -3455
rect -391 -3489 -357 -3455
rect -323 -3489 -289 -3455
rect -255 -3489 -221 -3455
rect -187 -3489 -153 -3455
rect -119 -3489 -85 -3455
rect -51 -3489 -17 -3455
rect 17 -3489 51 -3455
rect 85 -3489 119 -3455
rect 153 -3489 187 -3455
rect 221 -3489 255 -3455
rect 289 -3489 323 -3455
rect 357 -3489 391 -3455
rect 425 -3489 459 -3455
rect 493 -3489 527 -3455
rect 561 -3489 595 -3455
rect 629 -3489 663 -3455
rect 697 -3489 731 -3455
rect 765 -3489 799 -3455
rect 833 -3489 867 -3455
rect 901 -3489 935 -3455
rect 969 -3489 1003 -3455
rect 1037 -3489 1071 -3455
rect 1105 -3489 1139 -3455
rect 1173 -3489 1207 -3455
rect 1241 -3489 1275 -3455
rect 1309 -3489 1343 -3455
rect 1377 -3489 1411 -3455
rect 1445 -3489 1479 -3455
rect 1513 -3489 1547 -3455
rect 1581 -3489 1615 -3455
rect 1649 -3489 1683 -3455
rect 1717 -3489 1751 -3455
rect 1785 -3489 1819 -3455
rect 1853 -3489 1887 -3455
rect 1921 -3489 1955 -3455
rect 1989 -3489 2023 -3455
rect 2057 -3489 2091 -3455
rect 2125 -3489 2159 -3455
rect 2193 -3489 2227 -3455
rect 2261 -3489 2295 -3455
rect 2329 -3489 2363 -3455
rect 2397 -3489 2431 -3455
rect 2465 -3489 2499 -3455
rect 2533 -3489 2567 -3455
rect 2601 -3489 2635 -3455
rect 2669 -3489 2703 -3455
rect 2737 -3489 2771 -3455
rect 2805 -3489 2839 -3455
rect 2873 -3489 2907 -3455
rect 2941 -3489 2975 -3455
rect 3009 -3489 3043 -3455
rect 3077 -3489 3111 -3455
rect 3145 -3489 3322 -3455
rect -3322 -3522 3322 -3489
<< nsubdiff >>
rect -3322 3089 3322 3122
rect -3322 3055 -3145 3089
rect -3111 3055 -3077 3089
rect -3043 3055 -3009 3089
rect -2975 3055 -2941 3089
rect -2907 3055 -2873 3089
rect -2839 3055 -2805 3089
rect -2771 3055 -2737 3089
rect -2703 3055 -2669 3089
rect -2635 3055 -2601 3089
rect -2567 3055 -2533 3089
rect -2499 3055 -2465 3089
rect -2431 3055 -2397 3089
rect -2363 3055 -2329 3089
rect -2295 3055 -2261 3089
rect -2227 3055 -2193 3089
rect -2159 3055 -2125 3089
rect -2091 3055 -2057 3089
rect -2023 3055 -1989 3089
rect -1955 3055 -1921 3089
rect -1887 3055 -1853 3089
rect -1819 3055 -1785 3089
rect -1751 3055 -1717 3089
rect -1683 3055 -1649 3089
rect -1615 3055 -1581 3089
rect -1547 3055 -1513 3089
rect -1479 3055 -1445 3089
rect -1411 3055 -1377 3089
rect -1343 3055 -1309 3089
rect -1275 3055 -1241 3089
rect -1207 3055 -1173 3089
rect -1139 3055 -1105 3089
rect -1071 3055 -1037 3089
rect -1003 3055 -969 3089
rect -935 3055 -901 3089
rect -867 3055 -833 3089
rect -799 3055 -765 3089
rect -731 3055 -697 3089
rect -663 3055 -629 3089
rect -595 3055 -561 3089
rect -527 3055 -493 3089
rect -459 3055 -425 3089
rect -391 3055 -357 3089
rect -323 3055 -289 3089
rect -255 3055 -221 3089
rect -187 3055 -153 3089
rect -119 3055 -85 3089
rect -51 3055 -17 3089
rect 17 3055 51 3089
rect 85 3055 119 3089
rect 153 3055 187 3089
rect 221 3055 255 3089
rect 289 3055 323 3089
rect 357 3055 391 3089
rect 425 3055 459 3089
rect 493 3055 527 3089
rect 561 3055 595 3089
rect 629 3055 663 3089
rect 697 3055 731 3089
rect 765 3055 799 3089
rect 833 3055 867 3089
rect 901 3055 935 3089
rect 969 3055 1003 3089
rect 1037 3055 1071 3089
rect 1105 3055 1139 3089
rect 1173 3055 1207 3089
rect 1241 3055 1275 3089
rect 1309 3055 1343 3089
rect 1377 3055 1411 3089
rect 1445 3055 1479 3089
rect 1513 3055 1547 3089
rect 1581 3055 1615 3089
rect 1649 3055 1683 3089
rect 1717 3055 1751 3089
rect 1785 3055 1819 3089
rect 1853 3055 1887 3089
rect 1921 3055 1955 3089
rect 1989 3055 2023 3089
rect 2057 3055 2091 3089
rect 2125 3055 2159 3089
rect 2193 3055 2227 3089
rect 2261 3055 2295 3089
rect 2329 3055 2363 3089
rect 2397 3055 2431 3089
rect 2465 3055 2499 3089
rect 2533 3055 2567 3089
rect 2601 3055 2635 3089
rect 2669 3055 2703 3089
rect 2737 3055 2771 3089
rect 2805 3055 2839 3089
rect 2873 3055 2907 3089
rect 2941 3055 2975 3089
rect 3009 3055 3043 3089
rect 3077 3055 3111 3089
rect 3145 3055 3322 3089
rect -3322 3022 3322 3055
rect -3322 2941 -3222 3022
rect -3322 2907 -3289 2941
rect -3255 2907 -3222 2941
rect -3322 2873 -3222 2907
rect -3322 2839 -3289 2873
rect -3255 2839 -3222 2873
rect -3322 2805 -3222 2839
rect -3322 2771 -3289 2805
rect -3255 2771 -3222 2805
rect -3322 2737 -3222 2771
rect -3322 2703 -3289 2737
rect -3255 2703 -3222 2737
rect -3322 2669 -3222 2703
rect -3322 2635 -3289 2669
rect -3255 2635 -3222 2669
rect -3322 2601 -3222 2635
rect -3322 2567 -3289 2601
rect -3255 2567 -3222 2601
rect -3322 2533 -3222 2567
rect -3322 2499 -3289 2533
rect -3255 2499 -3222 2533
rect -3322 2465 -3222 2499
rect -3322 2431 -3289 2465
rect -3255 2431 -3222 2465
rect -3322 2397 -3222 2431
rect -3322 2363 -3289 2397
rect -3255 2363 -3222 2397
rect -3322 2329 -3222 2363
rect -3322 2295 -3289 2329
rect -3255 2295 -3222 2329
rect -3322 2261 -3222 2295
rect -3322 2227 -3289 2261
rect -3255 2227 -3222 2261
rect -3322 2193 -3222 2227
rect -3322 2159 -3289 2193
rect -3255 2159 -3222 2193
rect -3322 2125 -3222 2159
rect -3322 2091 -3289 2125
rect -3255 2091 -3222 2125
rect -3322 2057 -3222 2091
rect -3322 2023 -3289 2057
rect -3255 2023 -3222 2057
rect -3322 1989 -3222 2023
rect -3322 1955 -3289 1989
rect -3255 1955 -3222 1989
rect -3322 1921 -3222 1955
rect -3322 1887 -3289 1921
rect -3255 1887 -3222 1921
rect -3322 1853 -3222 1887
rect -3322 1819 -3289 1853
rect -3255 1819 -3222 1853
rect -3322 1785 -3222 1819
rect -3322 1751 -3289 1785
rect -3255 1751 -3222 1785
rect -3322 1717 -3222 1751
rect -3322 1683 -3289 1717
rect -3255 1683 -3222 1717
rect -3322 1649 -3222 1683
rect -3322 1615 -3289 1649
rect -3255 1615 -3222 1649
rect -3322 1581 -3222 1615
rect -3322 1547 -3289 1581
rect -3255 1547 -3222 1581
rect -3322 1513 -3222 1547
rect -3322 1479 -3289 1513
rect -3255 1479 -3222 1513
rect -3322 1445 -3222 1479
rect -3322 1411 -3289 1445
rect -3255 1411 -3222 1445
rect -3322 1377 -3222 1411
rect -3322 1343 -3289 1377
rect -3255 1343 -3222 1377
rect -3322 1309 -3222 1343
rect -3322 1275 -3289 1309
rect -3255 1275 -3222 1309
rect -3322 1241 -3222 1275
rect -3322 1207 -3289 1241
rect -3255 1207 -3222 1241
rect -3322 1173 -3222 1207
rect -3322 1139 -3289 1173
rect -3255 1139 -3222 1173
rect -3322 1105 -3222 1139
rect -3322 1071 -3289 1105
rect -3255 1071 -3222 1105
rect -3322 1037 -3222 1071
rect -3322 1003 -3289 1037
rect -3255 1003 -3222 1037
rect -3322 969 -3222 1003
rect -3322 935 -3289 969
rect -3255 935 -3222 969
rect -3322 901 -3222 935
rect -3322 867 -3289 901
rect -3255 867 -3222 901
rect -3322 833 -3222 867
rect -3322 799 -3289 833
rect -3255 799 -3222 833
rect -3322 718 -3222 799
rect 3222 2941 3322 3022
rect 3222 2907 3255 2941
rect 3289 2907 3322 2941
rect 3222 2873 3322 2907
rect 3222 2839 3255 2873
rect 3289 2839 3322 2873
rect 3222 2805 3322 2839
rect 3222 2771 3255 2805
rect 3289 2771 3322 2805
rect 3222 2737 3322 2771
rect 3222 2703 3255 2737
rect 3289 2703 3322 2737
rect 3222 2669 3322 2703
rect 3222 2635 3255 2669
rect 3289 2635 3322 2669
rect 3222 2601 3322 2635
rect 3222 2567 3255 2601
rect 3289 2567 3322 2601
rect 3222 2533 3322 2567
rect 3222 2499 3255 2533
rect 3289 2499 3322 2533
rect 3222 2465 3322 2499
rect 3222 2431 3255 2465
rect 3289 2431 3322 2465
rect 3222 2397 3322 2431
rect 3222 2363 3255 2397
rect 3289 2363 3322 2397
rect 3222 2329 3322 2363
rect 3222 2295 3255 2329
rect 3289 2295 3322 2329
rect 3222 2261 3322 2295
rect 3222 2227 3255 2261
rect 3289 2227 3322 2261
rect 3222 2193 3322 2227
rect 3222 2159 3255 2193
rect 3289 2159 3322 2193
rect 3222 2125 3322 2159
rect 3222 2091 3255 2125
rect 3289 2091 3322 2125
rect 3222 2057 3322 2091
rect 3222 2023 3255 2057
rect 3289 2023 3322 2057
rect 3222 1989 3322 2023
rect 3222 1955 3255 1989
rect 3289 1955 3322 1989
rect 3222 1921 3322 1955
rect 3222 1887 3255 1921
rect 3289 1887 3322 1921
rect 3222 1853 3322 1887
rect 3222 1819 3255 1853
rect 3289 1819 3322 1853
rect 3222 1785 3322 1819
rect 3222 1751 3255 1785
rect 3289 1751 3322 1785
rect 3222 1717 3322 1751
rect 3222 1683 3255 1717
rect 3289 1683 3322 1717
rect 3222 1649 3322 1683
rect 3222 1615 3255 1649
rect 3289 1615 3322 1649
rect 3222 1581 3322 1615
rect 3222 1547 3255 1581
rect 3289 1547 3322 1581
rect 3222 1513 3322 1547
rect 3222 1479 3255 1513
rect 3289 1479 3322 1513
rect 3222 1445 3322 1479
rect 3222 1411 3255 1445
rect 3289 1411 3322 1445
rect 3222 1377 3322 1411
rect 3222 1343 3255 1377
rect 3289 1343 3322 1377
rect 3222 1309 3322 1343
rect 3222 1275 3255 1309
rect 3289 1275 3322 1309
rect 3222 1241 3322 1275
rect 3222 1207 3255 1241
rect 3289 1207 3322 1241
rect 3222 1173 3322 1207
rect 3222 1139 3255 1173
rect 3289 1139 3322 1173
rect 3222 1105 3322 1139
rect 3222 1071 3255 1105
rect 3289 1071 3322 1105
rect 3222 1037 3322 1071
rect 3222 1003 3255 1037
rect 3289 1003 3322 1037
rect 3222 969 3322 1003
rect 3222 935 3255 969
rect 3289 935 3322 969
rect 3222 901 3322 935
rect 3222 867 3255 901
rect 3289 867 3322 901
rect 3222 833 3322 867
rect 3222 799 3255 833
rect 3289 799 3322 833
rect 3222 718 3322 799
rect -3322 685 3322 718
rect -3322 651 -3145 685
rect -3111 651 -3077 685
rect -3043 651 -3009 685
rect -2975 651 -2941 685
rect -2907 651 -2873 685
rect -2839 651 -2805 685
rect -2771 651 -2737 685
rect -2703 651 -2669 685
rect -2635 651 -2601 685
rect -2567 651 -2533 685
rect -2499 651 -2465 685
rect -2431 651 -2397 685
rect -2363 651 -2329 685
rect -2295 651 -2261 685
rect -2227 651 -2193 685
rect -2159 651 -2125 685
rect -2091 651 -2057 685
rect -2023 651 -1989 685
rect -1955 651 -1921 685
rect -1887 651 -1853 685
rect -1819 651 -1785 685
rect -1751 651 -1717 685
rect -1683 651 -1649 685
rect -1615 651 -1581 685
rect -1547 651 -1513 685
rect -1479 651 -1445 685
rect -1411 651 -1377 685
rect -1343 651 -1309 685
rect -1275 651 -1241 685
rect -1207 651 -1173 685
rect -1139 651 -1105 685
rect -1071 651 -1037 685
rect -1003 651 -969 685
rect -935 651 -901 685
rect -867 651 -833 685
rect -799 651 -765 685
rect -731 651 -697 685
rect -663 651 -629 685
rect -595 651 -561 685
rect -527 651 -493 685
rect -459 651 -425 685
rect -391 651 -357 685
rect -323 651 -289 685
rect -255 651 -221 685
rect -187 651 -153 685
rect -119 651 -85 685
rect -51 651 -17 685
rect 17 651 51 685
rect 85 651 119 685
rect 153 651 187 685
rect 221 651 255 685
rect 289 651 323 685
rect 357 651 391 685
rect 425 651 459 685
rect 493 651 527 685
rect 561 651 595 685
rect 629 651 663 685
rect 697 651 731 685
rect 765 651 799 685
rect 833 651 867 685
rect 901 651 935 685
rect 969 651 1003 685
rect 1037 651 1071 685
rect 1105 651 1139 685
rect 1173 651 1207 685
rect 1241 651 1275 685
rect 1309 651 1343 685
rect 1377 651 1411 685
rect 1445 651 1479 685
rect 1513 651 1547 685
rect 1581 651 1615 685
rect 1649 651 1683 685
rect 1717 651 1751 685
rect 1785 651 1819 685
rect 1853 651 1887 685
rect 1921 651 1955 685
rect 1989 651 2023 685
rect 2057 651 2091 685
rect 2125 651 2159 685
rect 2193 651 2227 685
rect 2261 651 2295 685
rect 2329 651 2363 685
rect 2397 651 2431 685
rect 2465 651 2499 685
rect 2533 651 2567 685
rect 2601 651 2635 685
rect 2669 651 2703 685
rect 2737 651 2771 685
rect 2805 651 2839 685
rect 2873 651 2907 685
rect 2941 651 2975 685
rect 3009 651 3043 685
rect 3077 651 3111 685
rect 3145 651 3322 685
rect -3322 618 3322 651
<< psubdiffcont >>
rect -3145 315 -3111 349
rect -3077 315 -3043 349
rect -3009 315 -2975 349
rect -2941 315 -2907 349
rect -2873 315 -2839 349
rect -2805 315 -2771 349
rect -2737 315 -2703 349
rect -2669 315 -2635 349
rect -2601 315 -2567 349
rect -2533 315 -2499 349
rect -2465 315 -2431 349
rect -2397 315 -2363 349
rect -2329 315 -2295 349
rect -2261 315 -2227 349
rect -2193 315 -2159 349
rect -2125 315 -2091 349
rect -2057 315 -2023 349
rect -1989 315 -1955 349
rect -1921 315 -1887 349
rect -1853 315 -1819 349
rect -1785 315 -1751 349
rect -1717 315 -1683 349
rect -1649 315 -1615 349
rect -1581 315 -1547 349
rect -1513 315 -1479 349
rect -1445 315 -1411 349
rect -1377 315 -1343 349
rect -1309 315 -1275 349
rect -1241 315 -1207 349
rect -1173 315 -1139 349
rect -1105 315 -1071 349
rect -1037 315 -1003 349
rect -969 315 -935 349
rect -901 315 -867 349
rect -833 315 -799 349
rect -765 315 -731 349
rect -697 315 -663 349
rect -629 315 -595 349
rect -561 315 -527 349
rect -493 315 -459 349
rect -425 315 -391 349
rect -357 315 -323 349
rect -289 315 -255 349
rect -221 315 -187 349
rect -153 315 -119 349
rect -85 315 -51 349
rect -17 315 17 349
rect 51 315 85 349
rect 119 315 153 349
rect 187 315 221 349
rect 255 315 289 349
rect 323 315 357 349
rect 391 315 425 349
rect 459 315 493 349
rect 527 315 561 349
rect 595 315 629 349
rect 663 315 697 349
rect 731 315 765 349
rect 799 315 833 349
rect 867 315 901 349
rect 935 315 969 349
rect 1003 315 1037 349
rect 1071 315 1105 349
rect 1139 315 1173 349
rect 1207 315 1241 349
rect 1275 315 1309 349
rect 1343 315 1377 349
rect 1411 315 1445 349
rect 1479 315 1513 349
rect 1547 315 1581 349
rect 1615 315 1649 349
rect 1683 315 1717 349
rect 1751 315 1785 349
rect 1819 315 1853 349
rect 1887 315 1921 349
rect 1955 315 1989 349
rect 2023 315 2057 349
rect 2091 315 2125 349
rect 2159 315 2193 349
rect 2227 315 2261 349
rect 2295 315 2329 349
rect 2363 315 2397 349
rect 2431 315 2465 349
rect 2499 315 2533 349
rect 2567 315 2601 349
rect 2635 315 2669 349
rect 2703 315 2737 349
rect 2771 315 2805 349
rect 2839 315 2873 349
rect 2907 315 2941 349
rect 2975 315 3009 349
rect 3043 315 3077 349
rect 3111 315 3145 349
rect -3289 181 -3255 215
rect -3289 113 -3255 147
rect -3289 45 -3255 79
rect -3289 -23 -3255 11
rect -3289 -91 -3255 -57
rect -3289 -159 -3255 -125
rect -3289 -227 -3255 -193
rect -3289 -295 -3255 -261
rect -3289 -363 -3255 -329
rect -3289 -431 -3255 -397
rect -3289 -499 -3255 -465
rect -3289 -567 -3255 -533
rect -3289 -635 -3255 -601
rect -3289 -703 -3255 -669
rect -3289 -771 -3255 -737
rect -3289 -839 -3255 -805
rect -3289 -907 -3255 -873
rect -3289 -975 -3255 -941
rect -3289 -1043 -3255 -1009
rect -3289 -1111 -3255 -1077
rect -2943 115 -2909 149
rect -2875 115 -2841 149
rect -2807 115 -2773 149
rect -2739 115 -2705 149
rect -2671 115 -2637 149
rect -2603 115 -2569 149
rect -2535 115 -2501 149
rect -2467 115 -2433 149
rect -2399 115 -2365 149
rect -2331 115 -2297 149
rect -2263 115 -2229 149
rect -2195 115 -2161 149
rect -2127 115 -2093 149
rect -2059 115 -2025 149
rect -1991 115 -1957 149
rect -1923 115 -1889 149
rect -1855 115 -1821 149
rect -1787 115 -1753 149
rect -1719 115 -1685 149
rect -1651 115 -1617 149
rect -1583 115 -1549 149
rect -1515 115 -1481 149
rect -1447 115 -1413 149
rect -1379 115 -1345 149
rect -1311 115 -1277 149
rect -1243 115 -1209 149
rect -1175 115 -1141 149
rect -1107 115 -1073 149
rect -1039 115 -1005 149
rect -971 115 -937 149
rect -903 115 -869 149
rect -835 115 -801 149
rect -767 115 -733 149
rect -699 115 -665 149
rect -631 115 -597 149
rect -563 115 -529 149
rect -495 115 -461 149
rect -427 115 -393 149
rect -359 115 -325 149
rect -291 115 -257 149
rect -3089 -35 -3055 -1
rect -3089 -103 -3055 -69
rect -3089 -171 -3055 -137
rect -3089 -239 -3055 -205
rect -3089 -307 -3055 -273
rect -3089 -375 -3055 -341
rect -3089 -443 -3055 -409
rect -3089 -511 -3055 -477
rect -3089 -579 -3055 -545
rect -3089 -647 -3055 -613
rect -3089 -715 -3055 -681
rect -3089 -783 -3055 -749
rect -3089 -851 -3055 -817
rect -3089 -919 -3055 -885
rect -145 -35 -111 -1
rect -145 -103 -111 -69
rect -145 -171 -111 -137
rect -145 -239 -111 -205
rect -145 -307 -111 -273
rect -145 -375 -111 -341
rect -145 -443 -111 -409
rect -145 -511 -111 -477
rect -145 -579 -111 -545
rect -145 -647 -111 -613
rect -145 -715 -111 -681
rect -145 -783 -111 -749
rect -145 -851 -111 -817
rect -145 -919 -111 -885
rect -2943 -1069 -2909 -1035
rect -2875 -1069 -2841 -1035
rect -2807 -1069 -2773 -1035
rect -2739 -1069 -2705 -1035
rect -2671 -1069 -2637 -1035
rect -2603 -1069 -2569 -1035
rect -2535 -1069 -2501 -1035
rect -2467 -1069 -2433 -1035
rect -2399 -1069 -2365 -1035
rect -2331 -1069 -2297 -1035
rect -2263 -1069 -2229 -1035
rect -2195 -1069 -2161 -1035
rect -2127 -1069 -2093 -1035
rect -2059 -1069 -2025 -1035
rect -1991 -1069 -1957 -1035
rect -1923 -1069 -1889 -1035
rect -1855 -1069 -1821 -1035
rect -1787 -1069 -1753 -1035
rect -1719 -1069 -1685 -1035
rect -1651 -1069 -1617 -1035
rect -1583 -1069 -1549 -1035
rect -1515 -1069 -1481 -1035
rect -1447 -1069 -1413 -1035
rect -1379 -1069 -1345 -1035
rect -1311 -1069 -1277 -1035
rect -1243 -1069 -1209 -1035
rect -1175 -1069 -1141 -1035
rect -1107 -1069 -1073 -1035
rect -1039 -1069 -1005 -1035
rect -971 -1069 -937 -1035
rect -903 -1069 -869 -1035
rect -835 -1069 -801 -1035
rect -767 -1069 -733 -1035
rect -699 -1069 -665 -1035
rect -631 -1069 -597 -1035
rect -563 -1069 -529 -1035
rect -495 -1069 -461 -1035
rect -427 -1069 -393 -1035
rect -359 -1069 -325 -1035
rect -291 -1069 -257 -1035
rect 3255 181 3289 215
rect 3255 113 3289 147
rect 3255 45 3289 79
rect 3255 -23 3289 11
rect 3255 -91 3289 -57
rect 3255 -159 3289 -125
rect 3255 -227 3289 -193
rect 3255 -295 3289 -261
rect 3255 -363 3289 -329
rect 3255 -431 3289 -397
rect 3255 -499 3289 -465
rect 3255 -567 3289 -533
rect 3255 -635 3289 -601
rect 3255 -703 3289 -669
rect 3255 -771 3289 -737
rect 3255 -839 3289 -805
rect 3255 -907 3289 -873
rect 3255 -975 3289 -941
rect 3255 -1043 3289 -1009
rect -3289 -1179 -3255 -1145
rect -3289 -1247 -3255 -1213
rect 3255 -1111 3289 -1077
rect 3255 -1179 3289 -1145
rect -3289 -1315 -3255 -1281
rect -3289 -1383 -3255 -1349
rect -3289 -1451 -3255 -1417
rect -3289 -1519 -3255 -1485
rect -3289 -1587 -3255 -1553
rect -3289 -1655 -3255 -1621
rect -3289 -1723 -3255 -1689
rect -3289 -1791 -3255 -1757
rect -3289 -1859 -3255 -1825
rect -3289 -1927 -3255 -1893
rect -3289 -1995 -3255 -1961
rect -3289 -2063 -3255 -2029
rect -3289 -2131 -3255 -2097
rect -3289 -2199 -3255 -2165
rect -3289 -2267 -3255 -2233
rect -3289 -2335 -3255 -2301
rect -3289 -2403 -3255 -2369
rect -3289 -2471 -3255 -2437
rect -3289 -2539 -3255 -2505
rect -3289 -2607 -3255 -2573
rect -3289 -2675 -3255 -2641
rect -3289 -2743 -3255 -2709
rect -2941 -1285 -2907 -1251
rect -2873 -1285 -2839 -1251
rect -2805 -1285 -2771 -1251
rect -2737 -1285 -2703 -1251
rect -2669 -1285 -2635 -1251
rect -2601 -1285 -2567 -1251
rect -2533 -1285 -2499 -1251
rect -2465 -1285 -2431 -1251
rect -2397 -1285 -2363 -1251
rect -2329 -1285 -2295 -1251
rect -2261 -1285 -2227 -1251
rect -2193 -1285 -2159 -1251
rect -2125 -1285 -2091 -1251
rect -2057 -1285 -2023 -1251
rect -1989 -1285 -1955 -1251
rect -1921 -1285 -1887 -1251
rect -1853 -1285 -1819 -1251
rect -1785 -1285 -1751 -1251
rect -1717 -1285 -1683 -1251
rect -1649 -1285 -1615 -1251
rect -1581 -1285 -1547 -1251
rect -1513 -1285 -1479 -1251
rect -1445 -1285 -1411 -1251
rect -1377 -1285 -1343 -1251
rect -1309 -1285 -1275 -1251
rect -1241 -1285 -1207 -1251
rect -1173 -1285 -1139 -1251
rect -1105 -1285 -1071 -1251
rect -1037 -1285 -1003 -1251
rect -969 -1285 -935 -1251
rect -901 -1285 -867 -1251
rect -833 -1285 -799 -1251
rect -765 -1285 -731 -1251
rect -697 -1285 -663 -1251
rect -629 -1285 -595 -1251
rect -561 -1285 -527 -1251
rect -493 -1285 -459 -1251
rect -425 -1285 -391 -1251
rect -357 -1285 -323 -1251
rect -289 -1285 -255 -1251
rect -221 -1285 -187 -1251
rect -153 -1285 -119 -1251
rect -85 -1285 -51 -1251
rect -17 -1285 17 -1251
rect 51 -1285 85 -1251
rect 119 -1285 153 -1251
rect 187 -1285 221 -1251
rect 255 -1285 289 -1251
rect 323 -1285 357 -1251
rect 391 -1285 425 -1251
rect 459 -1285 493 -1251
rect 527 -1285 561 -1251
rect 595 -1285 629 -1251
rect 663 -1285 697 -1251
rect 731 -1285 765 -1251
rect 799 -1285 833 -1251
rect 867 -1285 901 -1251
rect 935 -1285 969 -1251
rect 1003 -1285 1037 -1251
rect 1071 -1285 1105 -1251
rect 1139 -1285 1173 -1251
rect 1207 -1285 1241 -1251
rect 1275 -1285 1309 -1251
rect 1343 -1285 1377 -1251
rect 1411 -1285 1445 -1251
rect 1479 -1285 1513 -1251
rect 1547 -1285 1581 -1251
rect 1615 -1285 1649 -1251
rect 1683 -1285 1717 -1251
rect 1751 -1285 1785 -1251
rect 1819 -1285 1853 -1251
rect 1887 -1285 1921 -1251
rect 1955 -1285 1989 -1251
rect 2023 -1285 2057 -1251
rect 2091 -1285 2125 -1251
rect 2159 -1285 2193 -1251
rect 2227 -1285 2261 -1251
rect 2295 -1285 2329 -1251
rect 2363 -1285 2397 -1251
rect 2431 -1285 2465 -1251
rect 2499 -1285 2533 -1251
rect 2567 -1285 2601 -1251
rect 2635 -1285 2669 -1251
rect 2703 -1285 2737 -1251
rect 2771 -1285 2805 -1251
rect 2839 -1285 2873 -1251
rect 2907 -1285 2941 -1251
rect -3089 -1419 -3055 -1385
rect -3089 -1487 -3055 -1453
rect -3089 -1555 -3055 -1521
rect -3089 -1623 -3055 -1589
rect -3089 -1691 -3055 -1657
rect -3089 -1759 -3055 -1725
rect -3089 -1827 -3055 -1793
rect -3089 -1895 -3055 -1861
rect -3089 -1963 -3055 -1929
rect -3089 -2031 -3055 -1997
rect -3089 -2099 -3055 -2065
rect -3089 -2167 -3055 -2133
rect -3089 -2235 -3055 -2201
rect -3089 -2303 -3055 -2269
rect -3089 -2371 -3055 -2337
rect -3089 -2439 -3055 -2405
rect -3089 -2507 -3055 -2473
rect -3089 -2575 -3055 -2541
rect 3055 -1419 3089 -1385
rect 3055 -1487 3089 -1453
rect 3055 -1555 3089 -1521
rect 3055 -1623 3089 -1589
rect 3055 -1691 3089 -1657
rect 3055 -1759 3089 -1725
rect 3055 -1827 3089 -1793
rect 3055 -1895 3089 -1861
rect 3055 -1963 3089 -1929
rect 3055 -2031 3089 -1997
rect 3055 -2099 3089 -2065
rect 3055 -2167 3089 -2133
rect 3055 -2235 3089 -2201
rect 3055 -2303 3089 -2269
rect 3055 -2371 3089 -2337
rect 3055 -2439 3089 -2405
rect 3055 -2507 3089 -2473
rect 3055 -2575 3089 -2541
rect -2941 -2709 -2907 -2675
rect -2873 -2709 -2839 -2675
rect -2805 -2709 -2771 -2675
rect -2737 -2709 -2703 -2675
rect -2669 -2709 -2635 -2675
rect -2601 -2709 -2567 -2675
rect -2533 -2709 -2499 -2675
rect -2465 -2709 -2431 -2675
rect -2397 -2709 -2363 -2675
rect -2329 -2709 -2295 -2675
rect -2261 -2709 -2227 -2675
rect -2193 -2709 -2159 -2675
rect -2125 -2709 -2091 -2675
rect -2057 -2709 -2023 -2675
rect -1989 -2709 -1955 -2675
rect -1921 -2709 -1887 -2675
rect -1853 -2709 -1819 -2675
rect -1785 -2709 -1751 -2675
rect -1717 -2709 -1683 -2675
rect -1649 -2709 -1615 -2675
rect -1581 -2709 -1547 -2675
rect -1513 -2709 -1479 -2675
rect -1445 -2709 -1411 -2675
rect -1377 -2709 -1343 -2675
rect -1309 -2709 -1275 -2675
rect -1241 -2709 -1207 -2675
rect -1173 -2709 -1139 -2675
rect -1105 -2709 -1071 -2675
rect -1037 -2709 -1003 -2675
rect -969 -2709 -935 -2675
rect -901 -2709 -867 -2675
rect -833 -2709 -799 -2675
rect -765 -2709 -731 -2675
rect -697 -2709 -663 -2675
rect -629 -2709 -595 -2675
rect -561 -2709 -527 -2675
rect -493 -2709 -459 -2675
rect -425 -2709 -391 -2675
rect -357 -2709 -323 -2675
rect -289 -2709 -255 -2675
rect -221 -2709 -187 -2675
rect -153 -2709 -119 -2675
rect -85 -2709 -51 -2675
rect -17 -2709 17 -2675
rect 51 -2709 85 -2675
rect 119 -2709 153 -2675
rect 187 -2709 221 -2675
rect 255 -2709 289 -2675
rect 323 -2709 357 -2675
rect 391 -2709 425 -2675
rect 459 -2709 493 -2675
rect 527 -2709 561 -2675
rect 595 -2709 629 -2675
rect 663 -2709 697 -2675
rect 731 -2709 765 -2675
rect 799 -2709 833 -2675
rect 867 -2709 901 -2675
rect 935 -2709 969 -2675
rect 1003 -2709 1037 -2675
rect 1071 -2709 1105 -2675
rect 1139 -2709 1173 -2675
rect 1207 -2709 1241 -2675
rect 1275 -2709 1309 -2675
rect 1343 -2709 1377 -2675
rect 1411 -2709 1445 -2675
rect 1479 -2709 1513 -2675
rect 1547 -2709 1581 -2675
rect 1615 -2709 1649 -2675
rect 1683 -2709 1717 -2675
rect 1751 -2709 1785 -2675
rect 1819 -2709 1853 -2675
rect 1887 -2709 1921 -2675
rect 1955 -2709 1989 -2675
rect 2023 -2709 2057 -2675
rect 2091 -2709 2125 -2675
rect 2159 -2709 2193 -2675
rect 2227 -2709 2261 -2675
rect 2295 -2709 2329 -2675
rect 2363 -2709 2397 -2675
rect 2431 -2709 2465 -2675
rect 2499 -2709 2533 -2675
rect 2567 -2709 2601 -2675
rect 2635 -2709 2669 -2675
rect 2703 -2709 2737 -2675
rect 2771 -2709 2805 -2675
rect 2839 -2709 2873 -2675
rect 2907 -2709 2941 -2675
rect 3255 -1247 3289 -1213
rect 3255 -1315 3289 -1281
rect 3255 -1383 3289 -1349
rect 3255 -1451 3289 -1417
rect 3255 -1519 3289 -1485
rect 3255 -1587 3289 -1553
rect 3255 -1655 3289 -1621
rect 3255 -1723 3289 -1689
rect 3255 -1791 3289 -1757
rect 3255 -1859 3289 -1825
rect 3255 -1927 3289 -1893
rect 3255 -1995 3289 -1961
rect 3255 -2063 3289 -2029
rect 3255 -2131 3289 -2097
rect 3255 -2199 3289 -2165
rect 3255 -2267 3289 -2233
rect 3255 -2335 3289 -2301
rect 3255 -2403 3289 -2369
rect 3255 -2471 3289 -2437
rect 3255 -2539 3289 -2505
rect 3255 -2607 3289 -2573
rect 3255 -2675 3289 -2641
rect -3289 -2811 -3255 -2777
rect -3289 -2879 -3255 -2845
rect -3289 -2947 -3255 -2913
rect -3289 -3015 -3255 -2981
rect -3289 -3083 -3255 -3049
rect -3289 -3151 -3255 -3117
rect -3289 -3219 -3255 -3185
rect -3289 -3287 -3255 -3253
rect -3289 -3355 -3255 -3321
rect 3255 -2743 3289 -2709
rect 3255 -2811 3289 -2777
rect 3255 -2879 3289 -2845
rect 3255 -2947 3289 -2913
rect 3255 -3015 3289 -2981
rect 3255 -3083 3289 -3049
rect 3255 -3151 3289 -3117
rect 3255 -3219 3289 -3185
rect 3255 -3287 3289 -3253
rect 3255 -3355 3289 -3321
rect -3145 -3489 -3111 -3455
rect -3077 -3489 -3043 -3455
rect -3009 -3489 -2975 -3455
rect -2941 -3489 -2907 -3455
rect -2873 -3489 -2839 -3455
rect -2805 -3489 -2771 -3455
rect -2737 -3489 -2703 -3455
rect -2669 -3489 -2635 -3455
rect -2601 -3489 -2567 -3455
rect -2533 -3489 -2499 -3455
rect -2465 -3489 -2431 -3455
rect -2397 -3489 -2363 -3455
rect -2329 -3489 -2295 -3455
rect -2261 -3489 -2227 -3455
rect -2193 -3489 -2159 -3455
rect -2125 -3489 -2091 -3455
rect -2057 -3489 -2023 -3455
rect -1989 -3489 -1955 -3455
rect -1921 -3489 -1887 -3455
rect -1853 -3489 -1819 -3455
rect -1785 -3489 -1751 -3455
rect -1717 -3489 -1683 -3455
rect -1649 -3489 -1615 -3455
rect -1581 -3489 -1547 -3455
rect -1513 -3489 -1479 -3455
rect -1445 -3489 -1411 -3455
rect -1377 -3489 -1343 -3455
rect -1309 -3489 -1275 -3455
rect -1241 -3489 -1207 -3455
rect -1173 -3489 -1139 -3455
rect -1105 -3489 -1071 -3455
rect -1037 -3489 -1003 -3455
rect -969 -3489 -935 -3455
rect -901 -3489 -867 -3455
rect -833 -3489 -799 -3455
rect -765 -3489 -731 -3455
rect -697 -3489 -663 -3455
rect -629 -3489 -595 -3455
rect -561 -3489 -527 -3455
rect -493 -3489 -459 -3455
rect -425 -3489 -391 -3455
rect -357 -3489 -323 -3455
rect -289 -3489 -255 -3455
rect -221 -3489 -187 -3455
rect -153 -3489 -119 -3455
rect -85 -3489 -51 -3455
rect -17 -3489 17 -3455
rect 51 -3489 85 -3455
rect 119 -3489 153 -3455
rect 187 -3489 221 -3455
rect 255 -3489 289 -3455
rect 323 -3489 357 -3455
rect 391 -3489 425 -3455
rect 459 -3489 493 -3455
rect 527 -3489 561 -3455
rect 595 -3489 629 -3455
rect 663 -3489 697 -3455
rect 731 -3489 765 -3455
rect 799 -3489 833 -3455
rect 867 -3489 901 -3455
rect 935 -3489 969 -3455
rect 1003 -3489 1037 -3455
rect 1071 -3489 1105 -3455
rect 1139 -3489 1173 -3455
rect 1207 -3489 1241 -3455
rect 1275 -3489 1309 -3455
rect 1343 -3489 1377 -3455
rect 1411 -3489 1445 -3455
rect 1479 -3489 1513 -3455
rect 1547 -3489 1581 -3455
rect 1615 -3489 1649 -3455
rect 1683 -3489 1717 -3455
rect 1751 -3489 1785 -3455
rect 1819 -3489 1853 -3455
rect 1887 -3489 1921 -3455
rect 1955 -3489 1989 -3455
rect 2023 -3489 2057 -3455
rect 2091 -3489 2125 -3455
rect 2159 -3489 2193 -3455
rect 2227 -3489 2261 -3455
rect 2295 -3489 2329 -3455
rect 2363 -3489 2397 -3455
rect 2431 -3489 2465 -3455
rect 2499 -3489 2533 -3455
rect 2567 -3489 2601 -3455
rect 2635 -3489 2669 -3455
rect 2703 -3489 2737 -3455
rect 2771 -3489 2805 -3455
rect 2839 -3489 2873 -3455
rect 2907 -3489 2941 -3455
rect 2975 -3489 3009 -3455
rect 3043 -3489 3077 -3455
rect 3111 -3489 3145 -3455
<< nsubdiffcont >>
rect -3145 3055 -3111 3089
rect -3077 3055 -3043 3089
rect -3009 3055 -2975 3089
rect -2941 3055 -2907 3089
rect -2873 3055 -2839 3089
rect -2805 3055 -2771 3089
rect -2737 3055 -2703 3089
rect -2669 3055 -2635 3089
rect -2601 3055 -2567 3089
rect -2533 3055 -2499 3089
rect -2465 3055 -2431 3089
rect -2397 3055 -2363 3089
rect -2329 3055 -2295 3089
rect -2261 3055 -2227 3089
rect -2193 3055 -2159 3089
rect -2125 3055 -2091 3089
rect -2057 3055 -2023 3089
rect -1989 3055 -1955 3089
rect -1921 3055 -1887 3089
rect -1853 3055 -1819 3089
rect -1785 3055 -1751 3089
rect -1717 3055 -1683 3089
rect -1649 3055 -1615 3089
rect -1581 3055 -1547 3089
rect -1513 3055 -1479 3089
rect -1445 3055 -1411 3089
rect -1377 3055 -1343 3089
rect -1309 3055 -1275 3089
rect -1241 3055 -1207 3089
rect -1173 3055 -1139 3089
rect -1105 3055 -1071 3089
rect -1037 3055 -1003 3089
rect -969 3055 -935 3089
rect -901 3055 -867 3089
rect -833 3055 -799 3089
rect -765 3055 -731 3089
rect -697 3055 -663 3089
rect -629 3055 -595 3089
rect -561 3055 -527 3089
rect -493 3055 -459 3089
rect -425 3055 -391 3089
rect -357 3055 -323 3089
rect -289 3055 -255 3089
rect -221 3055 -187 3089
rect -153 3055 -119 3089
rect -85 3055 -51 3089
rect -17 3055 17 3089
rect 51 3055 85 3089
rect 119 3055 153 3089
rect 187 3055 221 3089
rect 255 3055 289 3089
rect 323 3055 357 3089
rect 391 3055 425 3089
rect 459 3055 493 3089
rect 527 3055 561 3089
rect 595 3055 629 3089
rect 663 3055 697 3089
rect 731 3055 765 3089
rect 799 3055 833 3089
rect 867 3055 901 3089
rect 935 3055 969 3089
rect 1003 3055 1037 3089
rect 1071 3055 1105 3089
rect 1139 3055 1173 3089
rect 1207 3055 1241 3089
rect 1275 3055 1309 3089
rect 1343 3055 1377 3089
rect 1411 3055 1445 3089
rect 1479 3055 1513 3089
rect 1547 3055 1581 3089
rect 1615 3055 1649 3089
rect 1683 3055 1717 3089
rect 1751 3055 1785 3089
rect 1819 3055 1853 3089
rect 1887 3055 1921 3089
rect 1955 3055 1989 3089
rect 2023 3055 2057 3089
rect 2091 3055 2125 3089
rect 2159 3055 2193 3089
rect 2227 3055 2261 3089
rect 2295 3055 2329 3089
rect 2363 3055 2397 3089
rect 2431 3055 2465 3089
rect 2499 3055 2533 3089
rect 2567 3055 2601 3089
rect 2635 3055 2669 3089
rect 2703 3055 2737 3089
rect 2771 3055 2805 3089
rect 2839 3055 2873 3089
rect 2907 3055 2941 3089
rect 2975 3055 3009 3089
rect 3043 3055 3077 3089
rect 3111 3055 3145 3089
rect -3289 2907 -3255 2941
rect -3289 2839 -3255 2873
rect -3289 2771 -3255 2805
rect -3289 2703 -3255 2737
rect -3289 2635 -3255 2669
rect -3289 2567 -3255 2601
rect -3289 2499 -3255 2533
rect -3289 2431 -3255 2465
rect -3289 2363 -3255 2397
rect -3289 2295 -3255 2329
rect -3289 2227 -3255 2261
rect -3289 2159 -3255 2193
rect -3289 2091 -3255 2125
rect -3289 2023 -3255 2057
rect -3289 1955 -3255 1989
rect -3289 1887 -3255 1921
rect -3289 1819 -3255 1853
rect -3289 1751 -3255 1785
rect -3289 1683 -3255 1717
rect -3289 1615 -3255 1649
rect -3289 1547 -3255 1581
rect -3289 1479 -3255 1513
rect -3289 1411 -3255 1445
rect -3289 1343 -3255 1377
rect -3289 1275 -3255 1309
rect -3289 1207 -3255 1241
rect -3289 1139 -3255 1173
rect -3289 1071 -3255 1105
rect -3289 1003 -3255 1037
rect -3289 935 -3255 969
rect -3289 867 -3255 901
rect -3289 799 -3255 833
rect 3255 2907 3289 2941
rect 3255 2839 3289 2873
rect 3255 2771 3289 2805
rect 3255 2703 3289 2737
rect 3255 2635 3289 2669
rect 3255 2567 3289 2601
rect 3255 2499 3289 2533
rect 3255 2431 3289 2465
rect 3255 2363 3289 2397
rect 3255 2295 3289 2329
rect 3255 2227 3289 2261
rect 3255 2159 3289 2193
rect 3255 2091 3289 2125
rect 3255 2023 3289 2057
rect 3255 1955 3289 1989
rect 3255 1887 3289 1921
rect 3255 1819 3289 1853
rect 3255 1751 3289 1785
rect 3255 1683 3289 1717
rect 3255 1615 3289 1649
rect 3255 1547 3289 1581
rect 3255 1479 3289 1513
rect 3255 1411 3289 1445
rect 3255 1343 3289 1377
rect 3255 1275 3289 1309
rect 3255 1207 3289 1241
rect 3255 1139 3289 1173
rect 3255 1071 3289 1105
rect 3255 1003 3289 1037
rect 3255 935 3289 969
rect 3255 867 3289 901
rect 3255 799 3289 833
rect -3145 651 -3111 685
rect -3077 651 -3043 685
rect -3009 651 -2975 685
rect -2941 651 -2907 685
rect -2873 651 -2839 685
rect -2805 651 -2771 685
rect -2737 651 -2703 685
rect -2669 651 -2635 685
rect -2601 651 -2567 685
rect -2533 651 -2499 685
rect -2465 651 -2431 685
rect -2397 651 -2363 685
rect -2329 651 -2295 685
rect -2261 651 -2227 685
rect -2193 651 -2159 685
rect -2125 651 -2091 685
rect -2057 651 -2023 685
rect -1989 651 -1955 685
rect -1921 651 -1887 685
rect -1853 651 -1819 685
rect -1785 651 -1751 685
rect -1717 651 -1683 685
rect -1649 651 -1615 685
rect -1581 651 -1547 685
rect -1513 651 -1479 685
rect -1445 651 -1411 685
rect -1377 651 -1343 685
rect -1309 651 -1275 685
rect -1241 651 -1207 685
rect -1173 651 -1139 685
rect -1105 651 -1071 685
rect -1037 651 -1003 685
rect -969 651 -935 685
rect -901 651 -867 685
rect -833 651 -799 685
rect -765 651 -731 685
rect -697 651 -663 685
rect -629 651 -595 685
rect -561 651 -527 685
rect -493 651 -459 685
rect -425 651 -391 685
rect -357 651 -323 685
rect -289 651 -255 685
rect -221 651 -187 685
rect -153 651 -119 685
rect -85 651 -51 685
rect -17 651 17 685
rect 51 651 85 685
rect 119 651 153 685
rect 187 651 221 685
rect 255 651 289 685
rect 323 651 357 685
rect 391 651 425 685
rect 459 651 493 685
rect 527 651 561 685
rect 595 651 629 685
rect 663 651 697 685
rect 731 651 765 685
rect 799 651 833 685
rect 867 651 901 685
rect 935 651 969 685
rect 1003 651 1037 685
rect 1071 651 1105 685
rect 1139 651 1173 685
rect 1207 651 1241 685
rect 1275 651 1309 685
rect 1343 651 1377 685
rect 1411 651 1445 685
rect 1479 651 1513 685
rect 1547 651 1581 685
rect 1615 651 1649 685
rect 1683 651 1717 685
rect 1751 651 1785 685
rect 1819 651 1853 685
rect 1887 651 1921 685
rect 1955 651 1989 685
rect 2023 651 2057 685
rect 2091 651 2125 685
rect 2159 651 2193 685
rect 2227 651 2261 685
rect 2295 651 2329 685
rect 2363 651 2397 685
rect 2431 651 2465 685
rect 2499 651 2533 685
rect 2567 651 2601 685
rect 2635 651 2669 685
rect 2703 651 2737 685
rect 2771 651 2805 685
rect 2839 651 2873 685
rect 2907 651 2941 685
rect 2975 651 3009 685
rect 3043 651 3077 685
rect 3111 651 3145 685
<< locali >>
rect -3322 3089 3322 3122
rect -3322 3055 -3221 3089
rect -3187 3055 -3149 3089
rect -3111 3055 -3077 3089
rect -3043 3055 -3009 3089
rect -2971 3055 -2941 3089
rect -2899 3055 -2873 3089
rect -2827 3055 -2805 3089
rect -2755 3055 -2737 3089
rect -2683 3055 -2669 3089
rect -2611 3055 -2601 3089
rect -2539 3055 -2533 3089
rect -2467 3055 -2465 3089
rect -2431 3055 -2429 3089
rect -2363 3055 -2357 3089
rect -2295 3055 -2285 3089
rect -2227 3055 -2213 3089
rect -2159 3055 -2141 3089
rect -2091 3055 -2069 3089
rect -2023 3055 -1997 3089
rect -1955 3055 -1925 3089
rect -1887 3055 -1853 3089
rect -1819 3055 -1785 3089
rect -1747 3055 -1717 3089
rect -1675 3055 -1649 3089
rect -1603 3055 -1581 3089
rect -1531 3055 -1513 3089
rect -1459 3055 -1445 3089
rect -1387 3055 -1377 3089
rect -1315 3055 -1309 3089
rect -1243 3055 -1241 3089
rect -1207 3055 -1205 3089
rect -1139 3055 -1133 3089
rect -1071 3055 -1061 3089
rect -1003 3055 -989 3089
rect -935 3055 -917 3089
rect -867 3055 -845 3089
rect -799 3055 -773 3089
rect -731 3055 -701 3089
rect -663 3055 -629 3089
rect -595 3055 -561 3089
rect -523 3055 -493 3089
rect -451 3055 -425 3089
rect -379 3055 -357 3089
rect -307 3055 -289 3089
rect -235 3055 -221 3089
rect -163 3055 -153 3089
rect -91 3055 -85 3089
rect -19 3055 -17 3089
rect 17 3055 19 3089
rect 85 3055 91 3089
rect 153 3055 163 3089
rect 221 3055 235 3089
rect 289 3055 307 3089
rect 357 3055 379 3089
rect 425 3055 451 3089
rect 493 3055 523 3089
rect 561 3055 595 3089
rect 629 3055 663 3089
rect 701 3055 731 3089
rect 773 3055 799 3089
rect 845 3055 867 3089
rect 917 3055 935 3089
rect 989 3055 1003 3089
rect 1061 3055 1071 3089
rect 1133 3055 1139 3089
rect 1205 3055 1207 3089
rect 1241 3055 1243 3089
rect 1309 3055 1315 3089
rect 1377 3055 1387 3089
rect 1445 3055 1459 3089
rect 1513 3055 1531 3089
rect 1581 3055 1603 3089
rect 1649 3055 1675 3089
rect 1717 3055 1747 3089
rect 1785 3055 1819 3089
rect 1853 3055 1887 3089
rect 1925 3055 1955 3089
rect 1997 3055 2023 3089
rect 2069 3055 2091 3089
rect 2141 3055 2159 3089
rect 2213 3055 2227 3089
rect 2285 3055 2295 3089
rect 2357 3055 2363 3089
rect 2429 3055 2431 3089
rect 2465 3055 2467 3089
rect 2533 3055 2539 3089
rect 2601 3055 2611 3089
rect 2669 3055 2683 3089
rect 2737 3055 2755 3089
rect 2805 3055 2827 3089
rect 2873 3055 2899 3089
rect 2941 3055 2971 3089
rect 3009 3055 3043 3089
rect 3077 3055 3111 3089
rect 3149 3055 3187 3089
rect 3221 3055 3322 3089
rect -3322 3022 3322 3055
rect -3322 2941 -3222 3022
rect -3322 2907 -3289 2941
rect -3255 2907 -3222 2941
rect -3322 2895 -3222 2907
rect -3322 2839 -3289 2895
rect -3255 2839 -3222 2895
rect -3322 2823 -3222 2839
rect -3322 2771 -3289 2823
rect -3255 2771 -3222 2823
rect -3322 2751 -3222 2771
rect -3322 2703 -3289 2751
rect -3255 2703 -3222 2751
rect -3322 2679 -3222 2703
rect -3322 2635 -3289 2679
rect -3255 2635 -3222 2679
rect -3322 2607 -3222 2635
rect -3322 2567 -3289 2607
rect -3255 2567 -3222 2607
rect -3322 2535 -3222 2567
rect -3322 2499 -3289 2535
rect -3255 2499 -3222 2535
rect -3322 2465 -3222 2499
rect -3322 2429 -3289 2465
rect -3255 2429 -3222 2465
rect -3322 2397 -3222 2429
rect -3322 2357 -3289 2397
rect -3255 2357 -3222 2397
rect -3322 2329 -3222 2357
rect -3322 2285 -3289 2329
rect -3255 2285 -3222 2329
rect -3322 2261 -3222 2285
rect -3322 2213 -3289 2261
rect -3255 2213 -3222 2261
rect -3322 2193 -3222 2213
rect -3322 2141 -3289 2193
rect -3255 2141 -3222 2193
rect -3322 2125 -3222 2141
rect -3322 2069 -3289 2125
rect -3255 2069 -3222 2125
rect -3322 2057 -3222 2069
rect -3322 1997 -3289 2057
rect -3255 1997 -3222 2057
rect -3322 1989 -3222 1997
rect -3322 1925 -3289 1989
rect -3255 1925 -3222 1989
rect -3322 1921 -3222 1925
rect -3322 1819 -3289 1921
rect -3255 1819 -3222 1921
rect -3322 1815 -3222 1819
rect -3322 1751 -3289 1815
rect -3255 1751 -3222 1815
rect -3322 1743 -3222 1751
rect -3322 1683 -3289 1743
rect -3255 1683 -3222 1743
rect -3322 1671 -3222 1683
rect -3322 1615 -3289 1671
rect -3255 1615 -3222 1671
rect -3322 1599 -3222 1615
rect -3322 1547 -3289 1599
rect -3255 1547 -3222 1599
rect -3322 1527 -3222 1547
rect -3322 1479 -3289 1527
rect -3255 1479 -3222 1527
rect -3322 1455 -3222 1479
rect -3322 1411 -3289 1455
rect -3255 1411 -3222 1455
rect -3322 1383 -3222 1411
rect -3322 1343 -3289 1383
rect -3255 1343 -3222 1383
rect -3322 1311 -3222 1343
rect -3322 1275 -3289 1311
rect -3255 1275 -3222 1311
rect -3322 1241 -3222 1275
rect -3322 1205 -3289 1241
rect -3255 1205 -3222 1241
rect -3322 1173 -3222 1205
rect -3322 1133 -3289 1173
rect -3255 1133 -3222 1173
rect -3322 1105 -3222 1133
rect -3322 1061 -3289 1105
rect -3255 1061 -3222 1105
rect -3322 1037 -3222 1061
rect -3322 989 -3289 1037
rect -3255 989 -3222 1037
rect -3322 969 -3222 989
rect -3322 917 -3289 969
rect -3255 917 -3222 969
rect -3322 901 -3222 917
rect -3322 845 -3289 901
rect -3255 845 -3222 901
rect -3322 833 -3222 845
rect -3322 799 -3289 833
rect -3255 799 -3222 833
rect -3322 718 -3222 799
rect 3222 2941 3322 3022
rect 3222 2907 3255 2941
rect 3289 2907 3322 2941
rect 3222 2895 3322 2907
rect 3222 2839 3255 2895
rect 3289 2839 3322 2895
rect 3222 2823 3322 2839
rect 3222 2771 3255 2823
rect 3289 2771 3322 2823
rect 3222 2751 3322 2771
rect 3222 2703 3255 2751
rect 3289 2703 3322 2751
rect 3222 2679 3322 2703
rect 3222 2635 3255 2679
rect 3289 2635 3322 2679
rect 3222 2607 3322 2635
rect 3222 2567 3255 2607
rect 3289 2567 3322 2607
rect 3222 2535 3322 2567
rect 3222 2499 3255 2535
rect 3289 2499 3322 2535
rect 3222 2465 3322 2499
rect 3222 2429 3255 2465
rect 3289 2429 3322 2465
rect 3222 2397 3322 2429
rect 3222 2357 3255 2397
rect 3289 2357 3322 2397
rect 3222 2329 3322 2357
rect 3222 2285 3255 2329
rect 3289 2285 3322 2329
rect 3222 2261 3322 2285
rect 3222 2213 3255 2261
rect 3289 2213 3322 2261
rect 3222 2193 3322 2213
rect 3222 2141 3255 2193
rect 3289 2141 3322 2193
rect 3222 2125 3322 2141
rect 3222 2069 3255 2125
rect 3289 2069 3322 2125
rect 3222 2057 3322 2069
rect 3222 1997 3255 2057
rect 3289 1997 3322 2057
rect 3222 1989 3322 1997
rect 3222 1925 3255 1989
rect 3289 1925 3322 1989
rect 3222 1921 3322 1925
rect 3222 1819 3255 1921
rect 3289 1819 3322 1921
rect 3222 1815 3322 1819
rect 3222 1751 3255 1815
rect 3289 1751 3322 1815
rect 3222 1743 3322 1751
rect 3222 1683 3255 1743
rect 3289 1683 3322 1743
rect 3222 1671 3322 1683
rect 3222 1615 3255 1671
rect 3289 1615 3322 1671
rect 3222 1599 3322 1615
rect 3222 1547 3255 1599
rect 3289 1547 3322 1599
rect 3222 1527 3322 1547
rect 3222 1479 3255 1527
rect 3289 1479 3322 1527
rect 3222 1455 3322 1479
rect 3222 1411 3255 1455
rect 3289 1411 3322 1455
rect 3222 1383 3322 1411
rect 3222 1343 3255 1383
rect 3289 1343 3322 1383
rect 3222 1311 3322 1343
rect 3222 1275 3255 1311
rect 3289 1275 3322 1311
rect 3222 1241 3322 1275
rect 3222 1205 3255 1241
rect 3289 1205 3322 1241
rect 3222 1173 3322 1205
rect 3222 1133 3255 1173
rect 3289 1133 3322 1173
rect 3222 1105 3322 1133
rect 3222 1061 3255 1105
rect 3289 1061 3322 1105
rect 3222 1037 3322 1061
rect 3222 989 3255 1037
rect 3289 989 3322 1037
rect 3222 969 3322 989
rect 3222 917 3255 969
rect 3289 917 3322 969
rect 3222 901 3322 917
rect 3222 845 3255 901
rect 3289 845 3322 901
rect 3222 833 3322 845
rect 3222 799 3255 833
rect 3289 799 3322 833
rect 3222 718 3322 799
rect -3322 685 3322 718
rect -3322 651 -3221 685
rect -3187 651 -3149 685
rect -3111 651 -3077 685
rect -3043 651 -3009 685
rect -2971 651 -2941 685
rect -2899 651 -2873 685
rect -2827 651 -2805 685
rect -2755 651 -2737 685
rect -2683 651 -2669 685
rect -2611 651 -2601 685
rect -2539 651 -2533 685
rect -2467 651 -2465 685
rect -2431 651 -2429 685
rect -2363 651 -2357 685
rect -2295 651 -2285 685
rect -2227 651 -2213 685
rect -2159 651 -2141 685
rect -2091 651 -2069 685
rect -2023 651 -1997 685
rect -1955 651 -1925 685
rect -1887 651 -1853 685
rect -1819 651 -1785 685
rect -1747 651 -1717 685
rect -1675 651 -1649 685
rect -1603 651 -1581 685
rect -1531 651 -1513 685
rect -1459 651 -1445 685
rect -1387 651 -1377 685
rect -1315 651 -1309 685
rect -1243 651 -1241 685
rect -1207 651 -1205 685
rect -1139 651 -1133 685
rect -1071 651 -1061 685
rect -1003 651 -989 685
rect -935 651 -917 685
rect -867 651 -845 685
rect -799 651 -773 685
rect -731 651 -701 685
rect -663 651 -629 685
rect -595 651 -561 685
rect -523 651 -493 685
rect -451 651 -425 685
rect -379 651 -357 685
rect -307 651 -289 685
rect -235 651 -221 685
rect -163 651 -153 685
rect -91 651 -85 685
rect -19 651 -17 685
rect 17 651 19 685
rect 85 651 91 685
rect 153 651 163 685
rect 221 651 235 685
rect 289 651 307 685
rect 357 651 379 685
rect 425 651 451 685
rect 493 651 523 685
rect 561 651 595 685
rect 629 651 663 685
rect 701 651 731 685
rect 773 651 799 685
rect 845 651 867 685
rect 917 651 935 685
rect 989 651 1003 685
rect 1061 651 1071 685
rect 1133 651 1139 685
rect 1205 651 1207 685
rect 1241 651 1243 685
rect 1309 651 1315 685
rect 1377 651 1387 685
rect 1445 651 1459 685
rect 1513 651 1531 685
rect 1581 651 1603 685
rect 1649 651 1675 685
rect 1717 651 1747 685
rect 1785 651 1819 685
rect 1853 651 1887 685
rect 1925 651 1955 685
rect 1997 651 2023 685
rect 2069 651 2091 685
rect 2141 651 2159 685
rect 2213 651 2227 685
rect 2285 651 2295 685
rect 2357 651 2363 685
rect 2429 651 2431 685
rect 2465 651 2467 685
rect 2533 651 2539 685
rect 2601 651 2611 685
rect 2669 651 2683 685
rect 2737 651 2755 685
rect 2805 651 2827 685
rect 2873 651 2899 685
rect 2941 651 2971 685
rect 3009 651 3043 685
rect 3077 651 3111 685
rect 3149 651 3187 685
rect 3221 651 3322 685
rect -3322 618 3322 651
rect -3322 349 3322 382
rect -3322 315 -3221 349
rect -3187 315 -3149 349
rect -3111 315 -3077 349
rect -3043 315 -3009 349
rect -2971 315 -2941 349
rect -2899 315 -2873 349
rect -2827 315 -2805 349
rect -2755 315 -2737 349
rect -2683 315 -2669 349
rect -2611 315 -2601 349
rect -2539 315 -2533 349
rect -2467 315 -2465 349
rect -2431 315 -2429 349
rect -2363 315 -2357 349
rect -2295 315 -2285 349
rect -2227 315 -2213 349
rect -2159 315 -2141 349
rect -2091 315 -2069 349
rect -2023 315 -1997 349
rect -1955 315 -1925 349
rect -1887 315 -1853 349
rect -1819 315 -1785 349
rect -1747 315 -1717 349
rect -1675 315 -1649 349
rect -1603 315 -1581 349
rect -1531 315 -1513 349
rect -1459 315 -1445 349
rect -1387 315 -1377 349
rect -1315 315 -1309 349
rect -1243 315 -1241 349
rect -1207 315 -1205 349
rect -1139 315 -1133 349
rect -1071 315 -1061 349
rect -1003 315 -989 349
rect -935 315 -917 349
rect -867 315 -845 349
rect -799 315 -773 349
rect -731 315 -701 349
rect -663 315 -629 349
rect -595 315 -561 349
rect -523 315 -493 349
rect -451 315 -425 349
rect -379 315 -357 349
rect -307 315 -289 349
rect -235 315 -221 349
rect -163 315 -153 349
rect -91 315 -85 349
rect -19 315 -17 349
rect 17 315 19 349
rect 85 315 91 349
rect 153 315 163 349
rect 221 315 235 349
rect 289 315 307 349
rect 357 315 379 349
rect 425 315 451 349
rect 493 315 523 349
rect 561 315 595 349
rect 629 315 663 349
rect 701 315 731 349
rect 773 315 799 349
rect 845 315 867 349
rect 917 315 935 349
rect 989 315 1003 349
rect 1061 315 1071 349
rect 1133 315 1139 349
rect 1205 315 1207 349
rect 1241 315 1243 349
rect 1309 315 1315 349
rect 1377 315 1387 349
rect 1445 315 1459 349
rect 1513 315 1531 349
rect 1581 315 1603 349
rect 1649 315 1675 349
rect 1717 315 1747 349
rect 1785 315 1819 349
rect 1853 315 1887 349
rect 1925 315 1955 349
rect 1997 315 2023 349
rect 2069 315 2091 349
rect 2141 315 2159 349
rect 2213 315 2227 349
rect 2285 315 2295 349
rect 2357 315 2363 349
rect 2429 315 2431 349
rect 2465 315 2467 349
rect 2533 315 2539 349
rect 2601 315 2611 349
rect 2669 315 2683 349
rect 2737 315 2755 349
rect 2805 315 2827 349
rect 2873 315 2899 349
rect 2941 315 2971 349
rect 3009 315 3043 349
rect 3077 315 3111 349
rect 3149 315 3187 349
rect 3221 315 3322 349
rect -3322 282 3322 315
rect -3322 215 -3222 282
rect -3322 181 -3289 215
rect -3255 181 -3222 215
rect 3222 215 3322 282
rect -3322 147 -3222 181
rect -3322 113 -3289 147
rect -3255 113 -3222 147
rect -3322 79 -3222 113
rect -3322 33 -3289 79
rect -3255 33 -3222 79
rect -3322 11 -3222 33
rect -3322 -39 -3289 11
rect -3255 -39 -3222 11
rect -3322 -57 -3222 -39
rect -3322 -111 -3289 -57
rect -3255 -111 -3222 -57
rect -3322 -125 -3222 -111
rect -3322 -183 -3289 -125
rect -3255 -183 -3222 -125
rect -3322 -193 -3222 -183
rect -3322 -255 -3289 -193
rect -3255 -255 -3222 -193
rect -3322 -261 -3222 -255
rect -3322 -327 -3289 -261
rect -3255 -327 -3222 -261
rect -3322 -329 -3222 -327
rect -3322 -363 -3289 -329
rect -3255 -363 -3222 -329
rect -3322 -365 -3222 -363
rect -3322 -431 -3289 -365
rect -3255 -431 -3222 -365
rect -3322 -437 -3222 -431
rect -3322 -499 -3289 -437
rect -3255 -499 -3222 -437
rect -3322 -509 -3222 -499
rect -3322 -567 -3289 -509
rect -3255 -567 -3222 -509
rect -3322 -581 -3222 -567
rect -3322 -635 -3289 -581
rect -3255 -635 -3222 -581
rect -3322 -653 -3222 -635
rect -3322 -703 -3289 -653
rect -3255 -703 -3222 -653
rect -3322 -725 -3222 -703
rect -3322 -771 -3289 -725
rect -3255 -771 -3222 -725
rect -3322 -797 -3222 -771
rect -3322 -839 -3289 -797
rect -3255 -839 -3222 -797
rect -3322 -869 -3222 -839
rect -3322 -907 -3289 -869
rect -3255 -907 -3222 -869
rect -3322 -941 -3222 -907
rect -3322 -975 -3289 -941
rect -3255 -975 -3222 -941
rect -3322 -1009 -3222 -975
rect -3322 -1047 -3289 -1009
rect -3255 -1047 -3222 -1009
rect -3322 -1077 -3222 -1047
rect -3322 -1119 -3289 -1077
rect -3255 -1119 -3222 -1077
rect -3122 149 -78 182
rect -3122 115 -3021 149
rect -2987 115 -2949 149
rect -2909 115 -2877 149
rect -2841 115 -2807 149
rect -2771 115 -2739 149
rect -2699 115 -2671 149
rect -2627 115 -2603 149
rect -2555 115 -2535 149
rect -2483 115 -2467 149
rect -2411 115 -2399 149
rect -2339 115 -2331 149
rect -2267 115 -2263 149
rect -2161 115 -2157 149
rect -2093 115 -2085 149
rect -2025 115 -2013 149
rect -1957 115 -1941 149
rect -1889 115 -1869 149
rect -1821 115 -1797 149
rect -1753 115 -1725 149
rect -1685 115 -1653 149
rect -1617 115 -1583 149
rect -1547 115 -1515 149
rect -1475 115 -1447 149
rect -1403 115 -1379 149
rect -1331 115 -1311 149
rect -1259 115 -1243 149
rect -1187 115 -1175 149
rect -1115 115 -1107 149
rect -1043 115 -1039 149
rect -937 115 -933 149
rect -869 115 -861 149
rect -801 115 -789 149
rect -733 115 -717 149
rect -665 115 -645 149
rect -597 115 -573 149
rect -529 115 -501 149
rect -461 115 -429 149
rect -393 115 -359 149
rect -323 115 -291 149
rect -251 115 -213 149
rect -179 115 -78 149
rect -3122 82 -78 115
rect -3122 25 -3022 82
rect -3122 -35 -3089 25
rect -3055 -35 -3022 25
rect -3122 -47 -3022 -35
rect -3122 -103 -3089 -47
rect -3055 -103 -3022 -47
rect -3122 -119 -3022 -103
rect -3122 -171 -3089 -119
rect -3055 -171 -3022 -119
rect -3122 -191 -3022 -171
rect -3122 -239 -3089 -191
rect -3055 -239 -3022 -191
rect -3122 -263 -3022 -239
rect -3122 -307 -3089 -263
rect -3055 -307 -3022 -263
rect -3122 -335 -3022 -307
rect -3122 -375 -3089 -335
rect -3055 -375 -3022 -335
rect -3122 -407 -3022 -375
rect -3122 -443 -3089 -407
rect -3055 -443 -3022 -407
rect -3122 -477 -3022 -443
rect -3122 -513 -3089 -477
rect -3055 -513 -3022 -477
rect -3122 -545 -3022 -513
rect -3122 -585 -3089 -545
rect -3055 -585 -3022 -545
rect -3122 -613 -3022 -585
rect -3122 -657 -3089 -613
rect -3055 -657 -3022 -613
rect -3122 -681 -3022 -657
rect -3122 -729 -3089 -681
rect -3055 -729 -3022 -681
rect -3122 -749 -3022 -729
rect -3122 -801 -3089 -749
rect -3055 -801 -3022 -749
rect -3122 -817 -3022 -801
rect -3122 -873 -3089 -817
rect -3055 -873 -3022 -817
rect -3122 -885 -3022 -873
rect -3122 -945 -3089 -885
rect -3055 -945 -3022 -885
rect -3122 -1002 -3022 -945
rect -178 25 -78 82
rect -178 -35 -145 25
rect -111 -35 -78 25
rect -178 -47 -78 -35
rect -178 -103 -145 -47
rect -111 -103 -78 -47
rect -178 -119 -78 -103
rect -178 -171 -145 -119
rect -111 -171 -78 -119
rect -178 -191 -78 -171
rect -178 -239 -145 -191
rect -111 -239 -78 -191
rect -178 -263 -78 -239
rect -178 -307 -145 -263
rect -111 -307 -78 -263
rect -178 -335 -78 -307
rect -178 -375 -145 -335
rect -111 -375 -78 -335
rect -178 -407 -78 -375
rect -178 -443 -145 -407
rect -111 -443 -78 -407
rect -178 -477 -78 -443
rect -178 -513 -145 -477
rect -111 -513 -78 -477
rect -178 -545 -78 -513
rect -178 -585 -145 -545
rect -111 -585 -78 -545
rect -178 -613 -78 -585
rect -178 -657 -145 -613
rect -111 -657 -78 -613
rect -178 -681 -78 -657
rect -178 -729 -145 -681
rect -111 -729 -78 -681
rect -178 -749 -78 -729
rect -178 -801 -145 -749
rect -111 -801 -78 -749
rect -178 -817 -78 -801
rect -178 -873 -145 -817
rect -111 -873 -78 -817
rect -178 -885 -78 -873
rect -178 -945 -145 -885
rect -111 -945 -78 -885
rect -178 -1002 -78 -945
rect -3122 -1035 -78 -1002
rect -3122 -1069 -3021 -1035
rect -2987 -1069 -2949 -1035
rect -2909 -1069 -2877 -1035
rect -2841 -1069 -2807 -1035
rect -2771 -1069 -2739 -1035
rect -2699 -1069 -2671 -1035
rect -2627 -1069 -2603 -1035
rect -2555 -1069 -2535 -1035
rect -2483 -1069 -2467 -1035
rect -2411 -1069 -2399 -1035
rect -2339 -1069 -2331 -1035
rect -2267 -1069 -2263 -1035
rect -2161 -1069 -2157 -1035
rect -2093 -1069 -2085 -1035
rect -2025 -1069 -2013 -1035
rect -1957 -1069 -1941 -1035
rect -1889 -1069 -1869 -1035
rect -1821 -1069 -1797 -1035
rect -1753 -1069 -1725 -1035
rect -1685 -1069 -1653 -1035
rect -1617 -1069 -1583 -1035
rect -1547 -1069 -1515 -1035
rect -1475 -1069 -1447 -1035
rect -1403 -1069 -1379 -1035
rect -1331 -1069 -1311 -1035
rect -1259 -1069 -1243 -1035
rect -1187 -1069 -1175 -1035
rect -1115 -1069 -1107 -1035
rect -1043 -1069 -1039 -1035
rect -937 -1069 -933 -1035
rect -869 -1069 -861 -1035
rect -801 -1069 -789 -1035
rect -733 -1069 -717 -1035
rect -665 -1069 -645 -1035
rect -597 -1069 -573 -1035
rect -529 -1069 -501 -1035
rect -461 -1069 -429 -1035
rect -393 -1069 -359 -1035
rect -323 -1069 -291 -1035
rect -251 -1069 -213 -1035
rect -179 -1069 -78 -1035
rect -3122 -1102 -78 -1069
rect 3222 181 3255 215
rect 3289 181 3322 215
rect 3222 147 3322 181
rect 3222 113 3255 147
rect 3289 113 3322 147
rect 3222 79 3322 113
rect 3222 33 3255 79
rect 3289 33 3322 79
rect 3222 11 3322 33
rect 3222 -39 3255 11
rect 3289 -39 3322 11
rect 3222 -57 3322 -39
rect 3222 -111 3255 -57
rect 3289 -111 3322 -57
rect 3222 -125 3322 -111
rect 3222 -183 3255 -125
rect 3289 -183 3322 -125
rect 3222 -193 3322 -183
rect 3222 -255 3255 -193
rect 3289 -255 3322 -193
rect 3222 -261 3322 -255
rect 3222 -327 3255 -261
rect 3289 -327 3322 -261
rect 3222 -329 3322 -327
rect 3222 -363 3255 -329
rect 3289 -363 3322 -329
rect 3222 -365 3322 -363
rect 3222 -431 3255 -365
rect 3289 -431 3322 -365
rect 3222 -437 3322 -431
rect 3222 -499 3255 -437
rect 3289 -499 3322 -437
rect 3222 -509 3322 -499
rect 3222 -567 3255 -509
rect 3289 -567 3322 -509
rect 3222 -581 3322 -567
rect 3222 -635 3255 -581
rect 3289 -635 3322 -581
rect 3222 -653 3322 -635
rect 3222 -703 3255 -653
rect 3289 -703 3322 -653
rect 3222 -725 3322 -703
rect 3222 -771 3255 -725
rect 3289 -771 3322 -725
rect 3222 -797 3322 -771
rect 3222 -839 3255 -797
rect 3289 -839 3322 -797
rect 3222 -869 3322 -839
rect 3222 -907 3255 -869
rect 3289 -907 3322 -869
rect 3222 -941 3322 -907
rect 3222 -975 3255 -941
rect 3289 -975 3322 -941
rect 3222 -1009 3322 -975
rect 3222 -1047 3255 -1009
rect 3289 -1047 3322 -1009
rect 3222 -1077 3322 -1047
rect -3322 -1145 -3222 -1119
rect -3322 -1191 -3289 -1145
rect -3255 -1191 -3222 -1145
rect -3322 -1213 -3222 -1191
rect -3322 -1263 -3289 -1213
rect -3255 -1263 -3222 -1213
rect 3222 -1119 3255 -1077
rect 3289 -1119 3322 -1077
rect 3222 -1145 3322 -1119
rect 3222 -1191 3255 -1145
rect 3289 -1191 3322 -1145
rect 3222 -1213 3322 -1191
rect -3322 -1281 -3222 -1263
rect -3322 -1335 -3289 -1281
rect -3255 -1335 -3222 -1281
rect -3322 -1349 -3222 -1335
rect -3322 -1407 -3289 -1349
rect -3255 -1407 -3222 -1349
rect -3322 -1417 -3222 -1407
rect -3322 -1479 -3289 -1417
rect -3255 -1479 -3222 -1417
rect -3322 -1485 -3222 -1479
rect -3322 -1551 -3289 -1485
rect -3255 -1551 -3222 -1485
rect -3322 -1553 -3222 -1551
rect -3322 -1587 -3289 -1553
rect -3255 -1587 -3222 -1553
rect -3322 -1589 -3222 -1587
rect -3322 -1655 -3289 -1589
rect -3255 -1655 -3222 -1589
rect -3322 -1661 -3222 -1655
rect -3322 -1723 -3289 -1661
rect -3255 -1723 -3222 -1661
rect -3322 -1733 -3222 -1723
rect -3322 -1791 -3289 -1733
rect -3255 -1791 -3222 -1733
rect -3322 -1805 -3222 -1791
rect -3322 -1859 -3289 -1805
rect -3255 -1859 -3222 -1805
rect -3322 -1877 -3222 -1859
rect -3322 -1927 -3289 -1877
rect -3255 -1927 -3222 -1877
rect -3322 -1949 -3222 -1927
rect -3322 -1995 -3289 -1949
rect -3255 -1995 -3222 -1949
rect -3322 -2021 -3222 -1995
rect -3322 -2063 -3289 -2021
rect -3255 -2063 -3222 -2021
rect -3322 -2093 -3222 -2063
rect -3322 -2131 -3289 -2093
rect -3255 -2131 -3222 -2093
rect -3322 -2165 -3222 -2131
rect -3322 -2199 -3289 -2165
rect -3255 -2199 -3222 -2165
rect -3322 -2233 -3222 -2199
rect -3322 -2271 -3289 -2233
rect -3255 -2271 -3222 -2233
rect -3322 -2301 -3222 -2271
rect -3322 -2343 -3289 -2301
rect -3255 -2343 -3222 -2301
rect -3322 -2369 -3222 -2343
rect -3322 -2415 -3289 -2369
rect -3255 -2415 -3222 -2369
rect -3322 -2437 -3222 -2415
rect -3322 -2487 -3289 -2437
rect -3255 -2487 -3222 -2437
rect -3322 -2505 -3222 -2487
rect -3322 -2559 -3289 -2505
rect -3255 -2559 -3222 -2505
rect -3322 -2573 -3222 -2559
rect -3322 -2631 -3289 -2573
rect -3255 -2631 -3222 -2573
rect -3322 -2641 -3222 -2631
rect -3322 -2703 -3289 -2641
rect -3255 -2703 -3222 -2641
rect -3322 -2709 -3222 -2703
rect -3322 -2775 -3289 -2709
rect -3255 -2775 -3222 -2709
rect -3122 -1251 3122 -1218
rect -3122 -1285 -3005 -1251
rect -2971 -1285 -2941 -1251
rect -2899 -1285 -2873 -1251
rect -2827 -1285 -2805 -1251
rect -2755 -1285 -2737 -1251
rect -2683 -1285 -2669 -1251
rect -2611 -1285 -2601 -1251
rect -2539 -1285 -2533 -1251
rect -2467 -1285 -2465 -1251
rect -2431 -1285 -2429 -1251
rect -2363 -1285 -2357 -1251
rect -2295 -1285 -2285 -1251
rect -2227 -1285 -2213 -1251
rect -2159 -1285 -2141 -1251
rect -2091 -1285 -2069 -1251
rect -2023 -1285 -1997 -1251
rect -1955 -1285 -1925 -1251
rect -1887 -1285 -1853 -1251
rect -1819 -1285 -1785 -1251
rect -1747 -1285 -1717 -1251
rect -1675 -1285 -1649 -1251
rect -1603 -1285 -1581 -1251
rect -1531 -1285 -1513 -1251
rect -1459 -1285 -1445 -1251
rect -1387 -1285 -1377 -1251
rect -1315 -1285 -1309 -1251
rect -1243 -1285 -1241 -1251
rect -1207 -1285 -1205 -1251
rect -1139 -1285 -1133 -1251
rect -1071 -1285 -1061 -1251
rect -1003 -1285 -989 -1251
rect -935 -1285 -917 -1251
rect -867 -1285 -845 -1251
rect -799 -1285 -773 -1251
rect -731 -1285 -701 -1251
rect -663 -1285 -629 -1251
rect -595 -1285 -561 -1251
rect -523 -1285 -493 -1251
rect -451 -1285 -425 -1251
rect -379 -1285 -357 -1251
rect -307 -1285 -289 -1251
rect -235 -1285 -221 -1251
rect -163 -1285 -153 -1251
rect -91 -1285 -85 -1251
rect -19 -1285 -17 -1251
rect 17 -1285 19 -1251
rect 85 -1285 91 -1251
rect 153 -1285 163 -1251
rect 221 -1285 235 -1251
rect 289 -1285 307 -1251
rect 357 -1285 379 -1251
rect 425 -1285 451 -1251
rect 493 -1285 523 -1251
rect 561 -1285 595 -1251
rect 629 -1285 663 -1251
rect 701 -1285 731 -1251
rect 773 -1285 799 -1251
rect 845 -1285 867 -1251
rect 917 -1285 935 -1251
rect 989 -1285 1003 -1251
rect 1061 -1285 1071 -1251
rect 1133 -1285 1139 -1251
rect 1205 -1285 1207 -1251
rect 1241 -1285 1243 -1251
rect 1309 -1285 1315 -1251
rect 1377 -1285 1387 -1251
rect 1445 -1285 1459 -1251
rect 1513 -1285 1531 -1251
rect 1581 -1285 1603 -1251
rect 1649 -1285 1675 -1251
rect 1717 -1285 1747 -1251
rect 1785 -1285 1819 -1251
rect 1853 -1285 1887 -1251
rect 1925 -1285 1955 -1251
rect 1997 -1285 2023 -1251
rect 2069 -1285 2091 -1251
rect 2141 -1285 2159 -1251
rect 2213 -1285 2227 -1251
rect 2285 -1285 2295 -1251
rect 2357 -1285 2363 -1251
rect 2429 -1285 2431 -1251
rect 2465 -1285 2467 -1251
rect 2533 -1285 2539 -1251
rect 2601 -1285 2611 -1251
rect 2669 -1285 2683 -1251
rect 2737 -1285 2755 -1251
rect 2805 -1285 2827 -1251
rect 2873 -1285 2899 -1251
rect 2941 -1285 2971 -1251
rect 3005 -1285 3122 -1251
rect -3122 -1318 3122 -1285
rect -3122 -1385 -3022 -1318
rect -3122 -1421 -3089 -1385
rect -3055 -1421 -3022 -1385
rect -3122 -1453 -3022 -1421
rect -3122 -1493 -3089 -1453
rect -3055 -1493 -3022 -1453
rect -3122 -1521 -3022 -1493
rect -3122 -1565 -3089 -1521
rect -3055 -1565 -3022 -1521
rect -3122 -1589 -3022 -1565
rect -3122 -1637 -3089 -1589
rect -3055 -1637 -3022 -1589
rect -3122 -1657 -3022 -1637
rect -3122 -1709 -3089 -1657
rect -3055 -1709 -3022 -1657
rect -3122 -1725 -3022 -1709
rect -3122 -1781 -3089 -1725
rect -3055 -1781 -3022 -1725
rect -3122 -1793 -3022 -1781
rect -3122 -1853 -3089 -1793
rect -3055 -1853 -3022 -1793
rect -3122 -1861 -3022 -1853
rect -3122 -1925 -3089 -1861
rect -3055 -1925 -3022 -1861
rect -3122 -1929 -3022 -1925
rect -3122 -2031 -3089 -1929
rect -3055 -2031 -3022 -1929
rect -3122 -2035 -3022 -2031
rect -3122 -2099 -3089 -2035
rect -3055 -2099 -3022 -2035
rect -3122 -2107 -3022 -2099
rect -3122 -2167 -3089 -2107
rect -3055 -2167 -3022 -2107
rect -3122 -2179 -3022 -2167
rect -3122 -2235 -3089 -2179
rect -3055 -2235 -3022 -2179
rect -3122 -2251 -3022 -2235
rect -3122 -2303 -3089 -2251
rect -3055 -2303 -3022 -2251
rect -3122 -2323 -3022 -2303
rect -3122 -2371 -3089 -2323
rect -3055 -2371 -3022 -2323
rect -3122 -2395 -3022 -2371
rect -3122 -2439 -3089 -2395
rect -3055 -2439 -3022 -2395
rect -3122 -2467 -3022 -2439
rect -3122 -2507 -3089 -2467
rect -3055 -2507 -3022 -2467
rect -3122 -2539 -3022 -2507
rect -3122 -2575 -3089 -2539
rect -3055 -2575 -3022 -2539
rect -3122 -2642 -3022 -2575
rect 3022 -1385 3122 -1318
rect 3022 -1421 3055 -1385
rect 3089 -1421 3122 -1385
rect 3022 -1453 3122 -1421
rect 3022 -1493 3055 -1453
rect 3089 -1493 3122 -1453
rect 3022 -1521 3122 -1493
rect 3022 -1565 3055 -1521
rect 3089 -1565 3122 -1521
rect 3022 -1589 3122 -1565
rect 3022 -1637 3055 -1589
rect 3089 -1637 3122 -1589
rect 3022 -1657 3122 -1637
rect 3022 -1709 3055 -1657
rect 3089 -1709 3122 -1657
rect 3022 -1725 3122 -1709
rect 3022 -1781 3055 -1725
rect 3089 -1781 3122 -1725
rect 3022 -1793 3122 -1781
rect 3022 -1853 3055 -1793
rect 3089 -1853 3122 -1793
rect 3022 -1861 3122 -1853
rect 3022 -1925 3055 -1861
rect 3089 -1925 3122 -1861
rect 3022 -1929 3122 -1925
rect 3022 -2031 3055 -1929
rect 3089 -2031 3122 -1929
rect 3022 -2035 3122 -2031
rect 3022 -2099 3055 -2035
rect 3089 -2099 3122 -2035
rect 3022 -2107 3122 -2099
rect 3022 -2167 3055 -2107
rect 3089 -2167 3122 -2107
rect 3022 -2179 3122 -2167
rect 3022 -2235 3055 -2179
rect 3089 -2235 3122 -2179
rect 3022 -2251 3122 -2235
rect 3022 -2303 3055 -2251
rect 3089 -2303 3122 -2251
rect 3022 -2323 3122 -2303
rect 3022 -2371 3055 -2323
rect 3089 -2371 3122 -2323
rect 3022 -2395 3122 -2371
rect 3022 -2439 3055 -2395
rect 3089 -2439 3122 -2395
rect 3022 -2467 3122 -2439
rect 3022 -2507 3055 -2467
rect 3089 -2507 3122 -2467
rect 3022 -2539 3122 -2507
rect 3022 -2575 3055 -2539
rect 3089 -2575 3122 -2539
rect 3022 -2642 3122 -2575
rect -3122 -2675 3122 -2642
rect -3122 -2709 -3005 -2675
rect -2971 -2709 -2941 -2675
rect -2899 -2709 -2873 -2675
rect -2827 -2709 -2805 -2675
rect -2755 -2709 -2737 -2675
rect -2683 -2709 -2669 -2675
rect -2611 -2709 -2601 -2675
rect -2539 -2709 -2533 -2675
rect -2467 -2709 -2465 -2675
rect -2431 -2709 -2429 -2675
rect -2363 -2709 -2357 -2675
rect -2295 -2709 -2285 -2675
rect -2227 -2709 -2213 -2675
rect -2159 -2709 -2141 -2675
rect -2091 -2709 -2069 -2675
rect -2023 -2709 -1997 -2675
rect -1955 -2709 -1925 -2675
rect -1887 -2709 -1853 -2675
rect -1819 -2709 -1785 -2675
rect -1747 -2709 -1717 -2675
rect -1675 -2709 -1649 -2675
rect -1603 -2709 -1581 -2675
rect -1531 -2709 -1513 -2675
rect -1459 -2709 -1445 -2675
rect -1387 -2709 -1377 -2675
rect -1315 -2709 -1309 -2675
rect -1243 -2709 -1241 -2675
rect -1207 -2709 -1205 -2675
rect -1139 -2709 -1133 -2675
rect -1071 -2709 -1061 -2675
rect -1003 -2709 -989 -2675
rect -935 -2709 -917 -2675
rect -867 -2709 -845 -2675
rect -799 -2709 -773 -2675
rect -731 -2709 -701 -2675
rect -663 -2709 -629 -2675
rect -595 -2709 -561 -2675
rect -523 -2709 -493 -2675
rect -451 -2709 -425 -2675
rect -379 -2709 -357 -2675
rect -307 -2709 -289 -2675
rect -235 -2709 -221 -2675
rect -163 -2709 -153 -2675
rect -91 -2709 -85 -2675
rect -19 -2709 -17 -2675
rect 17 -2709 19 -2675
rect 85 -2709 91 -2675
rect 153 -2709 163 -2675
rect 221 -2709 235 -2675
rect 289 -2709 307 -2675
rect 357 -2709 379 -2675
rect 425 -2709 451 -2675
rect 493 -2709 523 -2675
rect 561 -2709 595 -2675
rect 629 -2709 663 -2675
rect 701 -2709 731 -2675
rect 773 -2709 799 -2675
rect 845 -2709 867 -2675
rect 917 -2709 935 -2675
rect 989 -2709 1003 -2675
rect 1061 -2709 1071 -2675
rect 1133 -2709 1139 -2675
rect 1205 -2709 1207 -2675
rect 1241 -2709 1243 -2675
rect 1309 -2709 1315 -2675
rect 1377 -2709 1387 -2675
rect 1445 -2709 1459 -2675
rect 1513 -2709 1531 -2675
rect 1581 -2709 1603 -2675
rect 1649 -2709 1675 -2675
rect 1717 -2709 1747 -2675
rect 1785 -2709 1819 -2675
rect 1853 -2709 1887 -2675
rect 1925 -2709 1955 -2675
rect 1997 -2709 2023 -2675
rect 2069 -2709 2091 -2675
rect 2141 -2709 2159 -2675
rect 2213 -2709 2227 -2675
rect 2285 -2709 2295 -2675
rect 2357 -2709 2363 -2675
rect 2429 -2709 2431 -2675
rect 2465 -2709 2467 -2675
rect 2533 -2709 2539 -2675
rect 2601 -2709 2611 -2675
rect 2669 -2709 2683 -2675
rect 2737 -2709 2755 -2675
rect 2805 -2709 2827 -2675
rect 2873 -2709 2899 -2675
rect 2941 -2709 2971 -2675
rect 3005 -2709 3122 -2675
rect -3122 -2742 3122 -2709
rect 3222 -1263 3255 -1213
rect 3289 -1263 3322 -1213
rect 3222 -1281 3322 -1263
rect 3222 -1335 3255 -1281
rect 3289 -1335 3322 -1281
rect 3222 -1349 3322 -1335
rect 3222 -1407 3255 -1349
rect 3289 -1407 3322 -1349
rect 3222 -1417 3322 -1407
rect 3222 -1479 3255 -1417
rect 3289 -1479 3322 -1417
rect 3222 -1485 3322 -1479
rect 3222 -1551 3255 -1485
rect 3289 -1551 3322 -1485
rect 3222 -1553 3322 -1551
rect 3222 -1587 3255 -1553
rect 3289 -1587 3322 -1553
rect 3222 -1589 3322 -1587
rect 3222 -1655 3255 -1589
rect 3289 -1655 3322 -1589
rect 3222 -1661 3322 -1655
rect 3222 -1723 3255 -1661
rect 3289 -1723 3322 -1661
rect 3222 -1733 3322 -1723
rect 3222 -1791 3255 -1733
rect 3289 -1791 3322 -1733
rect 3222 -1805 3322 -1791
rect 3222 -1859 3255 -1805
rect 3289 -1859 3322 -1805
rect 3222 -1877 3322 -1859
rect 3222 -1927 3255 -1877
rect 3289 -1927 3322 -1877
rect 3222 -1949 3322 -1927
rect 3222 -1995 3255 -1949
rect 3289 -1995 3322 -1949
rect 3222 -2021 3322 -1995
rect 3222 -2063 3255 -2021
rect 3289 -2063 3322 -2021
rect 3222 -2093 3322 -2063
rect 3222 -2131 3255 -2093
rect 3289 -2131 3322 -2093
rect 3222 -2165 3322 -2131
rect 3222 -2199 3255 -2165
rect 3289 -2199 3322 -2165
rect 3222 -2233 3322 -2199
rect 3222 -2271 3255 -2233
rect 3289 -2271 3322 -2233
rect 3222 -2301 3322 -2271
rect 3222 -2343 3255 -2301
rect 3289 -2343 3322 -2301
rect 3222 -2369 3322 -2343
rect 3222 -2415 3255 -2369
rect 3289 -2415 3322 -2369
rect 3222 -2437 3322 -2415
rect 3222 -2487 3255 -2437
rect 3289 -2487 3322 -2437
rect 3222 -2505 3322 -2487
rect 3222 -2559 3255 -2505
rect 3289 -2559 3322 -2505
rect 3222 -2573 3322 -2559
rect 3222 -2631 3255 -2573
rect 3289 -2631 3322 -2573
rect 3222 -2641 3322 -2631
rect 3222 -2703 3255 -2641
rect 3289 -2703 3322 -2641
rect 3222 -2709 3322 -2703
rect -3322 -2777 -3222 -2775
rect -3322 -2811 -3289 -2777
rect -3255 -2811 -3222 -2777
rect -3322 -2813 -3222 -2811
rect -3322 -2879 -3289 -2813
rect -3255 -2879 -3222 -2813
rect -3322 -2885 -3222 -2879
rect -3322 -2947 -3289 -2885
rect -3255 -2947 -3222 -2885
rect -3322 -2957 -3222 -2947
rect -3322 -3015 -3289 -2957
rect -3255 -3015 -3222 -2957
rect -3322 -3029 -3222 -3015
rect -3322 -3083 -3289 -3029
rect -3255 -3083 -3222 -3029
rect -3322 -3101 -3222 -3083
rect -3322 -3151 -3289 -3101
rect -3255 -3151 -3222 -3101
rect -3322 -3173 -3222 -3151
rect -3322 -3219 -3289 -3173
rect -3255 -3219 -3222 -3173
rect -3322 -3253 -3222 -3219
rect -3322 -3287 -3289 -3253
rect -3255 -3287 -3222 -3253
rect -3322 -3321 -3222 -3287
rect -3322 -3355 -3289 -3321
rect -3255 -3355 -3222 -3321
rect -3322 -3422 -3222 -3355
rect 3222 -2775 3255 -2709
rect 3289 -2775 3322 -2709
rect 3222 -2777 3322 -2775
rect 3222 -2811 3255 -2777
rect 3289 -2811 3322 -2777
rect 3222 -2813 3322 -2811
rect 3222 -2879 3255 -2813
rect 3289 -2879 3322 -2813
rect 3222 -2885 3322 -2879
rect 3222 -2947 3255 -2885
rect 3289 -2947 3322 -2885
rect 3222 -2957 3322 -2947
rect 3222 -3015 3255 -2957
rect 3289 -3015 3322 -2957
rect 3222 -3029 3322 -3015
rect 3222 -3083 3255 -3029
rect 3289 -3083 3322 -3029
rect 3222 -3101 3322 -3083
rect 3222 -3151 3255 -3101
rect 3289 -3151 3322 -3101
rect 3222 -3173 3322 -3151
rect 3222 -3219 3255 -3173
rect 3289 -3219 3322 -3173
rect 3222 -3253 3322 -3219
rect 3222 -3287 3255 -3253
rect 3289 -3287 3322 -3253
rect 3222 -3321 3322 -3287
rect 3222 -3355 3255 -3321
rect 3289 -3355 3322 -3321
rect 3222 -3422 3322 -3355
rect -3322 -3455 3322 -3422
rect -3322 -3489 -3221 -3455
rect -3187 -3489 -3149 -3455
rect -3111 -3489 -3077 -3455
rect -3043 -3489 -3009 -3455
rect -2971 -3489 -2941 -3455
rect -2899 -3489 -2873 -3455
rect -2827 -3489 -2805 -3455
rect -2755 -3489 -2737 -3455
rect -2683 -3489 -2669 -3455
rect -2611 -3489 -2601 -3455
rect -2539 -3489 -2533 -3455
rect -2467 -3489 -2465 -3455
rect -2431 -3489 -2429 -3455
rect -2363 -3489 -2357 -3455
rect -2295 -3489 -2285 -3455
rect -2227 -3489 -2213 -3455
rect -2159 -3489 -2141 -3455
rect -2091 -3489 -2069 -3455
rect -2023 -3489 -1997 -3455
rect -1955 -3489 -1925 -3455
rect -1887 -3489 -1853 -3455
rect -1819 -3489 -1785 -3455
rect -1747 -3489 -1717 -3455
rect -1675 -3489 -1649 -3455
rect -1603 -3489 -1581 -3455
rect -1531 -3489 -1513 -3455
rect -1459 -3489 -1445 -3455
rect -1387 -3489 -1377 -3455
rect -1315 -3489 -1309 -3455
rect -1243 -3489 -1241 -3455
rect -1207 -3489 -1205 -3455
rect -1139 -3489 -1133 -3455
rect -1071 -3489 -1061 -3455
rect -1003 -3489 -989 -3455
rect -935 -3489 -917 -3455
rect -867 -3489 -845 -3455
rect -799 -3489 -773 -3455
rect -731 -3489 -701 -3455
rect -663 -3489 -629 -3455
rect -595 -3489 -561 -3455
rect -523 -3489 -493 -3455
rect -451 -3489 -425 -3455
rect -379 -3489 -357 -3455
rect -307 -3489 -289 -3455
rect -235 -3489 -221 -3455
rect -163 -3489 -153 -3455
rect -91 -3489 -85 -3455
rect -19 -3489 -17 -3455
rect 17 -3489 19 -3455
rect 85 -3489 91 -3455
rect 153 -3489 163 -3455
rect 221 -3489 235 -3455
rect 289 -3489 307 -3455
rect 357 -3489 379 -3455
rect 425 -3489 451 -3455
rect 493 -3489 523 -3455
rect 561 -3489 595 -3455
rect 629 -3489 663 -3455
rect 701 -3489 731 -3455
rect 773 -3489 799 -3455
rect 845 -3489 867 -3455
rect 917 -3489 935 -3455
rect 989 -3489 1003 -3455
rect 1061 -3489 1071 -3455
rect 1133 -3489 1139 -3455
rect 1205 -3489 1207 -3455
rect 1241 -3489 1243 -3455
rect 1309 -3489 1315 -3455
rect 1377 -3489 1387 -3455
rect 1445 -3489 1459 -3455
rect 1513 -3489 1531 -3455
rect 1581 -3489 1603 -3455
rect 1649 -3489 1675 -3455
rect 1717 -3489 1747 -3455
rect 1785 -3489 1819 -3455
rect 1853 -3489 1887 -3455
rect 1925 -3489 1955 -3455
rect 1997 -3489 2023 -3455
rect 2069 -3489 2091 -3455
rect 2141 -3489 2159 -3455
rect 2213 -3489 2227 -3455
rect 2285 -3489 2295 -3455
rect 2357 -3489 2363 -3455
rect 2429 -3489 2431 -3455
rect 2465 -3489 2467 -3455
rect 2533 -3489 2539 -3455
rect 2601 -3489 2611 -3455
rect 2669 -3489 2683 -3455
rect 2737 -3489 2755 -3455
rect 2805 -3489 2827 -3455
rect 2873 -3489 2899 -3455
rect 2941 -3489 2971 -3455
rect 3009 -3489 3043 -3455
rect 3077 -3489 3111 -3455
rect 3149 -3489 3187 -3455
rect 3221 -3489 3322 -3455
rect -3322 -3522 3322 -3489
<< viali >>
rect -3221 3055 -3187 3089
rect -3149 3055 -3145 3089
rect -3145 3055 -3115 3089
rect -3077 3055 -3043 3089
rect -3005 3055 -2975 3089
rect -2975 3055 -2971 3089
rect -2933 3055 -2907 3089
rect -2907 3055 -2899 3089
rect -2861 3055 -2839 3089
rect -2839 3055 -2827 3089
rect -2789 3055 -2771 3089
rect -2771 3055 -2755 3089
rect -2717 3055 -2703 3089
rect -2703 3055 -2683 3089
rect -2645 3055 -2635 3089
rect -2635 3055 -2611 3089
rect -2573 3055 -2567 3089
rect -2567 3055 -2539 3089
rect -2501 3055 -2499 3089
rect -2499 3055 -2467 3089
rect -2429 3055 -2397 3089
rect -2397 3055 -2395 3089
rect -2357 3055 -2329 3089
rect -2329 3055 -2323 3089
rect -2285 3055 -2261 3089
rect -2261 3055 -2251 3089
rect -2213 3055 -2193 3089
rect -2193 3055 -2179 3089
rect -2141 3055 -2125 3089
rect -2125 3055 -2107 3089
rect -2069 3055 -2057 3089
rect -2057 3055 -2035 3089
rect -1997 3055 -1989 3089
rect -1989 3055 -1963 3089
rect -1925 3055 -1921 3089
rect -1921 3055 -1891 3089
rect -1853 3055 -1819 3089
rect -1781 3055 -1751 3089
rect -1751 3055 -1747 3089
rect -1709 3055 -1683 3089
rect -1683 3055 -1675 3089
rect -1637 3055 -1615 3089
rect -1615 3055 -1603 3089
rect -1565 3055 -1547 3089
rect -1547 3055 -1531 3089
rect -1493 3055 -1479 3089
rect -1479 3055 -1459 3089
rect -1421 3055 -1411 3089
rect -1411 3055 -1387 3089
rect -1349 3055 -1343 3089
rect -1343 3055 -1315 3089
rect -1277 3055 -1275 3089
rect -1275 3055 -1243 3089
rect -1205 3055 -1173 3089
rect -1173 3055 -1171 3089
rect -1133 3055 -1105 3089
rect -1105 3055 -1099 3089
rect -1061 3055 -1037 3089
rect -1037 3055 -1027 3089
rect -989 3055 -969 3089
rect -969 3055 -955 3089
rect -917 3055 -901 3089
rect -901 3055 -883 3089
rect -845 3055 -833 3089
rect -833 3055 -811 3089
rect -773 3055 -765 3089
rect -765 3055 -739 3089
rect -701 3055 -697 3089
rect -697 3055 -667 3089
rect -629 3055 -595 3089
rect -557 3055 -527 3089
rect -527 3055 -523 3089
rect -485 3055 -459 3089
rect -459 3055 -451 3089
rect -413 3055 -391 3089
rect -391 3055 -379 3089
rect -341 3055 -323 3089
rect -323 3055 -307 3089
rect -269 3055 -255 3089
rect -255 3055 -235 3089
rect -197 3055 -187 3089
rect -187 3055 -163 3089
rect -125 3055 -119 3089
rect -119 3055 -91 3089
rect -53 3055 -51 3089
rect -51 3055 -19 3089
rect 19 3055 51 3089
rect 51 3055 53 3089
rect 91 3055 119 3089
rect 119 3055 125 3089
rect 163 3055 187 3089
rect 187 3055 197 3089
rect 235 3055 255 3089
rect 255 3055 269 3089
rect 307 3055 323 3089
rect 323 3055 341 3089
rect 379 3055 391 3089
rect 391 3055 413 3089
rect 451 3055 459 3089
rect 459 3055 485 3089
rect 523 3055 527 3089
rect 527 3055 557 3089
rect 595 3055 629 3089
rect 667 3055 697 3089
rect 697 3055 701 3089
rect 739 3055 765 3089
rect 765 3055 773 3089
rect 811 3055 833 3089
rect 833 3055 845 3089
rect 883 3055 901 3089
rect 901 3055 917 3089
rect 955 3055 969 3089
rect 969 3055 989 3089
rect 1027 3055 1037 3089
rect 1037 3055 1061 3089
rect 1099 3055 1105 3089
rect 1105 3055 1133 3089
rect 1171 3055 1173 3089
rect 1173 3055 1205 3089
rect 1243 3055 1275 3089
rect 1275 3055 1277 3089
rect 1315 3055 1343 3089
rect 1343 3055 1349 3089
rect 1387 3055 1411 3089
rect 1411 3055 1421 3089
rect 1459 3055 1479 3089
rect 1479 3055 1493 3089
rect 1531 3055 1547 3089
rect 1547 3055 1565 3089
rect 1603 3055 1615 3089
rect 1615 3055 1637 3089
rect 1675 3055 1683 3089
rect 1683 3055 1709 3089
rect 1747 3055 1751 3089
rect 1751 3055 1781 3089
rect 1819 3055 1853 3089
rect 1891 3055 1921 3089
rect 1921 3055 1925 3089
rect 1963 3055 1989 3089
rect 1989 3055 1997 3089
rect 2035 3055 2057 3089
rect 2057 3055 2069 3089
rect 2107 3055 2125 3089
rect 2125 3055 2141 3089
rect 2179 3055 2193 3089
rect 2193 3055 2213 3089
rect 2251 3055 2261 3089
rect 2261 3055 2285 3089
rect 2323 3055 2329 3089
rect 2329 3055 2357 3089
rect 2395 3055 2397 3089
rect 2397 3055 2429 3089
rect 2467 3055 2499 3089
rect 2499 3055 2501 3089
rect 2539 3055 2567 3089
rect 2567 3055 2573 3089
rect 2611 3055 2635 3089
rect 2635 3055 2645 3089
rect 2683 3055 2703 3089
rect 2703 3055 2717 3089
rect 2755 3055 2771 3089
rect 2771 3055 2789 3089
rect 2827 3055 2839 3089
rect 2839 3055 2861 3089
rect 2899 3055 2907 3089
rect 2907 3055 2933 3089
rect 2971 3055 2975 3089
rect 2975 3055 3005 3089
rect 3043 3055 3077 3089
rect 3115 3055 3145 3089
rect 3145 3055 3149 3089
rect 3187 3055 3221 3089
rect -3289 2873 -3255 2895
rect -3289 2861 -3255 2873
rect -3289 2805 -3255 2823
rect -3289 2789 -3255 2805
rect -3289 2737 -3255 2751
rect -3289 2717 -3255 2737
rect -3289 2669 -3255 2679
rect -3289 2645 -3255 2669
rect -3289 2601 -3255 2607
rect -3289 2573 -3255 2601
rect -3289 2533 -3255 2535
rect -3289 2501 -3255 2533
rect -3289 2431 -3255 2463
rect -3289 2429 -3255 2431
rect -3289 2363 -3255 2391
rect -3289 2357 -3255 2363
rect -3289 2295 -3255 2319
rect -3289 2285 -3255 2295
rect -3289 2227 -3255 2247
rect -3289 2213 -3255 2227
rect -3289 2159 -3255 2175
rect -3289 2141 -3255 2159
rect -3289 2091 -3255 2103
rect -3289 2069 -3255 2091
rect -3289 2023 -3255 2031
rect -3289 1997 -3255 2023
rect -3289 1955 -3255 1959
rect -3289 1925 -3255 1955
rect -3289 1853 -3255 1887
rect -3289 1785 -3255 1815
rect -3289 1781 -3255 1785
rect -3289 1717 -3255 1743
rect -3289 1709 -3255 1717
rect -3289 1649 -3255 1671
rect -3289 1637 -3255 1649
rect -3289 1581 -3255 1599
rect -3289 1565 -3255 1581
rect -3289 1513 -3255 1527
rect -3289 1493 -3255 1513
rect -3289 1445 -3255 1455
rect -3289 1421 -3255 1445
rect -3289 1377 -3255 1383
rect -3289 1349 -3255 1377
rect -3289 1309 -3255 1311
rect -3289 1277 -3255 1309
rect -3289 1207 -3255 1239
rect -3289 1205 -3255 1207
rect -3289 1139 -3255 1167
rect -3289 1133 -3255 1139
rect -3289 1071 -3255 1095
rect -3289 1061 -3255 1071
rect -3289 1003 -3255 1023
rect -3289 989 -3255 1003
rect -3289 935 -3255 951
rect -3289 917 -3255 935
rect -3289 867 -3255 879
rect -3289 845 -3255 867
rect 3255 2873 3289 2895
rect 3255 2861 3289 2873
rect 3255 2805 3289 2823
rect 3255 2789 3289 2805
rect 3255 2737 3289 2751
rect 3255 2717 3289 2737
rect 3255 2669 3289 2679
rect 3255 2645 3289 2669
rect 3255 2601 3289 2607
rect 3255 2573 3289 2601
rect 3255 2533 3289 2535
rect 3255 2501 3289 2533
rect 3255 2431 3289 2463
rect 3255 2429 3289 2431
rect 3255 2363 3289 2391
rect 3255 2357 3289 2363
rect 3255 2295 3289 2319
rect 3255 2285 3289 2295
rect 3255 2227 3289 2247
rect 3255 2213 3289 2227
rect 3255 2159 3289 2175
rect 3255 2141 3289 2159
rect 3255 2091 3289 2103
rect 3255 2069 3289 2091
rect 3255 2023 3289 2031
rect 3255 1997 3289 2023
rect 3255 1955 3289 1959
rect 3255 1925 3289 1955
rect 3255 1853 3289 1887
rect 3255 1785 3289 1815
rect 3255 1781 3289 1785
rect 3255 1717 3289 1743
rect 3255 1709 3289 1717
rect 3255 1649 3289 1671
rect 3255 1637 3289 1649
rect 3255 1581 3289 1599
rect 3255 1565 3289 1581
rect 3255 1513 3289 1527
rect 3255 1493 3289 1513
rect 3255 1445 3289 1455
rect 3255 1421 3289 1445
rect 3255 1377 3289 1383
rect 3255 1349 3289 1377
rect 3255 1309 3289 1311
rect 3255 1277 3289 1309
rect 3255 1207 3289 1239
rect 3255 1205 3289 1207
rect 3255 1139 3289 1167
rect 3255 1133 3289 1139
rect 3255 1071 3289 1095
rect 3255 1061 3289 1071
rect 3255 1003 3289 1023
rect 3255 989 3289 1003
rect 3255 935 3289 951
rect 3255 917 3289 935
rect 3255 867 3289 879
rect 3255 845 3289 867
rect -3221 651 -3187 685
rect -3149 651 -3145 685
rect -3145 651 -3115 685
rect -3077 651 -3043 685
rect -3005 651 -2975 685
rect -2975 651 -2971 685
rect -2933 651 -2907 685
rect -2907 651 -2899 685
rect -2861 651 -2839 685
rect -2839 651 -2827 685
rect -2789 651 -2771 685
rect -2771 651 -2755 685
rect -2717 651 -2703 685
rect -2703 651 -2683 685
rect -2645 651 -2635 685
rect -2635 651 -2611 685
rect -2573 651 -2567 685
rect -2567 651 -2539 685
rect -2501 651 -2499 685
rect -2499 651 -2467 685
rect -2429 651 -2397 685
rect -2397 651 -2395 685
rect -2357 651 -2329 685
rect -2329 651 -2323 685
rect -2285 651 -2261 685
rect -2261 651 -2251 685
rect -2213 651 -2193 685
rect -2193 651 -2179 685
rect -2141 651 -2125 685
rect -2125 651 -2107 685
rect -2069 651 -2057 685
rect -2057 651 -2035 685
rect -1997 651 -1989 685
rect -1989 651 -1963 685
rect -1925 651 -1921 685
rect -1921 651 -1891 685
rect -1853 651 -1819 685
rect -1781 651 -1751 685
rect -1751 651 -1747 685
rect -1709 651 -1683 685
rect -1683 651 -1675 685
rect -1637 651 -1615 685
rect -1615 651 -1603 685
rect -1565 651 -1547 685
rect -1547 651 -1531 685
rect -1493 651 -1479 685
rect -1479 651 -1459 685
rect -1421 651 -1411 685
rect -1411 651 -1387 685
rect -1349 651 -1343 685
rect -1343 651 -1315 685
rect -1277 651 -1275 685
rect -1275 651 -1243 685
rect -1205 651 -1173 685
rect -1173 651 -1171 685
rect -1133 651 -1105 685
rect -1105 651 -1099 685
rect -1061 651 -1037 685
rect -1037 651 -1027 685
rect -989 651 -969 685
rect -969 651 -955 685
rect -917 651 -901 685
rect -901 651 -883 685
rect -845 651 -833 685
rect -833 651 -811 685
rect -773 651 -765 685
rect -765 651 -739 685
rect -701 651 -697 685
rect -697 651 -667 685
rect -629 651 -595 685
rect -557 651 -527 685
rect -527 651 -523 685
rect -485 651 -459 685
rect -459 651 -451 685
rect -413 651 -391 685
rect -391 651 -379 685
rect -341 651 -323 685
rect -323 651 -307 685
rect -269 651 -255 685
rect -255 651 -235 685
rect -197 651 -187 685
rect -187 651 -163 685
rect -125 651 -119 685
rect -119 651 -91 685
rect -53 651 -51 685
rect -51 651 -19 685
rect 19 651 51 685
rect 51 651 53 685
rect 91 651 119 685
rect 119 651 125 685
rect 163 651 187 685
rect 187 651 197 685
rect 235 651 255 685
rect 255 651 269 685
rect 307 651 323 685
rect 323 651 341 685
rect 379 651 391 685
rect 391 651 413 685
rect 451 651 459 685
rect 459 651 485 685
rect 523 651 527 685
rect 527 651 557 685
rect 595 651 629 685
rect 667 651 697 685
rect 697 651 701 685
rect 739 651 765 685
rect 765 651 773 685
rect 811 651 833 685
rect 833 651 845 685
rect 883 651 901 685
rect 901 651 917 685
rect 955 651 969 685
rect 969 651 989 685
rect 1027 651 1037 685
rect 1037 651 1061 685
rect 1099 651 1105 685
rect 1105 651 1133 685
rect 1171 651 1173 685
rect 1173 651 1205 685
rect 1243 651 1275 685
rect 1275 651 1277 685
rect 1315 651 1343 685
rect 1343 651 1349 685
rect 1387 651 1411 685
rect 1411 651 1421 685
rect 1459 651 1479 685
rect 1479 651 1493 685
rect 1531 651 1547 685
rect 1547 651 1565 685
rect 1603 651 1615 685
rect 1615 651 1637 685
rect 1675 651 1683 685
rect 1683 651 1709 685
rect 1747 651 1751 685
rect 1751 651 1781 685
rect 1819 651 1853 685
rect 1891 651 1921 685
rect 1921 651 1925 685
rect 1963 651 1989 685
rect 1989 651 1997 685
rect 2035 651 2057 685
rect 2057 651 2069 685
rect 2107 651 2125 685
rect 2125 651 2141 685
rect 2179 651 2193 685
rect 2193 651 2213 685
rect 2251 651 2261 685
rect 2261 651 2285 685
rect 2323 651 2329 685
rect 2329 651 2357 685
rect 2395 651 2397 685
rect 2397 651 2429 685
rect 2467 651 2499 685
rect 2499 651 2501 685
rect 2539 651 2567 685
rect 2567 651 2573 685
rect 2611 651 2635 685
rect 2635 651 2645 685
rect 2683 651 2703 685
rect 2703 651 2717 685
rect 2755 651 2771 685
rect 2771 651 2789 685
rect 2827 651 2839 685
rect 2839 651 2861 685
rect 2899 651 2907 685
rect 2907 651 2933 685
rect 2971 651 2975 685
rect 2975 651 3005 685
rect 3043 651 3077 685
rect 3115 651 3145 685
rect 3145 651 3149 685
rect 3187 651 3221 685
rect -3221 315 -3187 349
rect -3149 315 -3145 349
rect -3145 315 -3115 349
rect -3077 315 -3043 349
rect -3005 315 -2975 349
rect -2975 315 -2971 349
rect -2933 315 -2907 349
rect -2907 315 -2899 349
rect -2861 315 -2839 349
rect -2839 315 -2827 349
rect -2789 315 -2771 349
rect -2771 315 -2755 349
rect -2717 315 -2703 349
rect -2703 315 -2683 349
rect -2645 315 -2635 349
rect -2635 315 -2611 349
rect -2573 315 -2567 349
rect -2567 315 -2539 349
rect -2501 315 -2499 349
rect -2499 315 -2467 349
rect -2429 315 -2397 349
rect -2397 315 -2395 349
rect -2357 315 -2329 349
rect -2329 315 -2323 349
rect -2285 315 -2261 349
rect -2261 315 -2251 349
rect -2213 315 -2193 349
rect -2193 315 -2179 349
rect -2141 315 -2125 349
rect -2125 315 -2107 349
rect -2069 315 -2057 349
rect -2057 315 -2035 349
rect -1997 315 -1989 349
rect -1989 315 -1963 349
rect -1925 315 -1921 349
rect -1921 315 -1891 349
rect -1853 315 -1819 349
rect -1781 315 -1751 349
rect -1751 315 -1747 349
rect -1709 315 -1683 349
rect -1683 315 -1675 349
rect -1637 315 -1615 349
rect -1615 315 -1603 349
rect -1565 315 -1547 349
rect -1547 315 -1531 349
rect -1493 315 -1479 349
rect -1479 315 -1459 349
rect -1421 315 -1411 349
rect -1411 315 -1387 349
rect -1349 315 -1343 349
rect -1343 315 -1315 349
rect -1277 315 -1275 349
rect -1275 315 -1243 349
rect -1205 315 -1173 349
rect -1173 315 -1171 349
rect -1133 315 -1105 349
rect -1105 315 -1099 349
rect -1061 315 -1037 349
rect -1037 315 -1027 349
rect -989 315 -969 349
rect -969 315 -955 349
rect -917 315 -901 349
rect -901 315 -883 349
rect -845 315 -833 349
rect -833 315 -811 349
rect -773 315 -765 349
rect -765 315 -739 349
rect -701 315 -697 349
rect -697 315 -667 349
rect -629 315 -595 349
rect -557 315 -527 349
rect -527 315 -523 349
rect -485 315 -459 349
rect -459 315 -451 349
rect -413 315 -391 349
rect -391 315 -379 349
rect -341 315 -323 349
rect -323 315 -307 349
rect -269 315 -255 349
rect -255 315 -235 349
rect -197 315 -187 349
rect -187 315 -163 349
rect -125 315 -119 349
rect -119 315 -91 349
rect -53 315 -51 349
rect -51 315 -19 349
rect 19 315 51 349
rect 51 315 53 349
rect 91 315 119 349
rect 119 315 125 349
rect 163 315 187 349
rect 187 315 197 349
rect 235 315 255 349
rect 255 315 269 349
rect 307 315 323 349
rect 323 315 341 349
rect 379 315 391 349
rect 391 315 413 349
rect 451 315 459 349
rect 459 315 485 349
rect 523 315 527 349
rect 527 315 557 349
rect 595 315 629 349
rect 667 315 697 349
rect 697 315 701 349
rect 739 315 765 349
rect 765 315 773 349
rect 811 315 833 349
rect 833 315 845 349
rect 883 315 901 349
rect 901 315 917 349
rect 955 315 969 349
rect 969 315 989 349
rect 1027 315 1037 349
rect 1037 315 1061 349
rect 1099 315 1105 349
rect 1105 315 1133 349
rect 1171 315 1173 349
rect 1173 315 1205 349
rect 1243 315 1275 349
rect 1275 315 1277 349
rect 1315 315 1343 349
rect 1343 315 1349 349
rect 1387 315 1411 349
rect 1411 315 1421 349
rect 1459 315 1479 349
rect 1479 315 1493 349
rect 1531 315 1547 349
rect 1547 315 1565 349
rect 1603 315 1615 349
rect 1615 315 1637 349
rect 1675 315 1683 349
rect 1683 315 1709 349
rect 1747 315 1751 349
rect 1751 315 1781 349
rect 1819 315 1853 349
rect 1891 315 1921 349
rect 1921 315 1925 349
rect 1963 315 1989 349
rect 1989 315 1997 349
rect 2035 315 2057 349
rect 2057 315 2069 349
rect 2107 315 2125 349
rect 2125 315 2141 349
rect 2179 315 2193 349
rect 2193 315 2213 349
rect 2251 315 2261 349
rect 2261 315 2285 349
rect 2323 315 2329 349
rect 2329 315 2357 349
rect 2395 315 2397 349
rect 2397 315 2429 349
rect 2467 315 2499 349
rect 2499 315 2501 349
rect 2539 315 2567 349
rect 2567 315 2573 349
rect 2611 315 2635 349
rect 2635 315 2645 349
rect 2683 315 2703 349
rect 2703 315 2717 349
rect 2755 315 2771 349
rect 2771 315 2789 349
rect 2827 315 2839 349
rect 2839 315 2861 349
rect 2899 315 2907 349
rect 2907 315 2933 349
rect 2971 315 2975 349
rect 2975 315 3005 349
rect 3043 315 3077 349
rect 3115 315 3145 349
rect 3145 315 3149 349
rect 3187 315 3221 349
rect -3289 45 -3255 67
rect -3289 33 -3255 45
rect -3289 -23 -3255 -5
rect -3289 -39 -3255 -23
rect -3289 -91 -3255 -77
rect -3289 -111 -3255 -91
rect -3289 -159 -3255 -149
rect -3289 -183 -3255 -159
rect -3289 -227 -3255 -221
rect -3289 -255 -3255 -227
rect -3289 -295 -3255 -293
rect -3289 -327 -3255 -295
rect -3289 -397 -3255 -365
rect -3289 -399 -3255 -397
rect -3289 -465 -3255 -437
rect -3289 -471 -3255 -465
rect -3289 -533 -3255 -509
rect -3289 -543 -3255 -533
rect -3289 -601 -3255 -581
rect -3289 -615 -3255 -601
rect -3289 -669 -3255 -653
rect -3289 -687 -3255 -669
rect -3289 -737 -3255 -725
rect -3289 -759 -3255 -737
rect -3289 -805 -3255 -797
rect -3289 -831 -3255 -805
rect -3289 -873 -3255 -869
rect -3289 -903 -3255 -873
rect -3289 -975 -3255 -941
rect -3289 -1043 -3255 -1013
rect -3289 -1047 -3255 -1043
rect -3289 -1111 -3255 -1085
rect -3289 -1119 -3255 -1111
rect -3021 115 -2987 149
rect -2949 115 -2943 149
rect -2943 115 -2915 149
rect -2877 115 -2875 149
rect -2875 115 -2843 149
rect -2805 115 -2773 149
rect -2773 115 -2771 149
rect -2733 115 -2705 149
rect -2705 115 -2699 149
rect -2661 115 -2637 149
rect -2637 115 -2627 149
rect -2589 115 -2569 149
rect -2569 115 -2555 149
rect -2517 115 -2501 149
rect -2501 115 -2483 149
rect -2445 115 -2433 149
rect -2433 115 -2411 149
rect -2373 115 -2365 149
rect -2365 115 -2339 149
rect -2301 115 -2297 149
rect -2297 115 -2267 149
rect -2229 115 -2195 149
rect -2157 115 -2127 149
rect -2127 115 -2123 149
rect -2085 115 -2059 149
rect -2059 115 -2051 149
rect -2013 115 -1991 149
rect -1991 115 -1979 149
rect -1941 115 -1923 149
rect -1923 115 -1907 149
rect -1869 115 -1855 149
rect -1855 115 -1835 149
rect -1797 115 -1787 149
rect -1787 115 -1763 149
rect -1725 115 -1719 149
rect -1719 115 -1691 149
rect -1653 115 -1651 149
rect -1651 115 -1619 149
rect -1581 115 -1549 149
rect -1549 115 -1547 149
rect -1509 115 -1481 149
rect -1481 115 -1475 149
rect -1437 115 -1413 149
rect -1413 115 -1403 149
rect -1365 115 -1345 149
rect -1345 115 -1331 149
rect -1293 115 -1277 149
rect -1277 115 -1259 149
rect -1221 115 -1209 149
rect -1209 115 -1187 149
rect -1149 115 -1141 149
rect -1141 115 -1115 149
rect -1077 115 -1073 149
rect -1073 115 -1043 149
rect -1005 115 -971 149
rect -933 115 -903 149
rect -903 115 -899 149
rect -861 115 -835 149
rect -835 115 -827 149
rect -789 115 -767 149
rect -767 115 -755 149
rect -717 115 -699 149
rect -699 115 -683 149
rect -645 115 -631 149
rect -631 115 -611 149
rect -573 115 -563 149
rect -563 115 -539 149
rect -501 115 -495 149
rect -495 115 -467 149
rect -429 115 -427 149
rect -427 115 -395 149
rect -357 115 -325 149
rect -325 115 -323 149
rect -285 115 -257 149
rect -257 115 -251 149
rect -213 115 -179 149
rect -3089 -1 -3055 25
rect -3089 -9 -3055 -1
rect -3089 -69 -3055 -47
rect -3089 -81 -3055 -69
rect -3089 -137 -3055 -119
rect -3089 -153 -3055 -137
rect -3089 -205 -3055 -191
rect -3089 -225 -3055 -205
rect -3089 -273 -3055 -263
rect -3089 -297 -3055 -273
rect -3089 -341 -3055 -335
rect -3089 -369 -3055 -341
rect -3089 -409 -3055 -407
rect -3089 -441 -3055 -409
rect -3089 -511 -3055 -479
rect -3089 -513 -3055 -511
rect -3089 -579 -3055 -551
rect -3089 -585 -3055 -579
rect -3089 -647 -3055 -623
rect -3089 -657 -3055 -647
rect -3089 -715 -3055 -695
rect -3089 -729 -3055 -715
rect -3089 -783 -3055 -767
rect -3089 -801 -3055 -783
rect -3089 -851 -3055 -839
rect -3089 -873 -3055 -851
rect -3089 -919 -3055 -911
rect -3089 -945 -3055 -919
rect -145 -1 -111 25
rect -145 -9 -111 -1
rect -145 -69 -111 -47
rect -145 -81 -111 -69
rect -145 -137 -111 -119
rect -145 -153 -111 -137
rect -145 -205 -111 -191
rect -145 -225 -111 -205
rect -145 -273 -111 -263
rect -145 -297 -111 -273
rect -145 -341 -111 -335
rect -145 -369 -111 -341
rect -145 -409 -111 -407
rect -145 -441 -111 -409
rect -145 -511 -111 -479
rect -145 -513 -111 -511
rect -145 -579 -111 -551
rect -145 -585 -111 -579
rect -145 -647 -111 -623
rect -145 -657 -111 -647
rect -145 -715 -111 -695
rect -145 -729 -111 -715
rect -145 -783 -111 -767
rect -145 -801 -111 -783
rect -145 -851 -111 -839
rect -145 -873 -111 -851
rect -145 -919 -111 -911
rect -145 -945 -111 -919
rect -3021 -1069 -2987 -1035
rect -2949 -1069 -2943 -1035
rect -2943 -1069 -2915 -1035
rect -2877 -1069 -2875 -1035
rect -2875 -1069 -2843 -1035
rect -2805 -1069 -2773 -1035
rect -2773 -1069 -2771 -1035
rect -2733 -1069 -2705 -1035
rect -2705 -1069 -2699 -1035
rect -2661 -1069 -2637 -1035
rect -2637 -1069 -2627 -1035
rect -2589 -1069 -2569 -1035
rect -2569 -1069 -2555 -1035
rect -2517 -1069 -2501 -1035
rect -2501 -1069 -2483 -1035
rect -2445 -1069 -2433 -1035
rect -2433 -1069 -2411 -1035
rect -2373 -1069 -2365 -1035
rect -2365 -1069 -2339 -1035
rect -2301 -1069 -2297 -1035
rect -2297 -1069 -2267 -1035
rect -2229 -1069 -2195 -1035
rect -2157 -1069 -2127 -1035
rect -2127 -1069 -2123 -1035
rect -2085 -1069 -2059 -1035
rect -2059 -1069 -2051 -1035
rect -2013 -1069 -1991 -1035
rect -1991 -1069 -1979 -1035
rect -1941 -1069 -1923 -1035
rect -1923 -1069 -1907 -1035
rect -1869 -1069 -1855 -1035
rect -1855 -1069 -1835 -1035
rect -1797 -1069 -1787 -1035
rect -1787 -1069 -1763 -1035
rect -1725 -1069 -1719 -1035
rect -1719 -1069 -1691 -1035
rect -1653 -1069 -1651 -1035
rect -1651 -1069 -1619 -1035
rect -1581 -1069 -1549 -1035
rect -1549 -1069 -1547 -1035
rect -1509 -1069 -1481 -1035
rect -1481 -1069 -1475 -1035
rect -1437 -1069 -1413 -1035
rect -1413 -1069 -1403 -1035
rect -1365 -1069 -1345 -1035
rect -1345 -1069 -1331 -1035
rect -1293 -1069 -1277 -1035
rect -1277 -1069 -1259 -1035
rect -1221 -1069 -1209 -1035
rect -1209 -1069 -1187 -1035
rect -1149 -1069 -1141 -1035
rect -1141 -1069 -1115 -1035
rect -1077 -1069 -1073 -1035
rect -1073 -1069 -1043 -1035
rect -1005 -1069 -971 -1035
rect -933 -1069 -903 -1035
rect -903 -1069 -899 -1035
rect -861 -1069 -835 -1035
rect -835 -1069 -827 -1035
rect -789 -1069 -767 -1035
rect -767 -1069 -755 -1035
rect -717 -1069 -699 -1035
rect -699 -1069 -683 -1035
rect -645 -1069 -631 -1035
rect -631 -1069 -611 -1035
rect -573 -1069 -563 -1035
rect -563 -1069 -539 -1035
rect -501 -1069 -495 -1035
rect -495 -1069 -467 -1035
rect -429 -1069 -427 -1035
rect -427 -1069 -395 -1035
rect -357 -1069 -325 -1035
rect -325 -1069 -323 -1035
rect -285 -1069 -257 -1035
rect -257 -1069 -251 -1035
rect -213 -1069 -179 -1035
rect 3255 45 3289 67
rect 3255 33 3289 45
rect 3255 -23 3289 -5
rect 3255 -39 3289 -23
rect 3255 -91 3289 -77
rect 3255 -111 3289 -91
rect 3255 -159 3289 -149
rect 3255 -183 3289 -159
rect 3255 -227 3289 -221
rect 3255 -255 3289 -227
rect 3255 -295 3289 -293
rect 3255 -327 3289 -295
rect 3255 -397 3289 -365
rect 3255 -399 3289 -397
rect 3255 -465 3289 -437
rect 3255 -471 3289 -465
rect 3255 -533 3289 -509
rect 3255 -543 3289 -533
rect 3255 -601 3289 -581
rect 3255 -615 3289 -601
rect 3255 -669 3289 -653
rect 3255 -687 3289 -669
rect 3255 -737 3289 -725
rect 3255 -759 3289 -737
rect 3255 -805 3289 -797
rect 3255 -831 3289 -805
rect 3255 -873 3289 -869
rect 3255 -903 3289 -873
rect 3255 -975 3289 -941
rect 3255 -1043 3289 -1013
rect 3255 -1047 3289 -1043
rect -3289 -1179 -3255 -1157
rect -3289 -1191 -3255 -1179
rect -3289 -1247 -3255 -1229
rect -3289 -1263 -3255 -1247
rect 3255 -1111 3289 -1085
rect 3255 -1119 3289 -1111
rect 3255 -1179 3289 -1157
rect 3255 -1191 3289 -1179
rect -3289 -1315 -3255 -1301
rect -3289 -1335 -3255 -1315
rect -3289 -1383 -3255 -1373
rect -3289 -1407 -3255 -1383
rect -3289 -1451 -3255 -1445
rect -3289 -1479 -3255 -1451
rect -3289 -1519 -3255 -1517
rect -3289 -1551 -3255 -1519
rect -3289 -1621 -3255 -1589
rect -3289 -1623 -3255 -1621
rect -3289 -1689 -3255 -1661
rect -3289 -1695 -3255 -1689
rect -3289 -1757 -3255 -1733
rect -3289 -1767 -3255 -1757
rect -3289 -1825 -3255 -1805
rect -3289 -1839 -3255 -1825
rect -3289 -1893 -3255 -1877
rect -3289 -1911 -3255 -1893
rect -3289 -1961 -3255 -1949
rect -3289 -1983 -3255 -1961
rect -3289 -2029 -3255 -2021
rect -3289 -2055 -3255 -2029
rect -3289 -2097 -3255 -2093
rect -3289 -2127 -3255 -2097
rect -3289 -2199 -3255 -2165
rect -3289 -2267 -3255 -2237
rect -3289 -2271 -3255 -2267
rect -3289 -2335 -3255 -2309
rect -3289 -2343 -3255 -2335
rect -3289 -2403 -3255 -2381
rect -3289 -2415 -3255 -2403
rect -3289 -2471 -3255 -2453
rect -3289 -2487 -3255 -2471
rect -3289 -2539 -3255 -2525
rect -3289 -2559 -3255 -2539
rect -3289 -2607 -3255 -2597
rect -3289 -2631 -3255 -2607
rect -3289 -2675 -3255 -2669
rect -3289 -2703 -3255 -2675
rect -3289 -2743 -3255 -2741
rect -3289 -2775 -3255 -2743
rect -3005 -1285 -2971 -1251
rect -2933 -1285 -2907 -1251
rect -2907 -1285 -2899 -1251
rect -2861 -1285 -2839 -1251
rect -2839 -1285 -2827 -1251
rect -2789 -1285 -2771 -1251
rect -2771 -1285 -2755 -1251
rect -2717 -1285 -2703 -1251
rect -2703 -1285 -2683 -1251
rect -2645 -1285 -2635 -1251
rect -2635 -1285 -2611 -1251
rect -2573 -1285 -2567 -1251
rect -2567 -1285 -2539 -1251
rect -2501 -1285 -2499 -1251
rect -2499 -1285 -2467 -1251
rect -2429 -1285 -2397 -1251
rect -2397 -1285 -2395 -1251
rect -2357 -1285 -2329 -1251
rect -2329 -1285 -2323 -1251
rect -2285 -1285 -2261 -1251
rect -2261 -1285 -2251 -1251
rect -2213 -1285 -2193 -1251
rect -2193 -1285 -2179 -1251
rect -2141 -1285 -2125 -1251
rect -2125 -1285 -2107 -1251
rect -2069 -1285 -2057 -1251
rect -2057 -1285 -2035 -1251
rect -1997 -1285 -1989 -1251
rect -1989 -1285 -1963 -1251
rect -1925 -1285 -1921 -1251
rect -1921 -1285 -1891 -1251
rect -1853 -1285 -1819 -1251
rect -1781 -1285 -1751 -1251
rect -1751 -1285 -1747 -1251
rect -1709 -1285 -1683 -1251
rect -1683 -1285 -1675 -1251
rect -1637 -1285 -1615 -1251
rect -1615 -1285 -1603 -1251
rect -1565 -1285 -1547 -1251
rect -1547 -1285 -1531 -1251
rect -1493 -1285 -1479 -1251
rect -1479 -1285 -1459 -1251
rect -1421 -1285 -1411 -1251
rect -1411 -1285 -1387 -1251
rect -1349 -1285 -1343 -1251
rect -1343 -1285 -1315 -1251
rect -1277 -1285 -1275 -1251
rect -1275 -1285 -1243 -1251
rect -1205 -1285 -1173 -1251
rect -1173 -1285 -1171 -1251
rect -1133 -1285 -1105 -1251
rect -1105 -1285 -1099 -1251
rect -1061 -1285 -1037 -1251
rect -1037 -1285 -1027 -1251
rect -989 -1285 -969 -1251
rect -969 -1285 -955 -1251
rect -917 -1285 -901 -1251
rect -901 -1285 -883 -1251
rect -845 -1285 -833 -1251
rect -833 -1285 -811 -1251
rect -773 -1285 -765 -1251
rect -765 -1285 -739 -1251
rect -701 -1285 -697 -1251
rect -697 -1285 -667 -1251
rect -629 -1285 -595 -1251
rect -557 -1285 -527 -1251
rect -527 -1285 -523 -1251
rect -485 -1285 -459 -1251
rect -459 -1285 -451 -1251
rect -413 -1285 -391 -1251
rect -391 -1285 -379 -1251
rect -341 -1285 -323 -1251
rect -323 -1285 -307 -1251
rect -269 -1285 -255 -1251
rect -255 -1285 -235 -1251
rect -197 -1285 -187 -1251
rect -187 -1285 -163 -1251
rect -125 -1285 -119 -1251
rect -119 -1285 -91 -1251
rect -53 -1285 -51 -1251
rect -51 -1285 -19 -1251
rect 19 -1285 51 -1251
rect 51 -1285 53 -1251
rect 91 -1285 119 -1251
rect 119 -1285 125 -1251
rect 163 -1285 187 -1251
rect 187 -1285 197 -1251
rect 235 -1285 255 -1251
rect 255 -1285 269 -1251
rect 307 -1285 323 -1251
rect 323 -1285 341 -1251
rect 379 -1285 391 -1251
rect 391 -1285 413 -1251
rect 451 -1285 459 -1251
rect 459 -1285 485 -1251
rect 523 -1285 527 -1251
rect 527 -1285 557 -1251
rect 595 -1285 629 -1251
rect 667 -1285 697 -1251
rect 697 -1285 701 -1251
rect 739 -1285 765 -1251
rect 765 -1285 773 -1251
rect 811 -1285 833 -1251
rect 833 -1285 845 -1251
rect 883 -1285 901 -1251
rect 901 -1285 917 -1251
rect 955 -1285 969 -1251
rect 969 -1285 989 -1251
rect 1027 -1285 1037 -1251
rect 1037 -1285 1061 -1251
rect 1099 -1285 1105 -1251
rect 1105 -1285 1133 -1251
rect 1171 -1285 1173 -1251
rect 1173 -1285 1205 -1251
rect 1243 -1285 1275 -1251
rect 1275 -1285 1277 -1251
rect 1315 -1285 1343 -1251
rect 1343 -1285 1349 -1251
rect 1387 -1285 1411 -1251
rect 1411 -1285 1421 -1251
rect 1459 -1285 1479 -1251
rect 1479 -1285 1493 -1251
rect 1531 -1285 1547 -1251
rect 1547 -1285 1565 -1251
rect 1603 -1285 1615 -1251
rect 1615 -1285 1637 -1251
rect 1675 -1285 1683 -1251
rect 1683 -1285 1709 -1251
rect 1747 -1285 1751 -1251
rect 1751 -1285 1781 -1251
rect 1819 -1285 1853 -1251
rect 1891 -1285 1921 -1251
rect 1921 -1285 1925 -1251
rect 1963 -1285 1989 -1251
rect 1989 -1285 1997 -1251
rect 2035 -1285 2057 -1251
rect 2057 -1285 2069 -1251
rect 2107 -1285 2125 -1251
rect 2125 -1285 2141 -1251
rect 2179 -1285 2193 -1251
rect 2193 -1285 2213 -1251
rect 2251 -1285 2261 -1251
rect 2261 -1285 2285 -1251
rect 2323 -1285 2329 -1251
rect 2329 -1285 2357 -1251
rect 2395 -1285 2397 -1251
rect 2397 -1285 2429 -1251
rect 2467 -1285 2499 -1251
rect 2499 -1285 2501 -1251
rect 2539 -1285 2567 -1251
rect 2567 -1285 2573 -1251
rect 2611 -1285 2635 -1251
rect 2635 -1285 2645 -1251
rect 2683 -1285 2703 -1251
rect 2703 -1285 2717 -1251
rect 2755 -1285 2771 -1251
rect 2771 -1285 2789 -1251
rect 2827 -1285 2839 -1251
rect 2839 -1285 2861 -1251
rect 2899 -1285 2907 -1251
rect 2907 -1285 2933 -1251
rect 2971 -1285 3005 -1251
rect -3089 -1419 -3055 -1387
rect -3089 -1421 -3055 -1419
rect -3089 -1487 -3055 -1459
rect -3089 -1493 -3055 -1487
rect -3089 -1555 -3055 -1531
rect -3089 -1565 -3055 -1555
rect -3089 -1623 -3055 -1603
rect -3089 -1637 -3055 -1623
rect -3089 -1691 -3055 -1675
rect -3089 -1709 -3055 -1691
rect -3089 -1759 -3055 -1747
rect -3089 -1781 -3055 -1759
rect -3089 -1827 -3055 -1819
rect -3089 -1853 -3055 -1827
rect -3089 -1895 -3055 -1891
rect -3089 -1925 -3055 -1895
rect -3089 -1997 -3055 -1963
rect -3089 -2065 -3055 -2035
rect -3089 -2069 -3055 -2065
rect -3089 -2133 -3055 -2107
rect -3089 -2141 -3055 -2133
rect -3089 -2201 -3055 -2179
rect -3089 -2213 -3055 -2201
rect -3089 -2269 -3055 -2251
rect -3089 -2285 -3055 -2269
rect -3089 -2337 -3055 -2323
rect -3089 -2357 -3055 -2337
rect -3089 -2405 -3055 -2395
rect -3089 -2429 -3055 -2405
rect -3089 -2473 -3055 -2467
rect -3089 -2501 -3055 -2473
rect -3089 -2541 -3055 -2539
rect -3089 -2573 -3055 -2541
rect 3055 -1419 3089 -1387
rect 3055 -1421 3089 -1419
rect 3055 -1487 3089 -1459
rect 3055 -1493 3089 -1487
rect 3055 -1555 3089 -1531
rect 3055 -1565 3089 -1555
rect 3055 -1623 3089 -1603
rect 3055 -1637 3089 -1623
rect 3055 -1691 3089 -1675
rect 3055 -1709 3089 -1691
rect 3055 -1759 3089 -1747
rect 3055 -1781 3089 -1759
rect 3055 -1827 3089 -1819
rect 3055 -1853 3089 -1827
rect 3055 -1895 3089 -1891
rect 3055 -1925 3089 -1895
rect 3055 -1997 3089 -1963
rect 3055 -2065 3089 -2035
rect 3055 -2069 3089 -2065
rect 3055 -2133 3089 -2107
rect 3055 -2141 3089 -2133
rect 3055 -2201 3089 -2179
rect 3055 -2213 3089 -2201
rect 3055 -2269 3089 -2251
rect 3055 -2285 3089 -2269
rect 3055 -2337 3089 -2323
rect 3055 -2357 3089 -2337
rect 3055 -2405 3089 -2395
rect 3055 -2429 3089 -2405
rect 3055 -2473 3089 -2467
rect 3055 -2501 3089 -2473
rect 3055 -2541 3089 -2539
rect 3055 -2573 3089 -2541
rect -3005 -2709 -2971 -2675
rect -2933 -2709 -2907 -2675
rect -2907 -2709 -2899 -2675
rect -2861 -2709 -2839 -2675
rect -2839 -2709 -2827 -2675
rect -2789 -2709 -2771 -2675
rect -2771 -2709 -2755 -2675
rect -2717 -2709 -2703 -2675
rect -2703 -2709 -2683 -2675
rect -2645 -2709 -2635 -2675
rect -2635 -2709 -2611 -2675
rect -2573 -2709 -2567 -2675
rect -2567 -2709 -2539 -2675
rect -2501 -2709 -2499 -2675
rect -2499 -2709 -2467 -2675
rect -2429 -2709 -2397 -2675
rect -2397 -2709 -2395 -2675
rect -2357 -2709 -2329 -2675
rect -2329 -2709 -2323 -2675
rect -2285 -2709 -2261 -2675
rect -2261 -2709 -2251 -2675
rect -2213 -2709 -2193 -2675
rect -2193 -2709 -2179 -2675
rect -2141 -2709 -2125 -2675
rect -2125 -2709 -2107 -2675
rect -2069 -2709 -2057 -2675
rect -2057 -2709 -2035 -2675
rect -1997 -2709 -1989 -2675
rect -1989 -2709 -1963 -2675
rect -1925 -2709 -1921 -2675
rect -1921 -2709 -1891 -2675
rect -1853 -2709 -1819 -2675
rect -1781 -2709 -1751 -2675
rect -1751 -2709 -1747 -2675
rect -1709 -2709 -1683 -2675
rect -1683 -2709 -1675 -2675
rect -1637 -2709 -1615 -2675
rect -1615 -2709 -1603 -2675
rect -1565 -2709 -1547 -2675
rect -1547 -2709 -1531 -2675
rect -1493 -2709 -1479 -2675
rect -1479 -2709 -1459 -2675
rect -1421 -2709 -1411 -2675
rect -1411 -2709 -1387 -2675
rect -1349 -2709 -1343 -2675
rect -1343 -2709 -1315 -2675
rect -1277 -2709 -1275 -2675
rect -1275 -2709 -1243 -2675
rect -1205 -2709 -1173 -2675
rect -1173 -2709 -1171 -2675
rect -1133 -2709 -1105 -2675
rect -1105 -2709 -1099 -2675
rect -1061 -2709 -1037 -2675
rect -1037 -2709 -1027 -2675
rect -989 -2709 -969 -2675
rect -969 -2709 -955 -2675
rect -917 -2709 -901 -2675
rect -901 -2709 -883 -2675
rect -845 -2709 -833 -2675
rect -833 -2709 -811 -2675
rect -773 -2709 -765 -2675
rect -765 -2709 -739 -2675
rect -701 -2709 -697 -2675
rect -697 -2709 -667 -2675
rect -629 -2709 -595 -2675
rect -557 -2709 -527 -2675
rect -527 -2709 -523 -2675
rect -485 -2709 -459 -2675
rect -459 -2709 -451 -2675
rect -413 -2709 -391 -2675
rect -391 -2709 -379 -2675
rect -341 -2709 -323 -2675
rect -323 -2709 -307 -2675
rect -269 -2709 -255 -2675
rect -255 -2709 -235 -2675
rect -197 -2709 -187 -2675
rect -187 -2709 -163 -2675
rect -125 -2709 -119 -2675
rect -119 -2709 -91 -2675
rect -53 -2709 -51 -2675
rect -51 -2709 -19 -2675
rect 19 -2709 51 -2675
rect 51 -2709 53 -2675
rect 91 -2709 119 -2675
rect 119 -2709 125 -2675
rect 163 -2709 187 -2675
rect 187 -2709 197 -2675
rect 235 -2709 255 -2675
rect 255 -2709 269 -2675
rect 307 -2709 323 -2675
rect 323 -2709 341 -2675
rect 379 -2709 391 -2675
rect 391 -2709 413 -2675
rect 451 -2709 459 -2675
rect 459 -2709 485 -2675
rect 523 -2709 527 -2675
rect 527 -2709 557 -2675
rect 595 -2709 629 -2675
rect 667 -2709 697 -2675
rect 697 -2709 701 -2675
rect 739 -2709 765 -2675
rect 765 -2709 773 -2675
rect 811 -2709 833 -2675
rect 833 -2709 845 -2675
rect 883 -2709 901 -2675
rect 901 -2709 917 -2675
rect 955 -2709 969 -2675
rect 969 -2709 989 -2675
rect 1027 -2709 1037 -2675
rect 1037 -2709 1061 -2675
rect 1099 -2709 1105 -2675
rect 1105 -2709 1133 -2675
rect 1171 -2709 1173 -2675
rect 1173 -2709 1205 -2675
rect 1243 -2709 1275 -2675
rect 1275 -2709 1277 -2675
rect 1315 -2709 1343 -2675
rect 1343 -2709 1349 -2675
rect 1387 -2709 1411 -2675
rect 1411 -2709 1421 -2675
rect 1459 -2709 1479 -2675
rect 1479 -2709 1493 -2675
rect 1531 -2709 1547 -2675
rect 1547 -2709 1565 -2675
rect 1603 -2709 1615 -2675
rect 1615 -2709 1637 -2675
rect 1675 -2709 1683 -2675
rect 1683 -2709 1709 -2675
rect 1747 -2709 1751 -2675
rect 1751 -2709 1781 -2675
rect 1819 -2709 1853 -2675
rect 1891 -2709 1921 -2675
rect 1921 -2709 1925 -2675
rect 1963 -2709 1989 -2675
rect 1989 -2709 1997 -2675
rect 2035 -2709 2057 -2675
rect 2057 -2709 2069 -2675
rect 2107 -2709 2125 -2675
rect 2125 -2709 2141 -2675
rect 2179 -2709 2193 -2675
rect 2193 -2709 2213 -2675
rect 2251 -2709 2261 -2675
rect 2261 -2709 2285 -2675
rect 2323 -2709 2329 -2675
rect 2329 -2709 2357 -2675
rect 2395 -2709 2397 -2675
rect 2397 -2709 2429 -2675
rect 2467 -2709 2499 -2675
rect 2499 -2709 2501 -2675
rect 2539 -2709 2567 -2675
rect 2567 -2709 2573 -2675
rect 2611 -2709 2635 -2675
rect 2635 -2709 2645 -2675
rect 2683 -2709 2703 -2675
rect 2703 -2709 2717 -2675
rect 2755 -2709 2771 -2675
rect 2771 -2709 2789 -2675
rect 2827 -2709 2839 -2675
rect 2839 -2709 2861 -2675
rect 2899 -2709 2907 -2675
rect 2907 -2709 2933 -2675
rect 2971 -2709 3005 -2675
rect 3255 -1247 3289 -1229
rect 3255 -1263 3289 -1247
rect 3255 -1315 3289 -1301
rect 3255 -1335 3289 -1315
rect 3255 -1383 3289 -1373
rect 3255 -1407 3289 -1383
rect 3255 -1451 3289 -1445
rect 3255 -1479 3289 -1451
rect 3255 -1519 3289 -1517
rect 3255 -1551 3289 -1519
rect 3255 -1621 3289 -1589
rect 3255 -1623 3289 -1621
rect 3255 -1689 3289 -1661
rect 3255 -1695 3289 -1689
rect 3255 -1757 3289 -1733
rect 3255 -1767 3289 -1757
rect 3255 -1825 3289 -1805
rect 3255 -1839 3289 -1825
rect 3255 -1893 3289 -1877
rect 3255 -1911 3289 -1893
rect 3255 -1961 3289 -1949
rect 3255 -1983 3289 -1961
rect 3255 -2029 3289 -2021
rect 3255 -2055 3289 -2029
rect 3255 -2097 3289 -2093
rect 3255 -2127 3289 -2097
rect 3255 -2199 3289 -2165
rect 3255 -2267 3289 -2237
rect 3255 -2271 3289 -2267
rect 3255 -2335 3289 -2309
rect 3255 -2343 3289 -2335
rect 3255 -2403 3289 -2381
rect 3255 -2415 3289 -2403
rect 3255 -2471 3289 -2453
rect 3255 -2487 3289 -2471
rect 3255 -2539 3289 -2525
rect 3255 -2559 3289 -2539
rect 3255 -2607 3289 -2597
rect 3255 -2631 3289 -2607
rect 3255 -2675 3289 -2669
rect 3255 -2703 3289 -2675
rect -3289 -2845 -3255 -2813
rect -3289 -2847 -3255 -2845
rect -3289 -2913 -3255 -2885
rect -3289 -2919 -3255 -2913
rect -3289 -2981 -3255 -2957
rect -3289 -2991 -3255 -2981
rect -3289 -3049 -3255 -3029
rect -3289 -3063 -3255 -3049
rect -3289 -3117 -3255 -3101
rect -3289 -3135 -3255 -3117
rect -3289 -3185 -3255 -3173
rect -3289 -3207 -3255 -3185
rect 3255 -2743 3289 -2741
rect 3255 -2775 3289 -2743
rect 3255 -2845 3289 -2813
rect 3255 -2847 3289 -2845
rect 3255 -2913 3289 -2885
rect 3255 -2919 3289 -2913
rect 3255 -2981 3289 -2957
rect 3255 -2991 3289 -2981
rect 3255 -3049 3289 -3029
rect 3255 -3063 3289 -3049
rect 3255 -3117 3289 -3101
rect 3255 -3135 3289 -3117
rect 3255 -3185 3289 -3173
rect 3255 -3207 3289 -3185
rect -3221 -3489 -3187 -3455
rect -3149 -3489 -3145 -3455
rect -3145 -3489 -3115 -3455
rect -3077 -3489 -3043 -3455
rect -3005 -3489 -2975 -3455
rect -2975 -3489 -2971 -3455
rect -2933 -3489 -2907 -3455
rect -2907 -3489 -2899 -3455
rect -2861 -3489 -2839 -3455
rect -2839 -3489 -2827 -3455
rect -2789 -3489 -2771 -3455
rect -2771 -3489 -2755 -3455
rect -2717 -3489 -2703 -3455
rect -2703 -3489 -2683 -3455
rect -2645 -3489 -2635 -3455
rect -2635 -3489 -2611 -3455
rect -2573 -3489 -2567 -3455
rect -2567 -3489 -2539 -3455
rect -2501 -3489 -2499 -3455
rect -2499 -3489 -2467 -3455
rect -2429 -3489 -2397 -3455
rect -2397 -3489 -2395 -3455
rect -2357 -3489 -2329 -3455
rect -2329 -3489 -2323 -3455
rect -2285 -3489 -2261 -3455
rect -2261 -3489 -2251 -3455
rect -2213 -3489 -2193 -3455
rect -2193 -3489 -2179 -3455
rect -2141 -3489 -2125 -3455
rect -2125 -3489 -2107 -3455
rect -2069 -3489 -2057 -3455
rect -2057 -3489 -2035 -3455
rect -1997 -3489 -1989 -3455
rect -1989 -3489 -1963 -3455
rect -1925 -3489 -1921 -3455
rect -1921 -3489 -1891 -3455
rect -1853 -3489 -1819 -3455
rect -1781 -3489 -1751 -3455
rect -1751 -3489 -1747 -3455
rect -1709 -3489 -1683 -3455
rect -1683 -3489 -1675 -3455
rect -1637 -3489 -1615 -3455
rect -1615 -3489 -1603 -3455
rect -1565 -3489 -1547 -3455
rect -1547 -3489 -1531 -3455
rect -1493 -3489 -1479 -3455
rect -1479 -3489 -1459 -3455
rect -1421 -3489 -1411 -3455
rect -1411 -3489 -1387 -3455
rect -1349 -3489 -1343 -3455
rect -1343 -3489 -1315 -3455
rect -1277 -3489 -1275 -3455
rect -1275 -3489 -1243 -3455
rect -1205 -3489 -1173 -3455
rect -1173 -3489 -1171 -3455
rect -1133 -3489 -1105 -3455
rect -1105 -3489 -1099 -3455
rect -1061 -3489 -1037 -3455
rect -1037 -3489 -1027 -3455
rect -989 -3489 -969 -3455
rect -969 -3489 -955 -3455
rect -917 -3489 -901 -3455
rect -901 -3489 -883 -3455
rect -845 -3489 -833 -3455
rect -833 -3489 -811 -3455
rect -773 -3489 -765 -3455
rect -765 -3489 -739 -3455
rect -701 -3489 -697 -3455
rect -697 -3489 -667 -3455
rect -629 -3489 -595 -3455
rect -557 -3489 -527 -3455
rect -527 -3489 -523 -3455
rect -485 -3489 -459 -3455
rect -459 -3489 -451 -3455
rect -413 -3489 -391 -3455
rect -391 -3489 -379 -3455
rect -341 -3489 -323 -3455
rect -323 -3489 -307 -3455
rect -269 -3489 -255 -3455
rect -255 -3489 -235 -3455
rect -197 -3489 -187 -3455
rect -187 -3489 -163 -3455
rect -125 -3489 -119 -3455
rect -119 -3489 -91 -3455
rect -53 -3489 -51 -3455
rect -51 -3489 -19 -3455
rect 19 -3489 51 -3455
rect 51 -3489 53 -3455
rect 91 -3489 119 -3455
rect 119 -3489 125 -3455
rect 163 -3489 187 -3455
rect 187 -3489 197 -3455
rect 235 -3489 255 -3455
rect 255 -3489 269 -3455
rect 307 -3489 323 -3455
rect 323 -3489 341 -3455
rect 379 -3489 391 -3455
rect 391 -3489 413 -3455
rect 451 -3489 459 -3455
rect 459 -3489 485 -3455
rect 523 -3489 527 -3455
rect 527 -3489 557 -3455
rect 595 -3489 629 -3455
rect 667 -3489 697 -3455
rect 697 -3489 701 -3455
rect 739 -3489 765 -3455
rect 765 -3489 773 -3455
rect 811 -3489 833 -3455
rect 833 -3489 845 -3455
rect 883 -3489 901 -3455
rect 901 -3489 917 -3455
rect 955 -3489 969 -3455
rect 969 -3489 989 -3455
rect 1027 -3489 1037 -3455
rect 1037 -3489 1061 -3455
rect 1099 -3489 1105 -3455
rect 1105 -3489 1133 -3455
rect 1171 -3489 1173 -3455
rect 1173 -3489 1205 -3455
rect 1243 -3489 1275 -3455
rect 1275 -3489 1277 -3455
rect 1315 -3489 1343 -3455
rect 1343 -3489 1349 -3455
rect 1387 -3489 1411 -3455
rect 1411 -3489 1421 -3455
rect 1459 -3489 1479 -3455
rect 1479 -3489 1493 -3455
rect 1531 -3489 1547 -3455
rect 1547 -3489 1565 -3455
rect 1603 -3489 1615 -3455
rect 1615 -3489 1637 -3455
rect 1675 -3489 1683 -3455
rect 1683 -3489 1709 -3455
rect 1747 -3489 1751 -3455
rect 1751 -3489 1781 -3455
rect 1819 -3489 1853 -3455
rect 1891 -3489 1921 -3455
rect 1921 -3489 1925 -3455
rect 1963 -3489 1989 -3455
rect 1989 -3489 1997 -3455
rect 2035 -3489 2057 -3455
rect 2057 -3489 2069 -3455
rect 2107 -3489 2125 -3455
rect 2125 -3489 2141 -3455
rect 2179 -3489 2193 -3455
rect 2193 -3489 2213 -3455
rect 2251 -3489 2261 -3455
rect 2261 -3489 2285 -3455
rect 2323 -3489 2329 -3455
rect 2329 -3489 2357 -3455
rect 2395 -3489 2397 -3455
rect 2397 -3489 2429 -3455
rect 2467 -3489 2499 -3455
rect 2499 -3489 2501 -3455
rect 2539 -3489 2567 -3455
rect 2567 -3489 2573 -3455
rect 2611 -3489 2635 -3455
rect 2635 -3489 2645 -3455
rect 2683 -3489 2703 -3455
rect 2703 -3489 2717 -3455
rect 2755 -3489 2771 -3455
rect 2771 -3489 2789 -3455
rect 2827 -3489 2839 -3455
rect 2839 -3489 2861 -3455
rect 2899 -3489 2907 -3455
rect 2907 -3489 2933 -3455
rect 2971 -3489 2975 -3455
rect 2975 -3489 3005 -3455
rect 3043 -3489 3077 -3455
rect 3115 -3489 3145 -3455
rect 3145 -3489 3149 -3455
rect 3187 -3489 3221 -3455
<< metal1 >>
rect -3328 3089 3328 3128
rect -3328 3055 -3221 3089
rect -3187 3055 -3149 3089
rect -3115 3055 -3077 3089
rect -3043 3055 -3005 3089
rect -2971 3055 -2933 3089
rect -2899 3055 -2861 3089
rect -2827 3055 -2789 3089
rect -2755 3055 -2717 3089
rect -2683 3055 -2645 3089
rect -2611 3055 -2573 3089
rect -2539 3055 -2501 3089
rect -2467 3055 -2429 3089
rect -2395 3055 -2357 3089
rect -2323 3055 -2285 3089
rect -2251 3055 -2213 3089
rect -2179 3055 -2141 3089
rect -2107 3055 -2069 3089
rect -2035 3055 -1997 3089
rect -1963 3055 -1925 3089
rect -1891 3055 -1853 3089
rect -1819 3055 -1781 3089
rect -1747 3055 -1709 3089
rect -1675 3055 -1637 3089
rect -1603 3055 -1565 3089
rect -1531 3055 -1493 3089
rect -1459 3055 -1421 3089
rect -1387 3055 -1349 3089
rect -1315 3055 -1277 3089
rect -1243 3055 -1205 3089
rect -1171 3055 -1133 3089
rect -1099 3055 -1061 3089
rect -1027 3055 -989 3089
rect -955 3055 -917 3089
rect -883 3055 -845 3089
rect -811 3055 -773 3089
rect -739 3055 -701 3089
rect -667 3055 -629 3089
rect -595 3055 -557 3089
rect -523 3055 -485 3089
rect -451 3055 -413 3089
rect -379 3055 -341 3089
rect -307 3055 -269 3089
rect -235 3055 -197 3089
rect -163 3055 -125 3089
rect -91 3055 -53 3089
rect -19 3055 19 3089
rect 53 3055 91 3089
rect 125 3055 163 3089
rect 197 3055 235 3089
rect 269 3055 307 3089
rect 341 3055 379 3089
rect 413 3055 451 3089
rect 485 3055 523 3089
rect 557 3055 595 3089
rect 629 3055 667 3089
rect 701 3055 739 3089
rect 773 3055 811 3089
rect 845 3055 883 3089
rect 917 3055 955 3089
rect 989 3055 1027 3089
rect 1061 3055 1099 3089
rect 1133 3055 1171 3089
rect 1205 3055 1243 3089
rect 1277 3055 1315 3089
rect 1349 3055 1387 3089
rect 1421 3055 1459 3089
rect 1493 3055 1531 3089
rect 1565 3055 1603 3089
rect 1637 3055 1675 3089
rect 1709 3055 1747 3089
rect 1781 3055 1819 3089
rect 1853 3055 1891 3089
rect 1925 3055 1963 3089
rect 1997 3055 2035 3089
rect 2069 3055 2107 3089
rect 2141 3055 2179 3089
rect 2213 3055 2251 3089
rect 2285 3055 2323 3089
rect 2357 3055 2395 3089
rect 2429 3055 2467 3089
rect 2501 3055 2539 3089
rect 2573 3055 2611 3089
rect 2645 3055 2683 3089
rect 2717 3055 2755 3089
rect 2789 3055 2827 3089
rect 2861 3055 2899 3089
rect 2933 3055 2971 3089
rect 3005 3055 3043 3089
rect 3077 3055 3115 3089
rect 3149 3055 3187 3089
rect 3221 3055 3328 3089
rect -3328 3016 3328 3055
rect -3328 2988 -2606 3016
rect -3328 2895 -3198 2988
rect -3328 2861 -3289 2895
rect -3255 2861 -3198 2895
rect -3328 2823 -3198 2861
rect -3328 2789 -3289 2823
rect -3255 2789 -3198 2823
rect -3328 2751 -3198 2789
rect -3328 2717 -3289 2751
rect -3255 2744 -3198 2751
rect -2634 2744 -2606 2988
rect -3255 2717 -2606 2744
rect -3328 2716 -2606 2717
rect 2606 2988 3328 3016
rect 2606 2744 2634 2988
rect 3198 2895 3328 2988
rect 3198 2861 3255 2895
rect 3289 2861 3328 2895
rect 3198 2823 3328 2861
rect 3198 2789 3255 2823
rect 3289 2789 3328 2823
rect 3198 2751 3328 2789
rect 3198 2744 3255 2751
rect 2606 2717 3255 2744
rect 3289 2717 3328 2751
rect 2606 2716 3328 2717
rect -3328 2679 -3216 2716
rect -3328 2645 -3289 2679
rect -3255 2645 -3216 2679
rect -3328 2607 -3216 2645
rect -3328 2573 -3289 2607
rect -3255 2573 -3216 2607
rect -3328 2535 -3216 2573
rect 3216 2679 3328 2716
rect 3216 2645 3255 2679
rect 3289 2645 3328 2679
rect 3216 2607 3328 2645
rect 3216 2573 3255 2607
rect 3289 2573 3328 2607
rect -3328 2501 -3289 2535
rect -3255 2501 -3216 2535
rect -3328 2463 -3216 2501
rect -3328 2429 -3289 2463
rect -3255 2429 -3216 2463
rect -2674 2518 2566 2562
rect -2674 2466 -2637 2518
rect -2585 2466 -2573 2518
rect -2521 2466 -2509 2518
rect -2457 2466 -2445 2518
rect -2393 2466 -2381 2518
rect -2329 2466 -2317 2518
rect -2265 2466 -2253 2518
rect -2201 2466 -2189 2518
rect -2137 2466 -2125 2518
rect -2073 2466 -2061 2518
rect -2009 2466 -1997 2518
rect -1945 2466 -1933 2518
rect -1881 2466 -1869 2518
rect -1817 2466 -1805 2518
rect -1753 2466 -1741 2518
rect -1689 2466 -1677 2518
rect -1625 2466 -1613 2518
rect -1561 2466 -1549 2518
rect -1497 2466 -1485 2518
rect -1433 2466 -1421 2518
rect -1369 2466 -1357 2518
rect -1305 2466 -1293 2518
rect -1241 2466 -1229 2518
rect -1177 2466 -1165 2518
rect -1113 2466 -1101 2518
rect -1049 2466 -1037 2518
rect -985 2466 -973 2518
rect -921 2466 -909 2518
rect -857 2466 -845 2518
rect -793 2466 -781 2518
rect -729 2466 -717 2518
rect -665 2466 -653 2518
rect -601 2466 -589 2518
rect -537 2466 -525 2518
rect -473 2466 -461 2518
rect -409 2466 -397 2518
rect -345 2466 -333 2518
rect -281 2466 -269 2518
rect -217 2466 -205 2518
rect -153 2466 -141 2518
rect -89 2466 -77 2518
rect -25 2466 -13 2518
rect 39 2466 51 2518
rect 103 2466 115 2518
rect 167 2466 179 2518
rect 231 2466 243 2518
rect 295 2466 307 2518
rect 359 2466 371 2518
rect 423 2466 435 2518
rect 487 2466 499 2518
rect 551 2466 563 2518
rect 615 2466 627 2518
rect 679 2466 691 2518
rect 743 2466 755 2518
rect 807 2466 819 2518
rect 871 2466 883 2518
rect 935 2466 947 2518
rect 999 2466 1011 2518
rect 1063 2466 1075 2518
rect 1127 2466 1139 2518
rect 1191 2466 1203 2518
rect 1255 2466 1267 2518
rect 1319 2466 1331 2518
rect 1383 2466 1395 2518
rect 1447 2466 1459 2518
rect 1511 2466 1523 2518
rect 1575 2466 1587 2518
rect 1639 2466 1651 2518
rect 1703 2466 1715 2518
rect 1767 2466 1779 2518
rect 1831 2466 1843 2518
rect 1895 2466 1907 2518
rect 1959 2466 1971 2518
rect 2023 2466 2035 2518
rect 2087 2466 2099 2518
rect 2151 2466 2163 2518
rect 2215 2466 2227 2518
rect 2279 2466 2291 2518
rect 2343 2466 2355 2518
rect 2407 2466 2419 2518
rect 2471 2466 2483 2518
rect 2535 2466 2566 2518
rect -2674 2430 2566 2466
rect 3216 2535 3328 2573
rect 3216 2501 3255 2535
rect 3289 2501 3328 2535
rect 3216 2463 3328 2501
rect -3328 2391 -3216 2429
rect -3328 2357 -3289 2391
rect -3255 2357 -3216 2391
rect -3328 2319 -3216 2357
rect -3328 2285 -3289 2319
rect -3255 2285 -3216 2319
rect -3328 2247 -3216 2285
rect -3328 2213 -3289 2247
rect -3255 2213 -3216 2247
rect -3328 2175 -3216 2213
rect -3328 2141 -3289 2175
rect -3255 2141 -3216 2175
rect -2782 2202 -2710 2206
rect -2782 2150 -2772 2202
rect -2720 2150 -2710 2202
rect -2782 2146 -2710 2150
rect -3328 2103 -3216 2141
rect -3328 2069 -3289 2103
rect -3255 2069 -3216 2103
rect -3328 2031 -3216 2069
rect -3328 1997 -3289 2031
rect -3255 1997 -3216 2031
rect -3328 1959 -3216 1997
rect -3328 1925 -3289 1959
rect -3255 1925 -3216 1959
rect -3328 1887 -3216 1925
rect -3328 1853 -3289 1887
rect -3255 1853 -3216 1887
rect -3328 1815 -3216 1853
rect -3328 1781 -3289 1815
rect -3255 1781 -3216 1815
rect -3328 1743 -3216 1781
rect -3328 1709 -3289 1743
rect -3255 1709 -3216 1743
rect -3328 1671 -3216 1709
rect -3328 1637 -3289 1671
rect -3255 1637 -3216 1671
rect -3328 1599 -3216 1637
rect -3328 1565 -3289 1599
rect -3255 1565 -3216 1599
rect -3328 1527 -3216 1565
rect -3328 1493 -3289 1527
rect -3255 1493 -3216 1527
rect -3328 1455 -3216 1493
rect -3328 1421 -3289 1455
rect -3255 1421 -3216 1455
rect -3328 1383 -3216 1421
rect -3328 1349 -3289 1383
rect -3255 1349 -3216 1383
rect -3328 1311 -3216 1349
rect -3328 1277 -3289 1311
rect -3255 1277 -3216 1311
rect -3328 1239 -3216 1277
rect -3328 1205 -3289 1239
rect -3255 1205 -3216 1239
rect -3328 1167 -3216 1205
rect -3328 1133 -3289 1167
rect -3255 1133 -3216 1167
rect -3328 1095 -3216 1133
rect -3328 1061 -3289 1095
rect -3255 1061 -3216 1095
rect -3328 1023 -3216 1061
rect -3328 989 -3289 1023
rect -3255 989 -3216 1023
rect -3328 951 -3216 989
rect -2776 978 -2716 2146
rect -2654 1602 -2594 2430
rect -2528 1602 -2468 1764
rect -2400 1602 -2340 2430
rect -2272 2202 -2200 2206
rect -2272 2150 -2262 2202
rect -2210 2150 -2200 2202
rect -2272 2146 -2200 2150
rect -2266 2056 -2206 2146
rect -2270 1664 -2210 1766
rect -2276 1660 -2204 1664
rect -2276 1608 -2266 1660
rect -2214 1608 -2204 1660
rect -2276 1604 -2204 1608
rect -2654 1542 -2340 1602
rect -2654 1318 -2594 1542
rect -2528 1390 -2468 1542
rect -2400 1284 -2340 1542
rect -2270 1388 -2210 1604
rect -2138 1530 -2078 1890
rect -2008 1530 -1948 1768
rect -2144 1526 -2072 1530
rect -2144 1474 -2134 1526
rect -2082 1474 -2072 1526
rect -2144 1470 -2072 1474
rect -2014 1526 -1942 1530
rect -2014 1474 -2004 1526
rect -1952 1474 -1942 1526
rect -2014 1470 -1942 1474
rect -2008 1392 -1948 1470
rect -1880 1292 -1820 2430
rect -1628 2202 -1556 2206
rect -1628 2150 -1618 2202
rect -1566 2150 -1556 2202
rect -1628 2146 -1556 2150
rect -1502 2202 -1430 2206
rect -1502 2150 -1492 2202
rect -1440 2150 -1430 2202
rect -1502 2146 -1430 2150
rect -1622 1966 -1562 2146
rect -1496 2060 -1436 2146
rect -1750 1530 -1690 1770
rect -1494 1664 -1434 1766
rect -1500 1660 -1428 1664
rect -1500 1608 -1490 1660
rect -1438 1608 -1428 1660
rect -1500 1604 -1428 1608
rect -1756 1526 -1684 1530
rect -1756 1474 -1746 1526
rect -1694 1474 -1684 1526
rect -1756 1470 -1684 1474
rect -1634 1526 -1562 1530
rect -1634 1474 -1624 1526
rect -1572 1474 -1562 1526
rect -1634 1470 -1562 1474
rect -1750 1386 -1690 1470
rect -1628 1280 -1568 1470
rect -1494 1388 -1434 1604
rect -1366 1298 -1306 2430
rect -1238 2202 -1166 2206
rect -1238 2150 -1228 2202
rect -1176 2150 -1166 2202
rect -1238 2146 -1166 2150
rect -1232 2060 -1172 2146
rect -1240 1664 -1180 1766
rect -1246 1660 -1174 1664
rect -1246 1608 -1236 1660
rect -1184 1608 -1174 1660
rect -1246 1604 -1174 1608
rect -1240 1392 -1180 1604
rect -1112 1530 -1052 1872
rect -980 1530 -920 1770
rect -1118 1526 -1046 1530
rect -1118 1474 -1108 1526
rect -1056 1474 -1046 1526
rect -1118 1470 -1046 1474
rect -986 1526 -914 1530
rect -986 1474 -976 1526
rect -924 1474 -914 1526
rect -986 1470 -914 1474
rect -980 1386 -920 1470
rect -846 1284 -786 2430
rect -602 2202 -530 2206
rect -602 2150 -592 2202
rect -540 2150 -530 2202
rect -602 2146 -530 2150
rect -470 2202 -398 2206
rect -470 2150 -460 2202
rect -408 2150 -398 2202
rect -470 2146 -398 2150
rect -596 1940 -536 2146
rect -464 2056 -404 2146
rect -720 1530 -660 1766
rect -464 1664 -404 1766
rect -470 1660 -398 1664
rect -470 1608 -460 1660
rect -408 1608 -398 1660
rect -470 1604 -398 1608
rect -726 1526 -654 1530
rect -726 1474 -716 1526
rect -664 1474 -654 1526
rect -726 1470 -654 1474
rect -602 1526 -530 1530
rect -602 1474 -592 1526
rect -540 1474 -530 1526
rect -602 1470 -530 1474
rect -720 1388 -660 1470
rect -596 1272 -536 1470
rect -464 1388 -404 1604
rect -334 1598 -274 2430
rect -210 1598 -150 1768
rect -76 1598 -16 2430
rect 210 2314 282 2318
rect 210 2262 220 2314
rect 272 2262 282 2314
rect 210 2258 282 2262
rect 594 2314 666 2318
rect 594 2262 604 2314
rect 656 2262 666 2314
rect 594 2258 666 2262
rect -334 1538 -16 1598
rect -334 1276 -274 1538
rect -210 1390 -150 1538
rect -76 1302 -16 1538
rect -2274 978 -2214 1088
rect -2142 978 -2082 1198
rect -3328 917 -3289 951
rect -3255 917 -3216 951
rect -2782 974 -2710 978
rect -2782 922 -2772 974
rect -2720 922 -2710 974
rect -2782 918 -2710 922
rect -2280 974 -2208 978
rect -2280 922 -2270 974
rect -2218 922 -2208 974
rect -2280 918 -2208 922
rect -2148 974 -2076 978
rect -2148 922 -2138 974
rect -2086 922 -2076 974
rect -2148 918 -2076 922
rect -3328 879 -3216 917
rect -3328 845 -3289 879
rect -3255 845 -3216 879
rect -2014 874 -1954 1090
rect -1500 978 -1440 1094
rect -1240 978 -1180 1092
rect -1108 978 -1048 1190
rect -1506 974 -1434 978
rect -1506 922 -1496 974
rect -1444 922 -1434 974
rect -1506 918 -1434 922
rect -1246 974 -1174 978
rect -1246 922 -1236 974
rect -1184 922 -1174 974
rect -1246 918 -1174 922
rect -1114 974 -1042 978
rect -1114 922 -1104 974
rect -1052 922 -1042 974
rect -1114 918 -1042 922
rect -3328 724 -3216 845
rect -2020 870 -1948 874
rect -2020 818 -2010 870
rect -1958 818 -1948 870
rect -2020 814 -1948 818
rect -724 862 -664 1088
rect -464 978 -404 1088
rect -470 974 -398 978
rect -470 922 -460 974
rect -408 922 -398 974
rect -470 918 -398 922
rect 216 874 276 2258
rect 344 1664 404 1858
rect 474 1664 534 1764
rect 600 1664 660 2258
rect 344 1604 660 1664
rect 730 1662 790 1764
rect 724 1658 796 1662
rect 724 1606 734 1658
rect 786 1606 796 1658
rect 724 1602 796 1606
rect 592 1534 664 1538
rect 592 1482 602 1534
rect 654 1482 664 1534
rect 592 1478 664 1482
rect 342 988 402 1192
rect 474 988 534 1088
rect 598 988 658 1478
rect 856 1292 916 2430
rect 982 2202 1054 2206
rect 982 2150 992 2202
rect 1044 2150 1054 2202
rect 982 2146 1054 2150
rect 1238 2202 1310 2206
rect 1238 2150 1248 2202
rect 1300 2150 1310 2202
rect 1238 2146 1310 2150
rect 988 2060 1048 2146
rect 1244 2060 1304 2146
rect 982 1658 1054 1662
rect 982 1606 992 1658
rect 1044 1606 1054 1658
rect 982 1602 1054 1606
rect 988 1386 1048 1602
rect 1116 1538 1176 1854
rect 1240 1658 1312 1662
rect 1240 1606 1250 1658
rect 1302 1606 1312 1658
rect 1240 1602 1312 1606
rect 1110 1534 1182 1538
rect 1110 1482 1120 1534
rect 1172 1482 1182 1534
rect 1110 1478 1182 1482
rect 1246 1386 1306 1602
rect 1374 1310 1434 2430
rect 1626 2314 1698 2318
rect 1626 2262 1636 2314
rect 1688 2262 1698 2314
rect 1626 2258 1698 2262
rect 1500 1662 1560 1764
rect 1632 1662 1692 2258
rect 1996 2202 2068 2206
rect 1996 2150 2006 2202
rect 2058 2150 2068 2202
rect 1996 2146 2068 2150
rect 1762 1662 1822 1764
rect 1892 1662 1952 1872
rect 1494 1658 1566 1662
rect 1494 1606 1504 1658
rect 1556 1606 1566 1658
rect 1494 1602 1566 1606
rect 1632 1602 1952 1662
rect 1624 1534 1950 1538
rect 1624 1482 1634 1534
rect 1686 1482 1950 1534
rect 1624 1478 1950 1482
rect 1630 1300 1690 1478
rect 1762 1390 1822 1478
rect 1890 1288 1950 1478
rect 342 928 658 988
rect 728 986 788 1088
rect 722 982 794 986
rect 722 930 732 982
rect 784 930 794 982
rect 722 926 794 930
rect 1114 874 1174 1186
rect 1502 986 1562 1088
rect 2002 986 2062 2146
rect 2304 1888 2364 2430
rect 3216 2429 3255 2463
rect 3289 2429 3328 2463
rect 3216 2391 3328 2429
rect 3216 2357 3255 2391
rect 3289 2357 3328 2391
rect 3216 2319 3328 2357
rect 3216 2285 3255 2319
rect 3289 2285 3328 2319
rect 3216 2247 3328 2285
rect 3216 2213 3255 2247
rect 3289 2213 3328 2247
rect 3216 2175 3328 2213
rect 2426 2150 2498 2154
rect 2426 2098 2436 2150
rect 2488 2098 2498 2150
rect 2426 2094 2498 2098
rect 3216 2141 3255 2175
rect 3289 2141 3328 2175
rect 3216 2103 3328 2141
rect 2432 1982 2492 2094
rect 3216 2069 3255 2103
rect 3289 2069 3328 2103
rect 3216 2031 3328 2069
rect 3216 1997 3255 2031
rect 3289 1997 3328 2031
rect 3216 1959 3328 1997
rect 3216 1925 3255 1959
rect 3289 1925 3328 1959
rect 3216 1887 3328 1925
rect 3216 1853 3255 1887
rect 3289 1853 3328 1887
rect 3216 1815 3328 1853
rect 3216 1781 3255 1815
rect 3289 1781 3328 1815
rect 3216 1743 3328 1781
rect 3216 1709 3255 1743
rect 3289 1709 3328 1743
rect 3216 1671 3328 1709
rect 3216 1637 3255 1671
rect 3289 1637 3328 1671
rect 3216 1599 3328 1637
rect 3216 1565 3255 1599
rect 3289 1565 3328 1599
rect 3216 1527 3328 1565
rect 3216 1493 3255 1527
rect 3289 1493 3328 1527
rect 3216 1455 3328 1493
rect 3216 1421 3255 1455
rect 3289 1421 3328 1455
rect 3216 1383 3328 1421
rect 3216 1349 3255 1383
rect 3289 1349 3328 1383
rect 3216 1311 3328 1349
rect 3216 1277 3255 1311
rect 3289 1277 3328 1311
rect 3216 1239 3328 1277
rect 3216 1205 3255 1239
rect 3289 1205 3328 1239
rect 1496 982 1568 986
rect 1496 930 1506 982
rect 1558 930 1568 982
rect 1496 926 1568 930
rect 1996 982 2068 986
rect 1996 930 2006 982
rect 2058 930 2068 982
rect 1996 926 2068 930
rect 2432 980 2492 1092
rect 2432 928 2436 980
rect 2488 928 2492 980
rect 2556 976 2616 1196
rect 3216 1167 3328 1205
rect 3216 1133 3255 1167
rect 3289 1133 3328 1167
rect 3216 1095 3328 1133
rect 3216 1061 3255 1095
rect 3289 1061 3328 1095
rect 3216 1023 3328 1061
rect 3216 989 3255 1023
rect 3289 989 3328 1023
rect 2432 918 2492 928
rect 2550 972 2622 976
rect 2550 920 2560 972
rect 2612 920 2622 972
rect 2550 916 2622 920
rect 3216 951 3328 989
rect 3216 917 3255 951
rect 3289 917 3328 951
rect 3216 879 3328 917
rect -724 810 -720 862
rect -668 810 -664 862
rect 210 870 282 874
rect 210 818 220 870
rect 272 818 282 870
rect 210 814 282 818
rect 1108 870 1180 874
rect 1108 818 1118 870
rect 1170 818 1180 870
rect 1108 814 1180 818
rect 3216 845 3255 879
rect 3289 845 3328 879
rect -724 800 -664 810
rect 3216 724 3328 845
rect -3328 685 3328 724
rect -3328 651 -3221 685
rect -3187 651 -3149 685
rect -3115 651 -3077 685
rect -3043 651 -3005 685
rect -2971 651 -2933 685
rect -2899 651 -2861 685
rect -2827 651 -2789 685
rect -2755 651 -2717 685
rect -2683 651 -2645 685
rect -2611 651 -2573 685
rect -2539 651 -2501 685
rect -2467 651 -2429 685
rect -2395 651 -2357 685
rect -2323 651 -2285 685
rect -2251 651 -2213 685
rect -2179 651 -2141 685
rect -2107 651 -2069 685
rect -2035 651 -1997 685
rect -1963 651 -1925 685
rect -1891 651 -1853 685
rect -1819 651 -1781 685
rect -1747 651 -1709 685
rect -1675 651 -1637 685
rect -1603 651 -1565 685
rect -1531 651 -1493 685
rect -1459 651 -1421 685
rect -1387 651 -1349 685
rect -1315 651 -1277 685
rect -1243 651 -1205 685
rect -1171 651 -1133 685
rect -1099 651 -1061 685
rect -1027 651 -989 685
rect -955 651 -917 685
rect -883 651 -845 685
rect -811 651 -773 685
rect -739 651 -701 685
rect -667 651 -629 685
rect -595 651 -557 685
rect -523 651 -485 685
rect -451 651 -413 685
rect -379 651 -341 685
rect -307 651 -269 685
rect -235 651 -197 685
rect -163 651 -125 685
rect -91 651 -53 685
rect -19 651 19 685
rect 53 651 91 685
rect 125 651 163 685
rect 197 651 235 685
rect 269 651 307 685
rect 341 651 379 685
rect 413 651 451 685
rect 485 651 523 685
rect 557 651 595 685
rect 629 651 667 685
rect 701 651 739 685
rect 773 651 811 685
rect 845 651 883 685
rect 917 651 955 685
rect 989 651 1027 685
rect 1061 651 1099 685
rect 1133 651 1171 685
rect 1205 651 1243 685
rect 1277 651 1315 685
rect 1349 651 1387 685
rect 1421 651 1459 685
rect 1493 651 1531 685
rect 1565 651 1603 685
rect 1637 651 1675 685
rect 1709 651 1747 685
rect 1781 651 1819 685
rect 1853 651 1891 685
rect 1925 651 1963 685
rect 1997 651 2035 685
rect 2069 651 2107 685
rect 2141 651 2179 685
rect 2213 651 2251 685
rect 2285 651 2323 685
rect 2357 651 2395 685
rect 2429 651 2467 685
rect 2501 651 2539 685
rect 2573 651 2611 685
rect 2645 651 2683 685
rect 2717 651 2755 685
rect 2789 651 2827 685
rect 2861 651 2899 685
rect 2933 651 2971 685
rect 3005 651 3043 685
rect 3077 651 3115 685
rect 3149 651 3187 685
rect 3221 651 3328 685
rect -3328 612 3328 651
rect -3328 349 3328 388
rect -3328 315 -3221 349
rect -3187 315 -3149 349
rect -3115 315 -3077 349
rect -3043 315 -3005 349
rect -2971 315 -2933 349
rect -2899 315 -2861 349
rect -2827 315 -2789 349
rect -2755 315 -2717 349
rect -2683 315 -2645 349
rect -2611 315 -2573 349
rect -2539 315 -2501 349
rect -2467 315 -2429 349
rect -2395 315 -2357 349
rect -2323 315 -2285 349
rect -2251 315 -2213 349
rect -2179 315 -2141 349
rect -2107 315 -2069 349
rect -2035 315 -1997 349
rect -1963 315 -1925 349
rect -1891 315 -1853 349
rect -1819 315 -1781 349
rect -1747 315 -1709 349
rect -1675 315 -1637 349
rect -1603 315 -1565 349
rect -1531 315 -1493 349
rect -1459 315 -1421 349
rect -1387 315 -1349 349
rect -1315 315 -1277 349
rect -1243 315 -1205 349
rect -1171 315 -1133 349
rect -1099 315 -1061 349
rect -1027 315 -989 349
rect -955 315 -917 349
rect -883 315 -845 349
rect -811 315 -773 349
rect -739 315 -701 349
rect -667 315 -629 349
rect -595 315 -557 349
rect -523 315 -485 349
rect -451 315 -413 349
rect -379 315 -341 349
rect -307 315 -269 349
rect -235 315 -197 349
rect -163 315 -125 349
rect -91 315 -53 349
rect -19 315 19 349
rect 53 315 91 349
rect 125 315 163 349
rect 197 315 235 349
rect 269 315 307 349
rect 341 315 379 349
rect 413 315 451 349
rect 485 315 523 349
rect 557 315 595 349
rect 629 315 667 349
rect 701 315 739 349
rect 773 315 811 349
rect 845 315 883 349
rect 917 315 955 349
rect 989 315 1027 349
rect 1061 315 1099 349
rect 1133 315 1171 349
rect 1205 315 1243 349
rect 1277 315 1315 349
rect 1349 315 1387 349
rect 1421 315 1459 349
rect 1493 315 1531 349
rect 1565 315 1603 349
rect 1637 315 1675 349
rect 1709 315 1747 349
rect 1781 315 1819 349
rect 1853 315 1891 349
rect 1925 315 1963 349
rect 1997 315 2035 349
rect 2069 315 2107 349
rect 2141 315 2179 349
rect 2213 315 2251 349
rect 2285 315 2323 349
rect 2357 315 2395 349
rect 2429 315 2467 349
rect 2501 315 2539 349
rect 2573 315 2611 349
rect 2645 315 2683 349
rect 2717 315 2755 349
rect 2789 315 2827 349
rect 2861 315 2899 349
rect 2933 315 2971 349
rect 3005 315 3043 349
rect 3077 315 3115 349
rect 3149 315 3187 349
rect 3221 315 3328 349
rect -3328 276 3328 315
rect -3328 67 -3216 276
rect -3328 33 -3289 67
rect -3255 33 -3216 67
rect -3328 -5 -3216 33
rect -3328 -39 -3289 -5
rect -3255 -39 -3216 -5
rect -3328 -77 -3216 -39
rect -3328 -111 -3289 -77
rect -3255 -111 -3216 -77
rect -3328 -149 -3216 -111
rect -3328 -183 -3289 -149
rect -3255 -183 -3216 -149
rect -3328 -221 -3216 -183
rect -3328 -255 -3289 -221
rect -3255 -255 -3216 -221
rect -3328 -293 -3216 -255
rect -3328 -327 -3289 -293
rect -3255 -327 -3216 -293
rect -3328 -365 -3216 -327
rect -3328 -399 -3289 -365
rect -3255 -399 -3216 -365
rect -3328 -437 -3216 -399
rect -3328 -471 -3289 -437
rect -3255 -471 -3216 -437
rect -3328 -509 -3216 -471
rect -3328 -543 -3289 -509
rect -3255 -543 -3216 -509
rect -3328 -581 -3216 -543
rect -3328 -615 -3289 -581
rect -3255 -615 -3216 -581
rect -3328 -653 -3216 -615
rect -3328 -687 -3289 -653
rect -3255 -687 -3216 -653
rect -3328 -725 -3216 -687
rect -3328 -759 -3289 -725
rect -3255 -759 -3216 -725
rect -3328 -797 -3216 -759
rect -3328 -831 -3289 -797
rect -3255 -831 -3216 -797
rect -3328 -869 -3216 -831
rect -3328 -903 -3289 -869
rect -3255 -903 -3216 -869
rect -3328 -941 -3216 -903
rect -3328 -975 -3289 -941
rect -3255 -975 -3216 -941
rect -3328 -1013 -3216 -975
rect -3328 -1047 -3289 -1013
rect -3255 -1047 -3216 -1013
rect -3328 -1085 -3216 -1047
rect -3328 -1119 -3289 -1085
rect -3255 -1119 -3216 -1085
rect -3128 149 -72 188
rect -3128 115 -3021 149
rect -2987 115 -2949 149
rect -2915 115 -2877 149
rect -2843 115 -2805 149
rect -2771 115 -2733 149
rect -2699 115 -2661 149
rect -2627 115 -2589 149
rect -2555 115 -2517 149
rect -2483 115 -2445 149
rect -2411 115 -2373 149
rect -2339 115 -2301 149
rect -2267 115 -2229 149
rect -2195 115 -2157 149
rect -2123 115 -2085 149
rect -2051 115 -2013 149
rect -1979 115 -1941 149
rect -1907 115 -1869 149
rect -1835 115 -1797 149
rect -1763 115 -1725 149
rect -1691 115 -1653 149
rect -1619 115 -1581 149
rect -1547 115 -1509 149
rect -1475 115 -1437 149
rect -1403 115 -1365 149
rect -1331 115 -1293 149
rect -1259 115 -1221 149
rect -1187 115 -1149 149
rect -1115 115 -1077 149
rect -1043 115 -1005 149
rect -971 115 -933 149
rect -899 115 -861 149
rect -827 115 -789 149
rect -755 115 -717 149
rect -683 115 -645 149
rect -611 115 -573 149
rect -539 115 -501 149
rect -467 115 -429 149
rect -395 115 -357 149
rect -323 115 -285 149
rect -251 115 -213 149
rect -179 115 -72 149
rect -3128 76 -72 115
rect -3128 25 -3016 76
rect -3128 -9 -3089 25
rect -3055 -9 -3016 25
rect -184 25 -72 76
rect -3128 -47 -3016 -9
rect -2112 10 -2040 14
rect -2112 -42 -2102 10
rect -2050 -42 -2040 10
rect -2112 -46 -2040 -42
rect -1078 10 -1006 14
rect -1078 -42 -1068 10
rect -1016 -42 -1006 10
rect -1078 -46 -1006 -42
rect -184 -9 -145 25
rect -111 -9 -72 25
rect -3128 -81 -3089 -47
rect -3055 -81 -3016 -47
rect -3128 -119 -3016 -81
rect -3128 -153 -3089 -119
rect -3055 -153 -3016 -119
rect -3128 -191 -3016 -153
rect -2628 -106 -2556 -102
rect -2628 -158 -2618 -106
rect -2566 -158 -2556 -106
rect -2628 -162 -2556 -158
rect -3128 -225 -3089 -191
rect -3055 -225 -3016 -191
rect -2622 -220 -2562 -162
rect -3128 -263 -3016 -225
rect -3128 -297 -3089 -263
rect -3055 -297 -3016 -263
rect -3128 -335 -3016 -297
rect -3128 -369 -3089 -335
rect -3055 -369 -3016 -335
rect -3128 -407 -3016 -369
rect -3128 -441 -3089 -407
rect -3055 -441 -3016 -407
rect -3128 -479 -3016 -441
rect -2876 -280 -2562 -220
rect -2496 -224 -2424 -220
rect -2496 -276 -2486 -224
rect -2434 -276 -2424 -224
rect -2496 -280 -2424 -276
rect -2876 -462 -2816 -280
rect -2750 -382 -2690 -280
rect -3128 -513 -3089 -479
rect -3055 -513 -3016 -479
rect -2622 -486 -2562 -280
rect -2490 -386 -2430 -280
rect -2106 -474 -2046 -46
rect -1592 -106 -1520 -102
rect -1592 -158 -1582 -106
rect -1530 -158 -1520 -106
rect -1592 -162 -1520 -158
rect -1720 -224 -1648 -220
rect -1720 -276 -1710 -224
rect -1658 -276 -1648 -224
rect -1720 -280 -1648 -276
rect -1714 -382 -1654 -280
rect -1586 -474 -1526 -162
rect -1466 -224 -1394 -220
rect -1466 -276 -1456 -224
rect -1404 -276 -1394 -224
rect -1466 -280 -1394 -276
rect -1460 -386 -1400 -280
rect -1072 -472 -1012 -46
rect -184 -47 -72 -9
rect -184 -81 -145 -47
rect -111 -81 -72 -47
rect 3216 67 3328 276
rect 3216 33 3255 67
rect 3289 33 3328 67
rect 3216 -5 3328 33
rect 3216 -39 3255 -5
rect 3289 -39 3328 -5
rect -562 -106 -490 -102
rect -562 -158 -552 -106
rect -500 -158 -490 -106
rect -562 -162 -490 -158
rect -184 -119 -72 -81
rect -184 -153 -145 -119
rect -111 -153 -72 -119
rect -556 -220 -496 -162
rect -184 -191 -72 -153
rect 1114 -70 1174 -60
rect 1114 -122 1118 -70
rect 1170 -122 1174 -70
rect 1114 -182 1174 -122
rect 2426 -68 2498 -64
rect 2426 -120 2436 -68
rect 2488 -120 2498 -68
rect 2426 -124 2498 -120
rect 2556 -76 2616 -66
rect -686 -224 -614 -220
rect -686 -276 -676 -224
rect -624 -276 -614 -224
rect -686 -280 -614 -276
rect -556 -280 -236 -220
rect -680 -386 -620 -280
rect -556 -480 -496 -280
rect -426 -382 -366 -280
rect -296 -480 -236 -280
rect -184 -225 -145 -191
rect -111 -225 -72 -191
rect -184 -263 -72 -225
rect -184 -297 -145 -263
rect -111 -297 -72 -263
rect -184 -335 -72 -297
rect -184 -369 -145 -335
rect -111 -369 -72 -335
rect 726 -242 1560 -182
rect 726 -346 786 -242
rect 988 -344 1048 -242
rect -184 -407 -72 -369
rect -184 -441 -145 -407
rect -111 -441 -72 -407
rect -184 -479 -72 -441
rect -3128 -551 -3016 -513
rect -3128 -585 -3089 -551
rect -3055 -585 -3016 -551
rect -184 -513 -145 -479
rect -111 -513 -72 -479
rect -184 -551 -72 -513
rect -3128 -623 -3016 -585
rect -3128 -657 -3089 -623
rect -3055 -657 -3016 -623
rect -3128 -695 -3016 -657
rect -3128 -729 -3089 -695
rect -3055 -729 -3016 -695
rect -3128 -767 -3016 -729
rect -3128 -801 -3089 -767
rect -3055 -801 -3016 -767
rect -3128 -839 -3016 -801
rect -3128 -873 -3089 -839
rect -3055 -873 -3016 -839
rect -3128 -911 -3016 -873
rect -2362 -874 -2302 -580
rect -2230 -756 -2170 -658
rect -1974 -756 -1914 -660
rect -2236 -760 -2164 -756
rect -2236 -812 -2226 -760
rect -2174 -812 -2164 -760
rect -2236 -816 -2164 -812
rect -1980 -760 -1908 -756
rect -1980 -812 -1970 -760
rect -1918 -812 -1908 -760
rect -1980 -816 -1908 -812
rect -1846 -874 -1786 -570
rect -1326 -874 -1266 -580
rect -1200 -756 -1140 -656
rect -942 -756 -882 -656
rect -1206 -760 -1134 -756
rect -1206 -812 -1196 -760
rect -1144 -812 -1134 -760
rect -1206 -816 -1134 -812
rect -948 -760 -876 -756
rect -948 -812 -938 -760
rect -886 -812 -876 -760
rect -948 -816 -876 -812
rect -814 -874 -754 -576
rect -184 -585 -145 -551
rect -111 -585 -72 -551
rect -184 -623 -72 -585
rect -184 -657 -145 -623
rect -111 -657 -72 -623
rect -184 -695 -72 -657
rect -184 -729 -145 -695
rect -111 -729 -72 -695
rect -184 -767 -72 -729
rect 344 -702 404 -542
rect 470 -702 530 -620
rect 596 -702 656 -524
rect 344 -706 662 -702
rect 344 -758 600 -706
rect 652 -758 662 -706
rect 344 -762 662 -758
rect -184 -801 -145 -767
rect -111 -801 -72 -767
rect -184 -839 -72 -801
rect -184 -873 -145 -839
rect -111 -873 -72 -839
rect -3128 -945 -3089 -911
rect -3055 -945 -3016 -911
rect -2368 -878 -2296 -874
rect -2368 -930 -2358 -878
rect -2306 -930 -2296 -878
rect -2368 -934 -2296 -930
rect -1852 -878 -1780 -874
rect -1852 -930 -1842 -878
rect -1790 -930 -1780 -878
rect -1852 -934 -1780 -930
rect -1332 -878 -1260 -874
rect -1332 -930 -1322 -878
rect -1270 -930 -1260 -878
rect -1332 -934 -1260 -930
rect -820 -878 -748 -874
rect -820 -930 -810 -878
rect -758 -930 -748 -878
rect -820 -934 -748 -930
rect -184 -911 -72 -873
rect -3128 -996 -3016 -945
rect -184 -945 -145 -911
rect -111 -945 -72 -911
rect -184 -996 -72 -945
rect -3128 -1035 -72 -996
rect -3128 -1069 -3021 -1035
rect -2987 -1069 -2949 -1035
rect -2915 -1069 -2877 -1035
rect -2843 -1069 -2805 -1035
rect -2771 -1069 -2733 -1035
rect -2699 -1069 -2661 -1035
rect -2627 -1069 -2589 -1035
rect -2555 -1069 -2517 -1035
rect -2483 -1069 -2445 -1035
rect -2411 -1069 -2373 -1035
rect -2339 -1069 -2301 -1035
rect -2267 -1069 -2229 -1035
rect -2195 -1069 -2157 -1035
rect -2123 -1069 -2085 -1035
rect -2051 -1069 -2013 -1035
rect -1979 -1069 -1941 -1035
rect -1907 -1069 -1869 -1035
rect -1835 -1069 -1797 -1035
rect -1763 -1069 -1725 -1035
rect -1691 -1069 -1653 -1035
rect -1619 -1069 -1581 -1035
rect -1547 -1069 -1509 -1035
rect -1475 -1069 -1437 -1035
rect -1403 -1069 -1365 -1035
rect -1331 -1069 -1293 -1035
rect -1259 -1069 -1221 -1035
rect -1187 -1069 -1149 -1035
rect -1115 -1069 -1077 -1035
rect -1043 -1069 -1005 -1035
rect -971 -1069 -933 -1035
rect -899 -1069 -861 -1035
rect -827 -1069 -789 -1035
rect -755 -1069 -717 -1035
rect -683 -1069 -645 -1035
rect -611 -1069 -573 -1035
rect -539 -1069 -501 -1035
rect -467 -1069 -429 -1035
rect -395 -1069 -357 -1035
rect -323 -1069 -285 -1035
rect -251 -1069 -213 -1035
rect -179 -1069 -72 -1035
rect -3128 -1108 -72 -1069
rect 854 -850 914 -526
rect 1114 -558 1174 -242
rect 1242 -346 1302 -242
rect 1500 -346 1560 -242
rect 2432 -322 2492 -124
rect 2556 -128 2560 -76
rect 2612 -128 2616 -76
rect 2556 -422 2616 -128
rect 3216 -77 3328 -39
rect 3216 -111 3255 -77
rect 3289 -111 3328 -77
rect 3216 -149 3328 -111
rect 3216 -183 3255 -149
rect 3289 -183 3328 -149
rect 3216 -221 3328 -183
rect 3216 -255 3255 -221
rect 3289 -255 3328 -221
rect 3216 -293 3328 -255
rect 3216 -327 3255 -293
rect 3289 -327 3328 -293
rect 3216 -365 3328 -327
rect 3216 -399 3255 -365
rect 3289 -399 3328 -365
rect 3216 -437 3328 -399
rect 3216 -471 3255 -437
rect 3289 -471 3328 -437
rect 3216 -509 3328 -471
rect 1370 -850 1430 -526
rect 1630 -702 1690 -530
rect 3216 -543 3255 -509
rect 3289 -543 3328 -509
rect 1760 -702 1820 -622
rect 1888 -702 1948 -546
rect 3216 -581 3328 -543
rect 3216 -615 3255 -581
rect 3289 -615 3328 -581
rect 3216 -653 3328 -615
rect 3216 -687 3255 -653
rect 3289 -687 3328 -653
rect 1624 -706 1948 -702
rect 1624 -758 1634 -706
rect 1686 -758 1948 -706
rect 1624 -762 1948 -758
rect 2296 -850 2356 -690
rect 3216 -725 3328 -687
rect 3216 -759 3255 -725
rect 3289 -759 3328 -725
rect 854 -910 2356 -850
rect 2432 -888 2492 -796
rect 3216 -797 3328 -759
rect 3216 -831 3255 -797
rect 3289 -831 3328 -797
rect 3216 -869 3328 -831
rect -3328 -1157 -3216 -1119
rect -3328 -1191 -3289 -1157
rect -3255 -1191 -3216 -1157
rect -3328 -1229 -3216 -1191
rect 854 -1212 914 -910
rect 2296 -1212 2356 -910
rect 2426 -892 2498 -888
rect 2426 -944 2436 -892
rect 2488 -944 2498 -892
rect 2426 -948 2498 -944
rect 3216 -903 3255 -869
rect 3289 -903 3328 -869
rect 3216 -941 3328 -903
rect 3216 -975 3255 -941
rect 3289 -975 3328 -941
rect 3216 -1013 3328 -975
rect 3216 -1047 3255 -1013
rect 3289 -1047 3328 -1013
rect 3216 -1085 3328 -1047
rect 3216 -1119 3255 -1085
rect 3289 -1119 3328 -1085
rect 3216 -1157 3328 -1119
rect 3216 -1191 3255 -1157
rect 3289 -1191 3328 -1157
rect -3328 -1263 -3289 -1229
rect -3255 -1263 -3216 -1229
rect -3328 -1301 -3216 -1263
rect -3328 -1335 -3289 -1301
rect -3255 -1335 -3216 -1301
rect -3328 -1373 -3216 -1335
rect -3328 -1407 -3289 -1373
rect -3255 -1407 -3216 -1373
rect -3328 -1445 -3216 -1407
rect -3328 -1479 -3289 -1445
rect -3255 -1479 -3216 -1445
rect -3328 -1517 -3216 -1479
rect -3328 -1551 -3289 -1517
rect -3255 -1551 -3216 -1517
rect -3328 -1589 -3216 -1551
rect -3328 -1623 -3289 -1589
rect -3255 -1623 -3216 -1589
rect -3328 -1661 -3216 -1623
rect -3328 -1695 -3289 -1661
rect -3255 -1695 -3216 -1661
rect -3328 -1733 -3216 -1695
rect -3328 -1767 -3289 -1733
rect -3255 -1767 -3216 -1733
rect -3328 -1805 -3216 -1767
rect -3328 -1839 -3289 -1805
rect -3255 -1839 -3216 -1805
rect -3328 -1877 -3216 -1839
rect -3328 -1911 -3289 -1877
rect -3255 -1911 -3216 -1877
rect -3328 -1949 -3216 -1911
rect -3328 -1983 -3289 -1949
rect -3255 -1983 -3216 -1949
rect -3328 -2021 -3216 -1983
rect -3328 -2055 -3289 -2021
rect -3255 -2055 -3216 -2021
rect -3328 -2093 -3216 -2055
rect -3328 -2127 -3289 -2093
rect -3255 -2127 -3216 -2093
rect -3328 -2165 -3216 -2127
rect -3328 -2199 -3289 -2165
rect -3255 -2199 -3216 -2165
rect -3328 -2237 -3216 -2199
rect -3328 -2271 -3289 -2237
rect -3255 -2271 -3216 -2237
rect -3328 -2309 -3216 -2271
rect -3328 -2343 -3289 -2309
rect -3255 -2343 -3216 -2309
rect -3328 -2381 -3216 -2343
rect -3328 -2415 -3289 -2381
rect -3255 -2415 -3216 -2381
rect -3328 -2453 -3216 -2415
rect -3328 -2487 -3289 -2453
rect -3255 -2487 -3216 -2453
rect -3328 -2525 -3216 -2487
rect -3328 -2559 -3289 -2525
rect -3255 -2559 -3216 -2525
rect -3328 -2597 -3216 -2559
rect -3328 -2631 -3289 -2597
rect -3255 -2631 -3216 -2597
rect -3328 -2669 -3216 -2631
rect -3328 -2703 -3289 -2669
rect -3255 -2703 -3216 -2669
rect -3328 -2741 -3216 -2703
rect -3328 -2775 -3289 -2741
rect -3255 -2775 -3216 -2741
rect -3128 -1251 3128 -1212
rect -3128 -1285 -3005 -1251
rect -2971 -1285 -2933 -1251
rect -2899 -1285 -2861 -1251
rect -2827 -1285 -2789 -1251
rect -2755 -1285 -2717 -1251
rect -2683 -1285 -2645 -1251
rect -2611 -1285 -2573 -1251
rect -2539 -1285 -2501 -1251
rect -2467 -1285 -2429 -1251
rect -2395 -1285 -2357 -1251
rect -2323 -1285 -2285 -1251
rect -2251 -1285 -2213 -1251
rect -2179 -1285 -2141 -1251
rect -2107 -1285 -2069 -1251
rect -2035 -1285 -1997 -1251
rect -1963 -1285 -1925 -1251
rect -1891 -1285 -1853 -1251
rect -1819 -1285 -1781 -1251
rect -1747 -1285 -1709 -1251
rect -1675 -1285 -1637 -1251
rect -1603 -1285 -1565 -1251
rect -1531 -1285 -1493 -1251
rect -1459 -1285 -1421 -1251
rect -1387 -1285 -1349 -1251
rect -1315 -1285 -1277 -1251
rect -1243 -1285 -1205 -1251
rect -1171 -1285 -1133 -1251
rect -1099 -1285 -1061 -1251
rect -1027 -1285 -989 -1251
rect -955 -1285 -917 -1251
rect -883 -1285 -845 -1251
rect -811 -1285 -773 -1251
rect -739 -1285 -701 -1251
rect -667 -1285 -629 -1251
rect -595 -1285 -557 -1251
rect -523 -1285 -485 -1251
rect -451 -1285 -413 -1251
rect -379 -1285 -341 -1251
rect -307 -1285 -269 -1251
rect -235 -1285 -197 -1251
rect -163 -1285 -125 -1251
rect -91 -1285 -53 -1251
rect -19 -1285 19 -1251
rect 53 -1285 91 -1251
rect 125 -1285 163 -1251
rect 197 -1285 235 -1251
rect 269 -1285 307 -1251
rect 341 -1285 379 -1251
rect 413 -1285 451 -1251
rect 485 -1285 523 -1251
rect 557 -1285 595 -1251
rect 629 -1285 667 -1251
rect 701 -1285 739 -1251
rect 773 -1285 811 -1251
rect 845 -1285 883 -1251
rect 917 -1285 955 -1251
rect 989 -1285 1027 -1251
rect 1061 -1285 1099 -1251
rect 1133 -1285 1171 -1251
rect 1205 -1285 1243 -1251
rect 1277 -1285 1315 -1251
rect 1349 -1285 1387 -1251
rect 1421 -1285 1459 -1251
rect 1493 -1285 1531 -1251
rect 1565 -1285 1603 -1251
rect 1637 -1285 1675 -1251
rect 1709 -1285 1747 -1251
rect 1781 -1285 1819 -1251
rect 1853 -1285 1891 -1251
rect 1925 -1285 1963 -1251
rect 1997 -1285 2035 -1251
rect 2069 -1285 2107 -1251
rect 2141 -1285 2179 -1251
rect 2213 -1285 2251 -1251
rect 2285 -1285 2323 -1251
rect 2357 -1285 2395 -1251
rect 2429 -1285 2467 -1251
rect 2501 -1285 2539 -1251
rect 2573 -1285 2611 -1251
rect 2645 -1285 2683 -1251
rect 2717 -1285 2755 -1251
rect 2789 -1285 2827 -1251
rect 2861 -1285 2899 -1251
rect 2933 -1285 2971 -1251
rect 3005 -1285 3128 -1251
rect -3128 -1324 3128 -1285
rect -3128 -1387 -3016 -1324
rect -3128 -1421 -3089 -1387
rect -3055 -1421 -3016 -1387
rect -3128 -1459 -3016 -1421
rect -3128 -1493 -3089 -1459
rect -3055 -1493 -3016 -1459
rect -2728 -1412 -2656 -1408
rect -2728 -1464 -2718 -1412
rect -2666 -1464 -2656 -1412
rect -1302 -1412 -1230 -1408
rect -2728 -1468 -2656 -1464
rect -3128 -1531 -3016 -1493
rect -3128 -1565 -3089 -1531
rect -3055 -1565 -3016 -1531
rect -3128 -1603 -3016 -1565
rect -3128 -1637 -3089 -1603
rect -3055 -1637 -3016 -1603
rect -3128 -1675 -3016 -1637
rect -3128 -1709 -3089 -1675
rect -3055 -1709 -3016 -1675
rect -3128 -1747 -3016 -1709
rect -3128 -1781 -3089 -1747
rect -3055 -1781 -3016 -1747
rect -3128 -1819 -3016 -1781
rect -3128 -1853 -3089 -1819
rect -3055 -1853 -3016 -1819
rect -3128 -1891 -3016 -1853
rect -3128 -1925 -3089 -1891
rect -3055 -1925 -3016 -1891
rect -3128 -1963 -3016 -1925
rect -3128 -1997 -3089 -1963
rect -3055 -1997 -3016 -1963
rect -3128 -2035 -3016 -1997
rect -3128 -2069 -3089 -2035
rect -3055 -2069 -3016 -2035
rect -3128 -2107 -3016 -2069
rect -3128 -2141 -3089 -2107
rect -3055 -2141 -3016 -2107
rect -3128 -2179 -3016 -2141
rect -3128 -2213 -3089 -2179
rect -3055 -2213 -3016 -2179
rect -3128 -2251 -3016 -2213
rect -3128 -2285 -3089 -2251
rect -3055 -2285 -3016 -2251
rect -3128 -2323 -3016 -2285
rect -3128 -2357 -3089 -2323
rect -3055 -2357 -3016 -2323
rect -3128 -2395 -3016 -2357
rect -3128 -2429 -3089 -2395
rect -3055 -2429 -3016 -2395
rect -2722 -2356 -2662 -1468
rect -2576 -1489 -1660 -1429
rect -1302 -1464 -1292 -1412
rect -1240 -1464 -1230 -1412
rect -1302 -1468 -1230 -1464
rect -434 -1412 -362 -1408
rect -434 -1464 -424 -1412
rect -372 -1464 -362 -1412
rect -434 -1468 -362 -1464
rect -8 -1412 64 -1408
rect -8 -1464 2 -1412
rect 54 -1464 64 -1412
rect -8 -1468 64 -1464
rect 418 -1412 490 -1408
rect 418 -1464 428 -1412
rect 480 -1464 490 -1412
rect 418 -1468 490 -1464
rect -2576 -1672 -2516 -1489
rect -2138 -1576 -2078 -1489
rect -1720 -1676 -1660 -1489
rect -1296 -1588 -1236 -1468
rect -428 -1582 -368 -1468
rect -2 -1674 58 -1468
rect 424 -1586 484 -1468
rect 854 -1680 914 -1324
rect 3016 -1387 3128 -1324
rect 1290 -1412 1362 -1408
rect 1290 -1464 1300 -1412
rect 1352 -1464 1362 -1412
rect 3016 -1421 3055 -1387
rect 3089 -1421 3128 -1387
rect 1290 -1468 1362 -1464
rect 1296 -1582 1356 -1468
rect 1712 -1489 2768 -1429
rect 1712 -1660 1772 -1489
rect 2132 -1576 2192 -1489
rect 2568 -1694 2628 -1489
rect -2582 -1892 -2522 -1742
rect -2588 -1896 -2516 -1892
rect -2588 -1948 -2578 -1896
rect -2526 -1948 -2516 -1896
rect -2588 -1952 -2516 -1948
rect -1286 -1998 -1226 -1851
rect -2576 -2356 -2516 -2160
rect -2138 -2356 -2078 -2269
rect -1720 -2356 -1660 -2166
rect -2722 -2416 -1660 -2356
rect -860 -2372 -800 -1765
rect -424 -1998 -364 -1851
rect 432 -1998 492 -1851
rect 852 -2088 912 -1761
rect 1284 -2002 1344 -1855
rect 2562 -1902 2634 -1898
rect 2562 -1954 2572 -1902
rect 2624 -1954 2634 -1902
rect 2562 -1958 2634 -1954
rect -866 -2376 -794 -2372
rect -3128 -2467 -3016 -2429
rect -866 -2428 -856 -2376
rect -804 -2428 -794 -2376
rect -866 -2432 -794 -2428
rect -3128 -2501 -3089 -2467
rect -3055 -2501 -3016 -2467
rect -3128 -2539 -3016 -2501
rect -3128 -2573 -3089 -2539
rect -3055 -2573 -3016 -2539
rect -3128 -2636 -3016 -2573
rect -860 -2636 -800 -2432
rect -2 -2486 58 -2178
rect 850 -2372 910 -2162
rect 1712 -2356 1772 -2160
rect 2150 -2356 2210 -2269
rect 2568 -2356 2628 -1958
rect 844 -2376 916 -2372
rect 844 -2428 854 -2376
rect 906 -2428 916 -2376
rect 1712 -2416 2628 -2356
rect 844 -2432 916 -2428
rect -8 -2490 64 -2486
rect -8 -2542 2 -2490
rect 54 -2542 64 -2490
rect -8 -2546 64 -2542
rect 850 -2636 910 -2432
rect 2708 -2486 2768 -1489
rect 3016 -1459 3128 -1421
rect 3016 -1493 3055 -1459
rect 3089 -1493 3128 -1459
rect 3016 -1531 3128 -1493
rect 3016 -1565 3055 -1531
rect 3089 -1565 3128 -1531
rect 3016 -1603 3128 -1565
rect 3016 -1637 3055 -1603
rect 3089 -1637 3128 -1603
rect 3016 -1675 3128 -1637
rect 3016 -1709 3055 -1675
rect 3089 -1709 3128 -1675
rect 3016 -1747 3128 -1709
rect 3016 -1781 3055 -1747
rect 3089 -1781 3128 -1747
rect 3016 -1819 3128 -1781
rect 3016 -1853 3055 -1819
rect 3089 -1853 3128 -1819
rect 3016 -1891 3128 -1853
rect 3016 -1925 3055 -1891
rect 3089 -1925 3128 -1891
rect 3016 -1963 3128 -1925
rect 3016 -1997 3055 -1963
rect 3089 -1997 3128 -1963
rect 3016 -2035 3128 -1997
rect 3016 -2069 3055 -2035
rect 3089 -2069 3128 -2035
rect 3016 -2107 3128 -2069
rect 3016 -2141 3055 -2107
rect 3089 -2141 3128 -2107
rect 3016 -2179 3128 -2141
rect 3016 -2213 3055 -2179
rect 3089 -2213 3128 -2179
rect 3016 -2251 3128 -2213
rect 3016 -2285 3055 -2251
rect 3089 -2285 3128 -2251
rect 3016 -2323 3128 -2285
rect 3016 -2357 3055 -2323
rect 3089 -2357 3128 -2323
rect 3016 -2395 3128 -2357
rect 3016 -2429 3055 -2395
rect 3089 -2429 3128 -2395
rect 3016 -2467 3128 -2429
rect 2702 -2490 2774 -2486
rect 2702 -2542 2712 -2490
rect 2764 -2542 2774 -2490
rect 2702 -2546 2774 -2542
rect 3016 -2501 3055 -2467
rect 3089 -2501 3128 -2467
rect 3016 -2539 3128 -2501
rect 3016 -2573 3055 -2539
rect 3089 -2573 3128 -2539
rect 3016 -2636 3128 -2573
rect -3128 -2675 3128 -2636
rect -3128 -2709 -3005 -2675
rect -2971 -2709 -2933 -2675
rect -2899 -2709 -2861 -2675
rect -2827 -2709 -2789 -2675
rect -2755 -2709 -2717 -2675
rect -2683 -2709 -2645 -2675
rect -2611 -2709 -2573 -2675
rect -2539 -2709 -2501 -2675
rect -2467 -2709 -2429 -2675
rect -2395 -2709 -2357 -2675
rect -2323 -2709 -2285 -2675
rect -2251 -2709 -2213 -2675
rect -2179 -2709 -2141 -2675
rect -2107 -2709 -2069 -2675
rect -2035 -2709 -1997 -2675
rect -1963 -2709 -1925 -2675
rect -1891 -2709 -1853 -2675
rect -1819 -2709 -1781 -2675
rect -1747 -2709 -1709 -2675
rect -1675 -2709 -1637 -2675
rect -1603 -2709 -1565 -2675
rect -1531 -2709 -1493 -2675
rect -1459 -2709 -1421 -2675
rect -1387 -2709 -1349 -2675
rect -1315 -2709 -1277 -2675
rect -1243 -2709 -1205 -2675
rect -1171 -2709 -1133 -2675
rect -1099 -2709 -1061 -2675
rect -1027 -2709 -989 -2675
rect -955 -2709 -917 -2675
rect -883 -2709 -845 -2675
rect -811 -2709 -773 -2675
rect -739 -2709 -701 -2675
rect -667 -2709 -629 -2675
rect -595 -2709 -557 -2675
rect -523 -2709 -485 -2675
rect -451 -2709 -413 -2675
rect -379 -2709 -341 -2675
rect -307 -2709 -269 -2675
rect -235 -2709 -197 -2675
rect -163 -2709 -125 -2675
rect -91 -2709 -53 -2675
rect -19 -2709 19 -2675
rect 53 -2709 91 -2675
rect 125 -2709 163 -2675
rect 197 -2709 235 -2675
rect 269 -2709 307 -2675
rect 341 -2709 379 -2675
rect 413 -2709 451 -2675
rect 485 -2709 523 -2675
rect 557 -2709 595 -2675
rect 629 -2709 667 -2675
rect 701 -2709 739 -2675
rect 773 -2709 811 -2675
rect 845 -2709 883 -2675
rect 917 -2709 955 -2675
rect 989 -2709 1027 -2675
rect 1061 -2709 1099 -2675
rect 1133 -2709 1171 -2675
rect 1205 -2709 1243 -2675
rect 1277 -2709 1315 -2675
rect 1349 -2709 1387 -2675
rect 1421 -2709 1459 -2675
rect 1493 -2709 1531 -2675
rect 1565 -2709 1603 -2675
rect 1637 -2709 1675 -2675
rect 1709 -2709 1747 -2675
rect 1781 -2709 1819 -2675
rect 1853 -2709 1891 -2675
rect 1925 -2709 1963 -2675
rect 1997 -2709 2035 -2675
rect 2069 -2709 2107 -2675
rect 2141 -2709 2179 -2675
rect 2213 -2709 2251 -2675
rect 2285 -2709 2323 -2675
rect 2357 -2709 2395 -2675
rect 2429 -2709 2467 -2675
rect 2501 -2709 2539 -2675
rect 2573 -2709 2611 -2675
rect 2645 -2709 2683 -2675
rect 2717 -2709 2755 -2675
rect 2789 -2709 2827 -2675
rect 2861 -2709 2899 -2675
rect 2933 -2709 2971 -2675
rect 3005 -2709 3128 -2675
rect -3128 -2748 3128 -2709
rect 3216 -1229 3328 -1191
rect 3216 -1263 3255 -1229
rect 3289 -1263 3328 -1229
rect 3216 -1301 3328 -1263
rect 3216 -1335 3255 -1301
rect 3289 -1335 3328 -1301
rect 3216 -1373 3328 -1335
rect 3216 -1407 3255 -1373
rect 3289 -1407 3328 -1373
rect 3216 -1445 3328 -1407
rect 3216 -1479 3255 -1445
rect 3289 -1479 3328 -1445
rect 3216 -1517 3328 -1479
rect 3216 -1551 3255 -1517
rect 3289 -1551 3328 -1517
rect 3216 -1589 3328 -1551
rect 3216 -1623 3255 -1589
rect 3289 -1623 3328 -1589
rect 3216 -1661 3328 -1623
rect 3216 -1695 3255 -1661
rect 3289 -1695 3328 -1661
rect 3216 -1733 3328 -1695
rect 3216 -1767 3255 -1733
rect 3289 -1767 3328 -1733
rect 3216 -1805 3328 -1767
rect 3216 -1839 3255 -1805
rect 3289 -1839 3328 -1805
rect 3216 -1877 3328 -1839
rect 3216 -1911 3255 -1877
rect 3289 -1911 3328 -1877
rect 3216 -1949 3328 -1911
rect 3216 -1983 3255 -1949
rect 3289 -1983 3328 -1949
rect 3216 -2021 3328 -1983
rect 3216 -2055 3255 -2021
rect 3289 -2055 3328 -2021
rect 3216 -2093 3328 -2055
rect 3216 -2127 3255 -2093
rect 3289 -2127 3328 -2093
rect 3216 -2165 3328 -2127
rect 3216 -2199 3255 -2165
rect 3289 -2199 3328 -2165
rect 3216 -2237 3328 -2199
rect 3216 -2271 3255 -2237
rect 3289 -2271 3328 -2237
rect 3216 -2309 3328 -2271
rect 3216 -2343 3255 -2309
rect 3289 -2343 3328 -2309
rect 3216 -2381 3328 -2343
rect 3216 -2415 3255 -2381
rect 3289 -2415 3328 -2381
rect 3216 -2453 3328 -2415
rect 3216 -2487 3255 -2453
rect 3289 -2487 3328 -2453
rect 3216 -2525 3328 -2487
rect 3216 -2559 3255 -2525
rect 3289 -2559 3328 -2525
rect 3216 -2597 3328 -2559
rect 3216 -2631 3255 -2597
rect 3289 -2631 3328 -2597
rect 3216 -2669 3328 -2631
rect 3216 -2703 3255 -2669
rect 3289 -2703 3328 -2669
rect 3216 -2741 3328 -2703
rect -3328 -2813 -3216 -2775
rect -3328 -2847 -3289 -2813
rect -3255 -2847 -3216 -2813
rect -860 -2836 -800 -2748
rect 850 -2836 910 -2748
rect 3216 -2775 3255 -2741
rect 3289 -2775 3328 -2741
rect 3216 -2813 3328 -2775
rect -3328 -2885 -3216 -2847
rect -3328 -2919 -3289 -2885
rect -3255 -2919 -3216 -2885
rect -3328 -2957 -3216 -2919
rect -3328 -2991 -3289 -2957
rect -3255 -2991 -3216 -2957
rect -3328 -3029 -3216 -2991
rect -928 -2893 970 -2836
rect -928 -2945 -868 -2893
rect -816 -2945 -804 -2893
rect -752 -2945 -740 -2893
rect -688 -2945 -676 -2893
rect -624 -2945 -612 -2893
rect -560 -2945 -548 -2893
rect -496 -2945 -484 -2893
rect -432 -2945 -420 -2893
rect -368 -2945 -356 -2893
rect -304 -2945 -292 -2893
rect -240 -2945 -228 -2893
rect -176 -2945 -164 -2893
rect -112 -2945 -100 -2893
rect -48 -2945 -36 -2893
rect 16 -2945 28 -2893
rect 80 -2945 92 -2893
rect 144 -2945 156 -2893
rect 208 -2945 220 -2893
rect 272 -2945 284 -2893
rect 336 -2945 348 -2893
rect 400 -2945 412 -2893
rect 464 -2945 476 -2893
rect 528 -2945 540 -2893
rect 592 -2945 604 -2893
rect 656 -2945 668 -2893
rect 720 -2945 732 -2893
rect 784 -2945 796 -2893
rect 848 -2945 860 -2893
rect 912 -2945 970 -2893
rect -928 -3002 970 -2945
rect 3216 -2847 3255 -2813
rect 3289 -2847 3328 -2813
rect 3216 -2885 3328 -2847
rect 3216 -2919 3255 -2885
rect 3289 -2919 3328 -2885
rect 3216 -2957 3328 -2919
rect 3216 -2991 3255 -2957
rect 3289 -2991 3328 -2957
rect -3328 -3063 -3289 -3029
rect -3255 -3063 -3216 -3029
rect -3328 -3101 -3216 -3063
rect -3328 -3135 -3289 -3101
rect -3255 -3116 -3216 -3101
rect 3216 -3029 3328 -2991
rect 3216 -3063 3255 -3029
rect 3289 -3063 3328 -3029
rect 3216 -3101 3328 -3063
rect 3216 -3116 3255 -3101
rect -3255 -3135 -2606 -3116
rect -3328 -3144 -2606 -3135
rect -3328 -3173 -3198 -3144
rect -3328 -3207 -3289 -3173
rect -3255 -3207 -3198 -3173
rect -3328 -3388 -3198 -3207
rect -2634 -3388 -2606 -3144
rect -3328 -3416 -2606 -3388
rect 2606 -3135 3255 -3116
rect 3289 -3135 3328 -3101
rect 2606 -3144 3328 -3135
rect 2606 -3388 2634 -3144
rect 3198 -3173 3328 -3144
rect 3198 -3207 3255 -3173
rect 3289 -3207 3328 -3173
rect 3198 -3388 3328 -3207
rect 2606 -3416 3328 -3388
rect -3328 -3455 3328 -3416
rect -3328 -3489 -3221 -3455
rect -3187 -3489 -3149 -3455
rect -3115 -3489 -3077 -3455
rect -3043 -3489 -3005 -3455
rect -2971 -3489 -2933 -3455
rect -2899 -3489 -2861 -3455
rect -2827 -3489 -2789 -3455
rect -2755 -3489 -2717 -3455
rect -2683 -3489 -2645 -3455
rect -2611 -3489 -2573 -3455
rect -2539 -3489 -2501 -3455
rect -2467 -3489 -2429 -3455
rect -2395 -3489 -2357 -3455
rect -2323 -3489 -2285 -3455
rect -2251 -3489 -2213 -3455
rect -2179 -3489 -2141 -3455
rect -2107 -3489 -2069 -3455
rect -2035 -3489 -1997 -3455
rect -1963 -3489 -1925 -3455
rect -1891 -3489 -1853 -3455
rect -1819 -3489 -1781 -3455
rect -1747 -3489 -1709 -3455
rect -1675 -3489 -1637 -3455
rect -1603 -3489 -1565 -3455
rect -1531 -3489 -1493 -3455
rect -1459 -3489 -1421 -3455
rect -1387 -3489 -1349 -3455
rect -1315 -3489 -1277 -3455
rect -1243 -3489 -1205 -3455
rect -1171 -3489 -1133 -3455
rect -1099 -3489 -1061 -3455
rect -1027 -3489 -989 -3455
rect -955 -3489 -917 -3455
rect -883 -3489 -845 -3455
rect -811 -3489 -773 -3455
rect -739 -3489 -701 -3455
rect -667 -3489 -629 -3455
rect -595 -3489 -557 -3455
rect -523 -3489 -485 -3455
rect -451 -3489 -413 -3455
rect -379 -3489 -341 -3455
rect -307 -3489 -269 -3455
rect -235 -3489 -197 -3455
rect -163 -3489 -125 -3455
rect -91 -3489 -53 -3455
rect -19 -3489 19 -3455
rect 53 -3489 91 -3455
rect 125 -3489 163 -3455
rect 197 -3489 235 -3455
rect 269 -3489 307 -3455
rect 341 -3489 379 -3455
rect 413 -3489 451 -3455
rect 485 -3489 523 -3455
rect 557 -3489 595 -3455
rect 629 -3489 667 -3455
rect 701 -3489 739 -3455
rect 773 -3489 811 -3455
rect 845 -3489 883 -3455
rect 917 -3489 955 -3455
rect 989 -3489 1027 -3455
rect 1061 -3489 1099 -3455
rect 1133 -3489 1171 -3455
rect 1205 -3489 1243 -3455
rect 1277 -3489 1315 -3455
rect 1349 -3489 1387 -3455
rect 1421 -3489 1459 -3455
rect 1493 -3489 1531 -3455
rect 1565 -3489 1603 -3455
rect 1637 -3489 1675 -3455
rect 1709 -3489 1747 -3455
rect 1781 -3489 1819 -3455
rect 1853 -3489 1891 -3455
rect 1925 -3489 1963 -3455
rect 1997 -3489 2035 -3455
rect 2069 -3489 2107 -3455
rect 2141 -3489 2179 -3455
rect 2213 -3489 2251 -3455
rect 2285 -3489 2323 -3455
rect 2357 -3489 2395 -3455
rect 2429 -3489 2467 -3455
rect 2501 -3489 2539 -3455
rect 2573 -3489 2611 -3455
rect 2645 -3489 2683 -3455
rect 2717 -3489 2755 -3455
rect 2789 -3489 2827 -3455
rect 2861 -3489 2899 -3455
rect 2933 -3489 2971 -3455
rect 3005 -3489 3043 -3455
rect 3077 -3489 3115 -3455
rect 3149 -3489 3187 -3455
rect 3221 -3489 3328 -3455
rect -3328 -3528 3328 -3489
<< via1 >>
rect -3198 2744 -2634 2988
rect 2634 2744 3198 2988
rect -2637 2466 -2585 2518
rect -2573 2466 -2521 2518
rect -2509 2466 -2457 2518
rect -2445 2466 -2393 2518
rect -2381 2466 -2329 2518
rect -2317 2466 -2265 2518
rect -2253 2466 -2201 2518
rect -2189 2466 -2137 2518
rect -2125 2466 -2073 2518
rect -2061 2466 -2009 2518
rect -1997 2466 -1945 2518
rect -1933 2466 -1881 2518
rect -1869 2466 -1817 2518
rect -1805 2466 -1753 2518
rect -1741 2466 -1689 2518
rect -1677 2466 -1625 2518
rect -1613 2466 -1561 2518
rect -1549 2466 -1497 2518
rect -1485 2466 -1433 2518
rect -1421 2466 -1369 2518
rect -1357 2466 -1305 2518
rect -1293 2466 -1241 2518
rect -1229 2466 -1177 2518
rect -1165 2466 -1113 2518
rect -1101 2466 -1049 2518
rect -1037 2466 -985 2518
rect -973 2466 -921 2518
rect -909 2466 -857 2518
rect -845 2466 -793 2518
rect -781 2466 -729 2518
rect -717 2466 -665 2518
rect -653 2466 -601 2518
rect -589 2466 -537 2518
rect -525 2466 -473 2518
rect -461 2466 -409 2518
rect -397 2466 -345 2518
rect -333 2466 -281 2518
rect -269 2466 -217 2518
rect -205 2466 -153 2518
rect -141 2466 -89 2518
rect -77 2466 -25 2518
rect -13 2466 39 2518
rect 51 2466 103 2518
rect 115 2466 167 2518
rect 179 2466 231 2518
rect 243 2466 295 2518
rect 307 2466 359 2518
rect 371 2466 423 2518
rect 435 2466 487 2518
rect 499 2466 551 2518
rect 563 2466 615 2518
rect 627 2466 679 2518
rect 691 2466 743 2518
rect 755 2466 807 2518
rect 819 2466 871 2518
rect 883 2466 935 2518
rect 947 2466 999 2518
rect 1011 2466 1063 2518
rect 1075 2466 1127 2518
rect 1139 2466 1191 2518
rect 1203 2466 1255 2518
rect 1267 2466 1319 2518
rect 1331 2466 1383 2518
rect 1395 2466 1447 2518
rect 1459 2466 1511 2518
rect 1523 2466 1575 2518
rect 1587 2466 1639 2518
rect 1651 2466 1703 2518
rect 1715 2466 1767 2518
rect 1779 2466 1831 2518
rect 1843 2466 1895 2518
rect 1907 2466 1959 2518
rect 1971 2466 2023 2518
rect 2035 2466 2087 2518
rect 2099 2466 2151 2518
rect 2163 2466 2215 2518
rect 2227 2466 2279 2518
rect 2291 2466 2343 2518
rect 2355 2466 2407 2518
rect 2419 2466 2471 2518
rect 2483 2466 2535 2518
rect -2772 2150 -2720 2202
rect -2262 2150 -2210 2202
rect -2266 1608 -2214 1660
rect -2134 1474 -2082 1526
rect -2004 1474 -1952 1526
rect -1618 2150 -1566 2202
rect -1492 2150 -1440 2202
rect -1490 1608 -1438 1660
rect -1746 1474 -1694 1526
rect -1624 1474 -1572 1526
rect -1228 2150 -1176 2202
rect -1236 1608 -1184 1660
rect -1108 1474 -1056 1526
rect -976 1474 -924 1526
rect -592 2150 -540 2202
rect -460 2150 -408 2202
rect -460 1608 -408 1660
rect -716 1474 -664 1526
rect -592 1474 -540 1526
rect 220 2262 272 2314
rect 604 2262 656 2314
rect -2772 922 -2720 974
rect -2270 922 -2218 974
rect -2138 922 -2086 974
rect -1496 922 -1444 974
rect -1236 922 -1184 974
rect -1104 922 -1052 974
rect -2010 818 -1958 870
rect -460 922 -408 974
rect 734 1606 786 1658
rect 602 1482 654 1534
rect 992 2150 1044 2202
rect 1248 2150 1300 2202
rect 992 1606 1044 1658
rect 1250 1606 1302 1658
rect 1120 1482 1172 1534
rect 1636 2262 1688 2314
rect 2006 2150 2058 2202
rect 1504 1606 1556 1658
rect 1634 1482 1686 1534
rect 732 930 784 982
rect 2436 2098 2488 2150
rect 1506 930 1558 982
rect 2006 930 2058 982
rect 2436 928 2488 980
rect 2560 920 2612 972
rect -720 810 -668 862
rect 220 818 272 870
rect 1118 818 1170 870
rect -2102 -42 -2050 10
rect -1068 -42 -1016 10
rect -2618 -158 -2566 -106
rect -2486 -276 -2434 -224
rect -1582 -158 -1530 -106
rect -1710 -276 -1658 -224
rect -1456 -276 -1404 -224
rect -552 -158 -500 -106
rect 1118 -122 1170 -70
rect 2436 -120 2488 -68
rect -676 -276 -624 -224
rect -2226 -812 -2174 -760
rect -1970 -812 -1918 -760
rect -1196 -812 -1144 -760
rect -938 -812 -886 -760
rect 600 -758 652 -706
rect -2358 -930 -2306 -878
rect -1842 -930 -1790 -878
rect -1322 -930 -1270 -878
rect -810 -930 -758 -878
rect 2560 -128 2612 -76
rect 1634 -758 1686 -706
rect 2436 -944 2488 -892
rect -2718 -1464 -2666 -1412
rect -1292 -1464 -1240 -1412
rect -424 -1464 -372 -1412
rect 2 -1464 54 -1412
rect 428 -1464 480 -1412
rect 1300 -1464 1352 -1412
rect -2578 -1948 -2526 -1896
rect 2572 -1954 2624 -1902
rect -856 -2428 -804 -2376
rect 854 -2428 906 -2376
rect 2 -2542 54 -2490
rect 2712 -2542 2764 -2490
rect -868 -2945 -816 -2893
rect -804 -2945 -752 -2893
rect -740 -2945 -688 -2893
rect -676 -2945 -624 -2893
rect -612 -2945 -560 -2893
rect -548 -2945 -496 -2893
rect -484 -2945 -432 -2893
rect -420 -2945 -368 -2893
rect -356 -2945 -304 -2893
rect -292 -2945 -240 -2893
rect -228 -2945 -176 -2893
rect -164 -2945 -112 -2893
rect -100 -2945 -48 -2893
rect -36 -2945 16 -2893
rect 28 -2945 80 -2893
rect 92 -2945 144 -2893
rect 156 -2945 208 -2893
rect 220 -2945 272 -2893
rect 284 -2945 336 -2893
rect 348 -2945 400 -2893
rect 412 -2945 464 -2893
rect 476 -2945 528 -2893
rect 540 -2945 592 -2893
rect 604 -2945 656 -2893
rect 668 -2945 720 -2893
rect 732 -2945 784 -2893
rect 796 -2945 848 -2893
rect 860 -2945 912 -2893
rect -3198 -3388 -2634 -3144
rect 2634 -3388 3198 -3144
<< metal2 >>
rect -3216 3014 -2616 3026
rect -3216 2988 -3184 3014
rect -2648 2988 -2616 3014
rect -3216 2744 -3198 2988
rect -2634 2744 -2616 2988
rect -3216 2718 -3184 2744
rect -2648 2718 -2616 2744
rect -3216 2706 -2616 2718
rect 2616 3014 3216 3026
rect 2616 2988 2648 3014
rect 3184 2988 3216 3014
rect 2616 2744 2634 2988
rect 3198 2744 3216 2988
rect 2616 2718 2648 2744
rect 3184 2718 3216 2744
rect 2616 2706 3216 2718
rect -2674 2520 2566 2562
rect -2674 2464 -2639 2520
rect -2583 2518 -2559 2520
rect -2503 2518 -2479 2520
rect -2423 2518 -2399 2520
rect -2343 2518 -2319 2520
rect -2263 2518 -2239 2520
rect -2183 2518 -2159 2520
rect -2103 2518 -2079 2520
rect -2023 2518 -1999 2520
rect -1943 2518 -1919 2520
rect -1863 2518 -1839 2520
rect -1783 2518 -1759 2520
rect -1703 2518 -1679 2520
rect -1623 2518 -1599 2520
rect -1543 2518 -1519 2520
rect -1463 2518 -1439 2520
rect -1383 2518 -1359 2520
rect -1303 2518 -1279 2520
rect -1223 2518 -1199 2520
rect -1143 2518 -1119 2520
rect -1063 2518 -1039 2520
rect -983 2518 -959 2520
rect -903 2518 -879 2520
rect -823 2518 -799 2520
rect -743 2518 -719 2520
rect -663 2518 -639 2520
rect -583 2518 -559 2520
rect -503 2518 -479 2520
rect -423 2518 -399 2520
rect -343 2518 -319 2520
rect -263 2518 -239 2520
rect -183 2518 -159 2520
rect -103 2518 -79 2520
rect -23 2518 1 2520
rect 57 2518 81 2520
rect 137 2518 161 2520
rect 217 2518 241 2520
rect 297 2518 321 2520
rect 377 2518 401 2520
rect 457 2518 481 2520
rect 537 2518 561 2520
rect 617 2518 641 2520
rect 697 2518 721 2520
rect 777 2518 801 2520
rect 857 2518 881 2520
rect 937 2518 961 2520
rect 1017 2518 1041 2520
rect 1097 2518 1121 2520
rect 1177 2518 1201 2520
rect 1257 2518 1281 2520
rect 1337 2518 1361 2520
rect 1417 2518 1441 2520
rect 1497 2518 1521 2520
rect 1577 2518 1601 2520
rect 1657 2518 1681 2520
rect 1737 2518 1761 2520
rect 1817 2518 1841 2520
rect 1897 2518 1921 2520
rect 1977 2518 2001 2520
rect 2057 2518 2081 2520
rect 2137 2518 2161 2520
rect 2217 2518 2241 2520
rect 2297 2518 2321 2520
rect 2377 2518 2401 2520
rect 2457 2518 2481 2520
rect -2583 2466 -2573 2518
rect -2329 2466 -2319 2518
rect -2263 2466 -2253 2518
rect -2009 2466 -1999 2518
rect -1943 2466 -1933 2518
rect -1689 2466 -1679 2518
rect -1623 2466 -1613 2518
rect -1369 2466 -1359 2518
rect -1303 2466 -1293 2518
rect -1049 2466 -1039 2518
rect -983 2466 -973 2518
rect -729 2466 -719 2518
rect -663 2466 -653 2518
rect -409 2466 -399 2518
rect -343 2466 -333 2518
rect -89 2466 -79 2518
rect -23 2466 -13 2518
rect 231 2466 241 2518
rect 297 2466 307 2518
rect 551 2466 561 2518
rect 617 2466 627 2518
rect 871 2466 881 2518
rect 937 2466 947 2518
rect 1191 2466 1201 2518
rect 1257 2466 1267 2518
rect 1511 2466 1521 2518
rect 1577 2466 1587 2518
rect 1831 2466 1841 2518
rect 1897 2466 1907 2518
rect 2151 2466 2161 2518
rect 2217 2466 2227 2518
rect 2471 2466 2481 2518
rect -2583 2464 -2559 2466
rect -2503 2464 -2479 2466
rect -2423 2464 -2399 2466
rect -2343 2464 -2319 2466
rect -2263 2464 -2239 2466
rect -2183 2464 -2159 2466
rect -2103 2464 -2079 2466
rect -2023 2464 -1999 2466
rect -1943 2464 -1919 2466
rect -1863 2464 -1839 2466
rect -1783 2464 -1759 2466
rect -1703 2464 -1679 2466
rect -1623 2464 -1599 2466
rect -1543 2464 -1519 2466
rect -1463 2464 -1439 2466
rect -1383 2464 -1359 2466
rect -1303 2464 -1279 2466
rect -1223 2464 -1199 2466
rect -1143 2464 -1119 2466
rect -1063 2464 -1039 2466
rect -983 2464 -959 2466
rect -903 2464 -879 2466
rect -823 2464 -799 2466
rect -743 2464 -719 2466
rect -663 2464 -639 2466
rect -583 2464 -559 2466
rect -503 2464 -479 2466
rect -423 2464 -399 2466
rect -343 2464 -319 2466
rect -263 2464 -239 2466
rect -183 2464 -159 2466
rect -103 2464 -79 2466
rect -23 2464 1 2466
rect 57 2464 81 2466
rect 137 2464 161 2466
rect 217 2464 241 2466
rect 297 2464 321 2466
rect 377 2464 401 2466
rect 457 2464 481 2466
rect 537 2464 561 2466
rect 617 2464 641 2466
rect 697 2464 721 2466
rect 777 2464 801 2466
rect 857 2464 881 2466
rect 937 2464 961 2466
rect 1017 2464 1041 2466
rect 1097 2464 1121 2466
rect 1177 2464 1201 2466
rect 1257 2464 1281 2466
rect 1337 2464 1361 2466
rect 1417 2464 1441 2466
rect 1497 2464 1521 2466
rect 1577 2464 1601 2466
rect 1657 2464 1681 2466
rect 1737 2464 1761 2466
rect 1817 2464 1841 2466
rect 1897 2464 1921 2466
rect 1977 2464 2001 2466
rect 2057 2464 2081 2466
rect 2137 2464 2161 2466
rect 2217 2464 2241 2466
rect 2297 2464 2321 2466
rect 2377 2464 2401 2466
rect 2457 2464 2481 2466
rect 2537 2464 2566 2520
rect -2674 2430 2566 2464
rect 216 2318 276 2324
rect 600 2318 660 2324
rect 1632 2318 1692 2324
rect 216 2314 1692 2318
rect 216 2262 220 2314
rect 272 2262 604 2314
rect 656 2262 1636 2314
rect 1688 2262 1692 2314
rect 216 2258 1692 2262
rect 216 2252 276 2258
rect 600 2252 660 2258
rect 1632 2252 1692 2258
rect -2776 2206 -2716 2212
rect -2266 2206 -2206 2212
rect -1622 2206 -1562 2212
rect -1496 2206 -1436 2212
rect -1232 2206 -1172 2212
rect -596 2206 -536 2212
rect -464 2206 -404 2212
rect 988 2206 1048 2212
rect 1244 2206 1304 2212
rect 2002 2206 2062 2212
rect -2776 2202 2062 2206
rect -2776 2150 -2772 2202
rect -2720 2150 -2262 2202
rect -2210 2150 -1618 2202
rect -1566 2150 -1492 2202
rect -1440 2150 -1228 2202
rect -1176 2150 -592 2202
rect -540 2150 -460 2202
rect -408 2150 992 2202
rect 1044 2150 1248 2202
rect 1300 2150 2006 2202
rect 2058 2150 2062 2202
rect 2432 2154 2492 2160
rect -2776 2146 2062 2150
rect -2776 2140 -2716 2146
rect -2266 2140 -2206 2146
rect -1622 2140 -1562 2146
rect -1496 2140 -1436 2146
rect -1232 2140 -1172 2146
rect -596 2140 -536 2146
rect -464 2140 -404 2146
rect 988 2140 1048 2146
rect 1244 2140 1304 2146
rect 2002 2140 2062 2146
rect 2132 2150 2492 2154
rect 2132 2098 2436 2150
rect 2488 2098 2492 2150
rect 2132 2094 2492 2098
rect -2270 1664 -2210 1670
rect -1494 1664 -1434 1670
rect -1240 1664 -1180 1670
rect -464 1664 -404 1670
rect -2270 1660 -404 1664
rect 730 1662 790 1668
rect 988 1662 1048 1668
rect 1246 1662 1306 1668
rect 1500 1662 1560 1668
rect -2270 1608 -2266 1660
rect -2214 1608 -1490 1660
rect -1438 1608 -1236 1660
rect -1184 1608 -460 1660
rect -408 1608 -404 1660
rect -2270 1604 -404 1608
rect -2270 1598 -2210 1604
rect -1494 1598 -1434 1604
rect -1240 1598 -1180 1604
rect -464 1598 -404 1604
rect 72 1658 1560 1662
rect 72 1606 734 1658
rect 786 1606 992 1658
rect 1044 1606 1250 1658
rect 1302 1606 1504 1658
rect 1556 1606 1560 1658
rect 72 1602 1560 1606
rect -2138 1530 -2078 1536
rect -2008 1530 -1948 1536
rect -1750 1530 -1690 1536
rect -1628 1530 -1568 1536
rect -1112 1530 -1052 1536
rect -980 1530 -920 1536
rect -720 1530 -660 1536
rect -596 1530 -536 1536
rect 72 1530 132 1602
rect 730 1596 790 1602
rect 988 1596 1048 1602
rect 1246 1596 1306 1602
rect 1500 1596 1560 1602
rect -2138 1526 132 1530
rect -2138 1474 -2134 1526
rect -2082 1474 -2004 1526
rect -1952 1474 -1746 1526
rect -1694 1474 -1624 1526
rect -1572 1474 -1108 1526
rect -1056 1474 -976 1526
rect -924 1474 -716 1526
rect -664 1474 -592 1526
rect -540 1474 132 1526
rect -2138 1470 132 1474
rect 598 1538 658 1544
rect 1116 1538 1176 1544
rect 1630 1538 1690 1544
rect 2132 1538 2192 2094
rect 2432 2088 2492 2094
rect 598 1534 2192 1538
rect 598 1482 602 1534
rect 654 1482 1120 1534
rect 1172 1482 1634 1534
rect 1686 1482 2192 1534
rect 598 1478 2192 1482
rect 598 1472 658 1478
rect 1116 1472 1176 1478
rect 1630 1472 1690 1478
rect -2138 1464 -2078 1470
rect -2008 1464 -1948 1470
rect -1750 1464 -1690 1470
rect -1628 1464 -1568 1470
rect -1112 1464 -1052 1470
rect -980 1464 -920 1470
rect -720 1464 -660 1470
rect -596 1464 -536 1470
rect 728 986 788 992
rect 1502 986 1562 992
rect 2002 986 2062 992
rect -2776 978 -2716 984
rect -2274 978 -2214 984
rect -2142 978 -2082 984
rect -1500 978 -1440 984
rect -1240 978 -1180 984
rect -1108 978 -1048 984
rect -464 978 -404 984
rect -2776 974 -404 978
rect -2776 922 -2772 974
rect -2720 922 -2270 974
rect -2218 922 -2138 974
rect -2086 922 -1496 974
rect -1444 922 -1236 974
rect -1184 922 -1104 974
rect -1052 922 -460 974
rect -408 922 -404 974
rect -2776 918 -404 922
rect 728 982 2062 986
rect 728 930 732 982
rect 784 930 1506 982
rect 1558 930 2006 982
rect 2058 930 2062 982
rect 728 926 2062 930
rect 728 920 788 926
rect 1502 920 1562 926
rect 2002 920 2062 926
rect -2776 912 -2716 918
rect -2274 912 -2214 918
rect -2142 912 -2082 918
rect -2014 870 -1954 880
rect -2014 818 -2010 870
rect -1958 818 -1954 870
rect -2014 534 -1954 818
rect -2234 474 -1954 534
rect -2622 -102 -2562 -96
rect -2234 -102 -2174 474
rect -2106 14 -2046 20
rect -1748 14 -1688 918
rect -1500 912 -1440 918
rect -1370 14 -1310 918
rect -1240 912 -1180 918
rect -1108 912 -1048 918
rect -464 912 -404 918
rect 216 874 276 880
rect 1114 874 1174 880
rect 216 870 1174 874
rect -730 862 -658 866
rect -730 810 -720 862
rect -668 810 -658 862
rect -730 806 -658 810
rect 216 818 220 870
rect 272 818 1118 870
rect 1170 818 1174 870
rect 216 814 1174 818
rect 216 808 276 814
rect -1072 14 -1012 20
rect -2106 10 -1012 14
rect -2106 -42 -2102 10
rect -2050 -42 -1068 10
rect -1016 -42 -1012 10
rect -2106 -46 -1012 -42
rect -2106 -52 -2046 -46
rect -1072 -52 -1012 -46
rect -1586 -102 -1526 -96
rect -724 -102 -664 806
rect 1114 -66 1174 814
rect 2132 254 2192 1478
rect 2426 980 2498 984
rect 2426 928 2436 980
rect 2488 928 2498 980
rect 2426 924 2498 928
rect 2556 972 2616 982
rect 2432 254 2492 924
rect 2132 194 2492 254
rect 1108 -70 1180 -66
rect -556 -102 -496 -96
rect -2622 -106 -496 -102
rect -2622 -158 -2618 -106
rect -2566 -158 -1582 -106
rect -1530 -158 -552 -106
rect -500 -158 -496 -106
rect 1108 -122 1118 -70
rect 1170 -122 1180 -70
rect 1108 -126 1180 -122
rect -2622 -162 -496 -158
rect -2622 -168 -2562 -162
rect -1586 -168 -1526 -162
rect -556 -168 -496 -162
rect -2490 -220 -2430 -214
rect -1714 -220 -1654 -214
rect -1460 -220 -1400 -214
rect -680 -220 -620 -214
rect -2490 -224 -620 -220
rect -2490 -276 -2486 -224
rect -2434 -276 -1710 -224
rect -1658 -276 -1456 -224
rect -1404 -276 -676 -224
rect -624 -276 -620 -224
rect -2490 -280 -620 -276
rect -2490 -286 -2430 -280
rect -1714 -286 -1654 -280
rect -1460 -286 -1400 -280
rect -680 -286 -620 -280
rect 596 -702 656 -696
rect 1630 -702 1690 -696
rect 2132 -702 2192 194
rect 2432 -68 2492 194
rect 2432 -120 2436 -68
rect 2488 -120 2492 -68
rect 2556 920 2560 972
rect 2612 920 2616 972
rect 2556 -72 2616 920
rect 2432 -130 2492 -120
rect 2550 -76 2622 -72
rect 2550 -128 2560 -76
rect 2612 -128 2622 -76
rect 2550 -132 2622 -128
rect 596 -706 2192 -702
rect -2230 -756 -2170 -750
rect -1974 -756 -1914 -750
rect -1200 -756 -1140 -750
rect -942 -756 -882 -750
rect -2230 -760 -882 -756
rect -2230 -812 -2226 -760
rect -2174 -812 -1970 -760
rect -1918 -812 -1196 -760
rect -1144 -812 -938 -760
rect -886 -812 -882 -760
rect 596 -758 600 -706
rect 652 -758 1634 -706
rect 1686 -758 2192 -706
rect 596 -762 2192 -758
rect 596 -768 656 -762
rect 1630 -768 1690 -762
rect -2230 -816 -882 -812
rect -2230 -822 -2170 -816
rect -1974 -822 -1914 -816
rect -1200 -822 -1140 -816
rect -942 -822 -882 -816
rect -2362 -874 -2302 -868
rect -1846 -874 -1786 -868
rect -1326 -874 -1266 -868
rect -814 -874 -754 -868
rect -2852 -878 -754 -874
rect -2852 -930 -2358 -878
rect -2306 -930 -1842 -878
rect -1790 -930 -1322 -878
rect -1270 -930 -810 -878
rect -758 -930 -754 -878
rect -2852 -934 -754 -930
rect -2852 -1892 -2792 -934
rect -2362 -940 -2302 -934
rect -1846 -940 -1786 -934
rect -1326 -940 -1266 -934
rect -814 -940 -754 -934
rect 2132 -888 2192 -762
rect 2432 -888 2492 -882
rect 2132 -892 2492 -888
rect 2132 -944 2436 -892
rect 2488 -944 2492 -892
rect 2132 -948 2492 -944
rect 2432 -954 2492 -948
rect -2722 -1408 -2662 -1402
rect -1296 -1408 -1236 -1402
rect -428 -1408 -368 -1402
rect -2 -1408 58 -1402
rect 424 -1408 484 -1402
rect 1296 -1408 1356 -1402
rect -2722 -1412 2908 -1408
rect -2722 -1464 -2718 -1412
rect -2666 -1464 -1292 -1412
rect -1240 -1464 -424 -1412
rect -372 -1464 2 -1412
rect 54 -1464 428 -1412
rect 480 -1464 1300 -1412
rect 1352 -1464 2908 -1412
rect -2722 -1468 2908 -1464
rect -2722 -1474 -2662 -1468
rect -1296 -1474 -1236 -1468
rect -428 -1474 -368 -1468
rect -2 -1474 58 -1468
rect 424 -1474 484 -1468
rect 1296 -1474 1356 -1468
rect -2582 -1892 -2522 -1886
rect -2852 -1896 -2522 -1892
rect -2852 -1948 -2578 -1896
rect -2526 -1948 -2522 -1896
rect -2852 -1952 -2522 -1948
rect -2852 -2486 -2792 -1952
rect -2582 -1958 -2522 -1952
rect 2568 -1898 2628 -1892
rect 2848 -1898 2908 -1468
rect 2568 -1902 2908 -1898
rect 2568 -1954 2572 -1902
rect 2624 -1954 2908 -1902
rect 2568 -1958 2908 -1954
rect 2568 -1964 2628 -1958
rect -860 -2372 -800 -2366
rect 850 -2372 910 -2366
rect -860 -2376 910 -2372
rect -860 -2428 -856 -2376
rect -804 -2428 854 -2376
rect 906 -2428 910 -2376
rect -860 -2432 910 -2428
rect -860 -2438 -800 -2432
rect 850 -2438 910 -2432
rect -2 -2486 58 -2480
rect 2708 -2486 2768 -2480
rect -2852 -2490 2768 -2486
rect -2852 -2542 2 -2490
rect 54 -2542 2712 -2490
rect 2764 -2542 2768 -2490
rect -2852 -2546 2768 -2542
rect -2 -2552 58 -2546
rect 2708 -2552 2768 -2546
rect -928 -2891 970 -2836
rect -928 -2947 -886 -2891
rect -830 -2893 -806 -2891
rect -750 -2893 -726 -2891
rect -670 -2893 -646 -2891
rect -590 -2893 -566 -2891
rect -510 -2893 -486 -2891
rect -430 -2893 -406 -2891
rect -350 -2893 -326 -2891
rect -270 -2893 -246 -2891
rect -190 -2893 -166 -2891
rect -110 -2893 -86 -2891
rect -30 -2893 -6 -2891
rect 50 -2893 74 -2891
rect 130 -2893 154 -2891
rect 210 -2893 234 -2891
rect 290 -2893 314 -2891
rect 370 -2893 394 -2891
rect 450 -2893 474 -2891
rect 530 -2893 554 -2891
rect 610 -2893 634 -2891
rect 690 -2893 714 -2891
rect 770 -2893 794 -2891
rect 850 -2893 874 -2891
rect -816 -2945 -806 -2893
rect -750 -2945 -740 -2893
rect -496 -2945 -486 -2893
rect -430 -2945 -420 -2893
rect -176 -2945 -166 -2893
rect -110 -2945 -100 -2893
rect 144 -2945 154 -2893
rect 210 -2945 220 -2893
rect 464 -2945 474 -2893
rect 530 -2945 540 -2893
rect 784 -2945 794 -2893
rect 850 -2945 860 -2893
rect -830 -2947 -806 -2945
rect -750 -2947 -726 -2945
rect -670 -2947 -646 -2945
rect -590 -2947 -566 -2945
rect -510 -2947 -486 -2945
rect -430 -2947 -406 -2945
rect -350 -2947 -326 -2945
rect -270 -2947 -246 -2945
rect -190 -2947 -166 -2945
rect -110 -2947 -86 -2945
rect -30 -2947 -6 -2945
rect 50 -2947 74 -2945
rect 130 -2947 154 -2945
rect 210 -2947 234 -2945
rect 290 -2947 314 -2945
rect 370 -2947 394 -2945
rect 450 -2947 474 -2945
rect 530 -2947 554 -2945
rect 610 -2947 634 -2945
rect 690 -2947 714 -2945
rect 770 -2947 794 -2945
rect 850 -2947 874 -2945
rect 930 -2947 970 -2891
rect -928 -3002 970 -2947
rect -3216 -3118 -2616 -3106
rect -3216 -3144 -3184 -3118
rect -2648 -3144 -2616 -3118
rect -3216 -3388 -3198 -3144
rect -2634 -3388 -2616 -3144
rect -3216 -3414 -3184 -3388
rect -2648 -3414 -2616 -3388
rect -3216 -3426 -2616 -3414
rect 2616 -3118 3216 -3106
rect 2616 -3144 2648 -3118
rect 3184 -3144 3216 -3118
rect 2616 -3388 2634 -3144
rect 3198 -3388 3216 -3144
rect 2616 -3414 2648 -3388
rect 3184 -3414 3216 -3388
rect 2616 -3426 3216 -3414
<< via2 >>
rect -3184 2988 -2648 3014
rect -3184 2744 -2648 2988
rect -3184 2718 -2648 2744
rect 2648 2988 3184 3014
rect 2648 2744 3184 2988
rect 2648 2718 3184 2744
rect -2639 2518 -2583 2520
rect -2559 2518 -2503 2520
rect -2479 2518 -2423 2520
rect -2399 2518 -2343 2520
rect -2319 2518 -2263 2520
rect -2239 2518 -2183 2520
rect -2159 2518 -2103 2520
rect -2079 2518 -2023 2520
rect -1999 2518 -1943 2520
rect -1919 2518 -1863 2520
rect -1839 2518 -1783 2520
rect -1759 2518 -1703 2520
rect -1679 2518 -1623 2520
rect -1599 2518 -1543 2520
rect -1519 2518 -1463 2520
rect -1439 2518 -1383 2520
rect -1359 2518 -1303 2520
rect -1279 2518 -1223 2520
rect -1199 2518 -1143 2520
rect -1119 2518 -1063 2520
rect -1039 2518 -983 2520
rect -959 2518 -903 2520
rect -879 2518 -823 2520
rect -799 2518 -743 2520
rect -719 2518 -663 2520
rect -639 2518 -583 2520
rect -559 2518 -503 2520
rect -479 2518 -423 2520
rect -399 2518 -343 2520
rect -319 2518 -263 2520
rect -239 2518 -183 2520
rect -159 2518 -103 2520
rect -79 2518 -23 2520
rect 1 2518 57 2520
rect 81 2518 137 2520
rect 161 2518 217 2520
rect 241 2518 297 2520
rect 321 2518 377 2520
rect 401 2518 457 2520
rect 481 2518 537 2520
rect 561 2518 617 2520
rect 641 2518 697 2520
rect 721 2518 777 2520
rect 801 2518 857 2520
rect 881 2518 937 2520
rect 961 2518 1017 2520
rect 1041 2518 1097 2520
rect 1121 2518 1177 2520
rect 1201 2518 1257 2520
rect 1281 2518 1337 2520
rect 1361 2518 1417 2520
rect 1441 2518 1497 2520
rect 1521 2518 1577 2520
rect 1601 2518 1657 2520
rect 1681 2518 1737 2520
rect 1761 2518 1817 2520
rect 1841 2518 1897 2520
rect 1921 2518 1977 2520
rect 2001 2518 2057 2520
rect 2081 2518 2137 2520
rect 2161 2518 2217 2520
rect 2241 2518 2297 2520
rect 2321 2518 2377 2520
rect 2401 2518 2457 2520
rect 2481 2518 2537 2520
rect -2639 2466 -2637 2518
rect -2637 2466 -2585 2518
rect -2585 2466 -2583 2518
rect -2559 2466 -2521 2518
rect -2521 2466 -2509 2518
rect -2509 2466 -2503 2518
rect -2479 2466 -2457 2518
rect -2457 2466 -2445 2518
rect -2445 2466 -2423 2518
rect -2399 2466 -2393 2518
rect -2393 2466 -2381 2518
rect -2381 2466 -2343 2518
rect -2319 2466 -2317 2518
rect -2317 2466 -2265 2518
rect -2265 2466 -2263 2518
rect -2239 2466 -2201 2518
rect -2201 2466 -2189 2518
rect -2189 2466 -2183 2518
rect -2159 2466 -2137 2518
rect -2137 2466 -2125 2518
rect -2125 2466 -2103 2518
rect -2079 2466 -2073 2518
rect -2073 2466 -2061 2518
rect -2061 2466 -2023 2518
rect -1999 2466 -1997 2518
rect -1997 2466 -1945 2518
rect -1945 2466 -1943 2518
rect -1919 2466 -1881 2518
rect -1881 2466 -1869 2518
rect -1869 2466 -1863 2518
rect -1839 2466 -1817 2518
rect -1817 2466 -1805 2518
rect -1805 2466 -1783 2518
rect -1759 2466 -1753 2518
rect -1753 2466 -1741 2518
rect -1741 2466 -1703 2518
rect -1679 2466 -1677 2518
rect -1677 2466 -1625 2518
rect -1625 2466 -1623 2518
rect -1599 2466 -1561 2518
rect -1561 2466 -1549 2518
rect -1549 2466 -1543 2518
rect -1519 2466 -1497 2518
rect -1497 2466 -1485 2518
rect -1485 2466 -1463 2518
rect -1439 2466 -1433 2518
rect -1433 2466 -1421 2518
rect -1421 2466 -1383 2518
rect -1359 2466 -1357 2518
rect -1357 2466 -1305 2518
rect -1305 2466 -1303 2518
rect -1279 2466 -1241 2518
rect -1241 2466 -1229 2518
rect -1229 2466 -1223 2518
rect -1199 2466 -1177 2518
rect -1177 2466 -1165 2518
rect -1165 2466 -1143 2518
rect -1119 2466 -1113 2518
rect -1113 2466 -1101 2518
rect -1101 2466 -1063 2518
rect -1039 2466 -1037 2518
rect -1037 2466 -985 2518
rect -985 2466 -983 2518
rect -959 2466 -921 2518
rect -921 2466 -909 2518
rect -909 2466 -903 2518
rect -879 2466 -857 2518
rect -857 2466 -845 2518
rect -845 2466 -823 2518
rect -799 2466 -793 2518
rect -793 2466 -781 2518
rect -781 2466 -743 2518
rect -719 2466 -717 2518
rect -717 2466 -665 2518
rect -665 2466 -663 2518
rect -639 2466 -601 2518
rect -601 2466 -589 2518
rect -589 2466 -583 2518
rect -559 2466 -537 2518
rect -537 2466 -525 2518
rect -525 2466 -503 2518
rect -479 2466 -473 2518
rect -473 2466 -461 2518
rect -461 2466 -423 2518
rect -399 2466 -397 2518
rect -397 2466 -345 2518
rect -345 2466 -343 2518
rect -319 2466 -281 2518
rect -281 2466 -269 2518
rect -269 2466 -263 2518
rect -239 2466 -217 2518
rect -217 2466 -205 2518
rect -205 2466 -183 2518
rect -159 2466 -153 2518
rect -153 2466 -141 2518
rect -141 2466 -103 2518
rect -79 2466 -77 2518
rect -77 2466 -25 2518
rect -25 2466 -23 2518
rect 1 2466 39 2518
rect 39 2466 51 2518
rect 51 2466 57 2518
rect 81 2466 103 2518
rect 103 2466 115 2518
rect 115 2466 137 2518
rect 161 2466 167 2518
rect 167 2466 179 2518
rect 179 2466 217 2518
rect 241 2466 243 2518
rect 243 2466 295 2518
rect 295 2466 297 2518
rect 321 2466 359 2518
rect 359 2466 371 2518
rect 371 2466 377 2518
rect 401 2466 423 2518
rect 423 2466 435 2518
rect 435 2466 457 2518
rect 481 2466 487 2518
rect 487 2466 499 2518
rect 499 2466 537 2518
rect 561 2466 563 2518
rect 563 2466 615 2518
rect 615 2466 617 2518
rect 641 2466 679 2518
rect 679 2466 691 2518
rect 691 2466 697 2518
rect 721 2466 743 2518
rect 743 2466 755 2518
rect 755 2466 777 2518
rect 801 2466 807 2518
rect 807 2466 819 2518
rect 819 2466 857 2518
rect 881 2466 883 2518
rect 883 2466 935 2518
rect 935 2466 937 2518
rect 961 2466 999 2518
rect 999 2466 1011 2518
rect 1011 2466 1017 2518
rect 1041 2466 1063 2518
rect 1063 2466 1075 2518
rect 1075 2466 1097 2518
rect 1121 2466 1127 2518
rect 1127 2466 1139 2518
rect 1139 2466 1177 2518
rect 1201 2466 1203 2518
rect 1203 2466 1255 2518
rect 1255 2466 1257 2518
rect 1281 2466 1319 2518
rect 1319 2466 1331 2518
rect 1331 2466 1337 2518
rect 1361 2466 1383 2518
rect 1383 2466 1395 2518
rect 1395 2466 1417 2518
rect 1441 2466 1447 2518
rect 1447 2466 1459 2518
rect 1459 2466 1497 2518
rect 1521 2466 1523 2518
rect 1523 2466 1575 2518
rect 1575 2466 1577 2518
rect 1601 2466 1639 2518
rect 1639 2466 1651 2518
rect 1651 2466 1657 2518
rect 1681 2466 1703 2518
rect 1703 2466 1715 2518
rect 1715 2466 1737 2518
rect 1761 2466 1767 2518
rect 1767 2466 1779 2518
rect 1779 2466 1817 2518
rect 1841 2466 1843 2518
rect 1843 2466 1895 2518
rect 1895 2466 1897 2518
rect 1921 2466 1959 2518
rect 1959 2466 1971 2518
rect 1971 2466 1977 2518
rect 2001 2466 2023 2518
rect 2023 2466 2035 2518
rect 2035 2466 2057 2518
rect 2081 2466 2087 2518
rect 2087 2466 2099 2518
rect 2099 2466 2137 2518
rect 2161 2466 2163 2518
rect 2163 2466 2215 2518
rect 2215 2466 2217 2518
rect 2241 2466 2279 2518
rect 2279 2466 2291 2518
rect 2291 2466 2297 2518
rect 2321 2466 2343 2518
rect 2343 2466 2355 2518
rect 2355 2466 2377 2518
rect 2401 2466 2407 2518
rect 2407 2466 2419 2518
rect 2419 2466 2457 2518
rect 2481 2466 2483 2518
rect 2483 2466 2535 2518
rect 2535 2466 2537 2518
rect -2639 2464 -2583 2466
rect -2559 2464 -2503 2466
rect -2479 2464 -2423 2466
rect -2399 2464 -2343 2466
rect -2319 2464 -2263 2466
rect -2239 2464 -2183 2466
rect -2159 2464 -2103 2466
rect -2079 2464 -2023 2466
rect -1999 2464 -1943 2466
rect -1919 2464 -1863 2466
rect -1839 2464 -1783 2466
rect -1759 2464 -1703 2466
rect -1679 2464 -1623 2466
rect -1599 2464 -1543 2466
rect -1519 2464 -1463 2466
rect -1439 2464 -1383 2466
rect -1359 2464 -1303 2466
rect -1279 2464 -1223 2466
rect -1199 2464 -1143 2466
rect -1119 2464 -1063 2466
rect -1039 2464 -983 2466
rect -959 2464 -903 2466
rect -879 2464 -823 2466
rect -799 2464 -743 2466
rect -719 2464 -663 2466
rect -639 2464 -583 2466
rect -559 2464 -503 2466
rect -479 2464 -423 2466
rect -399 2464 -343 2466
rect -319 2464 -263 2466
rect -239 2464 -183 2466
rect -159 2464 -103 2466
rect -79 2464 -23 2466
rect 1 2464 57 2466
rect 81 2464 137 2466
rect 161 2464 217 2466
rect 241 2464 297 2466
rect 321 2464 377 2466
rect 401 2464 457 2466
rect 481 2464 537 2466
rect 561 2464 617 2466
rect 641 2464 697 2466
rect 721 2464 777 2466
rect 801 2464 857 2466
rect 881 2464 937 2466
rect 961 2464 1017 2466
rect 1041 2464 1097 2466
rect 1121 2464 1177 2466
rect 1201 2464 1257 2466
rect 1281 2464 1337 2466
rect 1361 2464 1417 2466
rect 1441 2464 1497 2466
rect 1521 2464 1577 2466
rect 1601 2464 1657 2466
rect 1681 2464 1737 2466
rect 1761 2464 1817 2466
rect 1841 2464 1897 2466
rect 1921 2464 1977 2466
rect 2001 2464 2057 2466
rect 2081 2464 2137 2466
rect 2161 2464 2217 2466
rect 2241 2464 2297 2466
rect 2321 2464 2377 2466
rect 2401 2464 2457 2466
rect 2481 2464 2537 2466
rect -886 -2893 -830 -2891
rect -806 -2893 -750 -2891
rect -726 -2893 -670 -2891
rect -646 -2893 -590 -2891
rect -566 -2893 -510 -2891
rect -486 -2893 -430 -2891
rect -406 -2893 -350 -2891
rect -326 -2893 -270 -2891
rect -246 -2893 -190 -2891
rect -166 -2893 -110 -2891
rect -86 -2893 -30 -2891
rect -6 -2893 50 -2891
rect 74 -2893 130 -2891
rect 154 -2893 210 -2891
rect 234 -2893 290 -2891
rect 314 -2893 370 -2891
rect 394 -2893 450 -2891
rect 474 -2893 530 -2891
rect 554 -2893 610 -2891
rect 634 -2893 690 -2891
rect 714 -2893 770 -2891
rect 794 -2893 850 -2891
rect 874 -2893 930 -2891
rect -886 -2945 -868 -2893
rect -868 -2945 -830 -2893
rect -806 -2945 -804 -2893
rect -804 -2945 -752 -2893
rect -752 -2945 -750 -2893
rect -726 -2945 -688 -2893
rect -688 -2945 -676 -2893
rect -676 -2945 -670 -2893
rect -646 -2945 -624 -2893
rect -624 -2945 -612 -2893
rect -612 -2945 -590 -2893
rect -566 -2945 -560 -2893
rect -560 -2945 -548 -2893
rect -548 -2945 -510 -2893
rect -486 -2945 -484 -2893
rect -484 -2945 -432 -2893
rect -432 -2945 -430 -2893
rect -406 -2945 -368 -2893
rect -368 -2945 -356 -2893
rect -356 -2945 -350 -2893
rect -326 -2945 -304 -2893
rect -304 -2945 -292 -2893
rect -292 -2945 -270 -2893
rect -246 -2945 -240 -2893
rect -240 -2945 -228 -2893
rect -228 -2945 -190 -2893
rect -166 -2945 -164 -2893
rect -164 -2945 -112 -2893
rect -112 -2945 -110 -2893
rect -86 -2945 -48 -2893
rect -48 -2945 -36 -2893
rect -36 -2945 -30 -2893
rect -6 -2945 16 -2893
rect 16 -2945 28 -2893
rect 28 -2945 50 -2893
rect 74 -2945 80 -2893
rect 80 -2945 92 -2893
rect 92 -2945 130 -2893
rect 154 -2945 156 -2893
rect 156 -2945 208 -2893
rect 208 -2945 210 -2893
rect 234 -2945 272 -2893
rect 272 -2945 284 -2893
rect 284 -2945 290 -2893
rect 314 -2945 336 -2893
rect 336 -2945 348 -2893
rect 348 -2945 370 -2893
rect 394 -2945 400 -2893
rect 400 -2945 412 -2893
rect 412 -2945 450 -2893
rect 474 -2945 476 -2893
rect 476 -2945 528 -2893
rect 528 -2945 530 -2893
rect 554 -2945 592 -2893
rect 592 -2945 604 -2893
rect 604 -2945 610 -2893
rect 634 -2945 656 -2893
rect 656 -2945 668 -2893
rect 668 -2945 690 -2893
rect 714 -2945 720 -2893
rect 720 -2945 732 -2893
rect 732 -2945 770 -2893
rect 794 -2945 796 -2893
rect 796 -2945 848 -2893
rect 848 -2945 850 -2893
rect 874 -2945 912 -2893
rect 912 -2945 930 -2893
rect -886 -2947 -830 -2945
rect -806 -2947 -750 -2945
rect -726 -2947 -670 -2945
rect -646 -2947 -590 -2945
rect -566 -2947 -510 -2945
rect -486 -2947 -430 -2945
rect -406 -2947 -350 -2945
rect -326 -2947 -270 -2945
rect -246 -2947 -190 -2945
rect -166 -2947 -110 -2945
rect -86 -2947 -30 -2945
rect -6 -2947 50 -2945
rect 74 -2947 130 -2945
rect 154 -2947 210 -2945
rect 234 -2947 290 -2945
rect 314 -2947 370 -2945
rect 394 -2947 450 -2945
rect 474 -2947 530 -2945
rect 554 -2947 610 -2945
rect 634 -2947 690 -2945
rect 714 -2947 770 -2945
rect 794 -2947 850 -2945
rect 874 -2947 930 -2945
rect -3184 -3144 -2648 -3118
rect -3184 -3388 -2648 -3144
rect -3184 -3414 -2648 -3388
rect 2648 -3144 3184 -3118
rect 2648 -3388 3184 -3144
rect 2648 -3414 3184 -3388
<< metal3 >>
rect -3226 3014 -2606 3021
rect -3226 2978 -3184 3014
rect -2648 2978 -2606 3014
rect -3226 2754 -3188 2978
rect -2644 2754 -2606 2978
rect -3226 2718 -3184 2754
rect -2648 2718 -2606 2754
rect -3226 2711 -2606 2718
rect 2606 3014 3226 3021
rect 2606 2978 2648 3014
rect 3184 2978 3226 3014
rect 2606 2754 2644 2978
rect 3188 2754 3226 2978
rect 2606 2718 2648 2754
rect 3184 2718 3226 2754
rect 2606 2711 3226 2718
rect -2674 2524 2566 2562
rect -2674 2460 -2643 2524
rect -2579 2460 -2563 2524
rect -2499 2460 -2483 2524
rect -2419 2460 -2403 2524
rect -2339 2460 -2323 2524
rect -2259 2460 -2243 2524
rect -2179 2460 -2163 2524
rect -2099 2460 -2083 2524
rect -2019 2460 -2003 2524
rect -1939 2460 -1923 2524
rect -1859 2460 -1843 2524
rect -1779 2460 -1763 2524
rect -1699 2460 -1683 2524
rect -1619 2460 -1603 2524
rect -1539 2460 -1523 2524
rect -1459 2460 -1443 2524
rect -1379 2460 -1363 2524
rect -1299 2460 -1283 2524
rect -1219 2460 -1203 2524
rect -1139 2460 -1123 2524
rect -1059 2460 -1043 2524
rect -979 2460 -963 2524
rect -899 2460 -883 2524
rect -819 2460 -803 2524
rect -739 2460 -723 2524
rect -659 2460 -643 2524
rect -579 2460 -563 2524
rect -499 2460 -483 2524
rect -419 2460 -403 2524
rect -339 2460 -323 2524
rect -259 2460 -243 2524
rect -179 2460 -163 2524
rect -99 2460 -83 2524
rect -19 2460 -3 2524
rect 61 2460 77 2524
rect 141 2460 157 2524
rect 221 2460 237 2524
rect 301 2460 317 2524
rect 381 2460 397 2524
rect 461 2460 477 2524
rect 541 2460 557 2524
rect 621 2460 637 2524
rect 701 2460 717 2524
rect 781 2460 797 2524
rect 861 2460 877 2524
rect 941 2460 957 2524
rect 1021 2460 1037 2524
rect 1101 2460 1117 2524
rect 1181 2460 1197 2524
rect 1261 2460 1277 2524
rect 1341 2460 1357 2524
rect 1421 2460 1437 2524
rect 1501 2460 1517 2524
rect 1581 2460 1597 2524
rect 1661 2460 1677 2524
rect 1741 2460 1757 2524
rect 1821 2460 1837 2524
rect 1901 2460 1917 2524
rect 1981 2460 1997 2524
rect 2061 2460 2077 2524
rect 2141 2460 2157 2524
rect 2221 2460 2237 2524
rect 2301 2460 2317 2524
rect 2381 2460 2397 2524
rect 2461 2460 2477 2524
rect 2541 2460 2566 2524
rect -2674 2430 2566 2460
rect -928 -2887 970 -2836
rect -928 -2951 -890 -2887
rect -826 -2951 -810 -2887
rect -746 -2951 -730 -2887
rect -666 -2951 -650 -2887
rect -586 -2951 -570 -2887
rect -506 -2951 -490 -2887
rect -426 -2951 -410 -2887
rect -346 -2951 -330 -2887
rect -266 -2951 -250 -2887
rect -186 -2951 -170 -2887
rect -106 -2951 -90 -2887
rect -26 -2951 -10 -2887
rect 54 -2951 70 -2887
rect 134 -2951 150 -2887
rect 214 -2951 230 -2887
rect 294 -2951 310 -2887
rect 374 -2951 390 -2887
rect 454 -2951 470 -2887
rect 534 -2951 550 -2887
rect 614 -2951 630 -2887
rect 694 -2951 710 -2887
rect 774 -2951 790 -2887
rect 854 -2951 870 -2887
rect 934 -2951 970 -2887
rect -928 -3002 970 -2951
rect -3226 -3118 -2606 -3111
rect -3226 -3154 -3184 -3118
rect -2648 -3154 -2606 -3118
rect -3226 -3378 -3188 -3154
rect -2644 -3378 -2606 -3154
rect -3226 -3414 -3184 -3378
rect -2648 -3414 -2606 -3378
rect -3226 -3421 -2606 -3414
rect 2606 -3118 3226 -3111
rect 2606 -3154 2648 -3118
rect 3184 -3154 3226 -3118
rect 2606 -3378 2644 -3154
rect 3188 -3378 3226 -3154
rect 2606 -3414 2648 -3378
rect 3184 -3414 3226 -3378
rect 2606 -3421 3226 -3414
<< via3 >>
rect -3188 2754 -3184 2978
rect -3184 2754 -2648 2978
rect -2648 2754 -2644 2978
rect 2644 2754 2648 2978
rect 2648 2754 3184 2978
rect 3184 2754 3188 2978
rect -2643 2520 -2579 2524
rect -2643 2464 -2639 2520
rect -2639 2464 -2583 2520
rect -2583 2464 -2579 2520
rect -2643 2460 -2579 2464
rect -2563 2520 -2499 2524
rect -2563 2464 -2559 2520
rect -2559 2464 -2503 2520
rect -2503 2464 -2499 2520
rect -2563 2460 -2499 2464
rect -2483 2520 -2419 2524
rect -2483 2464 -2479 2520
rect -2479 2464 -2423 2520
rect -2423 2464 -2419 2520
rect -2483 2460 -2419 2464
rect -2403 2520 -2339 2524
rect -2403 2464 -2399 2520
rect -2399 2464 -2343 2520
rect -2343 2464 -2339 2520
rect -2403 2460 -2339 2464
rect -2323 2520 -2259 2524
rect -2323 2464 -2319 2520
rect -2319 2464 -2263 2520
rect -2263 2464 -2259 2520
rect -2323 2460 -2259 2464
rect -2243 2520 -2179 2524
rect -2243 2464 -2239 2520
rect -2239 2464 -2183 2520
rect -2183 2464 -2179 2520
rect -2243 2460 -2179 2464
rect -2163 2520 -2099 2524
rect -2163 2464 -2159 2520
rect -2159 2464 -2103 2520
rect -2103 2464 -2099 2520
rect -2163 2460 -2099 2464
rect -2083 2520 -2019 2524
rect -2083 2464 -2079 2520
rect -2079 2464 -2023 2520
rect -2023 2464 -2019 2520
rect -2083 2460 -2019 2464
rect -2003 2520 -1939 2524
rect -2003 2464 -1999 2520
rect -1999 2464 -1943 2520
rect -1943 2464 -1939 2520
rect -2003 2460 -1939 2464
rect -1923 2520 -1859 2524
rect -1923 2464 -1919 2520
rect -1919 2464 -1863 2520
rect -1863 2464 -1859 2520
rect -1923 2460 -1859 2464
rect -1843 2520 -1779 2524
rect -1843 2464 -1839 2520
rect -1839 2464 -1783 2520
rect -1783 2464 -1779 2520
rect -1843 2460 -1779 2464
rect -1763 2520 -1699 2524
rect -1763 2464 -1759 2520
rect -1759 2464 -1703 2520
rect -1703 2464 -1699 2520
rect -1763 2460 -1699 2464
rect -1683 2520 -1619 2524
rect -1683 2464 -1679 2520
rect -1679 2464 -1623 2520
rect -1623 2464 -1619 2520
rect -1683 2460 -1619 2464
rect -1603 2520 -1539 2524
rect -1603 2464 -1599 2520
rect -1599 2464 -1543 2520
rect -1543 2464 -1539 2520
rect -1603 2460 -1539 2464
rect -1523 2520 -1459 2524
rect -1523 2464 -1519 2520
rect -1519 2464 -1463 2520
rect -1463 2464 -1459 2520
rect -1523 2460 -1459 2464
rect -1443 2520 -1379 2524
rect -1443 2464 -1439 2520
rect -1439 2464 -1383 2520
rect -1383 2464 -1379 2520
rect -1443 2460 -1379 2464
rect -1363 2520 -1299 2524
rect -1363 2464 -1359 2520
rect -1359 2464 -1303 2520
rect -1303 2464 -1299 2520
rect -1363 2460 -1299 2464
rect -1283 2520 -1219 2524
rect -1283 2464 -1279 2520
rect -1279 2464 -1223 2520
rect -1223 2464 -1219 2520
rect -1283 2460 -1219 2464
rect -1203 2520 -1139 2524
rect -1203 2464 -1199 2520
rect -1199 2464 -1143 2520
rect -1143 2464 -1139 2520
rect -1203 2460 -1139 2464
rect -1123 2520 -1059 2524
rect -1123 2464 -1119 2520
rect -1119 2464 -1063 2520
rect -1063 2464 -1059 2520
rect -1123 2460 -1059 2464
rect -1043 2520 -979 2524
rect -1043 2464 -1039 2520
rect -1039 2464 -983 2520
rect -983 2464 -979 2520
rect -1043 2460 -979 2464
rect -963 2520 -899 2524
rect -963 2464 -959 2520
rect -959 2464 -903 2520
rect -903 2464 -899 2520
rect -963 2460 -899 2464
rect -883 2520 -819 2524
rect -883 2464 -879 2520
rect -879 2464 -823 2520
rect -823 2464 -819 2520
rect -883 2460 -819 2464
rect -803 2520 -739 2524
rect -803 2464 -799 2520
rect -799 2464 -743 2520
rect -743 2464 -739 2520
rect -803 2460 -739 2464
rect -723 2520 -659 2524
rect -723 2464 -719 2520
rect -719 2464 -663 2520
rect -663 2464 -659 2520
rect -723 2460 -659 2464
rect -643 2520 -579 2524
rect -643 2464 -639 2520
rect -639 2464 -583 2520
rect -583 2464 -579 2520
rect -643 2460 -579 2464
rect -563 2520 -499 2524
rect -563 2464 -559 2520
rect -559 2464 -503 2520
rect -503 2464 -499 2520
rect -563 2460 -499 2464
rect -483 2520 -419 2524
rect -483 2464 -479 2520
rect -479 2464 -423 2520
rect -423 2464 -419 2520
rect -483 2460 -419 2464
rect -403 2520 -339 2524
rect -403 2464 -399 2520
rect -399 2464 -343 2520
rect -343 2464 -339 2520
rect -403 2460 -339 2464
rect -323 2520 -259 2524
rect -323 2464 -319 2520
rect -319 2464 -263 2520
rect -263 2464 -259 2520
rect -323 2460 -259 2464
rect -243 2520 -179 2524
rect -243 2464 -239 2520
rect -239 2464 -183 2520
rect -183 2464 -179 2520
rect -243 2460 -179 2464
rect -163 2520 -99 2524
rect -163 2464 -159 2520
rect -159 2464 -103 2520
rect -103 2464 -99 2520
rect -163 2460 -99 2464
rect -83 2520 -19 2524
rect -83 2464 -79 2520
rect -79 2464 -23 2520
rect -23 2464 -19 2520
rect -83 2460 -19 2464
rect -3 2520 61 2524
rect -3 2464 1 2520
rect 1 2464 57 2520
rect 57 2464 61 2520
rect -3 2460 61 2464
rect 77 2520 141 2524
rect 77 2464 81 2520
rect 81 2464 137 2520
rect 137 2464 141 2520
rect 77 2460 141 2464
rect 157 2520 221 2524
rect 157 2464 161 2520
rect 161 2464 217 2520
rect 217 2464 221 2520
rect 157 2460 221 2464
rect 237 2520 301 2524
rect 237 2464 241 2520
rect 241 2464 297 2520
rect 297 2464 301 2520
rect 237 2460 301 2464
rect 317 2520 381 2524
rect 317 2464 321 2520
rect 321 2464 377 2520
rect 377 2464 381 2520
rect 317 2460 381 2464
rect 397 2520 461 2524
rect 397 2464 401 2520
rect 401 2464 457 2520
rect 457 2464 461 2520
rect 397 2460 461 2464
rect 477 2520 541 2524
rect 477 2464 481 2520
rect 481 2464 537 2520
rect 537 2464 541 2520
rect 477 2460 541 2464
rect 557 2520 621 2524
rect 557 2464 561 2520
rect 561 2464 617 2520
rect 617 2464 621 2520
rect 557 2460 621 2464
rect 637 2520 701 2524
rect 637 2464 641 2520
rect 641 2464 697 2520
rect 697 2464 701 2520
rect 637 2460 701 2464
rect 717 2520 781 2524
rect 717 2464 721 2520
rect 721 2464 777 2520
rect 777 2464 781 2520
rect 717 2460 781 2464
rect 797 2520 861 2524
rect 797 2464 801 2520
rect 801 2464 857 2520
rect 857 2464 861 2520
rect 797 2460 861 2464
rect 877 2520 941 2524
rect 877 2464 881 2520
rect 881 2464 937 2520
rect 937 2464 941 2520
rect 877 2460 941 2464
rect 957 2520 1021 2524
rect 957 2464 961 2520
rect 961 2464 1017 2520
rect 1017 2464 1021 2520
rect 957 2460 1021 2464
rect 1037 2520 1101 2524
rect 1037 2464 1041 2520
rect 1041 2464 1097 2520
rect 1097 2464 1101 2520
rect 1037 2460 1101 2464
rect 1117 2520 1181 2524
rect 1117 2464 1121 2520
rect 1121 2464 1177 2520
rect 1177 2464 1181 2520
rect 1117 2460 1181 2464
rect 1197 2520 1261 2524
rect 1197 2464 1201 2520
rect 1201 2464 1257 2520
rect 1257 2464 1261 2520
rect 1197 2460 1261 2464
rect 1277 2520 1341 2524
rect 1277 2464 1281 2520
rect 1281 2464 1337 2520
rect 1337 2464 1341 2520
rect 1277 2460 1341 2464
rect 1357 2520 1421 2524
rect 1357 2464 1361 2520
rect 1361 2464 1417 2520
rect 1417 2464 1421 2520
rect 1357 2460 1421 2464
rect 1437 2520 1501 2524
rect 1437 2464 1441 2520
rect 1441 2464 1497 2520
rect 1497 2464 1501 2520
rect 1437 2460 1501 2464
rect 1517 2520 1581 2524
rect 1517 2464 1521 2520
rect 1521 2464 1577 2520
rect 1577 2464 1581 2520
rect 1517 2460 1581 2464
rect 1597 2520 1661 2524
rect 1597 2464 1601 2520
rect 1601 2464 1657 2520
rect 1657 2464 1661 2520
rect 1597 2460 1661 2464
rect 1677 2520 1741 2524
rect 1677 2464 1681 2520
rect 1681 2464 1737 2520
rect 1737 2464 1741 2520
rect 1677 2460 1741 2464
rect 1757 2520 1821 2524
rect 1757 2464 1761 2520
rect 1761 2464 1817 2520
rect 1817 2464 1821 2520
rect 1757 2460 1821 2464
rect 1837 2520 1901 2524
rect 1837 2464 1841 2520
rect 1841 2464 1897 2520
rect 1897 2464 1901 2520
rect 1837 2460 1901 2464
rect 1917 2520 1981 2524
rect 1917 2464 1921 2520
rect 1921 2464 1977 2520
rect 1977 2464 1981 2520
rect 1917 2460 1981 2464
rect 1997 2520 2061 2524
rect 1997 2464 2001 2520
rect 2001 2464 2057 2520
rect 2057 2464 2061 2520
rect 1997 2460 2061 2464
rect 2077 2520 2141 2524
rect 2077 2464 2081 2520
rect 2081 2464 2137 2520
rect 2137 2464 2141 2520
rect 2077 2460 2141 2464
rect 2157 2520 2221 2524
rect 2157 2464 2161 2520
rect 2161 2464 2217 2520
rect 2217 2464 2221 2520
rect 2157 2460 2221 2464
rect 2237 2520 2301 2524
rect 2237 2464 2241 2520
rect 2241 2464 2297 2520
rect 2297 2464 2301 2520
rect 2237 2460 2301 2464
rect 2317 2520 2381 2524
rect 2317 2464 2321 2520
rect 2321 2464 2377 2520
rect 2377 2464 2381 2520
rect 2317 2460 2381 2464
rect 2397 2520 2461 2524
rect 2397 2464 2401 2520
rect 2401 2464 2457 2520
rect 2457 2464 2461 2520
rect 2397 2460 2461 2464
rect 2477 2520 2541 2524
rect 2477 2464 2481 2520
rect 2481 2464 2537 2520
rect 2537 2464 2541 2520
rect 2477 2460 2541 2464
rect -890 -2891 -826 -2887
rect -890 -2947 -886 -2891
rect -886 -2947 -830 -2891
rect -830 -2947 -826 -2891
rect -890 -2951 -826 -2947
rect -810 -2891 -746 -2887
rect -810 -2947 -806 -2891
rect -806 -2947 -750 -2891
rect -750 -2947 -746 -2891
rect -810 -2951 -746 -2947
rect -730 -2891 -666 -2887
rect -730 -2947 -726 -2891
rect -726 -2947 -670 -2891
rect -670 -2947 -666 -2891
rect -730 -2951 -666 -2947
rect -650 -2891 -586 -2887
rect -650 -2947 -646 -2891
rect -646 -2947 -590 -2891
rect -590 -2947 -586 -2891
rect -650 -2951 -586 -2947
rect -570 -2891 -506 -2887
rect -570 -2947 -566 -2891
rect -566 -2947 -510 -2891
rect -510 -2947 -506 -2891
rect -570 -2951 -506 -2947
rect -490 -2891 -426 -2887
rect -490 -2947 -486 -2891
rect -486 -2947 -430 -2891
rect -430 -2947 -426 -2891
rect -490 -2951 -426 -2947
rect -410 -2891 -346 -2887
rect -410 -2947 -406 -2891
rect -406 -2947 -350 -2891
rect -350 -2947 -346 -2891
rect -410 -2951 -346 -2947
rect -330 -2891 -266 -2887
rect -330 -2947 -326 -2891
rect -326 -2947 -270 -2891
rect -270 -2947 -266 -2891
rect -330 -2951 -266 -2947
rect -250 -2891 -186 -2887
rect -250 -2947 -246 -2891
rect -246 -2947 -190 -2891
rect -190 -2947 -186 -2891
rect -250 -2951 -186 -2947
rect -170 -2891 -106 -2887
rect -170 -2947 -166 -2891
rect -166 -2947 -110 -2891
rect -110 -2947 -106 -2891
rect -170 -2951 -106 -2947
rect -90 -2891 -26 -2887
rect -90 -2947 -86 -2891
rect -86 -2947 -30 -2891
rect -30 -2947 -26 -2891
rect -90 -2951 -26 -2947
rect -10 -2891 54 -2887
rect -10 -2947 -6 -2891
rect -6 -2947 50 -2891
rect 50 -2947 54 -2891
rect -10 -2951 54 -2947
rect 70 -2891 134 -2887
rect 70 -2947 74 -2891
rect 74 -2947 130 -2891
rect 130 -2947 134 -2891
rect 70 -2951 134 -2947
rect 150 -2891 214 -2887
rect 150 -2947 154 -2891
rect 154 -2947 210 -2891
rect 210 -2947 214 -2891
rect 150 -2951 214 -2947
rect 230 -2891 294 -2887
rect 230 -2947 234 -2891
rect 234 -2947 290 -2891
rect 290 -2947 294 -2891
rect 230 -2951 294 -2947
rect 310 -2891 374 -2887
rect 310 -2947 314 -2891
rect 314 -2947 370 -2891
rect 370 -2947 374 -2891
rect 310 -2951 374 -2947
rect 390 -2891 454 -2887
rect 390 -2947 394 -2891
rect 394 -2947 450 -2891
rect 450 -2947 454 -2891
rect 390 -2951 454 -2947
rect 470 -2891 534 -2887
rect 470 -2947 474 -2891
rect 474 -2947 530 -2891
rect 530 -2947 534 -2891
rect 470 -2951 534 -2947
rect 550 -2891 614 -2887
rect 550 -2947 554 -2891
rect 554 -2947 610 -2891
rect 610 -2947 614 -2891
rect 550 -2951 614 -2947
rect 630 -2891 694 -2887
rect 630 -2947 634 -2891
rect 634 -2947 690 -2891
rect 690 -2947 694 -2891
rect 630 -2951 694 -2947
rect 710 -2891 774 -2887
rect 710 -2947 714 -2891
rect 714 -2947 770 -2891
rect 770 -2947 774 -2891
rect 710 -2951 774 -2947
rect 790 -2891 854 -2887
rect 790 -2947 794 -2891
rect 794 -2947 850 -2891
rect 850 -2947 854 -2891
rect 790 -2951 854 -2947
rect 870 -2891 934 -2887
rect 870 -2947 874 -2891
rect 874 -2947 930 -2891
rect 930 -2947 934 -2891
rect 870 -2951 934 -2947
rect -3188 -3378 -3184 -3154
rect -3184 -3378 -2648 -3154
rect -2648 -3378 -2644 -3154
rect 2644 -3378 2648 -3154
rect 2648 -3378 3184 -3154
rect 3184 -3378 3188 -3154
<< metal4 >>
rect -3400 2978 3400 3200
rect -3400 2754 -3188 2978
rect -2644 2754 2644 2978
rect 3188 2754 3400 2978
rect -3400 2524 3400 2754
rect -3400 2460 -2643 2524
rect -2579 2460 -2563 2524
rect -2499 2460 -2483 2524
rect -2419 2460 -2403 2524
rect -2339 2460 -2323 2524
rect -2259 2460 -2243 2524
rect -2179 2460 -2163 2524
rect -2099 2460 -2083 2524
rect -2019 2460 -2003 2524
rect -1939 2460 -1923 2524
rect -1859 2460 -1843 2524
rect -1779 2460 -1763 2524
rect -1699 2460 -1683 2524
rect -1619 2460 -1603 2524
rect -1539 2460 -1523 2524
rect -1459 2460 -1443 2524
rect -1379 2460 -1363 2524
rect -1299 2460 -1283 2524
rect -1219 2460 -1203 2524
rect -1139 2460 -1123 2524
rect -1059 2460 -1043 2524
rect -979 2460 -963 2524
rect -899 2460 -883 2524
rect -819 2460 -803 2524
rect -739 2460 -723 2524
rect -659 2460 -643 2524
rect -579 2460 -563 2524
rect -499 2460 -483 2524
rect -419 2460 -403 2524
rect -339 2460 -323 2524
rect -259 2460 -243 2524
rect -179 2460 -163 2524
rect -99 2460 -83 2524
rect -19 2460 -3 2524
rect 61 2460 77 2524
rect 141 2460 157 2524
rect 221 2460 237 2524
rect 301 2460 317 2524
rect 381 2460 397 2524
rect 461 2460 477 2524
rect 541 2460 557 2524
rect 621 2460 637 2524
rect 701 2460 717 2524
rect 781 2460 797 2524
rect 861 2460 877 2524
rect 941 2460 957 2524
rect 1021 2460 1037 2524
rect 1101 2460 1117 2524
rect 1181 2460 1197 2524
rect 1261 2460 1277 2524
rect 1341 2460 1357 2524
rect 1421 2460 1437 2524
rect 1501 2460 1517 2524
rect 1581 2460 1597 2524
rect 1661 2460 1677 2524
rect 1741 2460 1757 2524
rect 1821 2460 1837 2524
rect 1901 2460 1917 2524
rect 1981 2460 1997 2524
rect 2061 2460 2077 2524
rect 2141 2460 2157 2524
rect 2221 2460 2237 2524
rect 2301 2460 2317 2524
rect 2381 2460 2397 2524
rect 2461 2460 2477 2524
rect 2541 2460 3400 2524
rect -3400 2400 3400 2460
rect -3400 -2887 3400 -2800
rect -3400 -2951 -890 -2887
rect -826 -2951 -810 -2887
rect -746 -2951 -730 -2887
rect -666 -2951 -650 -2887
rect -586 -2951 -570 -2887
rect -506 -2951 -490 -2887
rect -426 -2951 -410 -2887
rect -346 -2951 -330 -2887
rect -266 -2951 -250 -2887
rect -186 -2951 -170 -2887
rect -106 -2951 -90 -2887
rect -26 -2951 -10 -2887
rect 54 -2951 70 -2887
rect 134 -2951 150 -2887
rect 214 -2951 230 -2887
rect 294 -2951 310 -2887
rect 374 -2951 390 -2887
rect 454 -2951 470 -2887
rect 534 -2951 550 -2887
rect 614 -2951 630 -2887
rect 694 -2951 710 -2887
rect 774 -2951 790 -2887
rect 854 -2951 870 -2887
rect 934 -2951 3400 -2887
rect -3400 -3154 3400 -2951
rect -3400 -3378 -3188 -3154
rect -2644 -3378 2644 -3154
rect 3188 -3378 3400 -3154
rect -3400 -3600 3400 -3378
use sky130_fd_pr__nfet_01v8_lvt_G98Z6N  sky130_fd_pr__nfet_01v8_lvt_G98Z6N_0
timestamp 1626486988
transform 1 0 -1557 0 1 -522
box -1345 -188 1345 188
use sky130_fd_pr__nfet_01v8_JP3XZJ  sky130_fd_pr__nfet_01v8_JP3XZJ_0
timestamp 1626486988
transform 1 0 28 0 1 -1924
box -2629 -397 2629 397
use sky130_fd_pr__nfet_01v8_V7Q58M  sky130_fd_pr__nfet_01v8_V7Q58M_0
timestamp 1626486988
transform 1 0 2462 0 1 -558
box -184 -288 184 288
use sky130_fd_pr__nfet_01v8_8B5GXQ  sky130_fd_pr__nfet_01v8_8B5GXQ_0
timestamp 1626486988
transform 1 0 1145 0 1 -484
box -829 -188 829 188
use sky130_fd_pr__pfet_01v8_H2H4BB  sky130_fd_pr__pfet_01v8_H2H4BB_1
timestamp 1626486988
transform 1 0 -1336 0 1 1913
box -1355 -200 1355 200
use sky130_fd_pr__pfet_01v8_H2H4BB  sky130_fd_pr__pfet_01v8_H2H4BB_0
timestamp 1626486988
transform 1 0 -1336 0 1 1239
box -1355 -200 1355 200
use sky130_fd_pr__pfet_01v8_hvt_ATGTW6  sky130_fd_pr__pfet_01v8_hvt_ATGTW6_0
timestamp 1626486988
transform 1 0 2462 0 1 1538
box -194 -500 194 500
use sky130_fd_pr__pfet_01v8_RC2RSP  sky130_fd_pr__pfet_01v8_RC2RSP_1
timestamp 1626486988
transform 1 0 1147 0 1 1238
box -839 -200 839 200
use sky130_fd_pr__pfet_01v8_RC2RSP  sky130_fd_pr__pfet_01v8_RC2RSP_0
timestamp 1626486988
transform 1 0 1147 0 1 1912
box -839 -200 839 200
<< labels >>
flabel metal1 s 886 -216 900 -202 1 FreeSans 600 0 0 0 vmirror
flabel metal1 s 436 -744 448 -730 1 FreeSans 600 0 0 0 vo1
flabel metal1 s 2726 -2168 2748 -2144 1 FreeSans 600 0 0 0 vtail
flabel metal2 s -820 -1444 -780 -1426 1 FreeSans 600 0 0 0 ibiasn
flabel metal2 s -452 -2416 -440 -2394 1 FreeSans 600 0 0 0 VSS
flabel metal1 s -2766 -264 -2732 -234 1 FreeSans 600 0 0 0 vcompm
flabel metal2 s -2292 -262 -2260 -238 1 FreeSans 600 0 0 0 vip
flabel metal2 s -1592 -802 -1560 -774 1 FreeSans 600 0 0 0 vim
flabel metal2 s -1592 -914 -1566 -890 1 FreeSans 600 0 0 0 vtail
flabel metal2 s -1654 -28 -1634 -4 1 FreeSans 600 0 0 0 vcompp
flabel metal1 s 2026 1582 2042 1600 1 FreeSans 600 0 0 0 vcompp
flabel metal1 s 1522 1686 1534 1696 1 FreeSans 600 0 0 0 vcompm
flabel metal2 s 1500 1502 1516 1514 1 FreeSans 600 0 0 0 vo1
flabel metal2 s 824 832 836 848 1 FreeSans 600 0 0 0 vmirror
flabel metal1 s -2122 1544 -2104 1566 1 FreeSans 600 0 0 0 vcompm
flabel metal2 s 2586 472 2596 480 1 FreeSans 600 0 0 0 vo
flabel metal2 s -720 2168 -702 2188 1 FreeSans 600 0 0 0 vcompp
flabel metal4 s -1674 2724 -1612 2786 1 FreeSans 600 0 0 0 VDD
<< properties >>
string FIXED_BBOX -3272 -3472 3272 332
<< end >>
