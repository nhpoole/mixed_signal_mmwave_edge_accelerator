magic
tech sky130A
magscale 1 2
timestamp 1626065694
<< checkpaint >>
rect -1319 -1314 1469 2714
<< nwell >>
rect -54 -54 204 1454
<< scpmos >>
rect 60 0 90 1400
<< pdiff >>
rect 0 0 60 1400
rect 90 0 150 1400
<< poly >>
rect 60 1400 90 1426
rect 60 -26 90 0
<< locali >>
rect 8 667 42 733
rect 108 667 142 733
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_0
timestamp 1626065694
transform 1 0 100 0 1 667
box -59 -51 109 117
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_1
timestamp 1626065694
transform 1 0 0 0 1 667
box -59 -51 109 117
<< labels >>
rlabel locali s 25 700 25 700 4 S
rlabel locali s 125 700 125 700 4 D
rlabel poly s 75 700 75 700 4 G
<< properties >>
string FIXED_BBOX -54 -54 204 1454
<< end >>
