magic
tech sky130A
magscale 1 2
timestamp 1621983599
<< nwell >>
rect -5058 4282 5458 10358
<< pwell >>
rect -5058 1752 5458 4118
<< nmos >>
rect -4550 3512 -4150 3712
rect -4092 3512 -3692 3712
rect -3634 3512 -3234 3712
rect -3176 3512 -2776 3712
rect -2718 3512 -2318 3712
rect -2260 3512 -1860 3712
rect -1802 3512 -1402 3712
rect -1344 3512 -944 3712
rect -886 3512 -486 3712
rect -428 3512 -28 3712
rect 450 3512 850 3712
rect 908 3512 1308 3712
rect 1366 3512 1766 3712
rect 1824 3512 2224 3712
rect 2282 3512 2682 3712
rect 2740 3512 3140 3712
rect 3198 3512 3598 3712
rect 3656 3512 4056 3712
rect 4114 3512 4514 3712
rect 4572 3512 4972 3712
rect -4550 2844 -4150 3044
rect -4092 2844 -3692 3044
rect -3634 2844 -3234 3044
rect -3176 2844 -2776 3044
rect -2718 2844 -2318 3044
rect -2260 2844 -1860 3044
rect -1802 2844 -1402 3044
rect -1344 2844 -944 3044
rect -886 2844 -486 3044
rect -428 2844 -28 3044
<< pmoshvt >>
rect -3990 7270 -3590 8870
rect -3532 7270 -3132 8870
rect -3074 7270 -2674 8870
rect -2616 7270 -2216 8870
rect -2158 7270 -1758 8870
rect -1700 7270 -1300 8870
rect -1242 7270 -842 8870
rect -784 7270 -384 8870
rect -326 7270 74 8870
rect 132 7270 532 8870
rect 590 7270 990 8870
rect 1048 7270 1448 8870
rect 1506 7270 1906 8870
rect 1964 7270 2364 8870
rect 2422 7270 2822 8870
rect 2880 7270 3280 8870
rect 3338 7270 3738 8870
rect 3796 7270 4196 8870
rect -4549 5005 -4149 6205
rect -4091 5005 -3691 6205
rect -3633 5005 -3233 6205
rect -3175 5005 -2775 6205
rect -2717 5005 -2317 6205
rect -2259 5005 -1859 6205
rect -1801 5005 -1401 6205
rect -1343 5005 -943 6205
rect -885 5005 -485 6205
rect -427 5005 -27 6205
rect 451 5005 851 6205
rect 909 5005 1309 6205
rect 1367 5005 1767 6205
rect 1825 5005 2225 6205
rect 2283 5005 2683 6205
rect 2741 5005 3141 6205
rect 3199 5005 3599 6205
rect 3657 5005 4057 6205
rect 4115 5005 4515 6205
rect 4573 5005 4973 6205
<< ndiff >>
rect -4608 3700 -4550 3712
rect -4608 3524 -4596 3700
rect -4562 3524 -4550 3700
rect -4608 3512 -4550 3524
rect -4150 3700 -4092 3712
rect -4150 3524 -4138 3700
rect -4104 3524 -4092 3700
rect -4150 3512 -4092 3524
rect -3692 3700 -3634 3712
rect -3692 3524 -3680 3700
rect -3646 3524 -3634 3700
rect -3692 3512 -3634 3524
rect -3234 3700 -3176 3712
rect -3234 3524 -3222 3700
rect -3188 3524 -3176 3700
rect -3234 3512 -3176 3524
rect -2776 3700 -2718 3712
rect -2776 3524 -2764 3700
rect -2730 3524 -2718 3700
rect -2776 3512 -2718 3524
rect -2318 3700 -2260 3712
rect -2318 3524 -2306 3700
rect -2272 3524 -2260 3700
rect -2318 3512 -2260 3524
rect -1860 3700 -1802 3712
rect -1860 3524 -1848 3700
rect -1814 3524 -1802 3700
rect -1860 3512 -1802 3524
rect -1402 3700 -1344 3712
rect -1402 3524 -1390 3700
rect -1356 3524 -1344 3700
rect -1402 3512 -1344 3524
rect -944 3700 -886 3712
rect -944 3524 -932 3700
rect -898 3524 -886 3700
rect -944 3512 -886 3524
rect -486 3700 -428 3712
rect -486 3524 -474 3700
rect -440 3524 -428 3700
rect -486 3512 -428 3524
rect -28 3700 30 3712
rect -28 3524 -16 3700
rect 18 3524 30 3700
rect -28 3512 30 3524
rect 392 3700 450 3712
rect 392 3524 404 3700
rect 438 3524 450 3700
rect 392 3512 450 3524
rect 850 3700 908 3712
rect 850 3524 862 3700
rect 896 3524 908 3700
rect 850 3512 908 3524
rect 1308 3700 1366 3712
rect 1308 3524 1320 3700
rect 1354 3524 1366 3700
rect 1308 3512 1366 3524
rect 1766 3700 1824 3712
rect 1766 3524 1778 3700
rect 1812 3524 1824 3700
rect 1766 3512 1824 3524
rect 2224 3700 2282 3712
rect 2224 3524 2236 3700
rect 2270 3524 2282 3700
rect 2224 3512 2282 3524
rect 2682 3700 2740 3712
rect 2682 3524 2694 3700
rect 2728 3524 2740 3700
rect 2682 3512 2740 3524
rect 3140 3700 3198 3712
rect 3140 3524 3152 3700
rect 3186 3524 3198 3700
rect 3140 3512 3198 3524
rect 3598 3700 3656 3712
rect 3598 3524 3610 3700
rect 3644 3524 3656 3700
rect 3598 3512 3656 3524
rect 4056 3700 4114 3712
rect 4056 3524 4068 3700
rect 4102 3524 4114 3700
rect 4056 3512 4114 3524
rect 4514 3700 4572 3712
rect 4514 3524 4526 3700
rect 4560 3524 4572 3700
rect 4514 3512 4572 3524
rect 4972 3700 5030 3712
rect 4972 3524 4984 3700
rect 5018 3524 5030 3700
rect 4972 3512 5030 3524
rect -4608 3032 -4550 3044
rect -4608 2856 -4596 3032
rect -4562 2856 -4550 3032
rect -4608 2844 -4550 2856
rect -4150 3032 -4092 3044
rect -4150 2856 -4138 3032
rect -4104 2856 -4092 3032
rect -4150 2844 -4092 2856
rect -3692 3032 -3634 3044
rect -3692 2856 -3680 3032
rect -3646 2856 -3634 3032
rect -3692 2844 -3634 2856
rect -3234 3032 -3176 3044
rect -3234 2856 -3222 3032
rect -3188 2856 -3176 3032
rect -3234 2844 -3176 2856
rect -2776 3032 -2718 3044
rect -2776 2856 -2764 3032
rect -2730 2856 -2718 3032
rect -2776 2844 -2718 2856
rect -2318 3032 -2260 3044
rect -2318 2856 -2306 3032
rect -2272 2856 -2260 3032
rect -2318 2844 -2260 2856
rect -1860 3032 -1802 3044
rect -1860 2856 -1848 3032
rect -1814 2856 -1802 3032
rect -1860 2844 -1802 2856
rect -1402 3032 -1344 3044
rect -1402 2856 -1390 3032
rect -1356 2856 -1344 3032
rect -1402 2844 -1344 2856
rect -944 3032 -886 3044
rect -944 2856 -932 3032
rect -898 2856 -886 3032
rect -944 2844 -886 2856
rect -486 3032 -428 3044
rect -486 2856 -474 3032
rect -440 2856 -428 3032
rect -486 2844 -428 2856
rect -28 3032 30 3044
rect -28 2856 -16 3032
rect 18 2856 30 3032
rect -28 2844 30 2856
<< pdiff >>
rect -4048 8858 -3990 8870
rect -4048 7282 -4036 8858
rect -4002 7282 -3990 8858
rect -4048 7270 -3990 7282
rect -3590 8858 -3532 8870
rect -3590 7282 -3578 8858
rect -3544 7282 -3532 8858
rect -3590 7270 -3532 7282
rect -3132 8858 -3074 8870
rect -3132 7282 -3120 8858
rect -3086 7282 -3074 8858
rect -3132 7270 -3074 7282
rect -2674 8858 -2616 8870
rect -2674 7282 -2662 8858
rect -2628 7282 -2616 8858
rect -2674 7270 -2616 7282
rect -2216 8858 -2158 8870
rect -2216 7282 -2204 8858
rect -2170 7282 -2158 8858
rect -2216 7270 -2158 7282
rect -1758 8858 -1700 8870
rect -1758 7282 -1746 8858
rect -1712 7282 -1700 8858
rect -1758 7270 -1700 7282
rect -1300 8858 -1242 8870
rect -1300 7282 -1288 8858
rect -1254 7282 -1242 8858
rect -1300 7270 -1242 7282
rect -842 8858 -784 8870
rect -842 7282 -830 8858
rect -796 7282 -784 8858
rect -842 7270 -784 7282
rect -384 8858 -326 8870
rect -384 7282 -372 8858
rect -338 7282 -326 8858
rect -384 7270 -326 7282
rect 74 8858 132 8870
rect 74 7282 86 8858
rect 120 7282 132 8858
rect 74 7270 132 7282
rect 532 8858 590 8870
rect 532 7282 544 8858
rect 578 7282 590 8858
rect 532 7270 590 7282
rect 990 8858 1048 8870
rect 990 7282 1002 8858
rect 1036 7282 1048 8858
rect 990 7270 1048 7282
rect 1448 8858 1506 8870
rect 1448 7282 1460 8858
rect 1494 7282 1506 8858
rect 1448 7270 1506 7282
rect 1906 8858 1964 8870
rect 1906 7282 1918 8858
rect 1952 7282 1964 8858
rect 1906 7270 1964 7282
rect 2364 8858 2422 8870
rect 2364 7282 2376 8858
rect 2410 7282 2422 8858
rect 2364 7270 2422 7282
rect 2822 8858 2880 8870
rect 2822 7282 2834 8858
rect 2868 7282 2880 8858
rect 2822 7270 2880 7282
rect 3280 8858 3338 8870
rect 3280 7282 3292 8858
rect 3326 7282 3338 8858
rect 3280 7270 3338 7282
rect 3738 8858 3796 8870
rect 3738 7282 3750 8858
rect 3784 7282 3796 8858
rect 3738 7270 3796 7282
rect 4196 8858 4254 8870
rect 4196 7282 4208 8858
rect 4242 7282 4254 8858
rect 4196 7270 4254 7282
rect -4607 6193 -4549 6205
rect -4607 5017 -4595 6193
rect -4561 5017 -4549 6193
rect -4607 5005 -4549 5017
rect -4149 6193 -4091 6205
rect -4149 5017 -4137 6193
rect -4103 5017 -4091 6193
rect -4149 5005 -4091 5017
rect -3691 6193 -3633 6205
rect -3691 5017 -3679 6193
rect -3645 5017 -3633 6193
rect -3691 5005 -3633 5017
rect -3233 6193 -3175 6205
rect -3233 5017 -3221 6193
rect -3187 5017 -3175 6193
rect -3233 5005 -3175 5017
rect -2775 6193 -2717 6205
rect -2775 5017 -2763 6193
rect -2729 5017 -2717 6193
rect -2775 5005 -2717 5017
rect -2317 6193 -2259 6205
rect -2317 5017 -2305 6193
rect -2271 5017 -2259 6193
rect -2317 5005 -2259 5017
rect -1859 6193 -1801 6205
rect -1859 5017 -1847 6193
rect -1813 5017 -1801 6193
rect -1859 5005 -1801 5017
rect -1401 6193 -1343 6205
rect -1401 5017 -1389 6193
rect -1355 5017 -1343 6193
rect -1401 5005 -1343 5017
rect -943 6193 -885 6205
rect -943 5017 -931 6193
rect -897 5017 -885 6193
rect -943 5005 -885 5017
rect -485 6193 -427 6205
rect -485 5017 -473 6193
rect -439 5017 -427 6193
rect -485 5005 -427 5017
rect -27 6193 31 6205
rect -27 5017 -15 6193
rect 19 5017 31 6193
rect -27 5005 31 5017
rect 393 6193 451 6205
rect 393 5017 405 6193
rect 439 5017 451 6193
rect 393 5005 451 5017
rect 851 6193 909 6205
rect 851 5017 863 6193
rect 897 5017 909 6193
rect 851 5005 909 5017
rect 1309 6193 1367 6205
rect 1309 5017 1321 6193
rect 1355 5017 1367 6193
rect 1309 5005 1367 5017
rect 1767 6193 1825 6205
rect 1767 5017 1779 6193
rect 1813 5017 1825 6193
rect 1767 5005 1825 5017
rect 2225 6193 2283 6205
rect 2225 5017 2237 6193
rect 2271 5017 2283 6193
rect 2225 5005 2283 5017
rect 2683 6193 2741 6205
rect 2683 5017 2695 6193
rect 2729 5017 2741 6193
rect 2683 5005 2741 5017
rect 3141 6193 3199 6205
rect 3141 5017 3153 6193
rect 3187 5017 3199 6193
rect 3141 5005 3199 5017
rect 3599 6193 3657 6205
rect 3599 5017 3611 6193
rect 3645 5017 3657 6193
rect 3599 5005 3657 5017
rect 4057 6193 4115 6205
rect 4057 5017 4069 6193
rect 4103 5017 4115 6193
rect 4057 5005 4115 5017
rect 4515 6193 4573 6205
rect 4515 5017 4527 6193
rect 4561 5017 4573 6193
rect 4515 5005 4573 5017
rect 4973 6193 5031 6205
rect 4973 5017 4985 6193
rect 5019 5017 5031 6193
rect 4973 5005 5031 5017
<< ndiffc >>
rect -4596 3524 -4562 3700
rect -4138 3524 -4104 3700
rect -3680 3524 -3646 3700
rect -3222 3524 -3188 3700
rect -2764 3524 -2730 3700
rect -2306 3524 -2272 3700
rect -1848 3524 -1814 3700
rect -1390 3524 -1356 3700
rect -932 3524 -898 3700
rect -474 3524 -440 3700
rect -16 3524 18 3700
rect 404 3524 438 3700
rect 862 3524 896 3700
rect 1320 3524 1354 3700
rect 1778 3524 1812 3700
rect 2236 3524 2270 3700
rect 2694 3524 2728 3700
rect 3152 3524 3186 3700
rect 3610 3524 3644 3700
rect 4068 3524 4102 3700
rect 4526 3524 4560 3700
rect 4984 3524 5018 3700
rect -4596 2856 -4562 3032
rect -4138 2856 -4104 3032
rect -3680 2856 -3646 3032
rect -3222 2856 -3188 3032
rect -2764 2856 -2730 3032
rect -2306 2856 -2272 3032
rect -1848 2856 -1814 3032
rect -1390 2856 -1356 3032
rect -932 2856 -898 3032
rect -474 2856 -440 3032
rect -16 2856 18 3032
<< pdiffc >>
rect -4036 7282 -4002 8858
rect -3578 7282 -3544 8858
rect -3120 7282 -3086 8858
rect -2662 7282 -2628 8858
rect -2204 7282 -2170 8858
rect -1746 7282 -1712 8858
rect -1288 7282 -1254 8858
rect -830 7282 -796 8858
rect -372 7282 -338 8858
rect 86 7282 120 8858
rect 544 7282 578 8858
rect 1002 7282 1036 8858
rect 1460 7282 1494 8858
rect 1918 7282 1952 8858
rect 2376 7282 2410 8858
rect 2834 7282 2868 8858
rect 3292 7282 3326 8858
rect 3750 7282 3784 8858
rect 4208 7282 4242 8858
rect -4595 5017 -4561 6193
rect -4137 5017 -4103 6193
rect -3679 5017 -3645 6193
rect -3221 5017 -3187 6193
rect -2763 5017 -2729 6193
rect -2305 5017 -2271 6193
rect -1847 5017 -1813 6193
rect -1389 5017 -1355 6193
rect -931 5017 -897 6193
rect -473 5017 -439 6193
rect -15 5017 19 6193
rect 405 5017 439 6193
rect 863 5017 897 6193
rect 1321 5017 1355 6193
rect 1779 5017 1813 6193
rect 2237 5017 2271 6193
rect 2695 5017 2729 6193
rect 3153 5017 3187 6193
rect 3611 5017 3645 6193
rect 4069 5017 4103 6193
rect 4527 5017 4561 6193
rect 4985 5017 5019 6193
<< psubdiff >>
rect -5022 4142 -4860 4242
rect 5260 4142 5422 4242
rect -5022 4080 -4922 4142
rect 5322 4080 5422 4142
rect -5022 1878 -4922 1940
rect 5322 1878 5422 1940
rect -5022 1778 -4860 1878
rect 5260 1778 5422 1878
<< nsubdiff >>
rect -5022 10222 -4860 10322
rect 5260 10222 5422 10322
rect -5022 10160 -4922 10222
rect 5322 10160 5422 10222
rect -5022 4578 -4922 4640
rect 5322 4578 5422 4640
rect -5022 4478 -4860 4578
rect 5260 4478 5422 4578
<< psubdiffcont >>
rect -4860 4142 5260 4242
rect -5022 1940 -4922 4080
rect 5322 1940 5422 4080
rect -4860 1778 5260 1878
<< nsubdiffcont >>
rect -4860 10222 5260 10322
rect -5022 4640 -4922 10160
rect 5322 4640 5422 10160
rect -4860 4478 5260 4578
<< poly >>
rect -3916 8951 -3664 8967
rect -3916 8934 -3900 8951
rect -3990 8917 -3900 8934
rect -3680 8934 -3664 8951
rect -3458 8951 -3206 8967
rect -3458 8934 -3442 8951
rect -3680 8917 -3590 8934
rect -3990 8870 -3590 8917
rect -3532 8917 -3442 8934
rect -3222 8934 -3206 8951
rect -3000 8951 -2748 8967
rect -3000 8934 -2984 8951
rect -3222 8917 -3132 8934
rect -3532 8870 -3132 8917
rect -3074 8917 -2984 8934
rect -2764 8934 -2748 8951
rect -2542 8951 -2290 8967
rect -2542 8934 -2526 8951
rect -2764 8917 -2674 8934
rect -3074 8870 -2674 8917
rect -2616 8917 -2526 8934
rect -2306 8934 -2290 8951
rect -2084 8951 -1832 8967
rect -2084 8934 -2068 8951
rect -2306 8917 -2216 8934
rect -2616 8870 -2216 8917
rect -2158 8917 -2068 8934
rect -1848 8934 -1832 8951
rect -1626 8951 -1374 8967
rect -1626 8934 -1610 8951
rect -1848 8917 -1758 8934
rect -2158 8870 -1758 8917
rect -1700 8917 -1610 8934
rect -1390 8934 -1374 8951
rect -1168 8951 -916 8967
rect -1168 8934 -1152 8951
rect -1390 8917 -1300 8934
rect -1700 8870 -1300 8917
rect -1242 8917 -1152 8934
rect -932 8934 -916 8951
rect -710 8951 -458 8967
rect -710 8934 -694 8951
rect -932 8917 -842 8934
rect -1242 8870 -842 8917
rect -784 8917 -694 8934
rect -474 8934 -458 8951
rect -252 8951 0 8967
rect -252 8934 -236 8951
rect -474 8917 -384 8934
rect -784 8870 -384 8917
rect -326 8917 -236 8934
rect -16 8934 0 8951
rect 206 8951 458 8967
rect 206 8934 222 8951
rect -16 8917 74 8934
rect -326 8870 74 8917
rect 132 8917 222 8934
rect 442 8934 458 8951
rect 664 8951 916 8967
rect 664 8934 680 8951
rect 442 8917 532 8934
rect 132 8870 532 8917
rect 590 8917 680 8934
rect 900 8934 916 8951
rect 1122 8951 1374 8967
rect 1122 8934 1138 8951
rect 900 8917 990 8934
rect 590 8870 990 8917
rect 1048 8917 1138 8934
rect 1358 8934 1374 8951
rect 1580 8951 1832 8967
rect 1580 8934 1596 8951
rect 1358 8917 1448 8934
rect 1048 8870 1448 8917
rect 1506 8917 1596 8934
rect 1816 8934 1832 8951
rect 2038 8951 2290 8967
rect 2038 8934 2054 8951
rect 1816 8917 1906 8934
rect 1506 8870 1906 8917
rect 1964 8917 2054 8934
rect 2274 8934 2290 8951
rect 2496 8951 2748 8967
rect 2496 8934 2512 8951
rect 2274 8917 2364 8934
rect 1964 8870 2364 8917
rect 2422 8917 2512 8934
rect 2732 8934 2748 8951
rect 2954 8951 3206 8967
rect 2954 8934 2970 8951
rect 2732 8917 2822 8934
rect 2422 8870 2822 8917
rect 2880 8917 2970 8934
rect 3190 8934 3206 8951
rect 3412 8951 3664 8967
rect 3412 8934 3428 8951
rect 3190 8917 3280 8934
rect 2880 8870 3280 8917
rect 3338 8917 3428 8934
rect 3648 8934 3664 8951
rect 3870 8951 4122 8967
rect 3870 8934 3886 8951
rect 3648 8917 3738 8934
rect 3338 8870 3738 8917
rect 3796 8917 3886 8934
rect 4106 8934 4122 8951
rect 4106 8917 4196 8934
rect 3796 8870 4196 8917
rect -3990 7223 -3590 7270
rect -3990 7206 -3900 7223
rect -3916 7189 -3900 7206
rect -3680 7206 -3590 7223
rect -3532 7223 -3132 7270
rect -3532 7206 -3442 7223
rect -3680 7189 -3664 7206
rect -3916 7173 -3664 7189
rect -3458 7189 -3442 7206
rect -3222 7206 -3132 7223
rect -3074 7223 -2674 7270
rect -3074 7206 -2984 7223
rect -3222 7189 -3206 7206
rect -3458 7173 -3206 7189
rect -3000 7189 -2984 7206
rect -2764 7206 -2674 7223
rect -2616 7223 -2216 7270
rect -2616 7206 -2526 7223
rect -2764 7189 -2748 7206
rect -3000 7173 -2748 7189
rect -2542 7189 -2526 7206
rect -2306 7206 -2216 7223
rect -2158 7223 -1758 7270
rect -2158 7206 -2068 7223
rect -2306 7189 -2290 7206
rect -2542 7173 -2290 7189
rect -2084 7189 -2068 7206
rect -1848 7206 -1758 7223
rect -1700 7223 -1300 7270
rect -1700 7206 -1610 7223
rect -1848 7189 -1832 7206
rect -2084 7173 -1832 7189
rect -1626 7189 -1610 7206
rect -1390 7206 -1300 7223
rect -1242 7223 -842 7270
rect -1242 7206 -1152 7223
rect -1390 7189 -1374 7206
rect -1626 7173 -1374 7189
rect -1168 7189 -1152 7206
rect -932 7206 -842 7223
rect -784 7223 -384 7270
rect -784 7206 -694 7223
rect -932 7189 -916 7206
rect -1168 7173 -916 7189
rect -710 7189 -694 7206
rect -474 7206 -384 7223
rect -326 7223 74 7270
rect -326 7206 -236 7223
rect -474 7189 -458 7206
rect -710 7173 -458 7189
rect -252 7189 -236 7206
rect -16 7206 74 7223
rect 132 7223 532 7270
rect 132 7206 222 7223
rect -16 7189 0 7206
rect -252 7173 0 7189
rect 206 7189 222 7206
rect 442 7206 532 7223
rect 590 7223 990 7270
rect 590 7206 680 7223
rect 442 7189 458 7206
rect 206 7173 458 7189
rect 664 7189 680 7206
rect 900 7206 990 7223
rect 1048 7223 1448 7270
rect 1048 7206 1138 7223
rect 900 7189 916 7206
rect 664 7173 916 7189
rect 1122 7189 1138 7206
rect 1358 7206 1448 7223
rect 1506 7223 1906 7270
rect 1506 7206 1596 7223
rect 1358 7189 1374 7206
rect 1122 7173 1374 7189
rect 1580 7189 1596 7206
rect 1816 7206 1906 7223
rect 1964 7223 2364 7270
rect 1964 7206 2054 7223
rect 1816 7189 1832 7206
rect 1580 7173 1832 7189
rect 2038 7189 2054 7206
rect 2274 7206 2364 7223
rect 2422 7223 2822 7270
rect 2422 7206 2512 7223
rect 2274 7189 2290 7206
rect 2038 7173 2290 7189
rect 2496 7189 2512 7206
rect 2732 7206 2822 7223
rect 2880 7223 3280 7270
rect 2880 7206 2970 7223
rect 2732 7189 2748 7206
rect 2496 7173 2748 7189
rect 2954 7189 2970 7206
rect 3190 7206 3280 7223
rect 3338 7223 3738 7270
rect 3338 7206 3428 7223
rect 3190 7189 3206 7206
rect 2954 7173 3206 7189
rect 3412 7189 3428 7206
rect 3648 7206 3738 7223
rect 3796 7223 4196 7270
rect 3796 7206 3886 7223
rect 3648 7189 3664 7206
rect 3412 7173 3664 7189
rect 3870 7189 3886 7206
rect 4106 7206 4196 7223
rect 4106 7189 4122 7206
rect 3870 7173 4122 7189
rect -4475 6286 -4223 6302
rect -4475 6269 -4459 6286
rect -4549 6252 -4459 6269
rect -4239 6269 -4223 6286
rect -4017 6286 -3765 6302
rect -4017 6269 -4001 6286
rect -4239 6252 -4149 6269
rect -4549 6205 -4149 6252
rect -4091 6252 -4001 6269
rect -3781 6269 -3765 6286
rect -3559 6286 -3307 6302
rect -3559 6269 -3543 6286
rect -3781 6252 -3691 6269
rect -4091 6205 -3691 6252
rect -3633 6252 -3543 6269
rect -3323 6269 -3307 6286
rect -3101 6286 -2849 6302
rect -3101 6269 -3085 6286
rect -3323 6252 -3233 6269
rect -3633 6205 -3233 6252
rect -3175 6252 -3085 6269
rect -2865 6269 -2849 6286
rect -2643 6286 -2391 6302
rect -2643 6269 -2627 6286
rect -2865 6252 -2775 6269
rect -3175 6205 -2775 6252
rect -2717 6252 -2627 6269
rect -2407 6269 -2391 6286
rect -2185 6286 -1933 6302
rect -2185 6269 -2169 6286
rect -2407 6252 -2317 6269
rect -2717 6205 -2317 6252
rect -2259 6252 -2169 6269
rect -1949 6269 -1933 6286
rect -1727 6286 -1475 6302
rect -1727 6269 -1711 6286
rect -1949 6252 -1859 6269
rect -2259 6205 -1859 6252
rect -1801 6252 -1711 6269
rect -1491 6269 -1475 6286
rect -1269 6286 -1017 6302
rect -1269 6269 -1253 6286
rect -1491 6252 -1401 6269
rect -1801 6205 -1401 6252
rect -1343 6252 -1253 6269
rect -1033 6269 -1017 6286
rect -811 6286 -559 6302
rect -811 6269 -795 6286
rect -1033 6252 -943 6269
rect -1343 6205 -943 6252
rect -885 6252 -795 6269
rect -575 6269 -559 6286
rect -353 6286 -101 6302
rect -353 6269 -337 6286
rect -575 6252 -485 6269
rect -885 6205 -485 6252
rect -427 6252 -337 6269
rect -117 6269 -101 6286
rect 525 6286 777 6302
rect 525 6269 541 6286
rect -117 6252 -27 6269
rect -427 6205 -27 6252
rect 451 6252 541 6269
rect 761 6269 777 6286
rect 983 6286 1235 6302
rect 983 6269 999 6286
rect 761 6252 851 6269
rect 451 6205 851 6252
rect 909 6252 999 6269
rect 1219 6269 1235 6286
rect 1441 6286 1693 6302
rect 1441 6269 1457 6286
rect 1219 6252 1309 6269
rect 909 6205 1309 6252
rect 1367 6252 1457 6269
rect 1677 6269 1693 6286
rect 1899 6286 2151 6302
rect 1899 6269 1915 6286
rect 1677 6252 1767 6269
rect 1367 6205 1767 6252
rect 1825 6252 1915 6269
rect 2135 6269 2151 6286
rect 2357 6286 2609 6302
rect 2357 6269 2373 6286
rect 2135 6252 2225 6269
rect 1825 6205 2225 6252
rect 2283 6252 2373 6269
rect 2593 6269 2609 6286
rect 2815 6286 3067 6302
rect 2815 6269 2831 6286
rect 2593 6252 2683 6269
rect 2283 6205 2683 6252
rect 2741 6252 2831 6269
rect 3051 6269 3067 6286
rect 3273 6286 3525 6302
rect 3273 6269 3289 6286
rect 3051 6252 3141 6269
rect 2741 6205 3141 6252
rect 3199 6252 3289 6269
rect 3509 6269 3525 6286
rect 3731 6286 3983 6302
rect 3731 6269 3747 6286
rect 3509 6252 3599 6269
rect 3199 6205 3599 6252
rect 3657 6252 3747 6269
rect 3967 6269 3983 6286
rect 4189 6286 4441 6302
rect 4189 6269 4205 6286
rect 3967 6252 4057 6269
rect 3657 6205 4057 6252
rect 4115 6252 4205 6269
rect 4425 6269 4441 6286
rect 4647 6286 4899 6302
rect 4647 6269 4663 6286
rect 4425 6252 4515 6269
rect 4115 6205 4515 6252
rect 4573 6252 4663 6269
rect 4883 6269 4899 6286
rect 4883 6252 4973 6269
rect 4573 6205 4973 6252
rect -4549 4958 -4149 5005
rect -4549 4941 -4459 4958
rect -4475 4924 -4459 4941
rect -4239 4941 -4149 4958
rect -4091 4958 -3691 5005
rect -4091 4941 -4001 4958
rect -4239 4924 -4223 4941
rect -4475 4908 -4223 4924
rect -4017 4924 -4001 4941
rect -3781 4941 -3691 4958
rect -3633 4958 -3233 5005
rect -3633 4941 -3543 4958
rect -3781 4924 -3765 4941
rect -4017 4908 -3765 4924
rect -3559 4924 -3543 4941
rect -3323 4941 -3233 4958
rect -3175 4958 -2775 5005
rect -3175 4941 -3085 4958
rect -3323 4924 -3307 4941
rect -3559 4908 -3307 4924
rect -3101 4924 -3085 4941
rect -2865 4941 -2775 4958
rect -2717 4958 -2317 5005
rect -2717 4941 -2627 4958
rect -2865 4924 -2849 4941
rect -3101 4908 -2849 4924
rect -2643 4924 -2627 4941
rect -2407 4941 -2317 4958
rect -2259 4958 -1859 5005
rect -2259 4941 -2169 4958
rect -2407 4924 -2391 4941
rect -2643 4908 -2391 4924
rect -2185 4924 -2169 4941
rect -1949 4941 -1859 4958
rect -1801 4958 -1401 5005
rect -1801 4941 -1711 4958
rect -1949 4924 -1933 4941
rect -2185 4908 -1933 4924
rect -1727 4924 -1711 4941
rect -1491 4941 -1401 4958
rect -1343 4958 -943 5005
rect -1343 4941 -1253 4958
rect -1491 4924 -1475 4941
rect -1727 4908 -1475 4924
rect -1269 4924 -1253 4941
rect -1033 4941 -943 4958
rect -885 4958 -485 5005
rect -885 4941 -795 4958
rect -1033 4924 -1017 4941
rect -1269 4908 -1017 4924
rect -811 4924 -795 4941
rect -575 4941 -485 4958
rect -427 4958 -27 5005
rect -427 4941 -337 4958
rect -575 4924 -559 4941
rect -811 4908 -559 4924
rect -353 4924 -337 4941
rect -117 4941 -27 4958
rect 451 4958 851 5005
rect 451 4941 541 4958
rect -117 4924 -101 4941
rect -353 4908 -101 4924
rect 525 4924 541 4941
rect 761 4941 851 4958
rect 909 4958 1309 5005
rect 909 4941 999 4958
rect 761 4924 777 4941
rect 525 4908 777 4924
rect 983 4924 999 4941
rect 1219 4941 1309 4958
rect 1367 4958 1767 5005
rect 1367 4941 1457 4958
rect 1219 4924 1235 4941
rect 983 4908 1235 4924
rect 1441 4924 1457 4941
rect 1677 4941 1767 4958
rect 1825 4958 2225 5005
rect 1825 4941 1915 4958
rect 1677 4924 1693 4941
rect 1441 4908 1693 4924
rect 1899 4924 1915 4941
rect 2135 4941 2225 4958
rect 2283 4958 2683 5005
rect 2283 4941 2373 4958
rect 2135 4924 2151 4941
rect 1899 4908 2151 4924
rect 2357 4924 2373 4941
rect 2593 4941 2683 4958
rect 2741 4958 3141 5005
rect 2741 4941 2831 4958
rect 2593 4924 2609 4941
rect 2357 4908 2609 4924
rect 2815 4924 2831 4941
rect 3051 4941 3141 4958
rect 3199 4958 3599 5005
rect 3199 4941 3289 4958
rect 3051 4924 3067 4941
rect 2815 4908 3067 4924
rect 3273 4924 3289 4941
rect 3509 4941 3599 4958
rect 3657 4958 4057 5005
rect 3657 4941 3747 4958
rect 3509 4924 3525 4941
rect 3273 4908 3525 4924
rect 3731 4924 3747 4941
rect 3967 4941 4057 4958
rect 4115 4958 4515 5005
rect 4115 4941 4205 4958
rect 3967 4924 3983 4941
rect 3731 4908 3983 4924
rect 4189 4924 4205 4941
rect 4425 4941 4515 4958
rect 4573 4958 4973 5005
rect 4573 4941 4663 4958
rect 4425 4924 4441 4941
rect 4189 4908 4441 4924
rect 4647 4924 4663 4941
rect 4883 4941 4973 4958
rect 4883 4924 4899 4941
rect 4647 4908 4899 4924
rect -4476 3784 -4224 3800
rect -4476 3767 -4460 3784
rect -4550 3750 -4460 3767
rect -4240 3767 -4224 3784
rect -4018 3784 -3766 3800
rect -4018 3767 -4002 3784
rect -4240 3750 -4150 3767
rect -4550 3712 -4150 3750
rect -4092 3750 -4002 3767
rect -3782 3767 -3766 3784
rect -3560 3784 -3308 3800
rect -3560 3767 -3544 3784
rect -3782 3750 -3692 3767
rect -4092 3712 -3692 3750
rect -3634 3750 -3544 3767
rect -3324 3767 -3308 3784
rect -3102 3784 -2850 3800
rect -3102 3767 -3086 3784
rect -3324 3750 -3234 3767
rect -3634 3712 -3234 3750
rect -3176 3750 -3086 3767
rect -2866 3767 -2850 3784
rect -2644 3784 -2392 3800
rect -2644 3767 -2628 3784
rect -2866 3750 -2776 3767
rect -3176 3712 -2776 3750
rect -2718 3750 -2628 3767
rect -2408 3767 -2392 3784
rect -2186 3784 -1934 3800
rect -2186 3767 -2170 3784
rect -2408 3750 -2318 3767
rect -2718 3712 -2318 3750
rect -2260 3750 -2170 3767
rect -1950 3767 -1934 3784
rect -1728 3784 -1476 3800
rect -1728 3767 -1712 3784
rect -1950 3750 -1860 3767
rect -2260 3712 -1860 3750
rect -1802 3750 -1712 3767
rect -1492 3767 -1476 3784
rect -1270 3784 -1018 3800
rect -1270 3767 -1254 3784
rect -1492 3750 -1402 3767
rect -1802 3712 -1402 3750
rect -1344 3750 -1254 3767
rect -1034 3767 -1018 3784
rect -812 3784 -560 3800
rect -812 3767 -796 3784
rect -1034 3750 -944 3767
rect -1344 3712 -944 3750
rect -886 3750 -796 3767
rect -576 3767 -560 3784
rect -354 3784 -102 3800
rect -354 3767 -338 3784
rect -576 3750 -486 3767
rect -886 3712 -486 3750
rect -428 3750 -338 3767
rect -118 3767 -102 3784
rect 524 3784 776 3800
rect 524 3767 540 3784
rect -118 3750 -28 3767
rect -428 3712 -28 3750
rect 450 3750 540 3767
rect 760 3767 776 3784
rect 982 3784 1234 3800
rect 982 3767 998 3784
rect 760 3750 850 3767
rect 450 3712 850 3750
rect 908 3750 998 3767
rect 1218 3767 1234 3784
rect 1440 3784 1692 3800
rect 1440 3767 1456 3784
rect 1218 3750 1308 3767
rect 908 3712 1308 3750
rect 1366 3750 1456 3767
rect 1676 3767 1692 3784
rect 1898 3784 2150 3800
rect 1898 3767 1914 3784
rect 1676 3750 1766 3767
rect 1366 3712 1766 3750
rect 1824 3750 1914 3767
rect 2134 3767 2150 3784
rect 2356 3784 2608 3800
rect 2356 3767 2372 3784
rect 2134 3750 2224 3767
rect 1824 3712 2224 3750
rect 2282 3750 2372 3767
rect 2592 3767 2608 3784
rect 2814 3784 3066 3800
rect 2814 3767 2830 3784
rect 2592 3750 2682 3767
rect 2282 3712 2682 3750
rect 2740 3750 2830 3767
rect 3050 3767 3066 3784
rect 3272 3784 3524 3800
rect 3272 3767 3288 3784
rect 3050 3750 3140 3767
rect 2740 3712 3140 3750
rect 3198 3750 3288 3767
rect 3508 3767 3524 3784
rect 3730 3784 3982 3800
rect 3730 3767 3746 3784
rect 3508 3750 3598 3767
rect 3198 3712 3598 3750
rect 3656 3750 3746 3767
rect 3966 3767 3982 3784
rect 4188 3784 4440 3800
rect 4188 3767 4204 3784
rect 3966 3750 4056 3767
rect 3656 3712 4056 3750
rect 4114 3750 4204 3767
rect 4424 3767 4440 3784
rect 4646 3784 4898 3800
rect 4646 3767 4662 3784
rect 4424 3750 4514 3767
rect 4114 3712 4514 3750
rect 4572 3750 4662 3767
rect 4882 3767 4898 3784
rect 4882 3750 4972 3767
rect 4572 3712 4972 3750
rect -4550 3474 -4150 3512
rect -4550 3457 -4460 3474
rect -4476 3440 -4460 3457
rect -4240 3457 -4150 3474
rect -4092 3474 -3692 3512
rect -4092 3457 -4002 3474
rect -4240 3440 -4224 3457
rect -4476 3424 -4224 3440
rect -4018 3440 -4002 3457
rect -3782 3457 -3692 3474
rect -3634 3474 -3234 3512
rect -3634 3457 -3544 3474
rect -3782 3440 -3766 3457
rect -4018 3424 -3766 3440
rect -3560 3440 -3544 3457
rect -3324 3457 -3234 3474
rect -3176 3474 -2776 3512
rect -3176 3457 -3086 3474
rect -3324 3440 -3308 3457
rect -3560 3424 -3308 3440
rect -3102 3440 -3086 3457
rect -2866 3457 -2776 3474
rect -2718 3474 -2318 3512
rect -2718 3457 -2628 3474
rect -2866 3440 -2850 3457
rect -3102 3424 -2850 3440
rect -2644 3440 -2628 3457
rect -2408 3457 -2318 3474
rect -2260 3474 -1860 3512
rect -2260 3457 -2170 3474
rect -2408 3440 -2392 3457
rect -2644 3424 -2392 3440
rect -2186 3440 -2170 3457
rect -1950 3457 -1860 3474
rect -1802 3474 -1402 3512
rect -1802 3457 -1712 3474
rect -1950 3440 -1934 3457
rect -2186 3424 -1934 3440
rect -1728 3440 -1712 3457
rect -1492 3457 -1402 3474
rect -1344 3474 -944 3512
rect -1344 3457 -1254 3474
rect -1492 3440 -1476 3457
rect -1728 3424 -1476 3440
rect -1270 3440 -1254 3457
rect -1034 3457 -944 3474
rect -886 3474 -486 3512
rect -886 3457 -796 3474
rect -1034 3440 -1018 3457
rect -1270 3424 -1018 3440
rect -812 3440 -796 3457
rect -576 3457 -486 3474
rect -428 3474 -28 3512
rect -428 3457 -338 3474
rect -576 3440 -560 3457
rect -812 3424 -560 3440
rect -354 3440 -338 3457
rect -118 3457 -28 3474
rect 450 3474 850 3512
rect 450 3457 540 3474
rect -118 3440 -102 3457
rect -354 3424 -102 3440
rect 524 3440 540 3457
rect 760 3457 850 3474
rect 908 3474 1308 3512
rect 908 3457 998 3474
rect 760 3440 776 3457
rect 524 3424 776 3440
rect 982 3440 998 3457
rect 1218 3457 1308 3474
rect 1366 3474 1766 3512
rect 1366 3457 1456 3474
rect 1218 3440 1234 3457
rect 982 3424 1234 3440
rect 1440 3440 1456 3457
rect 1676 3457 1766 3474
rect 1824 3474 2224 3512
rect 1824 3457 1914 3474
rect 1676 3440 1692 3457
rect 1440 3424 1692 3440
rect 1898 3440 1914 3457
rect 2134 3457 2224 3474
rect 2282 3474 2682 3512
rect 2282 3457 2372 3474
rect 2134 3440 2150 3457
rect 1898 3424 2150 3440
rect 2356 3440 2372 3457
rect 2592 3457 2682 3474
rect 2740 3474 3140 3512
rect 2740 3457 2830 3474
rect 2592 3440 2608 3457
rect 2356 3424 2608 3440
rect 2814 3440 2830 3457
rect 3050 3457 3140 3474
rect 3198 3474 3598 3512
rect 3198 3457 3288 3474
rect 3050 3440 3066 3457
rect 2814 3424 3066 3440
rect 3272 3440 3288 3457
rect 3508 3457 3598 3474
rect 3656 3474 4056 3512
rect 3656 3457 3746 3474
rect 3508 3440 3524 3457
rect 3272 3424 3524 3440
rect 3730 3440 3746 3457
rect 3966 3457 4056 3474
rect 4114 3474 4514 3512
rect 4114 3457 4204 3474
rect 3966 3440 3982 3457
rect 3730 3424 3982 3440
rect 4188 3440 4204 3457
rect 4424 3457 4514 3474
rect 4572 3474 4972 3512
rect 4572 3457 4662 3474
rect 4424 3440 4440 3457
rect 4188 3424 4440 3440
rect 4646 3440 4662 3457
rect 4882 3457 4972 3474
rect 4882 3440 4898 3457
rect 4646 3424 4898 3440
rect -4476 3116 -4224 3132
rect -4476 3099 -4460 3116
rect -4550 3082 -4460 3099
rect -4240 3099 -4224 3116
rect -4018 3116 -3766 3132
rect -4018 3099 -4002 3116
rect -4240 3082 -4150 3099
rect -4550 3044 -4150 3082
rect -4092 3082 -4002 3099
rect -3782 3099 -3766 3116
rect -3560 3116 -3308 3132
rect -3560 3099 -3544 3116
rect -3782 3082 -3692 3099
rect -4092 3044 -3692 3082
rect -3634 3082 -3544 3099
rect -3324 3099 -3308 3116
rect -3102 3116 -2850 3132
rect -3102 3099 -3086 3116
rect -3324 3082 -3234 3099
rect -3634 3044 -3234 3082
rect -3176 3082 -3086 3099
rect -2866 3099 -2850 3116
rect -2644 3116 -2392 3132
rect -2644 3099 -2628 3116
rect -2866 3082 -2776 3099
rect -3176 3044 -2776 3082
rect -2718 3082 -2628 3099
rect -2408 3099 -2392 3116
rect -2186 3116 -1934 3132
rect -2186 3099 -2170 3116
rect -2408 3082 -2318 3099
rect -2718 3044 -2318 3082
rect -2260 3082 -2170 3099
rect -1950 3099 -1934 3116
rect -1728 3116 -1476 3132
rect -1728 3099 -1712 3116
rect -1950 3082 -1860 3099
rect -2260 3044 -1860 3082
rect -1802 3082 -1712 3099
rect -1492 3099 -1476 3116
rect -1270 3116 -1018 3132
rect -1270 3099 -1254 3116
rect -1492 3082 -1402 3099
rect -1802 3044 -1402 3082
rect -1344 3082 -1254 3099
rect -1034 3099 -1018 3116
rect -812 3116 -560 3132
rect -812 3099 -796 3116
rect -1034 3082 -944 3099
rect -1344 3044 -944 3082
rect -886 3082 -796 3099
rect -576 3099 -560 3116
rect -354 3116 -102 3132
rect -354 3099 -338 3116
rect -576 3082 -486 3099
rect -886 3044 -486 3082
rect -428 3082 -338 3099
rect -118 3099 -102 3116
rect -118 3082 -28 3099
rect -428 3044 -28 3082
rect -4550 2806 -4150 2844
rect -4550 2789 -4460 2806
rect -4476 2772 -4460 2789
rect -4240 2789 -4150 2806
rect -4092 2806 -3692 2844
rect -4092 2789 -4002 2806
rect -4240 2772 -4224 2789
rect -4476 2756 -4224 2772
rect -4018 2772 -4002 2789
rect -3782 2789 -3692 2806
rect -3634 2806 -3234 2844
rect -3634 2789 -3544 2806
rect -3782 2772 -3766 2789
rect -4018 2756 -3766 2772
rect -3560 2772 -3544 2789
rect -3324 2789 -3234 2806
rect -3176 2806 -2776 2844
rect -3176 2789 -3086 2806
rect -3324 2772 -3308 2789
rect -3560 2756 -3308 2772
rect -3102 2772 -3086 2789
rect -2866 2789 -2776 2806
rect -2718 2806 -2318 2844
rect -2718 2789 -2628 2806
rect -2866 2772 -2850 2789
rect -3102 2756 -2850 2772
rect -2644 2772 -2628 2789
rect -2408 2789 -2318 2806
rect -2260 2806 -1860 2844
rect -2260 2789 -2170 2806
rect -2408 2772 -2392 2789
rect -2644 2756 -2392 2772
rect -2186 2772 -2170 2789
rect -1950 2789 -1860 2806
rect -1802 2806 -1402 2844
rect -1802 2789 -1712 2806
rect -1950 2772 -1934 2789
rect -2186 2756 -1934 2772
rect -1728 2772 -1712 2789
rect -1492 2789 -1402 2806
rect -1344 2806 -944 2844
rect -1344 2789 -1254 2806
rect -1492 2772 -1476 2789
rect -1728 2756 -1476 2772
rect -1270 2772 -1254 2789
rect -1034 2789 -944 2806
rect -886 2806 -486 2844
rect -886 2789 -796 2806
rect -1034 2772 -1018 2789
rect -1270 2756 -1018 2772
rect -812 2772 -796 2789
rect -576 2789 -486 2806
rect -428 2806 -28 2844
rect -428 2789 -338 2806
rect -576 2772 -560 2789
rect -812 2756 -560 2772
rect -354 2772 -338 2789
rect -118 2789 -28 2806
rect -118 2772 -102 2789
rect -354 2756 -102 2772
<< polycont >>
rect -3900 8917 -3680 8951
rect -3442 8917 -3222 8951
rect -2984 8917 -2764 8951
rect -2526 8917 -2306 8951
rect -2068 8917 -1848 8951
rect -1610 8917 -1390 8951
rect -1152 8917 -932 8951
rect -694 8917 -474 8951
rect -236 8917 -16 8951
rect 222 8917 442 8951
rect 680 8917 900 8951
rect 1138 8917 1358 8951
rect 1596 8917 1816 8951
rect 2054 8917 2274 8951
rect 2512 8917 2732 8951
rect 2970 8917 3190 8951
rect 3428 8917 3648 8951
rect 3886 8917 4106 8951
rect -3900 7189 -3680 7223
rect -3442 7189 -3222 7223
rect -2984 7189 -2764 7223
rect -2526 7189 -2306 7223
rect -2068 7189 -1848 7223
rect -1610 7189 -1390 7223
rect -1152 7189 -932 7223
rect -694 7189 -474 7223
rect -236 7189 -16 7223
rect 222 7189 442 7223
rect 680 7189 900 7223
rect 1138 7189 1358 7223
rect 1596 7189 1816 7223
rect 2054 7189 2274 7223
rect 2512 7189 2732 7223
rect 2970 7189 3190 7223
rect 3428 7189 3648 7223
rect 3886 7189 4106 7223
rect -4459 6252 -4239 6286
rect -4001 6252 -3781 6286
rect -3543 6252 -3323 6286
rect -3085 6252 -2865 6286
rect -2627 6252 -2407 6286
rect -2169 6252 -1949 6286
rect -1711 6252 -1491 6286
rect -1253 6252 -1033 6286
rect -795 6252 -575 6286
rect -337 6252 -117 6286
rect 541 6252 761 6286
rect 999 6252 1219 6286
rect 1457 6252 1677 6286
rect 1915 6252 2135 6286
rect 2373 6252 2593 6286
rect 2831 6252 3051 6286
rect 3289 6252 3509 6286
rect 3747 6252 3967 6286
rect 4205 6252 4425 6286
rect 4663 6252 4883 6286
rect -4459 4924 -4239 4958
rect -4001 4924 -3781 4958
rect -3543 4924 -3323 4958
rect -3085 4924 -2865 4958
rect -2627 4924 -2407 4958
rect -2169 4924 -1949 4958
rect -1711 4924 -1491 4958
rect -1253 4924 -1033 4958
rect -795 4924 -575 4958
rect -337 4924 -117 4958
rect 541 4924 761 4958
rect 999 4924 1219 4958
rect 1457 4924 1677 4958
rect 1915 4924 2135 4958
rect 2373 4924 2593 4958
rect 2831 4924 3051 4958
rect 3289 4924 3509 4958
rect 3747 4924 3967 4958
rect 4205 4924 4425 4958
rect 4663 4924 4883 4958
rect -4460 3750 -4240 3784
rect -4002 3750 -3782 3784
rect -3544 3750 -3324 3784
rect -3086 3750 -2866 3784
rect -2628 3750 -2408 3784
rect -2170 3750 -1950 3784
rect -1712 3750 -1492 3784
rect -1254 3750 -1034 3784
rect -796 3750 -576 3784
rect -338 3750 -118 3784
rect 540 3750 760 3784
rect 998 3750 1218 3784
rect 1456 3750 1676 3784
rect 1914 3750 2134 3784
rect 2372 3750 2592 3784
rect 2830 3750 3050 3784
rect 3288 3750 3508 3784
rect 3746 3750 3966 3784
rect 4204 3750 4424 3784
rect 4662 3750 4882 3784
rect -4460 3440 -4240 3474
rect -4002 3440 -3782 3474
rect -3544 3440 -3324 3474
rect -3086 3440 -2866 3474
rect -2628 3440 -2408 3474
rect -2170 3440 -1950 3474
rect -1712 3440 -1492 3474
rect -1254 3440 -1034 3474
rect -796 3440 -576 3474
rect -338 3440 -118 3474
rect 540 3440 760 3474
rect 998 3440 1218 3474
rect 1456 3440 1676 3474
rect 1914 3440 2134 3474
rect 2372 3440 2592 3474
rect 2830 3440 3050 3474
rect 3288 3440 3508 3474
rect 3746 3440 3966 3474
rect 4204 3440 4424 3474
rect 4662 3440 4882 3474
rect -4460 3082 -4240 3116
rect -4002 3082 -3782 3116
rect -3544 3082 -3324 3116
rect -3086 3082 -2866 3116
rect -2628 3082 -2408 3116
rect -2170 3082 -1950 3116
rect -1712 3082 -1492 3116
rect -1254 3082 -1034 3116
rect -796 3082 -576 3116
rect -338 3082 -118 3116
rect -4460 2772 -4240 2806
rect -4002 2772 -3782 2806
rect -3544 2772 -3324 2806
rect -3086 2772 -2866 2806
rect -2628 2772 -2408 2806
rect -2170 2772 -1950 2806
rect -1712 2772 -1492 2806
rect -1254 2772 -1034 2806
rect -796 2772 -576 2806
rect -338 2772 -118 2806
<< locali >>
rect -5022 10160 -4922 10322
rect 5322 10160 5422 10322
rect -3916 8917 -3900 8951
rect -3680 8917 -3664 8951
rect -3458 8917 -3442 8951
rect -3222 8917 -3206 8951
rect -3000 8917 -2984 8951
rect -2764 8917 -2748 8951
rect -2542 8917 -2526 8951
rect -2306 8917 -2290 8951
rect -2084 8917 -2068 8951
rect -1848 8917 -1832 8951
rect -1626 8917 -1610 8951
rect -1390 8917 -1374 8951
rect -1168 8917 -1152 8951
rect -932 8917 -916 8951
rect -710 8917 -694 8951
rect -474 8917 -458 8951
rect -252 8917 -236 8951
rect -16 8917 0 8951
rect 206 8917 222 8951
rect 442 8917 458 8951
rect 664 8917 680 8951
rect 900 8917 916 8951
rect 1122 8917 1138 8951
rect 1358 8917 1374 8951
rect 1580 8917 1596 8951
rect 1816 8917 1832 8951
rect 2038 8917 2054 8951
rect 2274 8917 2290 8951
rect 2496 8917 2512 8951
rect 2732 8917 2748 8951
rect 2954 8917 2970 8951
rect 3190 8917 3206 8951
rect 3412 8917 3428 8951
rect 3648 8917 3664 8951
rect 3870 8917 3886 8951
rect 4106 8917 4122 8951
rect -4036 8858 -4002 8874
rect -4036 7266 -4002 7282
rect -3578 8858 -3544 8874
rect -3578 7266 -3544 7282
rect -3120 8858 -3086 8874
rect -3120 7266 -3086 7282
rect -2662 8858 -2628 8874
rect -2662 7266 -2628 7282
rect -2204 8858 -2170 8874
rect -2204 7266 -2170 7282
rect -1746 8858 -1712 8874
rect -1746 7266 -1712 7282
rect -1288 8858 -1254 8874
rect -1288 7266 -1254 7282
rect -830 8858 -796 8874
rect -830 7266 -796 7282
rect -372 8858 -338 8874
rect -372 7266 -338 7282
rect 86 8858 120 8874
rect 86 7266 120 7282
rect 544 8858 578 8874
rect 544 7266 578 7282
rect 1002 8858 1036 8874
rect 1002 7266 1036 7282
rect 1460 8858 1494 8874
rect 1460 7266 1494 7282
rect 1918 8858 1952 8874
rect 1918 7266 1952 7282
rect 2376 8858 2410 8874
rect 2376 7266 2410 7282
rect 2834 8858 2868 8874
rect 2834 7266 2868 7282
rect 3292 8858 3326 8874
rect 3292 7266 3326 7282
rect 3750 8858 3784 8874
rect 3750 7266 3784 7282
rect 4208 8858 4242 8874
rect 4208 7266 4242 7282
rect -3916 7189 -3900 7223
rect -3680 7189 -3664 7223
rect -3458 7189 -3442 7223
rect -3222 7189 -3206 7223
rect -3000 7189 -2984 7223
rect -2764 7189 -2748 7223
rect -2542 7189 -2526 7223
rect -2306 7189 -2290 7223
rect -2084 7189 -2068 7223
rect -1848 7189 -1832 7223
rect -1626 7189 -1610 7223
rect -1390 7189 -1374 7223
rect -1168 7189 -1152 7223
rect -932 7189 -916 7223
rect -710 7189 -694 7223
rect -474 7189 -458 7223
rect -252 7189 -236 7223
rect -16 7189 0 7223
rect 206 7189 222 7223
rect 442 7189 458 7223
rect 664 7189 680 7223
rect 900 7189 916 7223
rect 1122 7189 1138 7223
rect 1358 7189 1374 7223
rect 1580 7189 1596 7223
rect 1816 7189 1832 7223
rect 2038 7189 2054 7223
rect 2274 7189 2290 7223
rect 2496 7189 2512 7223
rect 2732 7189 2748 7223
rect 2954 7189 2970 7223
rect 3190 7189 3206 7223
rect 3412 7189 3428 7223
rect 3648 7189 3664 7223
rect 3870 7189 3886 7223
rect 4106 7189 4122 7223
rect -158 7106 302 7112
rect -158 7058 -152 7106
rect -104 7058 302 7106
rect -158 7052 302 7058
rect -4475 6252 -4459 6286
rect -4239 6252 -4223 6286
rect -4017 6252 -4001 6286
rect -3781 6252 -3765 6286
rect -3559 6252 -3543 6286
rect -3323 6252 -3307 6286
rect -3101 6252 -3085 6286
rect -2865 6252 -2849 6286
rect -2643 6252 -2627 6286
rect -2407 6252 -2391 6286
rect -2185 6252 -2169 6286
rect -1949 6252 -1933 6286
rect -1727 6252 -1711 6286
rect -1491 6252 -1475 6286
rect -1269 6252 -1253 6286
rect -1033 6252 -1017 6286
rect -811 6252 -795 6286
rect -575 6252 -559 6286
rect -353 6252 -337 6286
rect -117 6252 -101 6286
rect 525 6252 541 6286
rect 761 6252 777 6286
rect 983 6252 999 6286
rect 1219 6252 1235 6286
rect 1441 6252 1457 6286
rect 1677 6252 1693 6286
rect 1899 6252 1915 6286
rect 2135 6252 2151 6286
rect 2357 6252 2373 6286
rect 2593 6252 2609 6286
rect 2815 6252 2831 6286
rect 3051 6252 3067 6286
rect 3273 6252 3289 6286
rect 3509 6252 3525 6286
rect 3731 6252 3747 6286
rect 3967 6252 3983 6286
rect 4189 6252 4205 6286
rect 4425 6252 4441 6286
rect 4647 6252 4663 6286
rect 4883 6252 4899 6286
rect -4595 6193 -4561 6209
rect -4595 5001 -4561 5017
rect -4137 6193 -4103 6209
rect -4137 5001 -4103 5017
rect -3679 6193 -3645 6209
rect -3679 5001 -3645 5017
rect -3221 6193 -3187 6209
rect -3221 5001 -3187 5017
rect -2763 6193 -2729 6209
rect -2763 5001 -2729 5017
rect -2305 6193 -2271 6209
rect -2305 5001 -2271 5017
rect -1847 6193 -1813 6209
rect -1847 5001 -1813 5017
rect -1389 6193 -1355 6209
rect -1389 5001 -1355 5017
rect -931 6193 -897 6209
rect -931 5001 -897 5017
rect -473 6193 -439 6209
rect -473 5001 -439 5017
rect -15 6193 19 6209
rect -15 5001 19 5017
rect 405 6193 439 6209
rect 405 5001 439 5017
rect 863 6193 897 6209
rect 863 5001 897 5017
rect 1321 6193 1355 6209
rect 1321 5001 1355 5017
rect 1779 6193 1813 6209
rect 1779 5001 1813 5017
rect 2237 6193 2271 6209
rect 2237 5001 2271 5017
rect 2695 6193 2729 6209
rect 2695 5001 2729 5017
rect 3153 6193 3187 6209
rect 3153 5001 3187 5017
rect 3611 6193 3645 6209
rect 3611 5001 3645 5017
rect 4069 6193 4103 6209
rect 4069 5001 4103 5017
rect 4527 6193 4561 6209
rect 4527 5001 4561 5017
rect 4985 6193 5019 6209
rect 4985 5001 5019 5017
rect -4475 4924 -4459 4958
rect -4239 4924 -4223 4958
rect -4017 4924 -4001 4958
rect -3781 4924 -3765 4958
rect -3559 4924 -3543 4958
rect -3323 4924 -3307 4958
rect -3101 4924 -3085 4958
rect -2865 4924 -2849 4958
rect -2643 4924 -2627 4958
rect -2407 4924 -2391 4958
rect -2185 4924 -2169 4958
rect -1949 4924 -1933 4958
rect -1727 4924 -1711 4958
rect -1491 4924 -1475 4958
rect -1269 4924 -1253 4958
rect -1033 4924 -1017 4958
rect -811 4924 -795 4958
rect -575 4924 -559 4958
rect -353 4924 -337 4958
rect -117 4924 -101 4958
rect 525 4924 541 4958
rect 761 4924 777 4958
rect 983 4924 999 4958
rect 1219 4924 1235 4958
rect 1441 4924 1457 4958
rect 1677 4924 1693 4958
rect 1899 4924 1915 4958
rect 2135 4924 2151 4958
rect 2357 4924 2373 4958
rect 2593 4924 2609 4958
rect 2815 4924 2831 4958
rect 3051 4924 3067 4958
rect 3273 4924 3289 4958
rect 3509 4924 3525 4958
rect 3731 4924 3747 4958
rect 3967 4924 3983 4958
rect 4189 4924 4205 4958
rect 4425 4924 4441 4958
rect 4647 4924 4663 4958
rect 4883 4924 4899 4958
rect -5022 4478 -4922 4640
rect 5322 4478 5422 4640
rect -5022 4080 -4922 4242
rect 5322 4080 5422 4242
rect -4476 3750 -4460 3784
rect -4240 3750 -4224 3784
rect -4018 3750 -4002 3784
rect -3782 3750 -3766 3784
rect -3560 3750 -3544 3784
rect -3324 3750 -3308 3784
rect -3102 3750 -3086 3784
rect -2866 3750 -2850 3784
rect -2644 3750 -2628 3784
rect -2408 3750 -2392 3784
rect -2186 3750 -2170 3784
rect -1950 3750 -1934 3784
rect -1728 3750 -1712 3784
rect -1492 3750 -1476 3784
rect -1270 3750 -1254 3784
rect -1034 3750 -1018 3784
rect -812 3750 -796 3784
rect -576 3750 -560 3784
rect -354 3750 -338 3784
rect -118 3750 -102 3784
rect 524 3750 540 3784
rect 760 3750 776 3784
rect 982 3750 998 3784
rect 1218 3750 1234 3784
rect 1440 3750 1456 3784
rect 1676 3750 1692 3784
rect 1898 3750 1914 3784
rect 2134 3750 2150 3784
rect 2356 3750 2372 3784
rect 2592 3750 2608 3784
rect 2814 3750 2830 3784
rect 3050 3750 3066 3784
rect 3272 3750 3288 3784
rect 3508 3750 3524 3784
rect 3730 3750 3746 3784
rect 3966 3750 3982 3784
rect 4188 3750 4204 3784
rect 4424 3750 4440 3784
rect 4646 3750 4662 3784
rect 4882 3750 4898 3784
rect -4596 3700 -4562 3716
rect -4596 3508 -4562 3524
rect -4138 3700 -4104 3716
rect -4138 3508 -4104 3524
rect -3680 3700 -3646 3716
rect -3680 3508 -3646 3524
rect -3222 3700 -3188 3716
rect -3222 3508 -3188 3524
rect -2764 3700 -2730 3716
rect -2764 3508 -2730 3524
rect -2306 3700 -2272 3716
rect -2306 3508 -2272 3524
rect -1848 3700 -1814 3716
rect -1848 3508 -1814 3524
rect -1390 3700 -1356 3716
rect -1390 3508 -1356 3524
rect -932 3700 -898 3716
rect -932 3508 -898 3524
rect -474 3700 -440 3716
rect -474 3508 -440 3524
rect -16 3700 18 3716
rect -16 3508 18 3524
rect 404 3700 438 3716
rect 404 3508 438 3524
rect 862 3700 896 3716
rect 862 3508 896 3524
rect 1320 3700 1354 3716
rect 1320 3508 1354 3524
rect 1778 3700 1812 3716
rect 1778 3508 1812 3524
rect 2236 3700 2270 3716
rect 2236 3508 2270 3524
rect 2694 3700 2728 3716
rect 2694 3508 2728 3524
rect 3152 3700 3186 3716
rect 3152 3508 3186 3524
rect 3610 3700 3644 3716
rect 3610 3508 3644 3524
rect 4068 3700 4102 3716
rect 4068 3508 4102 3524
rect 4526 3700 4560 3716
rect 4526 3508 4560 3524
rect 4984 3700 5018 3716
rect 4984 3508 5018 3524
rect -4476 3440 -4460 3474
rect -4240 3440 -4224 3474
rect -4018 3440 -4002 3474
rect -3782 3440 -3766 3474
rect -3560 3440 -3544 3474
rect -3324 3440 -3308 3474
rect -3102 3440 -3086 3474
rect -2866 3440 -2850 3474
rect -2644 3440 -2628 3474
rect -2408 3440 -2392 3474
rect -2186 3440 -2170 3474
rect -1950 3440 -1934 3474
rect -1728 3440 -1712 3474
rect -1492 3440 -1476 3474
rect -1270 3440 -1254 3474
rect -1034 3440 -1018 3474
rect -812 3440 -796 3474
rect -576 3440 -560 3474
rect -354 3440 -338 3474
rect -118 3440 -102 3474
rect 524 3440 540 3474
rect 760 3440 776 3474
rect 982 3440 998 3474
rect 1218 3440 1234 3474
rect 1440 3440 1456 3474
rect 1676 3440 1692 3474
rect 1898 3440 1914 3474
rect 2134 3440 2150 3474
rect 2356 3440 2372 3474
rect 2592 3440 2608 3474
rect 2814 3440 2830 3474
rect 3050 3440 3066 3474
rect 3272 3440 3288 3474
rect 3508 3440 3524 3474
rect 3730 3440 3746 3474
rect 3966 3440 3982 3474
rect 4188 3440 4204 3474
rect 4424 3440 4440 3474
rect 4646 3440 4662 3474
rect 4882 3440 4898 3474
rect -4476 3082 -4460 3116
rect -4240 3082 -4224 3116
rect -4018 3082 -4002 3116
rect -3782 3082 -3766 3116
rect -3560 3082 -3544 3116
rect -3324 3082 -3308 3116
rect -3102 3082 -3086 3116
rect -2866 3082 -2850 3116
rect -2644 3082 -2628 3116
rect -2408 3082 -2392 3116
rect -2186 3082 -2170 3116
rect -1950 3082 -1934 3116
rect -1728 3082 -1712 3116
rect -1492 3082 -1476 3116
rect -1270 3082 -1254 3116
rect -1034 3082 -1018 3116
rect -812 3082 -796 3116
rect -576 3082 -560 3116
rect -354 3082 -338 3116
rect -118 3082 -102 3116
rect -4596 3032 -4562 3048
rect -4596 2840 -4562 2856
rect -4138 3032 -4104 3048
rect -4138 2840 -4104 2856
rect -3680 3032 -3646 3048
rect -3680 2840 -3646 2856
rect -3222 3032 -3188 3048
rect -3222 2840 -3188 2856
rect -2764 3032 -2730 3048
rect -2764 2840 -2730 2856
rect -2306 3032 -2272 3048
rect -2306 2840 -2272 2856
rect -1848 3032 -1814 3048
rect -1848 2840 -1814 2856
rect -1390 3032 -1356 3048
rect -1390 2840 -1356 2856
rect -932 3032 -898 3048
rect -932 2840 -898 2856
rect -474 3032 -440 3048
rect -474 2840 -440 2856
rect -16 3032 18 3048
rect -16 2840 18 2856
rect -4476 2772 -4460 2806
rect -4240 2772 -4224 2806
rect -4018 2772 -4002 2806
rect -3782 2772 -3766 2806
rect -3560 2772 -3544 2806
rect -3324 2772 -3308 2806
rect -3102 2772 -3086 2806
rect -2866 2772 -2850 2806
rect -2644 2772 -2628 2806
rect -2408 2772 -2392 2806
rect -2186 2772 -2170 2806
rect -1950 2772 -1934 2806
rect -1728 2772 -1712 2806
rect -1492 2772 -1476 2806
rect -1270 2772 -1254 2806
rect -1034 2772 -1018 2806
rect -812 2772 -796 2806
rect -576 2772 -560 2806
rect -354 2772 -338 2806
rect -118 2772 -102 2806
rect -5022 1778 -4922 1940
rect 5322 1778 5422 1940
<< viali >>
rect -4922 10222 -4860 10322
rect -4860 10222 5260 10322
rect 5260 10222 5322 10322
rect -5022 4760 -4922 9932
rect -3882 8917 -3698 8951
rect -3424 8917 -3240 8951
rect -2966 8917 -2782 8951
rect -2508 8917 -2324 8951
rect -2050 8917 -1866 8951
rect -1592 8917 -1408 8951
rect -1134 8917 -950 8951
rect -676 8917 -492 8951
rect -218 8917 -34 8951
rect 240 8917 424 8951
rect 698 8917 882 8951
rect 1156 8917 1340 8951
rect 1614 8917 1798 8951
rect 2072 8917 2256 8951
rect 2530 8917 2714 8951
rect 2988 8917 3172 8951
rect 3446 8917 3630 8951
rect 3904 8917 4088 8951
rect -4036 7282 -4002 8858
rect -3578 7282 -3544 8858
rect -3120 7282 -3086 8858
rect -2662 7282 -2628 8858
rect -2204 7282 -2170 8858
rect -1746 7282 -1712 8858
rect -1288 7282 -1254 8858
rect -830 7282 -796 8858
rect -372 7282 -338 8858
rect 86 7282 120 8858
rect 544 7282 578 8858
rect 1002 7282 1036 8858
rect 1460 7282 1494 8858
rect 1918 7282 1952 8858
rect 2376 7282 2410 8858
rect 2834 7282 2868 8858
rect 3292 7282 3326 8858
rect 3750 7282 3784 8858
rect 4208 7282 4242 8858
rect -3882 7189 -3698 7223
rect -3424 7189 -3240 7223
rect -2966 7189 -2782 7223
rect -2508 7189 -2324 7223
rect -2050 7189 -1866 7223
rect -1592 7189 -1408 7223
rect -1134 7189 -950 7223
rect -676 7189 -492 7223
rect -218 7189 -34 7223
rect 240 7189 424 7223
rect 698 7189 882 7223
rect 1156 7189 1340 7223
rect 1614 7189 1798 7223
rect 2072 7189 2256 7223
rect 2530 7189 2714 7223
rect 2988 7189 3172 7223
rect 3446 7189 3630 7223
rect 3904 7189 4088 7223
rect -152 7058 -104 7106
rect 302 7052 362 7112
rect -4441 6252 -4257 6286
rect -3983 6252 -3799 6286
rect -3525 6252 -3341 6286
rect -3067 6252 -2883 6286
rect -2609 6252 -2425 6286
rect -2151 6252 -1967 6286
rect -1693 6252 -1509 6286
rect -1235 6252 -1051 6286
rect -777 6252 -593 6286
rect -319 6252 -135 6286
rect 559 6252 743 6286
rect 1017 6252 1201 6286
rect 1475 6252 1659 6286
rect 1933 6252 2117 6286
rect 2391 6252 2575 6286
rect 2849 6252 3033 6286
rect 3307 6252 3491 6286
rect 3765 6252 3949 6286
rect 4223 6252 4407 6286
rect 4681 6252 4865 6286
rect -4595 5017 -4561 6193
rect -4137 5017 -4103 6193
rect -3679 5017 -3645 6193
rect -3221 5017 -3187 6193
rect -2763 5017 -2729 6193
rect -2305 5017 -2271 6193
rect -1847 5017 -1813 6193
rect -1389 5017 -1355 6193
rect -931 5017 -897 6193
rect -473 5017 -439 6193
rect -15 5017 19 6193
rect 405 5017 439 6193
rect 863 5017 897 6193
rect 1321 5017 1355 6193
rect 1779 5017 1813 6193
rect 2237 5017 2271 6193
rect 2695 5017 2729 6193
rect 3153 5017 3187 6193
rect 3611 5017 3645 6193
rect 4069 5017 4103 6193
rect 4527 5017 4561 6193
rect 4985 5017 5019 6193
rect -4441 4924 -4257 4958
rect -3983 4924 -3799 4958
rect -3525 4924 -3341 4958
rect -3067 4924 -2883 4958
rect -2609 4924 -2425 4958
rect -2151 4924 -1967 4958
rect -1693 4924 -1509 4958
rect -1235 4924 -1051 4958
rect -777 4924 -593 4958
rect -319 4924 -135 4958
rect 559 4924 743 4958
rect 1017 4924 1201 4958
rect 1475 4924 1659 4958
rect 1933 4924 2117 4958
rect 2391 4924 2575 4958
rect 2849 4924 3033 4958
rect 3307 4924 3491 4958
rect 3765 4924 3949 4958
rect 4223 4924 4407 4958
rect 4681 4924 4865 4958
rect 5322 4760 5422 9932
rect -4922 4478 -4860 4578
rect -4860 4478 5260 4578
rect 5260 4478 5322 4578
rect -4922 4142 -4860 4242
rect -4860 4142 5260 4242
rect 5260 4142 5322 4242
rect -5022 2008 -4922 4012
rect -4442 3750 -4258 3784
rect -3984 3750 -3800 3784
rect -3526 3750 -3342 3784
rect -3068 3750 -2884 3784
rect -2610 3750 -2426 3784
rect -2152 3750 -1968 3784
rect -1694 3750 -1510 3784
rect -1236 3750 -1052 3784
rect -778 3750 -594 3784
rect -320 3750 -136 3784
rect 558 3750 742 3784
rect 1016 3750 1200 3784
rect 1474 3750 1658 3784
rect 1932 3750 2116 3784
rect 2390 3750 2574 3784
rect 2848 3750 3032 3784
rect 3306 3750 3490 3784
rect 3764 3750 3948 3784
rect 4222 3750 4406 3784
rect 4680 3750 4864 3784
rect -4596 3524 -4562 3700
rect -4138 3524 -4104 3700
rect -3680 3524 -3646 3700
rect -3222 3524 -3188 3700
rect -2764 3524 -2730 3700
rect -2306 3524 -2272 3700
rect -1848 3524 -1814 3700
rect -1390 3524 -1356 3700
rect -932 3524 -898 3700
rect -474 3524 -440 3700
rect -16 3524 18 3700
rect 404 3524 438 3700
rect 862 3524 896 3700
rect 1320 3524 1354 3700
rect 1778 3524 1812 3700
rect 2236 3524 2270 3700
rect 2694 3524 2728 3700
rect 3152 3524 3186 3700
rect 3610 3524 3644 3700
rect 4068 3524 4102 3700
rect 4526 3524 4560 3700
rect 4984 3524 5018 3700
rect -4442 3440 -4258 3474
rect -3984 3440 -3800 3474
rect -3526 3440 -3342 3474
rect -3068 3440 -2884 3474
rect -2610 3440 -2426 3474
rect -2152 3440 -1968 3474
rect -1694 3440 -1510 3474
rect -1236 3440 -1052 3474
rect -778 3440 -594 3474
rect -320 3440 -136 3474
rect 558 3440 742 3474
rect 1016 3440 1200 3474
rect 1474 3440 1658 3474
rect 1932 3440 2116 3474
rect 2390 3440 2574 3474
rect 2848 3440 3032 3474
rect 3306 3440 3490 3474
rect 3764 3440 3948 3474
rect 4222 3440 4406 3474
rect 4680 3440 4864 3474
rect -4442 3082 -4258 3116
rect -3984 3082 -3800 3116
rect -3526 3082 -3342 3116
rect -3068 3082 -2884 3116
rect -2610 3082 -2426 3116
rect -2152 3082 -1968 3116
rect -1694 3082 -1510 3116
rect -1236 3082 -1052 3116
rect -778 3082 -594 3116
rect -320 3082 -136 3116
rect -4596 2856 -4562 3032
rect -4138 2856 -4104 3032
rect -3680 2856 -3646 3032
rect -3222 2856 -3188 3032
rect -2764 2856 -2730 3032
rect -2306 2856 -2272 3032
rect -1848 2856 -1814 3032
rect -1390 2856 -1356 3032
rect -932 2856 -898 3032
rect -474 2856 -440 3032
rect -16 2856 18 3032
rect -4442 2772 -4258 2806
rect -3984 2772 -3800 2806
rect -3526 2772 -3342 2806
rect -3068 2772 -2884 2806
rect -2610 2772 -2426 2806
rect -2152 2772 -1968 2806
rect -1694 2772 -1510 2806
rect -1236 2772 -1052 2806
rect -778 2772 -594 2806
rect -320 2772 -136 2806
rect 5322 2008 5422 4012
rect -4922 1778 -4860 1878
rect -4860 1778 5260 1878
rect 5260 1778 5322 1878
<< metal1 >>
rect -5028 10322 5428 10328
rect -5028 10222 -4922 10322
rect 5322 10222 5428 10322
rect -5028 10216 5428 10222
rect -5028 9932 -4916 10216
rect -5028 4760 -5022 9932
rect -4922 7110 -4916 9932
rect -4316 9916 -4306 10216
rect 4706 9916 4716 10216
rect 5316 9932 5428 10216
rect -4078 9742 4278 9756
rect -4078 9656 -4064 9742
rect -3968 9656 -3464 9742
rect -3368 9656 -2864 9742
rect -2768 9656 -2264 9742
rect -2168 9656 -1664 9742
rect -1568 9656 -1064 9742
rect -968 9656 -464 9742
rect -368 9656 136 9742
rect 232 9656 736 9742
rect 832 9656 1336 9742
rect 1432 9656 1936 9742
rect 2032 9656 2536 9742
rect 2632 9656 3136 9742
rect 3232 9656 3736 9742
rect 3832 9656 4156 9742
rect 4252 9656 4278 9742
rect -4078 9646 4278 9656
rect -4050 8858 -3990 9646
rect -3818 8957 -3758 9646
rect -3894 8951 -3686 8957
rect -3894 8917 -3882 8951
rect -3698 8917 -3686 8951
rect -3894 8911 -3686 8917
rect -4050 8826 -4036 8858
rect -4042 7342 -4036 8826
rect -4048 7282 -4036 7342
rect -4002 8826 -3990 8858
rect -3592 8858 -3532 9646
rect -2676 9392 2882 9452
rect -3366 9024 -3360 9084
rect -3300 9024 -3294 9084
rect -2910 9024 -2904 9084
rect -2844 9024 -2838 9084
rect -3360 8957 -3300 9024
rect -2904 8957 -2844 9024
rect -3436 8951 -3228 8957
rect -3436 8917 -3424 8951
rect -3240 8917 -3228 8951
rect -3436 8911 -3228 8917
rect -2978 8951 -2770 8957
rect -2978 8917 -2966 8951
rect -2782 8917 -2770 8951
rect -2978 8911 -2770 8917
rect -4002 7342 -3996 8826
rect -3592 8794 -3578 8858
rect -4002 7282 -3988 7342
rect -3584 7326 -3578 8794
rect -4048 7110 -3988 7282
rect -3594 7282 -3578 7326
rect -3544 8794 -3532 8858
rect -3126 8858 -3080 8870
rect -3544 7326 -3538 8794
rect -3126 7366 -3120 8858
rect -3544 7282 -3534 7326
rect -3894 7223 -3686 7229
rect -3894 7189 -3882 7223
rect -3698 7189 -3686 7223
rect -3894 7183 -3686 7189
rect -3820 7110 -3760 7183
rect -3594 7110 -3534 7282
rect -3136 7282 -3120 7366
rect -3086 7366 -3080 8858
rect -2676 8858 -2616 9392
rect -1760 9258 1962 9318
rect -2450 9024 -2444 9084
rect -2384 9024 -2378 9084
rect -1994 9024 -1988 9084
rect -1928 9024 -1922 9084
rect -2444 8957 -2384 9024
rect -1988 8957 -1928 9024
rect -2520 8951 -2312 8957
rect -2520 8917 -2508 8951
rect -2324 8917 -2312 8951
rect -2520 8911 -2312 8917
rect -2062 8951 -1854 8957
rect -2062 8917 -2050 8951
rect -1866 8917 -1854 8951
rect -2062 8911 -1854 8917
rect -2676 8800 -2662 8858
rect -3086 7282 -3076 7366
rect -3436 7223 -3228 7229
rect -3436 7189 -3424 7223
rect -3240 7189 -3228 7223
rect -3436 7183 -3228 7189
rect -3364 7110 -3304 7183
rect -4922 7050 -3534 7110
rect -3370 7050 -3364 7110
rect -3304 7050 -3298 7110
rect -4922 6678 -4916 7050
rect -4048 6678 -3988 7050
rect -4922 6618 -3988 6678
rect -3136 6630 -3076 7282
rect -2668 7282 -2662 8800
rect -2628 8800 -2616 8858
rect -2210 8858 -2164 8870
rect -2628 7282 -2622 8800
rect -2210 7360 -2204 8858
rect -2668 7270 -2622 7282
rect -2218 7282 -2204 7360
rect -2170 7360 -2164 8858
rect -1760 8858 -1700 9258
rect -844 9134 1046 9194
rect -1536 9024 -1530 9084
rect -1470 9024 -1464 9084
rect -1072 9024 -1066 9084
rect -1006 9024 -1000 9084
rect -1530 8957 -1470 9024
rect -1066 8957 -1006 9024
rect -1604 8951 -1396 8957
rect -1604 8917 -1592 8951
rect -1408 8917 -1396 8951
rect -1604 8911 -1396 8917
rect -1146 8951 -938 8957
rect -1146 8917 -1134 8951
rect -950 8917 -938 8951
rect -1146 8911 -938 8917
rect -1760 8798 -1746 8858
rect -2170 7282 -2158 7360
rect -2978 7223 -2770 7229
rect -2978 7189 -2966 7223
rect -2782 7189 -2770 7223
rect -2978 7183 -2770 7189
rect -2520 7223 -2312 7229
rect -2520 7189 -2508 7223
rect -2324 7189 -2312 7223
rect -2520 7183 -2312 7189
rect -2908 7110 -2848 7183
rect -2448 7110 -2388 7183
rect -2914 7050 -2908 7110
rect -2848 7050 -2842 7110
rect -2454 7050 -2448 7110
rect -2388 7050 -2382 7110
rect -2218 6760 -2158 7282
rect -1752 7282 -1746 8798
rect -1712 8798 -1700 8858
rect -1294 8858 -1248 8870
rect -1712 7282 -1706 8798
rect -1294 7354 -1288 8858
rect -1752 7270 -1706 7282
rect -1310 7282 -1288 7354
rect -1254 7282 -1248 8858
rect -844 8858 -784 9134
rect -622 9024 -616 9084
rect -556 9024 -550 9084
rect -166 9024 -160 9084
rect -100 9024 -94 9084
rect 302 9024 308 9084
rect 368 9024 374 9084
rect 760 9024 766 9084
rect 826 9024 832 9084
rect -616 8957 -556 9024
rect -160 8957 -100 9024
rect 308 8957 368 9024
rect 766 8957 826 9024
rect -688 8951 -480 8957
rect -688 8917 -676 8951
rect -492 8917 -480 8951
rect -688 8911 -480 8917
rect -230 8951 -22 8957
rect -230 8917 -218 8951
rect -34 8917 -22 8951
rect -230 8911 -22 8917
rect 228 8951 436 8957
rect 228 8917 240 8951
rect 424 8917 436 8951
rect 228 8911 436 8917
rect 686 8951 894 8957
rect 686 8917 698 8951
rect 882 8917 894 8951
rect 686 8911 894 8917
rect -844 8780 -830 8858
rect -1310 7270 -1248 7282
rect -836 7282 -830 8780
rect -796 8780 -784 8858
rect -378 8858 -332 8870
rect -796 7282 -790 8780
rect -378 7362 -372 8858
rect -836 7270 -790 7282
rect -386 7282 -372 7362
rect -338 7362 -332 8858
rect 80 8858 126 8870
rect -338 7282 -326 7362
rect 80 7304 86 8858
rect -2062 7223 -1854 7229
rect -2062 7189 -2050 7223
rect -1866 7189 -1854 7223
rect -2062 7183 -1854 7189
rect -1604 7223 -1396 7229
rect -1604 7189 -1592 7223
rect -1408 7189 -1396 7223
rect -1604 7183 -1396 7189
rect -1992 7110 -1932 7183
rect -1534 7110 -1474 7183
rect -1998 7050 -1992 7110
rect -1932 7050 -1926 7110
rect -1540 7050 -1534 7110
rect -1474 7050 -1468 7110
rect -1310 6886 -1250 7270
rect -1146 7223 -938 7229
rect -1146 7189 -1134 7223
rect -950 7189 -938 7223
rect -1146 7183 -938 7189
rect -688 7223 -480 7229
rect -688 7189 -676 7223
rect -492 7189 -480 7223
rect -688 7183 -480 7189
rect -1070 7110 -1010 7183
rect -616 7110 -556 7183
rect -1076 7050 -1070 7110
rect -1010 7050 -1004 7110
rect -622 7050 -616 7110
rect -556 7050 -550 7110
rect -386 7002 -326 7282
rect 76 7282 86 7304
rect 120 7304 126 8858
rect 538 8858 584 8870
rect 538 7310 544 8858
rect 120 7282 136 7304
rect -230 7223 -22 7229
rect -230 7189 -218 7223
rect -34 7189 -22 7223
rect -230 7183 -22 7189
rect -158 7112 -98 7183
rect 76 7122 136 7282
rect 532 7282 544 7310
rect 578 7310 584 8858
rect 986 8858 1046 9134
rect 1216 9024 1222 9084
rect 1282 9024 1288 9084
rect 1672 9024 1678 9084
rect 1738 9024 1744 9084
rect 1222 8957 1282 9024
rect 1678 8957 1738 9024
rect 1144 8951 1352 8957
rect 1144 8917 1156 8951
rect 1340 8917 1352 8951
rect 1144 8911 1352 8917
rect 1602 8951 1810 8957
rect 1602 8917 1614 8951
rect 1798 8917 1810 8951
rect 1602 8911 1810 8917
rect 986 8814 1002 8858
rect 578 7282 592 7310
rect 228 7223 436 7229
rect 228 7189 240 7223
rect 424 7189 436 7223
rect 228 7183 436 7189
rect -164 7110 -92 7112
rect -164 7050 -158 7110
rect -98 7050 -92 7110
rect 302 7118 362 7183
rect 76 7056 136 7062
rect 290 7112 374 7118
rect 290 7050 302 7112
rect 362 7050 374 7112
rect 290 7046 374 7050
rect 532 7002 592 7282
rect 996 7282 1002 8814
rect 1036 8814 1046 8858
rect 1454 8858 1500 8870
rect 1036 7282 1042 8814
rect 1454 7314 1460 8858
rect 996 7270 1042 7282
rect 1446 7282 1460 7314
rect 1494 7314 1500 8858
rect 1902 8858 1962 9258
rect 2128 9024 2134 9084
rect 2194 9024 2200 9084
rect 2584 9024 2590 9084
rect 2650 9024 2656 9084
rect 2134 8957 2194 9024
rect 2590 8957 2650 9024
rect 2060 8951 2268 8957
rect 2060 8917 2072 8951
rect 2256 8917 2268 8951
rect 2060 8911 2268 8917
rect 2518 8951 2726 8957
rect 2518 8917 2530 8951
rect 2714 8917 2726 8951
rect 2518 8911 2726 8917
rect 1902 8800 1918 8858
rect 1494 7282 1506 7314
rect 686 7223 894 7229
rect 686 7189 698 7223
rect 882 7189 894 7223
rect 686 7183 894 7189
rect 1144 7223 1352 7229
rect 1144 7189 1156 7223
rect 1340 7189 1352 7223
rect 1144 7183 1352 7189
rect 758 7110 818 7183
rect 1218 7110 1278 7183
rect 752 7050 758 7110
rect 818 7050 824 7110
rect 1212 7050 1218 7110
rect 1278 7050 1284 7110
rect -386 6942 592 7002
rect 1446 6886 1506 7282
rect 1912 7282 1918 8800
rect 1952 8800 1962 8858
rect 2370 8858 2416 8870
rect 1952 7282 1958 8800
rect 2370 7350 2376 8858
rect 1912 7270 1958 7282
rect 2366 7282 2376 7350
rect 2410 7350 2416 8858
rect 2822 8858 2882 9392
rect 3042 9024 3048 9084
rect 3108 9024 3114 9084
rect 3502 9024 3508 9084
rect 3568 9024 3574 9084
rect 3048 8957 3108 9024
rect 3508 8957 3568 9024
rect 2976 8951 3184 8957
rect 2976 8917 2988 8951
rect 3172 8917 3184 8951
rect 2976 8911 3184 8917
rect 3434 8951 3642 8957
rect 3434 8917 3446 8951
rect 3630 8917 3642 8951
rect 3434 8911 3642 8917
rect 2822 8802 2834 8858
rect 2410 7282 2426 7350
rect 1602 7223 1810 7229
rect 1602 7189 1614 7223
rect 1798 7189 1810 7223
rect 1602 7183 1810 7189
rect 2060 7223 2268 7229
rect 2060 7189 2072 7223
rect 2256 7189 2268 7223
rect 2060 7183 2268 7189
rect 1674 7110 1734 7183
rect 2130 7110 2190 7183
rect 1668 7050 1674 7110
rect 1734 7050 1740 7110
rect 2124 7050 2130 7110
rect 2190 7050 2196 7110
rect -1310 6826 1506 6886
rect 2366 6760 2426 7282
rect 2828 7282 2834 8802
rect 2868 8802 2882 8858
rect 3286 8858 3332 8870
rect 2868 7282 2874 8802
rect 3286 7342 3292 8858
rect 2828 7270 2874 7282
rect 3280 7282 3292 7342
rect 3326 7342 3332 8858
rect 3738 8858 3798 9646
rect 3968 8957 4028 9646
rect 3892 8951 4100 8957
rect 3892 8917 3904 8951
rect 4088 8917 4100 8951
rect 3892 8911 4100 8917
rect 3738 8782 3750 8858
rect 3744 7344 3750 8782
rect 3326 7282 3340 7342
rect 2518 7223 2726 7229
rect 2518 7189 2530 7223
rect 2714 7189 2726 7223
rect 2518 7183 2726 7189
rect 2976 7223 3184 7229
rect 2976 7189 2988 7223
rect 3172 7189 3184 7223
rect 2976 7183 3184 7189
rect 2586 7110 2646 7183
rect 3044 7110 3104 7183
rect 2580 7050 2586 7110
rect 2646 7050 2652 7110
rect 3038 7050 3044 7110
rect 3104 7050 3110 7110
rect -2218 6700 2426 6760
rect 3280 6630 3340 7282
rect 3734 7282 3750 7344
rect 3784 8782 3798 8858
rect 4196 8858 4256 9646
rect 4196 8788 4208 8858
rect 3784 7344 3790 8782
rect 3784 7282 3794 7344
rect 4202 7326 4208 8788
rect 3434 7223 3642 7229
rect 3434 7189 3446 7223
rect 3630 7189 3642 7223
rect 3434 7183 3642 7189
rect 3504 7110 3564 7183
rect 3498 7050 3504 7110
rect 3564 7050 3570 7110
rect 3734 7108 3794 7282
rect 4192 7282 4208 7326
rect 4242 8788 4256 8858
rect 4242 7326 4248 8788
rect 4242 7282 4252 7326
rect 3892 7223 4100 7229
rect 3892 7189 3904 7223
rect 4088 7189 4100 7223
rect 3892 7183 4100 7189
rect 3966 7108 4026 7183
rect 4192 7108 4252 7282
rect 5316 7108 5322 9932
rect 3734 7048 5322 7108
rect -4922 4760 -4916 6618
rect -4608 6193 -4548 6618
rect -4380 6292 -4320 6618
rect -3136 6570 3340 6630
rect 4192 6614 4252 7048
rect 5316 6614 5322 7048
rect 4192 6554 5322 6614
rect -4156 6464 -4150 6524
rect -4090 6464 -4084 6524
rect -4453 6286 -4245 6292
rect -4453 6252 -4441 6286
rect -4257 6252 -4245 6286
rect -4453 6246 -4245 6252
rect -4608 6146 -4595 6193
rect -4601 5038 -4595 6146
rect -5028 4584 -4916 4760
rect -4608 5017 -4595 5038
rect -4561 6146 -4548 6193
rect -4150 6193 -4090 6464
rect -3918 6362 -654 6422
rect -3918 6292 -3858 6362
rect -3456 6292 -3396 6362
rect -3002 6292 -2942 6362
rect -2540 6292 -2480 6362
rect -2086 6292 -2026 6362
rect -1636 6292 -1576 6362
rect -1170 6292 -1110 6362
rect -714 6292 -654 6362
rect -258 6344 910 6404
rect -258 6292 -198 6344
rect -3995 6286 -3787 6292
rect -3995 6252 -3983 6286
rect -3799 6252 -3787 6286
rect -3995 6246 -3787 6252
rect -3537 6286 -3329 6292
rect -3537 6252 -3525 6286
rect -3341 6252 -3329 6286
rect -3537 6246 -3329 6252
rect -3079 6286 -2871 6292
rect -3079 6252 -3067 6286
rect -2883 6252 -2871 6286
rect -3079 6246 -2871 6252
rect -2621 6286 -2413 6292
rect -2621 6252 -2609 6286
rect -2425 6252 -2413 6286
rect -2621 6246 -2413 6252
rect -2163 6286 -1955 6292
rect -2163 6252 -2151 6286
rect -1967 6252 -1955 6286
rect -2163 6246 -1955 6252
rect -1705 6286 -1497 6292
rect -1705 6252 -1693 6286
rect -1509 6252 -1497 6286
rect -1705 6246 -1497 6252
rect -1247 6286 -1039 6292
rect -1247 6252 -1235 6286
rect -1051 6252 -1039 6286
rect -1247 6246 -1039 6252
rect -789 6286 -581 6292
rect -789 6252 -777 6286
rect -593 6252 -581 6286
rect -789 6246 -581 6252
rect -331 6286 -123 6292
rect -331 6252 -319 6286
rect -135 6252 -123 6286
rect -331 6246 -123 6252
rect -4561 5038 -4555 6146
rect -4150 6126 -4137 6193
rect -4561 5017 -4548 5038
rect -4608 4584 -4548 5017
rect -4143 5017 -4137 6126
rect -4103 6126 -4090 6193
rect -3685 6193 -3639 6205
rect -4103 5017 -4097 6126
rect -4143 5005 -4097 5017
rect -3685 5017 -3679 6193
rect -3645 5017 -3639 6193
rect -3685 5005 -3639 5017
rect -3227 6193 -3181 6205
rect -3227 5017 -3221 6193
rect -3187 5017 -3181 6193
rect -3227 5005 -3181 5017
rect -2769 6193 -2723 6205
rect -2769 5017 -2763 6193
rect -2729 5017 -2723 6193
rect -2769 5005 -2723 5017
rect -2311 6193 -2265 6205
rect -2311 5017 -2305 6193
rect -2271 5017 -2265 6193
rect -2311 5005 -2265 5017
rect -1853 6193 -1807 6205
rect -1853 5017 -1847 6193
rect -1813 5017 -1807 6193
rect -1853 5005 -1807 5017
rect -1395 6193 -1349 6205
rect -1395 5017 -1389 6193
rect -1355 5017 -1349 6193
rect -1395 5005 -1349 5017
rect -937 6193 -891 6205
rect -937 5017 -931 6193
rect -897 5017 -891 6193
rect -479 6193 -433 6205
rect -479 5084 -473 6193
rect -937 5005 -891 5017
rect -488 5017 -473 5084
rect -439 5084 -433 6193
rect -28 6193 32 6344
rect -28 6178 -15 6193
rect -439 5017 -428 5084
rect -21 5052 -15 6178
rect -4453 4958 -4245 4964
rect -4453 4924 -4441 4958
rect -4257 4924 -4245 4958
rect -4453 4918 -4245 4924
rect -3995 4958 -3787 4964
rect -3995 4924 -3983 4958
rect -3799 4924 -3787 4958
rect -3995 4918 -3787 4924
rect -3537 4958 -3329 4964
rect -3537 4924 -3525 4958
rect -3341 4924 -3329 4958
rect -3537 4918 -3329 4924
rect -3079 4958 -2871 4964
rect -3079 4924 -3067 4958
rect -2883 4924 -2871 4958
rect -3079 4918 -2871 4924
rect -2621 4958 -2413 4964
rect -2621 4924 -2609 4958
rect -2425 4924 -2413 4958
rect -2621 4918 -2413 4924
rect -2163 4958 -1955 4964
rect -2163 4924 -2151 4958
rect -1967 4924 -1955 4958
rect -2163 4918 -1955 4924
rect -1705 4958 -1497 4964
rect -1705 4924 -1693 4958
rect -1509 4924 -1497 4958
rect -1705 4918 -1497 4924
rect -1247 4958 -1039 4964
rect -1247 4924 -1235 4958
rect -1051 4924 -1039 4958
rect -1247 4918 -1039 4924
rect -789 4958 -581 4964
rect -789 4924 -777 4958
rect -593 4924 -581 4958
rect -789 4918 -581 4924
rect -4380 4584 -4320 4918
rect -3926 4850 -3866 4918
rect -3464 4850 -3404 4918
rect -3010 4850 -2950 4918
rect -2548 4850 -2488 4918
rect -2094 4850 -2034 4918
rect -1644 4850 -1584 4918
rect -1178 4850 -1118 4918
rect -722 4850 -662 4918
rect -3926 4846 -3010 4850
rect -3866 4790 -3464 4846
rect -3926 4780 -3866 4786
rect -3404 4790 -3010 4846
rect -2950 4790 -2548 4850
rect -2488 4844 -1644 4850
rect -2488 4790 -2094 4844
rect -3464 4780 -3404 4786
rect -3010 4784 -2950 4790
rect -2548 4784 -2488 4790
rect -2034 4790 -1644 4844
rect -1584 4790 -1178 4850
rect -1118 4846 -662 4850
rect -1118 4790 -722 4846
rect -1644 4784 -1584 4790
rect -1178 4784 -1118 4790
rect -2094 4778 -2034 4784
rect -722 4780 -662 4786
rect -488 4724 -428 5017
rect -30 5017 -15 5052
rect 19 6178 32 6193
rect 392 6193 452 6344
rect 624 6292 684 6344
rect 547 6286 755 6292
rect 547 6252 559 6286
rect 743 6252 755 6286
rect 547 6246 755 6252
rect 19 5052 25 6178
rect 392 6172 405 6193
rect 399 5052 405 6172
rect 19 5017 30 5052
rect -331 4958 -123 4964
rect -331 4924 -319 4958
rect -135 4924 -123 4958
rect -331 4918 -123 4924
rect -494 4664 -488 4724
rect -428 4664 -422 4724
rect -258 4584 -198 4918
rect -30 4584 30 5017
rect 390 5017 405 5052
rect 439 6172 452 6193
rect 850 6193 910 6344
rect 1076 6362 4340 6422
rect 1076 6292 1136 6362
rect 1538 6292 1598 6362
rect 1992 6292 2052 6362
rect 2454 6292 2514 6362
rect 2908 6292 2968 6362
rect 3358 6292 3418 6362
rect 3824 6292 3884 6362
rect 4280 6292 4340 6362
rect 4742 6292 4802 6554
rect 1005 6286 1213 6292
rect 1005 6252 1017 6286
rect 1201 6252 1213 6286
rect 1005 6246 1213 6252
rect 1463 6286 1671 6292
rect 1463 6252 1475 6286
rect 1659 6252 1671 6286
rect 1463 6246 1671 6252
rect 1921 6286 2129 6292
rect 1921 6252 1933 6286
rect 2117 6252 2129 6286
rect 1921 6246 2129 6252
rect 2379 6286 2587 6292
rect 2379 6252 2391 6286
rect 2575 6252 2587 6286
rect 2379 6246 2587 6252
rect 2837 6286 3045 6292
rect 2837 6252 2849 6286
rect 3033 6252 3045 6286
rect 2837 6246 3045 6252
rect 3295 6286 3503 6292
rect 3295 6252 3307 6286
rect 3491 6252 3503 6286
rect 3295 6246 3503 6252
rect 3753 6286 3961 6292
rect 3753 6252 3765 6286
rect 3949 6252 3961 6286
rect 3753 6246 3961 6252
rect 4211 6286 4419 6292
rect 4211 6252 4223 6286
rect 4407 6252 4419 6286
rect 4211 6246 4419 6252
rect 4669 6286 4877 6292
rect 4669 6252 4681 6286
rect 4865 6252 4877 6286
rect 4669 6246 4877 6252
rect 439 5052 445 6172
rect 850 6150 863 6193
rect 857 5058 863 6150
rect 439 5017 450 5052
rect 390 4584 450 5017
rect 848 5017 863 5058
rect 897 6150 910 6193
rect 1315 6193 1361 6205
rect 897 5058 903 6150
rect 897 5017 908 5058
rect 547 4958 755 4964
rect 547 4924 559 4958
rect 743 4924 755 4958
rect 547 4918 755 4924
rect 618 4584 678 4918
rect 848 4584 908 5017
rect 1315 5017 1321 6193
rect 1355 5017 1361 6193
rect 1315 5005 1361 5017
rect 1773 6193 1819 6205
rect 1773 5017 1779 6193
rect 1813 5017 1819 6193
rect 1773 5005 1819 5017
rect 2231 6193 2277 6205
rect 2231 5017 2237 6193
rect 2271 5017 2277 6193
rect 2231 5005 2277 5017
rect 2689 6193 2735 6205
rect 2689 5017 2695 6193
rect 2729 5017 2735 6193
rect 2689 5005 2735 5017
rect 3147 6193 3193 6205
rect 3147 5017 3153 6193
rect 3187 5017 3193 6193
rect 3147 5005 3193 5017
rect 3605 6193 3651 6205
rect 3605 5017 3611 6193
rect 3645 5017 3651 6193
rect 3605 5005 3651 5017
rect 4063 6193 4109 6205
rect 4063 5017 4069 6193
rect 4103 5017 4109 6193
rect 4521 6193 4567 6205
rect 4521 5024 4527 6193
rect 4063 5005 4109 5017
rect 4512 5017 4527 5024
rect 4561 5024 4567 6193
rect 4968 6193 5028 6554
rect 4968 6140 4985 6193
rect 4979 5050 4985 6140
rect 4561 5017 4572 5024
rect 1005 4958 1213 4964
rect 1005 4924 1017 4958
rect 1201 4924 1213 4958
rect 1005 4918 1213 4924
rect 1463 4958 1671 4964
rect 1463 4924 1475 4958
rect 1659 4924 1671 4958
rect 1463 4918 1671 4924
rect 1921 4958 2129 4964
rect 1921 4924 1933 4958
rect 2117 4924 2129 4958
rect 1921 4918 2129 4924
rect 2379 4958 2587 4964
rect 2379 4924 2391 4958
rect 2575 4924 2587 4958
rect 2379 4918 2587 4924
rect 2837 4958 3045 4964
rect 2837 4924 2849 4958
rect 3033 4924 3045 4958
rect 2837 4918 3045 4924
rect 3295 4958 3503 4964
rect 3295 4924 3307 4958
rect 3491 4924 3503 4958
rect 3295 4918 3503 4924
rect 3753 4958 3961 4964
rect 3753 4924 3765 4958
rect 3949 4924 3961 4958
rect 3753 4918 3961 4924
rect 4211 4958 4419 4964
rect 4211 4924 4223 4958
rect 4407 4924 4419 4958
rect 4211 4918 4419 4924
rect 1076 4850 1136 4918
rect 1538 4854 1598 4918
rect 1076 4846 1538 4850
rect 1136 4794 1538 4846
rect 1992 4850 2052 4918
rect 2454 4850 2514 4918
rect 2908 4850 2968 4918
rect 3358 4854 3418 4918
rect 1598 4848 3358 4850
rect 1598 4794 1992 4848
rect 1136 4790 1992 4794
rect 1538 4788 1598 4790
rect 2052 4790 2454 4848
rect 1076 4780 1136 4786
rect 1992 4782 2052 4788
rect 2514 4790 2908 4848
rect 2454 4782 2514 4788
rect 2968 4794 3358 4848
rect 3824 4850 3884 4918
rect 4280 4850 4340 4918
rect 3418 4848 4340 4850
rect 3418 4794 3824 4848
rect 2968 4790 3824 4794
rect 3358 4788 3418 4790
rect 3884 4790 4280 4848
rect 2908 4782 2968 4788
rect 3824 4782 3884 4788
rect 4280 4782 4340 4788
rect 4512 4718 4572 5017
rect 4970 5017 4985 5050
rect 5019 6140 5028 6193
rect 5019 5050 5025 6140
rect 5019 5017 5030 5050
rect 4669 4958 4877 4964
rect 4669 4924 4681 4958
rect 4865 4924 4877 4958
rect 4669 4918 4877 4924
rect 4512 4652 4572 4658
rect 4742 4584 4802 4918
rect 4970 4584 5030 5017
rect 5316 4760 5322 6554
rect 5422 4760 5428 9932
rect 5316 4584 5428 4760
rect -5028 4578 5428 4584
rect -5028 4478 -4922 4578
rect 5322 4478 5428 4578
rect -5028 4472 5428 4478
rect -5028 4242 5428 4248
rect -5028 4142 -4922 4242
rect 5322 4142 5428 4242
rect -5028 4136 5428 4142
rect -5028 4012 -4916 4136
rect -5028 2008 -5022 4012
rect -4922 2008 -4916 4012
rect -4608 3700 -4548 4136
rect -4378 3790 -4318 4136
rect -488 4044 -428 4050
rect -3920 3910 -3464 3916
rect -3932 3850 -3926 3910
rect -3866 3856 -3464 3910
rect -3404 3910 -2548 3916
rect -3404 3856 -3010 3910
rect -3866 3850 -3860 3856
rect -3926 3790 -3860 3850
rect -3464 3790 -3398 3856
rect -3016 3850 -3010 3856
rect -2950 3856 -2548 3910
rect -2488 3856 -2094 3916
rect -2034 3856 -1644 3916
rect -1584 3910 -722 3916
rect -1584 3856 -1178 3910
rect -2950 3850 -2944 3856
rect -3010 3790 -2944 3850
rect -2548 3790 -2482 3856
rect -2094 3790 -2028 3856
rect -1644 3790 -1578 3856
rect -1184 3850 -1178 3856
rect -1118 3856 -722 3910
rect -662 3856 -656 3916
rect -1118 3850 -1112 3856
rect -1178 3790 -1112 3850
rect -722 3790 -656 3856
rect -4454 3784 -4246 3790
rect -4454 3750 -4442 3784
rect -4258 3750 -4246 3784
rect -4454 3744 -4246 3750
rect -3996 3784 -3788 3790
rect -3996 3750 -3984 3784
rect -3800 3750 -3788 3784
rect -3996 3744 -3788 3750
rect -3538 3784 -3330 3790
rect -3538 3750 -3526 3784
rect -3342 3750 -3330 3784
rect -3538 3744 -3330 3750
rect -3080 3784 -2872 3790
rect -3080 3750 -3068 3784
rect -2884 3750 -2872 3784
rect -3080 3744 -2872 3750
rect -2622 3784 -2414 3790
rect -2622 3750 -2610 3784
rect -2426 3750 -2414 3784
rect -2622 3744 -2414 3750
rect -2164 3784 -1956 3790
rect -2164 3750 -2152 3784
rect -1968 3750 -1956 3784
rect -2164 3744 -1956 3750
rect -1706 3784 -1498 3790
rect -1706 3750 -1694 3784
rect -1510 3750 -1498 3784
rect -1706 3744 -1498 3750
rect -1248 3784 -1040 3790
rect -1248 3750 -1236 3784
rect -1052 3750 -1040 3784
rect -1248 3744 -1040 3750
rect -790 3784 -582 3790
rect -790 3750 -778 3784
rect -594 3750 -582 3784
rect -790 3744 -582 3750
rect -4608 3660 -4596 3700
rect -4602 3564 -4596 3660
rect -4608 3524 -4596 3564
rect -4562 3660 -4548 3700
rect -4144 3700 -4098 3712
rect -4562 3564 -4556 3660
rect -4144 3566 -4138 3700
rect -4562 3524 -4548 3564
rect -4608 3308 -4548 3524
rect -4152 3524 -4138 3566
rect -4104 3566 -4098 3700
rect -3686 3700 -3640 3712
rect -4104 3524 -4092 3566
rect -4454 3474 -4246 3480
rect -4454 3440 -4442 3474
rect -4258 3440 -4246 3474
rect -4454 3434 -4246 3440
rect -4380 3308 -4320 3434
rect -4608 3248 -4320 3308
rect -4608 3032 -4548 3248
rect -4380 3122 -4320 3248
rect -4454 3116 -4246 3122
rect -4454 3082 -4442 3116
rect -4258 3082 -4246 3116
rect -4454 3076 -4246 3082
rect -4608 3012 -4596 3032
rect -4602 2886 -4596 3012
rect -4616 2856 -4596 2886
rect -4562 3012 -4548 3032
rect -4152 3032 -4092 3524
rect -3686 3524 -3680 3700
rect -3646 3524 -3640 3700
rect -3686 3512 -3640 3524
rect -3228 3700 -3182 3712
rect -3228 3524 -3222 3700
rect -3188 3524 -3182 3700
rect -3228 3512 -3182 3524
rect -2770 3700 -2724 3712
rect -2770 3524 -2764 3700
rect -2730 3524 -2724 3700
rect -2770 3512 -2724 3524
rect -2312 3700 -2266 3712
rect -2312 3524 -2306 3700
rect -2272 3524 -2266 3700
rect -2312 3512 -2266 3524
rect -1854 3700 -1808 3712
rect -1854 3524 -1848 3700
rect -1814 3524 -1808 3700
rect -1854 3512 -1808 3524
rect -1396 3700 -1350 3712
rect -1396 3524 -1390 3700
rect -1356 3524 -1350 3700
rect -1396 3512 -1350 3524
rect -938 3700 -892 3712
rect -938 3524 -932 3700
rect -898 3524 -892 3700
rect -488 3700 -428 3984
rect -260 3790 -200 4136
rect -332 3784 -124 3790
rect -332 3750 -320 3784
rect -136 3750 -124 3784
rect -332 3744 -124 3750
rect -488 3670 -474 3700
rect -938 3512 -892 3524
rect -480 3524 -474 3670
rect -440 3670 -428 3700
rect -28 3700 32 4136
rect -28 3672 -16 3700
rect -440 3524 -434 3670
rect -22 3580 -16 3672
rect -480 3512 -434 3524
rect -28 3524 -16 3580
rect 18 3672 32 3700
rect 392 3700 452 4136
rect 626 3790 686 4136
rect 546 3784 754 3790
rect 546 3750 558 3784
rect 742 3750 754 3784
rect 546 3744 754 3750
rect 18 3580 24 3672
rect 392 3664 404 3700
rect 18 3524 32 3580
rect 398 3560 404 3664
rect -3996 3474 -3788 3480
rect -3996 3440 -3984 3474
rect -3800 3440 -3788 3474
rect -3996 3434 -3788 3440
rect -3538 3474 -3330 3480
rect -3538 3440 -3526 3474
rect -3342 3440 -3330 3474
rect -3538 3434 -3330 3440
rect -3080 3474 -2872 3480
rect -3080 3440 -3068 3474
rect -2884 3440 -2872 3474
rect -3080 3434 -2872 3440
rect -2622 3474 -2414 3480
rect -2622 3440 -2610 3474
rect -2426 3440 -2414 3474
rect -2622 3434 -2414 3440
rect -2164 3474 -1956 3480
rect -2164 3440 -2152 3474
rect -1968 3440 -1956 3474
rect -2164 3434 -1956 3440
rect -1706 3474 -1498 3480
rect -1706 3440 -1694 3474
rect -1510 3440 -1498 3474
rect -1706 3434 -1498 3440
rect -1248 3474 -1040 3480
rect -1248 3440 -1236 3474
rect -1052 3440 -1040 3474
rect -1248 3434 -1040 3440
rect -790 3474 -582 3480
rect -790 3440 -778 3474
rect -594 3440 -582 3474
rect -790 3434 -582 3440
rect -332 3474 -124 3480
rect -332 3440 -320 3474
rect -136 3440 -124 3474
rect -332 3434 -124 3440
rect -3926 3368 -3866 3434
rect -3464 3368 -3404 3434
rect -3010 3368 -2950 3434
rect -2548 3368 -2488 3434
rect -2094 3368 -2034 3434
rect -1644 3368 -1584 3434
rect -1178 3368 -1118 3434
rect -722 3368 -662 3434
rect -3926 3308 -662 3368
rect -3920 3188 -656 3248
rect -3920 3122 -3860 3188
rect -3458 3122 -3398 3188
rect -3004 3122 -2944 3188
rect -2542 3122 -2482 3188
rect -2088 3122 -2028 3188
rect -1638 3122 -1578 3188
rect -1172 3122 -1112 3188
rect -716 3122 -656 3188
rect -260 3122 -200 3434
rect -3996 3116 -3788 3122
rect -3996 3082 -3984 3116
rect -3800 3082 -3788 3116
rect -3996 3076 -3788 3082
rect -3538 3116 -3330 3122
rect -3538 3082 -3526 3116
rect -3342 3082 -3330 3116
rect -3538 3076 -3330 3082
rect -3080 3116 -2872 3122
rect -3080 3082 -3068 3116
rect -2884 3082 -2872 3116
rect -3080 3076 -2872 3082
rect -2622 3116 -2414 3122
rect -2622 3082 -2610 3116
rect -2426 3082 -2414 3116
rect -2622 3076 -2414 3082
rect -2164 3116 -1956 3122
rect -2164 3082 -2152 3116
rect -1968 3082 -1956 3116
rect -2164 3076 -1956 3082
rect -1706 3116 -1498 3122
rect -1706 3082 -1694 3116
rect -1510 3082 -1498 3116
rect -1706 3076 -1498 3082
rect -1248 3116 -1040 3122
rect -1248 3082 -1236 3116
rect -1052 3082 -1040 3116
rect -1248 3076 -1040 3082
rect -790 3116 -582 3122
rect -790 3082 -778 3116
rect -594 3082 -582 3116
rect -790 3076 -582 3082
rect -332 3116 -124 3122
rect -332 3082 -320 3116
rect -136 3082 -124 3116
rect -332 3076 -124 3082
rect -4562 2856 -4556 3012
rect -4152 3004 -4138 3032
rect -4616 2476 -4556 2856
rect -4144 2856 -4138 3004
rect -4104 3004 -4092 3032
rect -3686 3032 -3640 3044
rect -4104 2856 -4098 3004
rect -4144 2844 -4098 2856
rect -3686 2856 -3680 3032
rect -3646 2856 -3640 3032
rect -3686 2844 -3640 2856
rect -3228 3032 -3182 3044
rect -3228 2856 -3222 3032
rect -3188 2856 -3182 3032
rect -3228 2844 -3182 2856
rect -2770 3032 -2724 3044
rect -2770 2856 -2764 3032
rect -2730 2856 -2724 3032
rect -2770 2844 -2724 2856
rect -2312 3032 -2266 3044
rect -2312 2856 -2306 3032
rect -2272 2856 -2266 3032
rect -2312 2844 -2266 2856
rect -1854 3032 -1808 3044
rect -1854 2856 -1848 3032
rect -1814 2856 -1808 3032
rect -1854 2844 -1808 2856
rect -1396 3032 -1350 3044
rect -1396 2856 -1390 3032
rect -1356 2856 -1350 3032
rect -1396 2844 -1350 2856
rect -938 3032 -892 3044
rect -938 2856 -932 3032
rect -898 2856 -892 3032
rect -480 3032 -434 3044
rect -480 2884 -474 3032
rect -938 2844 -892 2856
rect -488 2856 -474 2884
rect -440 2884 -434 3032
rect -28 3032 32 3524
rect -440 2856 -428 2884
rect -4454 2806 -4246 2812
rect -4454 2772 -4442 2806
rect -4258 2772 -4246 2806
rect -4454 2766 -4246 2772
rect -3996 2806 -3788 2812
rect -3996 2772 -3984 2806
rect -3800 2772 -3788 2806
rect -3996 2766 -3788 2772
rect -3538 2806 -3330 2812
rect -3538 2772 -3526 2806
rect -3342 2772 -3330 2806
rect -3538 2766 -3330 2772
rect -3080 2806 -2872 2812
rect -3080 2772 -3068 2806
rect -2884 2772 -2872 2806
rect -3080 2766 -2872 2772
rect -2622 2806 -2414 2812
rect -2622 2772 -2610 2806
rect -2426 2772 -2414 2806
rect -2622 2766 -2414 2772
rect -2164 2806 -1956 2812
rect -2164 2772 -2152 2806
rect -1968 2772 -1956 2806
rect -2164 2766 -1956 2772
rect -1706 2806 -1498 2812
rect -1706 2772 -1694 2806
rect -1510 2772 -1498 2806
rect -1706 2766 -1498 2772
rect -1248 2806 -1040 2812
rect -1248 2772 -1236 2806
rect -1052 2772 -1040 2806
rect -1248 2766 -1040 2772
rect -790 2806 -582 2812
rect -790 2772 -778 2806
rect -594 2772 -582 2806
rect -790 2766 -582 2772
rect -4376 2476 -4316 2766
rect -3926 2700 -3866 2766
rect -3464 2700 -3404 2766
rect -3010 2700 -2950 2766
rect -2548 2700 -2488 2766
rect -2094 2700 -2034 2766
rect -1644 2700 -1584 2766
rect -1178 2700 -1118 2766
rect -722 2700 -662 2766
rect -3926 2640 -662 2700
rect -488 2476 -428 2856
rect -28 2856 -16 3032
rect 18 2856 32 3032
rect -332 2806 -124 2812
rect -332 2772 -320 2806
rect -136 2772 -124 2806
rect -332 2766 -124 2772
rect -262 2476 -202 2766
rect -28 2476 32 2856
rect 388 3524 404 3560
rect 438 3664 452 3700
rect 848 3700 908 4136
rect 4506 3996 4512 4056
rect 4572 3996 4578 4056
rect 3352 3916 3358 3920
rect 1070 3856 1076 3916
rect 1136 3914 3358 3916
rect 1136 3856 1538 3914
rect 1076 3790 1140 3856
rect 1532 3854 1538 3856
rect 1598 3856 1992 3914
rect 1598 3854 1604 3856
rect 1986 3854 1992 3856
rect 2052 3856 2454 3914
rect 2052 3854 2058 3856
rect 2448 3854 2454 3856
rect 2514 3856 2908 3914
rect 2514 3854 2520 3856
rect 2902 3854 2908 3856
rect 2968 3860 3358 3914
rect 3418 3916 3424 3920
rect 3418 3860 3824 3916
rect 2968 3856 3824 3860
rect 3884 3856 4280 3916
rect 4340 3856 4346 3916
rect 2968 3854 2974 3856
rect 1538 3790 1602 3854
rect 1992 3790 2056 3854
rect 2454 3790 2518 3854
rect 2908 3790 2972 3854
rect 3358 3790 3422 3856
rect 3824 3790 3888 3856
rect 4280 3790 4344 3856
rect 1004 3784 1212 3790
rect 1004 3750 1016 3784
rect 1200 3750 1212 3784
rect 1004 3744 1212 3750
rect 1462 3784 1670 3790
rect 1462 3750 1474 3784
rect 1658 3750 1670 3784
rect 1462 3744 1670 3750
rect 1920 3784 2128 3790
rect 1920 3750 1932 3784
rect 2116 3750 2128 3784
rect 1920 3744 2128 3750
rect 2378 3784 2586 3790
rect 2378 3750 2390 3784
rect 2574 3750 2586 3784
rect 2378 3744 2586 3750
rect 2836 3784 3044 3790
rect 2836 3750 2848 3784
rect 3032 3750 3044 3784
rect 2836 3744 3044 3750
rect 3294 3784 3502 3790
rect 3294 3750 3306 3784
rect 3490 3750 3502 3784
rect 3294 3744 3502 3750
rect 3752 3784 3960 3790
rect 3752 3750 3764 3784
rect 3948 3750 3960 3784
rect 3752 3744 3960 3750
rect 4210 3784 4418 3790
rect 4210 3750 4222 3784
rect 4406 3750 4418 3784
rect 4210 3744 4418 3750
rect 438 3560 444 3664
rect 848 3636 862 3700
rect 856 3568 862 3636
rect 438 3524 448 3560
rect 388 3370 448 3524
rect 848 3524 862 3568
rect 896 3636 908 3700
rect 1314 3700 1360 3712
rect 896 3568 902 3636
rect 896 3524 908 3568
rect 546 3474 754 3480
rect 546 3440 558 3474
rect 742 3440 754 3474
rect 546 3434 754 3440
rect 616 3370 676 3434
rect 848 3370 908 3524
rect 1314 3524 1320 3700
rect 1354 3524 1360 3700
rect 1314 3512 1360 3524
rect 1772 3700 1818 3712
rect 1772 3524 1778 3700
rect 1812 3524 1818 3700
rect 1772 3512 1818 3524
rect 2230 3700 2276 3712
rect 2230 3524 2236 3700
rect 2270 3524 2276 3700
rect 2230 3512 2276 3524
rect 2688 3700 2734 3712
rect 2688 3524 2694 3700
rect 2728 3524 2734 3700
rect 2688 3512 2734 3524
rect 3146 3700 3192 3712
rect 3146 3524 3152 3700
rect 3186 3524 3192 3700
rect 3146 3512 3192 3524
rect 3604 3700 3650 3712
rect 3604 3524 3610 3700
rect 3644 3524 3650 3700
rect 3604 3512 3650 3524
rect 4062 3700 4108 3712
rect 4062 3524 4068 3700
rect 4102 3524 4108 3700
rect 4512 3700 4572 3996
rect 4752 3790 4812 4136
rect 4668 3784 4876 3790
rect 4668 3750 4680 3784
rect 4864 3750 4876 3784
rect 4668 3744 4876 3750
rect 4512 3658 4526 3700
rect 4062 3512 4108 3524
rect 4520 3524 4526 3658
rect 4560 3658 4572 3700
rect 4970 3700 5030 4136
rect 4970 3660 4984 3700
rect 4560 3524 4566 3658
rect 4978 3570 4984 3660
rect 4520 3512 4566 3524
rect 4968 3524 4984 3570
rect 5018 3660 5030 3700
rect 5316 4012 5428 4136
rect 5018 3570 5024 3660
rect 5018 3524 5028 3570
rect 1004 3474 1212 3480
rect 1004 3440 1016 3474
rect 1200 3440 1212 3474
rect 1004 3434 1212 3440
rect 1462 3474 1670 3480
rect 1462 3440 1474 3474
rect 1658 3440 1670 3474
rect 1462 3434 1670 3440
rect 1920 3474 2128 3480
rect 1920 3440 1932 3474
rect 2116 3440 2128 3474
rect 1920 3434 2128 3440
rect 2378 3474 2586 3480
rect 2378 3440 2390 3474
rect 2574 3440 2586 3474
rect 2378 3434 2586 3440
rect 2836 3474 3044 3480
rect 2836 3440 2848 3474
rect 3032 3440 3044 3474
rect 2836 3434 3044 3440
rect 3294 3474 3502 3480
rect 3294 3440 3306 3474
rect 3490 3440 3502 3474
rect 3294 3434 3502 3440
rect 3752 3474 3960 3480
rect 3752 3440 3764 3474
rect 3948 3440 3960 3474
rect 3752 3434 3960 3440
rect 4210 3474 4418 3480
rect 4210 3440 4222 3474
rect 4406 3440 4418 3474
rect 4210 3434 4418 3440
rect 4668 3474 4876 3480
rect 4668 3440 4680 3474
rect 4864 3440 4876 3474
rect 4668 3434 4876 3440
rect 388 3310 908 3370
rect 388 2476 448 3310
rect 616 2476 676 3310
rect 848 2476 908 3310
rect 1074 3368 1134 3434
rect 1536 3368 1596 3434
rect 1990 3368 2050 3434
rect 2452 3368 2512 3434
rect 2906 3368 2966 3434
rect 3356 3368 3416 3434
rect 3822 3368 3882 3434
rect 4278 3368 4338 3434
rect 1074 3308 4338 3368
rect 4742 2476 4802 3434
rect 4968 2476 5028 3524
rect -4680 2448 5090 2476
rect -4680 2362 -4630 2448
rect -4534 2362 -4050 2448
rect -3954 2362 -3450 2448
rect -3354 2362 -2850 2448
rect -2754 2362 -2250 2448
rect -2154 2362 -1650 2448
rect -1554 2362 -1050 2448
rect -954 2362 -450 2448
rect -354 2362 150 2448
rect 246 2362 750 2448
rect 846 2362 1350 2448
rect 1446 2362 1950 2448
rect 2046 2362 2550 2448
rect 2646 2362 3150 2448
rect 3246 2362 3750 2448
rect 3846 2362 4350 2448
rect 4446 2362 4950 2448
rect 5046 2362 5090 2448
rect -4680 2332 5090 2362
rect -5028 1884 -4916 2008
rect -4316 1884 -4306 2184
rect 4706 1884 4716 2184
rect 5316 2008 5322 4012
rect 5422 2008 5428 4012
rect 5316 1884 5428 2008
rect -5028 1878 5428 1884
rect -5028 1778 -4922 1878
rect 5322 1778 5428 1878
rect -5028 1772 5428 1778
<< via1 >>
rect -4916 9916 -4316 10216
rect 4716 9916 5316 10216
rect -4064 9656 -3968 9742
rect -3464 9656 -3368 9742
rect -2864 9656 -2768 9742
rect -2264 9656 -2168 9742
rect -1664 9656 -1568 9742
rect -1064 9656 -968 9742
rect -464 9656 -368 9742
rect 136 9656 232 9742
rect 736 9656 832 9742
rect 1336 9656 1432 9742
rect 1936 9656 2032 9742
rect 2536 9656 2632 9742
rect 3136 9656 3232 9742
rect 3736 9656 3832 9742
rect 4156 9656 4252 9742
rect -3360 9024 -3300 9084
rect -2904 9024 -2844 9084
rect -2444 9024 -2384 9084
rect -1988 9024 -1928 9084
rect -3364 7050 -3304 7110
rect -1530 9024 -1470 9084
rect -1066 9024 -1006 9084
rect -2908 7050 -2848 7110
rect -2448 7050 -2388 7110
rect -616 9024 -556 9084
rect -160 9024 -100 9084
rect 308 9024 368 9084
rect 766 9024 826 9084
rect -1992 7050 -1932 7110
rect -1534 7050 -1474 7110
rect -1070 7050 -1010 7110
rect -616 7050 -556 7110
rect 1222 9024 1282 9084
rect 1678 9024 1738 9084
rect -158 7106 -98 7110
rect -158 7058 -152 7106
rect -152 7058 -104 7106
rect -104 7058 -98 7106
rect -158 7050 -98 7058
rect 76 7062 136 7122
rect 302 7052 362 7110
rect 302 7050 362 7052
rect 2134 9024 2194 9084
rect 2590 9024 2650 9084
rect 758 7050 818 7110
rect 1218 7050 1278 7110
rect 3048 9024 3108 9084
rect 3508 9024 3568 9084
rect 1674 7050 1734 7110
rect 2130 7050 2190 7110
rect 2586 7050 2646 7110
rect 3044 7050 3104 7110
rect 3504 7050 3564 7110
rect -4150 6464 -4090 6524
rect -3926 4786 -3866 4846
rect -3464 4786 -3404 4846
rect -3010 4790 -2950 4850
rect -2548 4790 -2488 4850
rect -2094 4784 -2034 4844
rect -1644 4790 -1584 4850
rect -1178 4790 -1118 4850
rect -722 4786 -662 4846
rect -488 4664 -428 4724
rect 1076 4786 1136 4846
rect 1538 4794 1598 4854
rect 1992 4788 2052 4848
rect 2454 4788 2514 4848
rect 2908 4788 2968 4848
rect 3358 4794 3418 4854
rect 3824 4788 3884 4848
rect 4280 4788 4340 4848
rect 4512 4658 4572 4718
rect -488 3984 -428 4044
rect -3926 3850 -3866 3910
rect -3464 3856 -3404 3916
rect -3010 3850 -2950 3910
rect -2548 3856 -2488 3916
rect -2094 3856 -2034 3916
rect -1644 3856 -1584 3916
rect -1178 3850 -1118 3910
rect -722 3856 -662 3916
rect 4512 3996 4572 4056
rect 1076 3856 1136 3916
rect 1538 3854 1598 3914
rect 1992 3854 2052 3914
rect 2454 3854 2514 3914
rect 2908 3854 2968 3914
rect 3358 3860 3418 3920
rect 3824 3856 3884 3916
rect 4280 3856 4340 3916
rect -4630 2362 -4534 2448
rect -4050 2362 -3954 2448
rect -3450 2362 -3354 2448
rect -2850 2362 -2754 2448
rect -2250 2362 -2154 2448
rect -1650 2362 -1554 2448
rect -1050 2362 -954 2448
rect -450 2362 -354 2448
rect 150 2362 246 2448
rect 750 2362 846 2448
rect 1350 2362 1446 2448
rect 1950 2362 2046 2448
rect 2550 2362 2646 2448
rect 3150 2362 3246 2448
rect 3750 2362 3846 2448
rect 4350 2362 4446 2448
rect 4950 2362 5046 2448
rect -4916 1884 -4316 2184
rect 4716 1884 5316 2184
<< metal2 >>
rect -4916 10216 -4316 10226
rect -4916 9906 -4316 9916
rect 4716 10216 5316 10226
rect 4716 9906 5316 9916
rect -4078 9742 4278 9756
rect -4078 9656 -4064 9742
rect -3968 9656 -3464 9742
rect -3368 9656 -2864 9742
rect -2768 9656 -2264 9742
rect -2168 9656 -1664 9742
rect -1568 9656 -1064 9742
rect -968 9656 -464 9742
rect -368 9656 136 9742
rect 232 9656 736 9742
rect 832 9656 1336 9742
rect 1432 9656 1936 9742
rect 2032 9656 2536 9742
rect 2632 9656 3136 9742
rect 3232 9656 3736 9742
rect 3832 9656 4156 9742
rect 4252 9656 4278 9742
rect -4078 9646 4278 9656
rect -3360 9084 -3300 9090
rect -2904 9084 -2844 9090
rect -2444 9084 -2384 9090
rect -1988 9084 -1928 9090
rect -1530 9084 -1470 9090
rect -1066 9084 -1006 9090
rect -616 9084 -556 9090
rect -160 9084 -100 9090
rect 308 9084 368 9090
rect 766 9084 826 9090
rect 1222 9084 1282 9090
rect 1678 9084 1738 9090
rect 2134 9084 2194 9090
rect 2590 9084 2650 9090
rect 3048 9084 3108 9090
rect 3508 9084 3568 9090
rect -3300 9024 -2904 9084
rect -2844 9024 -2444 9084
rect -2384 9024 -1988 9084
rect -1928 9024 -1530 9084
rect -1470 9024 -1066 9084
rect -1006 9024 -616 9084
rect -556 9024 -160 9084
rect -100 9024 308 9084
rect 368 9024 766 9084
rect 826 9024 1222 9084
rect 1282 9024 1678 9084
rect 1738 9024 2134 9084
rect 2194 9024 2590 9084
rect 2650 9024 3048 9084
rect 3108 9024 3508 9084
rect -3360 9018 -3300 9024
rect -2904 9018 -2844 9024
rect -2444 9018 -2384 9024
rect -1988 9018 -1928 9024
rect -1530 9018 -1470 9024
rect -1066 9018 -1006 9024
rect -616 9018 -556 9024
rect -160 9018 -100 9024
rect 308 9018 368 9024
rect 766 9018 826 9024
rect 1222 9018 1282 9024
rect 1678 9018 1738 9024
rect 2134 9018 2194 9024
rect 2590 9018 2650 9024
rect 3048 9018 3108 9024
rect 3508 9018 3568 9024
rect -3364 7110 -3304 7116
rect -2908 7110 -2848 7116
rect -2448 7110 -2388 7116
rect -1992 7110 -1932 7116
rect -1534 7110 -1474 7116
rect -1070 7110 -1010 7116
rect -616 7110 -556 7116
rect -158 7110 -98 7116
rect -3304 7050 -2908 7110
rect -2848 7050 -2448 7110
rect -2388 7050 -1992 7110
rect -1932 7050 -1534 7110
rect -1474 7050 -1070 7110
rect -1010 7050 -616 7110
rect -556 7050 -158 7110
rect 70 7062 76 7122
rect 136 7062 142 7122
rect 302 7110 362 7116
rect 758 7110 818 7116
rect 1218 7110 1278 7116
rect 1674 7110 1734 7116
rect 2130 7110 2190 7116
rect 2586 7110 2646 7116
rect 3044 7110 3104 7116
rect 3504 7110 3564 7116
rect -3364 7044 -3304 7050
rect -2908 7044 -2848 7050
rect -2448 7044 -2388 7050
rect -1992 7044 -1932 7050
rect -1534 7044 -1474 7050
rect -1070 7044 -1010 7050
rect -616 7044 -556 7050
rect -158 7044 -98 7050
rect -4150 6524 -4090 6530
rect 76 6524 136 7062
rect 362 7050 758 7110
rect 818 7050 1218 7110
rect 1278 7050 1674 7110
rect 1734 7050 2130 7110
rect 2190 7050 2586 7110
rect 2646 7050 3044 7110
rect 3104 7050 3504 7110
rect 302 7044 362 7050
rect 758 7044 818 7050
rect 1218 7044 1278 7050
rect 1674 7044 1734 7050
rect 2130 7044 2190 7050
rect 2586 7044 2646 7050
rect 3044 7044 3104 7050
rect 3504 7044 3564 7050
rect -4090 6464 136 6524
rect -4150 6458 -4090 6464
rect -3932 4786 -3926 4846
rect -3866 4786 -3860 4846
rect -3470 4786 -3464 4846
rect -3404 4786 -3398 4846
rect -3016 4790 -3010 4850
rect -2950 4790 -2944 4850
rect -2554 4790 -2548 4850
rect -2488 4790 -2482 4850
rect -3926 4392 -3866 4786
rect -3464 4392 -3404 4786
rect -3010 4392 -2950 4790
rect -2548 4392 -2488 4790
rect -2100 4784 -2094 4844
rect -2034 4784 -2028 4844
rect -1650 4790 -1644 4850
rect -1584 4790 -1578 4850
rect -1184 4790 -1178 4850
rect -1118 4790 -1112 4850
rect -2094 4392 -2034 4784
rect -1644 4392 -1584 4790
rect -1178 4392 -1118 4790
rect -728 4786 -722 4846
rect -662 4786 -656 4846
rect 1070 4786 1076 4846
rect 1136 4786 1142 4846
rect 1532 4794 1538 4854
rect 1598 4794 1604 4854
rect -722 4392 -662 4786
rect -3928 4332 -662 4392
rect -3926 3910 -3866 4332
rect -3464 3916 -3404 4332
rect -3464 3850 -3404 3856
rect -3010 3910 -2950 4332
rect -2548 3916 -2488 4332
rect -2548 3850 -2488 3856
rect -2094 3916 -2034 4332
rect -2094 3850 -2034 3856
rect -1644 3916 -1584 4332
rect -1644 3850 -1584 3856
rect -1178 3910 -1118 4332
rect -722 3916 -662 4332
rect -488 4724 -428 4730
rect -488 4386 -428 4664
rect 1076 4386 1136 4786
rect 1538 4386 1598 4794
rect 1986 4788 1992 4848
rect 2052 4788 2058 4848
rect 2448 4788 2454 4848
rect 2514 4788 2520 4848
rect 2902 4788 2908 4848
rect 2968 4788 2974 4848
rect 3352 4794 3358 4854
rect 3418 4794 3424 4854
rect 1992 4386 2052 4788
rect 2454 4386 2514 4788
rect 2908 4386 2968 4788
rect 3358 4386 3418 4794
rect 3818 4788 3824 4848
rect 3884 4788 3890 4848
rect 4274 4788 4280 4848
rect 4340 4788 4346 4848
rect 3824 4386 3884 4788
rect 4280 4386 4340 4788
rect 4506 4658 4512 4718
rect 4572 4658 4578 4718
rect -488 4326 4340 4386
rect -488 4044 -428 4326
rect -494 3984 -488 4044
rect -428 3984 -422 4044
rect -722 3850 -662 3856
rect 1076 3916 1136 4326
rect 1076 3850 1136 3856
rect 1538 3914 1598 4326
rect -3926 3844 -3866 3850
rect -3010 3844 -2950 3850
rect -1178 3844 -1118 3850
rect 1538 3848 1598 3854
rect 1992 3914 2052 4326
rect 1992 3848 2052 3854
rect 2454 3914 2514 4326
rect 2454 3848 2514 3854
rect 2908 3914 2968 4326
rect 3358 3920 3418 4326
rect 3358 3854 3418 3860
rect 3824 3916 3884 4326
rect 2908 3848 2968 3854
rect 3824 3850 3884 3856
rect 4280 3916 4340 4326
rect 4512 4382 4572 4658
rect 4512 4322 5598 4382
rect 4512 4056 4572 4322
rect 5498 4193 5598 4322
rect 5494 4103 5503 4193
rect 5593 4103 5602 4193
rect 5498 4098 5598 4103
rect 4512 3990 4572 3996
rect 4280 3850 4340 3856
rect -4680 2448 5090 2476
rect -4680 2362 -4630 2448
rect -4534 2362 -4050 2448
rect -3954 2362 -3450 2448
rect -3354 2362 -2850 2448
rect -2754 2362 -2250 2448
rect -2154 2362 -1650 2448
rect -1554 2362 -1050 2448
rect -954 2362 -450 2448
rect -354 2362 150 2448
rect 246 2362 750 2448
rect 846 2362 1350 2448
rect 1446 2362 1950 2448
rect 2046 2362 2550 2448
rect 2646 2362 3150 2448
rect 3246 2362 3750 2448
rect 3846 2362 4350 2448
rect 4446 2362 4950 2448
rect 5046 2362 5090 2448
rect -4680 2332 5090 2362
rect -4916 2184 -4316 2194
rect -4916 1874 -4316 1884
rect 4716 2184 5316 2194
rect 4716 1874 5316 1884
<< via2 >>
rect -4916 9916 -4316 10216
rect 4716 9916 5316 10216
rect -4064 9656 -3968 9742
rect -3464 9656 -3368 9742
rect -2864 9656 -2768 9742
rect -2264 9656 -2168 9742
rect -1664 9656 -1568 9742
rect -1064 9656 -968 9742
rect -464 9656 -368 9742
rect 136 9656 232 9742
rect 736 9656 832 9742
rect 1336 9656 1432 9742
rect 1936 9656 2032 9742
rect 2536 9656 2632 9742
rect 3136 9656 3232 9742
rect 3736 9656 3832 9742
rect 4156 9656 4252 9742
rect 5503 4103 5593 4193
rect -4630 2362 -4534 2448
rect -4050 2362 -3954 2448
rect -3450 2362 -3354 2448
rect -2850 2362 -2754 2448
rect -2250 2362 -2154 2448
rect -1650 2362 -1554 2448
rect -1050 2362 -954 2448
rect -450 2362 -354 2448
rect 150 2362 246 2448
rect 750 2362 846 2448
rect 1350 2362 1446 2448
rect 1950 2362 2046 2448
rect 2550 2362 2646 2448
rect 3150 2362 3246 2448
rect 3750 2362 3846 2448
rect 4350 2362 4446 2448
rect 4950 2362 5046 2448
rect -4916 1884 -4316 2184
rect 4716 1884 5316 2184
<< metal3 >>
rect -4926 10216 -4306 10221
rect -4926 9916 -4916 10216
rect -4316 9916 -4306 10216
rect -4926 9911 -4306 9916
rect 4706 10216 5326 10221
rect 4706 9916 4716 10216
rect 5316 9916 5326 10216
rect 4706 9911 5326 9916
rect -4078 9742 4278 9756
rect -4078 9656 -4064 9742
rect -3968 9656 -3464 9742
rect -3368 9656 -2864 9742
rect -2768 9656 -2264 9742
rect -2168 9656 -1664 9742
rect -1568 9656 -1064 9742
rect -968 9656 -464 9742
rect -368 9656 136 9742
rect 232 9656 736 9742
rect 832 9656 1336 9742
rect 1432 9656 1936 9742
rect 2032 9656 2536 9742
rect 2632 9656 3136 9742
rect 3232 9656 3736 9742
rect 3832 9656 4156 9742
rect 4252 9656 4278 9742
rect -4078 9646 4278 9656
rect 5698 5384 9326 5518
rect 5698 5012 6335 5384
rect 6399 5382 9326 5384
rect 6399 5012 7054 5382
rect 7118 5012 7773 5382
rect 7837 5012 8492 5382
rect 8556 5012 9211 5382
rect 9275 5012 9326 5382
rect 5698 4682 9326 5012
rect 5698 4314 6335 4682
rect 6399 4314 7054 4682
rect 7118 4314 7773 4682
rect 7837 4314 8492 4682
rect 8556 4314 9211 4682
rect 9275 4314 9326 4682
rect 5498 4197 5598 4198
rect 5493 4099 5499 4197
rect 5597 4099 5603 4197
rect 5498 4098 5598 4099
rect 5698 3982 9326 4314
rect 5698 3614 6335 3982
rect 6399 3614 7054 3982
rect 7118 3614 7773 3982
rect 7837 3614 8492 3982
rect 8556 3614 9211 3982
rect 9275 3614 9326 3982
rect 5698 3282 9326 3614
rect 5698 2914 6335 3282
rect 6399 2914 7054 3282
rect 7118 2914 7773 3282
rect 7837 2914 8492 3282
rect 8556 2914 9211 3282
rect 9275 2914 9326 3282
rect 5698 2582 9326 2914
rect -4680 2448 5090 2476
rect -4680 2362 -4630 2448
rect -4534 2362 -4050 2448
rect -3954 2362 -3450 2448
rect -3354 2362 -2850 2448
rect -2754 2362 -2250 2448
rect -2154 2362 -1650 2448
rect -1554 2362 -1050 2448
rect -954 2362 -450 2448
rect -354 2362 150 2448
rect 246 2362 750 2448
rect 846 2362 1350 2448
rect 1446 2362 1950 2448
rect 2046 2362 2550 2448
rect 2646 2362 3150 2448
rect 3246 2362 3750 2448
rect 3846 2362 4350 2448
rect 4446 2362 4950 2448
rect 5046 2362 5090 2448
rect -4680 2332 5090 2362
rect 5698 2214 6335 2582
rect 6399 2214 7054 2582
rect 7118 2214 7773 2582
rect 7837 2214 8492 2582
rect 8556 2214 9211 2582
rect 9275 2214 9326 2582
rect -4926 2184 -4306 2189
rect -4926 1884 -4916 2184
rect -4316 1884 -4306 2184
rect -4926 1879 -4306 1884
rect 4706 2184 5326 2189
rect 4706 1884 4716 2184
rect 5316 1884 5326 2184
rect 5698 2064 9326 2214
rect 4706 1879 5326 1884
<< via3 >>
rect -4916 9916 -4316 10216
rect 4716 9916 5316 10216
rect -4064 9656 -3968 9742
rect -3464 9656 -3368 9742
rect -2864 9656 -2768 9742
rect -2264 9656 -2168 9742
rect -1664 9656 -1568 9742
rect -1064 9656 -968 9742
rect -464 9656 -368 9742
rect 136 9656 232 9742
rect 736 9656 832 9742
rect 1336 9656 1432 9742
rect 1936 9656 2032 9742
rect 2536 9656 2632 9742
rect 3136 9656 3232 9742
rect 3736 9656 3832 9742
rect 4156 9656 4252 9742
rect 6335 5012 6399 5384
rect 7054 5012 7118 5382
rect 7773 5012 7837 5382
rect 8492 5012 8556 5382
rect 9211 5012 9275 5382
rect 6335 4314 6399 4682
rect 7054 4314 7118 4682
rect 7773 4314 7837 4682
rect 8492 4314 8556 4682
rect 9211 4314 9275 4682
rect 5499 4193 5597 4197
rect 5499 4103 5503 4193
rect 5503 4103 5593 4193
rect 5593 4103 5597 4193
rect 5499 4099 5597 4103
rect 6335 3614 6399 3982
rect 7054 3614 7118 3982
rect 7773 3614 7837 3982
rect 8492 3614 8556 3982
rect 9211 3614 9275 3982
rect 6335 2914 6399 3282
rect 7054 2914 7118 3282
rect 7773 2914 7837 3282
rect 8492 2914 8556 3282
rect 9211 2914 9275 3282
rect -4630 2362 -4534 2448
rect -4050 2362 -3954 2448
rect -3450 2362 -3354 2448
rect -2850 2362 -2754 2448
rect -2250 2362 -2154 2448
rect -1650 2362 -1554 2448
rect -1050 2362 -954 2448
rect -450 2362 -354 2448
rect 150 2362 246 2448
rect 750 2362 846 2448
rect 1350 2362 1446 2448
rect 1950 2362 2046 2448
rect 2550 2362 2646 2448
rect 3150 2362 3246 2448
rect 3750 2362 3846 2448
rect 4350 2362 4446 2448
rect 4950 2362 5046 2448
rect 6335 2214 6399 2582
rect 7054 2214 7118 2582
rect 7773 2214 7837 2582
rect 8492 2214 8556 2582
rect 9211 2214 9275 2582
rect -4916 1884 -4316 2184
rect 4716 1884 5316 2184
<< mimcap >>
rect 5820 5360 6220 5400
rect 5820 5040 5860 5360
rect 6180 5040 6220 5360
rect 5820 5000 6220 5040
rect 6539 5360 6939 5400
rect 6539 5040 6579 5360
rect 6899 5040 6939 5360
rect 6539 5000 6939 5040
rect 7258 5360 7658 5400
rect 7258 5040 7298 5360
rect 7618 5040 7658 5360
rect 7258 5000 7658 5040
rect 7977 5360 8377 5400
rect 7977 5040 8017 5360
rect 8337 5040 8377 5360
rect 7977 5000 8377 5040
rect 8696 5360 9096 5400
rect 8696 5040 8736 5360
rect 9056 5040 9096 5360
rect 8696 5000 9096 5040
rect 5820 4660 6220 4700
rect 5820 4340 5860 4660
rect 6180 4340 6220 4660
rect 5820 4300 6220 4340
rect 6539 4660 6939 4700
rect 6539 4340 6579 4660
rect 6899 4340 6939 4660
rect 6539 4300 6939 4340
rect 7258 4660 7658 4700
rect 7258 4340 7298 4660
rect 7618 4340 7658 4660
rect 7258 4300 7658 4340
rect 7977 4660 8377 4700
rect 7977 4340 8017 4660
rect 8337 4340 8377 4660
rect 7977 4300 8377 4340
rect 8696 4660 9096 4700
rect 8696 4340 8736 4660
rect 9056 4340 9096 4660
rect 8696 4300 9096 4340
rect 5820 3960 6220 4000
rect 5820 3640 5860 3960
rect 6180 3640 6220 3960
rect 5820 3600 6220 3640
rect 6539 3960 6939 4000
rect 6539 3640 6579 3960
rect 6899 3640 6939 3960
rect 6539 3600 6939 3640
rect 7258 3960 7658 4000
rect 7258 3640 7298 3960
rect 7618 3640 7658 3960
rect 7258 3600 7658 3640
rect 7977 3960 8377 4000
rect 7977 3640 8017 3960
rect 8337 3640 8377 3960
rect 7977 3600 8377 3640
rect 8696 3960 9096 4000
rect 8696 3640 8736 3960
rect 9056 3640 9096 3960
rect 8696 3600 9096 3640
rect 5820 3260 6220 3300
rect 5820 2940 5860 3260
rect 6180 2940 6220 3260
rect 5820 2900 6220 2940
rect 6539 3260 6939 3300
rect 6539 2940 6579 3260
rect 6899 2940 6939 3260
rect 6539 2900 6939 2940
rect 7258 3260 7658 3300
rect 7258 2940 7298 3260
rect 7618 2940 7658 3260
rect 7258 2900 7658 2940
rect 7977 3260 8377 3300
rect 7977 2940 8017 3260
rect 8337 2940 8377 3260
rect 7977 2900 8377 2940
rect 8696 3260 9096 3300
rect 8696 2940 8736 3260
rect 9056 2940 9096 3260
rect 8696 2900 9096 2940
rect 5820 2560 6220 2600
rect 5820 2240 5860 2560
rect 6180 2240 6220 2560
rect 5820 2200 6220 2240
rect 6539 2560 6939 2600
rect 6539 2240 6579 2560
rect 6899 2240 6939 2560
rect 6539 2200 6939 2240
rect 7258 2560 7658 2600
rect 7258 2240 7298 2560
rect 7618 2240 7658 2560
rect 7258 2200 7658 2240
rect 7977 2560 8377 2600
rect 7977 2240 8017 2560
rect 8337 2240 8377 2560
rect 7977 2200 8377 2240
rect 8696 2560 9096 2600
rect 8696 2240 8736 2560
rect 9056 2240 9096 2560
rect 8696 2200 9096 2240
<< mimcapcontact >>
rect 5860 5040 6180 5360
rect 6579 5040 6899 5360
rect 7298 5040 7618 5360
rect 8017 5040 8337 5360
rect 8736 5040 9056 5360
rect 5860 4340 6180 4660
rect 6579 4340 6899 4660
rect 7298 4340 7618 4660
rect 8017 4340 8337 4660
rect 8736 4340 9056 4660
rect 5860 3640 6180 3960
rect 6579 3640 6899 3960
rect 7298 3640 7618 3960
rect 8017 3640 8337 3960
rect 8736 3640 9056 3960
rect 5860 2940 6180 3260
rect 6579 2940 6899 3260
rect 7298 2940 7618 3260
rect 8017 2940 8337 3260
rect 8736 2940 9056 3260
rect 5860 2240 6180 2560
rect 6579 2240 6899 2560
rect 7298 2240 7618 2560
rect 8017 2240 8337 2560
rect 8736 2240 9056 2560
<< metal4 >>
rect -5100 10216 9448 10400
rect -5100 9916 -4916 10216
rect -4316 9916 4716 10216
rect 5316 9916 9448 10216
rect -5100 9742 9448 9916
rect -5100 9656 -4064 9742
rect -3968 9656 -3464 9742
rect -3368 9656 -2864 9742
rect -2768 9656 -2264 9742
rect -2168 9656 -1664 9742
rect -1568 9656 -1064 9742
rect -968 9656 -464 9742
rect -368 9656 136 9742
rect 232 9656 736 9742
rect 832 9656 1336 9742
rect 1432 9656 1936 9742
rect 2032 9656 2536 9742
rect 2632 9656 3136 9742
rect 3232 9656 3736 9742
rect 3832 9656 4156 9742
rect 4252 9656 9448 9742
rect -5100 9600 9448 9656
rect 6319 5384 6415 5400
rect 5859 5360 6181 5361
rect 5859 5040 5860 5360
rect 6180 5244 6181 5360
rect 6319 5244 6335 5384
rect 6180 5144 6335 5244
rect 6180 5040 6181 5144
rect 5859 5039 6181 5040
rect 5974 4661 6074 5039
rect 6310 5012 6335 5144
rect 6399 5244 6415 5384
rect 7038 5382 7134 5398
rect 6578 5360 6900 5361
rect 6578 5244 6579 5360
rect 6399 5144 6579 5244
rect 6399 5012 6415 5144
rect 6578 5040 6579 5144
rect 6899 5244 6900 5360
rect 7038 5244 7054 5382
rect 6899 5144 7054 5244
rect 6899 5040 6900 5144
rect 6578 5039 6900 5040
rect 6310 4996 6415 5012
rect 7038 5012 7054 5144
rect 7118 5244 7134 5382
rect 7757 5382 7853 5398
rect 7297 5360 7619 5361
rect 7297 5244 7298 5360
rect 7118 5144 7298 5244
rect 7118 5012 7134 5144
rect 7297 5040 7298 5144
rect 7618 5244 7619 5360
rect 7757 5244 7773 5382
rect 7618 5144 7773 5244
rect 7618 5040 7619 5144
rect 7297 5039 7619 5040
rect 7038 4996 7134 5012
rect 7757 5012 7773 5144
rect 7837 5244 7853 5382
rect 8476 5382 8572 5398
rect 8016 5360 8338 5361
rect 8016 5244 8017 5360
rect 7837 5144 8017 5244
rect 7837 5012 7853 5144
rect 8016 5040 8017 5144
rect 8337 5244 8338 5360
rect 8476 5244 8492 5382
rect 8337 5144 8492 5244
rect 8337 5040 8338 5144
rect 8016 5039 8338 5040
rect 7757 4996 7853 5012
rect 8476 5012 8492 5144
rect 8556 5244 8572 5382
rect 9195 5382 9291 5398
rect 8735 5360 9057 5361
rect 8735 5244 8736 5360
rect 8556 5144 8736 5244
rect 8556 5012 8578 5144
rect 8735 5040 8736 5144
rect 9056 5244 9057 5360
rect 9195 5244 9211 5382
rect 9056 5144 9211 5244
rect 9056 5040 9057 5144
rect 8735 5039 9057 5040
rect 6310 4698 6410 4996
rect 6688 4790 8232 4890
rect 6310 4682 6415 4698
rect 5859 4660 6181 4661
rect 5859 4340 5860 4660
rect 6180 4554 6181 4660
rect 6310 4554 6335 4682
rect 6180 4454 6335 4554
rect 6180 4340 6181 4454
rect 6310 4340 6335 4454
rect 5859 4339 6181 4340
rect 6319 4314 6335 4340
rect 6399 4314 6415 4682
rect 6688 4661 6788 4790
rect 7038 4682 7134 4698
rect 6578 4660 6900 4661
rect 6578 4340 6579 4660
rect 6899 4340 6900 4660
rect 6578 4339 6900 4340
rect 6319 4294 6415 4314
rect 6688 4198 6788 4339
rect 7038 4314 7054 4682
rect 7118 4314 7134 4682
rect 7408 4661 7508 4790
rect 7757 4682 7853 4698
rect 7297 4660 7619 4661
rect 7297 4340 7298 4660
rect 7618 4340 7619 4660
rect 7297 4339 7619 4340
rect 7038 4294 7134 4314
rect 7408 4198 7508 4339
rect 7757 4314 7773 4682
rect 7837 4314 7853 4682
rect 8130 4661 8231 4790
rect 8476 4682 8578 5012
rect 8016 4660 8338 4661
rect 8016 4340 8017 4660
rect 8337 4340 8338 4660
rect 8016 4339 8338 4340
rect 7757 4294 7853 4314
rect 8130 4198 8231 4339
rect 8476 4314 8492 4682
rect 8556 4550 8578 4682
rect 8850 4661 8950 5039
rect 9188 5012 9211 5144
rect 9275 5012 9291 5382
rect 9188 4682 9291 5012
rect 8735 4660 9057 4661
rect 8735 4550 8736 4660
rect 8556 4450 8736 4550
rect 8556 4314 8578 4450
rect 8735 4340 8736 4450
rect 9056 4550 9057 4660
rect 9188 4550 9211 4682
rect 9056 4450 9211 4550
rect 9056 4340 9057 4450
rect 8735 4339 9057 4340
rect 8850 4338 8950 4339
rect 8476 4300 8578 4314
rect 9188 4314 9211 4450
rect 9275 4314 9291 4682
rect 9188 4300 9291 4314
rect 8476 4294 8572 4300
rect 9195 4294 9291 4300
rect 5498 4197 9450 4198
rect 5498 4099 5499 4197
rect 5597 4099 9450 4197
rect 5498 4098 9450 4099
rect 6319 3982 6415 3998
rect 6319 3962 6335 3982
rect 5974 3961 6074 3962
rect 5859 3960 6181 3961
rect 5859 3640 5860 3960
rect 6180 3852 6181 3960
rect 6310 3852 6335 3962
rect 6180 3752 6335 3852
rect 6180 3640 6181 3752
rect 5859 3639 6181 3640
rect 5974 3261 6074 3639
rect 6310 3614 6335 3752
rect 6399 3614 6415 3982
rect 6688 3961 6788 4098
rect 7038 3982 7134 3998
rect 6578 3960 6900 3961
rect 6578 3640 6579 3960
rect 6899 3640 6900 3960
rect 6578 3639 6900 3640
rect 6310 3596 6415 3614
rect 6310 3298 6410 3596
rect 6688 3496 6788 3639
rect 7038 3614 7054 3982
rect 7118 3614 7134 3982
rect 7408 3961 7508 4098
rect 7757 3982 7853 3998
rect 7297 3960 7619 3961
rect 7297 3640 7298 3960
rect 7618 3640 7619 3960
rect 7297 3639 7619 3640
rect 7038 3596 7134 3614
rect 7408 3496 7508 3639
rect 7757 3614 7773 3982
rect 7837 3614 7853 3982
rect 8130 3961 8231 4098
rect 8478 3998 8578 4000
rect 8476 3982 8578 3998
rect 8016 3960 8338 3961
rect 8016 3640 8017 3960
rect 8337 3640 8338 3960
rect 8016 3639 8338 3640
rect 7757 3596 7853 3614
rect 8130 3496 8231 3639
rect 8476 3614 8492 3982
rect 8556 3846 8578 3982
rect 9188 3998 9288 4000
rect 9188 3982 9291 3998
rect 8850 3961 8950 3962
rect 8735 3960 9057 3961
rect 8735 3846 8736 3960
rect 8556 3746 8736 3846
rect 8556 3614 8578 3746
rect 8735 3640 8736 3746
rect 9056 3846 9057 3960
rect 9188 3846 9211 3982
rect 9056 3746 9211 3846
rect 9056 3640 9057 3746
rect 8735 3639 9057 3640
rect 8476 3596 8578 3614
rect 6688 3396 8231 3496
rect 6310 3282 6415 3298
rect 5859 3260 6181 3261
rect 5859 2940 5860 3260
rect 6180 3146 6181 3260
rect 6310 3146 6335 3282
rect 6180 3046 6335 3146
rect 6180 2940 6181 3046
rect 5859 2939 6181 2940
rect 5974 2561 6074 2939
rect 6310 2914 6335 3046
rect 6399 2914 6415 3282
rect 6688 3261 6788 3396
rect 7038 3282 7134 3298
rect 6578 3260 6900 3261
rect 6578 2940 6579 3260
rect 6899 2940 6900 3260
rect 6578 2939 6900 2940
rect 6310 2896 6415 2914
rect 6310 2598 6410 2896
rect 6688 2796 6788 2939
rect 7038 2914 7054 3282
rect 7118 2914 7134 3282
rect 7408 3261 7508 3396
rect 7757 3282 7853 3298
rect 7297 3260 7619 3261
rect 7297 2940 7298 3260
rect 7618 2940 7619 3260
rect 7297 2939 7619 2940
rect 7038 2896 7134 2914
rect 7408 2796 7508 2939
rect 7757 2914 7773 3282
rect 7837 2914 7853 3282
rect 8130 3261 8231 3396
rect 8478 3298 8578 3596
rect 8476 3282 8578 3298
rect 8016 3260 8338 3261
rect 8016 2940 8017 3260
rect 8337 2940 8338 3260
rect 8016 2939 8338 2940
rect 7757 2896 7853 2914
rect 8130 2796 8231 2939
rect 8476 2914 8492 3282
rect 8556 3154 8578 3282
rect 8850 3261 8950 3639
rect 9188 3614 9211 3746
rect 9275 3614 9291 3982
rect 9188 3596 9291 3614
rect 9188 3298 9288 3596
rect 9188 3282 9291 3298
rect 8735 3260 9057 3261
rect 8735 3154 8736 3260
rect 8556 3054 8736 3154
rect 8556 2914 8578 3054
rect 8735 2940 8736 3054
rect 9056 3154 9057 3260
rect 9188 3154 9211 3282
rect 9056 3054 9211 3154
rect 9056 2940 9057 3054
rect 8735 2939 9057 2940
rect 6688 2696 8232 2796
rect 6310 2582 6415 2598
rect 5859 2560 6181 2561
rect 5859 2500 5860 2560
rect -5100 2448 5860 2500
rect -5100 2362 -4630 2448
rect -4534 2362 -4050 2448
rect -3954 2362 -3450 2448
rect -3354 2362 -2850 2448
rect -2754 2362 -2250 2448
rect -2154 2362 -1650 2448
rect -1554 2362 -1050 2448
rect -954 2362 -450 2448
rect -354 2362 150 2448
rect 246 2362 750 2448
rect 846 2362 1350 2448
rect 1446 2362 1950 2448
rect 2046 2362 2550 2448
rect 2646 2362 3150 2448
rect 3246 2362 3750 2448
rect 3846 2362 4350 2448
rect 4446 2362 4950 2448
rect 5046 2362 5860 2448
rect -5100 2240 5860 2362
rect 6180 2500 6181 2560
rect 6310 2500 6335 2582
rect 6180 2240 6335 2500
rect -5100 2214 6335 2240
rect 6399 2500 6415 2582
rect 7038 2582 7134 2598
rect 6578 2560 6900 2561
rect 6578 2500 6579 2560
rect 6399 2240 6579 2500
rect 6899 2500 6900 2560
rect 7038 2500 7054 2582
rect 6899 2240 7054 2500
rect 6399 2214 7054 2240
rect 7118 2500 7134 2582
rect 7757 2582 7853 2598
rect 7297 2560 7619 2561
rect 7297 2500 7298 2560
rect 7118 2240 7298 2500
rect 7618 2500 7619 2560
rect 7757 2500 7773 2582
rect 7618 2240 7773 2500
rect 7118 2214 7773 2240
rect 7837 2500 7853 2582
rect 8476 2582 8578 2914
rect 8016 2560 8338 2561
rect 8016 2500 8017 2560
rect 7837 2240 8017 2500
rect 8337 2500 8338 2560
rect 8476 2500 8492 2582
rect 8337 2240 8492 2500
rect 7837 2214 8492 2240
rect 8556 2500 8578 2582
rect 8850 2561 8950 2939
rect 9188 2914 9211 3054
rect 9275 2914 9291 3282
rect 9188 2582 9291 2914
rect 8735 2560 9057 2561
rect 8735 2500 8736 2560
rect 8556 2240 8736 2500
rect 9056 2500 9057 2560
rect 9188 2500 9211 2582
rect 9056 2240 9211 2500
rect 8556 2214 9211 2240
rect 9275 2500 9291 2582
rect 9275 2214 9448 2500
rect -5100 2184 9448 2214
rect -5100 1884 -4916 2184
rect -4316 1884 4716 2184
rect 5316 1884 9448 2184
rect -5100 1700 9448 1884
rect 8478 1696 8578 1700
<< labels >>
flabel metal4 -2300 2102 -2280 2122 1 FreeSans 480 0 0 0 VSS
port 6 n ground bidirectional
flabel metal4 -2534 10006 -2500 10030 1 FreeSans 480 0 0 0 VDD
port 5 n power bidirectional
flabel metal2 -3700 4356 -3686 4370 1 FreeSans 480 0 0 0 vin
port 2 n
flabel metal1 -3698 2662 -3690 2672 1 FreeSans 480 0 0 0 vbiasn
port 3 n
flabel metal2 -3228 7078 -3218 7084 1 FreeSans 480 0 0 0 vbiasp
port 4 n
flabel metal2 4126 4350 4138 4364 1 FreeSans 480 0 0 0 voutcs
flabel metal2 4532 4380 4544 4390 1 FreeSans 480 0 0 0 vout
port 1 n
flabel metal1 -4134 3252 -4122 3270 1 FreeSans 480 0 0 0 csinvn
flabel metal2 -3584 6480 -3574 6494 1 FreeSans 480 0 0 0 csinvp
<< end >>
