magic
tech sky130A
magscale 1 2
timestamp 1624494425
<< locali >>
rect 4857 101022 6363 101056
rect 7680 100983 8257 101017
rect 5497 100910 6253 100944
rect 6137 100820 6363 100854
rect 6137 100596 6363 100630
rect 5497 100506 6253 100540
rect 7680 100433 8257 100467
rect 4777 100394 6363 100428
rect 4697 100232 6363 100266
rect 7680 100193 8257 100227
rect 5497 100120 6253 100154
rect 6137 100030 6363 100064
rect 6137 99806 6363 99840
rect 5497 99716 6253 99750
rect 7680 99643 8257 99677
rect 4617 99604 6363 99638
rect 4857 99442 6363 99476
rect 7680 99403 8257 99437
rect 5417 99330 6253 99364
rect 6137 99240 6363 99274
rect 6137 99016 6363 99050
rect 5417 98926 6253 98960
rect 7680 98853 8257 98887
rect 4777 98814 6363 98848
rect 4697 98652 6363 98686
rect 7680 98613 8257 98647
rect 5417 98540 6253 98574
rect 6137 98450 6363 98484
rect 6137 98226 6363 98260
rect 5417 98136 6253 98170
rect 7680 98063 8257 98097
rect 4617 98024 6363 98058
rect 4857 97862 6363 97896
rect 7680 97823 8257 97857
rect 5337 97750 6253 97784
rect 6137 97660 6363 97694
rect 6137 97436 6363 97470
rect 5337 97346 6253 97380
rect 7680 97273 8257 97307
rect 4777 97234 6363 97268
rect 4697 97072 6363 97106
rect 7680 97033 8257 97067
rect 5337 96960 6253 96994
rect 6137 96870 6363 96904
rect 6137 96646 6363 96680
rect 5337 96556 6253 96590
rect 7680 96483 8257 96517
rect 4617 96444 6363 96478
rect 4857 96282 6363 96316
rect 7680 96243 8257 96277
rect 5257 96170 6253 96204
rect 6137 96080 6363 96114
rect 6137 95856 6363 95890
rect 5257 95766 6253 95800
rect 7680 95693 8257 95727
rect 4777 95654 6363 95688
rect 4697 95492 6363 95526
rect 7680 95453 8257 95487
rect 5257 95380 6253 95414
rect 6137 95290 6363 95324
rect 6137 95066 6363 95100
rect 5257 94976 6253 95010
rect 7680 94903 8257 94937
rect 4617 94864 6363 94898
rect 4857 94702 6363 94736
rect 7680 94663 8257 94697
rect 5177 94590 6253 94624
rect 6137 94500 6363 94534
rect 6137 94276 6363 94310
rect 5177 94186 6253 94220
rect 7680 94113 8257 94147
rect 4777 94074 6363 94108
rect 4697 93912 6363 93946
rect 7680 93873 8257 93907
rect 5177 93800 6253 93834
rect 6137 93710 6363 93744
rect 6137 93486 6363 93520
rect 5177 93396 6253 93430
rect 7680 93323 8257 93357
rect 4617 93284 6363 93318
rect 4857 93122 6363 93156
rect 7680 93083 8257 93117
rect 5097 93010 6253 93044
rect 6137 92920 6363 92954
rect 6137 92696 6363 92730
rect 5097 92606 6253 92640
rect 7680 92533 8257 92567
rect 4777 92494 6363 92528
rect 4697 92332 6363 92366
rect 7680 92293 8257 92327
rect 5097 92220 6253 92254
rect 6137 92130 6363 92164
rect 6137 91906 6363 91940
rect 5097 91816 6253 91850
rect 7680 91743 8257 91777
rect 4617 91704 6363 91738
rect 4857 91542 6363 91576
rect 7680 91503 8257 91537
rect 5017 91430 6253 91464
rect 6137 91340 6363 91374
rect 6137 91116 6363 91150
rect 5017 91026 6253 91060
rect 7680 90953 8257 90987
rect 4777 90914 6363 90948
rect 4697 90752 6363 90786
rect 7680 90713 8257 90747
rect 5017 90640 6253 90674
rect 6137 90550 6363 90584
rect 6137 90326 6363 90360
rect 5017 90236 6253 90270
rect 7680 90163 8257 90197
rect 4617 90124 6363 90158
rect 4857 89962 6363 89996
rect 7680 89923 8257 89957
rect 4937 89850 6253 89884
rect 6137 89760 6363 89794
rect 6137 89536 6363 89570
rect 4937 89446 6253 89480
rect 7680 89373 8257 89407
rect 4777 89334 6363 89368
rect 4697 89172 6363 89206
rect 7680 89133 8257 89167
rect 4937 89060 6253 89094
rect 6137 88970 6363 89004
rect 6137 88746 6363 88780
rect 4937 88656 6253 88690
rect 7680 88583 8257 88617
rect 4617 88544 6363 88578
rect 4857 88382 6363 88416
rect 7680 88343 8257 88377
rect 5497 88270 6253 88304
rect 6057 88180 6363 88214
rect 6057 87956 6363 87990
rect 5497 87866 6253 87900
rect 7680 87793 8257 87827
rect 4777 87754 6363 87788
rect 4697 87592 6363 87626
rect 7680 87553 8257 87587
rect 5497 87480 6253 87514
rect 6057 87390 6363 87424
rect 6057 87166 6363 87200
rect 5497 87076 6253 87110
rect 7680 87003 8257 87037
rect 4617 86964 6363 86998
rect 4857 86802 6363 86836
rect 7680 86763 8257 86797
rect 5417 86690 6253 86724
rect 6057 86600 6363 86634
rect 6057 86376 6363 86410
rect 5417 86286 6253 86320
rect 7680 86213 8257 86247
rect 4777 86174 6363 86208
rect 4697 86012 6363 86046
rect 7680 85973 8257 86007
rect 5417 85900 6253 85934
rect 6057 85810 6363 85844
rect 6057 85586 6363 85620
rect 5417 85496 6253 85530
rect 7680 85423 8257 85457
rect 4617 85384 6363 85418
rect 4857 85222 6363 85256
rect 7680 85183 8257 85217
rect 5337 85110 6253 85144
rect 6057 85020 6363 85054
rect 6057 84796 6363 84830
rect 5337 84706 6253 84740
rect 7680 84633 8257 84667
rect 4777 84594 6363 84628
rect 4697 84432 6363 84466
rect 7680 84393 8257 84427
rect 5337 84320 6253 84354
rect 6057 84230 6363 84264
rect 6057 84006 6363 84040
rect 5337 83916 6253 83950
rect 7680 83843 8257 83877
rect 4617 83804 6363 83838
rect 4857 83642 6363 83676
rect 7680 83603 8257 83637
rect 5257 83530 6253 83564
rect 6057 83440 6363 83474
rect 6057 83216 6363 83250
rect 5257 83126 6253 83160
rect 7680 83053 8257 83087
rect 4777 83014 6363 83048
rect 4697 82852 6363 82886
rect 7680 82813 8257 82847
rect 5257 82740 6253 82774
rect 6057 82650 6363 82684
rect 6057 82426 6363 82460
rect 5257 82336 6253 82370
rect 7680 82263 8257 82297
rect 4617 82224 6363 82258
rect 4857 82062 6363 82096
rect 7680 82023 8257 82057
rect 5177 81950 6253 81984
rect 6057 81860 6363 81894
rect 6057 81636 6363 81670
rect 5177 81546 6253 81580
rect 7680 81473 8257 81507
rect 4777 81434 6363 81468
rect 4697 81272 6363 81306
rect 7680 81233 8257 81267
rect 5177 81160 6253 81194
rect 6057 81070 6363 81104
rect 6057 80846 6363 80880
rect 5177 80756 6253 80790
rect 7680 80683 8257 80717
rect 4617 80644 6363 80678
rect 4857 80482 6363 80516
rect 7680 80443 8257 80477
rect 5097 80370 6253 80404
rect 6057 80280 6363 80314
rect 6057 80056 6363 80090
rect 5097 79966 6253 80000
rect 7680 79893 8257 79927
rect 4777 79854 6363 79888
rect 4697 79692 6363 79726
rect 7680 79653 8257 79687
rect 5097 79580 6253 79614
rect 6057 79490 6363 79524
rect 6057 79266 6363 79300
rect 5097 79176 6253 79210
rect 7680 79103 8257 79137
rect 4617 79064 6363 79098
rect 4857 78902 6363 78936
rect 7680 78863 8257 78897
rect 5017 78790 6253 78824
rect 6057 78700 6363 78734
rect 6057 78476 6363 78510
rect 5017 78386 6253 78420
rect 7680 78313 8257 78347
rect 4777 78274 6363 78308
rect 4697 78112 6363 78146
rect 7680 78073 8257 78107
rect 5017 78000 6253 78034
rect 6057 77910 6363 77944
rect 6057 77686 6363 77720
rect 5017 77596 6253 77630
rect 7680 77523 8257 77557
rect 4617 77484 6363 77518
rect 4857 77322 6363 77356
rect 7680 77283 8257 77317
rect 4937 77210 6253 77244
rect 6057 77120 6363 77154
rect 6057 76896 6363 76930
rect 4937 76806 6253 76840
rect 7680 76733 8257 76767
rect 4777 76694 6363 76728
rect 4697 76532 6363 76566
rect 7680 76493 8257 76527
rect 4937 76420 6253 76454
rect 6057 76330 6363 76364
rect 6057 76106 6363 76140
rect 4937 76016 6253 76050
rect 7680 75943 8257 75977
rect 4617 75904 6363 75938
rect 4857 75742 6363 75776
rect 7680 75703 8257 75737
rect 5497 75630 6253 75664
rect 5977 75540 6363 75574
rect 5977 75316 6363 75350
rect 5497 75226 6253 75260
rect 7680 75153 8257 75187
rect 4777 75114 6363 75148
rect 4697 74952 6363 74986
rect 7680 74913 8257 74947
rect 5497 74840 6253 74874
rect 5977 74750 6363 74784
rect 5977 74526 6363 74560
rect 5497 74436 6253 74470
rect 7680 74363 8257 74397
rect 4617 74324 6363 74358
rect 4857 74162 6363 74196
rect 7680 74123 8257 74157
rect 5417 74050 6253 74084
rect 5977 73960 6363 73994
rect 5977 73736 6363 73770
rect 5417 73646 6253 73680
rect 7680 73573 8257 73607
rect 4777 73534 6363 73568
rect 4697 73372 6363 73406
rect 7680 73333 8257 73367
rect 5417 73260 6253 73294
rect 5977 73170 6363 73204
rect 5977 72946 6363 72980
rect 5417 72856 6253 72890
rect 7680 72783 8257 72817
rect 4617 72744 6363 72778
rect 4857 72582 6363 72616
rect 7680 72543 8257 72577
rect 5337 72470 6253 72504
rect 5977 72380 6363 72414
rect 5977 72156 6363 72190
rect 5337 72066 6253 72100
rect 7680 71993 8257 72027
rect 4777 71954 6363 71988
rect 4697 71792 6363 71826
rect 7680 71753 8257 71787
rect 5337 71680 6253 71714
rect 5977 71590 6363 71624
rect 5977 71366 6363 71400
rect 5337 71276 6253 71310
rect 7680 71203 8257 71237
rect 4617 71164 6363 71198
rect 4857 71002 6363 71036
rect 7680 70963 8257 70997
rect 5257 70890 6253 70924
rect 5977 70800 6363 70834
rect 5977 70576 6363 70610
rect 5257 70486 6253 70520
rect 7680 70413 8257 70447
rect 4777 70374 6363 70408
rect 4697 70212 6363 70246
rect 7680 70173 8257 70207
rect 5257 70100 6253 70134
rect 5977 70010 6363 70044
rect 5977 69786 6363 69820
rect 5257 69696 6253 69730
rect 7680 69623 8257 69657
rect 4617 69584 6363 69618
rect 4857 69422 6363 69456
rect 7680 69383 8257 69417
rect 5177 69310 6253 69344
rect 5977 69220 6363 69254
rect 5977 68996 6363 69030
rect 5177 68906 6253 68940
rect 7680 68833 8257 68867
rect 4777 68794 6363 68828
rect 4697 68632 6363 68666
rect 7680 68593 8257 68627
rect 5177 68520 6253 68554
rect 5977 68430 6363 68464
rect 5977 68206 6363 68240
rect 5177 68116 6253 68150
rect 7680 68043 8257 68077
rect 4617 68004 6363 68038
rect 4857 67842 6363 67876
rect 7680 67803 8257 67837
rect 5097 67730 6253 67764
rect 5977 67640 6363 67674
rect 5977 67416 6363 67450
rect 5097 67326 6253 67360
rect 7680 67253 8257 67287
rect 4777 67214 6363 67248
rect 4697 67052 6363 67086
rect 7680 67013 8257 67047
rect 5097 66940 6253 66974
rect 5977 66850 6363 66884
rect 5977 66626 6363 66660
rect 5097 66536 6253 66570
rect 7680 66463 8257 66497
rect 4617 66424 6363 66458
rect 4857 66262 6363 66296
rect 7680 66223 8257 66257
rect 5017 66150 6253 66184
rect 5977 66060 6363 66094
rect 5977 65836 6363 65870
rect 5017 65746 6253 65780
rect 7680 65673 8257 65707
rect 4777 65634 6363 65668
rect 4697 65472 6363 65506
rect 7680 65433 8257 65467
rect 5017 65360 6253 65394
rect 5977 65270 6363 65304
rect 5977 65046 6363 65080
rect 5017 64956 6253 64990
rect 7680 64883 8257 64917
rect 4617 64844 6363 64878
rect 4857 64682 6363 64716
rect 7680 64643 8257 64677
rect 4937 64570 6253 64604
rect 5977 64480 6363 64514
rect 5977 64256 6363 64290
rect 4937 64166 6253 64200
rect 7680 64093 8257 64127
rect 4777 64054 6363 64088
rect 4697 63892 6363 63926
rect 7680 63853 8257 63887
rect 4937 63780 6253 63814
rect 5977 63690 6363 63724
rect 5977 63466 6363 63500
rect 4937 63376 6253 63410
rect 7680 63303 8257 63337
rect 4617 63264 6363 63298
rect 4857 63102 6363 63136
rect 7680 63063 8257 63097
rect 5497 62990 6253 63024
rect 5897 62900 6363 62934
rect 5897 62676 6363 62710
rect 5497 62586 6253 62620
rect 7680 62513 8257 62547
rect 4777 62474 6363 62508
rect 4697 62312 6363 62346
rect 7680 62273 8257 62307
rect 5497 62200 6253 62234
rect 5897 62110 6363 62144
rect 5897 61886 6363 61920
rect 5497 61796 6253 61830
rect 7680 61723 8257 61757
rect 4617 61684 6363 61718
rect 4857 61522 6363 61556
rect 7680 61483 8257 61517
rect 5417 61410 6253 61444
rect 5897 61320 6363 61354
rect 5897 61096 6363 61130
rect 5417 61006 6253 61040
rect 7680 60933 8257 60967
rect 4777 60894 6363 60928
rect 4697 60732 6363 60766
rect 7680 60693 8257 60727
rect 5417 60620 6253 60654
rect 5897 60530 6363 60564
rect 5897 60306 6363 60340
rect 5417 60216 6253 60250
rect 7680 60143 8257 60177
rect 4617 60104 6363 60138
rect 4857 59942 6363 59976
rect 7680 59903 8257 59937
rect 5337 59830 6253 59864
rect 5897 59740 6363 59774
rect 5897 59516 6363 59550
rect 5337 59426 6253 59460
rect 7680 59353 8257 59387
rect 4777 59314 6363 59348
rect 4697 59152 6363 59186
rect 7680 59113 8257 59147
rect 5337 59040 6253 59074
rect 5897 58950 6363 58984
rect 5897 58726 6363 58760
rect 5337 58636 6253 58670
rect 7680 58563 8257 58597
rect 4617 58524 6363 58558
rect 4857 58362 6363 58396
rect 7680 58323 8257 58357
rect 5257 58250 6253 58284
rect 5897 58160 6363 58194
rect 5897 57936 6363 57970
rect 5257 57846 6253 57880
rect 7680 57773 8257 57807
rect 4777 57734 6363 57768
rect 4697 57572 6363 57606
rect 7680 57533 8257 57567
rect 5257 57460 6253 57494
rect 5897 57370 6363 57404
rect 5897 57146 6363 57180
rect 5257 57056 6253 57090
rect 7680 56983 8257 57017
rect 4617 56944 6363 56978
rect 4857 56782 6363 56816
rect 7680 56743 8257 56777
rect 5177 56670 6253 56704
rect 5897 56580 6363 56614
rect 5897 56356 6363 56390
rect 5177 56266 6253 56300
rect 7680 56193 8257 56227
rect 4777 56154 6363 56188
rect 4697 55992 6363 56026
rect 7680 55953 8257 55987
rect 5177 55880 6253 55914
rect 5897 55790 6363 55824
rect 5897 55566 6363 55600
rect 5177 55476 6253 55510
rect 7680 55403 8257 55437
rect 4617 55364 6363 55398
rect 4857 55202 6363 55236
rect 7680 55163 8257 55197
rect 5097 55090 6253 55124
rect 5897 55000 6363 55034
rect 5897 54776 6363 54810
rect 5097 54686 6253 54720
rect 7680 54613 8257 54647
rect 4777 54574 6363 54608
rect 4697 54412 6363 54446
rect 7680 54373 8257 54407
rect 5097 54300 6253 54334
rect 5897 54210 6363 54244
rect 5897 53986 6363 54020
rect 5097 53896 6253 53930
rect 7680 53823 8257 53857
rect 4617 53784 6363 53818
rect 4857 53622 6363 53656
rect 7680 53583 8257 53617
rect 5017 53510 6253 53544
rect 5897 53420 6363 53454
rect 5897 53196 6363 53230
rect 5017 53106 6253 53140
rect 7680 53033 8257 53067
rect 4777 52994 6363 53028
rect 4697 52832 6363 52866
rect 7680 52793 8257 52827
rect 5017 52720 6253 52754
rect 5897 52630 6363 52664
rect 5897 52406 6363 52440
rect 5017 52316 6253 52350
rect 7680 52243 8257 52277
rect 4617 52204 6363 52238
rect 4857 52042 6363 52076
rect 7680 52003 8257 52037
rect 4937 51930 6253 51964
rect 5897 51840 6363 51874
rect 5897 51616 6363 51650
rect 4937 51526 6253 51560
rect 7680 51453 8257 51487
rect 4777 51414 6363 51448
rect 4697 51252 6363 51286
rect 7680 51213 8257 51247
rect 4937 51140 6253 51174
rect 5897 51050 6363 51084
rect 5897 50826 6363 50860
rect 4937 50736 6253 50770
rect 7680 50663 8257 50697
rect 4617 50624 6363 50658
rect 4857 50462 6363 50496
rect 7680 50423 8257 50457
rect 5497 50350 6253 50384
rect 5817 50260 6363 50294
rect 5817 50036 6363 50070
rect 5497 49946 6253 49980
rect 7680 49873 8257 49907
rect 4777 49834 6363 49868
rect 4697 49672 6363 49706
rect 7680 49633 8257 49667
rect 5497 49560 6253 49594
rect 5817 49470 6363 49504
rect 5817 49246 6363 49280
rect 5497 49156 6253 49190
rect 7680 49083 8257 49117
rect 4617 49044 6363 49078
rect 4857 48882 6363 48916
rect 7680 48843 8257 48877
rect 5417 48770 6253 48804
rect 5817 48680 6363 48714
rect 5817 48456 6363 48490
rect 5417 48366 6253 48400
rect 7680 48293 8257 48327
rect 4777 48254 6363 48288
rect 4697 48092 6363 48126
rect 7680 48053 8257 48087
rect 5417 47980 6253 48014
rect 5817 47890 6363 47924
rect 5817 47666 6363 47700
rect 5417 47576 6253 47610
rect 7680 47503 8257 47537
rect 4617 47464 6363 47498
rect 4857 47302 6363 47336
rect 7680 47263 8257 47297
rect 5337 47190 6253 47224
rect 5817 47100 6363 47134
rect 5817 46876 6363 46910
rect 5337 46786 6253 46820
rect 7680 46713 8257 46747
rect 4777 46674 6363 46708
rect 4697 46512 6363 46546
rect 7680 46473 8257 46507
rect 5337 46400 6253 46434
rect 5817 46310 6363 46344
rect 5817 46086 6363 46120
rect 5337 45996 6253 46030
rect 7680 45923 8257 45957
rect 4617 45884 6363 45918
rect 4857 45722 6363 45756
rect 7680 45683 8257 45717
rect 5257 45610 6253 45644
rect 5817 45520 6363 45554
rect 5817 45296 6363 45330
rect 5257 45206 6253 45240
rect 7680 45133 8257 45167
rect 4777 45094 6363 45128
rect 4697 44932 6363 44966
rect 7680 44893 8257 44927
rect 5257 44820 6253 44854
rect 5817 44730 6363 44764
rect 5817 44506 6363 44540
rect 5257 44416 6253 44450
rect 7680 44343 8257 44377
rect 4617 44304 6363 44338
rect 4857 44142 6363 44176
rect 7680 44103 8257 44137
rect 5177 44030 6253 44064
rect 5817 43940 6363 43974
rect 5817 43716 6363 43750
rect 5177 43626 6253 43660
rect 7680 43553 8257 43587
rect 4777 43514 6363 43548
rect 4697 43352 6363 43386
rect 7680 43313 8257 43347
rect 5177 43240 6253 43274
rect 5817 43150 6363 43184
rect 5817 42926 6363 42960
rect 5177 42836 6253 42870
rect 7680 42763 8257 42797
rect 4617 42724 6363 42758
rect 4857 42562 6363 42596
rect 7680 42523 8257 42557
rect 5097 42450 6253 42484
rect 5817 42360 6363 42394
rect 5817 42136 6363 42170
rect 5097 42046 6253 42080
rect 7680 41973 8257 42007
rect 4777 41934 6363 41968
rect 4697 41772 6363 41806
rect 7680 41733 8257 41767
rect 5097 41660 6253 41694
rect 5817 41570 6363 41604
rect 5817 41346 6363 41380
rect 5097 41256 6253 41290
rect 7680 41183 8257 41217
rect 4617 41144 6363 41178
rect 4857 40982 6363 41016
rect 7680 40943 8257 40977
rect 5017 40870 6253 40904
rect 5817 40780 6363 40814
rect 5817 40556 6363 40590
rect 5017 40466 6253 40500
rect 7680 40393 8257 40427
rect 4777 40354 6363 40388
rect 4697 40192 6363 40226
rect 7680 40153 8257 40187
rect 5017 40080 6253 40114
rect 5817 39990 6363 40024
rect 5817 39766 6363 39800
rect 5017 39676 6253 39710
rect 7680 39603 8257 39637
rect 4617 39564 6363 39598
rect 4857 39402 6363 39436
rect 7680 39363 8257 39397
rect 4937 39290 6253 39324
rect 5817 39200 6363 39234
rect 5817 38976 6363 39010
rect 4937 38886 6253 38920
rect 7680 38813 8257 38847
rect 4777 38774 6363 38808
rect 4697 38612 6363 38646
rect 7680 38573 8257 38607
rect 4937 38500 6253 38534
rect 5817 38410 6363 38444
rect 5817 38186 6363 38220
rect 4937 38096 6253 38130
rect 7680 38023 8257 38057
rect 4617 37984 6363 38018
rect 4857 37822 6363 37856
rect 7680 37783 8257 37817
rect 5497 37710 6253 37744
rect 5737 37620 6363 37654
rect 5737 37396 6363 37430
rect 5497 37306 6253 37340
rect 7680 37233 8257 37267
rect 4777 37194 6363 37228
rect 4697 37032 6363 37066
rect 7680 36993 8257 37027
rect 5497 36920 6253 36954
rect 5737 36830 6363 36864
rect 5737 36606 6363 36640
rect 5497 36516 6253 36550
rect 7680 36443 8257 36477
rect 4617 36404 6363 36438
rect 4857 36242 6363 36276
rect 7680 36203 8257 36237
rect 5417 36130 6253 36164
rect 5737 36040 6363 36074
rect 5737 35816 6363 35850
rect 5417 35726 6253 35760
rect 7680 35653 8257 35687
rect 4777 35614 6363 35648
rect 4697 35452 6363 35486
rect 7680 35413 8257 35447
rect 5417 35340 6253 35374
rect 5737 35250 6363 35284
rect 5737 35026 6363 35060
rect 5417 34936 6253 34970
rect 7680 34863 8257 34897
rect 4617 34824 6363 34858
rect 4857 34662 6363 34696
rect 7680 34623 8257 34657
rect 5337 34550 6253 34584
rect 5737 34460 6363 34494
rect 5737 34236 6363 34270
rect 5337 34146 6253 34180
rect 7680 34073 8257 34107
rect 4777 34034 6363 34068
rect 4697 33872 6363 33906
rect 7680 33833 8257 33867
rect 5337 33760 6253 33794
rect 5737 33670 6363 33704
rect 5737 33446 6363 33480
rect 5337 33356 6253 33390
rect 7680 33283 8257 33317
rect 4617 33244 6363 33278
rect 4857 33082 6363 33116
rect 7680 33043 8257 33077
rect 5257 32970 6253 33004
rect 5737 32880 6363 32914
rect 5737 32656 6363 32690
rect 5257 32566 6253 32600
rect 7680 32493 8257 32527
rect 4777 32454 6363 32488
rect 4697 32292 6363 32326
rect 7680 32253 8257 32287
rect 5257 32180 6253 32214
rect 5737 32090 6363 32124
rect 5737 31866 6363 31900
rect 5257 31776 6253 31810
rect 7680 31703 8257 31737
rect 4617 31664 6363 31698
rect 4857 31502 6363 31536
rect 7680 31463 8257 31497
rect 5177 31390 6253 31424
rect 5737 31300 6363 31334
rect 5737 31076 6363 31110
rect 5177 30986 6253 31020
rect 7680 30913 8257 30947
rect 4777 30874 6363 30908
rect 4697 30712 6363 30746
rect 7680 30673 8257 30707
rect 5177 30600 6253 30634
rect 5737 30510 6363 30544
rect 5737 30286 6363 30320
rect 5177 30196 6253 30230
rect 7680 30123 8257 30157
rect 4617 30084 6363 30118
rect 4857 29922 6363 29956
rect 7680 29883 8257 29917
rect 5097 29810 6253 29844
rect 5737 29720 6363 29754
rect 5737 29496 6363 29530
rect 5097 29406 6253 29440
rect 7680 29333 8257 29367
rect 4777 29294 6363 29328
rect 4697 29132 6363 29166
rect 7680 29093 8257 29127
rect 5097 29020 6253 29054
rect 5737 28930 6363 28964
rect 5737 28706 6363 28740
rect 5097 28616 6253 28650
rect 7680 28543 8257 28577
rect 4617 28504 6363 28538
rect 4857 28342 6363 28376
rect 7680 28303 8257 28337
rect 5017 28230 6253 28264
rect 5737 28140 6363 28174
rect 5737 27916 6363 27950
rect 5017 27826 6253 27860
rect 7680 27753 8257 27787
rect 4777 27714 6363 27748
rect 4697 27552 6363 27586
rect 7680 27513 8257 27547
rect 5017 27440 6253 27474
rect 5737 27350 6363 27384
rect 5737 27126 6363 27160
rect 5017 27036 6253 27070
rect 7680 26963 8257 26997
rect 4617 26924 6363 26958
rect 4857 26762 6363 26796
rect 7680 26723 8257 26757
rect 4937 26650 6253 26684
rect 5737 26560 6363 26594
rect 5737 26336 6363 26370
rect 4937 26246 6253 26280
rect 7680 26173 8257 26207
rect 4777 26134 6363 26168
rect 4697 25972 6363 26006
rect 7680 25933 8257 25967
rect 4937 25860 6253 25894
rect 5737 25770 6363 25804
rect 5737 25546 6363 25580
rect 4937 25456 6253 25490
rect 7680 25383 8257 25417
rect 4617 25344 6363 25378
rect 4857 25182 6363 25216
rect 7680 25143 8257 25177
rect 5497 25070 6253 25104
rect 5657 24980 6363 25014
rect 5657 24756 6363 24790
rect 5497 24666 6253 24700
rect 7680 24593 8257 24627
rect 4777 24554 6363 24588
rect 4697 24392 6363 24426
rect 7680 24353 8257 24387
rect 5497 24280 6253 24314
rect 5657 24190 6363 24224
rect 5657 23966 6363 24000
rect 5497 23876 6253 23910
rect 7680 23803 8257 23837
rect 4617 23764 6363 23798
rect 4857 23602 6363 23636
rect 7680 23563 8257 23597
rect 5417 23490 6253 23524
rect 5657 23400 6363 23434
rect 5657 23176 6363 23210
rect 5417 23086 6253 23120
rect 7680 23013 8257 23047
rect 4777 22974 6363 23008
rect 4697 22812 6363 22846
rect 7680 22773 8257 22807
rect 5417 22700 6253 22734
rect 5657 22610 6363 22644
rect 5657 22386 6363 22420
rect 5417 22296 6253 22330
rect 7680 22223 8257 22257
rect 4617 22184 6363 22218
rect 4857 22022 6363 22056
rect 7680 21983 8257 22017
rect 5337 21910 6253 21944
rect 5657 21820 6363 21854
rect 5657 21596 6363 21630
rect 5337 21506 6253 21540
rect 7680 21433 8257 21467
rect 4777 21394 6363 21428
rect 4697 21232 6363 21266
rect 7680 21193 8257 21227
rect 5337 21120 6253 21154
rect 5657 21030 6363 21064
rect 5657 20806 6363 20840
rect 5337 20716 6253 20750
rect 7680 20643 8257 20677
rect 4617 20604 6363 20638
rect 4857 20442 6363 20476
rect 7680 20403 8257 20437
rect 5257 20330 6253 20364
rect 5657 20240 6363 20274
rect 5657 20016 6363 20050
rect 5257 19926 6253 19960
rect 7680 19853 8257 19887
rect 4777 19814 6363 19848
rect 4697 19652 6363 19686
rect 7680 19613 8257 19647
rect 5257 19540 6253 19574
rect 5657 19450 6363 19484
rect 5657 19226 6363 19260
rect 5257 19136 6253 19170
rect 7680 19063 8257 19097
rect 4617 19024 6363 19058
rect 4857 18862 6363 18896
rect 7680 18823 8257 18857
rect 5177 18750 6253 18784
rect 5657 18660 6363 18694
rect 5657 18436 6363 18470
rect 5177 18346 6253 18380
rect 7680 18273 8257 18307
rect 4777 18234 6363 18268
rect 4697 18072 6363 18106
rect 7680 18033 8257 18067
rect 5177 17960 6253 17994
rect 5657 17870 6363 17904
rect 5657 17646 6363 17680
rect 5177 17556 6253 17590
rect 7680 17483 8257 17517
rect 4617 17444 6363 17478
rect 4857 17282 6363 17316
rect 7680 17243 8257 17277
rect 5097 17170 6253 17204
rect 5657 17080 6363 17114
rect 5657 16856 6363 16890
rect 5097 16766 6253 16800
rect 7680 16693 8257 16727
rect 4777 16654 6363 16688
rect 4697 16492 6363 16526
rect 7680 16453 8257 16487
rect 5097 16380 6253 16414
rect 5657 16290 6363 16324
rect 5657 16066 6363 16100
rect 5097 15976 6253 16010
rect 7680 15903 8257 15937
rect 4617 15864 6363 15898
rect 4857 15702 6363 15736
rect 7680 15663 8257 15697
rect 5017 15590 6253 15624
rect 5657 15500 6363 15534
rect 5657 15276 6363 15310
rect 5017 15186 6253 15220
rect 7680 15113 8257 15147
rect 4777 15074 6363 15108
rect 4697 14912 6363 14946
rect 7680 14873 8257 14907
rect 5017 14800 6253 14834
rect 5657 14710 6363 14744
rect 5657 14486 6363 14520
rect 5017 14396 6253 14430
rect 7680 14323 8257 14357
rect 4617 14284 6363 14318
rect 4857 14122 6363 14156
rect 7680 14083 8257 14117
rect 4937 14010 6253 14044
rect 5657 13920 6363 13954
rect 5657 13696 6363 13730
rect 4937 13606 6253 13640
rect 7680 13533 8257 13567
rect 4777 13494 6363 13528
rect 4697 13332 6363 13366
rect 7680 13293 8257 13327
rect 4937 13220 6253 13254
rect 5657 13130 6363 13164
rect 5657 12906 6363 12940
rect 4937 12816 6253 12850
rect 7680 12743 8257 12777
rect 4617 12704 6363 12738
rect 4857 12542 6363 12576
rect 7680 12503 8257 12537
rect 5497 12430 6253 12464
rect 5577 12340 6363 12374
rect 5577 12116 6363 12150
rect 5497 12026 6253 12060
rect 7680 11953 8257 11987
rect 4777 11914 6363 11948
rect 4697 11752 6363 11786
rect 7680 11713 8257 11747
rect 5497 11640 6253 11674
rect 5577 11550 6363 11584
rect 5577 11326 6363 11360
rect 5497 11236 6253 11270
rect 7680 11163 8257 11197
rect 4617 11124 6363 11158
rect 4857 10962 6363 10996
rect 7680 10923 8257 10957
rect 5417 10850 6253 10884
rect 5577 10760 6363 10794
rect 5577 10536 6363 10570
rect 5417 10446 6253 10480
rect 7680 10373 8257 10407
rect 4777 10334 6363 10368
rect 4697 10172 6363 10206
rect 7680 10133 8257 10167
rect 5417 10060 6253 10094
rect 5577 9970 6363 10004
rect 5577 9746 6363 9780
rect 5417 9656 6253 9690
rect 7680 9583 8257 9617
rect 4617 9544 6363 9578
rect 4857 9382 6363 9416
rect 7680 9343 8257 9377
rect 5337 9270 6253 9304
rect 5577 9180 6363 9214
rect 5577 8956 6363 8990
rect 5337 8866 6253 8900
rect 7680 8793 8257 8827
rect 4777 8754 6363 8788
rect 4697 8592 6363 8626
rect 7680 8553 8257 8587
rect 5337 8480 6253 8514
rect 5577 8390 6363 8424
rect 5577 8166 6363 8200
rect 5337 8076 6253 8110
rect 7680 8003 8257 8037
rect 4617 7964 6363 7998
rect 4857 7802 6363 7836
rect 7680 7763 8257 7797
rect 5257 7690 6253 7724
rect 5577 7600 6363 7634
rect 5577 7376 6363 7410
rect 593 7263 941 7297
rect 5257 7286 6253 7320
rect 7680 7213 8257 7247
rect 4777 7174 6363 7208
rect 4697 7012 6363 7046
rect 7680 6973 8257 7007
rect 513 6923 861 6957
rect 5257 6900 6253 6934
rect 5577 6810 6363 6844
rect 5577 6586 6363 6620
rect 433 6473 781 6507
rect 5257 6496 6253 6530
rect 7680 6423 8257 6457
rect 4617 6384 6363 6418
rect 4857 6222 6363 6256
rect 7680 6183 8257 6217
rect 5177 6110 6253 6144
rect 5577 6020 6363 6054
rect 5577 5796 6363 5830
rect 5177 5706 6253 5740
rect 7680 5633 8257 5667
rect 4777 5594 6363 5628
rect 4697 5432 6363 5466
rect 7680 5393 8257 5427
rect 5177 5320 6253 5354
rect 5577 5230 6363 5264
rect 5577 5006 6363 5040
rect 5177 4916 6253 4950
rect 7680 4843 8257 4877
rect 4617 4804 6363 4838
rect 4857 4642 6363 4676
rect 7680 4603 8257 4637
rect 5097 4530 6253 4564
rect 5577 4440 6363 4474
rect 5577 4216 6363 4250
rect 5097 4126 6253 4160
rect 7680 4053 8257 4087
rect 4777 4014 6363 4048
rect 4697 3852 6363 3886
rect 7680 3813 8257 3847
rect 5097 3740 6253 3774
rect 5577 3650 6363 3684
rect 5577 3426 6363 3460
rect 353 3313 941 3347
rect 5097 3336 6253 3370
rect 7680 3263 8257 3297
rect 4617 3224 6363 3258
rect 4857 3062 6363 3096
rect 7680 3023 8257 3057
rect 273 2973 861 3007
rect 5017 2950 6253 2984
rect 5577 2860 6363 2894
rect 5577 2636 6363 2670
rect 193 2523 781 2557
rect 5017 2546 6253 2580
rect 7680 2473 8257 2507
rect 4777 2434 6363 2468
rect 4697 2272 6363 2306
rect 7680 2233 8257 2267
rect 5017 2160 6253 2194
rect 5577 2070 6363 2104
rect 5577 1846 6363 1880
rect 5017 1756 6253 1790
rect 7680 1683 8257 1717
rect 4617 1644 6363 1678
rect 4857 1482 6363 1516
rect 7680 1443 8257 1477
rect 4937 1370 6253 1404
rect 5577 1280 6363 1314
rect 5577 1056 6363 1090
rect 4937 966 6253 1000
rect 7680 893 8257 927
rect 4777 854 6363 888
rect 4697 692 6363 726
rect 7680 653 8257 687
rect 113 603 1537 637
rect 4937 580 6253 614
rect 5577 490 6363 524
rect 5577 266 6363 300
rect 33 153 1457 187
rect 4937 176 6253 210
rect 7680 103 8257 137
rect 4617 64 6363 98
<< metal1 >>
rect 19 0 47 9480
rect 99 0 127 9480
rect 179 0 207 9480
rect 259 0 287 9480
rect 339 0 367 9480
rect 419 0 447 9480
rect 499 0 527 9480
rect 579 0 607 9480
rect 4491 9334 4555 9386
rect 4491 8784 4555 8836
rect 4491 8544 4555 8596
rect 4491 7994 4555 8046
rect 4491 7754 4555 7806
rect 4491 7204 4555 7256
rect 4491 6964 4555 7016
rect 4491 6414 4555 6466
rect 4491 5384 4555 5436
rect 4491 4834 4555 4886
rect 4491 4594 4555 4646
rect 4491 4044 4555 4096
rect 4491 3804 4555 3856
rect 4491 3254 4555 3306
rect 4491 3014 4555 3066
rect 4491 2464 4555 2516
rect 4491 1434 4555 1486
rect 4491 884 4555 936
rect 4491 644 4555 696
rect 4603 198 4631 101148
rect 4683 592 4711 101148
rect 4763 988 4791 101148
rect 4843 1382 4871 101148
rect 4923 2568 4951 101148
rect 5003 2962 5031 101148
rect 5083 3358 5111 101148
rect 5163 3752 5191 101148
rect 5243 4148 5271 101148
rect 5323 4542 5351 101148
rect 5403 4938 5431 101148
rect 5483 5332 5511 101148
rect 5563 6518 5591 101148
rect 5643 6912 5671 101148
rect 5723 7308 5751 101148
rect 5803 7702 5831 101148
rect 5883 8098 5911 101148
rect 5963 8492 5991 101148
rect 6043 8888 6071 101148
rect 6123 9282 6151 101148
rect 6114 9085 6160 9282
rect 6034 8690 6080 8888
rect 5954 8295 6000 8492
rect 5874 7900 5920 8098
rect 5794 7505 5840 7702
rect 5714 7110 5760 7308
rect 5634 6715 5680 6912
rect 5554 6320 5600 6518
rect 5474 5135 5520 5332
rect 5394 4740 5440 4938
rect 5314 4345 5360 4542
rect 5234 3950 5280 4148
rect 5154 3555 5200 3752
rect 5074 3160 5120 3358
rect 4994 2765 5040 2962
rect 4914 2370 4960 2568
rect 4834 1185 4880 1382
rect 4754 790 4800 988
rect 4674 395 4720 592
rect 4491 94 4555 146
rect 4594 0 4640 198
rect 4683 0 4711 395
rect 4763 0 4791 790
rect 4843 0 4871 1185
rect 4923 0 4951 2370
rect 5003 0 5031 2765
rect 5083 0 5111 3160
rect 5163 0 5191 3555
rect 5243 0 5271 3950
rect 5323 0 5351 4345
rect 5403 0 5431 4740
rect 5483 0 5511 5135
rect 5563 0 5591 6320
rect 5643 0 5671 6715
rect 5723 0 5751 7110
rect 5803 0 5831 7505
rect 5883 0 5911 7900
rect 5963 0 5991 8295
rect 6043 0 6071 8690
rect 6123 0 6151 9085
rect 6451 -16 6497 101076
rect 6875 42 6923 101134
rect 7307 42 7355 101134
rect 7699 28 7727 101120
rect 8095 28 8123 101120
<< metal2 >>
rect 6446 100724 6502 100772
rect 6871 100724 6927 100772
rect 7303 100724 7359 100772
rect 7685 100701 7741 100749
rect 8081 100701 8137 100749
rect 6446 100350 6502 100398
rect 6871 100292 6927 100340
rect 7303 100292 7359 100340
rect 7685 100306 7741 100354
rect 8081 100306 8137 100354
rect 6446 99934 6502 99982
rect 6871 99934 6927 99982
rect 7303 99934 7359 99982
rect 7685 99911 7741 99959
rect 8081 99911 8137 99959
rect 6446 99560 6502 99608
rect 6871 99502 6927 99550
rect 7303 99502 7359 99550
rect 7685 99516 7741 99564
rect 8081 99516 8137 99564
rect 6446 99144 6502 99192
rect 6871 99144 6927 99192
rect 7303 99144 7359 99192
rect 7685 99121 7741 99169
rect 8081 99121 8137 99169
rect 6446 98770 6502 98818
rect 6871 98712 6927 98760
rect 7303 98712 7359 98760
rect 7685 98726 7741 98774
rect 8081 98726 8137 98774
rect 6446 98354 6502 98402
rect 6871 98354 6927 98402
rect 7303 98354 7359 98402
rect 7685 98331 7741 98379
rect 8081 98331 8137 98379
rect 6446 97980 6502 98028
rect 6871 97922 6927 97970
rect 7303 97922 7359 97970
rect 7685 97936 7741 97984
rect 8081 97936 8137 97984
rect 6446 97564 6502 97612
rect 6871 97564 6927 97612
rect 7303 97564 7359 97612
rect 7685 97541 7741 97589
rect 8081 97541 8137 97589
rect 6446 97190 6502 97238
rect 6871 97132 6927 97180
rect 7303 97132 7359 97180
rect 7685 97146 7741 97194
rect 8081 97146 8137 97194
rect 6446 96774 6502 96822
rect 6871 96774 6927 96822
rect 7303 96774 7359 96822
rect 7685 96751 7741 96799
rect 8081 96751 8137 96799
rect 6446 96400 6502 96448
rect 6871 96342 6927 96390
rect 7303 96342 7359 96390
rect 7685 96356 7741 96404
rect 8081 96356 8137 96404
rect 6446 95984 6502 96032
rect 6871 95984 6927 96032
rect 7303 95984 7359 96032
rect 7685 95961 7741 96009
rect 8081 95961 8137 96009
rect 6446 95610 6502 95658
rect 6871 95552 6927 95600
rect 7303 95552 7359 95600
rect 7685 95566 7741 95614
rect 8081 95566 8137 95614
rect 6446 95194 6502 95242
rect 6871 95194 6927 95242
rect 7303 95194 7359 95242
rect 7685 95171 7741 95219
rect 8081 95171 8137 95219
rect 6446 94820 6502 94868
rect 6871 94762 6927 94810
rect 7303 94762 7359 94810
rect 7685 94776 7741 94824
rect 8081 94776 8137 94824
rect 6446 94404 6502 94452
rect 6871 94404 6927 94452
rect 7303 94404 7359 94452
rect 7685 94381 7741 94429
rect 8081 94381 8137 94429
rect 6446 94030 6502 94078
rect 6871 93972 6927 94020
rect 7303 93972 7359 94020
rect 7685 93986 7741 94034
rect 8081 93986 8137 94034
rect 6446 93614 6502 93662
rect 6871 93614 6927 93662
rect 7303 93614 7359 93662
rect 7685 93591 7741 93639
rect 8081 93591 8137 93639
rect 6446 93240 6502 93288
rect 6871 93182 6927 93230
rect 7303 93182 7359 93230
rect 7685 93196 7741 93244
rect 8081 93196 8137 93244
rect 6446 92824 6502 92872
rect 6871 92824 6927 92872
rect 7303 92824 7359 92872
rect 7685 92801 7741 92849
rect 8081 92801 8137 92849
rect 6446 92450 6502 92498
rect 6871 92392 6927 92440
rect 7303 92392 7359 92440
rect 7685 92406 7741 92454
rect 8081 92406 8137 92454
rect 6446 92034 6502 92082
rect 6871 92034 6927 92082
rect 7303 92034 7359 92082
rect 7685 92011 7741 92059
rect 8081 92011 8137 92059
rect 6446 91660 6502 91708
rect 6871 91602 6927 91650
rect 7303 91602 7359 91650
rect 7685 91616 7741 91664
rect 8081 91616 8137 91664
rect 6446 91244 6502 91292
rect 6871 91244 6927 91292
rect 7303 91244 7359 91292
rect 7685 91221 7741 91269
rect 8081 91221 8137 91269
rect 6446 90870 6502 90918
rect 6871 90812 6927 90860
rect 7303 90812 7359 90860
rect 7685 90826 7741 90874
rect 8081 90826 8137 90874
rect 6446 90454 6502 90502
rect 6871 90454 6927 90502
rect 7303 90454 7359 90502
rect 7685 90431 7741 90479
rect 8081 90431 8137 90479
rect 6446 90080 6502 90128
rect 6871 90022 6927 90070
rect 7303 90022 7359 90070
rect 7685 90036 7741 90084
rect 8081 90036 8137 90084
rect 6446 89664 6502 89712
rect 6871 89664 6927 89712
rect 7303 89664 7359 89712
rect 7685 89641 7741 89689
rect 8081 89641 8137 89689
rect 6446 89290 6502 89338
rect 6871 89232 6927 89280
rect 7303 89232 7359 89280
rect 7685 89246 7741 89294
rect 8081 89246 8137 89294
rect 6446 88874 6502 88922
rect 6871 88874 6927 88922
rect 7303 88874 7359 88922
rect 7685 88851 7741 88899
rect 8081 88851 8137 88899
rect 6446 88500 6502 88548
rect 6871 88442 6927 88490
rect 7303 88442 7359 88490
rect 7685 88456 7741 88504
rect 8081 88456 8137 88504
rect 6446 88084 6502 88132
rect 6871 88084 6927 88132
rect 7303 88084 7359 88132
rect 7685 88061 7741 88109
rect 8081 88061 8137 88109
rect 6446 87710 6502 87758
rect 6871 87652 6927 87700
rect 7303 87652 7359 87700
rect 7685 87666 7741 87714
rect 8081 87666 8137 87714
rect 6446 87294 6502 87342
rect 6871 87294 6927 87342
rect 7303 87294 7359 87342
rect 7685 87271 7741 87319
rect 8081 87271 8137 87319
rect 6446 86920 6502 86968
rect 6871 86862 6927 86910
rect 7303 86862 7359 86910
rect 7685 86876 7741 86924
rect 8081 86876 8137 86924
rect 6446 86504 6502 86552
rect 6871 86504 6927 86552
rect 7303 86504 7359 86552
rect 7685 86481 7741 86529
rect 8081 86481 8137 86529
rect 6446 86130 6502 86178
rect 6871 86072 6927 86120
rect 7303 86072 7359 86120
rect 7685 86086 7741 86134
rect 8081 86086 8137 86134
rect 6446 85714 6502 85762
rect 6871 85714 6927 85762
rect 7303 85714 7359 85762
rect 7685 85691 7741 85739
rect 8081 85691 8137 85739
rect 6446 85340 6502 85388
rect 6871 85282 6927 85330
rect 7303 85282 7359 85330
rect 7685 85296 7741 85344
rect 8081 85296 8137 85344
rect 6446 84924 6502 84972
rect 6871 84924 6927 84972
rect 7303 84924 7359 84972
rect 7685 84901 7741 84949
rect 8081 84901 8137 84949
rect 6446 84550 6502 84598
rect 6871 84492 6927 84540
rect 7303 84492 7359 84540
rect 7685 84506 7741 84554
rect 8081 84506 8137 84554
rect 6446 84134 6502 84182
rect 6871 84134 6927 84182
rect 7303 84134 7359 84182
rect 7685 84111 7741 84159
rect 8081 84111 8137 84159
rect 6446 83760 6502 83808
rect 6871 83702 6927 83750
rect 7303 83702 7359 83750
rect 7685 83716 7741 83764
rect 8081 83716 8137 83764
rect 6446 83344 6502 83392
rect 6871 83344 6927 83392
rect 7303 83344 7359 83392
rect 7685 83321 7741 83369
rect 8081 83321 8137 83369
rect 6446 82970 6502 83018
rect 6871 82912 6927 82960
rect 7303 82912 7359 82960
rect 7685 82926 7741 82974
rect 8081 82926 8137 82974
rect 6446 82554 6502 82602
rect 6871 82554 6927 82602
rect 7303 82554 7359 82602
rect 7685 82531 7741 82579
rect 8081 82531 8137 82579
rect 6446 82180 6502 82228
rect 6871 82122 6927 82170
rect 7303 82122 7359 82170
rect 7685 82136 7741 82184
rect 8081 82136 8137 82184
rect 6446 81764 6502 81812
rect 6871 81764 6927 81812
rect 7303 81764 7359 81812
rect 7685 81741 7741 81789
rect 8081 81741 8137 81789
rect 6446 81390 6502 81438
rect 6871 81332 6927 81380
rect 7303 81332 7359 81380
rect 7685 81346 7741 81394
rect 8081 81346 8137 81394
rect 6446 80974 6502 81022
rect 6871 80974 6927 81022
rect 7303 80974 7359 81022
rect 7685 80951 7741 80999
rect 8081 80951 8137 80999
rect 6446 80600 6502 80648
rect 6871 80542 6927 80590
rect 7303 80542 7359 80590
rect 7685 80556 7741 80604
rect 8081 80556 8137 80604
rect 6446 80184 6502 80232
rect 6871 80184 6927 80232
rect 7303 80184 7359 80232
rect 7685 80161 7741 80209
rect 8081 80161 8137 80209
rect 6446 79810 6502 79858
rect 6871 79752 6927 79800
rect 7303 79752 7359 79800
rect 7685 79766 7741 79814
rect 8081 79766 8137 79814
rect 6446 79394 6502 79442
rect 6871 79394 6927 79442
rect 7303 79394 7359 79442
rect 7685 79371 7741 79419
rect 8081 79371 8137 79419
rect 6446 79020 6502 79068
rect 6871 78962 6927 79010
rect 7303 78962 7359 79010
rect 7685 78976 7741 79024
rect 8081 78976 8137 79024
rect 6446 78604 6502 78652
rect 6871 78604 6927 78652
rect 7303 78604 7359 78652
rect 7685 78581 7741 78629
rect 8081 78581 8137 78629
rect 6446 78230 6502 78278
rect 6871 78172 6927 78220
rect 7303 78172 7359 78220
rect 7685 78186 7741 78234
rect 8081 78186 8137 78234
rect 6446 77814 6502 77862
rect 6871 77814 6927 77862
rect 7303 77814 7359 77862
rect 7685 77791 7741 77839
rect 8081 77791 8137 77839
rect 6446 77440 6502 77488
rect 6871 77382 6927 77430
rect 7303 77382 7359 77430
rect 7685 77396 7741 77444
rect 8081 77396 8137 77444
rect 6446 77024 6502 77072
rect 6871 77024 6927 77072
rect 7303 77024 7359 77072
rect 7685 77001 7741 77049
rect 8081 77001 8137 77049
rect 6446 76650 6502 76698
rect 6871 76592 6927 76640
rect 7303 76592 7359 76640
rect 7685 76606 7741 76654
rect 8081 76606 8137 76654
rect 6446 76234 6502 76282
rect 6871 76234 6927 76282
rect 7303 76234 7359 76282
rect 7685 76211 7741 76259
rect 8081 76211 8137 76259
rect 6446 75860 6502 75908
rect 6871 75802 6927 75850
rect 7303 75802 7359 75850
rect 7685 75816 7741 75864
rect 8081 75816 8137 75864
rect 6446 75444 6502 75492
rect 6871 75444 6927 75492
rect 7303 75444 7359 75492
rect 7685 75421 7741 75469
rect 8081 75421 8137 75469
rect 6446 75070 6502 75118
rect 6871 75012 6927 75060
rect 7303 75012 7359 75060
rect 7685 75026 7741 75074
rect 8081 75026 8137 75074
rect 6446 74654 6502 74702
rect 6871 74654 6927 74702
rect 7303 74654 7359 74702
rect 7685 74631 7741 74679
rect 8081 74631 8137 74679
rect 6446 74280 6502 74328
rect 6871 74222 6927 74270
rect 7303 74222 7359 74270
rect 7685 74236 7741 74284
rect 8081 74236 8137 74284
rect 6446 73864 6502 73912
rect 6871 73864 6927 73912
rect 7303 73864 7359 73912
rect 7685 73841 7741 73889
rect 8081 73841 8137 73889
rect 6446 73490 6502 73538
rect 6871 73432 6927 73480
rect 7303 73432 7359 73480
rect 7685 73446 7741 73494
rect 8081 73446 8137 73494
rect 6446 73074 6502 73122
rect 6871 73074 6927 73122
rect 7303 73074 7359 73122
rect 7685 73051 7741 73099
rect 8081 73051 8137 73099
rect 6446 72700 6502 72748
rect 6871 72642 6927 72690
rect 7303 72642 7359 72690
rect 7685 72656 7741 72704
rect 8081 72656 8137 72704
rect 6446 72284 6502 72332
rect 6871 72284 6927 72332
rect 7303 72284 7359 72332
rect 7685 72261 7741 72309
rect 8081 72261 8137 72309
rect 6446 71910 6502 71958
rect 6871 71852 6927 71900
rect 7303 71852 7359 71900
rect 7685 71866 7741 71914
rect 8081 71866 8137 71914
rect 6446 71494 6502 71542
rect 6871 71494 6927 71542
rect 7303 71494 7359 71542
rect 7685 71471 7741 71519
rect 8081 71471 8137 71519
rect 6446 71120 6502 71168
rect 6871 71062 6927 71110
rect 7303 71062 7359 71110
rect 7685 71076 7741 71124
rect 8081 71076 8137 71124
rect 6446 70704 6502 70752
rect 6871 70704 6927 70752
rect 7303 70704 7359 70752
rect 7685 70681 7741 70729
rect 8081 70681 8137 70729
rect 6446 70330 6502 70378
rect 6871 70272 6927 70320
rect 7303 70272 7359 70320
rect 7685 70286 7741 70334
rect 8081 70286 8137 70334
rect 6446 69914 6502 69962
rect 6871 69914 6927 69962
rect 7303 69914 7359 69962
rect 7685 69891 7741 69939
rect 8081 69891 8137 69939
rect 6446 69540 6502 69588
rect 6871 69482 6927 69530
rect 7303 69482 7359 69530
rect 7685 69496 7741 69544
rect 8081 69496 8137 69544
rect 6446 69124 6502 69172
rect 6871 69124 6927 69172
rect 7303 69124 7359 69172
rect 7685 69101 7741 69149
rect 8081 69101 8137 69149
rect 6446 68750 6502 68798
rect 6871 68692 6927 68740
rect 7303 68692 7359 68740
rect 7685 68706 7741 68754
rect 8081 68706 8137 68754
rect 6446 68334 6502 68382
rect 6871 68334 6927 68382
rect 7303 68334 7359 68382
rect 7685 68311 7741 68359
rect 8081 68311 8137 68359
rect 6446 67960 6502 68008
rect 6871 67902 6927 67950
rect 7303 67902 7359 67950
rect 7685 67916 7741 67964
rect 8081 67916 8137 67964
rect 6446 67544 6502 67592
rect 6871 67544 6927 67592
rect 7303 67544 7359 67592
rect 7685 67521 7741 67569
rect 8081 67521 8137 67569
rect 6446 67170 6502 67218
rect 6871 67112 6927 67160
rect 7303 67112 7359 67160
rect 7685 67126 7741 67174
rect 8081 67126 8137 67174
rect 6446 66754 6502 66802
rect 6871 66754 6927 66802
rect 7303 66754 7359 66802
rect 7685 66731 7741 66779
rect 8081 66731 8137 66779
rect 6446 66380 6502 66428
rect 6871 66322 6927 66370
rect 7303 66322 7359 66370
rect 7685 66336 7741 66384
rect 8081 66336 8137 66384
rect 6446 65964 6502 66012
rect 6871 65964 6927 66012
rect 7303 65964 7359 66012
rect 7685 65941 7741 65989
rect 8081 65941 8137 65989
rect 6446 65590 6502 65638
rect 6871 65532 6927 65580
rect 7303 65532 7359 65580
rect 7685 65546 7741 65594
rect 8081 65546 8137 65594
rect 6446 65174 6502 65222
rect 6871 65174 6927 65222
rect 7303 65174 7359 65222
rect 7685 65151 7741 65199
rect 8081 65151 8137 65199
rect 6446 64800 6502 64848
rect 6871 64742 6927 64790
rect 7303 64742 7359 64790
rect 7685 64756 7741 64804
rect 8081 64756 8137 64804
rect 6446 64384 6502 64432
rect 6871 64384 6927 64432
rect 7303 64384 7359 64432
rect 7685 64361 7741 64409
rect 8081 64361 8137 64409
rect 6446 64010 6502 64058
rect 6871 63952 6927 64000
rect 7303 63952 7359 64000
rect 7685 63966 7741 64014
rect 8081 63966 8137 64014
rect 6446 63594 6502 63642
rect 6871 63594 6927 63642
rect 7303 63594 7359 63642
rect 7685 63571 7741 63619
rect 8081 63571 8137 63619
rect 6446 63220 6502 63268
rect 6871 63162 6927 63210
rect 7303 63162 7359 63210
rect 7685 63176 7741 63224
rect 8081 63176 8137 63224
rect 6446 62804 6502 62852
rect 6871 62804 6927 62852
rect 7303 62804 7359 62852
rect 7685 62781 7741 62829
rect 8081 62781 8137 62829
rect 6446 62430 6502 62478
rect 6871 62372 6927 62420
rect 7303 62372 7359 62420
rect 7685 62386 7741 62434
rect 8081 62386 8137 62434
rect 6446 62014 6502 62062
rect 6871 62014 6927 62062
rect 7303 62014 7359 62062
rect 7685 61991 7741 62039
rect 8081 61991 8137 62039
rect 6446 61640 6502 61688
rect 6871 61582 6927 61630
rect 7303 61582 7359 61630
rect 7685 61596 7741 61644
rect 8081 61596 8137 61644
rect 6446 61224 6502 61272
rect 6871 61224 6927 61272
rect 7303 61224 7359 61272
rect 7685 61201 7741 61249
rect 8081 61201 8137 61249
rect 6446 60850 6502 60898
rect 6871 60792 6927 60840
rect 7303 60792 7359 60840
rect 7685 60806 7741 60854
rect 8081 60806 8137 60854
rect 6446 60434 6502 60482
rect 6871 60434 6927 60482
rect 7303 60434 7359 60482
rect 7685 60411 7741 60459
rect 8081 60411 8137 60459
rect 6446 60060 6502 60108
rect 6871 60002 6927 60050
rect 7303 60002 7359 60050
rect 7685 60016 7741 60064
rect 8081 60016 8137 60064
rect 6446 59644 6502 59692
rect 6871 59644 6927 59692
rect 7303 59644 7359 59692
rect 7685 59621 7741 59669
rect 8081 59621 8137 59669
rect 6446 59270 6502 59318
rect 6871 59212 6927 59260
rect 7303 59212 7359 59260
rect 7685 59226 7741 59274
rect 8081 59226 8137 59274
rect 6446 58854 6502 58902
rect 6871 58854 6927 58902
rect 7303 58854 7359 58902
rect 7685 58831 7741 58879
rect 8081 58831 8137 58879
rect 6446 58480 6502 58528
rect 6871 58422 6927 58470
rect 7303 58422 7359 58470
rect 7685 58436 7741 58484
rect 8081 58436 8137 58484
rect 6446 58064 6502 58112
rect 6871 58064 6927 58112
rect 7303 58064 7359 58112
rect 7685 58041 7741 58089
rect 8081 58041 8137 58089
rect 6446 57690 6502 57738
rect 6871 57632 6927 57680
rect 7303 57632 7359 57680
rect 7685 57646 7741 57694
rect 8081 57646 8137 57694
rect 6446 57274 6502 57322
rect 6871 57274 6927 57322
rect 7303 57274 7359 57322
rect 7685 57251 7741 57299
rect 8081 57251 8137 57299
rect 6446 56900 6502 56948
rect 6871 56842 6927 56890
rect 7303 56842 7359 56890
rect 7685 56856 7741 56904
rect 8081 56856 8137 56904
rect 6446 56484 6502 56532
rect 6871 56484 6927 56532
rect 7303 56484 7359 56532
rect 7685 56461 7741 56509
rect 8081 56461 8137 56509
rect 6446 56110 6502 56158
rect 6871 56052 6927 56100
rect 7303 56052 7359 56100
rect 7685 56066 7741 56114
rect 8081 56066 8137 56114
rect 6446 55694 6502 55742
rect 6871 55694 6927 55742
rect 7303 55694 7359 55742
rect 7685 55671 7741 55719
rect 8081 55671 8137 55719
rect 6446 55320 6502 55368
rect 6871 55262 6927 55310
rect 7303 55262 7359 55310
rect 7685 55276 7741 55324
rect 8081 55276 8137 55324
rect 6446 54904 6502 54952
rect 6871 54904 6927 54952
rect 7303 54904 7359 54952
rect 7685 54881 7741 54929
rect 8081 54881 8137 54929
rect 6446 54530 6502 54578
rect 6871 54472 6927 54520
rect 7303 54472 7359 54520
rect 7685 54486 7741 54534
rect 8081 54486 8137 54534
rect 6446 54114 6502 54162
rect 6871 54114 6927 54162
rect 7303 54114 7359 54162
rect 7685 54091 7741 54139
rect 8081 54091 8137 54139
rect 6446 53740 6502 53788
rect 6871 53682 6927 53730
rect 7303 53682 7359 53730
rect 7685 53696 7741 53744
rect 8081 53696 8137 53744
rect 6446 53324 6502 53372
rect 6871 53324 6927 53372
rect 7303 53324 7359 53372
rect 7685 53301 7741 53349
rect 8081 53301 8137 53349
rect 6446 52950 6502 52998
rect 6871 52892 6927 52940
rect 7303 52892 7359 52940
rect 7685 52906 7741 52954
rect 8081 52906 8137 52954
rect 6446 52534 6502 52582
rect 6871 52534 6927 52582
rect 7303 52534 7359 52582
rect 7685 52511 7741 52559
rect 8081 52511 8137 52559
rect 6446 52160 6502 52208
rect 6871 52102 6927 52150
rect 7303 52102 7359 52150
rect 7685 52116 7741 52164
rect 8081 52116 8137 52164
rect 6446 51744 6502 51792
rect 6871 51744 6927 51792
rect 7303 51744 7359 51792
rect 7685 51721 7741 51769
rect 8081 51721 8137 51769
rect 6446 51370 6502 51418
rect 6871 51312 6927 51360
rect 7303 51312 7359 51360
rect 7685 51326 7741 51374
rect 8081 51326 8137 51374
rect 6446 50954 6502 51002
rect 6871 50954 6927 51002
rect 7303 50954 7359 51002
rect 7685 50931 7741 50979
rect 8081 50931 8137 50979
rect 6446 50580 6502 50628
rect 6871 50522 6927 50570
rect 7303 50522 7359 50570
rect 7685 50536 7741 50584
rect 8081 50536 8137 50584
rect 6446 50164 6502 50212
rect 6871 50164 6927 50212
rect 7303 50164 7359 50212
rect 7685 50141 7741 50189
rect 8081 50141 8137 50189
rect 6446 49790 6502 49838
rect 6871 49732 6927 49780
rect 7303 49732 7359 49780
rect 7685 49746 7741 49794
rect 8081 49746 8137 49794
rect 6446 49374 6502 49422
rect 6871 49374 6927 49422
rect 7303 49374 7359 49422
rect 7685 49351 7741 49399
rect 8081 49351 8137 49399
rect 6446 49000 6502 49048
rect 6871 48942 6927 48990
rect 7303 48942 7359 48990
rect 7685 48956 7741 49004
rect 8081 48956 8137 49004
rect 6446 48584 6502 48632
rect 6871 48584 6927 48632
rect 7303 48584 7359 48632
rect 7685 48561 7741 48609
rect 8081 48561 8137 48609
rect 6446 48210 6502 48258
rect 6871 48152 6927 48200
rect 7303 48152 7359 48200
rect 7685 48166 7741 48214
rect 8081 48166 8137 48214
rect 6446 47794 6502 47842
rect 6871 47794 6927 47842
rect 7303 47794 7359 47842
rect 7685 47771 7741 47819
rect 8081 47771 8137 47819
rect 6446 47420 6502 47468
rect 6871 47362 6927 47410
rect 7303 47362 7359 47410
rect 7685 47376 7741 47424
rect 8081 47376 8137 47424
rect 6446 47004 6502 47052
rect 6871 47004 6927 47052
rect 7303 47004 7359 47052
rect 7685 46981 7741 47029
rect 8081 46981 8137 47029
rect 6446 46630 6502 46678
rect 6871 46572 6927 46620
rect 7303 46572 7359 46620
rect 7685 46586 7741 46634
rect 8081 46586 8137 46634
rect 6446 46214 6502 46262
rect 6871 46214 6927 46262
rect 7303 46214 7359 46262
rect 7685 46191 7741 46239
rect 8081 46191 8137 46239
rect 6446 45840 6502 45888
rect 6871 45782 6927 45830
rect 7303 45782 7359 45830
rect 7685 45796 7741 45844
rect 8081 45796 8137 45844
rect 6446 45424 6502 45472
rect 6871 45424 6927 45472
rect 7303 45424 7359 45472
rect 7685 45401 7741 45449
rect 8081 45401 8137 45449
rect 6446 45050 6502 45098
rect 6871 44992 6927 45040
rect 7303 44992 7359 45040
rect 7685 45006 7741 45054
rect 8081 45006 8137 45054
rect 6446 44634 6502 44682
rect 6871 44634 6927 44682
rect 7303 44634 7359 44682
rect 7685 44611 7741 44659
rect 8081 44611 8137 44659
rect 6446 44260 6502 44308
rect 6871 44202 6927 44250
rect 7303 44202 7359 44250
rect 7685 44216 7741 44264
rect 8081 44216 8137 44264
rect 6446 43844 6502 43892
rect 6871 43844 6927 43892
rect 7303 43844 7359 43892
rect 7685 43821 7741 43869
rect 8081 43821 8137 43869
rect 6446 43470 6502 43518
rect 6871 43412 6927 43460
rect 7303 43412 7359 43460
rect 7685 43426 7741 43474
rect 8081 43426 8137 43474
rect 6446 43054 6502 43102
rect 6871 43054 6927 43102
rect 7303 43054 7359 43102
rect 7685 43031 7741 43079
rect 8081 43031 8137 43079
rect 6446 42680 6502 42728
rect 6871 42622 6927 42670
rect 7303 42622 7359 42670
rect 7685 42636 7741 42684
rect 8081 42636 8137 42684
rect 6446 42264 6502 42312
rect 6871 42264 6927 42312
rect 7303 42264 7359 42312
rect 7685 42241 7741 42289
rect 8081 42241 8137 42289
rect 6446 41890 6502 41938
rect 6871 41832 6927 41880
rect 7303 41832 7359 41880
rect 7685 41846 7741 41894
rect 8081 41846 8137 41894
rect 6446 41474 6502 41522
rect 6871 41474 6927 41522
rect 7303 41474 7359 41522
rect 7685 41451 7741 41499
rect 8081 41451 8137 41499
rect 6446 41100 6502 41148
rect 6871 41042 6927 41090
rect 7303 41042 7359 41090
rect 7685 41056 7741 41104
rect 8081 41056 8137 41104
rect 6446 40684 6502 40732
rect 6871 40684 6927 40732
rect 7303 40684 7359 40732
rect 7685 40661 7741 40709
rect 8081 40661 8137 40709
rect 6446 40310 6502 40358
rect 6871 40252 6927 40300
rect 7303 40252 7359 40300
rect 7685 40266 7741 40314
rect 8081 40266 8137 40314
rect 6446 39894 6502 39942
rect 6871 39894 6927 39942
rect 7303 39894 7359 39942
rect 7685 39871 7741 39919
rect 8081 39871 8137 39919
rect 6446 39520 6502 39568
rect 6871 39462 6927 39510
rect 7303 39462 7359 39510
rect 7685 39476 7741 39524
rect 8081 39476 8137 39524
rect 6446 39104 6502 39152
rect 6871 39104 6927 39152
rect 7303 39104 7359 39152
rect 7685 39081 7741 39129
rect 8081 39081 8137 39129
rect 6446 38730 6502 38778
rect 6871 38672 6927 38720
rect 7303 38672 7359 38720
rect 7685 38686 7741 38734
rect 8081 38686 8137 38734
rect 6446 38314 6502 38362
rect 6871 38314 6927 38362
rect 7303 38314 7359 38362
rect 7685 38291 7741 38339
rect 8081 38291 8137 38339
rect 6446 37940 6502 37988
rect 6871 37882 6927 37930
rect 7303 37882 7359 37930
rect 7685 37896 7741 37944
rect 8081 37896 8137 37944
rect 6446 37524 6502 37572
rect 6871 37524 6927 37572
rect 7303 37524 7359 37572
rect 7685 37501 7741 37549
rect 8081 37501 8137 37549
rect 6446 37150 6502 37198
rect 6871 37092 6927 37140
rect 7303 37092 7359 37140
rect 7685 37106 7741 37154
rect 8081 37106 8137 37154
rect 6446 36734 6502 36782
rect 6871 36734 6927 36782
rect 7303 36734 7359 36782
rect 7685 36711 7741 36759
rect 8081 36711 8137 36759
rect 6446 36360 6502 36408
rect 6871 36302 6927 36350
rect 7303 36302 7359 36350
rect 7685 36316 7741 36364
rect 8081 36316 8137 36364
rect 6446 35944 6502 35992
rect 6871 35944 6927 35992
rect 7303 35944 7359 35992
rect 7685 35921 7741 35969
rect 8081 35921 8137 35969
rect 6446 35570 6502 35618
rect 6871 35512 6927 35560
rect 7303 35512 7359 35560
rect 7685 35526 7741 35574
rect 8081 35526 8137 35574
rect 6446 35154 6502 35202
rect 6871 35154 6927 35202
rect 7303 35154 7359 35202
rect 7685 35131 7741 35179
rect 8081 35131 8137 35179
rect 6446 34780 6502 34828
rect 6871 34722 6927 34770
rect 7303 34722 7359 34770
rect 7685 34736 7741 34784
rect 8081 34736 8137 34784
rect 6446 34364 6502 34412
rect 6871 34364 6927 34412
rect 7303 34364 7359 34412
rect 7685 34341 7741 34389
rect 8081 34341 8137 34389
rect 6446 33990 6502 34038
rect 6871 33932 6927 33980
rect 7303 33932 7359 33980
rect 7685 33946 7741 33994
rect 8081 33946 8137 33994
rect 6446 33574 6502 33622
rect 6871 33574 6927 33622
rect 7303 33574 7359 33622
rect 7685 33551 7741 33599
rect 8081 33551 8137 33599
rect 6446 33200 6502 33248
rect 6871 33142 6927 33190
rect 7303 33142 7359 33190
rect 7685 33156 7741 33204
rect 8081 33156 8137 33204
rect 6446 32784 6502 32832
rect 6871 32784 6927 32832
rect 7303 32784 7359 32832
rect 7685 32761 7741 32809
rect 8081 32761 8137 32809
rect 6446 32410 6502 32458
rect 6871 32352 6927 32400
rect 7303 32352 7359 32400
rect 7685 32366 7741 32414
rect 8081 32366 8137 32414
rect 6446 31994 6502 32042
rect 6871 31994 6927 32042
rect 7303 31994 7359 32042
rect 7685 31971 7741 32019
rect 8081 31971 8137 32019
rect 6446 31620 6502 31668
rect 6871 31562 6927 31610
rect 7303 31562 7359 31610
rect 7685 31576 7741 31624
rect 8081 31576 8137 31624
rect 6446 31204 6502 31252
rect 6871 31204 6927 31252
rect 7303 31204 7359 31252
rect 7685 31181 7741 31229
rect 8081 31181 8137 31229
rect 6446 30830 6502 30878
rect 6871 30772 6927 30820
rect 7303 30772 7359 30820
rect 7685 30786 7741 30834
rect 8081 30786 8137 30834
rect 6446 30414 6502 30462
rect 6871 30414 6927 30462
rect 7303 30414 7359 30462
rect 7685 30391 7741 30439
rect 8081 30391 8137 30439
rect 6446 30040 6502 30088
rect 6871 29982 6927 30030
rect 7303 29982 7359 30030
rect 7685 29996 7741 30044
rect 8081 29996 8137 30044
rect 6446 29624 6502 29672
rect 6871 29624 6927 29672
rect 7303 29624 7359 29672
rect 7685 29601 7741 29649
rect 8081 29601 8137 29649
rect 6446 29250 6502 29298
rect 6871 29192 6927 29240
rect 7303 29192 7359 29240
rect 7685 29206 7741 29254
rect 8081 29206 8137 29254
rect 6446 28834 6502 28882
rect 6871 28834 6927 28882
rect 7303 28834 7359 28882
rect 7685 28811 7741 28859
rect 8081 28811 8137 28859
rect 6446 28460 6502 28508
rect 6871 28402 6927 28450
rect 7303 28402 7359 28450
rect 7685 28416 7741 28464
rect 8081 28416 8137 28464
rect 6446 28044 6502 28092
rect 6871 28044 6927 28092
rect 7303 28044 7359 28092
rect 7685 28021 7741 28069
rect 8081 28021 8137 28069
rect 6446 27670 6502 27718
rect 6871 27612 6927 27660
rect 7303 27612 7359 27660
rect 7685 27626 7741 27674
rect 8081 27626 8137 27674
rect 6446 27254 6502 27302
rect 6871 27254 6927 27302
rect 7303 27254 7359 27302
rect 7685 27231 7741 27279
rect 8081 27231 8137 27279
rect 6446 26880 6502 26928
rect 6871 26822 6927 26870
rect 7303 26822 7359 26870
rect 7685 26836 7741 26884
rect 8081 26836 8137 26884
rect 6446 26464 6502 26512
rect 6871 26464 6927 26512
rect 7303 26464 7359 26512
rect 7685 26441 7741 26489
rect 8081 26441 8137 26489
rect 6446 26090 6502 26138
rect 6871 26032 6927 26080
rect 7303 26032 7359 26080
rect 7685 26046 7741 26094
rect 8081 26046 8137 26094
rect 6446 25674 6502 25722
rect 6871 25674 6927 25722
rect 7303 25674 7359 25722
rect 7685 25651 7741 25699
rect 8081 25651 8137 25699
rect 6446 25300 6502 25348
rect 6871 25242 6927 25290
rect 7303 25242 7359 25290
rect 7685 25256 7741 25304
rect 8081 25256 8137 25304
rect 6446 24884 6502 24932
rect 6871 24884 6927 24932
rect 7303 24884 7359 24932
rect 7685 24861 7741 24909
rect 8081 24861 8137 24909
rect 6446 24510 6502 24558
rect 6871 24452 6927 24500
rect 7303 24452 7359 24500
rect 7685 24466 7741 24514
rect 8081 24466 8137 24514
rect 6446 24094 6502 24142
rect 6871 24094 6927 24142
rect 7303 24094 7359 24142
rect 7685 24071 7741 24119
rect 8081 24071 8137 24119
rect 6446 23720 6502 23768
rect 6871 23662 6927 23710
rect 7303 23662 7359 23710
rect 7685 23676 7741 23724
rect 8081 23676 8137 23724
rect 6446 23304 6502 23352
rect 6871 23304 6927 23352
rect 7303 23304 7359 23352
rect 7685 23281 7741 23329
rect 8081 23281 8137 23329
rect 6446 22930 6502 22978
rect 6871 22872 6927 22920
rect 7303 22872 7359 22920
rect 7685 22886 7741 22934
rect 8081 22886 8137 22934
rect 6446 22514 6502 22562
rect 6871 22514 6927 22562
rect 7303 22514 7359 22562
rect 7685 22491 7741 22539
rect 8081 22491 8137 22539
rect 6446 22140 6502 22188
rect 6871 22082 6927 22130
rect 7303 22082 7359 22130
rect 7685 22096 7741 22144
rect 8081 22096 8137 22144
rect 6446 21724 6502 21772
rect 6871 21724 6927 21772
rect 7303 21724 7359 21772
rect 7685 21701 7741 21749
rect 8081 21701 8137 21749
rect 6446 21350 6502 21398
rect 6871 21292 6927 21340
rect 7303 21292 7359 21340
rect 7685 21306 7741 21354
rect 8081 21306 8137 21354
rect 6446 20934 6502 20982
rect 6871 20934 6927 20982
rect 7303 20934 7359 20982
rect 7685 20911 7741 20959
rect 8081 20911 8137 20959
rect 6446 20560 6502 20608
rect 6871 20502 6927 20550
rect 7303 20502 7359 20550
rect 7685 20516 7741 20564
rect 8081 20516 8137 20564
rect 6446 20144 6502 20192
rect 6871 20144 6927 20192
rect 7303 20144 7359 20192
rect 7685 20121 7741 20169
rect 8081 20121 8137 20169
rect 6446 19770 6502 19818
rect 6871 19712 6927 19760
rect 7303 19712 7359 19760
rect 7685 19726 7741 19774
rect 8081 19726 8137 19774
rect 6446 19354 6502 19402
rect 6871 19354 6927 19402
rect 7303 19354 7359 19402
rect 7685 19331 7741 19379
rect 8081 19331 8137 19379
rect 6446 18980 6502 19028
rect 6871 18922 6927 18970
rect 7303 18922 7359 18970
rect 7685 18936 7741 18984
rect 8081 18936 8137 18984
rect 6446 18564 6502 18612
rect 6871 18564 6927 18612
rect 7303 18564 7359 18612
rect 7685 18541 7741 18589
rect 8081 18541 8137 18589
rect 6446 18190 6502 18238
rect 6871 18132 6927 18180
rect 7303 18132 7359 18180
rect 7685 18146 7741 18194
rect 8081 18146 8137 18194
rect 6446 17774 6502 17822
rect 6871 17774 6927 17822
rect 7303 17774 7359 17822
rect 7685 17751 7741 17799
rect 8081 17751 8137 17799
rect 6446 17400 6502 17448
rect 6871 17342 6927 17390
rect 7303 17342 7359 17390
rect 7685 17356 7741 17404
rect 8081 17356 8137 17404
rect 6446 16984 6502 17032
rect 6871 16984 6927 17032
rect 7303 16984 7359 17032
rect 7685 16961 7741 17009
rect 8081 16961 8137 17009
rect 6446 16610 6502 16658
rect 6871 16552 6927 16600
rect 7303 16552 7359 16600
rect 7685 16566 7741 16614
rect 8081 16566 8137 16614
rect 6446 16194 6502 16242
rect 6871 16194 6927 16242
rect 7303 16194 7359 16242
rect 7685 16171 7741 16219
rect 8081 16171 8137 16219
rect 6446 15820 6502 15868
rect 6871 15762 6927 15810
rect 7303 15762 7359 15810
rect 7685 15776 7741 15824
rect 8081 15776 8137 15824
rect 6446 15404 6502 15452
rect 6871 15404 6927 15452
rect 7303 15404 7359 15452
rect 7685 15381 7741 15429
rect 8081 15381 8137 15429
rect 6446 15030 6502 15078
rect 6871 14972 6927 15020
rect 7303 14972 7359 15020
rect 7685 14986 7741 15034
rect 8081 14986 8137 15034
rect 6446 14614 6502 14662
rect 6871 14614 6927 14662
rect 7303 14614 7359 14662
rect 7685 14591 7741 14639
rect 8081 14591 8137 14639
rect 6446 14240 6502 14288
rect 6871 14182 6927 14230
rect 7303 14182 7359 14230
rect 7685 14196 7741 14244
rect 8081 14196 8137 14244
rect 6446 13824 6502 13872
rect 6871 13824 6927 13872
rect 7303 13824 7359 13872
rect 7685 13801 7741 13849
rect 8081 13801 8137 13849
rect 6446 13450 6502 13498
rect 6871 13392 6927 13440
rect 7303 13392 7359 13440
rect 7685 13406 7741 13454
rect 8081 13406 8137 13454
rect 6446 13034 6502 13082
rect 6871 13034 6927 13082
rect 7303 13034 7359 13082
rect 7685 13011 7741 13059
rect 8081 13011 8137 13059
rect 6446 12660 6502 12708
rect 6871 12602 6927 12650
rect 7303 12602 7359 12650
rect 7685 12616 7741 12664
rect 8081 12616 8137 12664
rect 6446 12244 6502 12292
rect 6871 12244 6927 12292
rect 7303 12244 7359 12292
rect 7685 12221 7741 12269
rect 8081 12221 8137 12269
rect 6446 11870 6502 11918
rect 6871 11812 6927 11860
rect 7303 11812 7359 11860
rect 7685 11826 7741 11874
rect 8081 11826 8137 11874
rect 6446 11454 6502 11502
rect 6871 11454 6927 11502
rect 7303 11454 7359 11502
rect 7685 11431 7741 11479
rect 8081 11431 8137 11479
rect 6446 11080 6502 11128
rect 6871 11022 6927 11070
rect 7303 11022 7359 11070
rect 7685 11036 7741 11084
rect 8081 11036 8137 11084
rect 6446 10664 6502 10712
rect 6871 10664 6927 10712
rect 7303 10664 7359 10712
rect 7685 10641 7741 10689
rect 8081 10641 8137 10689
rect 6446 10290 6502 10338
rect 6871 10232 6927 10280
rect 7303 10232 7359 10280
rect 7685 10246 7741 10294
rect 8081 10246 8137 10294
rect 6446 9874 6502 9922
rect 6871 9874 6927 9922
rect 7303 9874 7359 9922
rect 7685 9851 7741 9899
rect 8081 9851 8137 9899
rect 6446 9500 6502 9548
rect 6871 9442 6927 9490
rect 7303 9442 7359 9490
rect 7685 9456 7741 9504
rect 8081 9456 8137 9504
rect 4523 9346 4621 9374
rect 4593 9099 4621 9346
rect 4593 9071 6137 9099
rect 6446 9084 6502 9132
rect 6871 9084 6927 9132
rect 7303 9084 7359 9132
rect 7685 9061 7741 9109
rect 8081 9061 8137 9109
rect 4523 8796 4621 8824
rect 4593 8704 4621 8796
rect 6446 8710 6502 8758
rect 4593 8676 6057 8704
rect 6871 8652 6927 8700
rect 7303 8652 7359 8700
rect 7685 8666 7741 8714
rect 8081 8666 8137 8714
rect 4523 8556 4621 8584
rect 4593 8309 4621 8556
rect 4593 8281 5977 8309
rect 6446 8294 6502 8342
rect 6871 8294 6927 8342
rect 7303 8294 7359 8342
rect 7685 8271 7741 8319
rect 8081 8271 8137 8319
rect 4523 8006 4621 8034
rect 4593 7914 4621 8006
rect 6446 7920 6502 7968
rect 4593 7886 5897 7914
rect 6871 7862 6927 7910
rect 7303 7862 7359 7910
rect 7685 7876 7741 7924
rect 8081 7876 8137 7924
rect 4523 7766 4621 7794
rect 4593 7519 4621 7766
rect 4593 7491 5817 7519
rect 6446 7504 6502 7552
rect 6871 7504 6927 7552
rect 7303 7504 7359 7552
rect 7685 7481 7741 7529
rect 8081 7481 8137 7529
rect 4523 7216 4621 7244
rect 4593 7124 4621 7216
rect 6446 7130 6502 7178
rect 4593 7096 5737 7124
rect 6871 7072 6927 7120
rect 7303 7072 7359 7120
rect 7685 7086 7741 7134
rect 8081 7086 8137 7134
rect 4523 6976 4621 7004
rect 4593 6729 4621 6976
rect 4593 6701 5657 6729
rect 6446 6714 6502 6762
rect 6871 6714 6927 6762
rect 7303 6714 7359 6762
rect 7685 6691 7741 6739
rect 8081 6691 8137 6739
rect 4523 6426 4621 6454
rect 4593 6334 4621 6426
rect 6446 6340 6502 6388
rect 4593 6306 5577 6334
rect 6871 6282 6927 6330
rect 7303 6282 7359 6330
rect 7685 6296 7741 6344
rect 8081 6296 8137 6344
rect 6446 5924 6502 5972
rect 6871 5924 6927 5972
rect 7303 5924 7359 5972
rect 7685 5901 7741 5949
rect 8081 5901 8137 5949
rect 6446 5550 6502 5598
rect 6871 5492 6927 5540
rect 7303 5492 7359 5540
rect 7685 5506 7741 5554
rect 8081 5506 8137 5554
rect 4523 5396 4621 5424
rect 4593 5149 4621 5396
rect 4593 5121 5497 5149
rect 6446 5134 6502 5182
rect 6871 5134 6927 5182
rect 7303 5134 7359 5182
rect 7685 5111 7741 5159
rect 8081 5111 8137 5159
rect 4523 4846 4621 4874
rect 4593 4754 4621 4846
rect 6446 4760 6502 4808
rect 4593 4726 5417 4754
rect 6871 4702 6927 4750
rect 7303 4702 7359 4750
rect 7685 4716 7741 4764
rect 8081 4716 8137 4764
rect 4523 4606 4621 4634
rect 4593 4359 4621 4606
rect 4593 4331 5337 4359
rect 6446 4344 6502 4392
rect 6871 4344 6927 4392
rect 7303 4344 7359 4392
rect 7685 4321 7741 4369
rect 8081 4321 8137 4369
rect 4523 4056 4621 4084
rect 4593 3964 4621 4056
rect 6446 3970 6502 4018
rect 4593 3936 5257 3964
rect 6871 3912 6927 3960
rect 7303 3912 7359 3960
rect 7685 3926 7741 3974
rect 8081 3926 8137 3974
rect 4523 3816 4621 3844
rect 4593 3569 4621 3816
rect 4593 3541 5177 3569
rect 6446 3554 6502 3602
rect 6871 3554 6927 3602
rect 7303 3554 7359 3602
rect 7685 3531 7741 3579
rect 8081 3531 8137 3579
rect 4523 3266 4621 3294
rect 4593 3174 4621 3266
rect 6446 3180 6502 3228
rect 4593 3146 5097 3174
rect 6871 3122 6927 3170
rect 7303 3122 7359 3170
rect 7685 3136 7741 3184
rect 8081 3136 8137 3184
rect 4523 3026 4621 3054
rect 4593 2779 4621 3026
rect 4593 2751 5017 2779
rect 6446 2764 6502 2812
rect 6871 2764 6927 2812
rect 7303 2764 7359 2812
rect 7685 2741 7741 2789
rect 8081 2741 8137 2789
rect 4523 2476 4621 2504
rect 4593 2384 4621 2476
rect 6446 2390 6502 2438
rect 4593 2356 4937 2384
rect 6871 2332 6927 2380
rect 7303 2332 7359 2380
rect 7685 2346 7741 2394
rect 8081 2346 8137 2394
rect 6446 1974 6502 2022
rect 6871 1974 6927 2022
rect 7303 1974 7359 2022
rect 7685 1951 7741 1999
rect 8081 1951 8137 1999
rect 6446 1600 6502 1648
rect 6871 1542 6927 1590
rect 7303 1542 7359 1590
rect 7685 1556 7741 1604
rect 8081 1556 8137 1604
rect 4523 1446 4621 1474
rect 4593 1199 4621 1446
rect 4593 1171 4857 1199
rect 6446 1184 6502 1232
rect 6871 1184 6927 1232
rect 7303 1184 7359 1232
rect 7685 1161 7741 1209
rect 8081 1161 8137 1209
rect 4523 896 4621 924
rect 4593 804 4621 896
rect 6446 810 6502 858
rect 4593 776 4777 804
rect 6871 752 6927 800
rect 7303 752 7359 800
rect 7685 766 7741 814
rect 8081 766 8137 814
rect 4523 656 4621 684
rect 4593 409 4621 656
rect 4593 381 4697 409
rect 6446 394 6502 442
rect 6871 394 6927 442
rect 7303 394 7359 442
rect 7685 371 7741 419
rect 8081 371 8137 419
rect 4523 106 4621 134
rect 4593 -14 4621 106
<< metal3 >>
rect 6425 100699 6523 100797
rect 6850 100699 6948 100797
rect 7282 100699 7380 100797
rect 7664 100676 7762 100774
rect 8060 100676 8158 100774
rect 6425 100325 6523 100423
rect 6850 100267 6948 100365
rect 7282 100267 7380 100365
rect 7664 100281 7762 100379
rect 8060 100281 8158 100379
rect 6425 99909 6523 100007
rect 6850 99909 6948 100007
rect 7282 99909 7380 100007
rect 7664 99886 7762 99984
rect 8060 99886 8158 99984
rect 6425 99535 6523 99633
rect 6850 99477 6948 99575
rect 7282 99477 7380 99575
rect 7664 99491 7762 99589
rect 8060 99491 8158 99589
rect 6425 99119 6523 99217
rect 6850 99119 6948 99217
rect 7282 99119 7380 99217
rect 7664 99096 7762 99194
rect 8060 99096 8158 99194
rect 6425 98745 6523 98843
rect 6850 98687 6948 98785
rect 7282 98687 7380 98785
rect 7664 98701 7762 98799
rect 8060 98701 8158 98799
rect 6425 98329 6523 98427
rect 6850 98329 6948 98427
rect 7282 98329 7380 98427
rect 7664 98306 7762 98404
rect 8060 98306 8158 98404
rect 6425 97955 6523 98053
rect 6850 97897 6948 97995
rect 7282 97897 7380 97995
rect 7664 97911 7762 98009
rect 8060 97911 8158 98009
rect 6425 97539 6523 97637
rect 6850 97539 6948 97637
rect 7282 97539 7380 97637
rect 7664 97516 7762 97614
rect 8060 97516 8158 97614
rect 6425 97165 6523 97263
rect 6850 97107 6948 97205
rect 7282 97107 7380 97205
rect 7664 97121 7762 97219
rect 8060 97121 8158 97219
rect 6425 96749 6523 96847
rect 6850 96749 6948 96847
rect 7282 96749 7380 96847
rect 7664 96726 7762 96824
rect 8060 96726 8158 96824
rect 6425 96375 6523 96473
rect 6850 96317 6948 96415
rect 7282 96317 7380 96415
rect 7664 96331 7762 96429
rect 8060 96331 8158 96429
rect 6425 95959 6523 96057
rect 6850 95959 6948 96057
rect 7282 95959 7380 96057
rect 7664 95936 7762 96034
rect 8060 95936 8158 96034
rect 6425 95585 6523 95683
rect 6850 95527 6948 95625
rect 7282 95527 7380 95625
rect 7664 95541 7762 95639
rect 8060 95541 8158 95639
rect 6425 95169 6523 95267
rect 6850 95169 6948 95267
rect 7282 95169 7380 95267
rect 7664 95146 7762 95244
rect 8060 95146 8158 95244
rect 6425 94795 6523 94893
rect 6850 94737 6948 94835
rect 7282 94737 7380 94835
rect 7664 94751 7762 94849
rect 8060 94751 8158 94849
rect 6425 94379 6523 94477
rect 6850 94379 6948 94477
rect 7282 94379 7380 94477
rect 7664 94356 7762 94454
rect 8060 94356 8158 94454
rect 6425 94005 6523 94103
rect 6850 93947 6948 94045
rect 7282 93947 7380 94045
rect 7664 93961 7762 94059
rect 8060 93961 8158 94059
rect 6425 93589 6523 93687
rect 6850 93589 6948 93687
rect 7282 93589 7380 93687
rect 7664 93566 7762 93664
rect 8060 93566 8158 93664
rect 6425 93215 6523 93313
rect 6850 93157 6948 93255
rect 7282 93157 7380 93255
rect 7664 93171 7762 93269
rect 8060 93171 8158 93269
rect 6425 92799 6523 92897
rect 6850 92799 6948 92897
rect 7282 92799 7380 92897
rect 7664 92776 7762 92874
rect 8060 92776 8158 92874
rect 6425 92425 6523 92523
rect 6850 92367 6948 92465
rect 7282 92367 7380 92465
rect 7664 92381 7762 92479
rect 8060 92381 8158 92479
rect 6425 92009 6523 92107
rect 6850 92009 6948 92107
rect 7282 92009 7380 92107
rect 7664 91986 7762 92084
rect 8060 91986 8158 92084
rect 6425 91635 6523 91733
rect 6850 91577 6948 91675
rect 7282 91577 7380 91675
rect 7664 91591 7762 91689
rect 8060 91591 8158 91689
rect 6425 91219 6523 91317
rect 6850 91219 6948 91317
rect 7282 91219 7380 91317
rect 7664 91196 7762 91294
rect 8060 91196 8158 91294
rect 6425 90845 6523 90943
rect 6850 90787 6948 90885
rect 7282 90787 7380 90885
rect 7664 90801 7762 90899
rect 8060 90801 8158 90899
rect 6425 90429 6523 90527
rect 6850 90429 6948 90527
rect 7282 90429 7380 90527
rect 7664 90406 7762 90504
rect 8060 90406 8158 90504
rect 6425 90055 6523 90153
rect 6850 89997 6948 90095
rect 7282 89997 7380 90095
rect 7664 90011 7762 90109
rect 8060 90011 8158 90109
rect 6425 89639 6523 89737
rect 6850 89639 6948 89737
rect 7282 89639 7380 89737
rect 7664 89616 7762 89714
rect 8060 89616 8158 89714
rect 6425 89265 6523 89363
rect 6850 89207 6948 89305
rect 7282 89207 7380 89305
rect 7664 89221 7762 89319
rect 8060 89221 8158 89319
rect 6425 88849 6523 88947
rect 6850 88849 6948 88947
rect 7282 88849 7380 88947
rect 7664 88826 7762 88924
rect 8060 88826 8158 88924
rect 6425 88475 6523 88573
rect 6850 88417 6948 88515
rect 7282 88417 7380 88515
rect 7664 88431 7762 88529
rect 8060 88431 8158 88529
rect 6425 88059 6523 88157
rect 6850 88059 6948 88157
rect 7282 88059 7380 88157
rect 7664 88036 7762 88134
rect 8060 88036 8158 88134
rect 6425 87685 6523 87783
rect 6850 87627 6948 87725
rect 7282 87627 7380 87725
rect 7664 87641 7762 87739
rect 8060 87641 8158 87739
rect 6425 87269 6523 87367
rect 6850 87269 6948 87367
rect 7282 87269 7380 87367
rect 7664 87246 7762 87344
rect 8060 87246 8158 87344
rect 6425 86895 6523 86993
rect 6850 86837 6948 86935
rect 7282 86837 7380 86935
rect 7664 86851 7762 86949
rect 8060 86851 8158 86949
rect 6425 86479 6523 86577
rect 6850 86479 6948 86577
rect 7282 86479 7380 86577
rect 7664 86456 7762 86554
rect 8060 86456 8158 86554
rect 6425 86105 6523 86203
rect 6850 86047 6948 86145
rect 7282 86047 7380 86145
rect 7664 86061 7762 86159
rect 8060 86061 8158 86159
rect 6425 85689 6523 85787
rect 6850 85689 6948 85787
rect 7282 85689 7380 85787
rect 7664 85666 7762 85764
rect 8060 85666 8158 85764
rect 6425 85315 6523 85413
rect 6850 85257 6948 85355
rect 7282 85257 7380 85355
rect 7664 85271 7762 85369
rect 8060 85271 8158 85369
rect 6425 84899 6523 84997
rect 6850 84899 6948 84997
rect 7282 84899 7380 84997
rect 7664 84876 7762 84974
rect 8060 84876 8158 84974
rect 6425 84525 6523 84623
rect 6850 84467 6948 84565
rect 7282 84467 7380 84565
rect 7664 84481 7762 84579
rect 8060 84481 8158 84579
rect 6425 84109 6523 84207
rect 6850 84109 6948 84207
rect 7282 84109 7380 84207
rect 7664 84086 7762 84184
rect 8060 84086 8158 84184
rect 6425 83735 6523 83833
rect 6850 83677 6948 83775
rect 7282 83677 7380 83775
rect 7664 83691 7762 83789
rect 8060 83691 8158 83789
rect 6425 83319 6523 83417
rect 6850 83319 6948 83417
rect 7282 83319 7380 83417
rect 7664 83296 7762 83394
rect 8060 83296 8158 83394
rect 6425 82945 6523 83043
rect 6850 82887 6948 82985
rect 7282 82887 7380 82985
rect 7664 82901 7762 82999
rect 8060 82901 8158 82999
rect 6425 82529 6523 82627
rect 6850 82529 6948 82627
rect 7282 82529 7380 82627
rect 7664 82506 7762 82604
rect 8060 82506 8158 82604
rect 6425 82155 6523 82253
rect 6850 82097 6948 82195
rect 7282 82097 7380 82195
rect 7664 82111 7762 82209
rect 8060 82111 8158 82209
rect 6425 81739 6523 81837
rect 6850 81739 6948 81837
rect 7282 81739 7380 81837
rect 7664 81716 7762 81814
rect 8060 81716 8158 81814
rect 6425 81365 6523 81463
rect 6850 81307 6948 81405
rect 7282 81307 7380 81405
rect 7664 81321 7762 81419
rect 8060 81321 8158 81419
rect 6425 80949 6523 81047
rect 6850 80949 6948 81047
rect 7282 80949 7380 81047
rect 7664 80926 7762 81024
rect 8060 80926 8158 81024
rect 6425 80575 6523 80673
rect 6850 80517 6948 80615
rect 7282 80517 7380 80615
rect 7664 80531 7762 80629
rect 8060 80531 8158 80629
rect 6425 80159 6523 80257
rect 6850 80159 6948 80257
rect 7282 80159 7380 80257
rect 7664 80136 7762 80234
rect 8060 80136 8158 80234
rect 6425 79785 6523 79883
rect 6850 79727 6948 79825
rect 7282 79727 7380 79825
rect 7664 79741 7762 79839
rect 8060 79741 8158 79839
rect 6425 79369 6523 79467
rect 6850 79369 6948 79467
rect 7282 79369 7380 79467
rect 7664 79346 7762 79444
rect 8060 79346 8158 79444
rect 6425 78995 6523 79093
rect 6850 78937 6948 79035
rect 7282 78937 7380 79035
rect 7664 78951 7762 79049
rect 8060 78951 8158 79049
rect 6425 78579 6523 78677
rect 6850 78579 6948 78677
rect 7282 78579 7380 78677
rect 7664 78556 7762 78654
rect 8060 78556 8158 78654
rect 6425 78205 6523 78303
rect 6850 78147 6948 78245
rect 7282 78147 7380 78245
rect 7664 78161 7762 78259
rect 8060 78161 8158 78259
rect 6425 77789 6523 77887
rect 6850 77789 6948 77887
rect 7282 77789 7380 77887
rect 7664 77766 7762 77864
rect 8060 77766 8158 77864
rect 6425 77415 6523 77513
rect 6850 77357 6948 77455
rect 7282 77357 7380 77455
rect 7664 77371 7762 77469
rect 8060 77371 8158 77469
rect 6425 76999 6523 77097
rect 6850 76999 6948 77097
rect 7282 76999 7380 77097
rect 7664 76976 7762 77074
rect 8060 76976 8158 77074
rect 6425 76625 6523 76723
rect 6850 76567 6948 76665
rect 7282 76567 7380 76665
rect 7664 76581 7762 76679
rect 8060 76581 8158 76679
rect 6425 76209 6523 76307
rect 6850 76209 6948 76307
rect 7282 76209 7380 76307
rect 7664 76186 7762 76284
rect 8060 76186 8158 76284
rect 6425 75835 6523 75933
rect 6850 75777 6948 75875
rect 7282 75777 7380 75875
rect 7664 75791 7762 75889
rect 8060 75791 8158 75889
rect 6425 75419 6523 75517
rect 6850 75419 6948 75517
rect 7282 75419 7380 75517
rect 7664 75396 7762 75494
rect 8060 75396 8158 75494
rect 6425 75045 6523 75143
rect 6850 74987 6948 75085
rect 7282 74987 7380 75085
rect 7664 75001 7762 75099
rect 8060 75001 8158 75099
rect 6425 74629 6523 74727
rect 6850 74629 6948 74727
rect 7282 74629 7380 74727
rect 7664 74606 7762 74704
rect 8060 74606 8158 74704
rect 6425 74255 6523 74353
rect 6850 74197 6948 74295
rect 7282 74197 7380 74295
rect 7664 74211 7762 74309
rect 8060 74211 8158 74309
rect 6425 73839 6523 73937
rect 6850 73839 6948 73937
rect 7282 73839 7380 73937
rect 7664 73816 7762 73914
rect 8060 73816 8158 73914
rect 6425 73465 6523 73563
rect 6850 73407 6948 73505
rect 7282 73407 7380 73505
rect 7664 73421 7762 73519
rect 8060 73421 8158 73519
rect 6425 73049 6523 73147
rect 6850 73049 6948 73147
rect 7282 73049 7380 73147
rect 7664 73026 7762 73124
rect 8060 73026 8158 73124
rect 6425 72675 6523 72773
rect 6850 72617 6948 72715
rect 7282 72617 7380 72715
rect 7664 72631 7762 72729
rect 8060 72631 8158 72729
rect 6425 72259 6523 72357
rect 6850 72259 6948 72357
rect 7282 72259 7380 72357
rect 7664 72236 7762 72334
rect 8060 72236 8158 72334
rect 6425 71885 6523 71983
rect 6850 71827 6948 71925
rect 7282 71827 7380 71925
rect 7664 71841 7762 71939
rect 8060 71841 8158 71939
rect 6425 71469 6523 71567
rect 6850 71469 6948 71567
rect 7282 71469 7380 71567
rect 7664 71446 7762 71544
rect 8060 71446 8158 71544
rect 6425 71095 6523 71193
rect 6850 71037 6948 71135
rect 7282 71037 7380 71135
rect 7664 71051 7762 71149
rect 8060 71051 8158 71149
rect 6425 70679 6523 70777
rect 6850 70679 6948 70777
rect 7282 70679 7380 70777
rect 7664 70656 7762 70754
rect 8060 70656 8158 70754
rect 6425 70305 6523 70403
rect 6850 70247 6948 70345
rect 7282 70247 7380 70345
rect 7664 70261 7762 70359
rect 8060 70261 8158 70359
rect 6425 69889 6523 69987
rect 6850 69889 6948 69987
rect 7282 69889 7380 69987
rect 7664 69866 7762 69964
rect 8060 69866 8158 69964
rect 6425 69515 6523 69613
rect 6850 69457 6948 69555
rect 7282 69457 7380 69555
rect 7664 69471 7762 69569
rect 8060 69471 8158 69569
rect 6425 69099 6523 69197
rect 6850 69099 6948 69197
rect 7282 69099 7380 69197
rect 7664 69076 7762 69174
rect 8060 69076 8158 69174
rect 6425 68725 6523 68823
rect 6850 68667 6948 68765
rect 7282 68667 7380 68765
rect 7664 68681 7762 68779
rect 8060 68681 8158 68779
rect 6425 68309 6523 68407
rect 6850 68309 6948 68407
rect 7282 68309 7380 68407
rect 7664 68286 7762 68384
rect 8060 68286 8158 68384
rect 6425 67935 6523 68033
rect 6850 67877 6948 67975
rect 7282 67877 7380 67975
rect 7664 67891 7762 67989
rect 8060 67891 8158 67989
rect 6425 67519 6523 67617
rect 6850 67519 6948 67617
rect 7282 67519 7380 67617
rect 7664 67496 7762 67594
rect 8060 67496 8158 67594
rect 6425 67145 6523 67243
rect 6850 67087 6948 67185
rect 7282 67087 7380 67185
rect 7664 67101 7762 67199
rect 8060 67101 8158 67199
rect 6425 66729 6523 66827
rect 6850 66729 6948 66827
rect 7282 66729 7380 66827
rect 7664 66706 7762 66804
rect 8060 66706 8158 66804
rect 6425 66355 6523 66453
rect 6850 66297 6948 66395
rect 7282 66297 7380 66395
rect 7664 66311 7762 66409
rect 8060 66311 8158 66409
rect 6425 65939 6523 66037
rect 6850 65939 6948 66037
rect 7282 65939 7380 66037
rect 7664 65916 7762 66014
rect 8060 65916 8158 66014
rect 6425 65565 6523 65663
rect 6850 65507 6948 65605
rect 7282 65507 7380 65605
rect 7664 65521 7762 65619
rect 8060 65521 8158 65619
rect 6425 65149 6523 65247
rect 6850 65149 6948 65247
rect 7282 65149 7380 65247
rect 7664 65126 7762 65224
rect 8060 65126 8158 65224
rect 6425 64775 6523 64873
rect 6850 64717 6948 64815
rect 7282 64717 7380 64815
rect 7664 64731 7762 64829
rect 8060 64731 8158 64829
rect 6425 64359 6523 64457
rect 6850 64359 6948 64457
rect 7282 64359 7380 64457
rect 7664 64336 7762 64434
rect 8060 64336 8158 64434
rect 6425 63985 6523 64083
rect 6850 63927 6948 64025
rect 7282 63927 7380 64025
rect 7664 63941 7762 64039
rect 8060 63941 8158 64039
rect 6425 63569 6523 63667
rect 6850 63569 6948 63667
rect 7282 63569 7380 63667
rect 7664 63546 7762 63644
rect 8060 63546 8158 63644
rect 6425 63195 6523 63293
rect 6850 63137 6948 63235
rect 7282 63137 7380 63235
rect 7664 63151 7762 63249
rect 8060 63151 8158 63249
rect 6425 62779 6523 62877
rect 6850 62779 6948 62877
rect 7282 62779 7380 62877
rect 7664 62756 7762 62854
rect 8060 62756 8158 62854
rect 6425 62405 6523 62503
rect 6850 62347 6948 62445
rect 7282 62347 7380 62445
rect 7664 62361 7762 62459
rect 8060 62361 8158 62459
rect 6425 61989 6523 62087
rect 6850 61989 6948 62087
rect 7282 61989 7380 62087
rect 7664 61966 7762 62064
rect 8060 61966 8158 62064
rect 6425 61615 6523 61713
rect 6850 61557 6948 61655
rect 7282 61557 7380 61655
rect 7664 61571 7762 61669
rect 8060 61571 8158 61669
rect 6425 61199 6523 61297
rect 6850 61199 6948 61297
rect 7282 61199 7380 61297
rect 7664 61176 7762 61274
rect 8060 61176 8158 61274
rect 6425 60825 6523 60923
rect 6850 60767 6948 60865
rect 7282 60767 7380 60865
rect 7664 60781 7762 60879
rect 8060 60781 8158 60879
rect 6425 60409 6523 60507
rect 6850 60409 6948 60507
rect 7282 60409 7380 60507
rect 7664 60386 7762 60484
rect 8060 60386 8158 60484
rect 6425 60035 6523 60133
rect 6850 59977 6948 60075
rect 7282 59977 7380 60075
rect 7664 59991 7762 60089
rect 8060 59991 8158 60089
rect 6425 59619 6523 59717
rect 6850 59619 6948 59717
rect 7282 59619 7380 59717
rect 7664 59596 7762 59694
rect 8060 59596 8158 59694
rect 6425 59245 6523 59343
rect 6850 59187 6948 59285
rect 7282 59187 7380 59285
rect 7664 59201 7762 59299
rect 8060 59201 8158 59299
rect 6425 58829 6523 58927
rect 6850 58829 6948 58927
rect 7282 58829 7380 58927
rect 7664 58806 7762 58904
rect 8060 58806 8158 58904
rect 6425 58455 6523 58553
rect 6850 58397 6948 58495
rect 7282 58397 7380 58495
rect 7664 58411 7762 58509
rect 8060 58411 8158 58509
rect 6425 58039 6523 58137
rect 6850 58039 6948 58137
rect 7282 58039 7380 58137
rect 7664 58016 7762 58114
rect 8060 58016 8158 58114
rect 6425 57665 6523 57763
rect 6850 57607 6948 57705
rect 7282 57607 7380 57705
rect 7664 57621 7762 57719
rect 8060 57621 8158 57719
rect 6425 57249 6523 57347
rect 6850 57249 6948 57347
rect 7282 57249 7380 57347
rect 7664 57226 7762 57324
rect 8060 57226 8158 57324
rect 6425 56875 6523 56973
rect 6850 56817 6948 56915
rect 7282 56817 7380 56915
rect 7664 56831 7762 56929
rect 8060 56831 8158 56929
rect 6425 56459 6523 56557
rect 6850 56459 6948 56557
rect 7282 56459 7380 56557
rect 7664 56436 7762 56534
rect 8060 56436 8158 56534
rect 6425 56085 6523 56183
rect 6850 56027 6948 56125
rect 7282 56027 7380 56125
rect 7664 56041 7762 56139
rect 8060 56041 8158 56139
rect 6425 55669 6523 55767
rect 6850 55669 6948 55767
rect 7282 55669 7380 55767
rect 7664 55646 7762 55744
rect 8060 55646 8158 55744
rect 6425 55295 6523 55393
rect 6850 55237 6948 55335
rect 7282 55237 7380 55335
rect 7664 55251 7762 55349
rect 8060 55251 8158 55349
rect 6425 54879 6523 54977
rect 6850 54879 6948 54977
rect 7282 54879 7380 54977
rect 7664 54856 7762 54954
rect 8060 54856 8158 54954
rect 6425 54505 6523 54603
rect 6850 54447 6948 54545
rect 7282 54447 7380 54545
rect 7664 54461 7762 54559
rect 8060 54461 8158 54559
rect 6425 54089 6523 54187
rect 6850 54089 6948 54187
rect 7282 54089 7380 54187
rect 7664 54066 7762 54164
rect 8060 54066 8158 54164
rect 6425 53715 6523 53813
rect 6850 53657 6948 53755
rect 7282 53657 7380 53755
rect 7664 53671 7762 53769
rect 8060 53671 8158 53769
rect 6425 53299 6523 53397
rect 6850 53299 6948 53397
rect 7282 53299 7380 53397
rect 7664 53276 7762 53374
rect 8060 53276 8158 53374
rect 6425 52925 6523 53023
rect 6850 52867 6948 52965
rect 7282 52867 7380 52965
rect 7664 52881 7762 52979
rect 8060 52881 8158 52979
rect 6425 52509 6523 52607
rect 6850 52509 6948 52607
rect 7282 52509 7380 52607
rect 7664 52486 7762 52584
rect 8060 52486 8158 52584
rect 6425 52135 6523 52233
rect 6850 52077 6948 52175
rect 7282 52077 7380 52175
rect 7664 52091 7762 52189
rect 8060 52091 8158 52189
rect 6425 51719 6523 51817
rect 6850 51719 6948 51817
rect 7282 51719 7380 51817
rect 7664 51696 7762 51794
rect 8060 51696 8158 51794
rect 6425 51345 6523 51443
rect 6850 51287 6948 51385
rect 7282 51287 7380 51385
rect 7664 51301 7762 51399
rect 8060 51301 8158 51399
rect 6425 50929 6523 51027
rect 6850 50929 6948 51027
rect 7282 50929 7380 51027
rect 7664 50906 7762 51004
rect 8060 50906 8158 51004
rect 6425 50555 6523 50653
rect 6850 50497 6948 50595
rect 7282 50497 7380 50595
rect 7664 50511 7762 50609
rect 8060 50511 8158 50609
rect 6425 50139 6523 50237
rect 6850 50139 6948 50237
rect 7282 50139 7380 50237
rect 7664 50116 7762 50214
rect 8060 50116 8158 50214
rect 6425 49765 6523 49863
rect 6850 49707 6948 49805
rect 7282 49707 7380 49805
rect 7664 49721 7762 49819
rect 8060 49721 8158 49819
rect 6425 49349 6523 49447
rect 6850 49349 6948 49447
rect 7282 49349 7380 49447
rect 7664 49326 7762 49424
rect 8060 49326 8158 49424
rect 6425 48975 6523 49073
rect 6850 48917 6948 49015
rect 7282 48917 7380 49015
rect 7664 48931 7762 49029
rect 8060 48931 8158 49029
rect 6425 48559 6523 48657
rect 6850 48559 6948 48657
rect 7282 48559 7380 48657
rect 7664 48536 7762 48634
rect 8060 48536 8158 48634
rect 6425 48185 6523 48283
rect 6850 48127 6948 48225
rect 7282 48127 7380 48225
rect 7664 48141 7762 48239
rect 8060 48141 8158 48239
rect 6425 47769 6523 47867
rect 6850 47769 6948 47867
rect 7282 47769 7380 47867
rect 7664 47746 7762 47844
rect 8060 47746 8158 47844
rect 6425 47395 6523 47493
rect 6850 47337 6948 47435
rect 7282 47337 7380 47435
rect 7664 47351 7762 47449
rect 8060 47351 8158 47449
rect 6425 46979 6523 47077
rect 6850 46979 6948 47077
rect 7282 46979 7380 47077
rect 7664 46956 7762 47054
rect 8060 46956 8158 47054
rect 6425 46605 6523 46703
rect 6850 46547 6948 46645
rect 7282 46547 7380 46645
rect 7664 46561 7762 46659
rect 8060 46561 8158 46659
rect 6425 46189 6523 46287
rect 6850 46189 6948 46287
rect 7282 46189 7380 46287
rect 7664 46166 7762 46264
rect 8060 46166 8158 46264
rect 6425 45815 6523 45913
rect 6850 45757 6948 45855
rect 7282 45757 7380 45855
rect 7664 45771 7762 45869
rect 8060 45771 8158 45869
rect 6425 45399 6523 45497
rect 6850 45399 6948 45497
rect 7282 45399 7380 45497
rect 7664 45376 7762 45474
rect 8060 45376 8158 45474
rect 6425 45025 6523 45123
rect 6850 44967 6948 45065
rect 7282 44967 7380 45065
rect 7664 44981 7762 45079
rect 8060 44981 8158 45079
rect 6425 44609 6523 44707
rect 6850 44609 6948 44707
rect 7282 44609 7380 44707
rect 7664 44586 7762 44684
rect 8060 44586 8158 44684
rect 6425 44235 6523 44333
rect 6850 44177 6948 44275
rect 7282 44177 7380 44275
rect 7664 44191 7762 44289
rect 8060 44191 8158 44289
rect 6425 43819 6523 43917
rect 6850 43819 6948 43917
rect 7282 43819 7380 43917
rect 7664 43796 7762 43894
rect 8060 43796 8158 43894
rect 6425 43445 6523 43543
rect 6850 43387 6948 43485
rect 7282 43387 7380 43485
rect 7664 43401 7762 43499
rect 8060 43401 8158 43499
rect 6425 43029 6523 43127
rect 6850 43029 6948 43127
rect 7282 43029 7380 43127
rect 7664 43006 7762 43104
rect 8060 43006 8158 43104
rect 6425 42655 6523 42753
rect 6850 42597 6948 42695
rect 7282 42597 7380 42695
rect 7664 42611 7762 42709
rect 8060 42611 8158 42709
rect 6425 42239 6523 42337
rect 6850 42239 6948 42337
rect 7282 42239 7380 42337
rect 7664 42216 7762 42314
rect 8060 42216 8158 42314
rect 6425 41865 6523 41963
rect 6850 41807 6948 41905
rect 7282 41807 7380 41905
rect 7664 41821 7762 41919
rect 8060 41821 8158 41919
rect 6425 41449 6523 41547
rect 6850 41449 6948 41547
rect 7282 41449 7380 41547
rect 7664 41426 7762 41524
rect 8060 41426 8158 41524
rect 6425 41075 6523 41173
rect 6850 41017 6948 41115
rect 7282 41017 7380 41115
rect 7664 41031 7762 41129
rect 8060 41031 8158 41129
rect 6425 40659 6523 40757
rect 6850 40659 6948 40757
rect 7282 40659 7380 40757
rect 7664 40636 7762 40734
rect 8060 40636 8158 40734
rect 6425 40285 6523 40383
rect 6850 40227 6948 40325
rect 7282 40227 7380 40325
rect 7664 40241 7762 40339
rect 8060 40241 8158 40339
rect 6425 39869 6523 39967
rect 6850 39869 6948 39967
rect 7282 39869 7380 39967
rect 7664 39846 7762 39944
rect 8060 39846 8158 39944
rect 6425 39495 6523 39593
rect 6850 39437 6948 39535
rect 7282 39437 7380 39535
rect 7664 39451 7762 39549
rect 8060 39451 8158 39549
rect 6425 39079 6523 39177
rect 6850 39079 6948 39177
rect 7282 39079 7380 39177
rect 7664 39056 7762 39154
rect 8060 39056 8158 39154
rect 6425 38705 6523 38803
rect 6850 38647 6948 38745
rect 7282 38647 7380 38745
rect 7664 38661 7762 38759
rect 8060 38661 8158 38759
rect 6425 38289 6523 38387
rect 6850 38289 6948 38387
rect 7282 38289 7380 38387
rect 7664 38266 7762 38364
rect 8060 38266 8158 38364
rect 6425 37915 6523 38013
rect 6850 37857 6948 37955
rect 7282 37857 7380 37955
rect 7664 37871 7762 37969
rect 8060 37871 8158 37969
rect 6425 37499 6523 37597
rect 6850 37499 6948 37597
rect 7282 37499 7380 37597
rect 7664 37476 7762 37574
rect 8060 37476 8158 37574
rect 6425 37125 6523 37223
rect 6850 37067 6948 37165
rect 7282 37067 7380 37165
rect 7664 37081 7762 37179
rect 8060 37081 8158 37179
rect 6425 36709 6523 36807
rect 6850 36709 6948 36807
rect 7282 36709 7380 36807
rect 7664 36686 7762 36784
rect 8060 36686 8158 36784
rect 6425 36335 6523 36433
rect 6850 36277 6948 36375
rect 7282 36277 7380 36375
rect 7664 36291 7762 36389
rect 8060 36291 8158 36389
rect 6425 35919 6523 36017
rect 6850 35919 6948 36017
rect 7282 35919 7380 36017
rect 7664 35896 7762 35994
rect 8060 35896 8158 35994
rect 6425 35545 6523 35643
rect 6850 35487 6948 35585
rect 7282 35487 7380 35585
rect 7664 35501 7762 35599
rect 8060 35501 8158 35599
rect 6425 35129 6523 35227
rect 6850 35129 6948 35227
rect 7282 35129 7380 35227
rect 7664 35106 7762 35204
rect 8060 35106 8158 35204
rect 6425 34755 6523 34853
rect 6850 34697 6948 34795
rect 7282 34697 7380 34795
rect 7664 34711 7762 34809
rect 8060 34711 8158 34809
rect 6425 34339 6523 34437
rect 6850 34339 6948 34437
rect 7282 34339 7380 34437
rect 7664 34316 7762 34414
rect 8060 34316 8158 34414
rect 6425 33965 6523 34063
rect 6850 33907 6948 34005
rect 7282 33907 7380 34005
rect 7664 33921 7762 34019
rect 8060 33921 8158 34019
rect 6425 33549 6523 33647
rect 6850 33549 6948 33647
rect 7282 33549 7380 33647
rect 7664 33526 7762 33624
rect 8060 33526 8158 33624
rect 6425 33175 6523 33273
rect 6850 33117 6948 33215
rect 7282 33117 7380 33215
rect 7664 33131 7762 33229
rect 8060 33131 8158 33229
rect 6425 32759 6523 32857
rect 6850 32759 6948 32857
rect 7282 32759 7380 32857
rect 7664 32736 7762 32834
rect 8060 32736 8158 32834
rect 6425 32385 6523 32483
rect 6850 32327 6948 32425
rect 7282 32327 7380 32425
rect 7664 32341 7762 32439
rect 8060 32341 8158 32439
rect 6425 31969 6523 32067
rect 6850 31969 6948 32067
rect 7282 31969 7380 32067
rect 7664 31946 7762 32044
rect 8060 31946 8158 32044
rect 6425 31595 6523 31693
rect 6850 31537 6948 31635
rect 7282 31537 7380 31635
rect 7664 31551 7762 31649
rect 8060 31551 8158 31649
rect 6425 31179 6523 31277
rect 6850 31179 6948 31277
rect 7282 31179 7380 31277
rect 7664 31156 7762 31254
rect 8060 31156 8158 31254
rect 6425 30805 6523 30903
rect 6850 30747 6948 30845
rect 7282 30747 7380 30845
rect 7664 30761 7762 30859
rect 8060 30761 8158 30859
rect 6425 30389 6523 30487
rect 6850 30389 6948 30487
rect 7282 30389 7380 30487
rect 7664 30366 7762 30464
rect 8060 30366 8158 30464
rect 6425 30015 6523 30113
rect 6850 29957 6948 30055
rect 7282 29957 7380 30055
rect 7664 29971 7762 30069
rect 8060 29971 8158 30069
rect 6425 29599 6523 29697
rect 6850 29599 6948 29697
rect 7282 29599 7380 29697
rect 7664 29576 7762 29674
rect 8060 29576 8158 29674
rect 6425 29225 6523 29323
rect 6850 29167 6948 29265
rect 7282 29167 7380 29265
rect 7664 29181 7762 29279
rect 8060 29181 8158 29279
rect 6425 28809 6523 28907
rect 6850 28809 6948 28907
rect 7282 28809 7380 28907
rect 7664 28786 7762 28884
rect 8060 28786 8158 28884
rect 6425 28435 6523 28533
rect 6850 28377 6948 28475
rect 7282 28377 7380 28475
rect 7664 28391 7762 28489
rect 8060 28391 8158 28489
rect 6425 28019 6523 28117
rect 6850 28019 6948 28117
rect 7282 28019 7380 28117
rect 7664 27996 7762 28094
rect 8060 27996 8158 28094
rect 6425 27645 6523 27743
rect 6850 27587 6948 27685
rect 7282 27587 7380 27685
rect 7664 27601 7762 27699
rect 8060 27601 8158 27699
rect 6425 27229 6523 27327
rect 6850 27229 6948 27327
rect 7282 27229 7380 27327
rect 7664 27206 7762 27304
rect 8060 27206 8158 27304
rect 6425 26855 6523 26953
rect 6850 26797 6948 26895
rect 7282 26797 7380 26895
rect 7664 26811 7762 26909
rect 8060 26811 8158 26909
rect 6425 26439 6523 26537
rect 6850 26439 6948 26537
rect 7282 26439 7380 26537
rect 7664 26416 7762 26514
rect 8060 26416 8158 26514
rect 6425 26065 6523 26163
rect 6850 26007 6948 26105
rect 7282 26007 7380 26105
rect 7664 26021 7762 26119
rect 8060 26021 8158 26119
rect 6425 25649 6523 25747
rect 6850 25649 6948 25747
rect 7282 25649 7380 25747
rect 7664 25626 7762 25724
rect 8060 25626 8158 25724
rect 6425 25275 6523 25373
rect 6850 25217 6948 25315
rect 7282 25217 7380 25315
rect 7664 25231 7762 25329
rect 8060 25231 8158 25329
rect 6425 24859 6523 24957
rect 6850 24859 6948 24957
rect 7282 24859 7380 24957
rect 7664 24836 7762 24934
rect 8060 24836 8158 24934
rect 6425 24485 6523 24583
rect 6850 24427 6948 24525
rect 7282 24427 7380 24525
rect 7664 24441 7762 24539
rect 8060 24441 8158 24539
rect 6425 24069 6523 24167
rect 6850 24069 6948 24167
rect 7282 24069 7380 24167
rect 7664 24046 7762 24144
rect 8060 24046 8158 24144
rect 6425 23695 6523 23793
rect 6850 23637 6948 23735
rect 7282 23637 7380 23735
rect 7664 23651 7762 23749
rect 8060 23651 8158 23749
rect 6425 23279 6523 23377
rect 6850 23279 6948 23377
rect 7282 23279 7380 23377
rect 7664 23256 7762 23354
rect 8060 23256 8158 23354
rect 6425 22905 6523 23003
rect 6850 22847 6948 22945
rect 7282 22847 7380 22945
rect 7664 22861 7762 22959
rect 8060 22861 8158 22959
rect 6425 22489 6523 22587
rect 6850 22489 6948 22587
rect 7282 22489 7380 22587
rect 7664 22466 7762 22564
rect 8060 22466 8158 22564
rect 6425 22115 6523 22213
rect 6850 22057 6948 22155
rect 7282 22057 7380 22155
rect 7664 22071 7762 22169
rect 8060 22071 8158 22169
rect 6425 21699 6523 21797
rect 6850 21699 6948 21797
rect 7282 21699 7380 21797
rect 7664 21676 7762 21774
rect 8060 21676 8158 21774
rect 6425 21325 6523 21423
rect 6850 21267 6948 21365
rect 7282 21267 7380 21365
rect 7664 21281 7762 21379
rect 8060 21281 8158 21379
rect 6425 20909 6523 21007
rect 6850 20909 6948 21007
rect 7282 20909 7380 21007
rect 7664 20886 7762 20984
rect 8060 20886 8158 20984
rect 6425 20535 6523 20633
rect 6850 20477 6948 20575
rect 7282 20477 7380 20575
rect 7664 20491 7762 20589
rect 8060 20491 8158 20589
rect 6425 20119 6523 20217
rect 6850 20119 6948 20217
rect 7282 20119 7380 20217
rect 7664 20096 7762 20194
rect 8060 20096 8158 20194
rect 6425 19745 6523 19843
rect 6850 19687 6948 19785
rect 7282 19687 7380 19785
rect 7664 19701 7762 19799
rect 8060 19701 8158 19799
rect 6425 19329 6523 19427
rect 6850 19329 6948 19427
rect 7282 19329 7380 19427
rect 7664 19306 7762 19404
rect 8060 19306 8158 19404
rect 6425 18955 6523 19053
rect 6850 18897 6948 18995
rect 7282 18897 7380 18995
rect 7664 18911 7762 19009
rect 8060 18911 8158 19009
rect 6425 18539 6523 18637
rect 6850 18539 6948 18637
rect 7282 18539 7380 18637
rect 7664 18516 7762 18614
rect 8060 18516 8158 18614
rect 6425 18165 6523 18263
rect 6850 18107 6948 18205
rect 7282 18107 7380 18205
rect 7664 18121 7762 18219
rect 8060 18121 8158 18219
rect 6425 17749 6523 17847
rect 6850 17749 6948 17847
rect 7282 17749 7380 17847
rect 7664 17726 7762 17824
rect 8060 17726 8158 17824
rect 6425 17375 6523 17473
rect 6850 17317 6948 17415
rect 7282 17317 7380 17415
rect 7664 17331 7762 17429
rect 8060 17331 8158 17429
rect 6425 16959 6523 17057
rect 6850 16959 6948 17057
rect 7282 16959 7380 17057
rect 7664 16936 7762 17034
rect 8060 16936 8158 17034
rect 6425 16585 6523 16683
rect 6850 16527 6948 16625
rect 7282 16527 7380 16625
rect 7664 16541 7762 16639
rect 8060 16541 8158 16639
rect 6425 16169 6523 16267
rect 6850 16169 6948 16267
rect 7282 16169 7380 16267
rect 7664 16146 7762 16244
rect 8060 16146 8158 16244
rect 6425 15795 6523 15893
rect 6850 15737 6948 15835
rect 7282 15737 7380 15835
rect 7664 15751 7762 15849
rect 8060 15751 8158 15849
rect 6425 15379 6523 15477
rect 6850 15379 6948 15477
rect 7282 15379 7380 15477
rect 7664 15356 7762 15454
rect 8060 15356 8158 15454
rect 6425 15005 6523 15103
rect 6850 14947 6948 15045
rect 7282 14947 7380 15045
rect 7664 14961 7762 15059
rect 8060 14961 8158 15059
rect 6425 14589 6523 14687
rect 6850 14589 6948 14687
rect 7282 14589 7380 14687
rect 7664 14566 7762 14664
rect 8060 14566 8158 14664
rect 6425 14215 6523 14313
rect 6850 14157 6948 14255
rect 7282 14157 7380 14255
rect 7664 14171 7762 14269
rect 8060 14171 8158 14269
rect 6425 13799 6523 13897
rect 6850 13799 6948 13897
rect 7282 13799 7380 13897
rect 7664 13776 7762 13874
rect 8060 13776 8158 13874
rect 6425 13425 6523 13523
rect 6850 13367 6948 13465
rect 7282 13367 7380 13465
rect 7664 13381 7762 13479
rect 8060 13381 8158 13479
rect 6425 13009 6523 13107
rect 6850 13009 6948 13107
rect 7282 13009 7380 13107
rect 7664 12986 7762 13084
rect 8060 12986 8158 13084
rect 6425 12635 6523 12733
rect 6850 12577 6948 12675
rect 7282 12577 7380 12675
rect 7664 12591 7762 12689
rect 8060 12591 8158 12689
rect 6425 12219 6523 12317
rect 6850 12219 6948 12317
rect 7282 12219 7380 12317
rect 7664 12196 7762 12294
rect 8060 12196 8158 12294
rect 6425 11845 6523 11943
rect 6850 11787 6948 11885
rect 7282 11787 7380 11885
rect 7664 11801 7762 11899
rect 8060 11801 8158 11899
rect 6425 11429 6523 11527
rect 6850 11429 6948 11527
rect 7282 11429 7380 11527
rect 7664 11406 7762 11504
rect 8060 11406 8158 11504
rect 6425 11055 6523 11153
rect 6850 10997 6948 11095
rect 7282 10997 7380 11095
rect 7664 11011 7762 11109
rect 8060 11011 8158 11109
rect 6425 10639 6523 10737
rect 6850 10639 6948 10737
rect 7282 10639 7380 10737
rect 7664 10616 7762 10714
rect 8060 10616 8158 10714
rect 6425 10265 6523 10363
rect 6850 10207 6948 10305
rect 7282 10207 7380 10305
rect 7664 10221 7762 10319
rect 8060 10221 8158 10319
rect 6425 9849 6523 9947
rect 6850 9849 6948 9947
rect 7282 9849 7380 9947
rect 7664 9826 7762 9924
rect 8060 9826 8158 9924
rect 6425 9475 6523 9573
rect 6850 9417 6948 9515
rect 7282 9417 7380 9515
rect 7664 9431 7762 9529
rect 8060 9431 8158 9529
rect 2691 9059 2789 9157
rect 3116 9059 3214 9157
rect 3548 9059 3646 9157
rect 3930 9036 4028 9134
rect 4326 9036 4424 9134
rect 6425 9059 6523 9157
rect 6850 9059 6948 9157
rect 7282 9059 7380 9157
rect 7664 9036 7762 9134
rect 8060 9036 8158 9134
rect 6425 8685 6523 8783
rect 6850 8627 6948 8725
rect 7282 8627 7380 8725
rect 7664 8641 7762 8739
rect 8060 8641 8158 8739
rect 2691 8269 2789 8367
rect 3116 8269 3214 8367
rect 3548 8269 3646 8367
rect 3930 8246 4028 8344
rect 4326 8246 4424 8344
rect 6425 8269 6523 8367
rect 6850 8269 6948 8367
rect 7282 8269 7380 8367
rect 7664 8246 7762 8344
rect 8060 8246 8158 8344
rect 6425 7895 6523 7993
rect 6850 7837 6948 7935
rect 7282 7837 7380 7935
rect 7664 7851 7762 7949
rect 8060 7851 8158 7949
rect 2691 7479 2789 7577
rect 3116 7479 3214 7577
rect 3548 7479 3646 7577
rect 3930 7456 4028 7554
rect 4326 7456 4424 7554
rect 6425 7479 6523 7577
rect 6850 7479 6948 7577
rect 7282 7479 7380 7577
rect 7664 7456 7762 7554
rect 8060 7456 8158 7554
rect 6425 7105 6523 7203
rect 6850 7047 6948 7145
rect 7282 7047 7380 7145
rect 7664 7061 7762 7159
rect 8060 7061 8158 7159
rect 1236 6666 1334 6764
rect 1632 6666 1730 6764
rect 2691 6689 2789 6787
rect 3116 6689 3214 6787
rect 3548 6689 3646 6787
rect 3930 6666 4028 6764
rect 4326 6666 4424 6764
rect 6425 6689 6523 6787
rect 6850 6689 6948 6787
rect 7282 6689 7380 6787
rect 7664 6666 7762 6764
rect 8060 6666 8158 6764
rect 6425 6315 6523 6413
rect 6850 6257 6948 6355
rect 7282 6257 7380 6355
rect 7664 6271 7762 6369
rect 8060 6271 8158 6369
rect 6425 5899 6523 5997
rect 6850 5899 6948 5997
rect 7282 5899 7380 5997
rect 7664 5876 7762 5974
rect 8060 5876 8158 5974
rect 6425 5525 6523 5623
rect 6850 5467 6948 5565
rect 7282 5467 7380 5565
rect 7664 5481 7762 5579
rect 8060 5481 8158 5579
rect 2691 5109 2789 5207
rect 3116 5109 3214 5207
rect 3548 5109 3646 5207
rect 3930 5086 4028 5184
rect 4326 5086 4424 5184
rect 6425 5109 6523 5207
rect 6850 5109 6948 5207
rect 7282 5109 7380 5207
rect 7664 5086 7762 5184
rect 8060 5086 8158 5184
rect 6425 4735 6523 4833
rect 6850 4677 6948 4775
rect 7282 4677 7380 4775
rect 7664 4691 7762 4789
rect 8060 4691 8158 4789
rect 2691 4319 2789 4417
rect 3116 4319 3214 4417
rect 3548 4319 3646 4417
rect 3930 4296 4028 4394
rect 4326 4296 4424 4394
rect 6425 4319 6523 4417
rect 6850 4319 6948 4417
rect 7282 4319 7380 4417
rect 7664 4296 7762 4394
rect 8060 4296 8158 4394
rect 6425 3945 6523 4043
rect 6850 3887 6948 3985
rect 7282 3887 7380 3985
rect 7664 3901 7762 3999
rect 8060 3901 8158 3999
rect 2691 3529 2789 3627
rect 3116 3529 3214 3627
rect 3548 3529 3646 3627
rect 3930 3506 4028 3604
rect 4326 3506 4424 3604
rect 6425 3529 6523 3627
rect 6850 3529 6948 3627
rect 7282 3529 7380 3627
rect 7664 3506 7762 3604
rect 8060 3506 8158 3604
rect 6425 3155 6523 3253
rect 6850 3097 6948 3195
rect 7282 3097 7380 3195
rect 7664 3111 7762 3209
rect 8060 3111 8158 3209
rect 1236 2716 1334 2814
rect 1632 2716 1730 2814
rect 2691 2739 2789 2837
rect 3116 2739 3214 2837
rect 3548 2739 3646 2837
rect 3930 2716 4028 2814
rect 4326 2716 4424 2814
rect 6425 2739 6523 2837
rect 6850 2739 6948 2837
rect 7282 2739 7380 2837
rect 7664 2716 7762 2814
rect 8060 2716 8158 2814
rect 6425 2365 6523 2463
rect 6850 2307 6948 2405
rect 7282 2307 7380 2405
rect 7664 2321 7762 2419
rect 8060 2321 8158 2419
rect 6425 1949 6523 2047
rect 6850 1949 6948 2047
rect 7282 1949 7380 2047
rect 7664 1926 7762 2024
rect 8060 1926 8158 2024
rect 6425 1575 6523 1673
rect 6850 1517 6948 1615
rect 7282 1517 7380 1615
rect 7664 1531 7762 1629
rect 8060 1531 8158 1629
rect 3126 1143 3224 1241
rect 3551 1143 3649 1241
rect 3930 1136 4028 1234
rect 4326 1136 4424 1234
rect 6425 1159 6523 1257
rect 6850 1159 6948 1257
rect 7282 1159 7380 1257
rect 7664 1136 7762 1234
rect 8060 1136 8158 1234
rect 6425 785 6523 883
rect 6850 727 6948 825
rect 7282 727 7380 825
rect 7664 741 7762 839
rect 8060 741 8158 839
rect 1832 346 1930 444
rect 2228 346 2326 444
rect 3126 353 3224 451
rect 3551 353 3649 451
rect 3930 346 4028 444
rect 4326 346 4424 444
rect 6425 369 6523 467
rect 6850 369 6948 467
rect 7282 369 7380 467
rect 7664 346 7762 444
rect 8060 346 8158 444
use contact_16  contact_16_775
timestamp 1624494425
transform 1 0 0 0 1 141
box 0 0 66 58
use contact_16  contact_16_774
timestamp 1624494425
transform 1 0 80 0 1 591
box 0 0 66 58
use contact_7  contact_7_26
timestamp 1624494425
transform 1 0 1508 0 1 587
box 0 0 58 66
use contact_7  contact_7_27
timestamp 1624494425
transform 1 0 1428 0 1 137
box 0 0 58 66
use contact_16  contact_16_773
timestamp 1624494425
transform 1 0 160 0 1 2511
box 0 0 66 58
use contact_16  contact_16_772
timestamp 1624494425
transform 1 0 240 0 1 2961
box 0 0 66 58
use contact_7  contact_7_24
timestamp 1624494425
transform 1 0 832 0 1 2957
box 0 0 58 66
use contact_7  contact_7_25
timestamp 1624494425
transform 1 0 752 0 1 2507
box 0 0 58 66
use hierarchical_predecode3x8  hierarchical_predecode3x8_1
timestamp 1624494425
transform 1 0 687 0 1 2370
box 61 -60 3854 3220
use hierarchical_predecode2x4  hierarchical_predecode2x4_0
timestamp 1624494425
transform 1 0 1363 0 1 0
box 61 -56 3178 1636
use contact_7  contact_7_19
timestamp 1624494425
transform 1 0 4494 0 1 87
box 0 0 58 66
use contact_8  contact_8_1294
timestamp 1624494425
transform 1 0 4491 0 1 88
box 0 0 64 64
use contact_16  contact_16_766
timestamp 1624494425
transform 1 0 4904 0 1 164
box 0 0 66 58
use contact_16  contact_16_767
timestamp 1624494425
transform 1 0 4584 0 1 52
box 0 0 66 58
use contact_17  contact_17_19
timestamp 1624494425
transform 1 0 4585 0 1 -32
box 0 0 64 64
use contact_8  contact_8_1274
timestamp 1624494425
transform 1 0 7299 0 1 386
box 0 0 64 64
use contact_9  contact_9_1274
timestamp 1624494425
transform 1 0 7298 0 1 381
box 0 0 66 74
use contact_8  contact_8_1273
timestamp 1624494425
transform 1 0 6867 0 1 386
box 0 0 64 64
use contact_9  contact_9_1273
timestamp 1624494425
transform 1 0 6866 0 1 381
box 0 0 66 74
use contact_8  contact_8_509
timestamp 1624494425
transform 1 0 6442 0 1 386
box 0 0 64 64
use contact_9  contact_9_509
timestamp 1624494425
transform 1 0 6441 0 1 381
box 0 0 66 74
use contact_16  contact_16_762
timestamp 1624494425
transform 1 0 5544 0 1 478
box 0 0 66 58
use contact_16  contact_16_765
timestamp 1624494425
transform 1 0 5544 0 1 254
box 0 0 66 58
use contact_17  contact_17_18
timestamp 1624494425
transform 1 0 4665 0 1 363
box 0 0 64 64
use and3_dec  and3_dec_254
timestamp 1624494425
transform 1 0 6203 0 -1 790
box 0 -60 2072 490
use and3_dec  and3_dec_255
timestamp 1624494425
transform 1 0 6203 0 1 0
box 0 -60 2072 490
use contact_7  contact_7_18
timestamp 1624494425
transform 1 0 4494 0 1 637
box 0 0 58 66
use contact_8  contact_8_1293
timestamp 1624494425
transform 1 0 4491 0 1 638
box 0 0 64 64
use contact_8  contact_8_1271
timestamp 1624494425
transform 1 0 7299 0 1 744
box 0 0 64 64
use contact_9  contact_9_1271
timestamp 1624494425
transform 1 0 7298 0 1 739
box 0 0 66 74
use contact_8  contact_8_1270
timestamp 1624494425
transform 1 0 6867 0 1 744
box 0 0 64 64
use contact_9  contact_9_1270
timestamp 1624494425
transform 1 0 6866 0 1 739
box 0 0 66 74
use contact_16  contact_16_763
timestamp 1624494425
transform 1 0 4904 0 1 568
box 0 0 66 58
use contact_16  contact_16_764
timestamp 1624494425
transform 1 0 4664 0 1 680
box 0 0 66 58
use contact_17  contact_17_17
timestamp 1624494425
transform 1 0 4745 0 1 758
box 0 0 64 64
use contact_7  contact_7_17
timestamp 1624494425
transform 1 0 4494 0 1 877
box 0 0 58 66
use contact_8  contact_8_1292
timestamp 1624494425
transform 1 0 4491 0 1 878
box 0 0 64 64
use contact_8  contact_8_507
timestamp 1624494425
transform 1 0 6442 0 1 802
box 0 0 64 64
use contact_9  contact_9_507
timestamp 1624494425
transform 1 0 6441 0 1 797
box 0 0 66 74
use contact_16  contact_16_760
timestamp 1624494425
transform 1 0 4904 0 1 954
box 0 0 66 58
use contact_16  contact_16_761
timestamp 1624494425
transform 1 0 4744 0 1 842
box 0 0 66 58
use and3_dec  and3_dec_253
timestamp 1624494425
transform 1 0 6203 0 1 790
box 0 -60 2072 490
use contact_8  contact_8_1268
timestamp 1624494425
transform 1 0 7299 0 1 1176
box 0 0 64 64
use contact_9  contact_9_1268
timestamp 1624494425
transform 1 0 7298 0 1 1171
box 0 0 66 74
use contact_8  contact_8_1267
timestamp 1624494425
transform 1 0 6867 0 1 1176
box 0 0 64 64
use contact_9  contact_9_1267
timestamp 1624494425
transform 1 0 6866 0 1 1171
box 0 0 66 74
use contact_8  contact_8_505
timestamp 1624494425
transform 1 0 6442 0 1 1176
box 0 0 64 64
use contact_9  contact_9_505
timestamp 1624494425
transform 1 0 6441 0 1 1171
box 0 0 66 74
use contact_16  contact_16_756
timestamp 1624494425
transform 1 0 5544 0 1 1268
box 0 0 66 58
use contact_16  contact_16_759
timestamp 1624494425
transform 1 0 5544 0 1 1044
box 0 0 66 58
use contact_17  contact_17_16
timestamp 1624494425
transform 1 0 4825 0 1 1153
box 0 0 64 64
use contact_8  contact_8_1291
timestamp 1624494425
transform 1 0 4491 0 1 1428
box 0 0 64 64
use contact_7  contact_7_16
timestamp 1624494425
transform 1 0 4494 0 1 1427
box 0 0 58 66
use contact_16  contact_16_758
timestamp 1624494425
transform 1 0 4824 0 1 1470
box 0 0 66 58
use contact_16  contact_16_757
timestamp 1624494425
transform 1 0 4904 0 1 1358
box 0 0 66 58
use contact_9  contact_9_503
timestamp 1624494425
transform 1 0 6441 0 1 1587
box 0 0 66 74
use contact_8  contact_8_503
timestamp 1624494425
transform 1 0 6442 0 1 1592
box 0 0 64 64
use contact_9  contact_9_1264
timestamp 1624494425
transform 1 0 6866 0 1 1529
box 0 0 66 74
use contact_8  contact_8_1264
timestamp 1624494425
transform 1 0 6867 0 1 1534
box 0 0 64 64
use contact_9  contact_9_1265
timestamp 1624494425
transform 1 0 7298 0 1 1529
box 0 0 66 74
use contact_8  contact_8_1265
timestamp 1624494425
transform 1 0 7299 0 1 1534
box 0 0 64 64
use and3_dec  and3_dec_251
timestamp 1624494425
transform 1 0 6203 0 1 1580
box 0 -60 2072 490
use and3_dec  and3_dec_252
timestamp 1624494425
transform 1 0 6203 0 -1 1580
box 0 -60 2072 490
use contact_16  contact_16_753
timestamp 1624494425
transform 1 0 5544 0 1 1834
box 0 0 66 58
use contact_16  contact_16_754
timestamp 1624494425
transform 1 0 4984 0 1 1744
box 0 0 66 58
use contact_16  contact_16_755
timestamp 1624494425
transform 1 0 4584 0 1 1632
box 0 0 66 58
use contact_8  contact_8_1262
timestamp 1624494425
transform 1 0 7299 0 1 1966
box 0 0 64 64
use contact_9  contact_9_1262
timestamp 1624494425
transform 1 0 7298 0 1 1961
box 0 0 66 74
use contact_8  contact_8_1261
timestamp 1624494425
transform 1 0 6867 0 1 1966
box 0 0 64 64
use contact_9  contact_9_1261
timestamp 1624494425
transform 1 0 6866 0 1 1961
box 0 0 66 74
use contact_8  contact_8_501
timestamp 1624494425
transform 1 0 6442 0 1 1966
box 0 0 64 64
use contact_9  contact_9_501
timestamp 1624494425
transform 1 0 6441 0 1 1961
box 0 0 66 74
use contact_16  contact_16_750
timestamp 1624494425
transform 1 0 5544 0 1 2058
box 0 0 66 58
use and3_dec  and3_dec_250
timestamp 1624494425
transform 1 0 6203 0 -1 2370
box 0 -60 2072 490
use contact_8  contact_8_1259
timestamp 1624494425
transform 1 0 7299 0 1 2324
box 0 0 64 64
use contact_9  contact_9_1259
timestamp 1624494425
transform 1 0 7298 0 1 2319
box 0 0 66 74
use contact_8  contact_8_1258
timestamp 1624494425
transform 1 0 6867 0 1 2324
box 0 0 64 64
use contact_9  contact_9_1258
timestamp 1624494425
transform 1 0 6866 0 1 2319
box 0 0 66 74
use contact_8  contact_8_499
timestamp 1624494425
transform 1 0 6442 0 1 2382
box 0 0 64 64
use contact_9  contact_9_499
timestamp 1624494425
transform 1 0 6441 0 1 2377
box 0 0 66 74
use contact_16  contact_16_751
timestamp 1624494425
transform 1 0 4984 0 1 2148
box 0 0 66 58
use contact_16  contact_16_752
timestamp 1624494425
transform 1 0 4664 0 1 2260
box 0 0 66 58
use contact_17  contact_17_15
timestamp 1624494425
transform 1 0 4905 0 1 2338
box 0 0 64 64
use contact_7  contact_7_15
timestamp 1624494425
transform 1 0 4494 0 1 2457
box 0 0 58 66
use contact_8  contact_8_1290
timestamp 1624494425
transform 1 0 4491 0 1 2458
box 0 0 64 64
use contact_16  contact_16_747
timestamp 1624494425
transform 1 0 5544 0 1 2624
box 0 0 66 58
use contact_16  contact_16_748
timestamp 1624494425
transform 1 0 4984 0 1 2534
box 0 0 66 58
use contact_16  contact_16_749
timestamp 1624494425
transform 1 0 4744 0 1 2422
box 0 0 66 58
use and3_dec  and3_dec_248
timestamp 1624494425
transform 1 0 6203 0 -1 3160
box 0 -60 2072 490
use and3_dec  and3_dec_249
timestamp 1624494425
transform 1 0 6203 0 1 2370
box 0 -60 2072 490
use contact_8  contact_8_1256
timestamp 1624494425
transform 1 0 7299 0 1 2756
box 0 0 64 64
use contact_9  contact_9_1256
timestamp 1624494425
transform 1 0 7298 0 1 2751
box 0 0 66 74
use contact_8  contact_8_1255
timestamp 1624494425
transform 1 0 6867 0 1 2756
box 0 0 64 64
use contact_9  contact_9_1255
timestamp 1624494425
transform 1 0 6866 0 1 2751
box 0 0 66 74
use contact_8  contact_8_497
timestamp 1624494425
transform 1 0 6442 0 1 2756
box 0 0 64 64
use contact_9  contact_9_497
timestamp 1624494425
transform 1 0 6441 0 1 2751
box 0 0 66 74
use contact_16  contact_16_744
timestamp 1624494425
transform 1 0 5544 0 1 2848
box 0 0 66 58
use contact_16  contact_16_745
timestamp 1624494425
transform 1 0 4984 0 1 2938
box 0 0 66 58
use contact_17  contact_17_14
timestamp 1624494425
transform 1 0 4985 0 1 2733
box 0 0 64 64
use contact_16  contact_16_746
timestamp 1624494425
transform 1 0 4824 0 1 3050
box 0 0 66 58
use contact_16  contact_16_743
timestamp 1624494425
transform 1 0 4584 0 1 3212
box 0 0 66 58
use contact_8  contact_8_1289
timestamp 1624494425
transform 1 0 4491 0 1 3008
box 0 0 64 64
use contact_7  contact_7_14
timestamp 1624494425
transform 1 0 4494 0 1 3007
box 0 0 58 66
use contact_17  contact_17_13
timestamp 1624494425
transform 1 0 5065 0 1 3128
box 0 0 64 64
use contact_9  contact_9_495
timestamp 1624494425
transform 1 0 6441 0 1 3167
box 0 0 66 74
use contact_8  contact_8_495
timestamp 1624494425
transform 1 0 6442 0 1 3172
box 0 0 64 64
use contact_9  contact_9_1252
timestamp 1624494425
transform 1 0 6866 0 1 3109
box 0 0 66 74
use contact_8  contact_8_1252
timestamp 1624494425
transform 1 0 6867 0 1 3114
box 0 0 64 64
use contact_9  contact_9_1253
timestamp 1624494425
transform 1 0 7298 0 1 3109
box 0 0 66 74
use contact_8  contact_8_1253
timestamp 1624494425
transform 1 0 7299 0 1 3114
box 0 0 64 64
use and3_dec  and3_dec_247
timestamp 1624494425
transform 1 0 6203 0 1 3160
box 0 -60 2072 490
use contact_9  contact_9_508
timestamp 1624494425
transform 1 0 7680 0 1 358
box 0 0 66 74
use contact_8  contact_8_508
timestamp 1624494425
transform 1 0 7681 0 1 363
box 0 0 64 64
use contact_9  contact_9_1272
timestamp 1624494425
transform 1 0 8076 0 1 358
box 0 0 66 74
use contact_8  contact_8_1272
timestamp 1624494425
transform 1 0 8077 0 1 363
box 0 0 64 64
use contact_9  contact_9_504
timestamp 1624494425
transform 1 0 7680 0 1 1148
box 0 0 66 74
use contact_8  contact_8_504
timestamp 1624494425
transform 1 0 7681 0 1 1153
box 0 0 64 64
use contact_9  contact_9_506
timestamp 1624494425
transform 1 0 7680 0 1 753
box 0 0 66 74
use contact_8  contact_8_506
timestamp 1624494425
transform 1 0 7681 0 1 758
box 0 0 64 64
use contact_9  contact_9_1266
timestamp 1624494425
transform 1 0 8076 0 1 1148
box 0 0 66 74
use contact_8  contact_8_1266
timestamp 1624494425
transform 1 0 8077 0 1 1153
box 0 0 64 64
use contact_9  contact_9_1269
timestamp 1624494425
transform 1 0 8076 0 1 753
box 0 0 66 74
use contact_8  contact_8_1269
timestamp 1624494425
transform 1 0 8077 0 1 758
box 0 0 64 64
use contact_9  contact_9_502
timestamp 1624494425
transform 1 0 7680 0 1 1543
box 0 0 66 74
use contact_8  contact_8_502
timestamp 1624494425
transform 1 0 7681 0 1 1548
box 0 0 64 64
use contact_9  contact_9_1263
timestamp 1624494425
transform 1 0 8076 0 1 1543
box 0 0 66 74
use contact_8  contact_8_1263
timestamp 1624494425
transform 1 0 8077 0 1 1548
box 0 0 64 64
use contact_9  contact_9_498
timestamp 1624494425
transform 1 0 7680 0 1 2333
box 0 0 66 74
use contact_8  contact_8_498
timestamp 1624494425
transform 1 0 7681 0 1 2338
box 0 0 64 64
use contact_9  contact_9_500
timestamp 1624494425
transform 1 0 7680 0 1 1938
box 0 0 66 74
use contact_8  contact_8_500
timestamp 1624494425
transform 1 0 7681 0 1 1943
box 0 0 64 64
use contact_9  contact_9_1257
timestamp 1624494425
transform 1 0 8076 0 1 2333
box 0 0 66 74
use contact_8  contact_8_1257
timestamp 1624494425
transform 1 0 8077 0 1 2338
box 0 0 64 64
use contact_9  contact_9_1260
timestamp 1624494425
transform 1 0 8076 0 1 1938
box 0 0 66 74
use contact_8  contact_8_1260
timestamp 1624494425
transform 1 0 8077 0 1 1943
box 0 0 64 64
use contact_9  contact_9_496
timestamp 1624494425
transform 1 0 7680 0 1 2728
box 0 0 66 74
use contact_8  contact_8_496
timestamp 1624494425
transform 1 0 7681 0 1 2733
box 0 0 64 64
use contact_9  contact_9_1254
timestamp 1624494425
transform 1 0 8076 0 1 2728
box 0 0 66 74
use contact_8  contact_8_1254
timestamp 1624494425
transform 1 0 8077 0 1 2733
box 0 0 64 64
use contact_9  contact_9_494
timestamp 1624494425
transform 1 0 7680 0 1 3123
box 0 0 66 74
use contact_8  contact_8_494
timestamp 1624494425
transform 1 0 7681 0 1 3128
box 0 0 64 64
use contact_9  contact_9_1251
timestamp 1624494425
transform 1 0 8076 0 1 3123
box 0 0 66 74
use contact_8  contact_8_1251
timestamp 1624494425
transform 1 0 8077 0 1 3128
box 0 0 64 64
use contact_7  contact_7_23
timestamp 1624494425
transform 1 0 912 0 1 3297
box 0 0 58 66
use contact_7  contact_7_22
timestamp 1624494425
transform 1 0 752 0 1 6457
box 0 0 58 66
use contact_16  contact_16_770
timestamp 1624494425
transform 1 0 400 0 1 6461
box 0 0 66 58
use contact_16  contact_16_771
timestamp 1624494425
transform 1 0 320 0 1 3301
box 0 0 66 58
use hierarchical_predecode3x8  hierarchical_predecode3x8_0
timestamp 1624494425
transform 1 0 687 0 1 6320
box 61 -60 3854 3220
use contact_7  contact_7_13
timestamp 1624494425
transform 1 0 4494 0 1 3247
box 0 0 58 66
use contact_8  contact_8_1288
timestamp 1624494425
transform 1 0 4491 0 1 3248
box 0 0 64 64
use contact_16  contact_16_741
timestamp 1624494425
transform 1 0 5544 0 1 3414
box 0 0 66 58
use contact_16  contact_16_742
timestamp 1624494425
transform 1 0 5064 0 1 3324
box 0 0 66 58
use contact_8  contact_8_1250
timestamp 1624494425
transform 1 0 7299 0 1 3546
box 0 0 64 64
use contact_9  contact_9_1250
timestamp 1624494425
transform 1 0 7298 0 1 3541
box 0 0 66 74
use contact_8  contact_8_1249
timestamp 1624494425
transform 1 0 6867 0 1 3546
box 0 0 64 64
use contact_9  contact_9_1249
timestamp 1624494425
transform 1 0 6866 0 1 3541
box 0 0 66 74
use contact_8  contact_8_493
timestamp 1624494425
transform 1 0 6442 0 1 3546
box 0 0 64 64
use contact_9  contact_9_493
timestamp 1624494425
transform 1 0 6441 0 1 3541
box 0 0 66 74
use contact_16  contact_16_738
timestamp 1624494425
transform 1 0 5544 0 1 3638
box 0 0 66 58
use contact_16  contact_16_739
timestamp 1624494425
transform 1 0 5064 0 1 3728
box 0 0 66 58
use contact_17  contact_17_12
timestamp 1624494425
transform 1 0 5145 0 1 3523
box 0 0 64 64
use and3_dec  and3_dec_246
timestamp 1624494425
transform 1 0 6203 0 -1 3950
box 0 -60 2072 490
use contact_16  contact_16_740
timestamp 1624494425
transform 1 0 4664 0 1 3840
box 0 0 66 58
use contact_8  contact_8_1286
timestamp 1624494425
transform 1 0 4491 0 1 4038
box 0 0 64 64
use contact_7  contact_7_11
timestamp 1624494425
transform 1 0 4494 0 1 4037
box 0 0 58 66
use contact_8  contact_8_1287
timestamp 1624494425
transform 1 0 4491 0 1 3798
box 0 0 64 64
use contact_7  contact_7_12
timestamp 1624494425
transform 1 0 4494 0 1 3797
box 0 0 58 66
use contact_16  contact_16_737
timestamp 1624494425
transform 1 0 4744 0 1 4002
box 0 0 66 58
use contact_17  contact_17_11
timestamp 1624494425
transform 1 0 5225 0 1 3918
box 0 0 64 64
use contact_9  contact_9_491
timestamp 1624494425
transform 1 0 6441 0 1 3957
box 0 0 66 74
use contact_8  contact_8_491
timestamp 1624494425
transform 1 0 6442 0 1 3962
box 0 0 64 64
use contact_9  contact_9_1246
timestamp 1624494425
transform 1 0 6866 0 1 3899
box 0 0 66 74
use contact_8  contact_8_1246
timestamp 1624494425
transform 1 0 6867 0 1 3904
box 0 0 64 64
use contact_9  contact_9_1247
timestamp 1624494425
transform 1 0 7298 0 1 3899
box 0 0 66 74
use contact_8  contact_8_1247
timestamp 1624494425
transform 1 0 7299 0 1 3904
box 0 0 64 64
use contact_16  contact_16_735
timestamp 1624494425
transform 1 0 5544 0 1 4204
box 0 0 66 58
use contact_16  contact_16_736
timestamp 1624494425
transform 1 0 5064 0 1 4114
box 0 0 66 58
use contact_17  contact_17_10
timestamp 1624494425
transform 1 0 5305 0 1 4313
box 0 0 64 64
use and3_dec  and3_dec_244
timestamp 1624494425
transform 1 0 6203 0 -1 4740
box 0 -60 2072 490
use and3_dec  and3_dec_245
timestamp 1624494425
transform 1 0 6203 0 1 3950
box 0 -60 2072 490
use contact_8  contact_8_1285
timestamp 1624494425
transform 1 0 4491 0 1 4588
box 0 0 64 64
use contact_7  contact_7_10
timestamp 1624494425
transform 1 0 4494 0 1 4587
box 0 0 58 66
use contact_16  contact_16_733
timestamp 1624494425
transform 1 0 5064 0 1 4518
box 0 0 66 58
use contact_16  contact_16_732
timestamp 1624494425
transform 1 0 5544 0 1 4428
box 0 0 66 58
use contact_9  contact_9_489
timestamp 1624494425
transform 1 0 6441 0 1 4331
box 0 0 66 74
use contact_8  contact_8_489
timestamp 1624494425
transform 1 0 6442 0 1 4336
box 0 0 64 64
use contact_9  contact_9_1243
timestamp 1624494425
transform 1 0 6866 0 1 4331
box 0 0 66 74
use contact_8  contact_8_1243
timestamp 1624494425
transform 1 0 6867 0 1 4336
box 0 0 64 64
use contact_9  contact_9_1244
timestamp 1624494425
transform 1 0 7298 0 1 4331
box 0 0 66 74
use contact_8  contact_8_1244
timestamp 1624494425
transform 1 0 7299 0 1 4336
box 0 0 64 64
use contact_16  contact_16_734
timestamp 1624494425
transform 1 0 4824 0 1 4630
box 0 0 66 58
use contact_16  contact_16_731
timestamp 1624494425
transform 1 0 4584 0 1 4792
box 0 0 66 58
use contact_8  contact_8_1284
timestamp 1624494425
transform 1 0 4491 0 1 4828
box 0 0 64 64
use contact_7  contact_7_9
timestamp 1624494425
transform 1 0 4494 0 1 4827
box 0 0 58 66
use contact_17  contact_17_9
timestamp 1624494425
transform 1 0 5385 0 1 4708
box 0 0 64 64
use contact_9  contact_9_487
timestamp 1624494425
transform 1 0 6441 0 1 4747
box 0 0 66 74
use contact_8  contact_8_487
timestamp 1624494425
transform 1 0 6442 0 1 4752
box 0 0 64 64
use contact_9  contact_9_1240
timestamp 1624494425
transform 1 0 6866 0 1 4689
box 0 0 66 74
use contact_8  contact_8_1240
timestamp 1624494425
transform 1 0 6867 0 1 4694
box 0 0 64 64
use contact_9  contact_9_1241
timestamp 1624494425
transform 1 0 7298 0 1 4689
box 0 0 66 74
use contact_8  contact_8_1241
timestamp 1624494425
transform 1 0 7299 0 1 4694
box 0 0 64 64
use and3_dec  and3_dec_243
timestamp 1624494425
transform 1 0 6203 0 1 4740
box 0 -60 2072 490
use contact_8  contact_8_1238
timestamp 1624494425
transform 1 0 7299 0 1 5126
box 0 0 64 64
use contact_9  contact_9_1238
timestamp 1624494425
transform 1 0 7298 0 1 5121
box 0 0 66 74
use contact_8  contact_8_1237
timestamp 1624494425
transform 1 0 6867 0 1 5126
box 0 0 64 64
use contact_9  contact_9_1237
timestamp 1624494425
transform 1 0 6866 0 1 5121
box 0 0 66 74
use contact_8  contact_8_485
timestamp 1624494425
transform 1 0 6442 0 1 5126
box 0 0 64 64
use contact_9  contact_9_485
timestamp 1624494425
transform 1 0 6441 0 1 5121
box 0 0 66 74
use contact_16  contact_16_729
timestamp 1624494425
transform 1 0 5544 0 1 4994
box 0 0 66 58
use contact_16  contact_16_730
timestamp 1624494425
transform 1 0 5144 0 1 4904
box 0 0 66 58
use contact_17  contact_17_8
timestamp 1624494425
transform 1 0 5465 0 1 5103
box 0 0 64 64
use contact_7  contact_7_8
timestamp 1624494425
transform 1 0 4494 0 1 5377
box 0 0 58 66
use contact_8  contact_8_1283
timestamp 1624494425
transform 1 0 4491 0 1 5378
box 0 0 64 64
use contact_16  contact_16_726
timestamp 1624494425
transform 1 0 5544 0 1 5218
box 0 0 66 58
use contact_16  contact_16_727
timestamp 1624494425
transform 1 0 5144 0 1 5308
box 0 0 66 58
use contact_16  contact_16_728
timestamp 1624494425
transform 1 0 4664 0 1 5420
box 0 0 66 58
use and3_dec  and3_dec_242
timestamp 1624494425
transform 1 0 6203 0 -1 5530
box 0 -60 2072 490
use contact_8  contact_8_1235
timestamp 1624494425
transform 1 0 7299 0 1 5484
box 0 0 64 64
use contact_9  contact_9_1235
timestamp 1624494425
transform 1 0 7298 0 1 5479
box 0 0 66 74
use contact_8  contact_8_1234
timestamp 1624494425
transform 1 0 6867 0 1 5484
box 0 0 64 64
use contact_9  contact_9_1234
timestamp 1624494425
transform 1 0 6866 0 1 5479
box 0 0 66 74
use contact_8  contact_8_483
timestamp 1624494425
transform 1 0 6442 0 1 5542
box 0 0 64 64
use contact_9  contact_9_483
timestamp 1624494425
transform 1 0 6441 0 1 5537
box 0 0 66 74
use contact_16  contact_16_724
timestamp 1624494425
transform 1 0 5144 0 1 5694
box 0 0 66 58
use contact_16  contact_16_725
timestamp 1624494425
transform 1 0 4744 0 1 5582
box 0 0 66 58
use contact_8  contact_8_1232
timestamp 1624494425
transform 1 0 7299 0 1 5916
box 0 0 64 64
use contact_9  contact_9_1232
timestamp 1624494425
transform 1 0 7298 0 1 5911
box 0 0 66 74
use contact_8  contact_8_1231
timestamp 1624494425
transform 1 0 6867 0 1 5916
box 0 0 64 64
use contact_9  contact_9_1231
timestamp 1624494425
transform 1 0 6866 0 1 5911
box 0 0 66 74
use contact_8  contact_8_481
timestamp 1624494425
transform 1 0 6442 0 1 5916
box 0 0 64 64
use contact_9  contact_9_481
timestamp 1624494425
transform 1 0 6441 0 1 5911
box 0 0 66 74
use contact_16  contact_16_723
timestamp 1624494425
transform 1 0 5544 0 1 5784
box 0 0 66 58
use and3_dec  and3_dec_240
timestamp 1624494425
transform 1 0 6203 0 -1 6320
box 0 -60 2072 490
use and3_dec  and3_dec_241
timestamp 1624494425
transform 1 0 6203 0 1 5530
box 0 -60 2072 490
use contact_16  contact_16_720
timestamp 1624494425
transform 1 0 5544 0 1 6008
box 0 0 66 58
use contact_16  contact_16_721
timestamp 1624494425
transform 1 0 5144 0 1 6098
box 0 0 66 58
use contact_16  contact_16_722
timestamp 1624494425
transform 1 0 4824 0 1 6210
box 0 0 66 58
use contact_16  contact_16_719
timestamp 1624494425
transform 1 0 4584 0 1 6372
box 0 0 66 58
use contact_8  contact_8_1282
timestamp 1624494425
transform 1 0 4491 0 1 6408
box 0 0 64 64
use contact_7  contact_7_7
timestamp 1624494425
transform 1 0 4494 0 1 6407
box 0 0 58 66
use contact_16  contact_16_718
timestamp 1624494425
transform 1 0 5224 0 1 6484
box 0 0 66 58
use contact_17  contact_17_7
timestamp 1624494425
transform 1 0 5545 0 1 6288
box 0 0 64 64
use contact_9  contact_9_479
timestamp 1624494425
transform 1 0 6441 0 1 6327
box 0 0 66 74
use contact_8  contact_8_479
timestamp 1624494425
transform 1 0 6442 0 1 6332
box 0 0 64 64
use contact_9  contact_9_1228
timestamp 1624494425
transform 1 0 6866 0 1 6269
box 0 0 66 74
use contact_8  contact_8_1228
timestamp 1624494425
transform 1 0 6867 0 1 6274
box 0 0 64 64
use contact_9  contact_9_1229
timestamp 1624494425
transform 1 0 7298 0 1 6269
box 0 0 66 74
use contact_8  contact_8_1229
timestamp 1624494425
transform 1 0 7299 0 1 6274
box 0 0 64 64
use and3_dec  and3_dec_239
timestamp 1624494425
transform 1 0 6203 0 1 6320
box 0 -60 2072 490
use contact_9  contact_9_492
timestamp 1624494425
transform 1 0 7680 0 1 3518
box 0 0 66 74
use contact_8  contact_8_492
timestamp 1624494425
transform 1 0 7681 0 1 3523
box 0 0 64 64
use contact_9  contact_9_1248
timestamp 1624494425
transform 1 0 8076 0 1 3518
box 0 0 66 74
use contact_8  contact_8_1248
timestamp 1624494425
transform 1 0 8077 0 1 3523
box 0 0 64 64
use contact_9  contact_9_488
timestamp 1624494425
transform 1 0 7680 0 1 4308
box 0 0 66 74
use contact_8  contact_8_488
timestamp 1624494425
transform 1 0 7681 0 1 4313
box 0 0 64 64
use contact_9  contact_9_490
timestamp 1624494425
transform 1 0 7680 0 1 3913
box 0 0 66 74
use contact_8  contact_8_490
timestamp 1624494425
transform 1 0 7681 0 1 3918
box 0 0 64 64
use contact_9  contact_9_1242
timestamp 1624494425
transform 1 0 8076 0 1 4308
box 0 0 66 74
use contact_8  contact_8_1242
timestamp 1624494425
transform 1 0 8077 0 1 4313
box 0 0 64 64
use contact_9  contact_9_1245
timestamp 1624494425
transform 1 0 8076 0 1 3913
box 0 0 66 74
use contact_8  contact_8_1245
timestamp 1624494425
transform 1 0 8077 0 1 3918
box 0 0 64 64
use contact_9  contact_9_486
timestamp 1624494425
transform 1 0 7680 0 1 4703
box 0 0 66 74
use contact_8  contact_8_486
timestamp 1624494425
transform 1 0 7681 0 1 4708
box 0 0 64 64
use contact_9  contact_9_1239
timestamp 1624494425
transform 1 0 8076 0 1 4703
box 0 0 66 74
use contact_8  contact_8_1239
timestamp 1624494425
transform 1 0 8077 0 1 4708
box 0 0 64 64
use contact_9  contact_9_482
timestamp 1624494425
transform 1 0 7680 0 1 5493
box 0 0 66 74
use contact_8  contact_8_482
timestamp 1624494425
transform 1 0 7681 0 1 5498
box 0 0 64 64
use contact_9  contact_9_484
timestamp 1624494425
transform 1 0 7680 0 1 5098
box 0 0 66 74
use contact_8  contact_8_484
timestamp 1624494425
transform 1 0 7681 0 1 5103
box 0 0 64 64
use contact_9  contact_9_1233
timestamp 1624494425
transform 1 0 8076 0 1 5493
box 0 0 66 74
use contact_8  contact_8_1233
timestamp 1624494425
transform 1 0 8077 0 1 5498
box 0 0 64 64
use contact_9  contact_9_1236
timestamp 1624494425
transform 1 0 8076 0 1 5098
box 0 0 66 74
use contact_8  contact_8_1236
timestamp 1624494425
transform 1 0 8077 0 1 5103
box 0 0 64 64
use contact_9  contact_9_478
timestamp 1624494425
transform 1 0 7680 0 1 6283
box 0 0 66 74
use contact_8  contact_8_478
timestamp 1624494425
transform 1 0 7681 0 1 6288
box 0 0 64 64
use contact_9  contact_9_480
timestamp 1624494425
transform 1 0 7680 0 1 5888
box 0 0 66 74
use contact_8  contact_8_480
timestamp 1624494425
transform 1 0 7681 0 1 5893
box 0 0 64 64
use contact_9  contact_9_1227
timestamp 1624494425
transform 1 0 8076 0 1 6283
box 0 0 66 74
use contact_8  contact_8_1227
timestamp 1624494425
transform 1 0 8077 0 1 6288
box 0 0 64 64
use contact_9  contact_9_1230
timestamp 1624494425
transform 1 0 8076 0 1 5888
box 0 0 66 74
use contact_8  contact_8_1230
timestamp 1624494425
transform 1 0 8077 0 1 5893
box 0 0 64 64
use contact_7  contact_7_21
timestamp 1624494425
transform 1 0 832 0 1 6907
box 0 0 58 66
use contact_7  contact_7_20
timestamp 1624494425
transform 1 0 912 0 1 7247
box 0 0 58 66
use contact_16  contact_16_768
timestamp 1624494425
transform 1 0 560 0 1 7251
box 0 0 66 58
use contact_16  contact_16_769
timestamp 1624494425
transform 1 0 480 0 1 6911
box 0 0 66 58
use contact_8  contact_8_1226
timestamp 1624494425
transform 1 0 7299 0 1 6706
box 0 0 64 64
use contact_9  contact_9_1226
timestamp 1624494425
transform 1 0 7298 0 1 6701
box 0 0 66 74
use contact_8  contact_8_1225
timestamp 1624494425
transform 1 0 6867 0 1 6706
box 0 0 64 64
use contact_9  contact_9_1225
timestamp 1624494425
transform 1 0 6866 0 1 6701
box 0 0 66 74
use contact_8  contact_8_477
timestamp 1624494425
transform 1 0 6442 0 1 6706
box 0 0 64 64
use contact_9  contact_9_477
timestamp 1624494425
transform 1 0 6441 0 1 6701
box 0 0 66 74
use contact_16  contact_16_717
timestamp 1624494425
transform 1 0 5544 0 1 6574
box 0 0 66 58
use contact_17  contact_17_6
timestamp 1624494425
transform 1 0 5625 0 1 6683
box 0 0 64 64
use contact_7  contact_7_6
timestamp 1624494425
transform 1 0 4494 0 1 6957
box 0 0 58 66
use contact_8  contact_8_1281
timestamp 1624494425
transform 1 0 4491 0 1 6958
box 0 0 64 64
use contact_16  contact_16_714
timestamp 1624494425
transform 1 0 5544 0 1 6798
box 0 0 66 58
use contact_16  contact_16_715
timestamp 1624494425
transform 1 0 5224 0 1 6888
box 0 0 66 58
use contact_16  contact_16_716
timestamp 1624494425
transform 1 0 4664 0 1 7000
box 0 0 66 58
use and3_dec  and3_dec_237
timestamp 1624494425
transform 1 0 6203 0 1 7110
box 0 -60 2072 490
use and3_dec  and3_dec_238
timestamp 1624494425
transform 1 0 6203 0 -1 7110
box 0 -60 2072 490
use contact_16  contact_16_713
timestamp 1624494425
transform 1 0 4744 0 1 7162
box 0 0 66 58
use contact_8  contact_8_1280
timestamp 1624494425
transform 1 0 4491 0 1 7198
box 0 0 64 64
use contact_7  contact_7_5
timestamp 1624494425
transform 1 0 4494 0 1 7197
box 0 0 58 66
use contact_16  contact_16_712
timestamp 1624494425
transform 1 0 5224 0 1 7274
box 0 0 66 58
use contact_17  contact_17_5
timestamp 1624494425
transform 1 0 5705 0 1 7078
box 0 0 64 64
use contact_9  contact_9_475
timestamp 1624494425
transform 1 0 6441 0 1 7117
box 0 0 66 74
use contact_8  contact_8_475
timestamp 1624494425
transform 1 0 6442 0 1 7122
box 0 0 64 64
use contact_9  contact_9_1222
timestamp 1624494425
transform 1 0 6866 0 1 7059
box 0 0 66 74
use contact_8  contact_8_1222
timestamp 1624494425
transform 1 0 6867 0 1 7064
box 0 0 64 64
use contact_9  contact_9_1223
timestamp 1624494425
transform 1 0 7298 0 1 7059
box 0 0 66 74
use contact_8  contact_8_1223
timestamp 1624494425
transform 1 0 7299 0 1 7064
box 0 0 64 64
use contact_8  contact_8_1220
timestamp 1624494425
transform 1 0 7299 0 1 7496
box 0 0 64 64
use contact_9  contact_9_1220
timestamp 1624494425
transform 1 0 7298 0 1 7491
box 0 0 66 74
use contact_8  contact_8_1219
timestamp 1624494425
transform 1 0 6867 0 1 7496
box 0 0 64 64
use contact_9  contact_9_1219
timestamp 1624494425
transform 1 0 6866 0 1 7491
box 0 0 66 74
use contact_8  contact_8_473
timestamp 1624494425
transform 1 0 6442 0 1 7496
box 0 0 64 64
use contact_9  contact_9_473
timestamp 1624494425
transform 1 0 6441 0 1 7491
box 0 0 66 74
use contact_16  contact_16_708
timestamp 1624494425
transform 1 0 5544 0 1 7588
box 0 0 66 58
use contact_16  contact_16_711
timestamp 1624494425
transform 1 0 5544 0 1 7364
box 0 0 66 58
use contact_17  contact_17_4
timestamp 1624494425
transform 1 0 5785 0 1 7473
box 0 0 64 64
use and3_dec  and3_dec_236
timestamp 1624494425
transform 1 0 6203 0 -1 7900
box 0 -60 2072 490
use contact_7  contact_7_4
timestamp 1624494425
transform 1 0 4494 0 1 7747
box 0 0 58 66
use contact_8  contact_8_1279
timestamp 1624494425
transform 1 0 4491 0 1 7748
box 0 0 64 64
use contact_8  contact_8_1217
timestamp 1624494425
transform 1 0 7299 0 1 7854
box 0 0 64 64
use contact_9  contact_9_1217
timestamp 1624494425
transform 1 0 7298 0 1 7849
box 0 0 66 74
use contact_8  contact_8_1216
timestamp 1624494425
transform 1 0 6867 0 1 7854
box 0 0 64 64
use contact_9  contact_9_1216
timestamp 1624494425
transform 1 0 6866 0 1 7849
box 0 0 66 74
use contact_16  contact_16_709
timestamp 1624494425
transform 1 0 5224 0 1 7678
box 0 0 66 58
use contact_16  contact_16_710
timestamp 1624494425
transform 1 0 4824 0 1 7790
box 0 0 66 58
use contact_17  contact_17_3
timestamp 1624494425
transform 1 0 5865 0 1 7868
box 0 0 64 64
use contact_7  contact_7_3
timestamp 1624494425
transform 1 0 4494 0 1 7987
box 0 0 58 66
use contact_8  contact_8_1278
timestamp 1624494425
transform 1 0 4491 0 1 7988
box 0 0 64 64
use contact_8  contact_8_471
timestamp 1624494425
transform 1 0 6442 0 1 7912
box 0 0 64 64
use contact_9  contact_9_471
timestamp 1624494425
transform 1 0 6441 0 1 7907
box 0 0 66 74
use contact_16  contact_16_705
timestamp 1624494425
transform 1 0 5544 0 1 8154
box 0 0 66 58
use contact_16  contact_16_706
timestamp 1624494425
transform 1 0 5304 0 1 8064
box 0 0 66 58
use contact_16  contact_16_707
timestamp 1624494425
transform 1 0 4584 0 1 7952
box 0 0 66 58
use and3_dec  and3_dec_235
timestamp 1624494425
transform 1 0 6203 0 1 7900
box 0 -60 2072 490
use contact_8  contact_8_1214
timestamp 1624494425
transform 1 0 7299 0 1 8286
box 0 0 64 64
use contact_9  contact_9_1214
timestamp 1624494425
transform 1 0 7298 0 1 8281
box 0 0 66 74
use contact_8  contact_8_1213
timestamp 1624494425
transform 1 0 6867 0 1 8286
box 0 0 64 64
use contact_9  contact_9_1213
timestamp 1624494425
transform 1 0 6866 0 1 8281
box 0 0 66 74
use contact_8  contact_8_469
timestamp 1624494425
transform 1 0 6442 0 1 8286
box 0 0 64 64
use contact_9  contact_9_469
timestamp 1624494425
transform 1 0 6441 0 1 8281
box 0 0 66 74
use contact_16  contact_16_702
timestamp 1624494425
transform 1 0 5544 0 1 8378
box 0 0 66 58
use contact_17  contact_17_2
timestamp 1624494425
transform 1 0 5945 0 1 8263
box 0 0 64 64
use contact_16  contact_16_704
timestamp 1624494425
transform 1 0 4664 0 1 8580
box 0 0 66 58
use contact_8  contact_8_1277
timestamp 1624494425
transform 1 0 4491 0 1 8538
box 0 0 64 64
use contact_7  contact_7_2
timestamp 1624494425
transform 1 0 4494 0 1 8537
box 0 0 58 66
use contact_16  contact_16_703
timestamp 1624494425
transform 1 0 5304 0 1 8468
box 0 0 66 58
use contact_17  contact_17_1
timestamp 1624494425
transform 1 0 6025 0 1 8658
box 0 0 64 64
use contact_9  contact_9_467
timestamp 1624494425
transform 1 0 6441 0 1 8697
box 0 0 66 74
use contact_8  contact_8_467
timestamp 1624494425
transform 1 0 6442 0 1 8702
box 0 0 64 64
use contact_9  contact_9_1210
timestamp 1624494425
transform 1 0 6866 0 1 8639
box 0 0 66 74
use contact_8  contact_8_1210
timestamp 1624494425
transform 1 0 6867 0 1 8644
box 0 0 64 64
use contact_9  contact_9_1211
timestamp 1624494425
transform 1 0 7298 0 1 8639
box 0 0 66 74
use contact_8  contact_8_1211
timestamp 1624494425
transform 1 0 7299 0 1 8644
box 0 0 64 64
use and3_dec  and3_dec_233
timestamp 1624494425
transform 1 0 6203 0 1 8690
box 0 -60 2072 490
use and3_dec  and3_dec_234
timestamp 1624494425
transform 1 0 6203 0 -1 8690
box 0 -60 2072 490
use contact_7  contact_7_1
timestamp 1624494425
transform 1 0 4494 0 1 8777
box 0 0 58 66
use contact_8  contact_8_1276
timestamp 1624494425
transform 1 0 4491 0 1 8778
box 0 0 64 64
use contact_16  contact_16_699
timestamp 1624494425
transform 1 0 5544 0 1 8944
box 0 0 66 58
use contact_16  contact_16_700
timestamp 1624494425
transform 1 0 5304 0 1 8854
box 0 0 66 58
use contact_16  contact_16_701
timestamp 1624494425
transform 1 0 4744 0 1 8742
box 0 0 66 58
use contact_8  contact_8_1208
timestamp 1624494425
transform 1 0 7299 0 1 9076
box 0 0 64 64
use contact_9  contact_9_1208
timestamp 1624494425
transform 1 0 7298 0 1 9071
box 0 0 66 74
use contact_8  contact_8_1207
timestamp 1624494425
transform 1 0 6867 0 1 9076
box 0 0 64 64
use contact_9  contact_9_1207
timestamp 1624494425
transform 1 0 6866 0 1 9071
box 0 0 66 74
use contact_8  contact_8_465
timestamp 1624494425
transform 1 0 6442 0 1 9076
box 0 0 64 64
use contact_9  contact_9_465
timestamp 1624494425
transform 1 0 6441 0 1 9071
box 0 0 66 74
use contact_16  contact_16_696
timestamp 1624494425
transform 1 0 5544 0 1 9168
box 0 0 66 58
use contact_17  contact_17_0
timestamp 1624494425
transform 1 0 6105 0 1 9053
box 0 0 64 64
use and3_dec  and3_dec_232
timestamp 1624494425
transform 1 0 6203 0 -1 9480
box 0 -60 2072 490
use contact_16  contact_16_698
timestamp 1624494425
transform 1 0 4824 0 1 9370
box 0 0 66 58
use contact_16  contact_16_695
timestamp 1624494425
transform 1 0 4584 0 1 9532
box 0 0 66 58
use contact_8  contact_8_1275
timestamp 1624494425
transform 1 0 4491 0 1 9328
box 0 0 64 64
use contact_7  contact_7_0
timestamp 1624494425
transform 1 0 4494 0 1 9327
box 0 0 58 66
use contact_16  contact_16_697
timestamp 1624494425
transform 1 0 5304 0 1 9258
box 0 0 66 58
use contact_9  contact_9_463
timestamp 1624494425
transform 1 0 6441 0 1 9487
box 0 0 66 74
use contact_8  contact_8_463
timestamp 1624494425
transform 1 0 6442 0 1 9492
box 0 0 64 64
use contact_9  contact_9_1204
timestamp 1624494425
transform 1 0 6866 0 1 9429
box 0 0 66 74
use contact_8  contact_8_1204
timestamp 1624494425
transform 1 0 6867 0 1 9434
box 0 0 64 64
use contact_9  contact_9_1205
timestamp 1624494425
transform 1 0 7298 0 1 9429
box 0 0 66 74
use contact_8  contact_8_1205
timestamp 1624494425
transform 1 0 7299 0 1 9434
box 0 0 64 64
use contact_16  contact_16_693
timestamp 1624494425
transform 1 0 5544 0 1 9734
box 0 0 66 58
use contact_16  contact_16_694
timestamp 1624494425
transform 1 0 5384 0 1 9644
box 0 0 66 58
use and3_dec  and3_dec_230
timestamp 1624494425
transform 1 0 6203 0 -1 10270
box 0 -60 2072 490
use and3_dec  and3_dec_231
timestamp 1624494425
transform 1 0 6203 0 1 9480
box 0 -60 2072 490
use contact_9  contact_9_474
timestamp 1624494425
transform 1 0 7680 0 1 7073
box 0 0 66 74
use contact_8  contact_8_474
timestamp 1624494425
transform 1 0 7681 0 1 7078
box 0 0 64 64
use contact_9  contact_9_476
timestamp 1624494425
transform 1 0 7680 0 1 6678
box 0 0 66 74
use contact_8  contact_8_476
timestamp 1624494425
transform 1 0 7681 0 1 6683
box 0 0 64 64
use contact_9  contact_9_1221
timestamp 1624494425
transform 1 0 8076 0 1 7073
box 0 0 66 74
use contact_8  contact_8_1221
timestamp 1624494425
transform 1 0 8077 0 1 7078
box 0 0 64 64
use contact_9  contact_9_1224
timestamp 1624494425
transform 1 0 8076 0 1 6678
box 0 0 66 74
use contact_8  contact_8_1224
timestamp 1624494425
transform 1 0 8077 0 1 6683
box 0 0 64 64
use contact_9  contact_9_472
timestamp 1624494425
transform 1 0 7680 0 1 7468
box 0 0 66 74
use contact_8  contact_8_472
timestamp 1624494425
transform 1 0 7681 0 1 7473
box 0 0 64 64
use contact_9  contact_9_1218
timestamp 1624494425
transform 1 0 8076 0 1 7468
box 0 0 66 74
use contact_8  contact_8_1218
timestamp 1624494425
transform 1 0 8077 0 1 7473
box 0 0 64 64
use contact_9  contact_9_468
timestamp 1624494425
transform 1 0 7680 0 1 8258
box 0 0 66 74
use contact_8  contact_8_468
timestamp 1624494425
transform 1 0 7681 0 1 8263
box 0 0 64 64
use contact_9  contact_9_470
timestamp 1624494425
transform 1 0 7680 0 1 7863
box 0 0 66 74
use contact_8  contact_8_470
timestamp 1624494425
transform 1 0 7681 0 1 7868
box 0 0 64 64
use contact_9  contact_9_1212
timestamp 1624494425
transform 1 0 8076 0 1 8258
box 0 0 66 74
use contact_8  contact_8_1212
timestamp 1624494425
transform 1 0 8077 0 1 8263
box 0 0 64 64
use contact_9  contact_9_1215
timestamp 1624494425
transform 1 0 8076 0 1 7863
box 0 0 66 74
use contact_8  contact_8_1215
timestamp 1624494425
transform 1 0 8077 0 1 7868
box 0 0 64 64
use contact_9  contact_9_466
timestamp 1624494425
transform 1 0 7680 0 1 8653
box 0 0 66 74
use contact_8  contact_8_466
timestamp 1624494425
transform 1 0 7681 0 1 8658
box 0 0 64 64
use contact_9  contact_9_1209
timestamp 1624494425
transform 1 0 8076 0 1 8653
box 0 0 66 74
use contact_8  contact_8_1209
timestamp 1624494425
transform 1 0 8077 0 1 8658
box 0 0 64 64
use contact_9  contact_9_462
timestamp 1624494425
transform 1 0 7680 0 1 9443
box 0 0 66 74
use contact_8  contact_8_462
timestamp 1624494425
transform 1 0 7681 0 1 9448
box 0 0 64 64
use contact_9  contact_9_464
timestamp 1624494425
transform 1 0 7680 0 1 9048
box 0 0 66 74
use contact_8  contact_8_464
timestamp 1624494425
transform 1 0 7681 0 1 9053
box 0 0 64 64
use contact_9  contact_9_1203
timestamp 1624494425
transform 1 0 8076 0 1 9443
box 0 0 66 74
use contact_8  contact_8_1203
timestamp 1624494425
transform 1 0 8077 0 1 9448
box 0 0 64 64
use contact_9  contact_9_1206
timestamp 1624494425
transform 1 0 8076 0 1 9048
box 0 0 66 74
use contact_8  contact_8_1206
timestamp 1624494425
transform 1 0 8077 0 1 9053
box 0 0 64 64
use contact_8  contact_8_1202
timestamp 1624494425
transform 1 0 7299 0 1 9866
box 0 0 64 64
use contact_9  contact_9_1202
timestamp 1624494425
transform 1 0 7298 0 1 9861
box 0 0 66 74
use contact_8  contact_8_1201
timestamp 1624494425
transform 1 0 6867 0 1 9866
box 0 0 64 64
use contact_9  contact_9_1201
timestamp 1624494425
transform 1 0 6866 0 1 9861
box 0 0 66 74
use contact_8  contact_8_461
timestamp 1624494425
transform 1 0 6442 0 1 9866
box 0 0 64 64
use contact_9  contact_9_461
timestamp 1624494425
transform 1 0 6441 0 1 9861
box 0 0 66 74
use contact_16  contact_16_690
timestamp 1624494425
transform 1 0 5544 0 1 9958
box 0 0 66 58
use contact_16  contact_16_691
timestamp 1624494425
transform 1 0 5384 0 1 10048
box 0 0 66 58
use contact_8  contact_8_1199
timestamp 1624494425
transform 1 0 7299 0 1 10224
box 0 0 64 64
use contact_9  contact_9_1199
timestamp 1624494425
transform 1 0 7298 0 1 10219
box 0 0 66 74
use contact_8  contact_8_1198
timestamp 1624494425
transform 1 0 6867 0 1 10224
box 0 0 64 64
use contact_9  contact_9_1198
timestamp 1624494425
transform 1 0 6866 0 1 10219
box 0 0 66 74
use contact_8  contact_8_459
timestamp 1624494425
transform 1 0 6442 0 1 10282
box 0 0 64 64
use contact_9  contact_9_459
timestamp 1624494425
transform 1 0 6441 0 1 10277
box 0 0 66 74
use contact_16  contact_16_689
timestamp 1624494425
transform 1 0 4744 0 1 10322
box 0 0 66 58
use contact_16  contact_16_692
timestamp 1624494425
transform 1 0 4664 0 1 10160
box 0 0 66 58
use and3_dec  and3_dec_229
timestamp 1624494425
transform 1 0 6203 0 1 10270
box 0 -60 2072 490
use contact_16  contact_16_687
timestamp 1624494425
transform 1 0 5544 0 1 10524
box 0 0 66 58
use contact_16  contact_16_688
timestamp 1624494425
transform 1 0 5384 0 1 10434
box 0 0 66 58
use contact_8  contact_8_1196
timestamp 1624494425
transform 1 0 7299 0 1 10656
box 0 0 64 64
use contact_9  contact_9_1196
timestamp 1624494425
transform 1 0 7298 0 1 10651
box 0 0 66 74
use contact_8  contact_8_1195
timestamp 1624494425
transform 1 0 6867 0 1 10656
box 0 0 64 64
use contact_9  contact_9_1195
timestamp 1624494425
transform 1 0 6866 0 1 10651
box 0 0 66 74
use contact_8  contact_8_457
timestamp 1624494425
transform 1 0 6442 0 1 10656
box 0 0 64 64
use contact_9  contact_9_457
timestamp 1624494425
transform 1 0 6441 0 1 10651
box 0 0 66 74
use contact_16  contact_16_684
timestamp 1624494425
transform 1 0 5544 0 1 10748
box 0 0 66 58
use contact_16  contact_16_685
timestamp 1624494425
transform 1 0 5384 0 1 10838
box 0 0 66 58
use and3_dec  and3_dec_228
timestamp 1624494425
transform 1 0 6203 0 -1 11060
box 0 -60 2072 490
use contact_8  contact_8_1193
timestamp 1624494425
transform 1 0 7299 0 1 11014
box 0 0 64 64
use contact_9  contact_9_1193
timestamp 1624494425
transform 1 0 7298 0 1 11009
box 0 0 66 74
use contact_8  contact_8_1192
timestamp 1624494425
transform 1 0 6867 0 1 11014
box 0 0 64 64
use contact_9  contact_9_1192
timestamp 1624494425
transform 1 0 6866 0 1 11009
box 0 0 66 74
use contact_8  contact_8_455
timestamp 1624494425
transform 1 0 6442 0 1 11072
box 0 0 64 64
use contact_9  contact_9_455
timestamp 1624494425
transform 1 0 6441 0 1 11067
box 0 0 66 74
use contact_16  contact_16_683
timestamp 1624494425
transform 1 0 4584 0 1 11112
box 0 0 66 58
use contact_16  contact_16_686
timestamp 1624494425
transform 1 0 4824 0 1 10950
box 0 0 66 58
use contact_16  contact_16_681
timestamp 1624494425
transform 1 0 5544 0 1 11314
box 0 0 66 58
use contact_16  contact_16_682
timestamp 1624494425
transform 1 0 5464 0 1 11224
box 0 0 66 58
use and3_dec  and3_dec_226
timestamp 1624494425
transform 1 0 6203 0 -1 11850
box 0 -60 2072 490
use and3_dec  and3_dec_227
timestamp 1624494425
transform 1 0 6203 0 1 11060
box 0 -60 2072 490
use contact_8  contact_8_1190
timestamp 1624494425
transform 1 0 7299 0 1 11446
box 0 0 64 64
use contact_9  contact_9_1190
timestamp 1624494425
transform 1 0 7298 0 1 11441
box 0 0 66 74
use contact_8  contact_8_1189
timestamp 1624494425
transform 1 0 6867 0 1 11446
box 0 0 64 64
use contact_9  contact_9_1189
timestamp 1624494425
transform 1 0 6866 0 1 11441
box 0 0 66 74
use contact_8  contact_8_453
timestamp 1624494425
transform 1 0 6442 0 1 11446
box 0 0 64 64
use contact_9  contact_9_453
timestamp 1624494425
transform 1 0 6441 0 1 11441
box 0 0 66 74
use contact_16  contact_16_678
timestamp 1624494425
transform 1 0 5544 0 1 11538
box 0 0 66 58
use contact_16  contact_16_679
timestamp 1624494425
transform 1 0 5464 0 1 11628
box 0 0 66 58
use contact_8  contact_8_1187
timestamp 1624494425
transform 1 0 7299 0 1 11804
box 0 0 64 64
use contact_9  contact_9_1187
timestamp 1624494425
transform 1 0 7298 0 1 11799
box 0 0 66 74
use contact_8  contact_8_1186
timestamp 1624494425
transform 1 0 6867 0 1 11804
box 0 0 64 64
use contact_9  contact_9_1186
timestamp 1624494425
transform 1 0 6866 0 1 11799
box 0 0 66 74
use contact_8  contact_8_451
timestamp 1624494425
transform 1 0 6442 0 1 11862
box 0 0 64 64
use contact_9  contact_9_451
timestamp 1624494425
transform 1 0 6441 0 1 11857
box 0 0 66 74
use contact_16  contact_16_677
timestamp 1624494425
transform 1 0 4744 0 1 11902
box 0 0 66 58
use contact_16  contact_16_680
timestamp 1624494425
transform 1 0 4664 0 1 11740
box 0 0 66 58
use and3_dec  and3_dec_225
timestamp 1624494425
transform 1 0 6203 0 1 11850
box 0 -60 2072 490
use contact_8  contact_8_1184
timestamp 1624494425
transform 1 0 7299 0 1 12236
box 0 0 64 64
use contact_9  contact_9_1184
timestamp 1624494425
transform 1 0 7298 0 1 12231
box 0 0 66 74
use contact_8  contact_8_1183
timestamp 1624494425
transform 1 0 6867 0 1 12236
box 0 0 64 64
use contact_9  contact_9_1183
timestamp 1624494425
transform 1 0 6866 0 1 12231
box 0 0 66 74
use contact_8  contact_8_449
timestamp 1624494425
transform 1 0 6442 0 1 12236
box 0 0 64 64
use contact_9  contact_9_449
timestamp 1624494425
transform 1 0 6441 0 1 12231
box 0 0 66 74
use contact_16  contact_16_675
timestamp 1624494425
transform 1 0 5544 0 1 12104
box 0 0 66 58
use contact_16  contact_16_676
timestamp 1624494425
transform 1 0 5464 0 1 12014
box 0 0 66 58
use contact_16  contact_16_672
timestamp 1624494425
transform 1 0 5544 0 1 12328
box 0 0 66 58
use contact_16  contact_16_673
timestamp 1624494425
transform 1 0 5464 0 1 12418
box 0 0 66 58
use contact_16  contact_16_674
timestamp 1624494425
transform 1 0 4824 0 1 12530
box 0 0 66 58
use and3_dec  and3_dec_224
timestamp 1624494425
transform 1 0 6203 0 -1 12640
box 0 -60 2072 490
use contact_8  contact_8_1181
timestamp 1624494425
transform 1 0 7299 0 1 12594
box 0 0 64 64
use contact_9  contact_9_1181
timestamp 1624494425
transform 1 0 7298 0 1 12589
box 0 0 66 74
use contact_8  contact_8_1180
timestamp 1624494425
transform 1 0 6867 0 1 12594
box 0 0 64 64
use contact_9  contact_9_1180
timestamp 1624494425
transform 1 0 6866 0 1 12589
box 0 0 66 74
use contact_8  contact_8_447
timestamp 1624494425
transform 1 0 6442 0 1 12652
box 0 0 64 64
use contact_9  contact_9_447
timestamp 1624494425
transform 1 0 6441 0 1 12647
box 0 0 66 74
use contact_16  contact_16_670
timestamp 1624494425
transform 1 0 4904 0 1 12804
box 0 0 66 58
use contact_16  contact_16_671
timestamp 1624494425
transform 1 0 4584 0 1 12692
box 0 0 66 58
use contact_8  contact_8_1178
timestamp 1624494425
transform 1 0 7299 0 1 13026
box 0 0 64 64
use contact_9  contact_9_1178
timestamp 1624494425
transform 1 0 7298 0 1 13021
box 0 0 66 74
use contact_8  contact_8_1177
timestamp 1624494425
transform 1 0 6867 0 1 13026
box 0 0 64 64
use contact_9  contact_9_1177
timestamp 1624494425
transform 1 0 6866 0 1 13021
box 0 0 66 74
use contact_8  contact_8_445
timestamp 1624494425
transform 1 0 6442 0 1 13026
box 0 0 64 64
use contact_9  contact_9_445
timestamp 1624494425
transform 1 0 6441 0 1 13021
box 0 0 66 74
use contact_16  contact_16_669
timestamp 1624494425
transform 1 0 5624 0 1 12894
box 0 0 66 58
use and3_dec  and3_dec_222
timestamp 1624494425
transform 1 0 6203 0 -1 13430
box 0 -60 2072 490
use and3_dec  and3_dec_223
timestamp 1624494425
transform 1 0 6203 0 1 12640
box 0 -60 2072 490
use contact_9  contact_9_458
timestamp 1624494425
transform 1 0 7680 0 1 10233
box 0 0 66 74
use contact_8  contact_8_458
timestamp 1624494425
transform 1 0 7681 0 1 10238
box 0 0 64 64
use contact_9  contact_9_460
timestamp 1624494425
transform 1 0 7680 0 1 9838
box 0 0 66 74
use contact_8  contact_8_460
timestamp 1624494425
transform 1 0 7681 0 1 9843
box 0 0 64 64
use contact_9  contact_9_1197
timestamp 1624494425
transform 1 0 8076 0 1 10233
box 0 0 66 74
use contact_8  contact_8_1197
timestamp 1624494425
transform 1 0 8077 0 1 10238
box 0 0 64 64
use contact_9  contact_9_1200
timestamp 1624494425
transform 1 0 8076 0 1 9838
box 0 0 66 74
use contact_8  contact_8_1200
timestamp 1624494425
transform 1 0 8077 0 1 9843
box 0 0 64 64
use contact_9  contact_9_456
timestamp 1624494425
transform 1 0 7680 0 1 10628
box 0 0 66 74
use contact_8  contact_8_456
timestamp 1624494425
transform 1 0 7681 0 1 10633
box 0 0 64 64
use contact_9  contact_9_1194
timestamp 1624494425
transform 1 0 8076 0 1 10628
box 0 0 66 74
use contact_8  contact_8_1194
timestamp 1624494425
transform 1 0 8077 0 1 10633
box 0 0 64 64
use contact_9  contact_9_452
timestamp 1624494425
transform 1 0 7680 0 1 11418
box 0 0 66 74
use contact_8  contact_8_452
timestamp 1624494425
transform 1 0 7681 0 1 11423
box 0 0 64 64
use contact_9  contact_9_454
timestamp 1624494425
transform 1 0 7680 0 1 11023
box 0 0 66 74
use contact_8  contact_8_454
timestamp 1624494425
transform 1 0 7681 0 1 11028
box 0 0 64 64
use contact_9  contact_9_1188
timestamp 1624494425
transform 1 0 8076 0 1 11418
box 0 0 66 74
use contact_8  contact_8_1188
timestamp 1624494425
transform 1 0 8077 0 1 11423
box 0 0 64 64
use contact_9  contact_9_1191
timestamp 1624494425
transform 1 0 8076 0 1 11023
box 0 0 66 74
use contact_8  contact_8_1191
timestamp 1624494425
transform 1 0 8077 0 1 11028
box 0 0 64 64
use contact_9  contact_9_450
timestamp 1624494425
transform 1 0 7680 0 1 11813
box 0 0 66 74
use contact_8  contact_8_450
timestamp 1624494425
transform 1 0 7681 0 1 11818
box 0 0 64 64
use contact_9  contact_9_1185
timestamp 1624494425
transform 1 0 8076 0 1 11813
box 0 0 66 74
use contact_8  contact_8_1185
timestamp 1624494425
transform 1 0 8077 0 1 11818
box 0 0 64 64
use contact_9  contact_9_446
timestamp 1624494425
transform 1 0 7680 0 1 12603
box 0 0 66 74
use contact_8  contact_8_446
timestamp 1624494425
transform 1 0 7681 0 1 12608
box 0 0 64 64
use contact_9  contact_9_448
timestamp 1624494425
transform 1 0 7680 0 1 12208
box 0 0 66 74
use contact_8  contact_8_448
timestamp 1624494425
transform 1 0 7681 0 1 12213
box 0 0 64 64
use contact_9  contact_9_1179
timestamp 1624494425
transform 1 0 8076 0 1 12603
box 0 0 66 74
use contact_8  contact_8_1179
timestamp 1624494425
transform 1 0 8077 0 1 12608
box 0 0 64 64
use contact_9  contact_9_1182
timestamp 1624494425
transform 1 0 8076 0 1 12208
box 0 0 66 74
use contact_8  contact_8_1182
timestamp 1624494425
transform 1 0 8077 0 1 12213
box 0 0 64 64
use contact_9  contact_9_444
timestamp 1624494425
transform 1 0 7680 0 1 12998
box 0 0 66 74
use contact_8  contact_8_444
timestamp 1624494425
transform 1 0 7681 0 1 13003
box 0 0 64 64
use contact_9  contact_9_1176
timestamp 1624494425
transform 1 0 8076 0 1 12998
box 0 0 66 74
use contact_8  contact_8_1176
timestamp 1624494425
transform 1 0 8077 0 1 13003
box 0 0 64 64
use contact_16  contact_16_666
timestamp 1624494425
transform 1 0 5624 0 1 13118
box 0 0 66 58
use contact_16  contact_16_667
timestamp 1624494425
transform 1 0 4904 0 1 13208
box 0 0 66 58
use contact_16  contact_16_668
timestamp 1624494425
transform 1 0 4664 0 1 13320
box 0 0 66 58
use contact_8  contact_8_1175
timestamp 1624494425
transform 1 0 7299 0 1 13384
box 0 0 64 64
use contact_9  contact_9_1175
timestamp 1624494425
transform 1 0 7298 0 1 13379
box 0 0 66 74
use contact_8  contact_8_1174
timestamp 1624494425
transform 1 0 6867 0 1 13384
box 0 0 64 64
use contact_9  contact_9_1174
timestamp 1624494425
transform 1 0 6866 0 1 13379
box 0 0 66 74
use contact_8  contact_8_443
timestamp 1624494425
transform 1 0 6442 0 1 13442
box 0 0 64 64
use contact_9  contact_9_443
timestamp 1624494425
transform 1 0 6441 0 1 13437
box 0 0 66 74
use contact_16  contact_16_664
timestamp 1624494425
transform 1 0 4904 0 1 13594
box 0 0 66 58
use contact_16  contact_16_665
timestamp 1624494425
transform 1 0 4744 0 1 13482
box 0 0 66 58
use and3_dec  and3_dec_221
timestamp 1624494425
transform 1 0 6203 0 1 13430
box 0 -60 2072 490
use contact_8  contact_8_1172
timestamp 1624494425
transform 1 0 7299 0 1 13816
box 0 0 64 64
use contact_9  contact_9_1172
timestamp 1624494425
transform 1 0 7298 0 1 13811
box 0 0 66 74
use contact_8  contact_8_1171
timestamp 1624494425
transform 1 0 6867 0 1 13816
box 0 0 64 64
use contact_9  contact_9_1171
timestamp 1624494425
transform 1 0 6866 0 1 13811
box 0 0 66 74
use contact_8  contact_8_441
timestamp 1624494425
transform 1 0 6442 0 1 13816
box 0 0 64 64
use contact_9  contact_9_441
timestamp 1624494425
transform 1 0 6441 0 1 13811
box 0 0 66 74
use contact_16  contact_16_663
timestamp 1624494425
transform 1 0 5624 0 1 13684
box 0 0 66 58
use contact_16  contact_16_660
timestamp 1624494425
transform 1 0 5624 0 1 13908
box 0 0 66 58
use contact_16  contact_16_661
timestamp 1624494425
transform 1 0 4904 0 1 13998
box 0 0 66 58
use contact_16  contact_16_662
timestamp 1624494425
transform 1 0 4824 0 1 14110
box 0 0 66 58
use and3_dec  and3_dec_219
timestamp 1624494425
transform 1 0 6203 0 1 14220
box 0 -60 2072 490
use and3_dec  and3_dec_220
timestamp 1624494425
transform 1 0 6203 0 -1 14220
box 0 -60 2072 490
use contact_8  contact_8_1169
timestamp 1624494425
transform 1 0 7299 0 1 14174
box 0 0 64 64
use contact_9  contact_9_1169
timestamp 1624494425
transform 1 0 7298 0 1 14169
box 0 0 66 74
use contact_8  contact_8_1168
timestamp 1624494425
transform 1 0 6867 0 1 14174
box 0 0 64 64
use contact_9  contact_9_1168
timestamp 1624494425
transform 1 0 6866 0 1 14169
box 0 0 66 74
use contact_8  contact_8_439
timestamp 1624494425
transform 1 0 6442 0 1 14232
box 0 0 64 64
use contact_9  contact_9_439
timestamp 1624494425
transform 1 0 6441 0 1 14227
box 0 0 66 74
use contact_16  contact_16_658
timestamp 1624494425
transform 1 0 4984 0 1 14384
box 0 0 66 58
use contact_16  contact_16_659
timestamp 1624494425
transform 1 0 4584 0 1 14272
box 0 0 66 58
use contact_8  contact_8_1166
timestamp 1624494425
transform 1 0 7299 0 1 14606
box 0 0 64 64
use contact_9  contact_9_1166
timestamp 1624494425
transform 1 0 7298 0 1 14601
box 0 0 66 74
use contact_8  contact_8_1165
timestamp 1624494425
transform 1 0 6867 0 1 14606
box 0 0 64 64
use contact_9  contact_9_1165
timestamp 1624494425
transform 1 0 6866 0 1 14601
box 0 0 66 74
use contact_8  contact_8_437
timestamp 1624494425
transform 1 0 6442 0 1 14606
box 0 0 64 64
use contact_9  contact_9_437
timestamp 1624494425
transform 1 0 6441 0 1 14601
box 0 0 66 74
use contact_16  contact_16_654
timestamp 1624494425
transform 1 0 5624 0 1 14698
box 0 0 66 58
use contact_16  contact_16_657
timestamp 1624494425
transform 1 0 5624 0 1 14474
box 0 0 66 58
use and3_dec  and3_dec_218
timestamp 1624494425
transform 1 0 6203 0 -1 15010
box 0 -60 2072 490
use contact_8  contact_8_1163
timestamp 1624494425
transform 1 0 7299 0 1 14964
box 0 0 64 64
use contact_9  contact_9_1163
timestamp 1624494425
transform 1 0 7298 0 1 14959
box 0 0 66 74
use contact_8  contact_8_1162
timestamp 1624494425
transform 1 0 6867 0 1 14964
box 0 0 64 64
use contact_9  contact_9_1162
timestamp 1624494425
transform 1 0 6866 0 1 14959
box 0 0 66 74
use contact_16  contact_16_655
timestamp 1624494425
transform 1 0 4984 0 1 14788
box 0 0 66 58
use contact_16  contact_16_656
timestamp 1624494425
transform 1 0 4664 0 1 14900
box 0 0 66 58
use contact_8  contact_8_435
timestamp 1624494425
transform 1 0 6442 0 1 15022
box 0 0 64 64
use contact_9  contact_9_435
timestamp 1624494425
transform 1 0 6441 0 1 15017
box 0 0 66 74
use contact_16  contact_16_651
timestamp 1624494425
transform 1 0 5624 0 1 15264
box 0 0 66 58
use contact_16  contact_16_652
timestamp 1624494425
transform 1 0 4984 0 1 15174
box 0 0 66 58
use contact_16  contact_16_653
timestamp 1624494425
transform 1 0 4744 0 1 15062
box 0 0 66 58
use and3_dec  and3_dec_217
timestamp 1624494425
transform 1 0 6203 0 1 15010
box 0 -60 2072 490
use contact_8  contact_8_1160
timestamp 1624494425
transform 1 0 7299 0 1 15396
box 0 0 64 64
use contact_9  contact_9_1160
timestamp 1624494425
transform 1 0 7298 0 1 15391
box 0 0 66 74
use contact_8  contact_8_1159
timestamp 1624494425
transform 1 0 6867 0 1 15396
box 0 0 64 64
use contact_9  contact_9_1159
timestamp 1624494425
transform 1 0 6866 0 1 15391
box 0 0 66 74
use contact_8  contact_8_433
timestamp 1624494425
transform 1 0 6442 0 1 15396
box 0 0 64 64
use contact_9  contact_9_433
timestamp 1624494425
transform 1 0 6441 0 1 15391
box 0 0 66 74
use contact_16  contact_16_648
timestamp 1624494425
transform 1 0 5624 0 1 15488
box 0 0 66 58
use contact_8  contact_8_1157
timestamp 1624494425
transform 1 0 7299 0 1 15754
box 0 0 64 64
use contact_9  contact_9_1157
timestamp 1624494425
transform 1 0 7298 0 1 15749
box 0 0 66 74
use contact_8  contact_8_1156
timestamp 1624494425
transform 1 0 6867 0 1 15754
box 0 0 64 64
use contact_9  contact_9_1156
timestamp 1624494425
transform 1 0 6866 0 1 15749
box 0 0 66 74
use contact_8  contact_8_431
timestamp 1624494425
transform 1 0 6442 0 1 15812
box 0 0 64 64
use contact_9  contact_9_431
timestamp 1624494425
transform 1 0 6441 0 1 15807
box 0 0 66 74
use contact_16  contact_16_649
timestamp 1624494425
transform 1 0 4984 0 1 15578
box 0 0 66 58
use contact_16  contact_16_650
timestamp 1624494425
transform 1 0 4824 0 1 15690
box 0 0 66 58
use and3_dec  and3_dec_215
timestamp 1624494425
transform 1 0 6203 0 1 15800
box 0 -60 2072 490
use and3_dec  and3_dec_216
timestamp 1624494425
transform 1 0 6203 0 -1 15800
box 0 -60 2072 490
use contact_16  contact_16_645
timestamp 1624494425
transform 1 0 5624 0 1 16054
box 0 0 66 58
use contact_16  contact_16_646
timestamp 1624494425
transform 1 0 5064 0 1 15964
box 0 0 66 58
use contact_16  contact_16_647
timestamp 1624494425
transform 1 0 4584 0 1 15852
box 0 0 66 58
use contact_8  contact_8_1154
timestamp 1624494425
transform 1 0 7299 0 1 16186
box 0 0 64 64
use contact_9  contact_9_1154
timestamp 1624494425
transform 1 0 7298 0 1 16181
box 0 0 66 74
use contact_8  contact_8_1153
timestamp 1624494425
transform 1 0 6867 0 1 16186
box 0 0 64 64
use contact_9  contact_9_1153
timestamp 1624494425
transform 1 0 6866 0 1 16181
box 0 0 66 74
use contact_8  contact_8_429
timestamp 1624494425
transform 1 0 6442 0 1 16186
box 0 0 64 64
use contact_9  contact_9_429
timestamp 1624494425
transform 1 0 6441 0 1 16181
box 0 0 66 74
use contact_16  contact_16_642
timestamp 1624494425
transform 1 0 5624 0 1 16278
box 0 0 66 58
use and3_dec  and3_dec_214
timestamp 1624494425
transform 1 0 6203 0 -1 16590
box 0 -60 2072 490
use contact_9  contact_9_442
timestamp 1624494425
transform 1 0 7680 0 1 13393
box 0 0 66 74
use contact_8  contact_8_442
timestamp 1624494425
transform 1 0 7681 0 1 13398
box 0 0 64 64
use contact_9  contact_9_1173
timestamp 1624494425
transform 1 0 8076 0 1 13393
box 0 0 66 74
use contact_8  contact_8_1173
timestamp 1624494425
transform 1 0 8077 0 1 13398
box 0 0 64 64
use contact_9  contact_9_438
timestamp 1624494425
transform 1 0 7680 0 1 14183
box 0 0 66 74
use contact_8  contact_8_438
timestamp 1624494425
transform 1 0 7681 0 1 14188
box 0 0 64 64
use contact_9  contact_9_440
timestamp 1624494425
transform 1 0 7680 0 1 13788
box 0 0 66 74
use contact_8  contact_8_440
timestamp 1624494425
transform 1 0 7681 0 1 13793
box 0 0 64 64
use contact_9  contact_9_1167
timestamp 1624494425
transform 1 0 8076 0 1 14183
box 0 0 66 74
use contact_8  contact_8_1167
timestamp 1624494425
transform 1 0 8077 0 1 14188
box 0 0 64 64
use contact_9  contact_9_1170
timestamp 1624494425
transform 1 0 8076 0 1 13788
box 0 0 66 74
use contact_8  contact_8_1170
timestamp 1624494425
transform 1 0 8077 0 1 13793
box 0 0 64 64
use contact_9  contact_9_436
timestamp 1624494425
transform 1 0 7680 0 1 14578
box 0 0 66 74
use contact_8  contact_8_436
timestamp 1624494425
transform 1 0 7681 0 1 14583
box 0 0 64 64
use contact_9  contact_9_1164
timestamp 1624494425
transform 1 0 8076 0 1 14578
box 0 0 66 74
use contact_8  contact_8_1164
timestamp 1624494425
transform 1 0 8077 0 1 14583
box 0 0 64 64
use contact_9  contact_9_432
timestamp 1624494425
transform 1 0 7680 0 1 15368
box 0 0 66 74
use contact_8  contact_8_432
timestamp 1624494425
transform 1 0 7681 0 1 15373
box 0 0 64 64
use contact_9  contact_9_434
timestamp 1624494425
transform 1 0 7680 0 1 14973
box 0 0 66 74
use contact_8  contact_8_434
timestamp 1624494425
transform 1 0 7681 0 1 14978
box 0 0 64 64
use contact_9  contact_9_1158
timestamp 1624494425
transform 1 0 8076 0 1 15368
box 0 0 66 74
use contact_8  contact_8_1158
timestamp 1624494425
transform 1 0 8077 0 1 15373
box 0 0 64 64
use contact_9  contact_9_1161
timestamp 1624494425
transform 1 0 8076 0 1 14973
box 0 0 66 74
use contact_8  contact_8_1161
timestamp 1624494425
transform 1 0 8077 0 1 14978
box 0 0 64 64
use contact_9  contact_9_428
timestamp 1624494425
transform 1 0 7680 0 1 16158
box 0 0 66 74
use contact_8  contact_8_428
timestamp 1624494425
transform 1 0 7681 0 1 16163
box 0 0 64 64
use contact_9  contact_9_430
timestamp 1624494425
transform 1 0 7680 0 1 15763
box 0 0 66 74
use contact_8  contact_8_430
timestamp 1624494425
transform 1 0 7681 0 1 15768
box 0 0 64 64
use contact_9  contact_9_1152
timestamp 1624494425
transform 1 0 8076 0 1 16158
box 0 0 66 74
use contact_8  contact_8_1152
timestamp 1624494425
transform 1 0 8077 0 1 16163
box 0 0 64 64
use contact_9  contact_9_1155
timestamp 1624494425
transform 1 0 8076 0 1 15763
box 0 0 66 74
use contact_8  contact_8_1155
timestamp 1624494425
transform 1 0 8077 0 1 15768
box 0 0 64 64
use contact_8  contact_8_1151
timestamp 1624494425
transform 1 0 7299 0 1 16544
box 0 0 64 64
use contact_9  contact_9_1151
timestamp 1624494425
transform 1 0 7298 0 1 16539
box 0 0 66 74
use contact_8  contact_8_1150
timestamp 1624494425
transform 1 0 6867 0 1 16544
box 0 0 64 64
use contact_9  contact_9_1150
timestamp 1624494425
transform 1 0 6866 0 1 16539
box 0 0 66 74
use contact_8  contact_8_427
timestamp 1624494425
transform 1 0 6442 0 1 16602
box 0 0 64 64
use contact_9  contact_9_427
timestamp 1624494425
transform 1 0 6441 0 1 16597
box 0 0 66 74
use contact_16  contact_16_643
timestamp 1624494425
transform 1 0 5064 0 1 16368
box 0 0 66 58
use contact_16  contact_16_644
timestamp 1624494425
transform 1 0 4664 0 1 16480
box 0 0 66 58
use contact_16  contact_16_639
timestamp 1624494425
transform 1 0 5624 0 1 16844
box 0 0 66 58
use contact_16  contact_16_640
timestamp 1624494425
transform 1 0 5064 0 1 16754
box 0 0 66 58
use contact_16  contact_16_641
timestamp 1624494425
transform 1 0 4744 0 1 16642
box 0 0 66 58
use and3_dec  and3_dec_212
timestamp 1624494425
transform 1 0 6203 0 -1 17380
box 0 -60 2072 490
use and3_dec  and3_dec_213
timestamp 1624494425
transform 1 0 6203 0 1 16590
box 0 -60 2072 490
use contact_8  contact_8_1148
timestamp 1624494425
transform 1 0 7299 0 1 16976
box 0 0 64 64
use contact_9  contact_9_1148
timestamp 1624494425
transform 1 0 7298 0 1 16971
box 0 0 66 74
use contact_8  contact_8_1147
timestamp 1624494425
transform 1 0 6867 0 1 16976
box 0 0 64 64
use contact_9  contact_9_1147
timestamp 1624494425
transform 1 0 6866 0 1 16971
box 0 0 66 74
use contact_8  contact_8_425
timestamp 1624494425
transform 1 0 6442 0 1 16976
box 0 0 64 64
use contact_9  contact_9_425
timestamp 1624494425
transform 1 0 6441 0 1 16971
box 0 0 66 74
use contact_16  contact_16_636
timestamp 1624494425
transform 1 0 5624 0 1 17068
box 0 0 66 58
use contact_16  contact_16_637
timestamp 1624494425
transform 1 0 5064 0 1 17158
box 0 0 66 58
use contact_8  contact_8_1145
timestamp 1624494425
transform 1 0 7299 0 1 17334
box 0 0 64 64
use contact_9  contact_9_1145
timestamp 1624494425
transform 1 0 7298 0 1 17329
box 0 0 66 74
use contact_8  contact_8_1144
timestamp 1624494425
transform 1 0 6867 0 1 17334
box 0 0 64 64
use contact_9  contact_9_1144
timestamp 1624494425
transform 1 0 6866 0 1 17329
box 0 0 66 74
use contact_8  contact_8_423
timestamp 1624494425
transform 1 0 6442 0 1 17392
box 0 0 64 64
use contact_9  contact_9_423
timestamp 1624494425
transform 1 0 6441 0 1 17387
box 0 0 66 74
use contact_16  contact_16_635
timestamp 1624494425
transform 1 0 4584 0 1 17432
box 0 0 66 58
use contact_16  contact_16_638
timestamp 1624494425
transform 1 0 4824 0 1 17270
box 0 0 66 58
use and3_dec  and3_dec_211
timestamp 1624494425
transform 1 0 6203 0 1 17380
box 0 -60 2072 490
use contact_16  contact_16_633
timestamp 1624494425
transform 1 0 5624 0 1 17634
box 0 0 66 58
use contact_16  contact_16_634
timestamp 1624494425
transform 1 0 5144 0 1 17544
box 0 0 66 58
use contact_8  contact_8_1142
timestamp 1624494425
transform 1 0 7299 0 1 17766
box 0 0 64 64
use contact_9  contact_9_1142
timestamp 1624494425
transform 1 0 7298 0 1 17761
box 0 0 66 74
use contact_8  contact_8_1141
timestamp 1624494425
transform 1 0 6867 0 1 17766
box 0 0 64 64
use contact_9  contact_9_1141
timestamp 1624494425
transform 1 0 6866 0 1 17761
box 0 0 66 74
use contact_8  contact_8_421
timestamp 1624494425
transform 1 0 6442 0 1 17766
box 0 0 64 64
use contact_9  contact_9_421
timestamp 1624494425
transform 1 0 6441 0 1 17761
box 0 0 66 74
use contact_16  contact_16_630
timestamp 1624494425
transform 1 0 5624 0 1 17858
box 0 0 66 58
use contact_16  contact_16_631
timestamp 1624494425
transform 1 0 5144 0 1 17948
box 0 0 66 58
use and3_dec  and3_dec_210
timestamp 1624494425
transform 1 0 6203 0 -1 18170
box 0 -60 2072 490
use contact_8  contact_8_1139
timestamp 1624494425
transform 1 0 7299 0 1 18124
box 0 0 64 64
use contact_9  contact_9_1139
timestamp 1624494425
transform 1 0 7298 0 1 18119
box 0 0 66 74
use contact_8  contact_8_1138
timestamp 1624494425
transform 1 0 6867 0 1 18124
box 0 0 64 64
use contact_9  contact_9_1138
timestamp 1624494425
transform 1 0 6866 0 1 18119
box 0 0 66 74
use contact_8  contact_8_419
timestamp 1624494425
transform 1 0 6442 0 1 18182
box 0 0 64 64
use contact_9  contact_9_419
timestamp 1624494425
transform 1 0 6441 0 1 18177
box 0 0 66 74
use contact_16  contact_16_629
timestamp 1624494425
transform 1 0 4744 0 1 18222
box 0 0 66 58
use contact_16  contact_16_632
timestamp 1624494425
transform 1 0 4664 0 1 18060
box 0 0 66 58
use contact_16  contact_16_627
timestamp 1624494425
transform 1 0 5624 0 1 18424
box 0 0 66 58
use contact_16  contact_16_628
timestamp 1624494425
transform 1 0 5144 0 1 18334
box 0 0 66 58
use and3_dec  and3_dec_208
timestamp 1624494425
transform 1 0 6203 0 -1 18960
box 0 -60 2072 490
use and3_dec  and3_dec_209
timestamp 1624494425
transform 1 0 6203 0 1 18170
box 0 -60 2072 490
use contact_8  contact_8_1136
timestamp 1624494425
transform 1 0 7299 0 1 18556
box 0 0 64 64
use contact_9  contact_9_1136
timestamp 1624494425
transform 1 0 7298 0 1 18551
box 0 0 66 74
use contact_8  contact_8_1135
timestamp 1624494425
transform 1 0 6867 0 1 18556
box 0 0 64 64
use contact_9  contact_9_1135
timestamp 1624494425
transform 1 0 6866 0 1 18551
box 0 0 66 74
use contact_8  contact_8_417
timestamp 1624494425
transform 1 0 6442 0 1 18556
box 0 0 64 64
use contact_9  contact_9_417
timestamp 1624494425
transform 1 0 6441 0 1 18551
box 0 0 66 74
use contact_16  contact_16_624
timestamp 1624494425
transform 1 0 5624 0 1 18648
box 0 0 66 58
use contact_16  contact_16_625
timestamp 1624494425
transform 1 0 5144 0 1 18738
box 0 0 66 58
use contact_8  contact_8_1133
timestamp 1624494425
transform 1 0 7299 0 1 18914
box 0 0 64 64
use contact_9  contact_9_1133
timestamp 1624494425
transform 1 0 7298 0 1 18909
box 0 0 66 74
use contact_8  contact_8_1132
timestamp 1624494425
transform 1 0 6867 0 1 18914
box 0 0 64 64
use contact_9  contact_9_1132
timestamp 1624494425
transform 1 0 6866 0 1 18909
box 0 0 66 74
use contact_8  contact_8_415
timestamp 1624494425
transform 1 0 6442 0 1 18972
box 0 0 64 64
use contact_9  contact_9_415
timestamp 1624494425
transform 1 0 6441 0 1 18967
box 0 0 66 74
use contact_16  contact_16_623
timestamp 1624494425
transform 1 0 4584 0 1 19012
box 0 0 66 58
use contact_16  contact_16_626
timestamp 1624494425
transform 1 0 4824 0 1 18850
box 0 0 66 58
use and3_dec  and3_dec_207
timestamp 1624494425
transform 1 0 6203 0 1 18960
box 0 -60 2072 490
use contact_8  contact_8_1130
timestamp 1624494425
transform 1 0 7299 0 1 19346
box 0 0 64 64
use contact_9  contact_9_1130
timestamp 1624494425
transform 1 0 7298 0 1 19341
box 0 0 66 74
use contact_8  contact_8_1129
timestamp 1624494425
transform 1 0 6867 0 1 19346
box 0 0 64 64
use contact_9  contact_9_1129
timestamp 1624494425
transform 1 0 6866 0 1 19341
box 0 0 66 74
use contact_8  contact_8_413
timestamp 1624494425
transform 1 0 6442 0 1 19346
box 0 0 64 64
use contact_9  contact_9_413
timestamp 1624494425
transform 1 0 6441 0 1 19341
box 0 0 66 74
use contact_16  contact_16_621
timestamp 1624494425
transform 1 0 5624 0 1 19214
box 0 0 66 58
use contact_16  contact_16_622
timestamp 1624494425
transform 1 0 5224 0 1 19124
box 0 0 66 58
use contact_16  contact_16_618
timestamp 1624494425
transform 1 0 5624 0 1 19438
box 0 0 66 58
use contact_16  contact_16_619
timestamp 1624494425
transform 1 0 5224 0 1 19528
box 0 0 66 58
use and3_dec  and3_dec_206
timestamp 1624494425
transform 1 0 6203 0 -1 19750
box 0 -60 2072 490
use contact_9  contact_9_424
timestamp 1624494425
transform 1 0 7680 0 1 16948
box 0 0 66 74
use contact_8  contact_8_424
timestamp 1624494425
transform 1 0 7681 0 1 16953
box 0 0 64 64
use contact_9  contact_9_426
timestamp 1624494425
transform 1 0 7680 0 1 16553
box 0 0 66 74
use contact_8  contact_8_426
timestamp 1624494425
transform 1 0 7681 0 1 16558
box 0 0 64 64
use contact_9  contact_9_1146
timestamp 1624494425
transform 1 0 8076 0 1 16948
box 0 0 66 74
use contact_8  contact_8_1146
timestamp 1624494425
transform 1 0 8077 0 1 16953
box 0 0 64 64
use contact_9  contact_9_1149
timestamp 1624494425
transform 1 0 8076 0 1 16553
box 0 0 66 74
use contact_8  contact_8_1149
timestamp 1624494425
transform 1 0 8077 0 1 16558
box 0 0 64 64
use contact_9  contact_9_422
timestamp 1624494425
transform 1 0 7680 0 1 17343
box 0 0 66 74
use contact_8  contact_8_422
timestamp 1624494425
transform 1 0 7681 0 1 17348
box 0 0 64 64
use contact_9  contact_9_1143
timestamp 1624494425
transform 1 0 8076 0 1 17343
box 0 0 66 74
use contact_8  contact_8_1143
timestamp 1624494425
transform 1 0 8077 0 1 17348
box 0 0 64 64
use contact_9  contact_9_418
timestamp 1624494425
transform 1 0 7680 0 1 18133
box 0 0 66 74
use contact_8  contact_8_418
timestamp 1624494425
transform 1 0 7681 0 1 18138
box 0 0 64 64
use contact_9  contact_9_420
timestamp 1624494425
transform 1 0 7680 0 1 17738
box 0 0 66 74
use contact_8  contact_8_420
timestamp 1624494425
transform 1 0 7681 0 1 17743
box 0 0 64 64
use contact_9  contact_9_1137
timestamp 1624494425
transform 1 0 8076 0 1 18133
box 0 0 66 74
use contact_8  contact_8_1137
timestamp 1624494425
transform 1 0 8077 0 1 18138
box 0 0 64 64
use contact_9  contact_9_1140
timestamp 1624494425
transform 1 0 8076 0 1 17738
box 0 0 66 74
use contact_8  contact_8_1140
timestamp 1624494425
transform 1 0 8077 0 1 17743
box 0 0 64 64
use contact_9  contact_9_416
timestamp 1624494425
transform 1 0 7680 0 1 18528
box 0 0 66 74
use contact_8  contact_8_416
timestamp 1624494425
transform 1 0 7681 0 1 18533
box 0 0 64 64
use contact_9  contact_9_1134
timestamp 1624494425
transform 1 0 8076 0 1 18528
box 0 0 66 74
use contact_8  contact_8_1134
timestamp 1624494425
transform 1 0 8077 0 1 18533
box 0 0 64 64
use contact_9  contact_9_412
timestamp 1624494425
transform 1 0 7680 0 1 19318
box 0 0 66 74
use contact_8  contact_8_412
timestamp 1624494425
transform 1 0 7681 0 1 19323
box 0 0 64 64
use contact_9  contact_9_414
timestamp 1624494425
transform 1 0 7680 0 1 18923
box 0 0 66 74
use contact_8  contact_8_414
timestamp 1624494425
transform 1 0 7681 0 1 18928
box 0 0 64 64
use contact_9  contact_9_1128
timestamp 1624494425
transform 1 0 8076 0 1 19318
box 0 0 66 74
use contact_8  contact_8_1128
timestamp 1624494425
transform 1 0 8077 0 1 19323
box 0 0 64 64
use contact_9  contact_9_1131
timestamp 1624494425
transform 1 0 8076 0 1 18923
box 0 0 66 74
use contact_8  contact_8_1131
timestamp 1624494425
transform 1 0 8077 0 1 18928
box 0 0 64 64
use contact_8  contact_8_1127
timestamp 1624494425
transform 1 0 7299 0 1 19704
box 0 0 64 64
use contact_9  contact_9_1127
timestamp 1624494425
transform 1 0 7298 0 1 19699
box 0 0 66 74
use contact_8  contact_8_1126
timestamp 1624494425
transform 1 0 6867 0 1 19704
box 0 0 64 64
use contact_9  contact_9_1126
timestamp 1624494425
transform 1 0 6866 0 1 19699
box 0 0 66 74
use contact_8  contact_8_411
timestamp 1624494425
transform 1 0 6442 0 1 19762
box 0 0 64 64
use contact_9  contact_9_411
timestamp 1624494425
transform 1 0 6441 0 1 19757
box 0 0 66 74
use contact_16  contact_16_617
timestamp 1624494425
transform 1 0 4744 0 1 19802
box 0 0 66 58
use contact_16  contact_16_620
timestamp 1624494425
transform 1 0 4664 0 1 19640
box 0 0 66 58
use contact_8  contact_8_1124
timestamp 1624494425
transform 1 0 7299 0 1 20136
box 0 0 64 64
use contact_9  contact_9_1124
timestamp 1624494425
transform 1 0 7298 0 1 20131
box 0 0 66 74
use contact_8  contact_8_1123
timestamp 1624494425
transform 1 0 6867 0 1 20136
box 0 0 64 64
use contact_9  contact_9_1123
timestamp 1624494425
transform 1 0 6866 0 1 20131
box 0 0 66 74
use contact_8  contact_8_409
timestamp 1624494425
transform 1 0 6442 0 1 20136
box 0 0 64 64
use contact_9  contact_9_409
timestamp 1624494425
transform 1 0 6441 0 1 20131
box 0 0 66 74
use contact_16  contact_16_615
timestamp 1624494425
transform 1 0 5624 0 1 20004
box 0 0 66 58
use contact_16  contact_16_616
timestamp 1624494425
transform 1 0 5224 0 1 19914
box 0 0 66 58
use and3_dec  and3_dec_204
timestamp 1624494425
transform 1 0 6203 0 -1 20540
box 0 -60 2072 490
use and3_dec  and3_dec_205
timestamp 1624494425
transform 1 0 6203 0 1 19750
box 0 -60 2072 490
use contact_16  contact_16_612
timestamp 1624494425
transform 1 0 5624 0 1 20228
box 0 0 66 58
use contact_16  contact_16_613
timestamp 1624494425
transform 1 0 5224 0 1 20318
box 0 0 66 58
use contact_16  contact_16_614
timestamp 1624494425
transform 1 0 4824 0 1 20430
box 0 0 66 58
use contact_8  contact_8_1121
timestamp 1624494425
transform 1 0 7299 0 1 20494
box 0 0 64 64
use contact_9  contact_9_1121
timestamp 1624494425
transform 1 0 7298 0 1 20489
box 0 0 66 74
use contact_8  contact_8_1120
timestamp 1624494425
transform 1 0 6867 0 1 20494
box 0 0 64 64
use contact_9  contact_9_1120
timestamp 1624494425
transform 1 0 6866 0 1 20489
box 0 0 66 74
use contact_8  contact_8_407
timestamp 1624494425
transform 1 0 6442 0 1 20552
box 0 0 64 64
use contact_9  contact_9_407
timestamp 1624494425
transform 1 0 6441 0 1 20547
box 0 0 66 74
use contact_16  contact_16_610
timestamp 1624494425
transform 1 0 5304 0 1 20704
box 0 0 66 58
use contact_16  contact_16_611
timestamp 1624494425
transform 1 0 4584 0 1 20592
box 0 0 66 58
use and3_dec  and3_dec_203
timestamp 1624494425
transform 1 0 6203 0 1 20540
box 0 -60 2072 490
use contact_8  contact_8_1118
timestamp 1624494425
transform 1 0 7299 0 1 20926
box 0 0 64 64
use contact_9  contact_9_1118
timestamp 1624494425
transform 1 0 7298 0 1 20921
box 0 0 66 74
use contact_8  contact_8_1117
timestamp 1624494425
transform 1 0 6867 0 1 20926
box 0 0 64 64
use contact_9  contact_9_1117
timestamp 1624494425
transform 1 0 6866 0 1 20921
box 0 0 66 74
use contact_8  contact_8_405
timestamp 1624494425
transform 1 0 6442 0 1 20926
box 0 0 64 64
use contact_9  contact_9_405
timestamp 1624494425
transform 1 0 6441 0 1 20921
box 0 0 66 74
use contact_16  contact_16_609
timestamp 1624494425
transform 1 0 5624 0 1 20794
box 0 0 66 58
use contact_16  contact_16_606
timestamp 1624494425
transform 1 0 5624 0 1 21018
box 0 0 66 58
use contact_16  contact_16_607
timestamp 1624494425
transform 1 0 5304 0 1 21108
box 0 0 66 58
use contact_16  contact_16_608
timestamp 1624494425
transform 1 0 4664 0 1 21220
box 0 0 66 58
use and3_dec  and3_dec_201
timestamp 1624494425
transform 1 0 6203 0 1 21330
box 0 -60 2072 490
use and3_dec  and3_dec_202
timestamp 1624494425
transform 1 0 6203 0 -1 21330
box 0 -60 2072 490
use contact_8  contact_8_1115
timestamp 1624494425
transform 1 0 7299 0 1 21284
box 0 0 64 64
use contact_9  contact_9_1115
timestamp 1624494425
transform 1 0 7298 0 1 21279
box 0 0 66 74
use contact_8  contact_8_1114
timestamp 1624494425
transform 1 0 6867 0 1 21284
box 0 0 64 64
use contact_9  contact_9_1114
timestamp 1624494425
transform 1 0 6866 0 1 21279
box 0 0 66 74
use contact_8  contact_8_403
timestamp 1624494425
transform 1 0 6442 0 1 21342
box 0 0 64 64
use contact_9  contact_9_403
timestamp 1624494425
transform 1 0 6441 0 1 21337
box 0 0 66 74
use contact_16  contact_16_604
timestamp 1624494425
transform 1 0 5304 0 1 21494
box 0 0 66 58
use contact_16  contact_16_605
timestamp 1624494425
transform 1 0 4744 0 1 21382
box 0 0 66 58
use contact_8  contact_8_1112
timestamp 1624494425
transform 1 0 7299 0 1 21716
box 0 0 64 64
use contact_9  contact_9_1112
timestamp 1624494425
transform 1 0 7298 0 1 21711
box 0 0 66 74
use contact_8  contact_8_1111
timestamp 1624494425
transform 1 0 6867 0 1 21716
box 0 0 64 64
use contact_9  contact_9_1111
timestamp 1624494425
transform 1 0 6866 0 1 21711
box 0 0 66 74
use contact_8  contact_8_401
timestamp 1624494425
transform 1 0 6442 0 1 21716
box 0 0 64 64
use contact_9  contact_9_401
timestamp 1624494425
transform 1 0 6441 0 1 21711
box 0 0 66 74
use contact_16  contact_16_600
timestamp 1624494425
transform 1 0 5624 0 1 21808
box 0 0 66 58
use contact_16  contact_16_603
timestamp 1624494425
transform 1 0 5624 0 1 21584
box 0 0 66 58
use and3_dec  and3_dec_200
timestamp 1624494425
transform 1 0 6203 0 -1 22120
box 0 -60 2072 490
use contact_8  contact_8_1109
timestamp 1624494425
transform 1 0 7299 0 1 22074
box 0 0 64 64
use contact_9  contact_9_1109
timestamp 1624494425
transform 1 0 7298 0 1 22069
box 0 0 66 74
use contact_8  contact_8_1108
timestamp 1624494425
transform 1 0 6867 0 1 22074
box 0 0 64 64
use contact_9  contact_9_1108
timestamp 1624494425
transform 1 0 6866 0 1 22069
box 0 0 66 74
use contact_16  contact_16_601
timestamp 1624494425
transform 1 0 5304 0 1 21898
box 0 0 66 58
use contact_16  contact_16_602
timestamp 1624494425
transform 1 0 4824 0 1 22010
box 0 0 66 58
use contact_8  contact_8_399
timestamp 1624494425
transform 1 0 6442 0 1 22132
box 0 0 64 64
use contact_9  contact_9_399
timestamp 1624494425
transform 1 0 6441 0 1 22127
box 0 0 66 74
use contact_16  contact_16_597
timestamp 1624494425
transform 1 0 5624 0 1 22374
box 0 0 66 58
use contact_16  contact_16_598
timestamp 1624494425
transform 1 0 5384 0 1 22284
box 0 0 66 58
use contact_16  contact_16_599
timestamp 1624494425
transform 1 0 4584 0 1 22172
box 0 0 66 58
use and3_dec  and3_dec_199
timestamp 1624494425
transform 1 0 6203 0 1 22120
box 0 -60 2072 490
use contact_8  contact_8_1106
timestamp 1624494425
transform 1 0 7299 0 1 22506
box 0 0 64 64
use contact_9  contact_9_1106
timestamp 1624494425
transform 1 0 7298 0 1 22501
box 0 0 66 74
use contact_8  contact_8_1105
timestamp 1624494425
transform 1 0 6867 0 1 22506
box 0 0 64 64
use contact_9  contact_9_1105
timestamp 1624494425
transform 1 0 6866 0 1 22501
box 0 0 66 74
use contact_8  contact_8_397
timestamp 1624494425
transform 1 0 6442 0 1 22506
box 0 0 64 64
use contact_9  contact_9_397
timestamp 1624494425
transform 1 0 6441 0 1 22501
box 0 0 66 74
use contact_16  contact_16_594
timestamp 1624494425
transform 1 0 5624 0 1 22598
box 0 0 66 58
use contact_8  contact_8_1103
timestamp 1624494425
transform 1 0 7299 0 1 22864
box 0 0 64 64
use contact_9  contact_9_1103
timestamp 1624494425
transform 1 0 7298 0 1 22859
box 0 0 66 74
use contact_8  contact_8_1102
timestamp 1624494425
transform 1 0 6867 0 1 22864
box 0 0 64 64
use contact_9  contact_9_1102
timestamp 1624494425
transform 1 0 6866 0 1 22859
box 0 0 66 74
use contact_16  contact_16_595
timestamp 1624494425
transform 1 0 5384 0 1 22688
box 0 0 66 58
use contact_16  contact_16_596
timestamp 1624494425
transform 1 0 4664 0 1 22800
box 0 0 66 58
use and3_dec  and3_dec_197
timestamp 1624494425
transform 1 0 6203 0 1 22910
box 0 -60 2072 490
use and3_dec  and3_dec_198
timestamp 1624494425
transform 1 0 6203 0 -1 22910
box 0 -60 2072 490
use contact_9  contact_9_408
timestamp 1624494425
transform 1 0 7680 0 1 20108
box 0 0 66 74
use contact_8  contact_8_408
timestamp 1624494425
transform 1 0 7681 0 1 20113
box 0 0 64 64
use contact_9  contact_9_410
timestamp 1624494425
transform 1 0 7680 0 1 19713
box 0 0 66 74
use contact_8  contact_8_410
timestamp 1624494425
transform 1 0 7681 0 1 19718
box 0 0 64 64
use contact_9  contact_9_1122
timestamp 1624494425
transform 1 0 8076 0 1 20108
box 0 0 66 74
use contact_8  contact_8_1122
timestamp 1624494425
transform 1 0 8077 0 1 20113
box 0 0 64 64
use contact_9  contact_9_1125
timestamp 1624494425
transform 1 0 8076 0 1 19713
box 0 0 66 74
use contact_8  contact_8_1125
timestamp 1624494425
transform 1 0 8077 0 1 19718
box 0 0 64 64
use contact_9  contact_9_406
timestamp 1624494425
transform 1 0 7680 0 1 20503
box 0 0 66 74
use contact_8  contact_8_406
timestamp 1624494425
transform 1 0 7681 0 1 20508
box 0 0 64 64
use contact_9  contact_9_1119
timestamp 1624494425
transform 1 0 8076 0 1 20503
box 0 0 66 74
use contact_8  contact_8_1119
timestamp 1624494425
transform 1 0 8077 0 1 20508
box 0 0 64 64
use contact_9  contact_9_402
timestamp 1624494425
transform 1 0 7680 0 1 21293
box 0 0 66 74
use contact_8  contact_8_402
timestamp 1624494425
transform 1 0 7681 0 1 21298
box 0 0 64 64
use contact_9  contact_9_404
timestamp 1624494425
transform 1 0 7680 0 1 20898
box 0 0 66 74
use contact_8  contact_8_404
timestamp 1624494425
transform 1 0 7681 0 1 20903
box 0 0 64 64
use contact_9  contact_9_1113
timestamp 1624494425
transform 1 0 8076 0 1 21293
box 0 0 66 74
use contact_8  contact_8_1113
timestamp 1624494425
transform 1 0 8077 0 1 21298
box 0 0 64 64
use contact_9  contact_9_1116
timestamp 1624494425
transform 1 0 8076 0 1 20898
box 0 0 66 74
use contact_8  contact_8_1116
timestamp 1624494425
transform 1 0 8077 0 1 20903
box 0 0 64 64
use contact_9  contact_9_400
timestamp 1624494425
transform 1 0 7680 0 1 21688
box 0 0 66 74
use contact_8  contact_8_400
timestamp 1624494425
transform 1 0 7681 0 1 21693
box 0 0 64 64
use contact_9  contact_9_1110
timestamp 1624494425
transform 1 0 8076 0 1 21688
box 0 0 66 74
use contact_8  contact_8_1110
timestamp 1624494425
transform 1 0 8077 0 1 21693
box 0 0 64 64
use contact_9  contact_9_396
timestamp 1624494425
transform 1 0 7680 0 1 22478
box 0 0 66 74
use contact_8  contact_8_396
timestamp 1624494425
transform 1 0 7681 0 1 22483
box 0 0 64 64
use contact_9  contact_9_398
timestamp 1624494425
transform 1 0 7680 0 1 22083
box 0 0 66 74
use contact_8  contact_8_398
timestamp 1624494425
transform 1 0 7681 0 1 22088
box 0 0 64 64
use contact_9  contact_9_1104
timestamp 1624494425
transform 1 0 8076 0 1 22478
box 0 0 66 74
use contact_8  contact_8_1104
timestamp 1624494425
transform 1 0 8077 0 1 22483
box 0 0 64 64
use contact_9  contact_9_1107
timestamp 1624494425
transform 1 0 8076 0 1 22083
box 0 0 66 74
use contact_8  contact_8_1107
timestamp 1624494425
transform 1 0 8077 0 1 22088
box 0 0 64 64
use contact_9  contact_9_394
timestamp 1624494425
transform 1 0 7680 0 1 22873
box 0 0 66 74
use contact_8  contact_8_394
timestamp 1624494425
transform 1 0 7681 0 1 22878
box 0 0 64 64
use contact_9  contact_9_1101
timestamp 1624494425
transform 1 0 8076 0 1 22873
box 0 0 66 74
use contact_8  contact_8_1101
timestamp 1624494425
transform 1 0 8077 0 1 22878
box 0 0 64 64
use contact_8  contact_8_395
timestamp 1624494425
transform 1 0 6442 0 1 22922
box 0 0 64 64
use contact_9  contact_9_395
timestamp 1624494425
transform 1 0 6441 0 1 22917
box 0 0 66 74
use contact_16  contact_16_591
timestamp 1624494425
transform 1 0 5624 0 1 23164
box 0 0 66 58
use contact_16  contact_16_592
timestamp 1624494425
transform 1 0 5384 0 1 23074
box 0 0 66 58
use contact_16  contact_16_593
timestamp 1624494425
transform 1 0 4744 0 1 22962
box 0 0 66 58
use contact_8  contact_8_1100
timestamp 1624494425
transform 1 0 7299 0 1 23296
box 0 0 64 64
use contact_9  contact_9_1100
timestamp 1624494425
transform 1 0 7298 0 1 23291
box 0 0 66 74
use contact_8  contact_8_1099
timestamp 1624494425
transform 1 0 6867 0 1 23296
box 0 0 64 64
use contact_9  contact_9_1099
timestamp 1624494425
transform 1 0 6866 0 1 23291
box 0 0 66 74
use contact_8  contact_8_393
timestamp 1624494425
transform 1 0 6442 0 1 23296
box 0 0 64 64
use contact_9  contact_9_393
timestamp 1624494425
transform 1 0 6441 0 1 23291
box 0 0 66 74
use contact_16  contact_16_588
timestamp 1624494425
transform 1 0 5624 0 1 23388
box 0 0 66 58
use and3_dec  and3_dec_196
timestamp 1624494425
transform 1 0 6203 0 -1 23700
box 0 -60 2072 490
use contact_8  contact_8_1097
timestamp 1624494425
transform 1 0 7299 0 1 23654
box 0 0 64 64
use contact_9  contact_9_1097
timestamp 1624494425
transform 1 0 7298 0 1 23649
box 0 0 66 74
use contact_8  contact_8_1096
timestamp 1624494425
transform 1 0 6867 0 1 23654
box 0 0 64 64
use contact_9  contact_9_1096
timestamp 1624494425
transform 1 0 6866 0 1 23649
box 0 0 66 74
use contact_8  contact_8_391
timestamp 1624494425
transform 1 0 6442 0 1 23712
box 0 0 64 64
use contact_9  contact_9_391
timestamp 1624494425
transform 1 0 6441 0 1 23707
box 0 0 66 74
use contact_16  contact_16_589
timestamp 1624494425
transform 1 0 5384 0 1 23478
box 0 0 66 58
use contact_16  contact_16_590
timestamp 1624494425
transform 1 0 4824 0 1 23590
box 0 0 66 58
use contact_16  contact_16_585
timestamp 1624494425
transform 1 0 5624 0 1 23954
box 0 0 66 58
use contact_16  contact_16_586
timestamp 1624494425
transform 1 0 5464 0 1 23864
box 0 0 66 58
use contact_16  contact_16_587
timestamp 1624494425
transform 1 0 4584 0 1 23752
box 0 0 66 58
use and3_dec  and3_dec_194
timestamp 1624494425
transform 1 0 6203 0 -1 24490
box 0 -60 2072 490
use and3_dec  and3_dec_195
timestamp 1624494425
transform 1 0 6203 0 1 23700
box 0 -60 2072 490
use contact_8  contact_8_1094
timestamp 1624494425
transform 1 0 7299 0 1 24086
box 0 0 64 64
use contact_9  contact_9_1094
timestamp 1624494425
transform 1 0 7298 0 1 24081
box 0 0 66 74
use contact_8  contact_8_1093
timestamp 1624494425
transform 1 0 6867 0 1 24086
box 0 0 64 64
use contact_9  contact_9_1093
timestamp 1624494425
transform 1 0 6866 0 1 24081
box 0 0 66 74
use contact_8  contact_8_389
timestamp 1624494425
transform 1 0 6442 0 1 24086
box 0 0 64 64
use contact_9  contact_9_389
timestamp 1624494425
transform 1 0 6441 0 1 24081
box 0 0 66 74
use contact_16  contact_16_582
timestamp 1624494425
transform 1 0 5624 0 1 24178
box 0 0 66 58
use contact_16  contact_16_583
timestamp 1624494425
transform 1 0 5464 0 1 24268
box 0 0 66 58
use contact_8  contact_8_1091
timestamp 1624494425
transform 1 0 7299 0 1 24444
box 0 0 64 64
use contact_9  contact_9_1091
timestamp 1624494425
transform 1 0 7298 0 1 24439
box 0 0 66 74
use contact_8  contact_8_1090
timestamp 1624494425
transform 1 0 6867 0 1 24444
box 0 0 64 64
use contact_9  contact_9_1090
timestamp 1624494425
transform 1 0 6866 0 1 24439
box 0 0 66 74
use contact_8  contact_8_387
timestamp 1624494425
transform 1 0 6442 0 1 24502
box 0 0 64 64
use contact_9  contact_9_387
timestamp 1624494425
transform 1 0 6441 0 1 24497
box 0 0 66 74
use contact_16  contact_16_581
timestamp 1624494425
transform 1 0 4744 0 1 24542
box 0 0 66 58
use contact_16  contact_16_584
timestamp 1624494425
transform 1 0 4664 0 1 24380
box 0 0 66 58
use and3_dec  and3_dec_193
timestamp 1624494425
transform 1 0 6203 0 1 24490
box 0 -60 2072 490
use contact_16  contact_16_579
timestamp 1624494425
transform 1 0 5624 0 1 24744
box 0 0 66 58
use contact_16  contact_16_580
timestamp 1624494425
transform 1 0 5464 0 1 24654
box 0 0 66 58
use contact_8  contact_8_1088
timestamp 1624494425
transform 1 0 7299 0 1 24876
box 0 0 64 64
use contact_9  contact_9_1088
timestamp 1624494425
transform 1 0 7298 0 1 24871
box 0 0 66 74
use contact_8  contact_8_1087
timestamp 1624494425
transform 1 0 6867 0 1 24876
box 0 0 64 64
use contact_9  contact_9_1087
timestamp 1624494425
transform 1 0 6866 0 1 24871
box 0 0 66 74
use contact_8  contact_8_385
timestamp 1624494425
transform 1 0 6442 0 1 24876
box 0 0 64 64
use contact_9  contact_9_385
timestamp 1624494425
transform 1 0 6441 0 1 24871
box 0 0 66 74
use contact_16  contact_16_576
timestamp 1624494425
transform 1 0 5624 0 1 24968
box 0 0 66 58
use contact_16  contact_16_577
timestamp 1624494425
transform 1 0 5464 0 1 25058
box 0 0 66 58
use and3_dec  and3_dec_192
timestamp 1624494425
transform 1 0 6203 0 -1 25280
box 0 -60 2072 490
use contact_8  contact_8_1085
timestamp 1624494425
transform 1 0 7299 0 1 25234
box 0 0 64 64
use contact_9  contact_9_1085
timestamp 1624494425
transform 1 0 7298 0 1 25229
box 0 0 66 74
use contact_8  contact_8_1084
timestamp 1624494425
transform 1 0 6867 0 1 25234
box 0 0 64 64
use contact_9  contact_9_1084
timestamp 1624494425
transform 1 0 6866 0 1 25229
box 0 0 66 74
use contact_8  contact_8_383
timestamp 1624494425
transform 1 0 6442 0 1 25292
box 0 0 64 64
use contact_9  contact_9_383
timestamp 1624494425
transform 1 0 6441 0 1 25287
box 0 0 66 74
use contact_16  contact_16_575
timestamp 1624494425
transform 1 0 4584 0 1 25332
box 0 0 66 58
use contact_16  contact_16_578
timestamp 1624494425
transform 1 0 4824 0 1 25170
box 0 0 66 58
use contact_9  contact_9_1082
timestamp 1624494425
transform 1 0 7298 0 1 25661
box 0 0 66 74
use contact_9  contact_9_1081
timestamp 1624494425
transform 1 0 6866 0 1 25661
box 0 0 66 74
use contact_9  contact_9_381
timestamp 1624494425
transform 1 0 6441 0 1 25661
box 0 0 66 74
use contact_16  contact_16_573
timestamp 1624494425
transform 1 0 5704 0 1 25534
box 0 0 66 58
use contact_16  contact_16_574
timestamp 1624494425
transform 1 0 4904 0 1 25444
box 0 0 66 58
use and3_dec  and3_dec_190
timestamp 1624494425
transform 1 0 6203 0 -1 26070
box 0 -60 2072 490
use and3_dec  and3_dec_191
timestamp 1624494425
transform 1 0 6203 0 1 25280
box 0 -60 2072 490
use contact_8  contact_8_1082
timestamp 1624494425
transform 1 0 7299 0 1 25666
box 0 0 64 64
use contact_8  contact_8_1081
timestamp 1624494425
transform 1 0 6867 0 1 25666
box 0 0 64 64
use contact_8  contact_8_381
timestamp 1624494425
transform 1 0 6442 0 1 25666
box 0 0 64 64
use contact_16  contact_16_570
timestamp 1624494425
transform 1 0 5704 0 1 25758
box 0 0 66 58
use contact_16  contact_16_571
timestamp 1624494425
transform 1 0 4904 0 1 25848
box 0 0 66 58
use contact_8  contact_8_1079
timestamp 1624494425
transform 1 0 7299 0 1 26024
box 0 0 64 64
use contact_9  contact_9_1079
timestamp 1624494425
transform 1 0 7298 0 1 26019
box 0 0 66 74
use contact_8  contact_8_1078
timestamp 1624494425
transform 1 0 6867 0 1 26024
box 0 0 64 64
use contact_9  contact_9_1078
timestamp 1624494425
transform 1 0 6866 0 1 26019
box 0 0 66 74
use contact_8  contact_8_379
timestamp 1624494425
transform 1 0 6442 0 1 26082
box 0 0 64 64
use contact_9  contact_9_379
timestamp 1624494425
transform 1 0 6441 0 1 26077
box 0 0 66 74
use contact_16  contact_16_569
timestamp 1624494425
transform 1 0 4744 0 1 26122
box 0 0 66 58
use contact_16  contact_16_572
timestamp 1624494425
transform 1 0 4664 0 1 25960
box 0 0 66 58
use and3_dec  and3_dec_189
timestamp 1624494425
transform 1 0 6203 0 1 26070
box 0 -60 2072 490
use contact_9  contact_9_392
timestamp 1624494425
transform 1 0 7680 0 1 23268
box 0 0 66 74
use contact_8  contact_8_392
timestamp 1624494425
transform 1 0 7681 0 1 23273
box 0 0 64 64
use contact_9  contact_9_1098
timestamp 1624494425
transform 1 0 8076 0 1 23268
box 0 0 66 74
use contact_8  contact_8_1098
timestamp 1624494425
transform 1 0 8077 0 1 23273
box 0 0 64 64
use contact_9  contact_9_388
timestamp 1624494425
transform 1 0 7680 0 1 24058
box 0 0 66 74
use contact_8  contact_8_388
timestamp 1624494425
transform 1 0 7681 0 1 24063
box 0 0 64 64
use contact_9  contact_9_390
timestamp 1624494425
transform 1 0 7680 0 1 23663
box 0 0 66 74
use contact_8  contact_8_390
timestamp 1624494425
transform 1 0 7681 0 1 23668
box 0 0 64 64
use contact_9  contact_9_1092
timestamp 1624494425
transform 1 0 8076 0 1 24058
box 0 0 66 74
use contact_8  contact_8_1092
timestamp 1624494425
transform 1 0 8077 0 1 24063
box 0 0 64 64
use contact_9  contact_9_1095
timestamp 1624494425
transform 1 0 8076 0 1 23663
box 0 0 66 74
use contact_8  contact_8_1095
timestamp 1624494425
transform 1 0 8077 0 1 23668
box 0 0 64 64
use contact_9  contact_9_386
timestamp 1624494425
transform 1 0 7680 0 1 24453
box 0 0 66 74
use contact_8  contact_8_386
timestamp 1624494425
transform 1 0 7681 0 1 24458
box 0 0 64 64
use contact_9  contact_9_1089
timestamp 1624494425
transform 1 0 8076 0 1 24453
box 0 0 66 74
use contact_8  contact_8_1089
timestamp 1624494425
transform 1 0 8077 0 1 24458
box 0 0 64 64
use contact_9  contact_9_382
timestamp 1624494425
transform 1 0 7680 0 1 25243
box 0 0 66 74
use contact_8  contact_8_382
timestamp 1624494425
transform 1 0 7681 0 1 25248
box 0 0 64 64
use contact_9  contact_9_384
timestamp 1624494425
transform 1 0 7680 0 1 24848
box 0 0 66 74
use contact_8  contact_8_384
timestamp 1624494425
transform 1 0 7681 0 1 24853
box 0 0 64 64
use contact_9  contact_9_1083
timestamp 1624494425
transform 1 0 8076 0 1 25243
box 0 0 66 74
use contact_8  contact_8_1083
timestamp 1624494425
transform 1 0 8077 0 1 25248
box 0 0 64 64
use contact_9  contact_9_1086
timestamp 1624494425
transform 1 0 8076 0 1 24848
box 0 0 66 74
use contact_8  contact_8_1086
timestamp 1624494425
transform 1 0 8077 0 1 24853
box 0 0 64 64
use contact_9  contact_9_380
timestamp 1624494425
transform 1 0 7680 0 1 25638
box 0 0 66 74
use contact_8  contact_8_380
timestamp 1624494425
transform 1 0 7681 0 1 25643
box 0 0 64 64
use contact_9  contact_9_1080
timestamp 1624494425
transform 1 0 8076 0 1 25638
box 0 0 66 74
use contact_8  contact_8_1080
timestamp 1624494425
transform 1 0 8077 0 1 25643
box 0 0 64 64
use contact_9  contact_9_378
timestamp 1624494425
transform 1 0 7680 0 1 26033
box 0 0 66 74
use contact_8  contact_8_378
timestamp 1624494425
transform 1 0 7681 0 1 26038
box 0 0 64 64
use contact_9  contact_9_1077
timestamp 1624494425
transform 1 0 8076 0 1 26033
box 0 0 66 74
use contact_8  contact_8_1077
timestamp 1624494425
transform 1 0 8077 0 1 26038
box 0 0 64 64
use contact_8  contact_8_1076
timestamp 1624494425
transform 1 0 7299 0 1 26456
box 0 0 64 64
use contact_9  contact_9_1076
timestamp 1624494425
transform 1 0 7298 0 1 26451
box 0 0 66 74
use contact_8  contact_8_1075
timestamp 1624494425
transform 1 0 6867 0 1 26456
box 0 0 64 64
use contact_9  contact_9_1075
timestamp 1624494425
transform 1 0 6866 0 1 26451
box 0 0 66 74
use contact_8  contact_8_377
timestamp 1624494425
transform 1 0 6442 0 1 26456
box 0 0 64 64
use contact_9  contact_9_377
timestamp 1624494425
transform 1 0 6441 0 1 26451
box 0 0 66 74
use contact_16  contact_16_567
timestamp 1624494425
transform 1 0 5704 0 1 26324
box 0 0 66 58
use contact_16  contact_16_568
timestamp 1624494425
transform 1 0 4904 0 1 26234
box 0 0 66 58
use contact_16  contact_16_564
timestamp 1624494425
transform 1 0 5704 0 1 26548
box 0 0 66 58
use contact_16  contact_16_565
timestamp 1624494425
transform 1 0 4904 0 1 26638
box 0 0 66 58
use and3_dec  and3_dec_188
timestamp 1624494425
transform 1 0 6203 0 -1 26860
box 0 -60 2072 490
use contact_8  contact_8_1073
timestamp 1624494425
transform 1 0 7299 0 1 26814
box 0 0 64 64
use contact_9  contact_9_1073
timestamp 1624494425
transform 1 0 7298 0 1 26809
box 0 0 66 74
use contact_8  contact_8_1072
timestamp 1624494425
transform 1 0 6867 0 1 26814
box 0 0 64 64
use contact_9  contact_9_1072
timestamp 1624494425
transform 1 0 6866 0 1 26809
box 0 0 66 74
use contact_8  contact_8_375
timestamp 1624494425
transform 1 0 6442 0 1 26872
box 0 0 64 64
use contact_9  contact_9_375
timestamp 1624494425
transform 1 0 6441 0 1 26867
box 0 0 66 74
use contact_16  contact_16_563
timestamp 1624494425
transform 1 0 4584 0 1 26912
box 0 0 66 58
use contact_16  contact_16_566
timestamp 1624494425
transform 1 0 4824 0 1 26750
box 0 0 66 58
use contact_8  contact_8_1070
timestamp 1624494425
transform 1 0 7299 0 1 27246
box 0 0 64 64
use contact_9  contact_9_1070
timestamp 1624494425
transform 1 0 7298 0 1 27241
box 0 0 66 74
use contact_8  contact_8_1069
timestamp 1624494425
transform 1 0 6867 0 1 27246
box 0 0 64 64
use contact_9  contact_9_1069
timestamp 1624494425
transform 1 0 6866 0 1 27241
box 0 0 66 74
use contact_8  contact_8_373
timestamp 1624494425
transform 1 0 6442 0 1 27246
box 0 0 64 64
use contact_9  contact_9_373
timestamp 1624494425
transform 1 0 6441 0 1 27241
box 0 0 66 74
use contact_16  contact_16_561
timestamp 1624494425
transform 1 0 5704 0 1 27114
box 0 0 66 58
use contact_16  contact_16_562
timestamp 1624494425
transform 1 0 4984 0 1 27024
box 0 0 66 58
use and3_dec  and3_dec_186
timestamp 1624494425
transform 1 0 6203 0 -1 27650
box 0 -60 2072 490
use and3_dec  and3_dec_187
timestamp 1624494425
transform 1 0 6203 0 1 26860
box 0 -60 2072 490
use contact_16  contact_16_558
timestamp 1624494425
transform 1 0 5704 0 1 27338
box 0 0 66 58
use contact_16  contact_16_559
timestamp 1624494425
transform 1 0 4984 0 1 27428
box 0 0 66 58
use contact_16  contact_16_560
timestamp 1624494425
transform 1 0 4664 0 1 27540
box 0 0 66 58
use contact_8  contact_8_1067
timestamp 1624494425
transform 1 0 7299 0 1 27604
box 0 0 64 64
use contact_9  contact_9_1067
timestamp 1624494425
transform 1 0 7298 0 1 27599
box 0 0 66 74
use contact_8  contact_8_1066
timestamp 1624494425
transform 1 0 6867 0 1 27604
box 0 0 64 64
use contact_9  contact_9_1066
timestamp 1624494425
transform 1 0 6866 0 1 27599
box 0 0 66 74
use contact_8  contact_8_371
timestamp 1624494425
transform 1 0 6442 0 1 27662
box 0 0 64 64
use contact_9  contact_9_371
timestamp 1624494425
transform 1 0 6441 0 1 27657
box 0 0 66 74
use contact_16  contact_16_556
timestamp 1624494425
transform 1 0 4984 0 1 27814
box 0 0 66 58
use contact_16  contact_16_557
timestamp 1624494425
transform 1 0 4744 0 1 27702
box 0 0 66 58
use and3_dec  and3_dec_185
timestamp 1624494425
transform 1 0 6203 0 1 27650
box 0 -60 2072 490
use contact_8  contact_8_1064
timestamp 1624494425
transform 1 0 7299 0 1 28036
box 0 0 64 64
use contact_9  contact_9_1064
timestamp 1624494425
transform 1 0 7298 0 1 28031
box 0 0 66 74
use contact_8  contact_8_1063
timestamp 1624494425
transform 1 0 6867 0 1 28036
box 0 0 64 64
use contact_9  contact_9_1063
timestamp 1624494425
transform 1 0 6866 0 1 28031
box 0 0 66 74
use contact_8  contact_8_369
timestamp 1624494425
transform 1 0 6442 0 1 28036
box 0 0 64 64
use contact_9  contact_9_369
timestamp 1624494425
transform 1 0 6441 0 1 28031
box 0 0 66 74
use contact_16  contact_16_555
timestamp 1624494425
transform 1 0 5704 0 1 27904
box 0 0 66 58
use contact_9  contact_9_1061
timestamp 1624494425
transform 1 0 7298 0 1 28389
box 0 0 66 74
use contact_9  contact_9_1060
timestamp 1624494425
transform 1 0 6866 0 1 28389
box 0 0 66 74
use contact_16  contact_16_552
timestamp 1624494425
transform 1 0 5704 0 1 28128
box 0 0 66 58
use contact_16  contact_16_553
timestamp 1624494425
transform 1 0 4984 0 1 28218
box 0 0 66 58
use contact_16  contact_16_554
timestamp 1624494425
transform 1 0 4824 0 1 28330
box 0 0 66 58
use and3_dec  and3_dec_183
timestamp 1624494425
transform 1 0 6203 0 1 28440
box 0 -60 2072 490
use and3_dec  and3_dec_184
timestamp 1624494425
transform 1 0 6203 0 -1 28440
box 0 -60 2072 490
use contact_8  contact_8_1061
timestamp 1624494425
transform 1 0 7299 0 1 28394
box 0 0 64 64
use contact_8  contact_8_1060
timestamp 1624494425
transform 1 0 6867 0 1 28394
box 0 0 64 64
use contact_8  contact_8_367
timestamp 1624494425
transform 1 0 6442 0 1 28452
box 0 0 64 64
use contact_9  contact_9_367
timestamp 1624494425
transform 1 0 6441 0 1 28447
box 0 0 66 74
use contact_16  contact_16_550
timestamp 1624494425
transform 1 0 5064 0 1 28604
box 0 0 66 58
use contact_16  contact_16_551
timestamp 1624494425
transform 1 0 4584 0 1 28492
box 0 0 66 58
use contact_8  contact_8_1058
timestamp 1624494425
transform 1 0 7299 0 1 28826
box 0 0 64 64
use contact_9  contact_9_1058
timestamp 1624494425
transform 1 0 7298 0 1 28821
box 0 0 66 74
use contact_8  contact_8_1057
timestamp 1624494425
transform 1 0 6867 0 1 28826
box 0 0 64 64
use contact_9  contact_9_1057
timestamp 1624494425
transform 1 0 6866 0 1 28821
box 0 0 66 74
use contact_8  contact_8_365
timestamp 1624494425
transform 1 0 6442 0 1 28826
box 0 0 64 64
use contact_9  contact_9_365
timestamp 1624494425
transform 1 0 6441 0 1 28821
box 0 0 66 74
use contact_16  contact_16_546
timestamp 1624494425
transform 1 0 5704 0 1 28918
box 0 0 66 58
use contact_16  contact_16_549
timestamp 1624494425
transform 1 0 5704 0 1 28694
box 0 0 66 58
use and3_dec  and3_dec_182
timestamp 1624494425
transform 1 0 6203 0 -1 29230
box 0 -60 2072 490
use contact_8  contact_8_1055
timestamp 1624494425
transform 1 0 7299 0 1 29184
box 0 0 64 64
use contact_9  contact_9_1055
timestamp 1624494425
transform 1 0 7298 0 1 29179
box 0 0 66 74
use contact_8  contact_8_1054
timestamp 1624494425
transform 1 0 6867 0 1 29184
box 0 0 64 64
use contact_9  contact_9_1054
timestamp 1624494425
transform 1 0 6866 0 1 29179
box 0 0 66 74
use contact_16  contact_16_547
timestamp 1624494425
transform 1 0 5064 0 1 29008
box 0 0 66 58
use contact_16  contact_16_548
timestamp 1624494425
transform 1 0 4664 0 1 29120
box 0 0 66 58
use contact_8  contact_8_363
timestamp 1624494425
transform 1 0 6442 0 1 29242
box 0 0 64 64
use contact_9  contact_9_363
timestamp 1624494425
transform 1 0 6441 0 1 29237
box 0 0 66 74
use contact_16  contact_16_544
timestamp 1624494425
transform 1 0 5064 0 1 29394
box 0 0 66 58
use contact_16  contact_16_545
timestamp 1624494425
transform 1 0 4744 0 1 29282
box 0 0 66 58
use and3_dec  and3_dec_181
timestamp 1624494425
transform 1 0 6203 0 1 29230
box 0 -60 2072 490
use contact_9  contact_9_376
timestamp 1624494425
transform 1 0 7680 0 1 26428
box 0 0 66 74
use contact_8  contact_8_376
timestamp 1624494425
transform 1 0 7681 0 1 26433
box 0 0 64 64
use contact_9  contact_9_1074
timestamp 1624494425
transform 1 0 8076 0 1 26428
box 0 0 66 74
use contact_8  contact_8_1074
timestamp 1624494425
transform 1 0 8077 0 1 26433
box 0 0 64 64
use contact_9  contact_9_372
timestamp 1624494425
transform 1 0 7680 0 1 27218
box 0 0 66 74
use contact_8  contact_8_372
timestamp 1624494425
transform 1 0 7681 0 1 27223
box 0 0 64 64
use contact_9  contact_9_374
timestamp 1624494425
transform 1 0 7680 0 1 26823
box 0 0 66 74
use contact_8  contact_8_374
timestamp 1624494425
transform 1 0 7681 0 1 26828
box 0 0 64 64
use contact_9  contact_9_1068
timestamp 1624494425
transform 1 0 8076 0 1 27218
box 0 0 66 74
use contact_8  contact_8_1068
timestamp 1624494425
transform 1 0 8077 0 1 27223
box 0 0 64 64
use contact_9  contact_9_1071
timestamp 1624494425
transform 1 0 8076 0 1 26823
box 0 0 66 74
use contact_8  contact_8_1071
timestamp 1624494425
transform 1 0 8077 0 1 26828
box 0 0 64 64
use contact_9  contact_9_368
timestamp 1624494425
transform 1 0 7680 0 1 28008
box 0 0 66 74
use contact_8  contact_8_368
timestamp 1624494425
transform 1 0 7681 0 1 28013
box 0 0 64 64
use contact_9  contact_9_370
timestamp 1624494425
transform 1 0 7680 0 1 27613
box 0 0 66 74
use contact_8  contact_8_370
timestamp 1624494425
transform 1 0 7681 0 1 27618
box 0 0 64 64
use contact_9  contact_9_1062
timestamp 1624494425
transform 1 0 8076 0 1 28008
box 0 0 66 74
use contact_8  contact_8_1062
timestamp 1624494425
transform 1 0 8077 0 1 28013
box 0 0 64 64
use contact_9  contact_9_1065
timestamp 1624494425
transform 1 0 8076 0 1 27613
box 0 0 66 74
use contact_8  contact_8_1065
timestamp 1624494425
transform 1 0 8077 0 1 27618
box 0 0 64 64
use contact_9  contact_9_366
timestamp 1624494425
transform 1 0 7680 0 1 28403
box 0 0 66 74
use contact_8  contact_8_366
timestamp 1624494425
transform 1 0 7681 0 1 28408
box 0 0 64 64
use contact_9  contact_9_1059
timestamp 1624494425
transform 1 0 8076 0 1 28403
box 0 0 66 74
use contact_8  contact_8_1059
timestamp 1624494425
transform 1 0 8077 0 1 28408
box 0 0 64 64
use contact_9  contact_9_362
timestamp 1624494425
transform 1 0 7680 0 1 29193
box 0 0 66 74
use contact_8  contact_8_362
timestamp 1624494425
transform 1 0 7681 0 1 29198
box 0 0 64 64
use contact_9  contact_9_364
timestamp 1624494425
transform 1 0 7680 0 1 28798
box 0 0 66 74
use contact_8  contact_8_364
timestamp 1624494425
transform 1 0 7681 0 1 28803
box 0 0 64 64
use contact_9  contact_9_1053
timestamp 1624494425
transform 1 0 8076 0 1 29193
box 0 0 66 74
use contact_8  contact_8_1053
timestamp 1624494425
transform 1 0 8077 0 1 29198
box 0 0 64 64
use contact_9  contact_9_1056
timestamp 1624494425
transform 1 0 8076 0 1 28798
box 0 0 66 74
use contact_8  contact_8_1056
timestamp 1624494425
transform 1 0 8077 0 1 28803
box 0 0 64 64
use contact_8  contact_8_1052
timestamp 1624494425
transform 1 0 7299 0 1 29616
box 0 0 64 64
use contact_9  contact_9_1052
timestamp 1624494425
transform 1 0 7298 0 1 29611
box 0 0 66 74
use contact_8  contact_8_1051
timestamp 1624494425
transform 1 0 6867 0 1 29616
box 0 0 64 64
use contact_9  contact_9_1051
timestamp 1624494425
transform 1 0 6866 0 1 29611
box 0 0 66 74
use contact_8  contact_8_361
timestamp 1624494425
transform 1 0 6442 0 1 29616
box 0 0 64 64
use contact_9  contact_9_361
timestamp 1624494425
transform 1 0 6441 0 1 29611
box 0 0 66 74
use contact_16  contact_16_540
timestamp 1624494425
transform 1 0 5704 0 1 29708
box 0 0 66 58
use contact_16  contact_16_543
timestamp 1624494425
transform 1 0 5704 0 1 29484
box 0 0 66 58
use contact_8  contact_8_1049
timestamp 1624494425
transform 1 0 7299 0 1 29974
box 0 0 64 64
use contact_9  contact_9_1049
timestamp 1624494425
transform 1 0 7298 0 1 29969
box 0 0 66 74
use contact_8  contact_8_1048
timestamp 1624494425
transform 1 0 6867 0 1 29974
box 0 0 64 64
use contact_9  contact_9_1048
timestamp 1624494425
transform 1 0 6866 0 1 29969
box 0 0 66 74
use contact_16  contact_16_541
timestamp 1624494425
transform 1 0 5064 0 1 29798
box 0 0 66 58
use contact_16  contact_16_542
timestamp 1624494425
transform 1 0 4824 0 1 29910
box 0 0 66 58
use and3_dec  and3_dec_179
timestamp 1624494425
transform 1 0 6203 0 1 30020
box 0 -60 2072 490
use and3_dec  and3_dec_180
timestamp 1624494425
transform 1 0 6203 0 -1 30020
box 0 -60 2072 490
use contact_8  contact_8_359
timestamp 1624494425
transform 1 0 6442 0 1 30032
box 0 0 64 64
use contact_9  contact_9_359
timestamp 1624494425
transform 1 0 6441 0 1 30027
box 0 0 66 74
use contact_16  contact_16_537
timestamp 1624494425
transform 1 0 5704 0 1 30274
box 0 0 66 58
use contact_16  contact_16_538
timestamp 1624494425
transform 1 0 5144 0 1 30184
box 0 0 66 58
use contact_16  contact_16_539
timestamp 1624494425
transform 1 0 4584 0 1 30072
box 0 0 66 58
use contact_8  contact_8_1046
timestamp 1624494425
transform 1 0 7299 0 1 30406
box 0 0 64 64
use contact_9  contact_9_1046
timestamp 1624494425
transform 1 0 7298 0 1 30401
box 0 0 66 74
use contact_8  contact_8_1045
timestamp 1624494425
transform 1 0 6867 0 1 30406
box 0 0 64 64
use contact_9  contact_9_1045
timestamp 1624494425
transform 1 0 6866 0 1 30401
box 0 0 66 74
use contact_8  contact_8_357
timestamp 1624494425
transform 1 0 6442 0 1 30406
box 0 0 64 64
use contact_9  contact_9_357
timestamp 1624494425
transform 1 0 6441 0 1 30401
box 0 0 66 74
use contact_16  contact_16_534
timestamp 1624494425
transform 1 0 5704 0 1 30498
box 0 0 66 58
use and3_dec  and3_dec_178
timestamp 1624494425
transform 1 0 6203 0 -1 30810
box 0 -60 2072 490
use contact_8  contact_8_1043
timestamp 1624494425
transform 1 0 7299 0 1 30764
box 0 0 64 64
use contact_9  contact_9_1043
timestamp 1624494425
transform 1 0 7298 0 1 30759
box 0 0 66 74
use contact_8  contact_8_1042
timestamp 1624494425
transform 1 0 6867 0 1 30764
box 0 0 64 64
use contact_9  contact_9_1042
timestamp 1624494425
transform 1 0 6866 0 1 30759
box 0 0 66 74
use contact_8  contact_8_355
timestamp 1624494425
transform 1 0 6442 0 1 30822
box 0 0 64 64
use contact_9  contact_9_355
timestamp 1624494425
transform 1 0 6441 0 1 30817
box 0 0 66 74
use contact_16  contact_16_535
timestamp 1624494425
transform 1 0 5144 0 1 30588
box 0 0 66 58
use contact_16  contact_16_536
timestamp 1624494425
transform 1 0 4664 0 1 30700
box 0 0 66 58
use contact_16  contact_16_531
timestamp 1624494425
transform 1 0 5704 0 1 31064
box 0 0 66 58
use contact_16  contact_16_532
timestamp 1624494425
transform 1 0 5144 0 1 30974
box 0 0 66 58
use contact_16  contact_16_533
timestamp 1624494425
transform 1 0 4744 0 1 30862
box 0 0 66 58
use and3_dec  and3_dec_176
timestamp 1624494425
transform 1 0 6203 0 -1 31600
box 0 -60 2072 490
use and3_dec  and3_dec_177
timestamp 1624494425
transform 1 0 6203 0 1 30810
box 0 -60 2072 490
use contact_8  contact_8_1040
timestamp 1624494425
transform 1 0 7299 0 1 31196
box 0 0 64 64
use contact_9  contact_9_1040
timestamp 1624494425
transform 1 0 7298 0 1 31191
box 0 0 66 74
use contact_8  contact_8_1039
timestamp 1624494425
transform 1 0 6867 0 1 31196
box 0 0 64 64
use contact_9  contact_9_1039
timestamp 1624494425
transform 1 0 6866 0 1 31191
box 0 0 66 74
use contact_8  contact_8_353
timestamp 1624494425
transform 1 0 6442 0 1 31196
box 0 0 64 64
use contact_9  contact_9_353
timestamp 1624494425
transform 1 0 6441 0 1 31191
box 0 0 66 74
use contact_16  contact_16_528
timestamp 1624494425
transform 1 0 5704 0 1 31288
box 0 0 66 58
use contact_16  contact_16_529
timestamp 1624494425
transform 1 0 5144 0 1 31378
box 0 0 66 58
use contact_8  contact_8_1037
timestamp 1624494425
transform 1 0 7299 0 1 31554
box 0 0 64 64
use contact_9  contact_9_1037
timestamp 1624494425
transform 1 0 7298 0 1 31549
box 0 0 66 74
use contact_8  contact_8_1036
timestamp 1624494425
transform 1 0 6867 0 1 31554
box 0 0 64 64
use contact_9  contact_9_1036
timestamp 1624494425
transform 1 0 6866 0 1 31549
box 0 0 66 74
use contact_8  contact_8_351
timestamp 1624494425
transform 1 0 6442 0 1 31612
box 0 0 64 64
use contact_9  contact_9_351
timestamp 1624494425
transform 1 0 6441 0 1 31607
box 0 0 66 74
use contact_16  contact_16_527
timestamp 1624494425
transform 1 0 4584 0 1 31652
box 0 0 66 58
use contact_16  contact_16_530
timestamp 1624494425
transform 1 0 4824 0 1 31490
box 0 0 66 58
use and3_dec  and3_dec_175
timestamp 1624494425
transform 1 0 6203 0 1 31600
box 0 -60 2072 490
use contact_16  contact_16_525
timestamp 1624494425
transform 1 0 5704 0 1 31854
box 0 0 66 58
use contact_16  contact_16_526
timestamp 1624494425
transform 1 0 5224 0 1 31764
box 0 0 66 58
use contact_8  contact_8_1034
timestamp 1624494425
transform 1 0 7299 0 1 31986
box 0 0 64 64
use contact_9  contact_9_1034
timestamp 1624494425
transform 1 0 7298 0 1 31981
box 0 0 66 74
use contact_8  contact_8_1033
timestamp 1624494425
transform 1 0 6867 0 1 31986
box 0 0 64 64
use contact_9  contact_9_1033
timestamp 1624494425
transform 1 0 6866 0 1 31981
box 0 0 66 74
use contact_8  contact_8_349
timestamp 1624494425
transform 1 0 6442 0 1 31986
box 0 0 64 64
use contact_9  contact_9_349
timestamp 1624494425
transform 1 0 6441 0 1 31981
box 0 0 66 74
use contact_16  contact_16_522
timestamp 1624494425
transform 1 0 5704 0 1 32078
box 0 0 66 58
use contact_16  contact_16_523
timestamp 1624494425
transform 1 0 5224 0 1 32168
box 0 0 66 58
use and3_dec  and3_dec_174
timestamp 1624494425
transform 1 0 6203 0 -1 32390
box 0 -60 2072 490
use contact_8  contact_8_1031
timestamp 1624494425
transform 1 0 7299 0 1 32344
box 0 0 64 64
use contact_9  contact_9_1031
timestamp 1624494425
transform 1 0 7298 0 1 32339
box 0 0 66 74
use contact_8  contact_8_1030
timestamp 1624494425
transform 1 0 6867 0 1 32344
box 0 0 64 64
use contact_9  contact_9_1030
timestamp 1624494425
transform 1 0 6866 0 1 32339
box 0 0 66 74
use contact_8  contact_8_347
timestamp 1624494425
transform 1 0 6442 0 1 32402
box 0 0 64 64
use contact_9  contact_9_347
timestamp 1624494425
transform 1 0 6441 0 1 32397
box 0 0 66 74
use contact_16  contact_16_521
timestamp 1624494425
transform 1 0 4744 0 1 32442
box 0 0 66 58
use contact_16  contact_16_524
timestamp 1624494425
transform 1 0 4664 0 1 32280
box 0 0 66 58
use contact_16  contact_16_519
timestamp 1624494425
transform 1 0 5704 0 1 32644
box 0 0 66 58
use contact_16  contact_16_520
timestamp 1624494425
transform 1 0 5224 0 1 32554
box 0 0 66 58
use and3_dec  and3_dec_172
timestamp 1624494425
transform 1 0 6203 0 -1 33180
box 0 -60 2072 490
use and3_dec  and3_dec_173
timestamp 1624494425
transform 1 0 6203 0 1 32390
box 0 -60 2072 490
use contact_9  contact_9_358
timestamp 1624494425
transform 1 0 7680 0 1 29983
box 0 0 66 74
use contact_8  contact_8_358
timestamp 1624494425
transform 1 0 7681 0 1 29988
box 0 0 64 64
use contact_9  contact_9_360
timestamp 1624494425
transform 1 0 7680 0 1 29588
box 0 0 66 74
use contact_8  contact_8_360
timestamp 1624494425
transform 1 0 7681 0 1 29593
box 0 0 64 64
use contact_9  contact_9_1047
timestamp 1624494425
transform 1 0 8076 0 1 29983
box 0 0 66 74
use contact_8  contact_8_1047
timestamp 1624494425
transform 1 0 8077 0 1 29988
box 0 0 64 64
use contact_9  contact_9_1050
timestamp 1624494425
transform 1 0 8076 0 1 29588
box 0 0 66 74
use contact_8  contact_8_1050
timestamp 1624494425
transform 1 0 8077 0 1 29593
box 0 0 64 64
use contact_9  contact_9_356
timestamp 1624494425
transform 1 0 7680 0 1 30378
box 0 0 66 74
use contact_8  contact_8_356
timestamp 1624494425
transform 1 0 7681 0 1 30383
box 0 0 64 64
use contact_9  contact_9_1044
timestamp 1624494425
transform 1 0 8076 0 1 30378
box 0 0 66 74
use contact_8  contact_8_1044
timestamp 1624494425
transform 1 0 8077 0 1 30383
box 0 0 64 64
use contact_9  contact_9_352
timestamp 1624494425
transform 1 0 7680 0 1 31168
box 0 0 66 74
use contact_8  contact_8_352
timestamp 1624494425
transform 1 0 7681 0 1 31173
box 0 0 64 64
use contact_9  contact_9_354
timestamp 1624494425
transform 1 0 7680 0 1 30773
box 0 0 66 74
use contact_8  contact_8_354
timestamp 1624494425
transform 1 0 7681 0 1 30778
box 0 0 64 64
use contact_9  contact_9_1038
timestamp 1624494425
transform 1 0 8076 0 1 31168
box 0 0 66 74
use contact_8  contact_8_1038
timestamp 1624494425
transform 1 0 8077 0 1 31173
box 0 0 64 64
use contact_9  contact_9_1041
timestamp 1624494425
transform 1 0 8076 0 1 30773
box 0 0 66 74
use contact_8  contact_8_1041
timestamp 1624494425
transform 1 0 8077 0 1 30778
box 0 0 64 64
use contact_9  contact_9_350
timestamp 1624494425
transform 1 0 7680 0 1 31563
box 0 0 66 74
use contact_8  contact_8_350
timestamp 1624494425
transform 1 0 7681 0 1 31568
box 0 0 64 64
use contact_9  contact_9_1035
timestamp 1624494425
transform 1 0 8076 0 1 31563
box 0 0 66 74
use contact_8  contact_8_1035
timestamp 1624494425
transform 1 0 8077 0 1 31568
box 0 0 64 64
use contact_9  contact_9_346
timestamp 1624494425
transform 1 0 7680 0 1 32353
box 0 0 66 74
use contact_8  contact_8_346
timestamp 1624494425
transform 1 0 7681 0 1 32358
box 0 0 64 64
use contact_9  contact_9_348
timestamp 1624494425
transform 1 0 7680 0 1 31958
box 0 0 66 74
use contact_8  contact_8_348
timestamp 1624494425
transform 1 0 7681 0 1 31963
box 0 0 64 64
use contact_9  contact_9_1029
timestamp 1624494425
transform 1 0 8076 0 1 32353
box 0 0 66 74
use contact_8  contact_8_1029
timestamp 1624494425
transform 1 0 8077 0 1 32358
box 0 0 64 64
use contact_9  contact_9_1032
timestamp 1624494425
transform 1 0 8076 0 1 31958
box 0 0 66 74
use contact_8  contact_8_1032
timestamp 1624494425
transform 1 0 8077 0 1 31963
box 0 0 64 64
use contact_9  contact_9_344
timestamp 1624494425
transform 1 0 7680 0 1 32748
box 0 0 66 74
use contact_9  contact_9_1026
timestamp 1624494425
transform 1 0 8076 0 1 32748
box 0 0 66 74
use contact_8  contact_8_1028
timestamp 1624494425
transform 1 0 7299 0 1 32776
box 0 0 64 64
use contact_9  contact_9_1028
timestamp 1624494425
transform 1 0 7298 0 1 32771
box 0 0 66 74
use contact_8  contact_8_1027
timestamp 1624494425
transform 1 0 6867 0 1 32776
box 0 0 64 64
use contact_9  contact_9_1027
timestamp 1624494425
transform 1 0 6866 0 1 32771
box 0 0 66 74
use contact_8  contact_8_345
timestamp 1624494425
transform 1 0 6442 0 1 32776
box 0 0 64 64
use contact_9  contact_9_345
timestamp 1624494425
transform 1 0 6441 0 1 32771
box 0 0 66 74
use contact_16  contact_16_516
timestamp 1624494425
transform 1 0 5704 0 1 32868
box 0 0 66 58
use contact_16  contact_16_517
timestamp 1624494425
transform 1 0 5224 0 1 32958
box 0 0 66 58
use contact_8  contact_8_1025
timestamp 1624494425
transform 1 0 7299 0 1 33134
box 0 0 64 64
use contact_9  contact_9_1025
timestamp 1624494425
transform 1 0 7298 0 1 33129
box 0 0 66 74
use contact_8  contact_8_1024
timestamp 1624494425
transform 1 0 6867 0 1 33134
box 0 0 64 64
use contact_9  contact_9_1024
timestamp 1624494425
transform 1 0 6866 0 1 33129
box 0 0 66 74
use contact_8  contact_8_343
timestamp 1624494425
transform 1 0 6442 0 1 33192
box 0 0 64 64
use contact_9  contact_9_343
timestamp 1624494425
transform 1 0 6441 0 1 33187
box 0 0 66 74
use contact_16  contact_16_515
timestamp 1624494425
transform 1 0 4584 0 1 33232
box 0 0 66 58
use contact_16  contact_16_518
timestamp 1624494425
transform 1 0 4824 0 1 33070
box 0 0 66 58
use and3_dec  and3_dec_171
timestamp 1624494425
transform 1 0 6203 0 1 33180
box 0 -60 2072 490
use contact_8  contact_8_1022
timestamp 1624494425
transform 1 0 7299 0 1 33566
box 0 0 64 64
use contact_9  contact_9_1022
timestamp 1624494425
transform 1 0 7298 0 1 33561
box 0 0 66 74
use contact_8  contact_8_1021
timestamp 1624494425
transform 1 0 6867 0 1 33566
box 0 0 64 64
use contact_9  contact_9_1021
timestamp 1624494425
transform 1 0 6866 0 1 33561
box 0 0 66 74
use contact_8  contact_8_341
timestamp 1624494425
transform 1 0 6442 0 1 33566
box 0 0 64 64
use contact_9  contact_9_341
timestamp 1624494425
transform 1 0 6441 0 1 33561
box 0 0 66 74
use contact_16  contact_16_513
timestamp 1624494425
transform 1 0 5704 0 1 33434
box 0 0 66 58
use contact_16  contact_16_514
timestamp 1624494425
transform 1 0 5304 0 1 33344
box 0 0 66 58
use contact_16  contact_16_510
timestamp 1624494425
transform 1 0 5704 0 1 33658
box 0 0 66 58
use contact_16  contact_16_511
timestamp 1624494425
transform 1 0 5304 0 1 33748
box 0 0 66 58
use and3_dec  and3_dec_170
timestamp 1624494425
transform 1 0 6203 0 -1 33970
box 0 -60 2072 490
use contact_8  contact_8_1019
timestamp 1624494425
transform 1 0 7299 0 1 33924
box 0 0 64 64
use contact_9  contact_9_1019
timestamp 1624494425
transform 1 0 7298 0 1 33919
box 0 0 66 74
use contact_8  contact_8_1018
timestamp 1624494425
transform 1 0 6867 0 1 33924
box 0 0 64 64
use contact_9  contact_9_1018
timestamp 1624494425
transform 1 0 6866 0 1 33919
box 0 0 66 74
use contact_8  contact_8_339
timestamp 1624494425
transform 1 0 6442 0 1 33982
box 0 0 64 64
use contact_9  contact_9_339
timestamp 1624494425
transform 1 0 6441 0 1 33977
box 0 0 66 74
use contact_16  contact_16_509
timestamp 1624494425
transform 1 0 4744 0 1 34022
box 0 0 66 58
use contact_16  contact_16_512
timestamp 1624494425
transform 1 0 4664 0 1 33860
box 0 0 66 58
use contact_8  contact_8_1016
timestamp 1624494425
transform 1 0 7299 0 1 34356
box 0 0 64 64
use contact_9  contact_9_1016
timestamp 1624494425
transform 1 0 7298 0 1 34351
box 0 0 66 74
use contact_8  contact_8_1015
timestamp 1624494425
transform 1 0 6867 0 1 34356
box 0 0 64 64
use contact_9  contact_9_1015
timestamp 1624494425
transform 1 0 6866 0 1 34351
box 0 0 66 74
use contact_8  contact_8_337
timestamp 1624494425
transform 1 0 6442 0 1 34356
box 0 0 64 64
use contact_9  contact_9_337
timestamp 1624494425
transform 1 0 6441 0 1 34351
box 0 0 66 74
use contact_16  contact_16_507
timestamp 1624494425
transform 1 0 5704 0 1 34224
box 0 0 66 58
use contact_16  contact_16_508
timestamp 1624494425
transform 1 0 5304 0 1 34134
box 0 0 66 58
use and3_dec  and3_dec_168
timestamp 1624494425
transform 1 0 6203 0 -1 34760
box 0 -60 2072 490
use and3_dec  and3_dec_169
timestamp 1624494425
transform 1 0 6203 0 1 33970
box 0 -60 2072 490
use contact_16  contact_16_504
timestamp 1624494425
transform 1 0 5704 0 1 34448
box 0 0 66 58
use contact_16  contact_16_505
timestamp 1624494425
transform 1 0 5304 0 1 34538
box 0 0 66 58
use contact_16  contact_16_506
timestamp 1624494425
transform 1 0 4824 0 1 34650
box 0 0 66 58
use contact_8  contact_8_1013
timestamp 1624494425
transform 1 0 7299 0 1 34714
box 0 0 64 64
use contact_9  contact_9_1013
timestamp 1624494425
transform 1 0 7298 0 1 34709
box 0 0 66 74
use contact_8  contact_8_1012
timestamp 1624494425
transform 1 0 6867 0 1 34714
box 0 0 64 64
use contact_9  contact_9_1012
timestamp 1624494425
transform 1 0 6866 0 1 34709
box 0 0 66 74
use contact_8  contact_8_335
timestamp 1624494425
transform 1 0 6442 0 1 34772
box 0 0 64 64
use contact_9  contact_9_335
timestamp 1624494425
transform 1 0 6441 0 1 34767
box 0 0 66 74
use contact_16  contact_16_502
timestamp 1624494425
transform 1 0 5384 0 1 34924
box 0 0 66 58
use contact_16  contact_16_503
timestamp 1624494425
transform 1 0 4584 0 1 34812
box 0 0 66 58
use and3_dec  and3_dec_167
timestamp 1624494425
transform 1 0 6203 0 1 34760
box 0 -60 2072 490
use contact_8  contact_8_1010
timestamp 1624494425
transform 1 0 7299 0 1 35146
box 0 0 64 64
use contact_9  contact_9_1010
timestamp 1624494425
transform 1 0 7298 0 1 35141
box 0 0 66 74
use contact_8  contact_8_1009
timestamp 1624494425
transform 1 0 6867 0 1 35146
box 0 0 64 64
use contact_9  contact_9_1009
timestamp 1624494425
transform 1 0 6866 0 1 35141
box 0 0 66 74
use contact_8  contact_8_333
timestamp 1624494425
transform 1 0 6442 0 1 35146
box 0 0 64 64
use contact_9  contact_9_333
timestamp 1624494425
transform 1 0 6441 0 1 35141
box 0 0 66 74
use contact_16  contact_16_501
timestamp 1624494425
transform 1 0 5704 0 1 35014
box 0 0 66 58
use contact_8  contact_8_1007
timestamp 1624494425
transform 1 0 7299 0 1 35504
box 0 0 64 64
use contact_9  contact_9_1007
timestamp 1624494425
transform 1 0 7298 0 1 35499
box 0 0 66 74
use contact_8  contact_8_1006
timestamp 1624494425
transform 1 0 6867 0 1 35504
box 0 0 64 64
use contact_9  contact_9_1006
timestamp 1624494425
transform 1 0 6866 0 1 35499
box 0 0 66 74
use contact_16  contact_16_498
timestamp 1624494425
transform 1 0 5704 0 1 35238
box 0 0 66 58
use contact_16  contact_16_499
timestamp 1624494425
transform 1 0 5384 0 1 35328
box 0 0 66 58
use contact_16  contact_16_500
timestamp 1624494425
transform 1 0 4664 0 1 35440
box 0 0 66 58
use and3_dec  and3_dec_165
timestamp 1624494425
transform 1 0 6203 0 1 35550
box 0 -60 2072 490
use and3_dec  and3_dec_166
timestamp 1624494425
transform 1 0 6203 0 -1 35550
box 0 -60 2072 490
use contact_8  contact_8_331
timestamp 1624494425
transform 1 0 6442 0 1 35562
box 0 0 64 64
use contact_9  contact_9_331
timestamp 1624494425
transform 1 0 6441 0 1 35557
box 0 0 66 74
use contact_16  contact_16_496
timestamp 1624494425
transform 1 0 5384 0 1 35714
box 0 0 66 58
use contact_16  contact_16_497
timestamp 1624494425
transform 1 0 4744 0 1 35602
box 0 0 66 58
use contact_8  contact_8_1004
timestamp 1624494425
transform 1 0 7299 0 1 35936
box 0 0 64 64
use contact_9  contact_9_1004
timestamp 1624494425
transform 1 0 7298 0 1 35931
box 0 0 66 74
use contact_8  contact_8_1003
timestamp 1624494425
transform 1 0 6867 0 1 35936
box 0 0 64 64
use contact_9  contact_9_1003
timestamp 1624494425
transform 1 0 6866 0 1 35931
box 0 0 66 74
use contact_8  contact_8_329
timestamp 1624494425
transform 1 0 6442 0 1 35936
box 0 0 64 64
use contact_9  contact_9_329
timestamp 1624494425
transform 1 0 6441 0 1 35931
box 0 0 66 74
use contact_16  contact_16_492
timestamp 1624494425
transform 1 0 5704 0 1 36028
box 0 0 66 58
use contact_16  contact_16_495
timestamp 1624494425
transform 1 0 5704 0 1 35804
box 0 0 66 58
use and3_dec  and3_dec_164
timestamp 1624494425
transform 1 0 6203 0 -1 36340
box 0 -60 2072 490
use contact_9  contact_9_342
timestamp 1624494425
transform 1 0 7680 0 1 33143
box 0 0 66 74
use contact_8  contact_8_342
timestamp 1624494425
transform 1 0 7681 0 1 33148
box 0 0 64 64
use contact_8  contact_8_344
timestamp 1624494425
transform 1 0 7681 0 1 32753
box 0 0 64 64
use contact_9  contact_9_1023
timestamp 1624494425
transform 1 0 8076 0 1 33143
box 0 0 66 74
use contact_8  contact_8_1023
timestamp 1624494425
transform 1 0 8077 0 1 33148
box 0 0 64 64
use contact_8  contact_8_1026
timestamp 1624494425
transform 1 0 8077 0 1 32753
box 0 0 64 64
use contact_9  contact_9_338
timestamp 1624494425
transform 1 0 7680 0 1 33933
box 0 0 66 74
use contact_8  contact_8_338
timestamp 1624494425
transform 1 0 7681 0 1 33938
box 0 0 64 64
use contact_9  contact_9_340
timestamp 1624494425
transform 1 0 7680 0 1 33538
box 0 0 66 74
use contact_8  contact_8_340
timestamp 1624494425
transform 1 0 7681 0 1 33543
box 0 0 64 64
use contact_9  contact_9_1017
timestamp 1624494425
transform 1 0 8076 0 1 33933
box 0 0 66 74
use contact_8  contact_8_1017
timestamp 1624494425
transform 1 0 8077 0 1 33938
box 0 0 64 64
use contact_9  contact_9_1020
timestamp 1624494425
transform 1 0 8076 0 1 33538
box 0 0 66 74
use contact_8  contact_8_1020
timestamp 1624494425
transform 1 0 8077 0 1 33543
box 0 0 64 64
use contact_9  contact_9_336
timestamp 1624494425
transform 1 0 7680 0 1 34328
box 0 0 66 74
use contact_8  contact_8_336
timestamp 1624494425
transform 1 0 7681 0 1 34333
box 0 0 64 64
use contact_9  contact_9_1014
timestamp 1624494425
transform 1 0 8076 0 1 34328
box 0 0 66 74
use contact_8  contact_8_1014
timestamp 1624494425
transform 1 0 8077 0 1 34333
box 0 0 64 64
use contact_9  contact_9_332
timestamp 1624494425
transform 1 0 7680 0 1 35118
box 0 0 66 74
use contact_8  contact_8_332
timestamp 1624494425
transform 1 0 7681 0 1 35123
box 0 0 64 64
use contact_9  contact_9_334
timestamp 1624494425
transform 1 0 7680 0 1 34723
box 0 0 66 74
use contact_8  contact_8_334
timestamp 1624494425
transform 1 0 7681 0 1 34728
box 0 0 64 64
use contact_9  contact_9_1008
timestamp 1624494425
transform 1 0 8076 0 1 35118
box 0 0 66 74
use contact_8  contact_8_1008
timestamp 1624494425
transform 1 0 8077 0 1 35123
box 0 0 64 64
use contact_9  contact_9_1011
timestamp 1624494425
transform 1 0 8076 0 1 34723
box 0 0 66 74
use contact_8  contact_8_1011
timestamp 1624494425
transform 1 0 8077 0 1 34728
box 0 0 64 64
use contact_9  contact_9_330
timestamp 1624494425
transform 1 0 7680 0 1 35513
box 0 0 66 74
use contact_8  contact_8_330
timestamp 1624494425
transform 1 0 7681 0 1 35518
box 0 0 64 64
use contact_9  contact_9_1005
timestamp 1624494425
transform 1 0 8076 0 1 35513
box 0 0 66 74
use contact_8  contact_8_1005
timestamp 1624494425
transform 1 0 8077 0 1 35518
box 0 0 64 64
use contact_9  contact_9_328
timestamp 1624494425
transform 1 0 7680 0 1 35908
box 0 0 66 74
use contact_8  contact_8_328
timestamp 1624494425
transform 1 0 7681 0 1 35913
box 0 0 64 64
use contact_9  contact_9_1002
timestamp 1624494425
transform 1 0 8076 0 1 35908
box 0 0 66 74
use contact_8  contact_8_1002
timestamp 1624494425
transform 1 0 8077 0 1 35913
box 0 0 64 64
use contact_8  contact_8_1001
timestamp 1624494425
transform 1 0 7299 0 1 36294
box 0 0 64 64
use contact_9  contact_9_1001
timestamp 1624494425
transform 1 0 7298 0 1 36289
box 0 0 66 74
use contact_8  contact_8_1000
timestamp 1624494425
transform 1 0 6867 0 1 36294
box 0 0 64 64
use contact_9  contact_9_1000
timestamp 1624494425
transform 1 0 6866 0 1 36289
box 0 0 66 74
use contact_16  contact_16_493
timestamp 1624494425
transform 1 0 5384 0 1 36118
box 0 0 66 58
use contact_16  contact_16_494
timestamp 1624494425
transform 1 0 4824 0 1 36230
box 0 0 66 58
use contact_8  contact_8_327
timestamp 1624494425
transform 1 0 6442 0 1 36352
box 0 0 64 64
use contact_9  contact_9_327
timestamp 1624494425
transform 1 0 6441 0 1 36347
box 0 0 66 74
use contact_16  contact_16_490
timestamp 1624494425
transform 1 0 5464 0 1 36504
box 0 0 66 58
use contact_16  contact_16_491
timestamp 1624494425
transform 1 0 4584 0 1 36392
box 0 0 66 58
use and3_dec  and3_dec_163
timestamp 1624494425
transform 1 0 6203 0 1 36340
box 0 -60 2072 490
use contact_8  contact_8_998
timestamp 1624494425
transform 1 0 7299 0 1 36726
box 0 0 64 64
use contact_9  contact_9_998
timestamp 1624494425
transform 1 0 7298 0 1 36721
box 0 0 66 74
use contact_8  contact_8_997
timestamp 1624494425
transform 1 0 6867 0 1 36726
box 0 0 64 64
use contact_9  contact_9_997
timestamp 1624494425
transform 1 0 6866 0 1 36721
box 0 0 66 74
use contact_8  contact_8_325
timestamp 1624494425
transform 1 0 6442 0 1 36726
box 0 0 64 64
use contact_9  contact_9_325
timestamp 1624494425
transform 1 0 6441 0 1 36721
box 0 0 66 74
use contact_16  contact_16_486
timestamp 1624494425
transform 1 0 5704 0 1 36818
box 0 0 66 58
use contact_16  contact_16_489
timestamp 1624494425
transform 1 0 5704 0 1 36594
box 0 0 66 58
use contact_8  contact_8_995
timestamp 1624494425
transform 1 0 7299 0 1 37084
box 0 0 64 64
use contact_9  contact_9_995
timestamp 1624494425
transform 1 0 7298 0 1 37079
box 0 0 66 74
use contact_8  contact_8_994
timestamp 1624494425
transform 1 0 6867 0 1 37084
box 0 0 64 64
use contact_9  contact_9_994
timestamp 1624494425
transform 1 0 6866 0 1 37079
box 0 0 66 74
use contact_16  contact_16_487
timestamp 1624494425
transform 1 0 5464 0 1 36908
box 0 0 66 58
use contact_16  contact_16_488
timestamp 1624494425
transform 1 0 4664 0 1 37020
box 0 0 66 58
use and3_dec  and3_dec_161
timestamp 1624494425
transform 1 0 6203 0 1 37130
box 0 -60 2072 490
use and3_dec  and3_dec_162
timestamp 1624494425
transform 1 0 6203 0 -1 37130
box 0 -60 2072 490
use contact_8  contact_8_323
timestamp 1624494425
transform 1 0 6442 0 1 37142
box 0 0 64 64
use contact_9  contact_9_323
timestamp 1624494425
transform 1 0 6441 0 1 37137
box 0 0 66 74
use contact_16  contact_16_483
timestamp 1624494425
transform 1 0 5704 0 1 37384
box 0 0 66 58
use contact_16  contact_16_484
timestamp 1624494425
transform 1 0 5464 0 1 37294
box 0 0 66 58
use contact_16  contact_16_485
timestamp 1624494425
transform 1 0 4744 0 1 37182
box 0 0 66 58
use contact_8  contact_8_992
timestamp 1624494425
transform 1 0 7299 0 1 37516
box 0 0 64 64
use contact_9  contact_9_992
timestamp 1624494425
transform 1 0 7298 0 1 37511
box 0 0 66 74
use contact_8  contact_8_991
timestamp 1624494425
transform 1 0 6867 0 1 37516
box 0 0 64 64
use contact_9  contact_9_991
timestamp 1624494425
transform 1 0 6866 0 1 37511
box 0 0 66 74
use contact_8  contact_8_321
timestamp 1624494425
transform 1 0 6442 0 1 37516
box 0 0 64 64
use contact_9  contact_9_321
timestamp 1624494425
transform 1 0 6441 0 1 37511
box 0 0 66 74
use contact_16  contact_16_480
timestamp 1624494425
transform 1 0 5704 0 1 37608
box 0 0 66 58
use and3_dec  and3_dec_160
timestamp 1624494425
transform 1 0 6203 0 -1 37920
box 0 -60 2072 490
use contact_8  contact_8_989
timestamp 1624494425
transform 1 0 7299 0 1 37874
box 0 0 64 64
use contact_9  contact_9_989
timestamp 1624494425
transform 1 0 7298 0 1 37869
box 0 0 66 74
use contact_8  contact_8_988
timestamp 1624494425
transform 1 0 6867 0 1 37874
box 0 0 64 64
use contact_9  contact_9_988
timestamp 1624494425
transform 1 0 6866 0 1 37869
box 0 0 66 74
use contact_8  contact_8_319
timestamp 1624494425
transform 1 0 6442 0 1 37932
box 0 0 64 64
use contact_9  contact_9_319
timestamp 1624494425
transform 1 0 6441 0 1 37927
box 0 0 66 74
use contact_16  contact_16_481
timestamp 1624494425
transform 1 0 5464 0 1 37698
box 0 0 66 58
use contact_16  contact_16_482
timestamp 1624494425
transform 1 0 4824 0 1 37810
box 0 0 66 58
use contact_16  contact_16_477
timestamp 1624494425
transform 1 0 5784 0 1 38174
box 0 0 66 58
use contact_16  contact_16_478
timestamp 1624494425
transform 1 0 4904 0 1 38084
box 0 0 66 58
use contact_16  contact_16_479
timestamp 1624494425
transform 1 0 4584 0 1 37972
box 0 0 66 58
use and3_dec  and3_dec_158
timestamp 1624494425
transform 1 0 6203 0 -1 38710
box 0 -60 2072 490
use and3_dec  and3_dec_159
timestamp 1624494425
transform 1 0 6203 0 1 37920
box 0 -60 2072 490
use contact_8  contact_8_986
timestamp 1624494425
transform 1 0 7299 0 1 38306
box 0 0 64 64
use contact_9  contact_9_986
timestamp 1624494425
transform 1 0 7298 0 1 38301
box 0 0 66 74
use contact_8  contact_8_985
timestamp 1624494425
transform 1 0 6867 0 1 38306
box 0 0 64 64
use contact_9  contact_9_985
timestamp 1624494425
transform 1 0 6866 0 1 38301
box 0 0 66 74
use contact_8  contact_8_317
timestamp 1624494425
transform 1 0 6442 0 1 38306
box 0 0 64 64
use contact_9  contact_9_317
timestamp 1624494425
transform 1 0 6441 0 1 38301
box 0 0 66 74
use contact_16  contact_16_474
timestamp 1624494425
transform 1 0 5784 0 1 38398
box 0 0 66 58
use contact_16  contact_16_475
timestamp 1624494425
transform 1 0 4904 0 1 38488
box 0 0 66 58
use contact_8  contact_8_983
timestamp 1624494425
transform 1 0 7299 0 1 38664
box 0 0 64 64
use contact_9  contact_9_983
timestamp 1624494425
transform 1 0 7298 0 1 38659
box 0 0 66 74
use contact_8  contact_8_982
timestamp 1624494425
transform 1 0 6867 0 1 38664
box 0 0 64 64
use contact_9  contact_9_982
timestamp 1624494425
transform 1 0 6866 0 1 38659
box 0 0 66 74
use contact_8  contact_8_315
timestamp 1624494425
transform 1 0 6442 0 1 38722
box 0 0 64 64
use contact_9  contact_9_315
timestamp 1624494425
transform 1 0 6441 0 1 38717
box 0 0 66 74
use contact_16  contact_16_473
timestamp 1624494425
transform 1 0 4744 0 1 38762
box 0 0 66 58
use contact_16  contact_16_476
timestamp 1624494425
transform 1 0 4664 0 1 38600
box 0 0 66 58
use and3_dec  and3_dec_157
timestamp 1624494425
transform 1 0 6203 0 1 38710
box 0 -60 2072 490
use contact_16  contact_16_471
timestamp 1624494425
transform 1 0 5784 0 1 38964
box 0 0 66 58
use contact_16  contact_16_472
timestamp 1624494425
transform 1 0 4904 0 1 38874
box 0 0 66 58
use contact_8  contact_8_980
timestamp 1624494425
transform 1 0 7299 0 1 39096
box 0 0 64 64
use contact_9  contact_9_980
timestamp 1624494425
transform 1 0 7298 0 1 39091
box 0 0 66 74
use contact_8  contact_8_979
timestamp 1624494425
transform 1 0 6867 0 1 39096
box 0 0 64 64
use contact_9  contact_9_979
timestamp 1624494425
transform 1 0 6866 0 1 39091
box 0 0 66 74
use contact_8  contact_8_313
timestamp 1624494425
transform 1 0 6442 0 1 39096
box 0 0 64 64
use contact_9  contact_9_313
timestamp 1624494425
transform 1 0 6441 0 1 39091
box 0 0 66 74
use contact_16  contact_16_468
timestamp 1624494425
transform 1 0 5784 0 1 39188
box 0 0 66 58
use contact_16  contact_16_469
timestamp 1624494425
transform 1 0 4904 0 1 39278
box 0 0 66 58
use and3_dec  and3_dec_156
timestamp 1624494425
transform 1 0 6203 0 -1 39500
box 0 -60 2072 490
use contact_9  contact_9_326
timestamp 1624494425
transform 1 0 7680 0 1 36303
box 0 0 66 74
use contact_8  contact_8_326
timestamp 1624494425
transform 1 0 7681 0 1 36308
box 0 0 64 64
use contact_9  contact_9_999
timestamp 1624494425
transform 1 0 8076 0 1 36303
box 0 0 66 74
use contact_8  contact_8_999
timestamp 1624494425
transform 1 0 8077 0 1 36308
box 0 0 64 64
use contact_9  contact_9_322
timestamp 1624494425
transform 1 0 7680 0 1 37093
box 0 0 66 74
use contact_8  contact_8_322
timestamp 1624494425
transform 1 0 7681 0 1 37098
box 0 0 64 64
use contact_9  contact_9_324
timestamp 1624494425
transform 1 0 7680 0 1 36698
box 0 0 66 74
use contact_8  contact_8_324
timestamp 1624494425
transform 1 0 7681 0 1 36703
box 0 0 64 64
use contact_9  contact_9_993
timestamp 1624494425
transform 1 0 8076 0 1 37093
box 0 0 66 74
use contact_8  contact_8_993
timestamp 1624494425
transform 1 0 8077 0 1 37098
box 0 0 64 64
use contact_9  contact_9_996
timestamp 1624494425
transform 1 0 8076 0 1 36698
box 0 0 66 74
use contact_8  contact_8_996
timestamp 1624494425
transform 1 0 8077 0 1 36703
box 0 0 64 64
use contact_9  contact_9_318
timestamp 1624494425
transform 1 0 7680 0 1 37883
box 0 0 66 74
use contact_8  contact_8_318
timestamp 1624494425
transform 1 0 7681 0 1 37888
box 0 0 64 64
use contact_9  contact_9_320
timestamp 1624494425
transform 1 0 7680 0 1 37488
box 0 0 66 74
use contact_8  contact_8_320
timestamp 1624494425
transform 1 0 7681 0 1 37493
box 0 0 64 64
use contact_9  contact_9_987
timestamp 1624494425
transform 1 0 8076 0 1 37883
box 0 0 66 74
use contact_8  contact_8_987
timestamp 1624494425
transform 1 0 8077 0 1 37888
box 0 0 64 64
use contact_9  contact_9_990
timestamp 1624494425
transform 1 0 8076 0 1 37488
box 0 0 66 74
use contact_8  contact_8_990
timestamp 1624494425
transform 1 0 8077 0 1 37493
box 0 0 64 64
use contact_9  contact_9_316
timestamp 1624494425
transform 1 0 7680 0 1 38278
box 0 0 66 74
use contact_8  contact_8_316
timestamp 1624494425
transform 1 0 7681 0 1 38283
box 0 0 64 64
use contact_9  contact_9_984
timestamp 1624494425
transform 1 0 8076 0 1 38278
box 0 0 66 74
use contact_8  contact_8_984
timestamp 1624494425
transform 1 0 8077 0 1 38283
box 0 0 64 64
use contact_9  contact_9_312
timestamp 1624494425
transform 1 0 7680 0 1 39068
box 0 0 66 74
use contact_8  contact_8_312
timestamp 1624494425
transform 1 0 7681 0 1 39073
box 0 0 64 64
use contact_9  contact_9_314
timestamp 1624494425
transform 1 0 7680 0 1 38673
box 0 0 66 74
use contact_8  contact_8_314
timestamp 1624494425
transform 1 0 7681 0 1 38678
box 0 0 64 64
use contact_9  contact_9_978
timestamp 1624494425
transform 1 0 8076 0 1 39068
box 0 0 66 74
use contact_8  contact_8_978
timestamp 1624494425
transform 1 0 8077 0 1 39073
box 0 0 64 64
use contact_9  contact_9_981
timestamp 1624494425
transform 1 0 8076 0 1 38673
box 0 0 66 74
use contact_8  contact_8_981
timestamp 1624494425
transform 1 0 8077 0 1 38678
box 0 0 64 64
use contact_8  contact_8_977
timestamp 1624494425
transform 1 0 7299 0 1 39454
box 0 0 64 64
use contact_9  contact_9_977
timestamp 1624494425
transform 1 0 7298 0 1 39449
box 0 0 66 74
use contact_8  contact_8_976
timestamp 1624494425
transform 1 0 6867 0 1 39454
box 0 0 64 64
use contact_9  contact_9_976
timestamp 1624494425
transform 1 0 6866 0 1 39449
box 0 0 66 74
use contact_8  contact_8_311
timestamp 1624494425
transform 1 0 6442 0 1 39512
box 0 0 64 64
use contact_9  contact_9_311
timestamp 1624494425
transform 1 0 6441 0 1 39507
box 0 0 66 74
use contact_16  contact_16_467
timestamp 1624494425
transform 1 0 4584 0 1 39552
box 0 0 66 58
use contact_16  contact_16_470
timestamp 1624494425
transform 1 0 4824 0 1 39390
box 0 0 66 58
use contact_16  contact_16_465
timestamp 1624494425
transform 1 0 5784 0 1 39754
box 0 0 66 58
use contact_16  contact_16_466
timestamp 1624494425
transform 1 0 4984 0 1 39664
box 0 0 66 58
use and3_dec  and3_dec_154
timestamp 1624494425
transform 1 0 6203 0 -1 40290
box 0 -60 2072 490
use and3_dec  and3_dec_155
timestamp 1624494425
transform 1 0 6203 0 1 39500
box 0 -60 2072 490
use contact_8  contact_8_974
timestamp 1624494425
transform 1 0 7299 0 1 39886
box 0 0 64 64
use contact_9  contact_9_974
timestamp 1624494425
transform 1 0 7298 0 1 39881
box 0 0 66 74
use contact_8  contact_8_973
timestamp 1624494425
transform 1 0 6867 0 1 39886
box 0 0 64 64
use contact_9  contact_9_973
timestamp 1624494425
transform 1 0 6866 0 1 39881
box 0 0 66 74
use contact_8  contact_8_309
timestamp 1624494425
transform 1 0 6442 0 1 39886
box 0 0 64 64
use contact_9  contact_9_309
timestamp 1624494425
transform 1 0 6441 0 1 39881
box 0 0 66 74
use contact_16  contact_16_462
timestamp 1624494425
transform 1 0 5784 0 1 39978
box 0 0 66 58
use contact_16  contact_16_463
timestamp 1624494425
transform 1 0 4984 0 1 40068
box 0 0 66 58
use contact_8  contact_8_971
timestamp 1624494425
transform 1 0 7299 0 1 40244
box 0 0 64 64
use contact_9  contact_9_971
timestamp 1624494425
transform 1 0 7298 0 1 40239
box 0 0 66 74
use contact_8  contact_8_970
timestamp 1624494425
transform 1 0 6867 0 1 40244
box 0 0 64 64
use contact_9  contact_9_970
timestamp 1624494425
transform 1 0 6866 0 1 40239
box 0 0 66 74
use contact_8  contact_8_307
timestamp 1624494425
transform 1 0 6442 0 1 40302
box 0 0 64 64
use contact_9  contact_9_307
timestamp 1624494425
transform 1 0 6441 0 1 40297
box 0 0 66 74
use contact_16  contact_16_461
timestamp 1624494425
transform 1 0 4744 0 1 40342
box 0 0 66 58
use contact_16  contact_16_464
timestamp 1624494425
transform 1 0 4664 0 1 40180
box 0 0 66 58
use and3_dec  and3_dec_153
timestamp 1624494425
transform 1 0 6203 0 1 40290
box 0 -60 2072 490
use contact_8  contact_8_968
timestamp 1624494425
transform 1 0 7299 0 1 40676
box 0 0 64 64
use contact_9  contact_9_968
timestamp 1624494425
transform 1 0 7298 0 1 40671
box 0 0 66 74
use contact_8  contact_8_967
timestamp 1624494425
transform 1 0 6867 0 1 40676
box 0 0 64 64
use contact_9  contact_9_967
timestamp 1624494425
transform 1 0 6866 0 1 40671
box 0 0 66 74
use contact_8  contact_8_305
timestamp 1624494425
transform 1 0 6442 0 1 40676
box 0 0 64 64
use contact_9  contact_9_305
timestamp 1624494425
transform 1 0 6441 0 1 40671
box 0 0 66 74
use contact_16  contact_16_459
timestamp 1624494425
transform 1 0 5784 0 1 40544
box 0 0 66 58
use contact_16  contact_16_460
timestamp 1624494425
transform 1 0 4984 0 1 40454
box 0 0 66 58
use contact_16  contact_16_456
timestamp 1624494425
transform 1 0 5784 0 1 40768
box 0 0 66 58
use contact_16  contact_16_457
timestamp 1624494425
transform 1 0 4984 0 1 40858
box 0 0 66 58
use and3_dec  and3_dec_152
timestamp 1624494425
transform 1 0 6203 0 -1 41080
box 0 -60 2072 490
use contact_8  contact_8_965
timestamp 1624494425
transform 1 0 7299 0 1 41034
box 0 0 64 64
use contact_9  contact_9_965
timestamp 1624494425
transform 1 0 7298 0 1 41029
box 0 0 66 74
use contact_8  contact_8_964
timestamp 1624494425
transform 1 0 6867 0 1 41034
box 0 0 64 64
use contact_9  contact_9_964
timestamp 1624494425
transform 1 0 6866 0 1 41029
box 0 0 66 74
use contact_8  contact_8_303
timestamp 1624494425
transform 1 0 6442 0 1 41092
box 0 0 64 64
use contact_9  contact_9_303
timestamp 1624494425
transform 1 0 6441 0 1 41087
box 0 0 66 74
use contact_16  contact_16_455
timestamp 1624494425
transform 1 0 4584 0 1 41132
box 0 0 66 58
use contact_16  contact_16_458
timestamp 1624494425
transform 1 0 4824 0 1 40970
box 0 0 66 58
use contact_8  contact_8_962
timestamp 1624494425
transform 1 0 7299 0 1 41466
box 0 0 64 64
use contact_9  contact_9_962
timestamp 1624494425
transform 1 0 7298 0 1 41461
box 0 0 66 74
use contact_8  contact_8_961
timestamp 1624494425
transform 1 0 6867 0 1 41466
box 0 0 64 64
use contact_9  contact_9_961
timestamp 1624494425
transform 1 0 6866 0 1 41461
box 0 0 66 74
use contact_8  contact_8_301
timestamp 1624494425
transform 1 0 6442 0 1 41466
box 0 0 64 64
use contact_9  contact_9_301
timestamp 1624494425
transform 1 0 6441 0 1 41461
box 0 0 66 74
use contact_16  contact_16_453
timestamp 1624494425
transform 1 0 5784 0 1 41334
box 0 0 66 58
use contact_16  contact_16_454
timestamp 1624494425
transform 1 0 5064 0 1 41244
box 0 0 66 58
use and3_dec  and3_dec_150
timestamp 1624494425
transform 1 0 6203 0 -1 41870
box 0 -60 2072 490
use and3_dec  and3_dec_151
timestamp 1624494425
transform 1 0 6203 0 1 41080
box 0 -60 2072 490
use contact_16  contact_16_450
timestamp 1624494425
transform 1 0 5784 0 1 41558
box 0 0 66 58
use contact_16  contact_16_451
timestamp 1624494425
transform 1 0 5064 0 1 41648
box 0 0 66 58
use contact_16  contact_16_452
timestamp 1624494425
transform 1 0 4664 0 1 41760
box 0 0 66 58
use contact_8  contact_8_959
timestamp 1624494425
transform 1 0 7299 0 1 41824
box 0 0 64 64
use contact_9  contact_9_959
timestamp 1624494425
transform 1 0 7298 0 1 41819
box 0 0 66 74
use contact_8  contact_8_958
timestamp 1624494425
transform 1 0 6867 0 1 41824
box 0 0 64 64
use contact_9  contact_9_958
timestamp 1624494425
transform 1 0 6866 0 1 41819
box 0 0 66 74
use contact_8  contact_8_299
timestamp 1624494425
transform 1 0 6442 0 1 41882
box 0 0 64 64
use contact_9  contact_9_299
timestamp 1624494425
transform 1 0 6441 0 1 41877
box 0 0 66 74
use contact_16  contact_16_448
timestamp 1624494425
transform 1 0 5064 0 1 42034
box 0 0 66 58
use contact_16  contact_16_449
timestamp 1624494425
transform 1 0 4744 0 1 41922
box 0 0 66 58
use and3_dec  and3_dec_149
timestamp 1624494425
transform 1 0 6203 0 1 41870
box 0 -60 2072 490
use contact_8  contact_8_956
timestamp 1624494425
transform 1 0 7299 0 1 42256
box 0 0 64 64
use contact_9  contact_9_956
timestamp 1624494425
transform 1 0 7298 0 1 42251
box 0 0 66 74
use contact_8  contact_8_955
timestamp 1624494425
transform 1 0 6867 0 1 42256
box 0 0 64 64
use contact_9  contact_9_955
timestamp 1624494425
transform 1 0 6866 0 1 42251
box 0 0 66 74
use contact_8  contact_8_297
timestamp 1624494425
transform 1 0 6442 0 1 42256
box 0 0 64 64
use contact_9  contact_9_297
timestamp 1624494425
transform 1 0 6441 0 1 42251
box 0 0 66 74
use contact_16  contact_16_447
timestamp 1624494425
transform 1 0 5784 0 1 42124
box 0 0 66 58
use contact_16  contact_16_444
timestamp 1624494425
transform 1 0 5784 0 1 42348
box 0 0 66 58
use contact_16  contact_16_445
timestamp 1624494425
transform 1 0 5064 0 1 42438
box 0 0 66 58
use contact_16  contact_16_446
timestamp 1624494425
transform 1 0 4824 0 1 42550
box 0 0 66 58
use and3_dec  and3_dec_148
timestamp 1624494425
transform 1 0 6203 0 -1 42660
box 0 -60 2072 490
use contact_9  contact_9_308
timestamp 1624494425
transform 1 0 7680 0 1 39858
box 0 0 66 74
use contact_8  contact_8_308
timestamp 1624494425
transform 1 0 7681 0 1 39863
box 0 0 64 64
use contact_9  contact_9_310
timestamp 1624494425
transform 1 0 7680 0 1 39463
box 0 0 66 74
use contact_8  contact_8_310
timestamp 1624494425
transform 1 0 7681 0 1 39468
box 0 0 64 64
use contact_9  contact_9_972
timestamp 1624494425
transform 1 0 8076 0 1 39858
box 0 0 66 74
use contact_8  contact_8_972
timestamp 1624494425
transform 1 0 8077 0 1 39863
box 0 0 64 64
use contact_9  contact_9_975
timestamp 1624494425
transform 1 0 8076 0 1 39463
box 0 0 66 74
use contact_8  contact_8_975
timestamp 1624494425
transform 1 0 8077 0 1 39468
box 0 0 64 64
use contact_9  contact_9_306
timestamp 1624494425
transform 1 0 7680 0 1 40253
box 0 0 66 74
use contact_8  contact_8_306
timestamp 1624494425
transform 1 0 7681 0 1 40258
box 0 0 64 64
use contact_9  contact_9_969
timestamp 1624494425
transform 1 0 8076 0 1 40253
box 0 0 66 74
use contact_8  contact_8_969
timestamp 1624494425
transform 1 0 8077 0 1 40258
box 0 0 64 64
use contact_9  contact_9_302
timestamp 1624494425
transform 1 0 7680 0 1 41043
box 0 0 66 74
use contact_8  contact_8_302
timestamp 1624494425
transform 1 0 7681 0 1 41048
box 0 0 64 64
use contact_9  contact_9_304
timestamp 1624494425
transform 1 0 7680 0 1 40648
box 0 0 66 74
use contact_8  contact_8_304
timestamp 1624494425
transform 1 0 7681 0 1 40653
box 0 0 64 64
use contact_9  contact_9_963
timestamp 1624494425
transform 1 0 8076 0 1 41043
box 0 0 66 74
use contact_8  contact_8_963
timestamp 1624494425
transform 1 0 8077 0 1 41048
box 0 0 64 64
use contact_9  contact_9_966
timestamp 1624494425
transform 1 0 8076 0 1 40648
box 0 0 66 74
use contact_8  contact_8_966
timestamp 1624494425
transform 1 0 8077 0 1 40653
box 0 0 64 64
use contact_9  contact_9_300
timestamp 1624494425
transform 1 0 7680 0 1 41438
box 0 0 66 74
use contact_8  contact_8_300
timestamp 1624494425
transform 1 0 7681 0 1 41443
box 0 0 64 64
use contact_9  contact_9_960
timestamp 1624494425
transform 1 0 8076 0 1 41438
box 0 0 66 74
use contact_8  contact_8_960
timestamp 1624494425
transform 1 0 8077 0 1 41443
box 0 0 64 64
use contact_9  contact_9_296
timestamp 1624494425
transform 1 0 7680 0 1 42228
box 0 0 66 74
use contact_8  contact_8_296
timestamp 1624494425
transform 1 0 7681 0 1 42233
box 0 0 64 64
use contact_9  contact_9_298
timestamp 1624494425
transform 1 0 7680 0 1 41833
box 0 0 66 74
use contact_8  contact_8_298
timestamp 1624494425
transform 1 0 7681 0 1 41838
box 0 0 64 64
use contact_9  contact_9_954
timestamp 1624494425
transform 1 0 8076 0 1 42228
box 0 0 66 74
use contact_8  contact_8_954
timestamp 1624494425
transform 1 0 8077 0 1 42233
box 0 0 64 64
use contact_9  contact_9_957
timestamp 1624494425
transform 1 0 8076 0 1 41833
box 0 0 66 74
use contact_8  contact_8_957
timestamp 1624494425
transform 1 0 8077 0 1 41838
box 0 0 64 64
use contact_8  contact_8_953
timestamp 1624494425
transform 1 0 7299 0 1 42614
box 0 0 64 64
use contact_9  contact_9_953
timestamp 1624494425
transform 1 0 7298 0 1 42609
box 0 0 66 74
use contact_8  contact_8_952
timestamp 1624494425
transform 1 0 6867 0 1 42614
box 0 0 64 64
use contact_9  contact_9_952
timestamp 1624494425
transform 1 0 6866 0 1 42609
box 0 0 66 74
use contact_8  contact_8_295
timestamp 1624494425
transform 1 0 6442 0 1 42672
box 0 0 64 64
use contact_9  contact_9_295
timestamp 1624494425
transform 1 0 6441 0 1 42667
box 0 0 66 74
use contact_16  contact_16_442
timestamp 1624494425
transform 1 0 5144 0 1 42824
box 0 0 66 58
use contact_16  contact_16_443
timestamp 1624494425
transform 1 0 4584 0 1 42712
box 0 0 66 58
use contact_8  contact_8_950
timestamp 1624494425
transform 1 0 7299 0 1 43046
box 0 0 64 64
use contact_9  contact_9_950
timestamp 1624494425
transform 1 0 7298 0 1 43041
box 0 0 66 74
use contact_8  contact_8_949
timestamp 1624494425
transform 1 0 6867 0 1 43046
box 0 0 64 64
use contact_9  contact_9_949
timestamp 1624494425
transform 1 0 6866 0 1 43041
box 0 0 66 74
use contact_8  contact_8_293
timestamp 1624494425
transform 1 0 6442 0 1 43046
box 0 0 64 64
use contact_9  contact_9_293
timestamp 1624494425
transform 1 0 6441 0 1 43041
box 0 0 66 74
use contact_16  contact_16_438
timestamp 1624494425
transform 1 0 5784 0 1 43138
box 0 0 66 58
use contact_16  contact_16_441
timestamp 1624494425
transform 1 0 5784 0 1 42914
box 0 0 66 58
use and3_dec  and3_dec_146
timestamp 1624494425
transform 1 0 6203 0 -1 43450
box 0 -60 2072 490
use and3_dec  and3_dec_147
timestamp 1624494425
transform 1 0 6203 0 1 42660
box 0 -60 2072 490
use contact_8  contact_8_947
timestamp 1624494425
transform 1 0 7299 0 1 43404
box 0 0 64 64
use contact_9  contact_9_947
timestamp 1624494425
transform 1 0 7298 0 1 43399
box 0 0 66 74
use contact_8  contact_8_946
timestamp 1624494425
transform 1 0 6867 0 1 43404
box 0 0 64 64
use contact_9  contact_9_946
timestamp 1624494425
transform 1 0 6866 0 1 43399
box 0 0 66 74
use contact_16  contact_16_439
timestamp 1624494425
transform 1 0 5144 0 1 43228
box 0 0 66 58
use contact_16  contact_16_440
timestamp 1624494425
transform 1 0 4664 0 1 43340
box 0 0 66 58
use contact_8  contact_8_291
timestamp 1624494425
transform 1 0 6442 0 1 43462
box 0 0 64 64
use contact_9  contact_9_291
timestamp 1624494425
transform 1 0 6441 0 1 43457
box 0 0 66 74
use contact_16  contact_16_436
timestamp 1624494425
transform 1 0 5144 0 1 43614
box 0 0 66 58
use contact_16  contact_16_437
timestamp 1624494425
transform 1 0 4744 0 1 43502
box 0 0 66 58
use and3_dec  and3_dec_145
timestamp 1624494425
transform 1 0 6203 0 1 43450
box 0 -60 2072 490
use contact_8  contact_8_944
timestamp 1624494425
transform 1 0 7299 0 1 43836
box 0 0 64 64
use contact_9  contact_9_944
timestamp 1624494425
transform 1 0 7298 0 1 43831
box 0 0 66 74
use contact_8  contact_8_943
timestamp 1624494425
transform 1 0 6867 0 1 43836
box 0 0 64 64
use contact_9  contact_9_943
timestamp 1624494425
transform 1 0 6866 0 1 43831
box 0 0 66 74
use contact_8  contact_8_289
timestamp 1624494425
transform 1 0 6442 0 1 43836
box 0 0 64 64
use contact_9  contact_9_289
timestamp 1624494425
transform 1 0 6441 0 1 43831
box 0 0 66 74
use contact_16  contact_16_432
timestamp 1624494425
transform 1 0 5784 0 1 43928
box 0 0 66 58
use contact_16  contact_16_435
timestamp 1624494425
transform 1 0 5784 0 1 43704
box 0 0 66 58
use contact_8  contact_8_941
timestamp 1624494425
transform 1 0 7299 0 1 44194
box 0 0 64 64
use contact_9  contact_9_941
timestamp 1624494425
transform 1 0 7298 0 1 44189
box 0 0 66 74
use contact_8  contact_8_940
timestamp 1624494425
transform 1 0 6867 0 1 44194
box 0 0 64 64
use contact_9  contact_9_940
timestamp 1624494425
transform 1 0 6866 0 1 44189
box 0 0 66 74
use contact_16  contact_16_433
timestamp 1624494425
transform 1 0 5144 0 1 44018
box 0 0 66 58
use contact_16  contact_16_434
timestamp 1624494425
transform 1 0 4824 0 1 44130
box 0 0 66 58
use and3_dec  and3_dec_143
timestamp 1624494425
transform 1 0 6203 0 1 44240
box 0 -60 2072 490
use and3_dec  and3_dec_144
timestamp 1624494425
transform 1 0 6203 0 -1 44240
box 0 -60 2072 490
use contact_8  contact_8_287
timestamp 1624494425
transform 1 0 6442 0 1 44252
box 0 0 64 64
use contact_9  contact_9_287
timestamp 1624494425
transform 1 0 6441 0 1 44247
box 0 0 66 74
use contact_16  contact_16_429
timestamp 1624494425
transform 1 0 5784 0 1 44494
box 0 0 66 58
use contact_16  contact_16_430
timestamp 1624494425
transform 1 0 5224 0 1 44404
box 0 0 66 58
use contact_16  contact_16_431
timestamp 1624494425
transform 1 0 4584 0 1 44292
box 0 0 66 58
use contact_8  contact_8_938
timestamp 1624494425
transform 1 0 7299 0 1 44626
box 0 0 64 64
use contact_9  contact_9_938
timestamp 1624494425
transform 1 0 7298 0 1 44621
box 0 0 66 74
use contact_8  contact_8_937
timestamp 1624494425
transform 1 0 6867 0 1 44626
box 0 0 64 64
use contact_9  contact_9_937
timestamp 1624494425
transform 1 0 6866 0 1 44621
box 0 0 66 74
use contact_8  contact_8_285
timestamp 1624494425
transform 1 0 6442 0 1 44626
box 0 0 64 64
use contact_9  contact_9_285
timestamp 1624494425
transform 1 0 6441 0 1 44621
box 0 0 66 74
use contact_16  contact_16_426
timestamp 1624494425
transform 1 0 5784 0 1 44718
box 0 0 66 58
use and3_dec  and3_dec_142
timestamp 1624494425
transform 1 0 6203 0 -1 45030
box 0 -60 2072 490
use contact_8  contact_8_935
timestamp 1624494425
transform 1 0 7299 0 1 44984
box 0 0 64 64
use contact_9  contact_9_935
timestamp 1624494425
transform 1 0 7298 0 1 44979
box 0 0 66 74
use contact_8  contact_8_934
timestamp 1624494425
transform 1 0 6867 0 1 44984
box 0 0 64 64
use contact_9  contact_9_934
timestamp 1624494425
transform 1 0 6866 0 1 44979
box 0 0 66 74
use contact_8  contact_8_283
timestamp 1624494425
transform 1 0 6442 0 1 45042
box 0 0 64 64
use contact_9  contact_9_283
timestamp 1624494425
transform 1 0 6441 0 1 45037
box 0 0 66 74
use contact_16  contact_16_427
timestamp 1624494425
transform 1 0 5224 0 1 44808
box 0 0 66 58
use contact_16  contact_16_428
timestamp 1624494425
transform 1 0 4664 0 1 44920
box 0 0 66 58
use contact_16  contact_16_423
timestamp 1624494425
transform 1 0 5784 0 1 45284
box 0 0 66 58
use contact_16  contact_16_424
timestamp 1624494425
transform 1 0 5224 0 1 45194
box 0 0 66 58
use contact_16  contact_16_425
timestamp 1624494425
transform 1 0 4744 0 1 45082
box 0 0 66 58
use and3_dec  and3_dec_140
timestamp 1624494425
transform 1 0 6203 0 -1 45820
box 0 -60 2072 490
use and3_dec  and3_dec_141
timestamp 1624494425
transform 1 0 6203 0 1 45030
box 0 -60 2072 490
use contact_8  contact_8_932
timestamp 1624494425
transform 1 0 7299 0 1 45416
box 0 0 64 64
use contact_9  contact_9_932
timestamp 1624494425
transform 1 0 7298 0 1 45411
box 0 0 66 74
use contact_8  contact_8_931
timestamp 1624494425
transform 1 0 6867 0 1 45416
box 0 0 64 64
use contact_9  contact_9_931
timestamp 1624494425
transform 1 0 6866 0 1 45411
box 0 0 66 74
use contact_8  contact_8_281
timestamp 1624494425
transform 1 0 6442 0 1 45416
box 0 0 64 64
use contact_9  contact_9_281
timestamp 1624494425
transform 1 0 6441 0 1 45411
box 0 0 66 74
use contact_16  contact_16_420
timestamp 1624494425
transform 1 0 5784 0 1 45508
box 0 0 66 58
use contact_16  contact_16_421
timestamp 1624494425
transform 1 0 5224 0 1 45598
box 0 0 66 58
use contact_8  contact_8_929
timestamp 1624494425
transform 1 0 7299 0 1 45774
box 0 0 64 64
use contact_9  contact_9_929
timestamp 1624494425
transform 1 0 7298 0 1 45769
box 0 0 66 74
use contact_8  contact_8_928
timestamp 1624494425
transform 1 0 6867 0 1 45774
box 0 0 64 64
use contact_9  contact_9_928
timestamp 1624494425
transform 1 0 6866 0 1 45769
box 0 0 66 74
use contact_8  contact_8_279
timestamp 1624494425
transform 1 0 6442 0 1 45832
box 0 0 64 64
use contact_9  contact_9_279
timestamp 1624494425
transform 1 0 6441 0 1 45827
box 0 0 66 74
use contact_16  contact_16_419
timestamp 1624494425
transform 1 0 4584 0 1 45872
box 0 0 66 58
use contact_16  contact_16_422
timestamp 1624494425
transform 1 0 4824 0 1 45710
box 0 0 66 58
use and3_dec  and3_dec_139
timestamp 1624494425
transform 1 0 6203 0 1 45820
box 0 -60 2072 490
use contact_9  contact_9_292
timestamp 1624494425
transform 1 0 7680 0 1 43018
box 0 0 66 74
use contact_8  contact_8_292
timestamp 1624494425
transform 1 0 7681 0 1 43023
box 0 0 64 64
use contact_9  contact_9_294
timestamp 1624494425
transform 1 0 7680 0 1 42623
box 0 0 66 74
use contact_8  contact_8_294
timestamp 1624494425
transform 1 0 7681 0 1 42628
box 0 0 64 64
use contact_9  contact_9_948
timestamp 1624494425
transform 1 0 8076 0 1 43018
box 0 0 66 74
use contact_8  contact_8_948
timestamp 1624494425
transform 1 0 8077 0 1 43023
box 0 0 64 64
use contact_9  contact_9_951
timestamp 1624494425
transform 1 0 8076 0 1 42623
box 0 0 66 74
use contact_8  contact_8_951
timestamp 1624494425
transform 1 0 8077 0 1 42628
box 0 0 64 64
use contact_9  contact_9_290
timestamp 1624494425
transform 1 0 7680 0 1 43413
box 0 0 66 74
use contact_8  contact_8_290
timestamp 1624494425
transform 1 0 7681 0 1 43418
box 0 0 64 64
use contact_9  contact_9_945
timestamp 1624494425
transform 1 0 8076 0 1 43413
box 0 0 66 74
use contact_8  contact_8_945
timestamp 1624494425
transform 1 0 8077 0 1 43418
box 0 0 64 64
use contact_9  contact_9_286
timestamp 1624494425
transform 1 0 7680 0 1 44203
box 0 0 66 74
use contact_8  contact_8_286
timestamp 1624494425
transform 1 0 7681 0 1 44208
box 0 0 64 64
use contact_9  contact_9_288
timestamp 1624494425
transform 1 0 7680 0 1 43808
box 0 0 66 74
use contact_8  contact_8_288
timestamp 1624494425
transform 1 0 7681 0 1 43813
box 0 0 64 64
use contact_9  contact_9_939
timestamp 1624494425
transform 1 0 8076 0 1 44203
box 0 0 66 74
use contact_8  contact_8_939
timestamp 1624494425
transform 1 0 8077 0 1 44208
box 0 0 64 64
use contact_9  contact_9_942
timestamp 1624494425
transform 1 0 8076 0 1 43808
box 0 0 66 74
use contact_8  contact_8_942
timestamp 1624494425
transform 1 0 8077 0 1 43813
box 0 0 64 64
use contact_9  contact_9_284
timestamp 1624494425
transform 1 0 7680 0 1 44598
box 0 0 66 74
use contact_8  contact_8_284
timestamp 1624494425
transform 1 0 7681 0 1 44603
box 0 0 64 64
use contact_9  contact_9_936
timestamp 1624494425
transform 1 0 8076 0 1 44598
box 0 0 66 74
use contact_8  contact_8_936
timestamp 1624494425
transform 1 0 8077 0 1 44603
box 0 0 64 64
use contact_9  contact_9_280
timestamp 1624494425
transform 1 0 7680 0 1 45388
box 0 0 66 74
use contact_8  contact_8_280
timestamp 1624494425
transform 1 0 7681 0 1 45393
box 0 0 64 64
use contact_9  contact_9_282
timestamp 1624494425
transform 1 0 7680 0 1 44993
box 0 0 66 74
use contact_8  contact_8_282
timestamp 1624494425
transform 1 0 7681 0 1 44998
box 0 0 64 64
use contact_9  contact_9_930
timestamp 1624494425
transform 1 0 8076 0 1 45388
box 0 0 66 74
use contact_8  contact_8_930
timestamp 1624494425
transform 1 0 8077 0 1 45393
box 0 0 64 64
use contact_9  contact_9_933
timestamp 1624494425
transform 1 0 8076 0 1 44993
box 0 0 66 74
use contact_8  contact_8_933
timestamp 1624494425
transform 1 0 8077 0 1 44998
box 0 0 64 64
use contact_9  contact_9_278
timestamp 1624494425
transform 1 0 7680 0 1 45783
box 0 0 66 74
use contact_8  contact_8_278
timestamp 1624494425
transform 1 0 7681 0 1 45788
box 0 0 64 64
use contact_9  contact_9_927
timestamp 1624494425
transform 1 0 8076 0 1 45783
box 0 0 66 74
use contact_8  contact_8_927
timestamp 1624494425
transform 1 0 8077 0 1 45788
box 0 0 64 64
use contact_16  contact_16_417
timestamp 1624494425
transform 1 0 5784 0 1 46074
box 0 0 66 58
use contact_16  contact_16_418
timestamp 1624494425
transform 1 0 5304 0 1 45984
box 0 0 66 58
use contact_8  contact_8_926
timestamp 1624494425
transform 1 0 7299 0 1 46206
box 0 0 64 64
use contact_9  contact_9_926
timestamp 1624494425
transform 1 0 7298 0 1 46201
box 0 0 66 74
use contact_8  contact_8_925
timestamp 1624494425
transform 1 0 6867 0 1 46206
box 0 0 64 64
use contact_9  contact_9_925
timestamp 1624494425
transform 1 0 6866 0 1 46201
box 0 0 66 74
use contact_8  contact_8_277
timestamp 1624494425
transform 1 0 6442 0 1 46206
box 0 0 64 64
use contact_9  contact_9_277
timestamp 1624494425
transform 1 0 6441 0 1 46201
box 0 0 66 74
use contact_16  contact_16_414
timestamp 1624494425
transform 1 0 5784 0 1 46298
box 0 0 66 58
use contact_16  contact_16_415
timestamp 1624494425
transform 1 0 5304 0 1 46388
box 0 0 66 58
use and3_dec  and3_dec_138
timestamp 1624494425
transform 1 0 6203 0 -1 46610
box 0 -60 2072 490
use contact_8  contact_8_923
timestamp 1624494425
transform 1 0 7299 0 1 46564
box 0 0 64 64
use contact_9  contact_9_923
timestamp 1624494425
transform 1 0 7298 0 1 46559
box 0 0 66 74
use contact_8  contact_8_922
timestamp 1624494425
transform 1 0 6867 0 1 46564
box 0 0 64 64
use contact_9  contact_9_922
timestamp 1624494425
transform 1 0 6866 0 1 46559
box 0 0 66 74
use contact_8  contact_8_275
timestamp 1624494425
transform 1 0 6442 0 1 46622
box 0 0 64 64
use contact_9  contact_9_275
timestamp 1624494425
transform 1 0 6441 0 1 46617
box 0 0 66 74
use contact_16  contact_16_413
timestamp 1624494425
transform 1 0 4744 0 1 46662
box 0 0 66 58
use contact_16  contact_16_416
timestamp 1624494425
transform 1 0 4664 0 1 46500
box 0 0 66 58
use contact_16  contact_16_411
timestamp 1624494425
transform 1 0 5784 0 1 46864
box 0 0 66 58
use contact_16  contact_16_412
timestamp 1624494425
transform 1 0 5304 0 1 46774
box 0 0 66 58
use and3_dec  and3_dec_136
timestamp 1624494425
transform 1 0 6203 0 -1 47400
box 0 -60 2072 490
use and3_dec  and3_dec_137
timestamp 1624494425
transform 1 0 6203 0 1 46610
box 0 -60 2072 490
use contact_8  contact_8_920
timestamp 1624494425
transform 1 0 7299 0 1 46996
box 0 0 64 64
use contact_9  contact_9_920
timestamp 1624494425
transform 1 0 7298 0 1 46991
box 0 0 66 74
use contact_8  contact_8_919
timestamp 1624494425
transform 1 0 6867 0 1 46996
box 0 0 64 64
use contact_9  contact_9_919
timestamp 1624494425
transform 1 0 6866 0 1 46991
box 0 0 66 74
use contact_8  contact_8_273
timestamp 1624494425
transform 1 0 6442 0 1 46996
box 0 0 64 64
use contact_9  contact_9_273
timestamp 1624494425
transform 1 0 6441 0 1 46991
box 0 0 66 74
use contact_16  contact_16_408
timestamp 1624494425
transform 1 0 5784 0 1 47088
box 0 0 66 58
use contact_16  contact_16_409
timestamp 1624494425
transform 1 0 5304 0 1 47178
box 0 0 66 58
use contact_8  contact_8_917
timestamp 1624494425
transform 1 0 7299 0 1 47354
box 0 0 64 64
use contact_9  contact_9_917
timestamp 1624494425
transform 1 0 7298 0 1 47349
box 0 0 66 74
use contact_8  contact_8_916
timestamp 1624494425
transform 1 0 6867 0 1 47354
box 0 0 64 64
use contact_9  contact_9_916
timestamp 1624494425
transform 1 0 6866 0 1 47349
box 0 0 66 74
use contact_8  contact_8_271
timestamp 1624494425
transform 1 0 6442 0 1 47412
box 0 0 64 64
use contact_9  contact_9_271
timestamp 1624494425
transform 1 0 6441 0 1 47407
box 0 0 66 74
use contact_16  contact_16_407
timestamp 1624494425
transform 1 0 4584 0 1 47452
box 0 0 66 58
use contact_16  contact_16_410
timestamp 1624494425
transform 1 0 4824 0 1 47290
box 0 0 66 58
use and3_dec  and3_dec_135
timestamp 1624494425
transform 1 0 6203 0 1 47400
box 0 -60 2072 490
use contact_8  contact_8_914
timestamp 1624494425
transform 1 0 7299 0 1 47786
box 0 0 64 64
use contact_9  contact_9_914
timestamp 1624494425
transform 1 0 7298 0 1 47781
box 0 0 66 74
use contact_8  contact_8_913
timestamp 1624494425
transform 1 0 6867 0 1 47786
box 0 0 64 64
use contact_9  contact_9_913
timestamp 1624494425
transform 1 0 6866 0 1 47781
box 0 0 66 74
use contact_8  contact_8_269
timestamp 1624494425
transform 1 0 6442 0 1 47786
box 0 0 64 64
use contact_9  contact_9_269
timestamp 1624494425
transform 1 0 6441 0 1 47781
box 0 0 66 74
use contact_16  contact_16_405
timestamp 1624494425
transform 1 0 5784 0 1 47654
box 0 0 66 58
use contact_16  contact_16_406
timestamp 1624494425
transform 1 0 5384 0 1 47564
box 0 0 66 58
use contact_16  contact_16_402
timestamp 1624494425
transform 1 0 5784 0 1 47878
box 0 0 66 58
use contact_16  contact_16_403
timestamp 1624494425
transform 1 0 5384 0 1 47968
box 0 0 66 58
use and3_dec  and3_dec_134
timestamp 1624494425
transform 1 0 6203 0 -1 48190
box 0 -60 2072 490
use contact_8  contact_8_911
timestamp 1624494425
transform 1 0 7299 0 1 48144
box 0 0 64 64
use contact_9  contact_9_911
timestamp 1624494425
transform 1 0 7298 0 1 48139
box 0 0 66 74
use contact_8  contact_8_910
timestamp 1624494425
transform 1 0 6867 0 1 48144
box 0 0 64 64
use contact_9  contact_9_910
timestamp 1624494425
transform 1 0 6866 0 1 48139
box 0 0 66 74
use contact_8  contact_8_267
timestamp 1624494425
transform 1 0 6442 0 1 48202
box 0 0 64 64
use contact_9  contact_9_267
timestamp 1624494425
transform 1 0 6441 0 1 48197
box 0 0 66 74
use contact_16  contact_16_401
timestamp 1624494425
transform 1 0 4744 0 1 48242
box 0 0 66 58
use contact_16  contact_16_404
timestamp 1624494425
transform 1 0 4664 0 1 48080
box 0 0 66 58
use contact_8  contact_8_908
timestamp 1624494425
transform 1 0 7299 0 1 48576
box 0 0 64 64
use contact_9  contact_9_908
timestamp 1624494425
transform 1 0 7298 0 1 48571
box 0 0 66 74
use contact_8  contact_8_907
timestamp 1624494425
transform 1 0 6867 0 1 48576
box 0 0 64 64
use contact_9  contact_9_907
timestamp 1624494425
transform 1 0 6866 0 1 48571
box 0 0 66 74
use contact_8  contact_8_265
timestamp 1624494425
transform 1 0 6442 0 1 48576
box 0 0 64 64
use contact_9  contact_9_265
timestamp 1624494425
transform 1 0 6441 0 1 48571
box 0 0 66 74
use contact_16  contact_16_399
timestamp 1624494425
transform 1 0 5784 0 1 48444
box 0 0 66 58
use contact_16  contact_16_400
timestamp 1624494425
transform 1 0 5384 0 1 48354
box 0 0 66 58
use and3_dec  and3_dec_132
timestamp 1624494425
transform 1 0 6203 0 -1 48980
box 0 -60 2072 490
use and3_dec  and3_dec_133
timestamp 1624494425
transform 1 0 6203 0 1 48190
box 0 -60 2072 490
use contact_16  contact_16_396
timestamp 1624494425
transform 1 0 5784 0 1 48668
box 0 0 66 58
use contact_16  contact_16_397
timestamp 1624494425
transform 1 0 5384 0 1 48758
box 0 0 66 58
use contact_16  contact_16_398
timestamp 1624494425
transform 1 0 4824 0 1 48870
box 0 0 66 58
use contact_8  contact_8_905
timestamp 1624494425
transform 1 0 7299 0 1 48934
box 0 0 64 64
use contact_9  contact_9_905
timestamp 1624494425
transform 1 0 7298 0 1 48929
box 0 0 66 74
use contact_8  contact_8_904
timestamp 1624494425
transform 1 0 6867 0 1 48934
box 0 0 64 64
use contact_9  contact_9_904
timestamp 1624494425
transform 1 0 6866 0 1 48929
box 0 0 66 74
use contact_8  contact_8_263
timestamp 1624494425
transform 1 0 6442 0 1 48992
box 0 0 64 64
use contact_9  contact_9_263
timestamp 1624494425
transform 1 0 6441 0 1 48987
box 0 0 66 74
use contact_16  contact_16_394
timestamp 1624494425
transform 1 0 5464 0 1 49144
box 0 0 66 58
use contact_16  contact_16_395
timestamp 1624494425
transform 1 0 4584 0 1 49032
box 0 0 66 58
use and3_dec  and3_dec_131
timestamp 1624494425
transform 1 0 6203 0 1 48980
box 0 -60 2072 490
use contact_9  contact_9_276
timestamp 1624494425
transform 1 0 7680 0 1 46178
box 0 0 66 74
use contact_8  contact_8_276
timestamp 1624494425
transform 1 0 7681 0 1 46183
box 0 0 64 64
use contact_9  contact_9_924
timestamp 1624494425
transform 1 0 8076 0 1 46178
box 0 0 66 74
use contact_8  contact_8_924
timestamp 1624494425
transform 1 0 8077 0 1 46183
box 0 0 64 64
use contact_9  contact_9_272
timestamp 1624494425
transform 1 0 7680 0 1 46968
box 0 0 66 74
use contact_8  contact_8_272
timestamp 1624494425
transform 1 0 7681 0 1 46973
box 0 0 64 64
use contact_9  contact_9_274
timestamp 1624494425
transform 1 0 7680 0 1 46573
box 0 0 66 74
use contact_8  contact_8_274
timestamp 1624494425
transform 1 0 7681 0 1 46578
box 0 0 64 64
use contact_9  contact_9_918
timestamp 1624494425
transform 1 0 8076 0 1 46968
box 0 0 66 74
use contact_8  contact_8_918
timestamp 1624494425
transform 1 0 8077 0 1 46973
box 0 0 64 64
use contact_9  contact_9_921
timestamp 1624494425
transform 1 0 8076 0 1 46573
box 0 0 66 74
use contact_8  contact_8_921
timestamp 1624494425
transform 1 0 8077 0 1 46578
box 0 0 64 64
use contact_9  contact_9_270
timestamp 1624494425
transform 1 0 7680 0 1 47363
box 0 0 66 74
use contact_8  contact_8_270
timestamp 1624494425
transform 1 0 7681 0 1 47368
box 0 0 64 64
use contact_9  contact_9_915
timestamp 1624494425
transform 1 0 8076 0 1 47363
box 0 0 66 74
use contact_8  contact_8_915
timestamp 1624494425
transform 1 0 8077 0 1 47368
box 0 0 64 64
use contact_9  contact_9_266
timestamp 1624494425
transform 1 0 7680 0 1 48153
box 0 0 66 74
use contact_8  contact_8_266
timestamp 1624494425
transform 1 0 7681 0 1 48158
box 0 0 64 64
use contact_9  contact_9_268
timestamp 1624494425
transform 1 0 7680 0 1 47758
box 0 0 66 74
use contact_8  contact_8_268
timestamp 1624494425
transform 1 0 7681 0 1 47763
box 0 0 64 64
use contact_9  contact_9_909
timestamp 1624494425
transform 1 0 8076 0 1 48153
box 0 0 66 74
use contact_8  contact_8_909
timestamp 1624494425
transform 1 0 8077 0 1 48158
box 0 0 64 64
use contact_9  contact_9_912
timestamp 1624494425
transform 1 0 8076 0 1 47758
box 0 0 66 74
use contact_8  contact_8_912
timestamp 1624494425
transform 1 0 8077 0 1 47763
box 0 0 64 64
use contact_9  contact_9_262
timestamp 1624494425
transform 1 0 7680 0 1 48943
box 0 0 66 74
use contact_8  contact_8_262
timestamp 1624494425
transform 1 0 7681 0 1 48948
box 0 0 64 64
use contact_9  contact_9_264
timestamp 1624494425
transform 1 0 7680 0 1 48548
box 0 0 66 74
use contact_8  contact_8_264
timestamp 1624494425
transform 1 0 7681 0 1 48553
box 0 0 64 64
use contact_9  contact_9_903
timestamp 1624494425
transform 1 0 8076 0 1 48943
box 0 0 66 74
use contact_8  contact_8_903
timestamp 1624494425
transform 1 0 8077 0 1 48948
box 0 0 64 64
use contact_9  contact_9_906
timestamp 1624494425
transform 1 0 8076 0 1 48548
box 0 0 66 74
use contact_8  contact_8_906
timestamp 1624494425
transform 1 0 8077 0 1 48553
box 0 0 64 64
use contact_8  contact_8_902
timestamp 1624494425
transform 1 0 7299 0 1 49366
box 0 0 64 64
use contact_9  contact_9_902
timestamp 1624494425
transform 1 0 7298 0 1 49361
box 0 0 66 74
use contact_8  contact_8_901
timestamp 1624494425
transform 1 0 6867 0 1 49366
box 0 0 64 64
use contact_9  contact_9_901
timestamp 1624494425
transform 1 0 6866 0 1 49361
box 0 0 66 74
use contact_8  contact_8_261
timestamp 1624494425
transform 1 0 6442 0 1 49366
box 0 0 64 64
use contact_9  contact_9_261
timestamp 1624494425
transform 1 0 6441 0 1 49361
box 0 0 66 74
use contact_16  contact_16_393
timestamp 1624494425
transform 1 0 5784 0 1 49234
box 0 0 66 58
use contact_16  contact_16_390
timestamp 1624494425
transform 1 0 5784 0 1 49458
box 0 0 66 58
use contact_16  contact_16_391
timestamp 1624494425
transform 1 0 5464 0 1 49548
box 0 0 66 58
use contact_16  contact_16_392
timestamp 1624494425
transform 1 0 4664 0 1 49660
box 0 0 66 58
use and3_dec  and3_dec_130
timestamp 1624494425
transform 1 0 6203 0 -1 49770
box 0 -60 2072 490
use contact_8  contact_8_899
timestamp 1624494425
transform 1 0 7299 0 1 49724
box 0 0 64 64
use contact_9  contact_9_899
timestamp 1624494425
transform 1 0 7298 0 1 49719
box 0 0 66 74
use contact_8  contact_8_898
timestamp 1624494425
transform 1 0 6867 0 1 49724
box 0 0 64 64
use contact_9  contact_9_898
timestamp 1624494425
transform 1 0 6866 0 1 49719
box 0 0 66 74
use contact_8  contact_8_259
timestamp 1624494425
transform 1 0 6442 0 1 49782
box 0 0 64 64
use contact_9  contact_9_259
timestamp 1624494425
transform 1 0 6441 0 1 49777
box 0 0 66 74
use contact_16  contact_16_388
timestamp 1624494425
transform 1 0 5464 0 1 49934
box 0 0 66 58
use contact_16  contact_16_389
timestamp 1624494425
transform 1 0 4744 0 1 49822
box 0 0 66 58
use contact_8  contact_8_896
timestamp 1624494425
transform 1 0 7299 0 1 50156
box 0 0 64 64
use contact_9  contact_9_896
timestamp 1624494425
transform 1 0 7298 0 1 50151
box 0 0 66 74
use contact_8  contact_8_895
timestamp 1624494425
transform 1 0 6867 0 1 50156
box 0 0 64 64
use contact_9  contact_9_895
timestamp 1624494425
transform 1 0 6866 0 1 50151
box 0 0 66 74
use contact_8  contact_8_257
timestamp 1624494425
transform 1 0 6442 0 1 50156
box 0 0 64 64
use contact_9  contact_9_257
timestamp 1624494425
transform 1 0 6441 0 1 50151
box 0 0 66 74
use contact_16  contact_16_384
timestamp 1624494425
transform 1 0 5784 0 1 50248
box 0 0 66 58
use contact_16  contact_16_387
timestamp 1624494425
transform 1 0 5784 0 1 50024
box 0 0 66 58
use and3_dec  and3_dec_128
timestamp 1624494425
transform 1 0 6203 0 -1 50560
box 0 -60 2072 490
use and3_dec  and3_dec_129
timestamp 1624494425
transform 1 0 6203 0 1 49770
box 0 -60 2072 490
use contact_8  contact_8_893
timestamp 1624494425
transform 1 0 7299 0 1 50514
box 0 0 64 64
use contact_9  contact_9_893
timestamp 1624494425
transform 1 0 7298 0 1 50509
box 0 0 66 74
use contact_8  contact_8_892
timestamp 1624494425
transform 1 0 6867 0 1 50514
box 0 0 64 64
use contact_9  contact_9_892
timestamp 1624494425
transform 1 0 6866 0 1 50509
box 0 0 66 74
use contact_16  contact_16_385
timestamp 1624494425
transform 1 0 5464 0 1 50338
box 0 0 66 58
use contact_16  contact_16_386
timestamp 1624494425
transform 1 0 4824 0 1 50450
box 0 0 66 58
use contact_8  contact_8_255
timestamp 1624494425
transform 1 0 6442 0 1 50572
box 0 0 64 64
use contact_9  contact_9_255
timestamp 1624494425
transform 1 0 6441 0 1 50567
box 0 0 66 74
use contact_16  contact_16_382
timestamp 1624494425
transform 1 0 4904 0 1 50724
box 0 0 66 58
use contact_16  contact_16_383
timestamp 1624494425
transform 1 0 4584 0 1 50612
box 0 0 66 58
use and3_dec  and3_dec_127
timestamp 1624494425
transform 1 0 6203 0 1 50560
box 0 -60 2072 490
use contact_8  contact_8_890
timestamp 1624494425
transform 1 0 7299 0 1 50946
box 0 0 64 64
use contact_9  contact_9_890
timestamp 1624494425
transform 1 0 7298 0 1 50941
box 0 0 66 74
use contact_8  contact_8_889
timestamp 1624494425
transform 1 0 6867 0 1 50946
box 0 0 64 64
use contact_9  contact_9_889
timestamp 1624494425
transform 1 0 6866 0 1 50941
box 0 0 66 74
use contact_8  contact_8_253
timestamp 1624494425
transform 1 0 6442 0 1 50946
box 0 0 64 64
use contact_9  contact_9_253
timestamp 1624494425
transform 1 0 6441 0 1 50941
box 0 0 66 74
use contact_16  contact_16_378
timestamp 1624494425
transform 1 0 5864 0 1 51038
box 0 0 66 58
use contact_16  contact_16_381
timestamp 1624494425
transform 1 0 5864 0 1 50814
box 0 0 66 58
use contact_8  contact_8_887
timestamp 1624494425
transform 1 0 7299 0 1 51304
box 0 0 64 64
use contact_9  contact_9_887
timestamp 1624494425
transform 1 0 7298 0 1 51299
box 0 0 66 74
use contact_8  contact_8_886
timestamp 1624494425
transform 1 0 6867 0 1 51304
box 0 0 64 64
use contact_9  contact_9_886
timestamp 1624494425
transform 1 0 6866 0 1 51299
box 0 0 66 74
use contact_9  contact_9_251
timestamp 1624494425
transform 1 0 6441 0 1 51357
box 0 0 66 74
use contact_16  contact_16_379
timestamp 1624494425
transform 1 0 4904 0 1 51128
box 0 0 66 58
use contact_16  contact_16_380
timestamp 1624494425
transform 1 0 4664 0 1 51240
box 0 0 66 58
use and3_dec  and3_dec_125
timestamp 1624494425
transform 1 0 6203 0 1 51350
box 0 -60 2072 490
use and3_dec  and3_dec_126
timestamp 1624494425
transform 1 0 6203 0 -1 51350
box 0 -60 2072 490
use contact_8  contact_8_251
timestamp 1624494425
transform 1 0 6442 0 1 51362
box 0 0 64 64
use contact_16  contact_16_375
timestamp 1624494425
transform 1 0 5864 0 1 51604
box 0 0 66 58
use contact_16  contact_16_376
timestamp 1624494425
transform 1 0 4904 0 1 51514
box 0 0 66 58
use contact_16  contact_16_377
timestamp 1624494425
transform 1 0 4744 0 1 51402
box 0 0 66 58
use contact_8  contact_8_884
timestamp 1624494425
transform 1 0 7299 0 1 51736
box 0 0 64 64
use contact_9  contact_9_884
timestamp 1624494425
transform 1 0 7298 0 1 51731
box 0 0 66 74
use contact_8  contact_8_883
timestamp 1624494425
transform 1 0 6867 0 1 51736
box 0 0 64 64
use contact_9  contact_9_883
timestamp 1624494425
transform 1 0 6866 0 1 51731
box 0 0 66 74
use contact_8  contact_8_249
timestamp 1624494425
transform 1 0 6442 0 1 51736
box 0 0 64 64
use contact_9  contact_9_249
timestamp 1624494425
transform 1 0 6441 0 1 51731
box 0 0 66 74
use contact_16  contact_16_372
timestamp 1624494425
transform 1 0 5864 0 1 51828
box 0 0 66 58
use and3_dec  and3_dec_124
timestamp 1624494425
transform 1 0 6203 0 -1 52140
box 0 -60 2072 490
use contact_8  contact_8_881
timestamp 1624494425
transform 1 0 7299 0 1 52094
box 0 0 64 64
use contact_9  contact_9_881
timestamp 1624494425
transform 1 0 7298 0 1 52089
box 0 0 66 74
use contact_8  contact_8_880
timestamp 1624494425
transform 1 0 6867 0 1 52094
box 0 0 64 64
use contact_9  contact_9_880
timestamp 1624494425
transform 1 0 6866 0 1 52089
box 0 0 66 74
use contact_8  contact_8_247
timestamp 1624494425
transform 1 0 6442 0 1 52152
box 0 0 64 64
use contact_9  contact_9_247
timestamp 1624494425
transform 1 0 6441 0 1 52147
box 0 0 66 74
use contact_16  contact_16_373
timestamp 1624494425
transform 1 0 4904 0 1 51918
box 0 0 66 58
use contact_16  contact_16_374
timestamp 1624494425
transform 1 0 4824 0 1 52030
box 0 0 66 58
use contact_16  contact_16_369
timestamp 1624494425
transform 1 0 5864 0 1 52394
box 0 0 66 58
use contact_16  contact_16_370
timestamp 1624494425
transform 1 0 4984 0 1 52304
box 0 0 66 58
use contact_16  contact_16_371
timestamp 1624494425
transform 1 0 4584 0 1 52192
box 0 0 66 58
use and3_dec  and3_dec_123
timestamp 1624494425
transform 1 0 6203 0 1 52140
box 0 -60 2072 490
use contact_9  contact_9_258
timestamp 1624494425
transform 1 0 7680 0 1 49733
box 0 0 66 74
use contact_8  contact_8_258
timestamp 1624494425
transform 1 0 7681 0 1 49738
box 0 0 64 64
use contact_9  contact_9_260
timestamp 1624494425
transform 1 0 7680 0 1 49338
box 0 0 66 74
use contact_8  contact_8_260
timestamp 1624494425
transform 1 0 7681 0 1 49343
box 0 0 64 64
use contact_9  contact_9_897
timestamp 1624494425
transform 1 0 8076 0 1 49733
box 0 0 66 74
use contact_8  contact_8_897
timestamp 1624494425
transform 1 0 8077 0 1 49738
box 0 0 64 64
use contact_9  contact_9_900
timestamp 1624494425
transform 1 0 8076 0 1 49338
box 0 0 66 74
use contact_8  contact_8_900
timestamp 1624494425
transform 1 0 8077 0 1 49343
box 0 0 64 64
use contact_9  contact_9_256
timestamp 1624494425
transform 1 0 7680 0 1 50128
box 0 0 66 74
use contact_8  contact_8_256
timestamp 1624494425
transform 1 0 7681 0 1 50133
box 0 0 64 64
use contact_9  contact_9_894
timestamp 1624494425
transform 1 0 8076 0 1 50128
box 0 0 66 74
use contact_8  contact_8_894
timestamp 1624494425
transform 1 0 8077 0 1 50133
box 0 0 64 64
use contact_9  contact_9_252
timestamp 1624494425
transform 1 0 7680 0 1 50918
box 0 0 66 74
use contact_8  contact_8_252
timestamp 1624494425
transform 1 0 7681 0 1 50923
box 0 0 64 64
use contact_9  contact_9_254
timestamp 1624494425
transform 1 0 7680 0 1 50523
box 0 0 66 74
use contact_8  contact_8_254
timestamp 1624494425
transform 1 0 7681 0 1 50528
box 0 0 64 64
use contact_9  contact_9_888
timestamp 1624494425
transform 1 0 8076 0 1 50918
box 0 0 66 74
use contact_8  contact_8_888
timestamp 1624494425
transform 1 0 8077 0 1 50923
box 0 0 64 64
use contact_9  contact_9_891
timestamp 1624494425
transform 1 0 8076 0 1 50523
box 0 0 66 74
use contact_8  contact_8_891
timestamp 1624494425
transform 1 0 8077 0 1 50528
box 0 0 64 64
use contact_9  contact_9_250
timestamp 1624494425
transform 1 0 7680 0 1 51313
box 0 0 66 74
use contact_8  contact_8_250
timestamp 1624494425
transform 1 0 7681 0 1 51318
box 0 0 64 64
use contact_9  contact_9_885
timestamp 1624494425
transform 1 0 8076 0 1 51313
box 0 0 66 74
use contact_8  contact_8_885
timestamp 1624494425
transform 1 0 8077 0 1 51318
box 0 0 64 64
use contact_9  contact_9_246
timestamp 1624494425
transform 1 0 7680 0 1 52103
box 0 0 66 74
use contact_8  contact_8_246
timestamp 1624494425
transform 1 0 7681 0 1 52108
box 0 0 64 64
use contact_9  contact_9_248
timestamp 1624494425
transform 1 0 7680 0 1 51708
box 0 0 66 74
use contact_8  contact_8_248
timestamp 1624494425
transform 1 0 7681 0 1 51713
box 0 0 64 64
use contact_9  contact_9_879
timestamp 1624494425
transform 1 0 8076 0 1 52103
box 0 0 66 74
use contact_8  contact_8_879
timestamp 1624494425
transform 1 0 8077 0 1 52108
box 0 0 64 64
use contact_9  contact_9_882
timestamp 1624494425
transform 1 0 8076 0 1 51708
box 0 0 66 74
use contact_8  contact_8_882
timestamp 1624494425
transform 1 0 8077 0 1 51713
box 0 0 64 64
use contact_8  contact_8_878
timestamp 1624494425
transform 1 0 7299 0 1 52526
box 0 0 64 64
use contact_9  contact_9_878
timestamp 1624494425
transform 1 0 7298 0 1 52521
box 0 0 66 74
use contact_8  contact_8_877
timestamp 1624494425
transform 1 0 6867 0 1 52526
box 0 0 64 64
use contact_9  contact_9_877
timestamp 1624494425
transform 1 0 6866 0 1 52521
box 0 0 66 74
use contact_8  contact_8_245
timestamp 1624494425
transform 1 0 6442 0 1 52526
box 0 0 64 64
use contact_9  contact_9_245
timestamp 1624494425
transform 1 0 6441 0 1 52521
box 0 0 66 74
use contact_16  contact_16_366
timestamp 1624494425
transform 1 0 5864 0 1 52618
box 0 0 66 58
use contact_16  contact_16_367
timestamp 1624494425
transform 1 0 4984 0 1 52708
box 0 0 66 58
use contact_8  contact_8_875
timestamp 1624494425
transform 1 0 7299 0 1 52884
box 0 0 64 64
use contact_9  contact_9_875
timestamp 1624494425
transform 1 0 7298 0 1 52879
box 0 0 66 74
use contact_8  contact_8_874
timestamp 1624494425
transform 1 0 6867 0 1 52884
box 0 0 64 64
use contact_9  contact_9_874
timestamp 1624494425
transform 1 0 6866 0 1 52879
box 0 0 66 74
use contact_8  contact_8_243
timestamp 1624494425
transform 1 0 6442 0 1 52942
box 0 0 64 64
use contact_9  contact_9_243
timestamp 1624494425
transform 1 0 6441 0 1 52937
box 0 0 66 74
use contact_16  contact_16_365
timestamp 1624494425
transform 1 0 4744 0 1 52982
box 0 0 66 58
use contact_16  contact_16_368
timestamp 1624494425
transform 1 0 4664 0 1 52820
box 0 0 66 58
use and3_dec  and3_dec_121
timestamp 1624494425
transform 1 0 6203 0 1 52930
box 0 -60 2072 490
use and3_dec  and3_dec_122
timestamp 1624494425
transform 1 0 6203 0 -1 52930
box 0 -60 2072 490
use contact_16  contact_16_363
timestamp 1624494425
transform 1 0 5864 0 1 53184
box 0 0 66 58
use contact_16  contact_16_364
timestamp 1624494425
transform 1 0 4984 0 1 53094
box 0 0 66 58
use contact_8  contact_8_872
timestamp 1624494425
transform 1 0 7299 0 1 53316
box 0 0 64 64
use contact_9  contact_9_872
timestamp 1624494425
transform 1 0 7298 0 1 53311
box 0 0 66 74
use contact_8  contact_8_871
timestamp 1624494425
transform 1 0 6867 0 1 53316
box 0 0 64 64
use contact_9  contact_9_871
timestamp 1624494425
transform 1 0 6866 0 1 53311
box 0 0 66 74
use contact_8  contact_8_241
timestamp 1624494425
transform 1 0 6442 0 1 53316
box 0 0 64 64
use contact_9  contact_9_241
timestamp 1624494425
transform 1 0 6441 0 1 53311
box 0 0 66 74
use contact_16  contact_16_360
timestamp 1624494425
transform 1 0 5864 0 1 53408
box 0 0 66 58
use contact_16  contact_16_361
timestamp 1624494425
transform 1 0 4984 0 1 53498
box 0 0 66 58
use and3_dec  and3_dec_120
timestamp 1624494425
transform 1 0 6203 0 -1 53720
box 0 -60 2072 490
use contact_8  contact_8_869
timestamp 1624494425
transform 1 0 7299 0 1 53674
box 0 0 64 64
use contact_9  contact_9_869
timestamp 1624494425
transform 1 0 7298 0 1 53669
box 0 0 66 74
use contact_8  contact_8_868
timestamp 1624494425
transform 1 0 6867 0 1 53674
box 0 0 64 64
use contact_9  contact_9_868
timestamp 1624494425
transform 1 0 6866 0 1 53669
box 0 0 66 74
use contact_8  contact_8_239
timestamp 1624494425
transform 1 0 6442 0 1 53732
box 0 0 64 64
use contact_9  contact_9_239
timestamp 1624494425
transform 1 0 6441 0 1 53727
box 0 0 66 74
use contact_16  contact_16_359
timestamp 1624494425
transform 1 0 4584 0 1 53772
box 0 0 66 58
use contact_16  contact_16_362
timestamp 1624494425
transform 1 0 4824 0 1 53610
box 0 0 66 58
use contact_16  contact_16_357
timestamp 1624494425
transform 1 0 5864 0 1 53974
box 0 0 66 58
use contact_16  contact_16_358
timestamp 1624494425
transform 1 0 5064 0 1 53884
box 0 0 66 58
use and3_dec  and3_dec_118
timestamp 1624494425
transform 1 0 6203 0 -1 54510
box 0 -60 2072 490
use and3_dec  and3_dec_119
timestamp 1624494425
transform 1 0 6203 0 1 53720
box 0 -60 2072 490
use contact_8  contact_8_866
timestamp 1624494425
transform 1 0 7299 0 1 54106
box 0 0 64 64
use contact_9  contact_9_866
timestamp 1624494425
transform 1 0 7298 0 1 54101
box 0 0 66 74
use contact_8  contact_8_865
timestamp 1624494425
transform 1 0 6867 0 1 54106
box 0 0 64 64
use contact_9  contact_9_865
timestamp 1624494425
transform 1 0 6866 0 1 54101
box 0 0 66 74
use contact_8  contact_8_237
timestamp 1624494425
transform 1 0 6442 0 1 54106
box 0 0 64 64
use contact_9  contact_9_237
timestamp 1624494425
transform 1 0 6441 0 1 54101
box 0 0 66 74
use contact_16  contact_16_354
timestamp 1624494425
transform 1 0 5864 0 1 54198
box 0 0 66 58
use contact_16  contact_16_355
timestamp 1624494425
transform 1 0 5064 0 1 54288
box 0 0 66 58
use contact_8  contact_8_863
timestamp 1624494425
transform 1 0 7299 0 1 54464
box 0 0 64 64
use contact_9  contact_9_863
timestamp 1624494425
transform 1 0 7298 0 1 54459
box 0 0 66 74
use contact_8  contact_8_862
timestamp 1624494425
transform 1 0 6867 0 1 54464
box 0 0 64 64
use contact_9  contact_9_862
timestamp 1624494425
transform 1 0 6866 0 1 54459
box 0 0 66 74
use contact_8  contact_8_235
timestamp 1624494425
transform 1 0 6442 0 1 54522
box 0 0 64 64
use contact_9  contact_9_235
timestamp 1624494425
transform 1 0 6441 0 1 54517
box 0 0 66 74
use contact_16  contact_16_353
timestamp 1624494425
transform 1 0 4744 0 1 54562
box 0 0 66 58
use contact_16  contact_16_356
timestamp 1624494425
transform 1 0 4664 0 1 54400
box 0 0 66 58
use and3_dec  and3_dec_117
timestamp 1624494425
transform 1 0 6203 0 1 54510
box 0 -60 2072 490
use contact_8  contact_8_860
timestamp 1624494425
transform 1 0 7299 0 1 54896
box 0 0 64 64
use contact_9  contact_9_860
timestamp 1624494425
transform 1 0 7298 0 1 54891
box 0 0 66 74
use contact_8  contact_8_859
timestamp 1624494425
transform 1 0 6867 0 1 54896
box 0 0 64 64
use contact_9  contact_9_859
timestamp 1624494425
transform 1 0 6866 0 1 54891
box 0 0 66 74
use contact_8  contact_8_233
timestamp 1624494425
transform 1 0 6442 0 1 54896
box 0 0 64 64
use contact_9  contact_9_233
timestamp 1624494425
transform 1 0 6441 0 1 54891
box 0 0 66 74
use contact_16  contact_16_351
timestamp 1624494425
transform 1 0 5864 0 1 54764
box 0 0 66 58
use contact_16  contact_16_352
timestamp 1624494425
transform 1 0 5064 0 1 54674
box 0 0 66 58
use contact_16  contact_16_348
timestamp 1624494425
transform 1 0 5864 0 1 54988
box 0 0 66 58
use contact_16  contact_16_349
timestamp 1624494425
transform 1 0 5064 0 1 55078
box 0 0 66 58
use contact_16  contact_16_350
timestamp 1624494425
transform 1 0 4824 0 1 55190
box 0 0 66 58
use and3_dec  and3_dec_116
timestamp 1624494425
transform 1 0 6203 0 -1 55300
box 0 -60 2072 490
use contact_8  contact_8_857
timestamp 1624494425
transform 1 0 7299 0 1 55254
box 0 0 64 64
use contact_9  contact_9_857
timestamp 1624494425
transform 1 0 7298 0 1 55249
box 0 0 66 74
use contact_8  contact_8_856
timestamp 1624494425
transform 1 0 6867 0 1 55254
box 0 0 64 64
use contact_9  contact_9_856
timestamp 1624494425
transform 1 0 6866 0 1 55249
box 0 0 66 74
use contact_8  contact_8_231
timestamp 1624494425
transform 1 0 6442 0 1 55312
box 0 0 64 64
use contact_9  contact_9_231
timestamp 1624494425
transform 1 0 6441 0 1 55307
box 0 0 66 74
use contact_16  contact_16_346
timestamp 1624494425
transform 1 0 5144 0 1 55464
box 0 0 66 58
use contact_16  contact_16_347
timestamp 1624494425
transform 1 0 4584 0 1 55352
box 0 0 66 58
use contact_8  contact_8_854
timestamp 1624494425
transform 1 0 7299 0 1 55686
box 0 0 64 64
use contact_9  contact_9_854
timestamp 1624494425
transform 1 0 7298 0 1 55681
box 0 0 66 74
use contact_8  contact_8_853
timestamp 1624494425
transform 1 0 6867 0 1 55686
box 0 0 64 64
use contact_9  contact_9_853
timestamp 1624494425
transform 1 0 6866 0 1 55681
box 0 0 66 74
use contact_8  contact_8_229
timestamp 1624494425
transform 1 0 6442 0 1 55686
box 0 0 64 64
use contact_9  contact_9_229
timestamp 1624494425
transform 1 0 6441 0 1 55681
box 0 0 66 74
use contact_16  contact_16_345
timestamp 1624494425
transform 1 0 5864 0 1 55554
box 0 0 66 58
use and3_dec  and3_dec_114
timestamp 1624494425
transform 1 0 6203 0 -1 56090
box 0 -60 2072 490
use and3_dec  and3_dec_115
timestamp 1624494425
transform 1 0 6203 0 1 55300
box 0 -60 2072 490
use contact_9  contact_9_242
timestamp 1624494425
transform 1 0 7680 0 1 52893
box 0 0 66 74
use contact_8  contact_8_242
timestamp 1624494425
transform 1 0 7681 0 1 52898
box 0 0 64 64
use contact_9  contact_9_244
timestamp 1624494425
transform 1 0 7680 0 1 52498
box 0 0 66 74
use contact_8  contact_8_244
timestamp 1624494425
transform 1 0 7681 0 1 52503
box 0 0 64 64
use contact_9  contact_9_873
timestamp 1624494425
transform 1 0 8076 0 1 52893
box 0 0 66 74
use contact_8  contact_8_873
timestamp 1624494425
transform 1 0 8077 0 1 52898
box 0 0 64 64
use contact_9  contact_9_876
timestamp 1624494425
transform 1 0 8076 0 1 52498
box 0 0 66 74
use contact_8  contact_8_876
timestamp 1624494425
transform 1 0 8077 0 1 52503
box 0 0 64 64
use contact_9  contact_9_240
timestamp 1624494425
transform 1 0 7680 0 1 53288
box 0 0 66 74
use contact_8  contact_8_240
timestamp 1624494425
transform 1 0 7681 0 1 53293
box 0 0 64 64
use contact_9  contact_9_870
timestamp 1624494425
transform 1 0 8076 0 1 53288
box 0 0 66 74
use contact_8  contact_8_870
timestamp 1624494425
transform 1 0 8077 0 1 53293
box 0 0 64 64
use contact_9  contact_9_236
timestamp 1624494425
transform 1 0 7680 0 1 54078
box 0 0 66 74
use contact_8  contact_8_236
timestamp 1624494425
transform 1 0 7681 0 1 54083
box 0 0 64 64
use contact_9  contact_9_238
timestamp 1624494425
transform 1 0 7680 0 1 53683
box 0 0 66 74
use contact_8  contact_8_238
timestamp 1624494425
transform 1 0 7681 0 1 53688
box 0 0 64 64
use contact_9  contact_9_864
timestamp 1624494425
transform 1 0 8076 0 1 54078
box 0 0 66 74
use contact_8  contact_8_864
timestamp 1624494425
transform 1 0 8077 0 1 54083
box 0 0 64 64
use contact_9  contact_9_867
timestamp 1624494425
transform 1 0 8076 0 1 53683
box 0 0 66 74
use contact_8  contact_8_867
timestamp 1624494425
transform 1 0 8077 0 1 53688
box 0 0 64 64
use contact_9  contact_9_234
timestamp 1624494425
transform 1 0 7680 0 1 54473
box 0 0 66 74
use contact_8  contact_8_234
timestamp 1624494425
transform 1 0 7681 0 1 54478
box 0 0 64 64
use contact_9  contact_9_861
timestamp 1624494425
transform 1 0 8076 0 1 54473
box 0 0 66 74
use contact_8  contact_8_861
timestamp 1624494425
transform 1 0 8077 0 1 54478
box 0 0 64 64
use contact_9  contact_9_230
timestamp 1624494425
transform 1 0 7680 0 1 55263
box 0 0 66 74
use contact_8  contact_8_230
timestamp 1624494425
transform 1 0 7681 0 1 55268
box 0 0 64 64
use contact_9  contact_9_232
timestamp 1624494425
transform 1 0 7680 0 1 54868
box 0 0 66 74
use contact_8  contact_8_232
timestamp 1624494425
transform 1 0 7681 0 1 54873
box 0 0 64 64
use contact_9  contact_9_855
timestamp 1624494425
transform 1 0 8076 0 1 55263
box 0 0 66 74
use contact_8  contact_8_855
timestamp 1624494425
transform 1 0 8077 0 1 55268
box 0 0 64 64
use contact_9  contact_9_858
timestamp 1624494425
transform 1 0 8076 0 1 54868
box 0 0 66 74
use contact_8  contact_8_858
timestamp 1624494425
transform 1 0 8077 0 1 54873
box 0 0 64 64
use contact_9  contact_9_228
timestamp 1624494425
transform 1 0 7680 0 1 55658
box 0 0 66 74
use contact_8  contact_8_228
timestamp 1624494425
transform 1 0 7681 0 1 55663
box 0 0 64 64
use contact_9  contact_9_852
timestamp 1624494425
transform 1 0 8076 0 1 55658
box 0 0 66 74
use contact_8  contact_8_852
timestamp 1624494425
transform 1 0 8077 0 1 55663
box 0 0 64 64
use contact_16  contact_16_342
timestamp 1624494425
transform 1 0 5864 0 1 55778
box 0 0 66 58
use contact_16  contact_16_343
timestamp 1624494425
transform 1 0 5144 0 1 55868
box 0 0 66 58
use contact_16  contact_16_344
timestamp 1624494425
transform 1 0 4664 0 1 55980
box 0 0 66 58
use contact_8  contact_8_851
timestamp 1624494425
transform 1 0 7299 0 1 56044
box 0 0 64 64
use contact_9  contact_9_851
timestamp 1624494425
transform 1 0 7298 0 1 56039
box 0 0 66 74
use contact_8  contact_8_850
timestamp 1624494425
transform 1 0 6867 0 1 56044
box 0 0 64 64
use contact_9  contact_9_850
timestamp 1624494425
transform 1 0 6866 0 1 56039
box 0 0 66 74
use contact_8  contact_8_227
timestamp 1624494425
transform 1 0 6442 0 1 56102
box 0 0 64 64
use contact_9  contact_9_227
timestamp 1624494425
transform 1 0 6441 0 1 56097
box 0 0 66 74
use contact_16  contact_16_340
timestamp 1624494425
transform 1 0 5144 0 1 56254
box 0 0 66 58
use contact_16  contact_16_341
timestamp 1624494425
transform 1 0 4744 0 1 56142
box 0 0 66 58
use and3_dec  and3_dec_113
timestamp 1624494425
transform 1 0 6203 0 1 56090
box 0 -60 2072 490
use contact_8  contact_8_848
timestamp 1624494425
transform 1 0 7299 0 1 56476
box 0 0 64 64
use contact_9  contact_9_848
timestamp 1624494425
transform 1 0 7298 0 1 56471
box 0 0 66 74
use contact_8  contact_8_847
timestamp 1624494425
transform 1 0 6867 0 1 56476
box 0 0 64 64
use contact_9  contact_9_847
timestamp 1624494425
transform 1 0 6866 0 1 56471
box 0 0 66 74
use contact_8  contact_8_225
timestamp 1624494425
transform 1 0 6442 0 1 56476
box 0 0 64 64
use contact_9  contact_9_225
timestamp 1624494425
transform 1 0 6441 0 1 56471
box 0 0 66 74
use contact_16  contact_16_339
timestamp 1624494425
transform 1 0 5864 0 1 56344
box 0 0 66 58
use contact_16  contact_16_336
timestamp 1624494425
transform 1 0 5864 0 1 56568
box 0 0 66 58
use contact_16  contact_16_337
timestamp 1624494425
transform 1 0 5144 0 1 56658
box 0 0 66 58
use contact_16  contact_16_338
timestamp 1624494425
transform 1 0 4824 0 1 56770
box 0 0 66 58
use and3_dec  and3_dec_112
timestamp 1624494425
transform 1 0 6203 0 -1 56880
box 0 -60 2072 490
use contact_8  contact_8_845
timestamp 1624494425
transform 1 0 7299 0 1 56834
box 0 0 64 64
use contact_9  contact_9_845
timestamp 1624494425
transform 1 0 7298 0 1 56829
box 0 0 66 74
use contact_8  contact_8_844
timestamp 1624494425
transform 1 0 6867 0 1 56834
box 0 0 64 64
use contact_9  contact_9_844
timestamp 1624494425
transform 1 0 6866 0 1 56829
box 0 0 66 74
use contact_8  contact_8_223
timestamp 1624494425
transform 1 0 6442 0 1 56892
box 0 0 64 64
use contact_9  contact_9_223
timestamp 1624494425
transform 1 0 6441 0 1 56887
box 0 0 66 74
use contact_16  contact_16_334
timestamp 1624494425
transform 1 0 5224 0 1 57044
box 0 0 66 58
use contact_16  contact_16_335
timestamp 1624494425
transform 1 0 4584 0 1 56932
box 0 0 66 58
use contact_8  contact_8_842
timestamp 1624494425
transform 1 0 7299 0 1 57266
box 0 0 64 64
use contact_9  contact_9_842
timestamp 1624494425
transform 1 0 7298 0 1 57261
box 0 0 66 74
use contact_8  contact_8_841
timestamp 1624494425
transform 1 0 6867 0 1 57266
box 0 0 64 64
use contact_9  contact_9_841
timestamp 1624494425
transform 1 0 6866 0 1 57261
box 0 0 66 74
use contact_8  contact_8_221
timestamp 1624494425
transform 1 0 6442 0 1 57266
box 0 0 64 64
use contact_9  contact_9_221
timestamp 1624494425
transform 1 0 6441 0 1 57261
box 0 0 66 74
use contact_16  contact_16_330
timestamp 1624494425
transform 1 0 5864 0 1 57358
box 0 0 66 58
use contact_16  contact_16_333
timestamp 1624494425
transform 1 0 5864 0 1 57134
box 0 0 66 58
use and3_dec  and3_dec_110
timestamp 1624494425
transform 1 0 6203 0 -1 57670
box 0 -60 2072 490
use and3_dec  and3_dec_111
timestamp 1624494425
transform 1 0 6203 0 1 56880
box 0 -60 2072 490
use contact_8  contact_8_839
timestamp 1624494425
transform 1 0 7299 0 1 57624
box 0 0 64 64
use contact_9  contact_9_839
timestamp 1624494425
transform 1 0 7298 0 1 57619
box 0 0 66 74
use contact_8  contact_8_838
timestamp 1624494425
transform 1 0 6867 0 1 57624
box 0 0 64 64
use contact_9  contact_9_838
timestamp 1624494425
transform 1 0 6866 0 1 57619
box 0 0 66 74
use contact_16  contact_16_331
timestamp 1624494425
transform 1 0 5224 0 1 57448
box 0 0 66 58
use contact_16  contact_16_332
timestamp 1624494425
transform 1 0 4664 0 1 57560
box 0 0 66 58
use contact_8  contact_8_219
timestamp 1624494425
transform 1 0 6442 0 1 57682
box 0 0 64 64
use contact_9  contact_9_219
timestamp 1624494425
transform 1 0 6441 0 1 57677
box 0 0 66 74
use contact_16  contact_16_328
timestamp 1624494425
transform 1 0 5224 0 1 57834
box 0 0 66 58
use contact_16  contact_16_329
timestamp 1624494425
transform 1 0 4744 0 1 57722
box 0 0 66 58
use and3_dec  and3_dec_109
timestamp 1624494425
transform 1 0 6203 0 1 57670
box 0 -60 2072 490
use contact_8  contact_8_836
timestamp 1624494425
transform 1 0 7299 0 1 58056
box 0 0 64 64
use contact_9  contact_9_836
timestamp 1624494425
transform 1 0 7298 0 1 58051
box 0 0 66 74
use contact_8  contact_8_835
timestamp 1624494425
transform 1 0 6867 0 1 58056
box 0 0 64 64
use contact_9  contact_9_835
timestamp 1624494425
transform 1 0 6866 0 1 58051
box 0 0 66 74
use contact_8  contact_8_217
timestamp 1624494425
transform 1 0 6442 0 1 58056
box 0 0 64 64
use contact_9  contact_9_217
timestamp 1624494425
transform 1 0 6441 0 1 58051
box 0 0 66 74
use contact_16  contact_16_324
timestamp 1624494425
transform 1 0 5864 0 1 58148
box 0 0 66 58
use contact_16  contact_16_327
timestamp 1624494425
transform 1 0 5864 0 1 57924
box 0 0 66 58
use contact_8  contact_8_833
timestamp 1624494425
transform 1 0 7299 0 1 58414
box 0 0 64 64
use contact_9  contact_9_833
timestamp 1624494425
transform 1 0 7298 0 1 58409
box 0 0 66 74
use contact_8  contact_8_832
timestamp 1624494425
transform 1 0 6867 0 1 58414
box 0 0 64 64
use contact_9  contact_9_832
timestamp 1624494425
transform 1 0 6866 0 1 58409
box 0 0 66 74
use contact_9  contact_9_215
timestamp 1624494425
transform 1 0 6441 0 1 58467
box 0 0 66 74
use contact_16  contact_16_325
timestamp 1624494425
transform 1 0 5224 0 1 58238
box 0 0 66 58
use contact_16  contact_16_326
timestamp 1624494425
transform 1 0 4824 0 1 58350
box 0 0 66 58
use and3_dec  and3_dec_107
timestamp 1624494425
transform 1 0 6203 0 1 58460
box 0 -60 2072 490
use and3_dec  and3_dec_108
timestamp 1624494425
transform 1 0 6203 0 -1 58460
box 0 -60 2072 490
use contact_8  contact_8_215
timestamp 1624494425
transform 1 0 6442 0 1 58472
box 0 0 64 64
use contact_16  contact_16_321
timestamp 1624494425
transform 1 0 5864 0 1 58714
box 0 0 66 58
use contact_16  contact_16_322
timestamp 1624494425
transform 1 0 5304 0 1 58624
box 0 0 66 58
use contact_16  contact_16_323
timestamp 1624494425
transform 1 0 4584 0 1 58512
box 0 0 66 58
use contact_8  contact_8_830
timestamp 1624494425
transform 1 0 7299 0 1 58846
box 0 0 64 64
use contact_9  contact_9_830
timestamp 1624494425
transform 1 0 7298 0 1 58841
box 0 0 66 74
use contact_8  contact_8_829
timestamp 1624494425
transform 1 0 6867 0 1 58846
box 0 0 64 64
use contact_9  contact_9_829
timestamp 1624494425
transform 1 0 6866 0 1 58841
box 0 0 66 74
use contact_8  contact_8_213
timestamp 1624494425
transform 1 0 6442 0 1 58846
box 0 0 64 64
use contact_9  contact_9_213
timestamp 1624494425
transform 1 0 6441 0 1 58841
box 0 0 66 74
use contact_16  contact_16_318
timestamp 1624494425
transform 1 0 5864 0 1 58938
box 0 0 66 58
use and3_dec  and3_dec_106
timestamp 1624494425
transform 1 0 6203 0 -1 59250
box 0 -60 2072 490
use contact_9  contact_9_226
timestamp 1624494425
transform 1 0 7680 0 1 56053
box 0 0 66 74
use contact_8  contact_8_226
timestamp 1624494425
transform 1 0 7681 0 1 56058
box 0 0 64 64
use contact_9  contact_9_849
timestamp 1624494425
transform 1 0 8076 0 1 56053
box 0 0 66 74
use contact_8  contact_8_849
timestamp 1624494425
transform 1 0 8077 0 1 56058
box 0 0 64 64
use contact_9  contact_9_222
timestamp 1624494425
transform 1 0 7680 0 1 56843
box 0 0 66 74
use contact_8  contact_8_222
timestamp 1624494425
transform 1 0 7681 0 1 56848
box 0 0 64 64
use contact_9  contact_9_224
timestamp 1624494425
transform 1 0 7680 0 1 56448
box 0 0 66 74
use contact_8  contact_8_224
timestamp 1624494425
transform 1 0 7681 0 1 56453
box 0 0 64 64
use contact_9  contact_9_843
timestamp 1624494425
transform 1 0 8076 0 1 56843
box 0 0 66 74
use contact_8  contact_8_843
timestamp 1624494425
transform 1 0 8077 0 1 56848
box 0 0 64 64
use contact_9  contact_9_846
timestamp 1624494425
transform 1 0 8076 0 1 56448
box 0 0 66 74
use contact_8  contact_8_846
timestamp 1624494425
transform 1 0 8077 0 1 56453
box 0 0 64 64
use contact_9  contact_9_220
timestamp 1624494425
transform 1 0 7680 0 1 57238
box 0 0 66 74
use contact_8  contact_8_220
timestamp 1624494425
transform 1 0 7681 0 1 57243
box 0 0 64 64
use contact_9  contact_9_840
timestamp 1624494425
transform 1 0 8076 0 1 57238
box 0 0 66 74
use contact_8  contact_8_840
timestamp 1624494425
transform 1 0 8077 0 1 57243
box 0 0 64 64
use contact_9  contact_9_216
timestamp 1624494425
transform 1 0 7680 0 1 58028
box 0 0 66 74
use contact_8  contact_8_216
timestamp 1624494425
transform 1 0 7681 0 1 58033
box 0 0 64 64
use contact_9  contact_9_218
timestamp 1624494425
transform 1 0 7680 0 1 57633
box 0 0 66 74
use contact_8  contact_8_218
timestamp 1624494425
transform 1 0 7681 0 1 57638
box 0 0 64 64
use contact_9  contact_9_834
timestamp 1624494425
transform 1 0 8076 0 1 58028
box 0 0 66 74
use contact_8  contact_8_834
timestamp 1624494425
transform 1 0 8077 0 1 58033
box 0 0 64 64
use contact_9  contact_9_837
timestamp 1624494425
transform 1 0 8076 0 1 57633
box 0 0 66 74
use contact_8  contact_8_837
timestamp 1624494425
transform 1 0 8077 0 1 57638
box 0 0 64 64
use contact_9  contact_9_212
timestamp 1624494425
transform 1 0 7680 0 1 58818
box 0 0 66 74
use contact_8  contact_8_212
timestamp 1624494425
transform 1 0 7681 0 1 58823
box 0 0 64 64
use contact_9  contact_9_214
timestamp 1624494425
transform 1 0 7680 0 1 58423
box 0 0 66 74
use contact_8  contact_8_214
timestamp 1624494425
transform 1 0 7681 0 1 58428
box 0 0 64 64
use contact_9  contact_9_828
timestamp 1624494425
transform 1 0 8076 0 1 58818
box 0 0 66 74
use contact_8  contact_8_828
timestamp 1624494425
transform 1 0 8077 0 1 58823
box 0 0 64 64
use contact_9  contact_9_831
timestamp 1624494425
transform 1 0 8076 0 1 58423
box 0 0 66 74
use contact_8  contact_8_831
timestamp 1624494425
transform 1 0 8077 0 1 58428
box 0 0 64 64
use contact_8  contact_8_827
timestamp 1624494425
transform 1 0 7299 0 1 59204
box 0 0 64 64
use contact_9  contact_9_827
timestamp 1624494425
transform 1 0 7298 0 1 59199
box 0 0 66 74
use contact_8  contact_8_826
timestamp 1624494425
transform 1 0 6867 0 1 59204
box 0 0 64 64
use contact_9  contact_9_826
timestamp 1624494425
transform 1 0 6866 0 1 59199
box 0 0 66 74
use contact_8  contact_8_211
timestamp 1624494425
transform 1 0 6442 0 1 59262
box 0 0 64 64
use contact_9  contact_9_211
timestamp 1624494425
transform 1 0 6441 0 1 59257
box 0 0 66 74
use contact_16  contact_16_319
timestamp 1624494425
transform 1 0 5304 0 1 59028
box 0 0 66 58
use contact_16  contact_16_320
timestamp 1624494425
transform 1 0 4664 0 1 59140
box 0 0 66 58
use contact_16  contact_16_315
timestamp 1624494425
transform 1 0 5864 0 1 59504
box 0 0 66 58
use contact_16  contact_16_316
timestamp 1624494425
transform 1 0 5304 0 1 59414
box 0 0 66 58
use contact_16  contact_16_317
timestamp 1624494425
transform 1 0 4744 0 1 59302
box 0 0 66 58
use and3_dec  and3_dec_105
timestamp 1624494425
transform 1 0 6203 0 1 59250
box 0 -60 2072 490
use contact_8  contact_8_824
timestamp 1624494425
transform 1 0 7299 0 1 59636
box 0 0 64 64
use contact_9  contact_9_824
timestamp 1624494425
transform 1 0 7298 0 1 59631
box 0 0 66 74
use contact_8  contact_8_823
timestamp 1624494425
transform 1 0 6867 0 1 59636
box 0 0 64 64
use contact_9  contact_9_823
timestamp 1624494425
transform 1 0 6866 0 1 59631
box 0 0 66 74
use contact_8  contact_8_209
timestamp 1624494425
transform 1 0 6442 0 1 59636
box 0 0 64 64
use contact_9  contact_9_209
timestamp 1624494425
transform 1 0 6441 0 1 59631
box 0 0 66 74
use contact_16  contact_16_312
timestamp 1624494425
transform 1 0 5864 0 1 59728
box 0 0 66 58
use contact_16  contact_16_313
timestamp 1624494425
transform 1 0 5304 0 1 59818
box 0 0 66 58
use contact_8  contact_8_821
timestamp 1624494425
transform 1 0 7299 0 1 59994
box 0 0 64 64
use contact_9  contact_9_821
timestamp 1624494425
transform 1 0 7298 0 1 59989
box 0 0 66 74
use contact_8  contact_8_820
timestamp 1624494425
transform 1 0 6867 0 1 59994
box 0 0 64 64
use contact_9  contact_9_820
timestamp 1624494425
transform 1 0 6866 0 1 59989
box 0 0 66 74
use contact_8  contact_8_207
timestamp 1624494425
transform 1 0 6442 0 1 60052
box 0 0 64 64
use contact_9  contact_9_207
timestamp 1624494425
transform 1 0 6441 0 1 60047
box 0 0 66 74
use contact_16  contact_16_311
timestamp 1624494425
transform 1 0 4584 0 1 60092
box 0 0 66 58
use contact_16  contact_16_314
timestamp 1624494425
transform 1 0 4824 0 1 59930
box 0 0 66 58
use and3_dec  and3_dec_103
timestamp 1624494425
transform 1 0 6203 0 1 60040
box 0 -60 2072 490
use and3_dec  and3_dec_104
timestamp 1624494425
transform 1 0 6203 0 -1 60040
box 0 -60 2072 490
use contact_16  contact_16_309
timestamp 1624494425
transform 1 0 5864 0 1 60294
box 0 0 66 58
use contact_16  contact_16_310
timestamp 1624494425
transform 1 0 5384 0 1 60204
box 0 0 66 58
use contact_8  contact_8_818
timestamp 1624494425
transform 1 0 7299 0 1 60426
box 0 0 64 64
use contact_9  contact_9_818
timestamp 1624494425
transform 1 0 7298 0 1 60421
box 0 0 66 74
use contact_8  contact_8_817
timestamp 1624494425
transform 1 0 6867 0 1 60426
box 0 0 64 64
use contact_9  contact_9_817
timestamp 1624494425
transform 1 0 6866 0 1 60421
box 0 0 66 74
use contact_8  contact_8_205
timestamp 1624494425
transform 1 0 6442 0 1 60426
box 0 0 64 64
use contact_9  contact_9_205
timestamp 1624494425
transform 1 0 6441 0 1 60421
box 0 0 66 74
use contact_16  contact_16_306
timestamp 1624494425
transform 1 0 5864 0 1 60518
box 0 0 66 58
use contact_16  contact_16_307
timestamp 1624494425
transform 1 0 5384 0 1 60608
box 0 0 66 58
use and3_dec  and3_dec_102
timestamp 1624494425
transform 1 0 6203 0 -1 60830
box 0 -60 2072 490
use contact_8  contact_8_815
timestamp 1624494425
transform 1 0 7299 0 1 60784
box 0 0 64 64
use contact_9  contact_9_815
timestamp 1624494425
transform 1 0 7298 0 1 60779
box 0 0 66 74
use contact_8  contact_8_814
timestamp 1624494425
transform 1 0 6867 0 1 60784
box 0 0 64 64
use contact_9  contact_9_814
timestamp 1624494425
transform 1 0 6866 0 1 60779
box 0 0 66 74
use contact_8  contact_8_203
timestamp 1624494425
transform 1 0 6442 0 1 60842
box 0 0 64 64
use contact_9  contact_9_203
timestamp 1624494425
transform 1 0 6441 0 1 60837
box 0 0 66 74
use contact_16  contact_16_305
timestamp 1624494425
transform 1 0 4744 0 1 60882
box 0 0 66 58
use contact_16  contact_16_308
timestamp 1624494425
transform 1 0 4664 0 1 60720
box 0 0 66 58
use contact_16  contact_16_303
timestamp 1624494425
transform 1 0 5864 0 1 61084
box 0 0 66 58
use contact_16  contact_16_304
timestamp 1624494425
transform 1 0 5384 0 1 60994
box 0 0 66 58
use and3_dec  and3_dec_100
timestamp 1624494425
transform 1 0 6203 0 -1 61620
box 0 -60 2072 490
use and3_dec  and3_dec_101
timestamp 1624494425
transform 1 0 6203 0 1 60830
box 0 -60 2072 490
use contact_8  contact_8_812
timestamp 1624494425
transform 1 0 7299 0 1 61216
box 0 0 64 64
use contact_9  contact_9_812
timestamp 1624494425
transform 1 0 7298 0 1 61211
box 0 0 66 74
use contact_8  contact_8_811
timestamp 1624494425
transform 1 0 6867 0 1 61216
box 0 0 64 64
use contact_9  contact_9_811
timestamp 1624494425
transform 1 0 6866 0 1 61211
box 0 0 66 74
use contact_8  contact_8_201
timestamp 1624494425
transform 1 0 6442 0 1 61216
box 0 0 64 64
use contact_9  contact_9_201
timestamp 1624494425
transform 1 0 6441 0 1 61211
box 0 0 66 74
use contact_16  contact_16_300
timestamp 1624494425
transform 1 0 5864 0 1 61308
box 0 0 66 58
use contact_16  contact_16_301
timestamp 1624494425
transform 1 0 5384 0 1 61398
box 0 0 66 58
use contact_8  contact_8_809
timestamp 1624494425
transform 1 0 7299 0 1 61574
box 0 0 64 64
use contact_9  contact_9_809
timestamp 1624494425
transform 1 0 7298 0 1 61569
box 0 0 66 74
use contact_8  contact_8_808
timestamp 1624494425
transform 1 0 6867 0 1 61574
box 0 0 64 64
use contact_9  contact_9_808
timestamp 1624494425
transform 1 0 6866 0 1 61569
box 0 0 66 74
use contact_8  contact_8_199
timestamp 1624494425
transform 1 0 6442 0 1 61632
box 0 0 64 64
use contact_9  contact_9_199
timestamp 1624494425
transform 1 0 6441 0 1 61627
box 0 0 66 74
use contact_16  contact_16_299
timestamp 1624494425
transform 1 0 4584 0 1 61672
box 0 0 66 58
use contact_16  contact_16_302
timestamp 1624494425
transform 1 0 4824 0 1 61510
box 0 0 66 58
use and3_dec  and3_dec_99
timestamp 1624494425
transform 1 0 6203 0 1 61620
box 0 -60 2072 490
use contact_8  contact_8_806
timestamp 1624494425
transform 1 0 7299 0 1 62006
box 0 0 64 64
use contact_9  contact_9_806
timestamp 1624494425
transform 1 0 7298 0 1 62001
box 0 0 66 74
use contact_8  contact_8_805
timestamp 1624494425
transform 1 0 6867 0 1 62006
box 0 0 64 64
use contact_9  contact_9_805
timestamp 1624494425
transform 1 0 6866 0 1 62001
box 0 0 66 74
use contact_8  contact_8_197
timestamp 1624494425
transform 1 0 6442 0 1 62006
box 0 0 64 64
use contact_9  contact_9_197
timestamp 1624494425
transform 1 0 6441 0 1 62001
box 0 0 66 74
use contact_16  contact_16_297
timestamp 1624494425
transform 1 0 5864 0 1 61874
box 0 0 66 58
use contact_16  contact_16_298
timestamp 1624494425
transform 1 0 5464 0 1 61784
box 0 0 66 58
use contact_16  contact_16_294
timestamp 1624494425
transform 1 0 5864 0 1 62098
box 0 0 66 58
use contact_16  contact_16_295
timestamp 1624494425
transform 1 0 5464 0 1 62188
box 0 0 66 58
use and3_dec  and3_dec_98
timestamp 1624494425
transform 1 0 6203 0 -1 62410
box 0 -60 2072 490
use contact_9  contact_9_208
timestamp 1624494425
transform 1 0 7680 0 1 59608
box 0 0 66 74
use contact_8  contact_8_208
timestamp 1624494425
transform 1 0 7681 0 1 59613
box 0 0 64 64
use contact_9  contact_9_210
timestamp 1624494425
transform 1 0 7680 0 1 59213
box 0 0 66 74
use contact_8  contact_8_210
timestamp 1624494425
transform 1 0 7681 0 1 59218
box 0 0 64 64
use contact_9  contact_9_822
timestamp 1624494425
transform 1 0 8076 0 1 59608
box 0 0 66 74
use contact_8  contact_8_822
timestamp 1624494425
transform 1 0 8077 0 1 59613
box 0 0 64 64
use contact_9  contact_9_825
timestamp 1624494425
transform 1 0 8076 0 1 59213
box 0 0 66 74
use contact_8  contact_8_825
timestamp 1624494425
transform 1 0 8077 0 1 59218
box 0 0 64 64
use contact_9  contact_9_206
timestamp 1624494425
transform 1 0 7680 0 1 60003
box 0 0 66 74
use contact_8  contact_8_206
timestamp 1624494425
transform 1 0 7681 0 1 60008
box 0 0 64 64
use contact_9  contact_9_819
timestamp 1624494425
transform 1 0 8076 0 1 60003
box 0 0 66 74
use contact_8  contact_8_819
timestamp 1624494425
transform 1 0 8077 0 1 60008
box 0 0 64 64
use contact_9  contact_9_202
timestamp 1624494425
transform 1 0 7680 0 1 60793
box 0 0 66 74
use contact_8  contact_8_202
timestamp 1624494425
transform 1 0 7681 0 1 60798
box 0 0 64 64
use contact_9  contact_9_204
timestamp 1624494425
transform 1 0 7680 0 1 60398
box 0 0 66 74
use contact_8  contact_8_204
timestamp 1624494425
transform 1 0 7681 0 1 60403
box 0 0 64 64
use contact_9  contact_9_813
timestamp 1624494425
transform 1 0 8076 0 1 60793
box 0 0 66 74
use contact_8  contact_8_813
timestamp 1624494425
transform 1 0 8077 0 1 60798
box 0 0 64 64
use contact_9  contact_9_816
timestamp 1624494425
transform 1 0 8076 0 1 60398
box 0 0 66 74
use contact_8  contact_8_816
timestamp 1624494425
transform 1 0 8077 0 1 60403
box 0 0 64 64
use contact_9  contact_9_200
timestamp 1624494425
transform 1 0 7680 0 1 61188
box 0 0 66 74
use contact_8  contact_8_200
timestamp 1624494425
transform 1 0 7681 0 1 61193
box 0 0 64 64
use contact_9  contact_9_810
timestamp 1624494425
transform 1 0 8076 0 1 61188
box 0 0 66 74
use contact_8  contact_8_810
timestamp 1624494425
transform 1 0 8077 0 1 61193
box 0 0 64 64
use contact_9  contact_9_196
timestamp 1624494425
transform 1 0 7680 0 1 61978
box 0 0 66 74
use contact_8  contact_8_196
timestamp 1624494425
transform 1 0 7681 0 1 61983
box 0 0 64 64
use contact_9  contact_9_198
timestamp 1624494425
transform 1 0 7680 0 1 61583
box 0 0 66 74
use contact_8  contact_8_198
timestamp 1624494425
transform 1 0 7681 0 1 61588
box 0 0 64 64
use contact_9  contact_9_804
timestamp 1624494425
transform 1 0 8076 0 1 61978
box 0 0 66 74
use contact_8  contact_8_804
timestamp 1624494425
transform 1 0 8077 0 1 61983
box 0 0 64 64
use contact_9  contact_9_807
timestamp 1624494425
transform 1 0 8076 0 1 61583
box 0 0 66 74
use contact_8  contact_8_807
timestamp 1624494425
transform 1 0 8077 0 1 61588
box 0 0 64 64
use contact_8  contact_8_803
timestamp 1624494425
transform 1 0 7299 0 1 62364
box 0 0 64 64
use contact_9  contact_9_803
timestamp 1624494425
transform 1 0 7298 0 1 62359
box 0 0 66 74
use contact_8  contact_8_802
timestamp 1624494425
transform 1 0 6867 0 1 62364
box 0 0 64 64
use contact_9  contact_9_802
timestamp 1624494425
transform 1 0 6866 0 1 62359
box 0 0 66 74
use contact_8  contact_8_195
timestamp 1624494425
transform 1 0 6442 0 1 62422
box 0 0 64 64
use contact_9  contact_9_195
timestamp 1624494425
transform 1 0 6441 0 1 62417
box 0 0 66 74
use contact_16  contact_16_293
timestamp 1624494425
transform 1 0 4744 0 1 62462
box 0 0 66 58
use contact_16  contact_16_296
timestamp 1624494425
transform 1 0 4664 0 1 62300
box 0 0 66 58
use contact_8  contact_8_800
timestamp 1624494425
transform 1 0 7299 0 1 62796
box 0 0 64 64
use contact_9  contact_9_800
timestamp 1624494425
transform 1 0 7298 0 1 62791
box 0 0 66 74
use contact_8  contact_8_799
timestamp 1624494425
transform 1 0 6867 0 1 62796
box 0 0 64 64
use contact_9  contact_9_799
timestamp 1624494425
transform 1 0 6866 0 1 62791
box 0 0 66 74
use contact_8  contact_8_193
timestamp 1624494425
transform 1 0 6442 0 1 62796
box 0 0 64 64
use contact_9  contact_9_193
timestamp 1624494425
transform 1 0 6441 0 1 62791
box 0 0 66 74
use contact_16  contact_16_291
timestamp 1624494425
transform 1 0 5864 0 1 62664
box 0 0 66 58
use contact_16  contact_16_292
timestamp 1624494425
transform 1 0 5464 0 1 62574
box 0 0 66 58
use and3_dec  and3_dec_96
timestamp 1624494425
transform 1 0 6203 0 -1 63200
box 0 -60 2072 490
use and3_dec  and3_dec_97
timestamp 1624494425
transform 1 0 6203 0 1 62410
box 0 -60 2072 490
use contact_16  contact_16_288
timestamp 1624494425
transform 1 0 5864 0 1 62888
box 0 0 66 58
use contact_16  contact_16_289
timestamp 1624494425
transform 1 0 5464 0 1 62978
box 0 0 66 58
use contact_16  contact_16_290
timestamp 1624494425
transform 1 0 4824 0 1 63090
box 0 0 66 58
use contact_8  contact_8_797
timestamp 1624494425
transform 1 0 7299 0 1 63154
box 0 0 64 64
use contact_9  contact_9_797
timestamp 1624494425
transform 1 0 7298 0 1 63149
box 0 0 66 74
use contact_8  contact_8_796
timestamp 1624494425
transform 1 0 6867 0 1 63154
box 0 0 64 64
use contact_9  contact_9_796
timestamp 1624494425
transform 1 0 6866 0 1 63149
box 0 0 66 74
use contact_8  contact_8_191
timestamp 1624494425
transform 1 0 6442 0 1 63212
box 0 0 64 64
use contact_9  contact_9_191
timestamp 1624494425
transform 1 0 6441 0 1 63207
box 0 0 66 74
use contact_16  contact_16_286
timestamp 1624494425
transform 1 0 4904 0 1 63364
box 0 0 66 58
use contact_16  contact_16_287
timestamp 1624494425
transform 1 0 4584 0 1 63252
box 0 0 66 58
use and3_dec  and3_dec_95
timestamp 1624494425
transform 1 0 6203 0 1 63200
box 0 -60 2072 490
use contact_8  contact_8_794
timestamp 1624494425
transform 1 0 7299 0 1 63586
box 0 0 64 64
use contact_9  contact_9_794
timestamp 1624494425
transform 1 0 7298 0 1 63581
box 0 0 66 74
use contact_8  contact_8_793
timestamp 1624494425
transform 1 0 6867 0 1 63586
box 0 0 64 64
use contact_9  contact_9_793
timestamp 1624494425
transform 1 0 6866 0 1 63581
box 0 0 66 74
use contact_8  contact_8_189
timestamp 1624494425
transform 1 0 6442 0 1 63586
box 0 0 64 64
use contact_9  contact_9_189
timestamp 1624494425
transform 1 0 6441 0 1 63581
box 0 0 66 74
use contact_16  contact_16_285
timestamp 1624494425
transform 1 0 5944 0 1 63454
box 0 0 66 58
use contact_16  contact_16_282
timestamp 1624494425
transform 1 0 5944 0 1 63678
box 0 0 66 58
use contact_16  contact_16_283
timestamp 1624494425
transform 1 0 4904 0 1 63768
box 0 0 66 58
use contact_16  contact_16_284
timestamp 1624494425
transform 1 0 4664 0 1 63880
box 0 0 66 58
use and3_dec  and3_dec_93
timestamp 1624494425
transform 1 0 6203 0 1 63990
box 0 -60 2072 490
use and3_dec  and3_dec_94
timestamp 1624494425
transform 1 0 6203 0 -1 63990
box 0 -60 2072 490
use contact_8  contact_8_791
timestamp 1624494425
transform 1 0 7299 0 1 63944
box 0 0 64 64
use contact_9  contact_9_791
timestamp 1624494425
transform 1 0 7298 0 1 63939
box 0 0 66 74
use contact_8  contact_8_790
timestamp 1624494425
transform 1 0 6867 0 1 63944
box 0 0 64 64
use contact_9  contact_9_790
timestamp 1624494425
transform 1 0 6866 0 1 63939
box 0 0 66 74
use contact_8  contact_8_187
timestamp 1624494425
transform 1 0 6442 0 1 64002
box 0 0 64 64
use contact_9  contact_9_187
timestamp 1624494425
transform 1 0 6441 0 1 63997
box 0 0 66 74
use contact_16  contact_16_280
timestamp 1624494425
transform 1 0 4904 0 1 64154
box 0 0 66 58
use contact_16  contact_16_281
timestamp 1624494425
transform 1 0 4744 0 1 64042
box 0 0 66 58
use contact_8  contact_8_788
timestamp 1624494425
transform 1 0 7299 0 1 64376
box 0 0 64 64
use contact_9  contact_9_788
timestamp 1624494425
transform 1 0 7298 0 1 64371
box 0 0 66 74
use contact_8  contact_8_787
timestamp 1624494425
transform 1 0 6867 0 1 64376
box 0 0 64 64
use contact_9  contact_9_787
timestamp 1624494425
transform 1 0 6866 0 1 64371
box 0 0 66 74
use contact_8  contact_8_185
timestamp 1624494425
transform 1 0 6442 0 1 64376
box 0 0 64 64
use contact_9  contact_9_185
timestamp 1624494425
transform 1 0 6441 0 1 64371
box 0 0 66 74
use contact_16  contact_16_276
timestamp 1624494425
transform 1 0 5944 0 1 64468
box 0 0 66 58
use contact_16  contact_16_279
timestamp 1624494425
transform 1 0 5944 0 1 64244
box 0 0 66 58
use and3_dec  and3_dec_92
timestamp 1624494425
transform 1 0 6203 0 -1 64780
box 0 -60 2072 490
use contact_8  contact_8_785
timestamp 1624494425
transform 1 0 7299 0 1 64734
box 0 0 64 64
use contact_9  contact_9_785
timestamp 1624494425
transform 1 0 7298 0 1 64729
box 0 0 66 74
use contact_8  contact_8_784
timestamp 1624494425
transform 1 0 6867 0 1 64734
box 0 0 64 64
use contact_9  contact_9_784
timestamp 1624494425
transform 1 0 6866 0 1 64729
box 0 0 66 74
use contact_16  contact_16_277
timestamp 1624494425
transform 1 0 4904 0 1 64558
box 0 0 66 58
use contact_16  contact_16_278
timestamp 1624494425
transform 1 0 4824 0 1 64670
box 0 0 66 58
use contact_8  contact_8_183
timestamp 1624494425
transform 1 0 6442 0 1 64792
box 0 0 64 64
use contact_9  contact_9_183
timestamp 1624494425
transform 1 0 6441 0 1 64787
box 0 0 66 74
use contact_16  contact_16_274
timestamp 1624494425
transform 1 0 4984 0 1 64944
box 0 0 66 58
use contact_16  contact_16_275
timestamp 1624494425
transform 1 0 4584 0 1 64832
box 0 0 66 58
use and3_dec  and3_dec_91
timestamp 1624494425
transform 1 0 6203 0 1 64780
box 0 -60 2072 490
use contact_8  contact_8_782
timestamp 1624494425
transform 1 0 7299 0 1 65166
box 0 0 64 64
use contact_9  contact_9_782
timestamp 1624494425
transform 1 0 7298 0 1 65161
box 0 0 66 74
use contact_8  contact_8_781
timestamp 1624494425
transform 1 0 6867 0 1 65166
box 0 0 64 64
use contact_9  contact_9_781
timestamp 1624494425
transform 1 0 6866 0 1 65161
box 0 0 66 74
use contact_8  contact_8_181
timestamp 1624494425
transform 1 0 6442 0 1 65166
box 0 0 64 64
use contact_9  contact_9_181
timestamp 1624494425
transform 1 0 6441 0 1 65161
box 0 0 66 74
use contact_16  contact_16_270
timestamp 1624494425
transform 1 0 5944 0 1 65258
box 0 0 66 58
use contact_16  contact_16_273
timestamp 1624494425
transform 1 0 5944 0 1 65034
box 0 0 66 58
use contact_8  contact_8_779
timestamp 1624494425
transform 1 0 7299 0 1 65524
box 0 0 64 64
use contact_9  contact_9_779
timestamp 1624494425
transform 1 0 7298 0 1 65519
box 0 0 66 74
use contact_8  contact_8_778
timestamp 1624494425
transform 1 0 6867 0 1 65524
box 0 0 64 64
use contact_9  contact_9_778
timestamp 1624494425
transform 1 0 6866 0 1 65519
box 0 0 66 74
use contact_16  contact_16_271
timestamp 1624494425
transform 1 0 4984 0 1 65348
box 0 0 66 58
use contact_16  contact_16_272
timestamp 1624494425
transform 1 0 4664 0 1 65460
box 0 0 66 58
use and3_dec  and3_dec_89
timestamp 1624494425
transform 1 0 6203 0 1 65570
box 0 -60 2072 490
use and3_dec  and3_dec_90
timestamp 1624494425
transform 1 0 6203 0 -1 65570
box 0 -60 2072 490
use contact_9  contact_9_192
timestamp 1624494425
transform 1 0 7680 0 1 62768
box 0 0 66 74
use contact_8  contact_8_192
timestamp 1624494425
transform 1 0 7681 0 1 62773
box 0 0 64 64
use contact_9  contact_9_194
timestamp 1624494425
transform 1 0 7680 0 1 62373
box 0 0 66 74
use contact_8  contact_8_194
timestamp 1624494425
transform 1 0 7681 0 1 62378
box 0 0 64 64
use contact_9  contact_9_798
timestamp 1624494425
transform 1 0 8076 0 1 62768
box 0 0 66 74
use contact_8  contact_8_798
timestamp 1624494425
transform 1 0 8077 0 1 62773
box 0 0 64 64
use contact_9  contact_9_801
timestamp 1624494425
transform 1 0 8076 0 1 62373
box 0 0 66 74
use contact_8  contact_8_801
timestamp 1624494425
transform 1 0 8077 0 1 62378
box 0 0 64 64
use contact_9  contact_9_190
timestamp 1624494425
transform 1 0 7680 0 1 63163
box 0 0 66 74
use contact_8  contact_8_190
timestamp 1624494425
transform 1 0 7681 0 1 63168
box 0 0 64 64
use contact_9  contact_9_795
timestamp 1624494425
transform 1 0 8076 0 1 63163
box 0 0 66 74
use contact_8  contact_8_795
timestamp 1624494425
transform 1 0 8077 0 1 63168
box 0 0 64 64
use contact_9  contact_9_186
timestamp 1624494425
transform 1 0 7680 0 1 63953
box 0 0 66 74
use contact_8  contact_8_186
timestamp 1624494425
transform 1 0 7681 0 1 63958
box 0 0 64 64
use contact_9  contact_9_188
timestamp 1624494425
transform 1 0 7680 0 1 63558
box 0 0 66 74
use contact_8  contact_8_188
timestamp 1624494425
transform 1 0 7681 0 1 63563
box 0 0 64 64
use contact_9  contact_9_789
timestamp 1624494425
transform 1 0 8076 0 1 63953
box 0 0 66 74
use contact_8  contact_8_789
timestamp 1624494425
transform 1 0 8077 0 1 63958
box 0 0 64 64
use contact_9  contact_9_792
timestamp 1624494425
transform 1 0 8076 0 1 63558
box 0 0 66 74
use contact_8  contact_8_792
timestamp 1624494425
transform 1 0 8077 0 1 63563
box 0 0 64 64
use contact_9  contact_9_184
timestamp 1624494425
transform 1 0 7680 0 1 64348
box 0 0 66 74
use contact_8  contact_8_184
timestamp 1624494425
transform 1 0 7681 0 1 64353
box 0 0 64 64
use contact_9  contact_9_786
timestamp 1624494425
transform 1 0 8076 0 1 64348
box 0 0 66 74
use contact_8  contact_8_786
timestamp 1624494425
transform 1 0 8077 0 1 64353
box 0 0 64 64
use contact_9  contact_9_180
timestamp 1624494425
transform 1 0 7680 0 1 65138
box 0 0 66 74
use contact_8  contact_8_180
timestamp 1624494425
transform 1 0 7681 0 1 65143
box 0 0 64 64
use contact_9  contact_9_182
timestamp 1624494425
transform 1 0 7680 0 1 64743
box 0 0 66 74
use contact_8  contact_8_182
timestamp 1624494425
transform 1 0 7681 0 1 64748
box 0 0 64 64
use contact_9  contact_9_780
timestamp 1624494425
transform 1 0 8076 0 1 65138
box 0 0 66 74
use contact_8  contact_8_780
timestamp 1624494425
transform 1 0 8077 0 1 65143
box 0 0 64 64
use contact_9  contact_9_783
timestamp 1624494425
transform 1 0 8076 0 1 64743
box 0 0 66 74
use contact_8  contact_8_783
timestamp 1624494425
transform 1 0 8077 0 1 64748
box 0 0 64 64
use contact_9  contact_9_178
timestamp 1624494425
transform 1 0 7680 0 1 65533
box 0 0 66 74
use contact_8  contact_8_178
timestamp 1624494425
transform 1 0 7681 0 1 65538
box 0 0 64 64
use contact_9  contact_9_777
timestamp 1624494425
transform 1 0 8076 0 1 65533
box 0 0 66 74
use contact_8  contact_8_777
timestamp 1624494425
transform 1 0 8077 0 1 65538
box 0 0 64 64
use contact_8  contact_8_179
timestamp 1624494425
transform 1 0 6442 0 1 65582
box 0 0 64 64
use contact_9  contact_9_179
timestamp 1624494425
transform 1 0 6441 0 1 65577
box 0 0 66 74
use contact_16  contact_16_267
timestamp 1624494425
transform 1 0 5944 0 1 65824
box 0 0 66 58
use contact_16  contact_16_268
timestamp 1624494425
transform 1 0 4984 0 1 65734
box 0 0 66 58
use contact_16  contact_16_269
timestamp 1624494425
transform 1 0 4744 0 1 65622
box 0 0 66 58
use contact_8  contact_8_776
timestamp 1624494425
transform 1 0 7299 0 1 65956
box 0 0 64 64
use contact_9  contact_9_776
timestamp 1624494425
transform 1 0 7298 0 1 65951
box 0 0 66 74
use contact_8  contact_8_775
timestamp 1624494425
transform 1 0 6867 0 1 65956
box 0 0 64 64
use contact_9  contact_9_775
timestamp 1624494425
transform 1 0 6866 0 1 65951
box 0 0 66 74
use contact_8  contact_8_177
timestamp 1624494425
transform 1 0 6442 0 1 65956
box 0 0 64 64
use contact_9  contact_9_177
timestamp 1624494425
transform 1 0 6441 0 1 65951
box 0 0 66 74
use contact_16  contact_16_264
timestamp 1624494425
transform 1 0 5944 0 1 66048
box 0 0 66 58
use and3_dec  and3_dec_88
timestamp 1624494425
transform 1 0 6203 0 -1 66360
box 0 -60 2072 490
use contact_8  contact_8_773
timestamp 1624494425
transform 1 0 7299 0 1 66314
box 0 0 64 64
use contact_9  contact_9_773
timestamp 1624494425
transform 1 0 7298 0 1 66309
box 0 0 66 74
use contact_8  contact_8_772
timestamp 1624494425
transform 1 0 6867 0 1 66314
box 0 0 64 64
use contact_9  contact_9_772
timestamp 1624494425
transform 1 0 6866 0 1 66309
box 0 0 66 74
use contact_8  contact_8_175
timestamp 1624494425
transform 1 0 6442 0 1 66372
box 0 0 64 64
use contact_9  contact_9_175
timestamp 1624494425
transform 1 0 6441 0 1 66367
box 0 0 66 74
use contact_16  contact_16_265
timestamp 1624494425
transform 1 0 4984 0 1 66138
box 0 0 66 58
use contact_16  contact_16_266
timestamp 1624494425
transform 1 0 4824 0 1 66250
box 0 0 66 58
use contact_16  contact_16_261
timestamp 1624494425
transform 1 0 5944 0 1 66614
box 0 0 66 58
use contact_16  contact_16_262
timestamp 1624494425
transform 1 0 5064 0 1 66524
box 0 0 66 58
use contact_16  contact_16_263
timestamp 1624494425
transform 1 0 4584 0 1 66412
box 0 0 66 58
use and3_dec  and3_dec_86
timestamp 1624494425
transform 1 0 6203 0 -1 67150
box 0 -60 2072 490
use and3_dec  and3_dec_87
timestamp 1624494425
transform 1 0 6203 0 1 66360
box 0 -60 2072 490
use contact_8  contact_8_770
timestamp 1624494425
transform 1 0 7299 0 1 66746
box 0 0 64 64
use contact_9  contact_9_770
timestamp 1624494425
transform 1 0 7298 0 1 66741
box 0 0 66 74
use contact_8  contact_8_769
timestamp 1624494425
transform 1 0 6867 0 1 66746
box 0 0 64 64
use contact_9  contact_9_769
timestamp 1624494425
transform 1 0 6866 0 1 66741
box 0 0 66 74
use contact_8  contact_8_173
timestamp 1624494425
transform 1 0 6442 0 1 66746
box 0 0 64 64
use contact_9  contact_9_173
timestamp 1624494425
transform 1 0 6441 0 1 66741
box 0 0 66 74
use contact_16  contact_16_258
timestamp 1624494425
transform 1 0 5944 0 1 66838
box 0 0 66 58
use contact_16  contact_16_259
timestamp 1624494425
transform 1 0 5064 0 1 66928
box 0 0 66 58
use contact_8  contact_8_767
timestamp 1624494425
transform 1 0 7299 0 1 67104
box 0 0 64 64
use contact_9  contact_9_767
timestamp 1624494425
transform 1 0 7298 0 1 67099
box 0 0 66 74
use contact_8  contact_8_766
timestamp 1624494425
transform 1 0 6867 0 1 67104
box 0 0 64 64
use contact_9  contact_9_766
timestamp 1624494425
transform 1 0 6866 0 1 67099
box 0 0 66 74
use contact_8  contact_8_171
timestamp 1624494425
transform 1 0 6442 0 1 67162
box 0 0 64 64
use contact_9  contact_9_171
timestamp 1624494425
transform 1 0 6441 0 1 67157
box 0 0 66 74
use contact_16  contact_16_257
timestamp 1624494425
transform 1 0 4744 0 1 67202
box 0 0 66 58
use contact_16  contact_16_260
timestamp 1624494425
transform 1 0 4664 0 1 67040
box 0 0 66 58
use and3_dec  and3_dec_85
timestamp 1624494425
transform 1 0 6203 0 1 67150
box 0 -60 2072 490
use contact_16  contact_16_255
timestamp 1624494425
transform 1 0 5944 0 1 67404
box 0 0 66 58
use contact_16  contact_16_256
timestamp 1624494425
transform 1 0 5064 0 1 67314
box 0 0 66 58
use contact_8  contact_8_764
timestamp 1624494425
transform 1 0 7299 0 1 67536
box 0 0 64 64
use contact_9  contact_9_764
timestamp 1624494425
transform 1 0 7298 0 1 67531
box 0 0 66 74
use contact_8  contact_8_763
timestamp 1624494425
transform 1 0 6867 0 1 67536
box 0 0 64 64
use contact_9  contact_9_763
timestamp 1624494425
transform 1 0 6866 0 1 67531
box 0 0 66 74
use contact_8  contact_8_169
timestamp 1624494425
transform 1 0 6442 0 1 67536
box 0 0 64 64
use contact_9  contact_9_169
timestamp 1624494425
transform 1 0 6441 0 1 67531
box 0 0 66 74
use contact_16  contact_16_252
timestamp 1624494425
transform 1 0 5944 0 1 67628
box 0 0 66 58
use contact_16  contact_16_253
timestamp 1624494425
transform 1 0 5064 0 1 67718
box 0 0 66 58
use and3_dec  and3_dec_84
timestamp 1624494425
transform 1 0 6203 0 -1 67940
box 0 -60 2072 490
use contact_8  contact_8_761
timestamp 1624494425
transform 1 0 7299 0 1 67894
box 0 0 64 64
use contact_9  contact_9_761
timestamp 1624494425
transform 1 0 7298 0 1 67889
box 0 0 66 74
use contact_8  contact_8_760
timestamp 1624494425
transform 1 0 6867 0 1 67894
box 0 0 64 64
use contact_9  contact_9_760
timestamp 1624494425
transform 1 0 6866 0 1 67889
box 0 0 66 74
use contact_8  contact_8_167
timestamp 1624494425
transform 1 0 6442 0 1 67952
box 0 0 64 64
use contact_9  contact_9_167
timestamp 1624494425
transform 1 0 6441 0 1 67947
box 0 0 66 74
use contact_16  contact_16_251
timestamp 1624494425
transform 1 0 4584 0 1 67992
box 0 0 66 58
use contact_16  contact_16_254
timestamp 1624494425
transform 1 0 4824 0 1 67830
box 0 0 66 58
use contact_16  contact_16_249
timestamp 1624494425
transform 1 0 5944 0 1 68194
box 0 0 66 58
use contact_16  contact_16_250
timestamp 1624494425
transform 1 0 5144 0 1 68104
box 0 0 66 58
use and3_dec  and3_dec_82
timestamp 1624494425
transform 1 0 6203 0 -1 68730
box 0 -60 2072 490
use and3_dec  and3_dec_83
timestamp 1624494425
transform 1 0 6203 0 1 67940
box 0 -60 2072 490
use contact_8  contact_8_758
timestamp 1624494425
transform 1 0 7299 0 1 68326
box 0 0 64 64
use contact_9  contact_9_758
timestamp 1624494425
transform 1 0 7298 0 1 68321
box 0 0 66 74
use contact_8  contact_8_757
timestamp 1624494425
transform 1 0 6867 0 1 68326
box 0 0 64 64
use contact_9  contact_9_757
timestamp 1624494425
transform 1 0 6866 0 1 68321
box 0 0 66 74
use contact_8  contact_8_165
timestamp 1624494425
transform 1 0 6442 0 1 68326
box 0 0 64 64
use contact_9  contact_9_165
timestamp 1624494425
transform 1 0 6441 0 1 68321
box 0 0 66 74
use contact_16  contact_16_246
timestamp 1624494425
transform 1 0 5944 0 1 68418
box 0 0 66 58
use contact_16  contact_16_247
timestamp 1624494425
transform 1 0 5144 0 1 68508
box 0 0 66 58
use contact_8  contact_8_755
timestamp 1624494425
transform 1 0 7299 0 1 68684
box 0 0 64 64
use contact_9  contact_9_755
timestamp 1624494425
transform 1 0 7298 0 1 68679
box 0 0 66 74
use contact_8  contact_8_754
timestamp 1624494425
transform 1 0 6867 0 1 68684
box 0 0 64 64
use contact_9  contact_9_754
timestamp 1624494425
transform 1 0 6866 0 1 68679
box 0 0 66 74
use contact_8  contact_8_163
timestamp 1624494425
transform 1 0 6442 0 1 68742
box 0 0 64 64
use contact_9  contact_9_163
timestamp 1624494425
transform 1 0 6441 0 1 68737
box 0 0 66 74
use contact_16  contact_16_245
timestamp 1624494425
transform 1 0 4744 0 1 68782
box 0 0 66 58
use contact_16  contact_16_248
timestamp 1624494425
transform 1 0 4664 0 1 68620
box 0 0 66 58
use and3_dec  and3_dec_81
timestamp 1624494425
transform 1 0 6203 0 1 68730
box 0 -60 2072 490
use contact_9  contact_9_176
timestamp 1624494425
transform 1 0 7680 0 1 65928
box 0 0 66 74
use contact_8  contact_8_176
timestamp 1624494425
transform 1 0 7681 0 1 65933
box 0 0 64 64
use contact_9  contact_9_774
timestamp 1624494425
transform 1 0 8076 0 1 65928
box 0 0 66 74
use contact_8  contact_8_774
timestamp 1624494425
transform 1 0 8077 0 1 65933
box 0 0 64 64
use contact_9  contact_9_172
timestamp 1624494425
transform 1 0 7680 0 1 66718
box 0 0 66 74
use contact_8  contact_8_172
timestamp 1624494425
transform 1 0 7681 0 1 66723
box 0 0 64 64
use contact_9  contact_9_174
timestamp 1624494425
transform 1 0 7680 0 1 66323
box 0 0 66 74
use contact_8  contact_8_174
timestamp 1624494425
transform 1 0 7681 0 1 66328
box 0 0 64 64
use contact_9  contact_9_768
timestamp 1624494425
transform 1 0 8076 0 1 66718
box 0 0 66 74
use contact_8  contact_8_768
timestamp 1624494425
transform 1 0 8077 0 1 66723
box 0 0 64 64
use contact_9  contact_9_771
timestamp 1624494425
transform 1 0 8076 0 1 66323
box 0 0 66 74
use contact_8  contact_8_771
timestamp 1624494425
transform 1 0 8077 0 1 66328
box 0 0 64 64
use contact_9  contact_9_170
timestamp 1624494425
transform 1 0 7680 0 1 67113
box 0 0 66 74
use contact_8  contact_8_170
timestamp 1624494425
transform 1 0 7681 0 1 67118
box 0 0 64 64
use contact_9  contact_9_765
timestamp 1624494425
transform 1 0 8076 0 1 67113
box 0 0 66 74
use contact_8  contact_8_765
timestamp 1624494425
transform 1 0 8077 0 1 67118
box 0 0 64 64
use contact_9  contact_9_166
timestamp 1624494425
transform 1 0 7680 0 1 67903
box 0 0 66 74
use contact_8  contact_8_166
timestamp 1624494425
transform 1 0 7681 0 1 67908
box 0 0 64 64
use contact_9  contact_9_168
timestamp 1624494425
transform 1 0 7680 0 1 67508
box 0 0 66 74
use contact_8  contact_8_168
timestamp 1624494425
transform 1 0 7681 0 1 67513
box 0 0 64 64
use contact_9  contact_9_759
timestamp 1624494425
transform 1 0 8076 0 1 67903
box 0 0 66 74
use contact_8  contact_8_759
timestamp 1624494425
transform 1 0 8077 0 1 67908
box 0 0 64 64
use contact_9  contact_9_762
timestamp 1624494425
transform 1 0 8076 0 1 67508
box 0 0 66 74
use contact_8  contact_8_762
timestamp 1624494425
transform 1 0 8077 0 1 67513
box 0 0 64 64
use contact_9  contact_9_164
timestamp 1624494425
transform 1 0 7680 0 1 68298
box 0 0 66 74
use contact_8  contact_8_164
timestamp 1624494425
transform 1 0 7681 0 1 68303
box 0 0 64 64
use contact_9  contact_9_756
timestamp 1624494425
transform 1 0 8076 0 1 68298
box 0 0 66 74
use contact_8  contact_8_756
timestamp 1624494425
transform 1 0 8077 0 1 68303
box 0 0 64 64
use contact_9  contact_9_162
timestamp 1624494425
transform 1 0 7680 0 1 68693
box 0 0 66 74
use contact_8  contact_8_162
timestamp 1624494425
transform 1 0 7681 0 1 68698
box 0 0 64 64
use contact_9  contact_9_753
timestamp 1624494425
transform 1 0 8076 0 1 68693
box 0 0 66 74
use contact_8  contact_8_753
timestamp 1624494425
transform 1 0 8077 0 1 68698
box 0 0 64 64
use contact_8  contact_8_752
timestamp 1624494425
transform 1 0 7299 0 1 69116
box 0 0 64 64
use contact_9  contact_9_752
timestamp 1624494425
transform 1 0 7298 0 1 69111
box 0 0 66 74
use contact_8  contact_8_751
timestamp 1624494425
transform 1 0 6867 0 1 69116
box 0 0 64 64
use contact_9  contact_9_751
timestamp 1624494425
transform 1 0 6866 0 1 69111
box 0 0 66 74
use contact_8  contact_8_161
timestamp 1624494425
transform 1 0 6442 0 1 69116
box 0 0 64 64
use contact_9  contact_9_161
timestamp 1624494425
transform 1 0 6441 0 1 69111
box 0 0 66 74
use contact_16  contact_16_243
timestamp 1624494425
transform 1 0 5944 0 1 68984
box 0 0 66 58
use contact_16  contact_16_244
timestamp 1624494425
transform 1 0 5144 0 1 68894
box 0 0 66 58
use contact_16  contact_16_240
timestamp 1624494425
transform 1 0 5944 0 1 69208
box 0 0 66 58
use contact_16  contact_16_241
timestamp 1624494425
transform 1 0 5144 0 1 69298
box 0 0 66 58
use and3_dec  and3_dec_80
timestamp 1624494425
transform 1 0 6203 0 -1 69520
box 0 -60 2072 490
use contact_8  contact_8_749
timestamp 1624494425
transform 1 0 7299 0 1 69474
box 0 0 64 64
use contact_9  contact_9_749
timestamp 1624494425
transform 1 0 7298 0 1 69469
box 0 0 66 74
use contact_8  contact_8_748
timestamp 1624494425
transform 1 0 6867 0 1 69474
box 0 0 64 64
use contact_9  contact_9_748
timestamp 1624494425
transform 1 0 6866 0 1 69469
box 0 0 66 74
use contact_8  contact_8_159
timestamp 1624494425
transform 1 0 6442 0 1 69532
box 0 0 64 64
use contact_9  contact_9_159
timestamp 1624494425
transform 1 0 6441 0 1 69527
box 0 0 66 74
use contact_16  contact_16_239
timestamp 1624494425
transform 1 0 4584 0 1 69572
box 0 0 66 58
use contact_16  contact_16_242
timestamp 1624494425
transform 1 0 4824 0 1 69410
box 0 0 66 58
use contact_8  contact_8_746
timestamp 1624494425
transform 1 0 7299 0 1 69906
box 0 0 64 64
use contact_9  contact_9_746
timestamp 1624494425
transform 1 0 7298 0 1 69901
box 0 0 66 74
use contact_8  contact_8_745
timestamp 1624494425
transform 1 0 6867 0 1 69906
box 0 0 64 64
use contact_9  contact_9_745
timestamp 1624494425
transform 1 0 6866 0 1 69901
box 0 0 66 74
use contact_8  contact_8_157
timestamp 1624494425
transform 1 0 6442 0 1 69906
box 0 0 64 64
use contact_9  contact_9_157
timestamp 1624494425
transform 1 0 6441 0 1 69901
box 0 0 66 74
use contact_16  contact_16_237
timestamp 1624494425
transform 1 0 5944 0 1 69774
box 0 0 66 58
use contact_16  contact_16_238
timestamp 1624494425
transform 1 0 5224 0 1 69684
box 0 0 66 58
use and3_dec  and3_dec_78
timestamp 1624494425
transform 1 0 6203 0 -1 70310
box 0 -60 2072 490
use and3_dec  and3_dec_79
timestamp 1624494425
transform 1 0 6203 0 1 69520
box 0 -60 2072 490
use contact_16  contact_16_234
timestamp 1624494425
transform 1 0 5944 0 1 69998
box 0 0 66 58
use contact_16  contact_16_235
timestamp 1624494425
transform 1 0 5224 0 1 70088
box 0 0 66 58
use contact_16  contact_16_236
timestamp 1624494425
transform 1 0 4664 0 1 70200
box 0 0 66 58
use contact_8  contact_8_743
timestamp 1624494425
transform 1 0 7299 0 1 70264
box 0 0 64 64
use contact_9  contact_9_743
timestamp 1624494425
transform 1 0 7298 0 1 70259
box 0 0 66 74
use contact_8  contact_8_742
timestamp 1624494425
transform 1 0 6867 0 1 70264
box 0 0 64 64
use contact_9  contact_9_742
timestamp 1624494425
transform 1 0 6866 0 1 70259
box 0 0 66 74
use contact_8  contact_8_155
timestamp 1624494425
transform 1 0 6442 0 1 70322
box 0 0 64 64
use contact_9  contact_9_155
timestamp 1624494425
transform 1 0 6441 0 1 70317
box 0 0 66 74
use contact_16  contact_16_232
timestamp 1624494425
transform 1 0 5224 0 1 70474
box 0 0 66 58
use contact_16  contact_16_233
timestamp 1624494425
transform 1 0 4744 0 1 70362
box 0 0 66 58
use and3_dec  and3_dec_77
timestamp 1624494425
transform 1 0 6203 0 1 70310
box 0 -60 2072 490
use contact_8  contact_8_740
timestamp 1624494425
transform 1 0 7299 0 1 70696
box 0 0 64 64
use contact_9  contact_9_740
timestamp 1624494425
transform 1 0 7298 0 1 70691
box 0 0 66 74
use contact_8  contact_8_739
timestamp 1624494425
transform 1 0 6867 0 1 70696
box 0 0 64 64
use contact_9  contact_9_739
timestamp 1624494425
transform 1 0 6866 0 1 70691
box 0 0 66 74
use contact_8  contact_8_153
timestamp 1624494425
transform 1 0 6442 0 1 70696
box 0 0 64 64
use contact_9  contact_9_153
timestamp 1624494425
transform 1 0 6441 0 1 70691
box 0 0 66 74
use contact_16  contact_16_231
timestamp 1624494425
transform 1 0 5944 0 1 70564
box 0 0 66 58
use contact_16  contact_16_228
timestamp 1624494425
transform 1 0 5944 0 1 70788
box 0 0 66 58
use contact_16  contact_16_229
timestamp 1624494425
transform 1 0 5224 0 1 70878
box 0 0 66 58
use contact_16  contact_16_230
timestamp 1624494425
transform 1 0 4824 0 1 70990
box 0 0 66 58
use and3_dec  and3_dec_75
timestamp 1624494425
transform 1 0 6203 0 1 71100
box 0 -60 2072 490
use and3_dec  and3_dec_76
timestamp 1624494425
transform 1 0 6203 0 -1 71100
box 0 -60 2072 490
use contact_8  contact_8_737
timestamp 1624494425
transform 1 0 7299 0 1 71054
box 0 0 64 64
use contact_9  contact_9_737
timestamp 1624494425
transform 1 0 7298 0 1 71049
box 0 0 66 74
use contact_8  contact_8_736
timestamp 1624494425
transform 1 0 6867 0 1 71054
box 0 0 64 64
use contact_9  contact_9_736
timestamp 1624494425
transform 1 0 6866 0 1 71049
box 0 0 66 74
use contact_8  contact_8_151
timestamp 1624494425
transform 1 0 6442 0 1 71112
box 0 0 64 64
use contact_9  contact_9_151
timestamp 1624494425
transform 1 0 6441 0 1 71107
box 0 0 66 74
use contact_16  contact_16_226
timestamp 1624494425
transform 1 0 5304 0 1 71264
box 0 0 66 58
use contact_16  contact_16_227
timestamp 1624494425
transform 1 0 4584 0 1 71152
box 0 0 66 58
use contact_8  contact_8_734
timestamp 1624494425
transform 1 0 7299 0 1 71486
box 0 0 64 64
use contact_9  contact_9_734
timestamp 1624494425
transform 1 0 7298 0 1 71481
box 0 0 66 74
use contact_8  contact_8_733
timestamp 1624494425
transform 1 0 6867 0 1 71486
box 0 0 64 64
use contact_9  contact_9_733
timestamp 1624494425
transform 1 0 6866 0 1 71481
box 0 0 66 74
use contact_8  contact_8_149
timestamp 1624494425
transform 1 0 6442 0 1 71486
box 0 0 64 64
use contact_9  contact_9_149
timestamp 1624494425
transform 1 0 6441 0 1 71481
box 0 0 66 74
use contact_16  contact_16_222
timestamp 1624494425
transform 1 0 5944 0 1 71578
box 0 0 66 58
use contact_16  contact_16_225
timestamp 1624494425
transform 1 0 5944 0 1 71354
box 0 0 66 58
use and3_dec  and3_dec_74
timestamp 1624494425
transform 1 0 6203 0 -1 71890
box 0 -60 2072 490
use contact_8  contact_8_731
timestamp 1624494425
transform 1 0 7299 0 1 71844
box 0 0 64 64
use contact_9  contact_9_731
timestamp 1624494425
transform 1 0 7298 0 1 71839
box 0 0 66 74
use contact_8  contact_8_730
timestamp 1624494425
transform 1 0 6867 0 1 71844
box 0 0 64 64
use contact_9  contact_9_730
timestamp 1624494425
transform 1 0 6866 0 1 71839
box 0 0 66 74
use contact_16  contact_16_223
timestamp 1624494425
transform 1 0 5304 0 1 71668
box 0 0 66 58
use contact_16  contact_16_224
timestamp 1624494425
transform 1 0 4664 0 1 71780
box 0 0 66 58
use contact_8  contact_8_147
timestamp 1624494425
transform 1 0 6442 0 1 71902
box 0 0 64 64
use contact_9  contact_9_147
timestamp 1624494425
transform 1 0 6441 0 1 71897
box 0 0 66 74
use contact_16  contact_16_220
timestamp 1624494425
transform 1 0 5304 0 1 72054
box 0 0 66 58
use contact_16  contact_16_221
timestamp 1624494425
transform 1 0 4744 0 1 71942
box 0 0 66 58
use and3_dec  and3_dec_73
timestamp 1624494425
transform 1 0 6203 0 1 71890
box 0 -60 2072 490
use contact_9  contact_9_160
timestamp 1624494425
transform 1 0 7680 0 1 69088
box 0 0 66 74
use contact_8  contact_8_160
timestamp 1624494425
transform 1 0 7681 0 1 69093
box 0 0 64 64
use contact_9  contact_9_750
timestamp 1624494425
transform 1 0 8076 0 1 69088
box 0 0 66 74
use contact_8  contact_8_750
timestamp 1624494425
transform 1 0 8077 0 1 69093
box 0 0 64 64
use contact_9  contact_9_156
timestamp 1624494425
transform 1 0 7680 0 1 69878
box 0 0 66 74
use contact_8  contact_8_156
timestamp 1624494425
transform 1 0 7681 0 1 69883
box 0 0 64 64
use contact_9  contact_9_158
timestamp 1624494425
transform 1 0 7680 0 1 69483
box 0 0 66 74
use contact_8  contact_8_158
timestamp 1624494425
transform 1 0 7681 0 1 69488
box 0 0 64 64
use contact_9  contact_9_744
timestamp 1624494425
transform 1 0 8076 0 1 69878
box 0 0 66 74
use contact_8  contact_8_744
timestamp 1624494425
transform 1 0 8077 0 1 69883
box 0 0 64 64
use contact_9  contact_9_747
timestamp 1624494425
transform 1 0 8076 0 1 69483
box 0 0 66 74
use contact_8  contact_8_747
timestamp 1624494425
transform 1 0 8077 0 1 69488
box 0 0 64 64
use contact_9  contact_9_152
timestamp 1624494425
transform 1 0 7680 0 1 70668
box 0 0 66 74
use contact_8  contact_8_152
timestamp 1624494425
transform 1 0 7681 0 1 70673
box 0 0 64 64
use contact_9  contact_9_154
timestamp 1624494425
transform 1 0 7680 0 1 70273
box 0 0 66 74
use contact_8  contact_8_154
timestamp 1624494425
transform 1 0 7681 0 1 70278
box 0 0 64 64
use contact_9  contact_9_738
timestamp 1624494425
transform 1 0 8076 0 1 70668
box 0 0 66 74
use contact_8  contact_8_738
timestamp 1624494425
transform 1 0 8077 0 1 70673
box 0 0 64 64
use contact_9  contact_9_741
timestamp 1624494425
transform 1 0 8076 0 1 70273
box 0 0 66 74
use contact_8  contact_8_741
timestamp 1624494425
transform 1 0 8077 0 1 70278
box 0 0 64 64
use contact_9  contact_9_150
timestamp 1624494425
transform 1 0 7680 0 1 71063
box 0 0 66 74
use contact_8  contact_8_150
timestamp 1624494425
transform 1 0 7681 0 1 71068
box 0 0 64 64
use contact_9  contact_9_735
timestamp 1624494425
transform 1 0 8076 0 1 71063
box 0 0 66 74
use contact_8  contact_8_735
timestamp 1624494425
transform 1 0 8077 0 1 71068
box 0 0 64 64
use contact_9  contact_9_146
timestamp 1624494425
transform 1 0 7680 0 1 71853
box 0 0 66 74
use contact_8  contact_8_146
timestamp 1624494425
transform 1 0 7681 0 1 71858
box 0 0 64 64
use contact_9  contact_9_148
timestamp 1624494425
transform 1 0 7680 0 1 71458
box 0 0 66 74
use contact_8  contact_8_148
timestamp 1624494425
transform 1 0 7681 0 1 71463
box 0 0 64 64
use contact_9  contact_9_729
timestamp 1624494425
transform 1 0 8076 0 1 71853
box 0 0 66 74
use contact_8  contact_8_729
timestamp 1624494425
transform 1 0 8077 0 1 71858
box 0 0 64 64
use contact_9  contact_9_732
timestamp 1624494425
transform 1 0 8076 0 1 71458
box 0 0 66 74
use contact_8  contact_8_732
timestamp 1624494425
transform 1 0 8077 0 1 71463
box 0 0 64 64
use contact_8  contact_8_728
timestamp 1624494425
transform 1 0 7299 0 1 72276
box 0 0 64 64
use contact_9  contact_9_728
timestamp 1624494425
transform 1 0 7298 0 1 72271
box 0 0 66 74
use contact_8  contact_8_727
timestamp 1624494425
transform 1 0 6867 0 1 72276
box 0 0 64 64
use contact_9  contact_9_727
timestamp 1624494425
transform 1 0 6866 0 1 72271
box 0 0 66 74
use contact_8  contact_8_145
timestamp 1624494425
transform 1 0 6442 0 1 72276
box 0 0 64 64
use contact_9  contact_9_145
timestamp 1624494425
transform 1 0 6441 0 1 72271
box 0 0 66 74
use contact_16  contact_16_216
timestamp 1624494425
transform 1 0 5944 0 1 72368
box 0 0 66 58
use contact_16  contact_16_219
timestamp 1624494425
transform 1 0 5944 0 1 72144
box 0 0 66 58
use contact_8  contact_8_725
timestamp 1624494425
transform 1 0 7299 0 1 72634
box 0 0 64 64
use contact_9  contact_9_725
timestamp 1624494425
transform 1 0 7298 0 1 72629
box 0 0 66 74
use contact_8  contact_8_724
timestamp 1624494425
transform 1 0 6867 0 1 72634
box 0 0 64 64
use contact_9  contact_9_724
timestamp 1624494425
transform 1 0 6866 0 1 72629
box 0 0 66 74
use contact_16  contact_16_217
timestamp 1624494425
transform 1 0 5304 0 1 72458
box 0 0 66 58
use contact_16  contact_16_218
timestamp 1624494425
transform 1 0 4824 0 1 72570
box 0 0 66 58
use and3_dec  and3_dec_71
timestamp 1624494425
transform 1 0 6203 0 1 72680
box 0 -60 2072 490
use and3_dec  and3_dec_72
timestamp 1624494425
transform 1 0 6203 0 -1 72680
box 0 -60 2072 490
use contact_8  contact_8_143
timestamp 1624494425
transform 1 0 6442 0 1 72692
box 0 0 64 64
use contact_9  contact_9_143
timestamp 1624494425
transform 1 0 6441 0 1 72687
box 0 0 66 74
use contact_16  contact_16_213
timestamp 1624494425
transform 1 0 5944 0 1 72934
box 0 0 66 58
use contact_16  contact_16_214
timestamp 1624494425
transform 1 0 5384 0 1 72844
box 0 0 66 58
use contact_16  contact_16_215
timestamp 1624494425
transform 1 0 4584 0 1 72732
box 0 0 66 58
use contact_8  contact_8_722
timestamp 1624494425
transform 1 0 7299 0 1 73066
box 0 0 64 64
use contact_9  contact_9_722
timestamp 1624494425
transform 1 0 7298 0 1 73061
box 0 0 66 74
use contact_8  contact_8_721
timestamp 1624494425
transform 1 0 6867 0 1 73066
box 0 0 64 64
use contact_9  contact_9_721
timestamp 1624494425
transform 1 0 6866 0 1 73061
box 0 0 66 74
use contact_8  contact_8_141
timestamp 1624494425
transform 1 0 6442 0 1 73066
box 0 0 64 64
use contact_9  contact_9_141
timestamp 1624494425
transform 1 0 6441 0 1 73061
box 0 0 66 74
use contact_16  contact_16_210
timestamp 1624494425
transform 1 0 5944 0 1 73158
box 0 0 66 58
use and3_dec  and3_dec_70
timestamp 1624494425
transform 1 0 6203 0 -1 73470
box 0 -60 2072 490
use contact_8  contact_8_719
timestamp 1624494425
transform 1 0 7299 0 1 73424
box 0 0 64 64
use contact_9  contact_9_719
timestamp 1624494425
transform 1 0 7298 0 1 73419
box 0 0 66 74
use contact_8  contact_8_718
timestamp 1624494425
transform 1 0 6867 0 1 73424
box 0 0 64 64
use contact_9  contact_9_718
timestamp 1624494425
transform 1 0 6866 0 1 73419
box 0 0 66 74
use contact_8  contact_8_139
timestamp 1624494425
transform 1 0 6442 0 1 73482
box 0 0 64 64
use contact_9  contact_9_139
timestamp 1624494425
transform 1 0 6441 0 1 73477
box 0 0 66 74
use contact_16  contact_16_211
timestamp 1624494425
transform 1 0 5384 0 1 73248
box 0 0 66 58
use contact_16  contact_16_212
timestamp 1624494425
transform 1 0 4664 0 1 73360
box 0 0 66 58
use contact_16  contact_16_207
timestamp 1624494425
transform 1 0 5944 0 1 73724
box 0 0 66 58
use contact_16  contact_16_208
timestamp 1624494425
transform 1 0 5384 0 1 73634
box 0 0 66 58
use contact_16  contact_16_209
timestamp 1624494425
transform 1 0 4744 0 1 73522
box 0 0 66 58
use and3_dec  and3_dec_68
timestamp 1624494425
transform 1 0 6203 0 -1 74260
box 0 -60 2072 490
use and3_dec  and3_dec_69
timestamp 1624494425
transform 1 0 6203 0 1 73470
box 0 -60 2072 490
use contact_8  contact_8_716
timestamp 1624494425
transform 1 0 7299 0 1 73856
box 0 0 64 64
use contact_9  contact_9_716
timestamp 1624494425
transform 1 0 7298 0 1 73851
box 0 0 66 74
use contact_8  contact_8_715
timestamp 1624494425
transform 1 0 6867 0 1 73856
box 0 0 64 64
use contact_9  contact_9_715
timestamp 1624494425
transform 1 0 6866 0 1 73851
box 0 0 66 74
use contact_8  contact_8_137
timestamp 1624494425
transform 1 0 6442 0 1 73856
box 0 0 64 64
use contact_9  contact_9_137
timestamp 1624494425
transform 1 0 6441 0 1 73851
box 0 0 66 74
use contact_16  contact_16_204
timestamp 1624494425
transform 1 0 5944 0 1 73948
box 0 0 66 58
use contact_16  contact_16_205
timestamp 1624494425
transform 1 0 5384 0 1 74038
box 0 0 66 58
use contact_8  contact_8_713
timestamp 1624494425
transform 1 0 7299 0 1 74214
box 0 0 64 64
use contact_9  contact_9_713
timestamp 1624494425
transform 1 0 7298 0 1 74209
box 0 0 66 74
use contact_8  contact_8_712
timestamp 1624494425
transform 1 0 6867 0 1 74214
box 0 0 64 64
use contact_9  contact_9_712
timestamp 1624494425
transform 1 0 6866 0 1 74209
box 0 0 66 74
use contact_8  contact_8_135
timestamp 1624494425
transform 1 0 6442 0 1 74272
box 0 0 64 64
use contact_9  contact_9_135
timestamp 1624494425
transform 1 0 6441 0 1 74267
box 0 0 66 74
use contact_16  contact_16_203
timestamp 1624494425
transform 1 0 4584 0 1 74312
box 0 0 66 58
use contact_16  contact_16_206
timestamp 1624494425
transform 1 0 4824 0 1 74150
box 0 0 66 58
use and3_dec  and3_dec_67
timestamp 1624494425
transform 1 0 6203 0 1 74260
box 0 -60 2072 490
use contact_16  contact_16_201
timestamp 1624494425
transform 1 0 5944 0 1 74514
box 0 0 66 58
use contact_16  contact_16_202
timestamp 1624494425
transform 1 0 5464 0 1 74424
box 0 0 66 58
use contact_8  contact_8_710
timestamp 1624494425
transform 1 0 7299 0 1 74646
box 0 0 64 64
use contact_9  contact_9_710
timestamp 1624494425
transform 1 0 7298 0 1 74641
box 0 0 66 74
use contact_8  contact_8_709
timestamp 1624494425
transform 1 0 6867 0 1 74646
box 0 0 64 64
use contact_9  contact_9_709
timestamp 1624494425
transform 1 0 6866 0 1 74641
box 0 0 66 74
use contact_8  contact_8_133
timestamp 1624494425
transform 1 0 6442 0 1 74646
box 0 0 64 64
use contact_9  contact_9_133
timestamp 1624494425
transform 1 0 6441 0 1 74641
box 0 0 66 74
use contact_16  contact_16_198
timestamp 1624494425
transform 1 0 5944 0 1 74738
box 0 0 66 58
use contact_16  contact_16_199
timestamp 1624494425
transform 1 0 5464 0 1 74828
box 0 0 66 58
use and3_dec  and3_dec_66
timestamp 1624494425
transform 1 0 6203 0 -1 75050
box 0 -60 2072 490
use contact_8  contact_8_707
timestamp 1624494425
transform 1 0 7299 0 1 75004
box 0 0 64 64
use contact_9  contact_9_707
timestamp 1624494425
transform 1 0 7298 0 1 74999
box 0 0 66 74
use contact_8  contact_8_706
timestamp 1624494425
transform 1 0 6867 0 1 75004
box 0 0 64 64
use contact_9  contact_9_706
timestamp 1624494425
transform 1 0 6866 0 1 74999
box 0 0 66 74
use contact_8  contact_8_131
timestamp 1624494425
transform 1 0 6442 0 1 75062
box 0 0 64 64
use contact_9  contact_9_131
timestamp 1624494425
transform 1 0 6441 0 1 75057
box 0 0 66 74
use contact_16  contact_16_197
timestamp 1624494425
transform 1 0 4744 0 1 75102
box 0 0 66 58
use contact_16  contact_16_200
timestamp 1624494425
transform 1 0 4664 0 1 74940
box 0 0 66 58
use contact_16  contact_16_195
timestamp 1624494425
transform 1 0 5944 0 1 75304
box 0 0 66 58
use contact_16  contact_16_196
timestamp 1624494425
transform 1 0 5464 0 1 75214
box 0 0 66 58
use and3_dec  and3_dec_64
timestamp 1624494425
transform 1 0 6203 0 -1 75840
box 0 -60 2072 490
use and3_dec  and3_dec_65
timestamp 1624494425
transform 1 0 6203 0 1 75050
box 0 -60 2072 490
use contact_9  contact_9_142
timestamp 1624494425
transform 1 0 7680 0 1 72643
box 0 0 66 74
use contact_8  contact_8_142
timestamp 1624494425
transform 1 0 7681 0 1 72648
box 0 0 64 64
use contact_9  contact_9_144
timestamp 1624494425
transform 1 0 7680 0 1 72248
box 0 0 66 74
use contact_8  contact_8_144
timestamp 1624494425
transform 1 0 7681 0 1 72253
box 0 0 64 64
use contact_9  contact_9_723
timestamp 1624494425
transform 1 0 8076 0 1 72643
box 0 0 66 74
use contact_8  contact_8_723
timestamp 1624494425
transform 1 0 8077 0 1 72648
box 0 0 64 64
use contact_9  contact_9_726
timestamp 1624494425
transform 1 0 8076 0 1 72248
box 0 0 66 74
use contact_8  contact_8_726
timestamp 1624494425
transform 1 0 8077 0 1 72253
box 0 0 64 64
use contact_9  contact_9_140
timestamp 1624494425
transform 1 0 7680 0 1 73038
box 0 0 66 74
use contact_8  contact_8_140
timestamp 1624494425
transform 1 0 7681 0 1 73043
box 0 0 64 64
use contact_9  contact_9_720
timestamp 1624494425
transform 1 0 8076 0 1 73038
box 0 0 66 74
use contact_8  contact_8_720
timestamp 1624494425
transform 1 0 8077 0 1 73043
box 0 0 64 64
use contact_9  contact_9_136
timestamp 1624494425
transform 1 0 7680 0 1 73828
box 0 0 66 74
use contact_8  contact_8_136
timestamp 1624494425
transform 1 0 7681 0 1 73833
box 0 0 64 64
use contact_9  contact_9_138
timestamp 1624494425
transform 1 0 7680 0 1 73433
box 0 0 66 74
use contact_8  contact_8_138
timestamp 1624494425
transform 1 0 7681 0 1 73438
box 0 0 64 64
use contact_9  contact_9_714
timestamp 1624494425
transform 1 0 8076 0 1 73828
box 0 0 66 74
use contact_8  contact_8_714
timestamp 1624494425
transform 1 0 8077 0 1 73833
box 0 0 64 64
use contact_9  contact_9_717
timestamp 1624494425
transform 1 0 8076 0 1 73433
box 0 0 66 74
use contact_8  contact_8_717
timestamp 1624494425
transform 1 0 8077 0 1 73438
box 0 0 64 64
use contact_9  contact_9_134
timestamp 1624494425
transform 1 0 7680 0 1 74223
box 0 0 66 74
use contact_8  contact_8_134
timestamp 1624494425
transform 1 0 7681 0 1 74228
box 0 0 64 64
use contact_9  contact_9_711
timestamp 1624494425
transform 1 0 8076 0 1 74223
box 0 0 66 74
use contact_8  contact_8_711
timestamp 1624494425
transform 1 0 8077 0 1 74228
box 0 0 64 64
use contact_9  contact_9_130
timestamp 1624494425
transform 1 0 7680 0 1 75013
box 0 0 66 74
use contact_8  contact_8_130
timestamp 1624494425
transform 1 0 7681 0 1 75018
box 0 0 64 64
use contact_9  contact_9_132
timestamp 1624494425
transform 1 0 7680 0 1 74618
box 0 0 66 74
use contact_8  contact_8_132
timestamp 1624494425
transform 1 0 7681 0 1 74623
box 0 0 64 64
use contact_9  contact_9_705
timestamp 1624494425
transform 1 0 8076 0 1 75013
box 0 0 66 74
use contact_8  contact_8_705
timestamp 1624494425
transform 1 0 8077 0 1 75018
box 0 0 64 64
use contact_9  contact_9_708
timestamp 1624494425
transform 1 0 8076 0 1 74618
box 0 0 66 74
use contact_8  contact_8_708
timestamp 1624494425
transform 1 0 8077 0 1 74623
box 0 0 64 64
use contact_8  contact_8_704
timestamp 1624494425
transform 1 0 7299 0 1 75436
box 0 0 64 64
use contact_9  contact_9_704
timestamp 1624494425
transform 1 0 7298 0 1 75431
box 0 0 66 74
use contact_8  contact_8_703
timestamp 1624494425
transform 1 0 6867 0 1 75436
box 0 0 64 64
use contact_9  contact_9_703
timestamp 1624494425
transform 1 0 6866 0 1 75431
box 0 0 66 74
use contact_8  contact_8_129
timestamp 1624494425
transform 1 0 6442 0 1 75436
box 0 0 64 64
use contact_9  contact_9_129
timestamp 1624494425
transform 1 0 6441 0 1 75431
box 0 0 66 74
use contact_16  contact_16_192
timestamp 1624494425
transform 1 0 5944 0 1 75528
box 0 0 66 58
use contact_16  contact_16_193
timestamp 1624494425
transform 1 0 5464 0 1 75618
box 0 0 66 58
use contact_8  contact_8_701
timestamp 1624494425
transform 1 0 7299 0 1 75794
box 0 0 64 64
use contact_9  contact_9_701
timestamp 1624494425
transform 1 0 7298 0 1 75789
box 0 0 66 74
use contact_8  contact_8_700
timestamp 1624494425
transform 1 0 6867 0 1 75794
box 0 0 64 64
use contact_9  contact_9_700
timestamp 1624494425
transform 1 0 6866 0 1 75789
box 0 0 66 74
use contact_8  contact_8_127
timestamp 1624494425
transform 1 0 6442 0 1 75852
box 0 0 64 64
use contact_9  contact_9_127
timestamp 1624494425
transform 1 0 6441 0 1 75847
box 0 0 66 74
use contact_16  contact_16_191
timestamp 1624494425
transform 1 0 4584 0 1 75892
box 0 0 66 58
use contact_16  contact_16_194
timestamp 1624494425
transform 1 0 4824 0 1 75730
box 0 0 66 58
use and3_dec  and3_dec_63
timestamp 1624494425
transform 1 0 6203 0 1 75840
box 0 -60 2072 490
use contact_8  contact_8_698
timestamp 1624494425
transform 1 0 7299 0 1 76226
box 0 0 64 64
use contact_9  contact_9_698
timestamp 1624494425
transform 1 0 7298 0 1 76221
box 0 0 66 74
use contact_8  contact_8_697
timestamp 1624494425
transform 1 0 6867 0 1 76226
box 0 0 64 64
use contact_9  contact_9_697
timestamp 1624494425
transform 1 0 6866 0 1 76221
box 0 0 66 74
use contact_8  contact_8_125
timestamp 1624494425
transform 1 0 6442 0 1 76226
box 0 0 64 64
use contact_9  contact_9_125
timestamp 1624494425
transform 1 0 6441 0 1 76221
box 0 0 66 74
use contact_16  contact_16_189
timestamp 1624494425
transform 1 0 6024 0 1 76094
box 0 0 66 58
use contact_16  contact_16_190
timestamp 1624494425
transform 1 0 4904 0 1 76004
box 0 0 66 58
use contact_16  contact_16_186
timestamp 1624494425
transform 1 0 6024 0 1 76318
box 0 0 66 58
use contact_16  contact_16_187
timestamp 1624494425
transform 1 0 4904 0 1 76408
box 0 0 66 58
use and3_dec  and3_dec_62
timestamp 1624494425
transform 1 0 6203 0 -1 76630
box 0 -60 2072 490
use contact_8  contact_8_695
timestamp 1624494425
transform 1 0 7299 0 1 76584
box 0 0 64 64
use contact_9  contact_9_695
timestamp 1624494425
transform 1 0 7298 0 1 76579
box 0 0 66 74
use contact_8  contact_8_694
timestamp 1624494425
transform 1 0 6867 0 1 76584
box 0 0 64 64
use contact_9  contact_9_694
timestamp 1624494425
transform 1 0 6866 0 1 76579
box 0 0 66 74
use contact_8  contact_8_123
timestamp 1624494425
transform 1 0 6442 0 1 76642
box 0 0 64 64
use contact_9  contact_9_123
timestamp 1624494425
transform 1 0 6441 0 1 76637
box 0 0 66 74
use contact_16  contact_16_185
timestamp 1624494425
transform 1 0 4744 0 1 76682
box 0 0 66 58
use contact_16  contact_16_188
timestamp 1624494425
transform 1 0 4664 0 1 76520
box 0 0 66 58
use contact_8  contact_8_692
timestamp 1624494425
transform 1 0 7299 0 1 77016
box 0 0 64 64
use contact_9  contact_9_692
timestamp 1624494425
transform 1 0 7298 0 1 77011
box 0 0 66 74
use contact_8  contact_8_691
timestamp 1624494425
transform 1 0 6867 0 1 77016
box 0 0 64 64
use contact_9  contact_9_691
timestamp 1624494425
transform 1 0 6866 0 1 77011
box 0 0 66 74
use contact_8  contact_8_121
timestamp 1624494425
transform 1 0 6442 0 1 77016
box 0 0 64 64
use contact_9  contact_9_121
timestamp 1624494425
transform 1 0 6441 0 1 77011
box 0 0 66 74
use contact_16  contact_16_183
timestamp 1624494425
transform 1 0 6024 0 1 76884
box 0 0 66 58
use contact_16  contact_16_184
timestamp 1624494425
transform 1 0 4904 0 1 76794
box 0 0 66 58
use and3_dec  and3_dec_60
timestamp 1624494425
transform 1 0 6203 0 -1 77420
box 0 -60 2072 490
use and3_dec  and3_dec_61
timestamp 1624494425
transform 1 0 6203 0 1 76630
box 0 -60 2072 490
use contact_16  contact_16_180
timestamp 1624494425
transform 1 0 6024 0 1 77108
box 0 0 66 58
use contact_16  contact_16_181
timestamp 1624494425
transform 1 0 4904 0 1 77198
box 0 0 66 58
use contact_16  contact_16_182
timestamp 1624494425
transform 1 0 4824 0 1 77310
box 0 0 66 58
use contact_8  contact_8_689
timestamp 1624494425
transform 1 0 7299 0 1 77374
box 0 0 64 64
use contact_9  contact_9_689
timestamp 1624494425
transform 1 0 7298 0 1 77369
box 0 0 66 74
use contact_8  contact_8_688
timestamp 1624494425
transform 1 0 6867 0 1 77374
box 0 0 64 64
use contact_9  contact_9_688
timestamp 1624494425
transform 1 0 6866 0 1 77369
box 0 0 66 74
use contact_8  contact_8_119
timestamp 1624494425
transform 1 0 6442 0 1 77432
box 0 0 64 64
use contact_9  contact_9_119
timestamp 1624494425
transform 1 0 6441 0 1 77427
box 0 0 66 74
use contact_16  contact_16_178
timestamp 1624494425
transform 1 0 4984 0 1 77584
box 0 0 66 58
use contact_16  contact_16_179
timestamp 1624494425
transform 1 0 4584 0 1 77472
box 0 0 66 58
use and3_dec  and3_dec_59
timestamp 1624494425
transform 1 0 6203 0 1 77420
box 0 -60 2072 490
use contact_8  contact_8_686
timestamp 1624494425
transform 1 0 7299 0 1 77806
box 0 0 64 64
use contact_9  contact_9_686
timestamp 1624494425
transform 1 0 7298 0 1 77801
box 0 0 66 74
use contact_8  contact_8_685
timestamp 1624494425
transform 1 0 6867 0 1 77806
box 0 0 64 64
use contact_9  contact_9_685
timestamp 1624494425
transform 1 0 6866 0 1 77801
box 0 0 66 74
use contact_8  contact_8_117
timestamp 1624494425
transform 1 0 6442 0 1 77806
box 0 0 64 64
use contact_9  contact_9_117
timestamp 1624494425
transform 1 0 6441 0 1 77801
box 0 0 66 74
use contact_16  contact_16_177
timestamp 1624494425
transform 1 0 6024 0 1 77674
box 0 0 66 58
use contact_16  contact_16_174
timestamp 1624494425
transform 1 0 6024 0 1 77898
box 0 0 66 58
use contact_16  contact_16_175
timestamp 1624494425
transform 1 0 4984 0 1 77988
box 0 0 66 58
use contact_16  contact_16_176
timestamp 1624494425
transform 1 0 4664 0 1 78100
box 0 0 66 58
use and3_dec  and3_dec_57
timestamp 1624494425
transform 1 0 6203 0 1 78210
box 0 -60 2072 490
use and3_dec  and3_dec_58
timestamp 1624494425
transform 1 0 6203 0 -1 78210
box 0 -60 2072 490
use contact_8  contact_8_683
timestamp 1624494425
transform 1 0 7299 0 1 78164
box 0 0 64 64
use contact_9  contact_9_683
timestamp 1624494425
transform 1 0 7298 0 1 78159
box 0 0 66 74
use contact_8  contact_8_682
timestamp 1624494425
transform 1 0 6867 0 1 78164
box 0 0 64 64
use contact_9  contact_9_682
timestamp 1624494425
transform 1 0 6866 0 1 78159
box 0 0 66 74
use contact_8  contact_8_115
timestamp 1624494425
transform 1 0 6442 0 1 78222
box 0 0 64 64
use contact_9  contact_9_115
timestamp 1624494425
transform 1 0 6441 0 1 78217
box 0 0 66 74
use contact_16  contact_16_172
timestamp 1624494425
transform 1 0 4984 0 1 78374
box 0 0 66 58
use contact_16  contact_16_173
timestamp 1624494425
transform 1 0 4744 0 1 78262
box 0 0 66 58
use contact_8  contact_8_680
timestamp 1624494425
transform 1 0 7299 0 1 78596
box 0 0 64 64
use contact_9  contact_9_680
timestamp 1624494425
transform 1 0 7298 0 1 78591
box 0 0 66 74
use contact_8  contact_8_679
timestamp 1624494425
transform 1 0 6867 0 1 78596
box 0 0 64 64
use contact_9  contact_9_679
timestamp 1624494425
transform 1 0 6866 0 1 78591
box 0 0 66 74
use contact_8  contact_8_113
timestamp 1624494425
transform 1 0 6442 0 1 78596
box 0 0 64 64
use contact_9  contact_9_113
timestamp 1624494425
transform 1 0 6441 0 1 78591
box 0 0 66 74
use contact_16  contact_16_171
timestamp 1624494425
transform 1 0 6024 0 1 78464
box 0 0 66 58
use and3_dec  and3_dec_56
timestamp 1624494425
transform 1 0 6203 0 -1 79000
box 0 -60 2072 490
use contact_9  contact_9_126
timestamp 1624494425
transform 1 0 7680 0 1 75803
box 0 0 66 74
use contact_8  contact_8_126
timestamp 1624494425
transform 1 0 7681 0 1 75808
box 0 0 64 64
use contact_9  contact_9_128
timestamp 1624494425
transform 1 0 7680 0 1 75408
box 0 0 66 74
use contact_8  contact_8_128
timestamp 1624494425
transform 1 0 7681 0 1 75413
box 0 0 64 64
use contact_9  contact_9_699
timestamp 1624494425
transform 1 0 8076 0 1 75803
box 0 0 66 74
use contact_8  contact_8_699
timestamp 1624494425
transform 1 0 8077 0 1 75808
box 0 0 64 64
use contact_9  contact_9_702
timestamp 1624494425
transform 1 0 8076 0 1 75408
box 0 0 66 74
use contact_8  contact_8_702
timestamp 1624494425
transform 1 0 8077 0 1 75413
box 0 0 64 64
use contact_9  contact_9_124
timestamp 1624494425
transform 1 0 7680 0 1 76198
box 0 0 66 74
use contact_8  contact_8_124
timestamp 1624494425
transform 1 0 7681 0 1 76203
box 0 0 64 64
use contact_9  contact_9_696
timestamp 1624494425
transform 1 0 8076 0 1 76198
box 0 0 66 74
use contact_8  contact_8_696
timestamp 1624494425
transform 1 0 8077 0 1 76203
box 0 0 64 64
use contact_9  contact_9_120
timestamp 1624494425
transform 1 0 7680 0 1 76988
box 0 0 66 74
use contact_8  contact_8_120
timestamp 1624494425
transform 1 0 7681 0 1 76993
box 0 0 64 64
use contact_9  contact_9_122
timestamp 1624494425
transform 1 0 7680 0 1 76593
box 0 0 66 74
use contact_8  contact_8_122
timestamp 1624494425
transform 1 0 7681 0 1 76598
box 0 0 64 64
use contact_9  contact_9_690
timestamp 1624494425
transform 1 0 8076 0 1 76988
box 0 0 66 74
use contact_8  contact_8_690
timestamp 1624494425
transform 1 0 8077 0 1 76993
box 0 0 64 64
use contact_9  contact_9_693
timestamp 1624494425
transform 1 0 8076 0 1 76593
box 0 0 66 74
use contact_8  contact_8_693
timestamp 1624494425
transform 1 0 8077 0 1 76598
box 0 0 64 64
use contact_9  contact_9_118
timestamp 1624494425
transform 1 0 7680 0 1 77383
box 0 0 66 74
use contact_8  contact_8_118
timestamp 1624494425
transform 1 0 7681 0 1 77388
box 0 0 64 64
use contact_9  contact_9_687
timestamp 1624494425
transform 1 0 8076 0 1 77383
box 0 0 66 74
use contact_8  contact_8_687
timestamp 1624494425
transform 1 0 8077 0 1 77388
box 0 0 64 64
use contact_9  contact_9_114
timestamp 1624494425
transform 1 0 7680 0 1 78173
box 0 0 66 74
use contact_8  contact_8_114
timestamp 1624494425
transform 1 0 7681 0 1 78178
box 0 0 64 64
use contact_9  contact_9_116
timestamp 1624494425
transform 1 0 7680 0 1 77778
box 0 0 66 74
use contact_8  contact_8_116
timestamp 1624494425
transform 1 0 7681 0 1 77783
box 0 0 64 64
use contact_9  contact_9_681
timestamp 1624494425
transform 1 0 8076 0 1 78173
box 0 0 66 74
use contact_8  contact_8_681
timestamp 1624494425
transform 1 0 8077 0 1 78178
box 0 0 64 64
use contact_9  contact_9_684
timestamp 1624494425
transform 1 0 8076 0 1 77778
box 0 0 66 74
use contact_8  contact_8_684
timestamp 1624494425
transform 1 0 8077 0 1 77783
box 0 0 64 64
use contact_9  contact_9_112
timestamp 1624494425
transform 1 0 7680 0 1 78568
box 0 0 66 74
use contact_8  contact_8_112
timestamp 1624494425
transform 1 0 7681 0 1 78573
box 0 0 64 64
use contact_9  contact_9_678
timestamp 1624494425
transform 1 0 8076 0 1 78568
box 0 0 66 74
use contact_8  contact_8_678
timestamp 1624494425
transform 1 0 8077 0 1 78573
box 0 0 64 64
use contact_8  contact_8_677
timestamp 1624494425
transform 1 0 7299 0 1 78954
box 0 0 64 64
use contact_9  contact_9_677
timestamp 1624494425
transform 1 0 7298 0 1 78949
box 0 0 66 74
use contact_8  contact_8_676
timestamp 1624494425
transform 1 0 6867 0 1 78954
box 0 0 64 64
use contact_9  contact_9_676
timestamp 1624494425
transform 1 0 6866 0 1 78949
box 0 0 66 74
use contact_16  contact_16_168
timestamp 1624494425
transform 1 0 6024 0 1 78688
box 0 0 66 58
use contact_16  contact_16_169
timestamp 1624494425
transform 1 0 4984 0 1 78778
box 0 0 66 58
use contact_16  contact_16_170
timestamp 1624494425
transform 1 0 4824 0 1 78890
box 0 0 66 58
use contact_8  contact_8_111
timestamp 1624494425
transform 1 0 6442 0 1 79012
box 0 0 64 64
use contact_9  contact_9_111
timestamp 1624494425
transform 1 0 6441 0 1 79007
box 0 0 66 74
use contact_16  contact_16_166
timestamp 1624494425
transform 1 0 5064 0 1 79164
box 0 0 66 58
use contact_16  contact_16_167
timestamp 1624494425
transform 1 0 4584 0 1 79052
box 0 0 66 58
use and3_dec  and3_dec_55
timestamp 1624494425
transform 1 0 6203 0 1 79000
box 0 -60 2072 490
use contact_8  contact_8_674
timestamp 1624494425
transform 1 0 7299 0 1 79386
box 0 0 64 64
use contact_9  contact_9_674
timestamp 1624494425
transform 1 0 7298 0 1 79381
box 0 0 66 74
use contact_8  contact_8_673
timestamp 1624494425
transform 1 0 6867 0 1 79386
box 0 0 64 64
use contact_9  contact_9_673
timestamp 1624494425
transform 1 0 6866 0 1 79381
box 0 0 66 74
use contact_8  contact_8_109
timestamp 1624494425
transform 1 0 6442 0 1 79386
box 0 0 64 64
use contact_9  contact_9_109
timestamp 1624494425
transform 1 0 6441 0 1 79381
box 0 0 66 74
use contact_16  contact_16_162
timestamp 1624494425
transform 1 0 6024 0 1 79478
box 0 0 66 58
use contact_16  contact_16_165
timestamp 1624494425
transform 1 0 6024 0 1 79254
box 0 0 66 58
use contact_8  contact_8_671
timestamp 1624494425
transform 1 0 7299 0 1 79744
box 0 0 64 64
use contact_9  contact_9_671
timestamp 1624494425
transform 1 0 7298 0 1 79739
box 0 0 66 74
use contact_8  contact_8_670
timestamp 1624494425
transform 1 0 6867 0 1 79744
box 0 0 64 64
use contact_9  contact_9_670
timestamp 1624494425
transform 1 0 6866 0 1 79739
box 0 0 66 74
use contact_16  contact_16_163
timestamp 1624494425
transform 1 0 5064 0 1 79568
box 0 0 66 58
use contact_16  contact_16_164
timestamp 1624494425
transform 1 0 4664 0 1 79680
box 0 0 66 58
use and3_dec  and3_dec_53
timestamp 1624494425
transform 1 0 6203 0 1 79790
box 0 -60 2072 490
use and3_dec  and3_dec_54
timestamp 1624494425
transform 1 0 6203 0 -1 79790
box 0 -60 2072 490
use contact_8  contact_8_107
timestamp 1624494425
transform 1 0 6442 0 1 79802
box 0 0 64 64
use contact_9  contact_9_107
timestamp 1624494425
transform 1 0 6441 0 1 79797
box 0 0 66 74
use contact_16  contact_16_159
timestamp 1624494425
transform 1 0 6024 0 1 80044
box 0 0 66 58
use contact_16  contact_16_160
timestamp 1624494425
transform 1 0 5064 0 1 79954
box 0 0 66 58
use contact_16  contact_16_161
timestamp 1624494425
transform 1 0 4744 0 1 79842
box 0 0 66 58
use contact_8  contact_8_668
timestamp 1624494425
transform 1 0 7299 0 1 80176
box 0 0 64 64
use contact_9  contact_9_668
timestamp 1624494425
transform 1 0 7298 0 1 80171
box 0 0 66 74
use contact_8  contact_8_667
timestamp 1624494425
transform 1 0 6867 0 1 80176
box 0 0 64 64
use contact_9  contact_9_667
timestamp 1624494425
transform 1 0 6866 0 1 80171
box 0 0 66 74
use contact_8  contact_8_105
timestamp 1624494425
transform 1 0 6442 0 1 80176
box 0 0 64 64
use contact_9  contact_9_105
timestamp 1624494425
transform 1 0 6441 0 1 80171
box 0 0 66 74
use contact_16  contact_16_156
timestamp 1624494425
transform 1 0 6024 0 1 80268
box 0 0 66 58
use and3_dec  and3_dec_52
timestamp 1624494425
transform 1 0 6203 0 -1 80580
box 0 -60 2072 490
use contact_8  contact_8_665
timestamp 1624494425
transform 1 0 7299 0 1 80534
box 0 0 64 64
use contact_9  contact_9_665
timestamp 1624494425
transform 1 0 7298 0 1 80529
box 0 0 66 74
use contact_8  contact_8_664
timestamp 1624494425
transform 1 0 6867 0 1 80534
box 0 0 64 64
use contact_9  contact_9_664
timestamp 1624494425
transform 1 0 6866 0 1 80529
box 0 0 66 74
use contact_8  contact_8_103
timestamp 1624494425
transform 1 0 6442 0 1 80592
box 0 0 64 64
use contact_9  contact_9_103
timestamp 1624494425
transform 1 0 6441 0 1 80587
box 0 0 66 74
use contact_16  contact_16_157
timestamp 1624494425
transform 1 0 5064 0 1 80358
box 0 0 66 58
use contact_16  contact_16_158
timestamp 1624494425
transform 1 0 4824 0 1 80470
box 0 0 66 58
use contact_16  contact_16_153
timestamp 1624494425
transform 1 0 6024 0 1 80834
box 0 0 66 58
use contact_16  contact_16_154
timestamp 1624494425
transform 1 0 5144 0 1 80744
box 0 0 66 58
use contact_16  contact_16_155
timestamp 1624494425
transform 1 0 4584 0 1 80632
box 0 0 66 58
use and3_dec  and3_dec_50
timestamp 1624494425
transform 1 0 6203 0 -1 81370
box 0 -60 2072 490
use and3_dec  and3_dec_51
timestamp 1624494425
transform 1 0 6203 0 1 80580
box 0 -60 2072 490
use contact_8  contact_8_662
timestamp 1624494425
transform 1 0 7299 0 1 80966
box 0 0 64 64
use contact_9  contact_9_662
timestamp 1624494425
transform 1 0 7298 0 1 80961
box 0 0 66 74
use contact_8  contact_8_661
timestamp 1624494425
transform 1 0 6867 0 1 80966
box 0 0 64 64
use contact_9  contact_9_661
timestamp 1624494425
transform 1 0 6866 0 1 80961
box 0 0 66 74
use contact_8  contact_8_101
timestamp 1624494425
transform 1 0 6442 0 1 80966
box 0 0 64 64
use contact_9  contact_9_101
timestamp 1624494425
transform 1 0 6441 0 1 80961
box 0 0 66 74
use contact_16  contact_16_150
timestamp 1624494425
transform 1 0 6024 0 1 81058
box 0 0 66 58
use contact_16  contact_16_151
timestamp 1624494425
transform 1 0 5144 0 1 81148
box 0 0 66 58
use contact_8  contact_8_659
timestamp 1624494425
transform 1 0 7299 0 1 81324
box 0 0 64 64
use contact_9  contact_9_659
timestamp 1624494425
transform 1 0 7298 0 1 81319
box 0 0 66 74
use contact_8  contact_8_658
timestamp 1624494425
transform 1 0 6867 0 1 81324
box 0 0 64 64
use contact_9  contact_9_658
timestamp 1624494425
transform 1 0 6866 0 1 81319
box 0 0 66 74
use contact_8  contact_8_99
timestamp 1624494425
transform 1 0 6442 0 1 81382
box 0 0 64 64
use contact_9  contact_9_99
timestamp 1624494425
transform 1 0 6441 0 1 81377
box 0 0 66 74
use contact_16  contact_16_149
timestamp 1624494425
transform 1 0 4744 0 1 81422
box 0 0 66 58
use contact_16  contact_16_152
timestamp 1624494425
transform 1 0 4664 0 1 81260
box 0 0 66 58
use and3_dec  and3_dec_49
timestamp 1624494425
transform 1 0 6203 0 1 81370
box 0 -60 2072 490
use contact_16  contact_16_147
timestamp 1624494425
transform 1 0 6024 0 1 81624
box 0 0 66 58
use contact_16  contact_16_148
timestamp 1624494425
transform 1 0 5144 0 1 81534
box 0 0 66 58
use contact_8  contact_8_656
timestamp 1624494425
transform 1 0 7299 0 1 81756
box 0 0 64 64
use contact_9  contact_9_656
timestamp 1624494425
transform 1 0 7298 0 1 81751
box 0 0 66 74
use contact_8  contact_8_655
timestamp 1624494425
transform 1 0 6867 0 1 81756
box 0 0 64 64
use contact_9  contact_9_655
timestamp 1624494425
transform 1 0 6866 0 1 81751
box 0 0 66 74
use contact_8  contact_8_97
timestamp 1624494425
transform 1 0 6442 0 1 81756
box 0 0 64 64
use contact_9  contact_9_97
timestamp 1624494425
transform 1 0 6441 0 1 81751
box 0 0 66 74
use contact_16  contact_16_144
timestamp 1624494425
transform 1 0 6024 0 1 81848
box 0 0 66 58
use contact_16  contact_16_145
timestamp 1624494425
transform 1 0 5144 0 1 81938
box 0 0 66 58
use and3_dec  and3_dec_48
timestamp 1624494425
transform 1 0 6203 0 -1 82160
box 0 -60 2072 490
use contact_9  contact_9_110
timestamp 1624494425
transform 1 0 7680 0 1 78963
box 0 0 66 74
use contact_8  contact_8_110
timestamp 1624494425
transform 1 0 7681 0 1 78968
box 0 0 64 64
use contact_9  contact_9_675
timestamp 1624494425
transform 1 0 8076 0 1 78963
box 0 0 66 74
use contact_8  contact_8_675
timestamp 1624494425
transform 1 0 8077 0 1 78968
box 0 0 64 64
use contact_9  contact_9_106
timestamp 1624494425
transform 1 0 7680 0 1 79753
box 0 0 66 74
use contact_8  contact_8_106
timestamp 1624494425
transform 1 0 7681 0 1 79758
box 0 0 64 64
use contact_9  contact_9_108
timestamp 1624494425
transform 1 0 7680 0 1 79358
box 0 0 66 74
use contact_8  contact_8_108
timestamp 1624494425
transform 1 0 7681 0 1 79363
box 0 0 64 64
use contact_9  contact_9_669
timestamp 1624494425
transform 1 0 8076 0 1 79753
box 0 0 66 74
use contact_8  contact_8_669
timestamp 1624494425
transform 1 0 8077 0 1 79758
box 0 0 64 64
use contact_9  contact_9_672
timestamp 1624494425
transform 1 0 8076 0 1 79358
box 0 0 66 74
use contact_8  contact_8_672
timestamp 1624494425
transform 1 0 8077 0 1 79363
box 0 0 64 64
use contact_9  contact_9_102
timestamp 1624494425
transform 1 0 7680 0 1 80543
box 0 0 66 74
use contact_8  contact_8_102
timestamp 1624494425
transform 1 0 7681 0 1 80548
box 0 0 64 64
use contact_9  contact_9_104
timestamp 1624494425
transform 1 0 7680 0 1 80148
box 0 0 66 74
use contact_8  contact_8_104
timestamp 1624494425
transform 1 0 7681 0 1 80153
box 0 0 64 64
use contact_9  contact_9_663
timestamp 1624494425
transform 1 0 8076 0 1 80543
box 0 0 66 74
use contact_8  contact_8_663
timestamp 1624494425
transform 1 0 8077 0 1 80548
box 0 0 64 64
use contact_9  contact_9_666
timestamp 1624494425
transform 1 0 8076 0 1 80148
box 0 0 66 74
use contact_8  contact_8_666
timestamp 1624494425
transform 1 0 8077 0 1 80153
box 0 0 64 64
use contact_9  contact_9_100
timestamp 1624494425
transform 1 0 7680 0 1 80938
box 0 0 66 74
use contact_8  contact_8_100
timestamp 1624494425
transform 1 0 7681 0 1 80943
box 0 0 64 64
use contact_9  contact_9_660
timestamp 1624494425
transform 1 0 8076 0 1 80938
box 0 0 66 74
use contact_8  contact_8_660
timestamp 1624494425
transform 1 0 8077 0 1 80943
box 0 0 64 64
use contact_9  contact_9_96
timestamp 1624494425
transform 1 0 7680 0 1 81728
box 0 0 66 74
use contact_8  contact_8_96
timestamp 1624494425
transform 1 0 7681 0 1 81733
box 0 0 64 64
use contact_9  contact_9_98
timestamp 1624494425
transform 1 0 7680 0 1 81333
box 0 0 66 74
use contact_8  contact_8_98
timestamp 1624494425
transform 1 0 7681 0 1 81338
box 0 0 64 64
use contact_9  contact_9_654
timestamp 1624494425
transform 1 0 8076 0 1 81728
box 0 0 66 74
use contact_8  contact_8_654
timestamp 1624494425
transform 1 0 8077 0 1 81733
box 0 0 64 64
use contact_9  contact_9_657
timestamp 1624494425
transform 1 0 8076 0 1 81333
box 0 0 66 74
use contact_8  contact_8_657
timestamp 1624494425
transform 1 0 8077 0 1 81338
box 0 0 64 64
use contact_8  contact_8_653
timestamp 1624494425
transform 1 0 7299 0 1 82114
box 0 0 64 64
use contact_9  contact_9_653
timestamp 1624494425
transform 1 0 7298 0 1 82109
box 0 0 66 74
use contact_8  contact_8_652
timestamp 1624494425
transform 1 0 6867 0 1 82114
box 0 0 64 64
use contact_9  contact_9_652
timestamp 1624494425
transform 1 0 6866 0 1 82109
box 0 0 66 74
use contact_8  contact_8_95
timestamp 1624494425
transform 1 0 6442 0 1 82172
box 0 0 64 64
use contact_9  contact_9_95
timestamp 1624494425
transform 1 0 6441 0 1 82167
box 0 0 66 74
use contact_16  contact_16_143
timestamp 1624494425
transform 1 0 4584 0 1 82212
box 0 0 66 58
use contact_16  contact_16_146
timestamp 1624494425
transform 1 0 4824 0 1 82050
box 0 0 66 58
use contact_16  contact_16_141
timestamp 1624494425
transform 1 0 6024 0 1 82414
box 0 0 66 58
use contact_16  contact_16_142
timestamp 1624494425
transform 1 0 5224 0 1 82324
box 0 0 66 58
use and3_dec  and3_dec_46
timestamp 1624494425
transform 1 0 6203 0 -1 82950
box 0 -60 2072 490
use and3_dec  and3_dec_47
timestamp 1624494425
transform 1 0 6203 0 1 82160
box 0 -60 2072 490
use contact_8  contact_8_650
timestamp 1624494425
transform 1 0 7299 0 1 82546
box 0 0 64 64
use contact_9  contact_9_650
timestamp 1624494425
transform 1 0 7298 0 1 82541
box 0 0 66 74
use contact_8  contact_8_649
timestamp 1624494425
transform 1 0 6867 0 1 82546
box 0 0 64 64
use contact_9  contact_9_649
timestamp 1624494425
transform 1 0 6866 0 1 82541
box 0 0 66 74
use contact_8  contact_8_93
timestamp 1624494425
transform 1 0 6442 0 1 82546
box 0 0 64 64
use contact_9  contact_9_93
timestamp 1624494425
transform 1 0 6441 0 1 82541
box 0 0 66 74
use contact_16  contact_16_138
timestamp 1624494425
transform 1 0 6024 0 1 82638
box 0 0 66 58
use contact_16  contact_16_139
timestamp 1624494425
transform 1 0 5224 0 1 82728
box 0 0 66 58
use contact_8  contact_8_647
timestamp 1624494425
transform 1 0 7299 0 1 82904
box 0 0 64 64
use contact_9  contact_9_647
timestamp 1624494425
transform 1 0 7298 0 1 82899
box 0 0 66 74
use contact_8  contact_8_646
timestamp 1624494425
transform 1 0 6867 0 1 82904
box 0 0 64 64
use contact_9  contact_9_646
timestamp 1624494425
transform 1 0 6866 0 1 82899
box 0 0 66 74
use contact_8  contact_8_91
timestamp 1624494425
transform 1 0 6442 0 1 82962
box 0 0 64 64
use contact_9  contact_9_91
timestamp 1624494425
transform 1 0 6441 0 1 82957
box 0 0 66 74
use contact_16  contact_16_137
timestamp 1624494425
transform 1 0 4744 0 1 83002
box 0 0 66 58
use contact_16  contact_16_140
timestamp 1624494425
transform 1 0 4664 0 1 82840
box 0 0 66 58
use and3_dec  and3_dec_45
timestamp 1624494425
transform 1 0 6203 0 1 82950
box 0 -60 2072 490
use contact_8  contact_8_644
timestamp 1624494425
transform 1 0 7299 0 1 83336
box 0 0 64 64
use contact_9  contact_9_644
timestamp 1624494425
transform 1 0 7298 0 1 83331
box 0 0 66 74
use contact_8  contact_8_643
timestamp 1624494425
transform 1 0 6867 0 1 83336
box 0 0 64 64
use contact_9  contact_9_643
timestamp 1624494425
transform 1 0 6866 0 1 83331
box 0 0 66 74
use contact_8  contact_8_89
timestamp 1624494425
transform 1 0 6442 0 1 83336
box 0 0 64 64
use contact_9  contact_9_89
timestamp 1624494425
transform 1 0 6441 0 1 83331
box 0 0 66 74
use contact_16  contact_16_135
timestamp 1624494425
transform 1 0 6024 0 1 83204
box 0 0 66 58
use contact_16  contact_16_136
timestamp 1624494425
transform 1 0 5224 0 1 83114
box 0 0 66 58
use contact_16  contact_16_132
timestamp 1624494425
transform 1 0 6024 0 1 83428
box 0 0 66 58
use contact_16  contact_16_133
timestamp 1624494425
transform 1 0 5224 0 1 83518
box 0 0 66 58
use and3_dec  and3_dec_44
timestamp 1624494425
transform 1 0 6203 0 -1 83740
box 0 -60 2072 490
use contact_8  contact_8_641
timestamp 1624494425
transform 1 0 7299 0 1 83694
box 0 0 64 64
use contact_9  contact_9_641
timestamp 1624494425
transform 1 0 7298 0 1 83689
box 0 0 66 74
use contact_8  contact_8_640
timestamp 1624494425
transform 1 0 6867 0 1 83694
box 0 0 64 64
use contact_9  contact_9_640
timestamp 1624494425
transform 1 0 6866 0 1 83689
box 0 0 66 74
use contact_8  contact_8_87
timestamp 1624494425
transform 1 0 6442 0 1 83752
box 0 0 64 64
use contact_9  contact_9_87
timestamp 1624494425
transform 1 0 6441 0 1 83747
box 0 0 66 74
use contact_16  contact_16_131
timestamp 1624494425
transform 1 0 4584 0 1 83792
box 0 0 66 58
use contact_16  contact_16_134
timestamp 1624494425
transform 1 0 4824 0 1 83630
box 0 0 66 58
use contact_8  contact_8_638
timestamp 1624494425
transform 1 0 7299 0 1 84126
box 0 0 64 64
use contact_9  contact_9_638
timestamp 1624494425
transform 1 0 7298 0 1 84121
box 0 0 66 74
use contact_8  contact_8_637
timestamp 1624494425
transform 1 0 6867 0 1 84126
box 0 0 64 64
use contact_9  contact_9_637
timestamp 1624494425
transform 1 0 6866 0 1 84121
box 0 0 66 74
use contact_8  contact_8_85
timestamp 1624494425
transform 1 0 6442 0 1 84126
box 0 0 64 64
use contact_9  contact_9_85
timestamp 1624494425
transform 1 0 6441 0 1 84121
box 0 0 66 74
use contact_16  contact_16_129
timestamp 1624494425
transform 1 0 6024 0 1 83994
box 0 0 66 58
use contact_16  contact_16_130
timestamp 1624494425
transform 1 0 5304 0 1 83904
box 0 0 66 58
use and3_dec  and3_dec_42
timestamp 1624494425
transform 1 0 6203 0 -1 84530
box 0 -60 2072 490
use and3_dec  and3_dec_43
timestamp 1624494425
transform 1 0 6203 0 1 83740
box 0 -60 2072 490
use contact_16  contact_16_126
timestamp 1624494425
transform 1 0 6024 0 1 84218
box 0 0 66 58
use contact_16  contact_16_127
timestamp 1624494425
transform 1 0 5304 0 1 84308
box 0 0 66 58
use contact_16  contact_16_128
timestamp 1624494425
transform 1 0 4664 0 1 84420
box 0 0 66 58
use contact_8  contact_8_635
timestamp 1624494425
transform 1 0 7299 0 1 84484
box 0 0 64 64
use contact_9  contact_9_635
timestamp 1624494425
transform 1 0 7298 0 1 84479
box 0 0 66 74
use contact_8  contact_8_634
timestamp 1624494425
transform 1 0 6867 0 1 84484
box 0 0 64 64
use contact_9  contact_9_634
timestamp 1624494425
transform 1 0 6866 0 1 84479
box 0 0 66 74
use contact_8  contact_8_83
timestamp 1624494425
transform 1 0 6442 0 1 84542
box 0 0 64 64
use contact_9  contact_9_83
timestamp 1624494425
transform 1 0 6441 0 1 84537
box 0 0 66 74
use contact_16  contact_16_124
timestamp 1624494425
transform 1 0 5304 0 1 84694
box 0 0 66 58
use contact_16  contact_16_125
timestamp 1624494425
transform 1 0 4744 0 1 84582
box 0 0 66 58
use and3_dec  and3_dec_41
timestamp 1624494425
transform 1 0 6203 0 1 84530
box 0 -60 2072 490
use contact_8  contact_8_632
timestamp 1624494425
transform 1 0 7299 0 1 84916
box 0 0 64 64
use contact_9  contact_9_632
timestamp 1624494425
transform 1 0 7298 0 1 84911
box 0 0 66 74
use contact_8  contact_8_631
timestamp 1624494425
transform 1 0 6867 0 1 84916
box 0 0 64 64
use contact_9  contact_9_631
timestamp 1624494425
transform 1 0 6866 0 1 84911
box 0 0 66 74
use contact_8  contact_8_81
timestamp 1624494425
transform 1 0 6442 0 1 84916
box 0 0 64 64
use contact_9  contact_9_81
timestamp 1624494425
transform 1 0 6441 0 1 84911
box 0 0 66 74
use contact_16  contact_16_123
timestamp 1624494425
transform 1 0 6024 0 1 84784
box 0 0 66 58
use contact_16  contact_16_120
timestamp 1624494425
transform 1 0 6024 0 1 85008
box 0 0 66 58
use contact_16  contact_16_121
timestamp 1624494425
transform 1 0 5304 0 1 85098
box 0 0 66 58
use contact_16  contact_16_122
timestamp 1624494425
transform 1 0 4824 0 1 85210
box 0 0 66 58
use and3_dec  and3_dec_40
timestamp 1624494425
transform 1 0 6203 0 -1 85320
box 0 -60 2072 490
use contact_9  contact_9_92
timestamp 1624494425
transform 1 0 7680 0 1 82518
box 0 0 66 74
use contact_8  contact_8_92
timestamp 1624494425
transform 1 0 7681 0 1 82523
box 0 0 64 64
use contact_9  contact_9_94
timestamp 1624494425
transform 1 0 7680 0 1 82123
box 0 0 66 74
use contact_8  contact_8_94
timestamp 1624494425
transform 1 0 7681 0 1 82128
box 0 0 64 64
use contact_9  contact_9_648
timestamp 1624494425
transform 1 0 8076 0 1 82518
box 0 0 66 74
use contact_8  contact_8_648
timestamp 1624494425
transform 1 0 8077 0 1 82523
box 0 0 64 64
use contact_9  contact_9_651
timestamp 1624494425
transform 1 0 8076 0 1 82123
box 0 0 66 74
use contact_8  contact_8_651
timestamp 1624494425
transform 1 0 8077 0 1 82128
box 0 0 64 64
use contact_9  contact_9_90
timestamp 1624494425
transform 1 0 7680 0 1 82913
box 0 0 66 74
use contact_8  contact_8_90
timestamp 1624494425
transform 1 0 7681 0 1 82918
box 0 0 64 64
use contact_9  contact_9_645
timestamp 1624494425
transform 1 0 8076 0 1 82913
box 0 0 66 74
use contact_8  contact_8_645
timestamp 1624494425
transform 1 0 8077 0 1 82918
box 0 0 64 64
use contact_9  contact_9_86
timestamp 1624494425
transform 1 0 7680 0 1 83703
box 0 0 66 74
use contact_8  contact_8_86
timestamp 1624494425
transform 1 0 7681 0 1 83708
box 0 0 64 64
use contact_9  contact_9_88
timestamp 1624494425
transform 1 0 7680 0 1 83308
box 0 0 66 74
use contact_8  contact_8_88
timestamp 1624494425
transform 1 0 7681 0 1 83313
box 0 0 64 64
use contact_9  contact_9_639
timestamp 1624494425
transform 1 0 8076 0 1 83703
box 0 0 66 74
use contact_8  contact_8_639
timestamp 1624494425
transform 1 0 8077 0 1 83708
box 0 0 64 64
use contact_9  contact_9_642
timestamp 1624494425
transform 1 0 8076 0 1 83308
box 0 0 66 74
use contact_8  contact_8_642
timestamp 1624494425
transform 1 0 8077 0 1 83313
box 0 0 64 64
use contact_9  contact_9_84
timestamp 1624494425
transform 1 0 7680 0 1 84098
box 0 0 66 74
use contact_8  contact_8_84
timestamp 1624494425
transform 1 0 7681 0 1 84103
box 0 0 64 64
use contact_9  contact_9_636
timestamp 1624494425
transform 1 0 8076 0 1 84098
box 0 0 66 74
use contact_8  contact_8_636
timestamp 1624494425
transform 1 0 8077 0 1 84103
box 0 0 64 64
use contact_9  contact_9_80
timestamp 1624494425
transform 1 0 7680 0 1 84888
box 0 0 66 74
use contact_8  contact_8_80
timestamp 1624494425
transform 1 0 7681 0 1 84893
box 0 0 64 64
use contact_9  contact_9_82
timestamp 1624494425
transform 1 0 7680 0 1 84493
box 0 0 66 74
use contact_8  contact_8_82
timestamp 1624494425
transform 1 0 7681 0 1 84498
box 0 0 64 64
use contact_9  contact_9_630
timestamp 1624494425
transform 1 0 8076 0 1 84888
box 0 0 66 74
use contact_8  contact_8_630
timestamp 1624494425
transform 1 0 8077 0 1 84893
box 0 0 64 64
use contact_9  contact_9_633
timestamp 1624494425
transform 1 0 8076 0 1 84493
box 0 0 66 74
use contact_8  contact_8_633
timestamp 1624494425
transform 1 0 8077 0 1 84498
box 0 0 64 64
use contact_8  contact_8_629
timestamp 1624494425
transform 1 0 7299 0 1 85274
box 0 0 64 64
use contact_9  contact_9_629
timestamp 1624494425
transform 1 0 7298 0 1 85269
box 0 0 66 74
use contact_8  contact_8_628
timestamp 1624494425
transform 1 0 6867 0 1 85274
box 0 0 64 64
use contact_9  contact_9_628
timestamp 1624494425
transform 1 0 6866 0 1 85269
box 0 0 66 74
use contact_8  contact_8_79
timestamp 1624494425
transform 1 0 6442 0 1 85332
box 0 0 64 64
use contact_9  contact_9_79
timestamp 1624494425
transform 1 0 6441 0 1 85327
box 0 0 66 74
use contact_16  contact_16_118
timestamp 1624494425
transform 1 0 5384 0 1 85484
box 0 0 66 58
use contact_16  contact_16_119
timestamp 1624494425
transform 1 0 4584 0 1 85372
box 0 0 66 58
use contact_8  contact_8_626
timestamp 1624494425
transform 1 0 7299 0 1 85706
box 0 0 64 64
use contact_9  contact_9_626
timestamp 1624494425
transform 1 0 7298 0 1 85701
box 0 0 66 74
use contact_8  contact_8_625
timestamp 1624494425
transform 1 0 6867 0 1 85706
box 0 0 64 64
use contact_9  contact_9_625
timestamp 1624494425
transform 1 0 6866 0 1 85701
box 0 0 66 74
use contact_8  contact_8_77
timestamp 1624494425
transform 1 0 6442 0 1 85706
box 0 0 64 64
use contact_9  contact_9_77
timestamp 1624494425
transform 1 0 6441 0 1 85701
box 0 0 66 74
use contact_16  contact_16_117
timestamp 1624494425
transform 1 0 6024 0 1 85574
box 0 0 66 58
use and3_dec  and3_dec_38
timestamp 1624494425
transform 1 0 6203 0 -1 86110
box 0 -60 2072 490
use and3_dec  and3_dec_39
timestamp 1624494425
transform 1 0 6203 0 1 85320
box 0 -60 2072 490
use contact_8  contact_8_623
timestamp 1624494425
transform 1 0 7299 0 1 86064
box 0 0 64 64
use contact_9  contact_9_623
timestamp 1624494425
transform 1 0 7298 0 1 86059
box 0 0 66 74
use contact_8  contact_8_622
timestamp 1624494425
transform 1 0 6867 0 1 86064
box 0 0 64 64
use contact_9  contact_9_622
timestamp 1624494425
transform 1 0 6866 0 1 86059
box 0 0 66 74
use contact_16  contact_16_114
timestamp 1624494425
transform 1 0 6024 0 1 85798
box 0 0 66 58
use contact_16  contact_16_115
timestamp 1624494425
transform 1 0 5384 0 1 85888
box 0 0 66 58
use contact_16  contact_16_116
timestamp 1624494425
transform 1 0 4664 0 1 86000
box 0 0 66 58
use contact_8  contact_8_75
timestamp 1624494425
transform 1 0 6442 0 1 86122
box 0 0 64 64
use contact_9  contact_9_75
timestamp 1624494425
transform 1 0 6441 0 1 86117
box 0 0 66 74
use contact_16  contact_16_112
timestamp 1624494425
transform 1 0 5384 0 1 86274
box 0 0 66 58
use contact_16  contact_16_113
timestamp 1624494425
transform 1 0 4744 0 1 86162
box 0 0 66 58
use and3_dec  and3_dec_37
timestamp 1624494425
transform 1 0 6203 0 1 86110
box 0 -60 2072 490
use contact_8  contact_8_620
timestamp 1624494425
transform 1 0 7299 0 1 86496
box 0 0 64 64
use contact_9  contact_9_620
timestamp 1624494425
transform 1 0 7298 0 1 86491
box 0 0 66 74
use contact_8  contact_8_619
timestamp 1624494425
transform 1 0 6867 0 1 86496
box 0 0 64 64
use contact_9  contact_9_619
timestamp 1624494425
transform 1 0 6866 0 1 86491
box 0 0 66 74
use contact_8  contact_8_73
timestamp 1624494425
transform 1 0 6442 0 1 86496
box 0 0 64 64
use contact_9  contact_9_73
timestamp 1624494425
transform 1 0 6441 0 1 86491
box 0 0 66 74
use contact_16  contact_16_108
timestamp 1624494425
transform 1 0 6024 0 1 86588
box 0 0 66 58
use contact_16  contact_16_111
timestamp 1624494425
transform 1 0 6024 0 1 86364
box 0 0 66 58
use contact_8  contact_8_617
timestamp 1624494425
transform 1 0 7299 0 1 86854
box 0 0 64 64
use contact_9  contact_9_617
timestamp 1624494425
transform 1 0 7298 0 1 86849
box 0 0 66 74
use contact_8  contact_8_616
timestamp 1624494425
transform 1 0 6867 0 1 86854
box 0 0 64 64
use contact_9  contact_9_616
timestamp 1624494425
transform 1 0 6866 0 1 86849
box 0 0 66 74
use contact_16  contact_16_109
timestamp 1624494425
transform 1 0 5384 0 1 86678
box 0 0 66 58
use contact_16  contact_16_110
timestamp 1624494425
transform 1 0 4824 0 1 86790
box 0 0 66 58
use and3_dec  and3_dec_35
timestamp 1624494425
transform 1 0 6203 0 1 86900
box 0 -60 2072 490
use and3_dec  and3_dec_36
timestamp 1624494425
transform 1 0 6203 0 -1 86900
box 0 -60 2072 490
use contact_8  contact_8_71
timestamp 1624494425
transform 1 0 6442 0 1 86912
box 0 0 64 64
use contact_9  contact_9_71
timestamp 1624494425
transform 1 0 6441 0 1 86907
box 0 0 66 74
use contact_16  contact_16_105
timestamp 1624494425
transform 1 0 6024 0 1 87154
box 0 0 66 58
use contact_16  contact_16_106
timestamp 1624494425
transform 1 0 5464 0 1 87064
box 0 0 66 58
use contact_16  contact_16_107
timestamp 1624494425
transform 1 0 4584 0 1 86952
box 0 0 66 58
use contact_8  contact_8_614
timestamp 1624494425
transform 1 0 7299 0 1 87286
box 0 0 64 64
use contact_9  contact_9_614
timestamp 1624494425
transform 1 0 7298 0 1 87281
box 0 0 66 74
use contact_8  contact_8_613
timestamp 1624494425
transform 1 0 6867 0 1 87286
box 0 0 64 64
use contact_9  contact_9_613
timestamp 1624494425
transform 1 0 6866 0 1 87281
box 0 0 66 74
use contact_8  contact_8_69
timestamp 1624494425
transform 1 0 6442 0 1 87286
box 0 0 64 64
use contact_9  contact_9_69
timestamp 1624494425
transform 1 0 6441 0 1 87281
box 0 0 66 74
use contact_16  contact_16_102
timestamp 1624494425
transform 1 0 6024 0 1 87378
box 0 0 66 58
use and3_dec  and3_dec_34
timestamp 1624494425
transform 1 0 6203 0 -1 87690
box 0 -60 2072 490
use contact_8  contact_8_611
timestamp 1624494425
transform 1 0 7299 0 1 87644
box 0 0 64 64
use contact_9  contact_9_611
timestamp 1624494425
transform 1 0 7298 0 1 87639
box 0 0 66 74
use contact_8  contact_8_610
timestamp 1624494425
transform 1 0 6867 0 1 87644
box 0 0 64 64
use contact_9  contact_9_610
timestamp 1624494425
transform 1 0 6866 0 1 87639
box 0 0 66 74
use contact_8  contact_8_67
timestamp 1624494425
transform 1 0 6442 0 1 87702
box 0 0 64 64
use contact_9  contact_9_67
timestamp 1624494425
transform 1 0 6441 0 1 87697
box 0 0 66 74
use contact_16  contact_16_103
timestamp 1624494425
transform 1 0 5464 0 1 87468
box 0 0 66 58
use contact_16  contact_16_104
timestamp 1624494425
transform 1 0 4664 0 1 87580
box 0 0 66 58
use contact_16  contact_16_99
timestamp 1624494425
transform 1 0 6024 0 1 87944
box 0 0 66 58
use contact_16  contact_16_100
timestamp 1624494425
transform 1 0 5464 0 1 87854
box 0 0 66 58
use contact_16  contact_16_101
timestamp 1624494425
transform 1 0 4744 0 1 87742
box 0 0 66 58
use and3_dec  and3_dec_32
timestamp 1624494425
transform 1 0 6203 0 -1 88480
box 0 -60 2072 490
use and3_dec  and3_dec_33
timestamp 1624494425
transform 1 0 6203 0 1 87690
box 0 -60 2072 490
use contact_8  contact_8_608
timestamp 1624494425
transform 1 0 7299 0 1 88076
box 0 0 64 64
use contact_9  contact_9_608
timestamp 1624494425
transform 1 0 7298 0 1 88071
box 0 0 66 74
use contact_8  contact_8_607
timestamp 1624494425
transform 1 0 6867 0 1 88076
box 0 0 64 64
use contact_9  contact_9_607
timestamp 1624494425
transform 1 0 6866 0 1 88071
box 0 0 66 74
use contact_8  contact_8_65
timestamp 1624494425
transform 1 0 6442 0 1 88076
box 0 0 64 64
use contact_9  contact_9_65
timestamp 1624494425
transform 1 0 6441 0 1 88071
box 0 0 66 74
use contact_16  contact_16_96
timestamp 1624494425
transform 1 0 6024 0 1 88168
box 0 0 66 58
use contact_16  contact_16_97
timestamp 1624494425
transform 1 0 5464 0 1 88258
box 0 0 66 58
use contact_8  contact_8_605
timestamp 1624494425
transform 1 0 7299 0 1 88434
box 0 0 64 64
use contact_9  contact_9_605
timestamp 1624494425
transform 1 0 7298 0 1 88429
box 0 0 66 74
use contact_8  contact_8_604
timestamp 1624494425
transform 1 0 6867 0 1 88434
box 0 0 64 64
use contact_9  contact_9_604
timestamp 1624494425
transform 1 0 6866 0 1 88429
box 0 0 66 74
use contact_8  contact_8_63
timestamp 1624494425
transform 1 0 6442 0 1 88492
box 0 0 64 64
use contact_9  contact_9_63
timestamp 1624494425
transform 1 0 6441 0 1 88487
box 0 0 66 74
use contact_16  contact_16_98
timestamp 1624494425
transform 1 0 4824 0 1 88370
box 0 0 66 58
use and3_dec  and3_dec_31
timestamp 1624494425
transform 1 0 6203 0 1 88480
box 0 -60 2072 490
use contact_9  contact_9_76
timestamp 1624494425
transform 1 0 7680 0 1 85678
box 0 0 66 74
use contact_8  contact_8_76
timestamp 1624494425
transform 1 0 7681 0 1 85683
box 0 0 64 64
use contact_9  contact_9_78
timestamp 1624494425
transform 1 0 7680 0 1 85283
box 0 0 66 74
use contact_8  contact_8_78
timestamp 1624494425
transform 1 0 7681 0 1 85288
box 0 0 64 64
use contact_9  contact_9_624
timestamp 1624494425
transform 1 0 8076 0 1 85678
box 0 0 66 74
use contact_8  contact_8_624
timestamp 1624494425
transform 1 0 8077 0 1 85683
box 0 0 64 64
use contact_9  contact_9_627
timestamp 1624494425
transform 1 0 8076 0 1 85283
box 0 0 66 74
use contact_8  contact_8_627
timestamp 1624494425
transform 1 0 8077 0 1 85288
box 0 0 64 64
use contact_9  contact_9_74
timestamp 1624494425
transform 1 0 7680 0 1 86073
box 0 0 66 74
use contact_8  contact_8_74
timestamp 1624494425
transform 1 0 7681 0 1 86078
box 0 0 64 64
use contact_9  contact_9_621
timestamp 1624494425
transform 1 0 8076 0 1 86073
box 0 0 66 74
use contact_8  contact_8_621
timestamp 1624494425
transform 1 0 8077 0 1 86078
box 0 0 64 64
use contact_9  contact_9_70
timestamp 1624494425
transform 1 0 7680 0 1 86863
box 0 0 66 74
use contact_8  contact_8_70
timestamp 1624494425
transform 1 0 7681 0 1 86868
box 0 0 64 64
use contact_9  contact_9_72
timestamp 1624494425
transform 1 0 7680 0 1 86468
box 0 0 66 74
use contact_8  contact_8_72
timestamp 1624494425
transform 1 0 7681 0 1 86473
box 0 0 64 64
use contact_9  contact_9_615
timestamp 1624494425
transform 1 0 8076 0 1 86863
box 0 0 66 74
use contact_8  contact_8_615
timestamp 1624494425
transform 1 0 8077 0 1 86868
box 0 0 64 64
use contact_9  contact_9_618
timestamp 1624494425
transform 1 0 8076 0 1 86468
box 0 0 66 74
use contact_8  contact_8_618
timestamp 1624494425
transform 1 0 8077 0 1 86473
box 0 0 64 64
use contact_9  contact_9_68
timestamp 1624494425
transform 1 0 7680 0 1 87258
box 0 0 66 74
use contact_8  contact_8_68
timestamp 1624494425
transform 1 0 7681 0 1 87263
box 0 0 64 64
use contact_9  contact_9_612
timestamp 1624494425
transform 1 0 8076 0 1 87258
box 0 0 66 74
use contact_8  contact_8_612
timestamp 1624494425
transform 1 0 8077 0 1 87263
box 0 0 64 64
use contact_9  contact_9_64
timestamp 1624494425
transform 1 0 7680 0 1 88048
box 0 0 66 74
use contact_8  contact_8_64
timestamp 1624494425
transform 1 0 7681 0 1 88053
box 0 0 64 64
use contact_9  contact_9_66
timestamp 1624494425
transform 1 0 7680 0 1 87653
box 0 0 66 74
use contact_8  contact_8_66
timestamp 1624494425
transform 1 0 7681 0 1 87658
box 0 0 64 64
use contact_9  contact_9_606
timestamp 1624494425
transform 1 0 8076 0 1 88048
box 0 0 66 74
use contact_8  contact_8_606
timestamp 1624494425
transform 1 0 8077 0 1 88053
box 0 0 64 64
use contact_9  contact_9_609
timestamp 1624494425
transform 1 0 8076 0 1 87653
box 0 0 66 74
use contact_8  contact_8_609
timestamp 1624494425
transform 1 0 8077 0 1 87658
box 0 0 64 64
use contact_9  contact_9_62
timestamp 1624494425
transform 1 0 7680 0 1 88443
box 0 0 66 74
use contact_8  contact_8_62
timestamp 1624494425
transform 1 0 7681 0 1 88448
box 0 0 64 64
use contact_9  contact_9_603
timestamp 1624494425
transform 1 0 8076 0 1 88443
box 0 0 66 74
use contact_8  contact_8_603
timestamp 1624494425
transform 1 0 8077 0 1 88448
box 0 0 64 64
use contact_16  contact_16_93
timestamp 1624494425
transform 1 0 6104 0 1 88734
box 0 0 66 58
use contact_16  contact_16_94
timestamp 1624494425
transform 1 0 4904 0 1 88644
box 0 0 66 58
use contact_16  contact_16_95
timestamp 1624494425
transform 1 0 4584 0 1 88532
box 0 0 66 58
use contact_8  contact_8_602
timestamp 1624494425
transform 1 0 7299 0 1 88866
box 0 0 64 64
use contact_9  contact_9_602
timestamp 1624494425
transform 1 0 7298 0 1 88861
box 0 0 66 74
use contact_8  contact_8_601
timestamp 1624494425
transform 1 0 6867 0 1 88866
box 0 0 64 64
use contact_9  contact_9_601
timestamp 1624494425
transform 1 0 6866 0 1 88861
box 0 0 66 74
use contact_8  contact_8_61
timestamp 1624494425
transform 1 0 6442 0 1 88866
box 0 0 64 64
use contact_9  contact_9_61
timestamp 1624494425
transform 1 0 6441 0 1 88861
box 0 0 66 74
use contact_16  contact_16_90
timestamp 1624494425
transform 1 0 6104 0 1 88958
box 0 0 66 58
use contact_16  contact_16_91
timestamp 1624494425
transform 1 0 4904 0 1 89048
box 0 0 66 58
use and3_dec  and3_dec_30
timestamp 1624494425
transform 1 0 6203 0 -1 89270
box 0 -60 2072 490
use contact_8  contact_8_599
timestamp 1624494425
transform 1 0 7299 0 1 89224
box 0 0 64 64
use contact_9  contact_9_599
timestamp 1624494425
transform 1 0 7298 0 1 89219
box 0 0 66 74
use contact_8  contact_8_598
timestamp 1624494425
transform 1 0 6867 0 1 89224
box 0 0 64 64
use contact_9  contact_9_598
timestamp 1624494425
transform 1 0 6866 0 1 89219
box 0 0 66 74
use contact_8  contact_8_59
timestamp 1624494425
transform 1 0 6442 0 1 89282
box 0 0 64 64
use contact_9  contact_9_59
timestamp 1624494425
transform 1 0 6441 0 1 89277
box 0 0 66 74
use contact_16  contact_16_89
timestamp 1624494425
transform 1 0 4744 0 1 89322
box 0 0 66 58
use contact_16  contact_16_92
timestamp 1624494425
transform 1 0 4664 0 1 89160
box 0 0 66 58
use contact_16  contact_16_87
timestamp 1624494425
transform 1 0 6104 0 1 89524
box 0 0 66 58
use contact_16  contact_16_88
timestamp 1624494425
transform 1 0 4904 0 1 89434
box 0 0 66 58
use and3_dec  and3_dec_28
timestamp 1624494425
transform 1 0 6203 0 -1 90060
box 0 -60 2072 490
use and3_dec  and3_dec_29
timestamp 1624494425
transform 1 0 6203 0 1 89270
box 0 -60 2072 490
use contact_8  contact_8_596
timestamp 1624494425
transform 1 0 7299 0 1 89656
box 0 0 64 64
use contact_9  contact_9_596
timestamp 1624494425
transform 1 0 7298 0 1 89651
box 0 0 66 74
use contact_8  contact_8_595
timestamp 1624494425
transform 1 0 6867 0 1 89656
box 0 0 64 64
use contact_9  contact_9_595
timestamp 1624494425
transform 1 0 6866 0 1 89651
box 0 0 66 74
use contact_8  contact_8_57
timestamp 1624494425
transform 1 0 6442 0 1 89656
box 0 0 64 64
use contact_9  contact_9_57
timestamp 1624494425
transform 1 0 6441 0 1 89651
box 0 0 66 74
use contact_16  contact_16_84
timestamp 1624494425
transform 1 0 6104 0 1 89748
box 0 0 66 58
use contact_16  contact_16_85
timestamp 1624494425
transform 1 0 4904 0 1 89838
box 0 0 66 58
use contact_8  contact_8_593
timestamp 1624494425
transform 1 0 7299 0 1 90014
box 0 0 64 64
use contact_9  contact_9_593
timestamp 1624494425
transform 1 0 7298 0 1 90009
box 0 0 66 74
use contact_8  contact_8_592
timestamp 1624494425
transform 1 0 6867 0 1 90014
box 0 0 64 64
use contact_9  contact_9_592
timestamp 1624494425
transform 1 0 6866 0 1 90009
box 0 0 66 74
use contact_8  contact_8_55
timestamp 1624494425
transform 1 0 6442 0 1 90072
box 0 0 64 64
use contact_9  contact_9_55
timestamp 1624494425
transform 1 0 6441 0 1 90067
box 0 0 66 74
use contact_16  contact_16_83
timestamp 1624494425
transform 1 0 4584 0 1 90112
box 0 0 66 58
use contact_16  contact_16_86
timestamp 1624494425
transform 1 0 4824 0 1 89950
box 0 0 66 58
use and3_dec  and3_dec_27
timestamp 1624494425
transform 1 0 6203 0 1 90060
box 0 -60 2072 490
use contact_8  contact_8_590
timestamp 1624494425
transform 1 0 7299 0 1 90446
box 0 0 64 64
use contact_9  contact_9_590
timestamp 1624494425
transform 1 0 7298 0 1 90441
box 0 0 66 74
use contact_8  contact_8_589
timestamp 1624494425
transform 1 0 6867 0 1 90446
box 0 0 64 64
use contact_9  contact_9_589
timestamp 1624494425
transform 1 0 6866 0 1 90441
box 0 0 66 74
use contact_8  contact_8_53
timestamp 1624494425
transform 1 0 6442 0 1 90446
box 0 0 64 64
use contact_9  contact_9_53
timestamp 1624494425
transform 1 0 6441 0 1 90441
box 0 0 66 74
use contact_16  contact_16_81
timestamp 1624494425
transform 1 0 6104 0 1 90314
box 0 0 66 58
use contact_16  contact_16_82
timestamp 1624494425
transform 1 0 4984 0 1 90224
box 0 0 66 58
use contact_16  contact_16_78
timestamp 1624494425
transform 1 0 6104 0 1 90538
box 0 0 66 58
use contact_16  contact_16_79
timestamp 1624494425
transform 1 0 4984 0 1 90628
box 0 0 66 58
use and3_dec  and3_dec_26
timestamp 1624494425
transform 1 0 6203 0 -1 90850
box 0 -60 2072 490
use contact_8  contact_8_587
timestamp 1624494425
transform 1 0 7299 0 1 90804
box 0 0 64 64
use contact_9  contact_9_587
timestamp 1624494425
transform 1 0 7298 0 1 90799
box 0 0 66 74
use contact_8  contact_8_586
timestamp 1624494425
transform 1 0 6867 0 1 90804
box 0 0 64 64
use contact_9  contact_9_586
timestamp 1624494425
transform 1 0 6866 0 1 90799
box 0 0 66 74
use contact_8  contact_8_51
timestamp 1624494425
transform 1 0 6442 0 1 90862
box 0 0 64 64
use contact_9  contact_9_51
timestamp 1624494425
transform 1 0 6441 0 1 90857
box 0 0 66 74
use contact_16  contact_16_77
timestamp 1624494425
transform 1 0 4744 0 1 90902
box 0 0 66 58
use contact_16  contact_16_80
timestamp 1624494425
transform 1 0 4664 0 1 90740
box 0 0 66 58
use contact_8  contact_8_584
timestamp 1624494425
transform 1 0 7299 0 1 91236
box 0 0 64 64
use contact_9  contact_9_584
timestamp 1624494425
transform 1 0 7298 0 1 91231
box 0 0 66 74
use contact_8  contact_8_583
timestamp 1624494425
transform 1 0 6867 0 1 91236
box 0 0 64 64
use contact_9  contact_9_583
timestamp 1624494425
transform 1 0 6866 0 1 91231
box 0 0 66 74
use contact_8  contact_8_49
timestamp 1624494425
transform 1 0 6442 0 1 91236
box 0 0 64 64
use contact_9  contact_9_49
timestamp 1624494425
transform 1 0 6441 0 1 91231
box 0 0 66 74
use contact_16  contact_16_75
timestamp 1624494425
transform 1 0 6104 0 1 91104
box 0 0 66 58
use contact_16  contact_16_76
timestamp 1624494425
transform 1 0 4984 0 1 91014
box 0 0 66 58
use and3_dec  and3_dec_24
timestamp 1624494425
transform 1 0 6203 0 -1 91640
box 0 -60 2072 490
use and3_dec  and3_dec_25
timestamp 1624494425
transform 1 0 6203 0 1 90850
box 0 -60 2072 490
use contact_16  contact_16_72
timestamp 1624494425
transform 1 0 6104 0 1 91328
box 0 0 66 58
use contact_16  contact_16_73
timestamp 1624494425
transform 1 0 4984 0 1 91418
box 0 0 66 58
use contact_16  contact_16_74
timestamp 1624494425
transform 1 0 4824 0 1 91530
box 0 0 66 58
use contact_8  contact_8_581
timestamp 1624494425
transform 1 0 7299 0 1 91594
box 0 0 64 64
use contact_9  contact_9_581
timestamp 1624494425
transform 1 0 7298 0 1 91589
box 0 0 66 74
use contact_8  contact_8_580
timestamp 1624494425
transform 1 0 6867 0 1 91594
box 0 0 64 64
use contact_9  contact_9_580
timestamp 1624494425
transform 1 0 6866 0 1 91589
box 0 0 66 74
use contact_8  contact_8_47
timestamp 1624494425
transform 1 0 6442 0 1 91652
box 0 0 64 64
use contact_9  contact_9_47
timestamp 1624494425
transform 1 0 6441 0 1 91647
box 0 0 66 74
use contact_16  contact_16_70
timestamp 1624494425
transform 1 0 5064 0 1 91804
box 0 0 66 58
use contact_16  contact_16_71
timestamp 1624494425
transform 1 0 4584 0 1 91692
box 0 0 66 58
use and3_dec  and3_dec_23
timestamp 1624494425
transform 1 0 6203 0 1 91640
box 0 -60 2072 490
use contact_9  contact_9_60
timestamp 1624494425
transform 1 0 7680 0 1 88838
box 0 0 66 74
use contact_8  contact_8_60
timestamp 1624494425
transform 1 0 7681 0 1 88843
box 0 0 64 64
use contact_9  contact_9_600
timestamp 1624494425
transform 1 0 8076 0 1 88838
box 0 0 66 74
use contact_8  contact_8_600
timestamp 1624494425
transform 1 0 8077 0 1 88843
box 0 0 64 64
use contact_9  contact_9_56
timestamp 1624494425
transform 1 0 7680 0 1 89628
box 0 0 66 74
use contact_8  contact_8_56
timestamp 1624494425
transform 1 0 7681 0 1 89633
box 0 0 64 64
use contact_9  contact_9_58
timestamp 1624494425
transform 1 0 7680 0 1 89233
box 0 0 66 74
use contact_8  contact_8_58
timestamp 1624494425
transform 1 0 7681 0 1 89238
box 0 0 64 64
use contact_9  contact_9_594
timestamp 1624494425
transform 1 0 8076 0 1 89628
box 0 0 66 74
use contact_8  contact_8_594
timestamp 1624494425
transform 1 0 8077 0 1 89633
box 0 0 64 64
use contact_9  contact_9_597
timestamp 1624494425
transform 1 0 8076 0 1 89233
box 0 0 66 74
use contact_8  contact_8_597
timestamp 1624494425
transform 1 0 8077 0 1 89238
box 0 0 64 64
use contact_9  contact_9_54
timestamp 1624494425
transform 1 0 7680 0 1 90023
box 0 0 66 74
use contact_8  contact_8_54
timestamp 1624494425
transform 1 0 7681 0 1 90028
box 0 0 64 64
use contact_9  contact_9_591
timestamp 1624494425
transform 1 0 8076 0 1 90023
box 0 0 66 74
use contact_8  contact_8_591
timestamp 1624494425
transform 1 0 8077 0 1 90028
box 0 0 64 64
use contact_9  contact_9_50
timestamp 1624494425
transform 1 0 7680 0 1 90813
box 0 0 66 74
use contact_8  contact_8_50
timestamp 1624494425
transform 1 0 7681 0 1 90818
box 0 0 64 64
use contact_9  contact_9_52
timestamp 1624494425
transform 1 0 7680 0 1 90418
box 0 0 66 74
use contact_8  contact_8_52
timestamp 1624494425
transform 1 0 7681 0 1 90423
box 0 0 64 64
use contact_9  contact_9_585
timestamp 1624494425
transform 1 0 8076 0 1 90813
box 0 0 66 74
use contact_8  contact_8_585
timestamp 1624494425
transform 1 0 8077 0 1 90818
box 0 0 64 64
use contact_9  contact_9_588
timestamp 1624494425
transform 1 0 8076 0 1 90418
box 0 0 66 74
use contact_8  contact_8_588
timestamp 1624494425
transform 1 0 8077 0 1 90423
box 0 0 64 64
use contact_9  contact_9_46
timestamp 1624494425
transform 1 0 7680 0 1 91603
box 0 0 66 74
use contact_8  contact_8_46
timestamp 1624494425
transform 1 0 7681 0 1 91608
box 0 0 64 64
use contact_9  contact_9_48
timestamp 1624494425
transform 1 0 7680 0 1 91208
box 0 0 66 74
use contact_8  contact_8_48
timestamp 1624494425
transform 1 0 7681 0 1 91213
box 0 0 64 64
use contact_9  contact_9_579
timestamp 1624494425
transform 1 0 8076 0 1 91603
box 0 0 66 74
use contact_8  contact_8_579
timestamp 1624494425
transform 1 0 8077 0 1 91608
box 0 0 64 64
use contact_9  contact_9_582
timestamp 1624494425
transform 1 0 8076 0 1 91208
box 0 0 66 74
use contact_8  contact_8_582
timestamp 1624494425
transform 1 0 8077 0 1 91213
box 0 0 64 64
use contact_8  contact_8_578
timestamp 1624494425
transform 1 0 7299 0 1 92026
box 0 0 64 64
use contact_9  contact_9_578
timestamp 1624494425
transform 1 0 7298 0 1 92021
box 0 0 66 74
use contact_8  contact_8_577
timestamp 1624494425
transform 1 0 6867 0 1 92026
box 0 0 64 64
use contact_9  contact_9_577
timestamp 1624494425
transform 1 0 6866 0 1 92021
box 0 0 66 74
use contact_8  contact_8_45
timestamp 1624494425
transform 1 0 6442 0 1 92026
box 0 0 64 64
use contact_9  contact_9_45
timestamp 1624494425
transform 1 0 6441 0 1 92021
box 0 0 66 74
use contact_16  contact_16_69
timestamp 1624494425
transform 1 0 6104 0 1 91894
box 0 0 66 58
use contact_16  contact_16_66
timestamp 1624494425
transform 1 0 6104 0 1 92118
box 0 0 66 58
use contact_16  contact_16_67
timestamp 1624494425
transform 1 0 5064 0 1 92208
box 0 0 66 58
use contact_16  contact_16_68
timestamp 1624494425
transform 1 0 4664 0 1 92320
box 0 0 66 58
use and3_dec  and3_dec_22
timestamp 1624494425
transform 1 0 6203 0 -1 92430
box 0 -60 2072 490
use contact_8  contact_8_575
timestamp 1624494425
transform 1 0 7299 0 1 92384
box 0 0 64 64
use contact_9  contact_9_575
timestamp 1624494425
transform 1 0 7298 0 1 92379
box 0 0 66 74
use contact_8  contact_8_574
timestamp 1624494425
transform 1 0 6867 0 1 92384
box 0 0 64 64
use contact_9  contact_9_574
timestamp 1624494425
transform 1 0 6866 0 1 92379
box 0 0 66 74
use contact_8  contact_8_43
timestamp 1624494425
transform 1 0 6442 0 1 92442
box 0 0 64 64
use contact_9  contact_9_43
timestamp 1624494425
transform 1 0 6441 0 1 92437
box 0 0 66 74
use contact_16  contact_16_64
timestamp 1624494425
transform 1 0 5064 0 1 92594
box 0 0 66 58
use contact_16  contact_16_65
timestamp 1624494425
transform 1 0 4744 0 1 92482
box 0 0 66 58
use contact_8  contact_8_572
timestamp 1624494425
transform 1 0 7299 0 1 92816
box 0 0 64 64
use contact_9  contact_9_572
timestamp 1624494425
transform 1 0 7298 0 1 92811
box 0 0 66 74
use contact_8  contact_8_571
timestamp 1624494425
transform 1 0 6867 0 1 92816
box 0 0 64 64
use contact_9  contact_9_571
timestamp 1624494425
transform 1 0 6866 0 1 92811
box 0 0 66 74
use contact_8  contact_8_41
timestamp 1624494425
transform 1 0 6442 0 1 92816
box 0 0 64 64
use contact_9  contact_9_41
timestamp 1624494425
transform 1 0 6441 0 1 92811
box 0 0 66 74
use contact_16  contact_16_60
timestamp 1624494425
transform 1 0 6104 0 1 92908
box 0 0 66 58
use contact_16  contact_16_63
timestamp 1624494425
transform 1 0 6104 0 1 92684
box 0 0 66 58
use and3_dec  and3_dec_20
timestamp 1624494425
transform 1 0 6203 0 -1 93220
box 0 -60 2072 490
use and3_dec  and3_dec_21
timestamp 1624494425
transform 1 0 6203 0 1 92430
box 0 -60 2072 490
use contact_8  contact_8_569
timestamp 1624494425
transform 1 0 7299 0 1 93174
box 0 0 64 64
use contact_9  contact_9_569
timestamp 1624494425
transform 1 0 7298 0 1 93169
box 0 0 66 74
use contact_8  contact_8_568
timestamp 1624494425
transform 1 0 6867 0 1 93174
box 0 0 64 64
use contact_9  contact_9_568
timestamp 1624494425
transform 1 0 6866 0 1 93169
box 0 0 66 74
use contact_16  contact_16_61
timestamp 1624494425
transform 1 0 5064 0 1 92998
box 0 0 66 58
use contact_16  contact_16_62
timestamp 1624494425
transform 1 0 4824 0 1 93110
box 0 0 66 58
use contact_8  contact_8_39
timestamp 1624494425
transform 1 0 6442 0 1 93232
box 0 0 64 64
use contact_9  contact_9_39
timestamp 1624494425
transform 1 0 6441 0 1 93227
box 0 0 66 74
use contact_16  contact_16_58
timestamp 1624494425
transform 1 0 5144 0 1 93384
box 0 0 66 58
use contact_16  contact_16_59
timestamp 1624494425
transform 1 0 4584 0 1 93272
box 0 0 66 58
use and3_dec  and3_dec_19
timestamp 1624494425
transform 1 0 6203 0 1 93220
box 0 -60 2072 490
use contact_8  contact_8_566
timestamp 1624494425
transform 1 0 7299 0 1 93606
box 0 0 64 64
use contact_9  contact_9_566
timestamp 1624494425
transform 1 0 7298 0 1 93601
box 0 0 66 74
use contact_8  contact_8_565
timestamp 1624494425
transform 1 0 6867 0 1 93606
box 0 0 64 64
use contact_9  contact_9_565
timestamp 1624494425
transform 1 0 6866 0 1 93601
box 0 0 66 74
use contact_8  contact_8_37
timestamp 1624494425
transform 1 0 6442 0 1 93606
box 0 0 64 64
use contact_9  contact_9_37
timestamp 1624494425
transform 1 0 6441 0 1 93601
box 0 0 66 74
use contact_16  contact_16_54
timestamp 1624494425
transform 1 0 6104 0 1 93698
box 0 0 66 58
use contact_16  contact_16_57
timestamp 1624494425
transform 1 0 6104 0 1 93474
box 0 0 66 58
use contact_8  contact_8_563
timestamp 1624494425
transform 1 0 7299 0 1 93964
box 0 0 64 64
use contact_9  contact_9_563
timestamp 1624494425
transform 1 0 7298 0 1 93959
box 0 0 66 74
use contact_8  contact_8_562
timestamp 1624494425
transform 1 0 6867 0 1 93964
box 0 0 64 64
use contact_9  contact_9_562
timestamp 1624494425
transform 1 0 6866 0 1 93959
box 0 0 66 74
use contact_16  contact_16_55
timestamp 1624494425
transform 1 0 5144 0 1 93788
box 0 0 66 58
use contact_16  contact_16_56
timestamp 1624494425
transform 1 0 4664 0 1 93900
box 0 0 66 58
use and3_dec  and3_dec_17
timestamp 1624494425
transform 1 0 6203 0 1 94010
box 0 -60 2072 490
use and3_dec  and3_dec_18
timestamp 1624494425
transform 1 0 6203 0 -1 94010
box 0 -60 2072 490
use contact_8  contact_8_35
timestamp 1624494425
transform 1 0 6442 0 1 94022
box 0 0 64 64
use contact_9  contact_9_35
timestamp 1624494425
transform 1 0 6441 0 1 94017
box 0 0 66 74
use contact_16  contact_16_51
timestamp 1624494425
transform 1 0 6104 0 1 94264
box 0 0 66 58
use contact_16  contact_16_52
timestamp 1624494425
transform 1 0 5144 0 1 94174
box 0 0 66 58
use contact_16  contact_16_53
timestamp 1624494425
transform 1 0 4744 0 1 94062
box 0 0 66 58
use contact_8  contact_8_560
timestamp 1624494425
transform 1 0 7299 0 1 94396
box 0 0 64 64
use contact_9  contact_9_560
timestamp 1624494425
transform 1 0 7298 0 1 94391
box 0 0 66 74
use contact_8  contact_8_559
timestamp 1624494425
transform 1 0 6867 0 1 94396
box 0 0 64 64
use contact_9  contact_9_559
timestamp 1624494425
transform 1 0 6866 0 1 94391
box 0 0 66 74
use contact_8  contact_8_33
timestamp 1624494425
transform 1 0 6442 0 1 94396
box 0 0 64 64
use contact_9  contact_9_33
timestamp 1624494425
transform 1 0 6441 0 1 94391
box 0 0 66 74
use contact_16  contact_16_48
timestamp 1624494425
transform 1 0 6104 0 1 94488
box 0 0 66 58
use and3_dec  and3_dec_16
timestamp 1624494425
transform 1 0 6203 0 -1 94800
box 0 -60 2072 490
use contact_8  contact_8_557
timestamp 1624494425
transform 1 0 7299 0 1 94754
box 0 0 64 64
use contact_9  contact_9_557
timestamp 1624494425
transform 1 0 7298 0 1 94749
box 0 0 66 74
use contact_8  contact_8_556
timestamp 1624494425
transform 1 0 6867 0 1 94754
box 0 0 64 64
use contact_9  contact_9_556
timestamp 1624494425
transform 1 0 6866 0 1 94749
box 0 0 66 74
use contact_8  contact_8_31
timestamp 1624494425
transform 1 0 6442 0 1 94812
box 0 0 64 64
use contact_9  contact_9_31
timestamp 1624494425
transform 1 0 6441 0 1 94807
box 0 0 66 74
use contact_16  contact_16_49
timestamp 1624494425
transform 1 0 5144 0 1 94578
box 0 0 66 58
use contact_16  contact_16_50
timestamp 1624494425
transform 1 0 4824 0 1 94690
box 0 0 66 58
use contact_16  contact_16_45
timestamp 1624494425
transform 1 0 6104 0 1 95054
box 0 0 66 58
use contact_16  contact_16_46
timestamp 1624494425
transform 1 0 5224 0 1 94964
box 0 0 66 58
use contact_16  contact_16_47
timestamp 1624494425
transform 1 0 4584 0 1 94852
box 0 0 66 58
use and3_dec  and3_dec_15
timestamp 1624494425
transform 1 0 6203 0 1 94800
box 0 -60 2072 490
use contact_9  contact_9_42
timestamp 1624494425
transform 1 0 7680 0 1 92393
box 0 0 66 74
use contact_8  contact_8_42
timestamp 1624494425
transform 1 0 7681 0 1 92398
box 0 0 64 64
use contact_9  contact_9_44
timestamp 1624494425
transform 1 0 7680 0 1 91998
box 0 0 66 74
use contact_8  contact_8_44
timestamp 1624494425
transform 1 0 7681 0 1 92003
box 0 0 64 64
use contact_9  contact_9_573
timestamp 1624494425
transform 1 0 8076 0 1 92393
box 0 0 66 74
use contact_8  contact_8_573
timestamp 1624494425
transform 1 0 8077 0 1 92398
box 0 0 64 64
use contact_9  contact_9_576
timestamp 1624494425
transform 1 0 8076 0 1 91998
box 0 0 66 74
use contact_8  contact_8_576
timestamp 1624494425
transform 1 0 8077 0 1 92003
box 0 0 64 64
use contact_9  contact_9_40
timestamp 1624494425
transform 1 0 7680 0 1 92788
box 0 0 66 74
use contact_8  contact_8_40
timestamp 1624494425
transform 1 0 7681 0 1 92793
box 0 0 64 64
use contact_9  contact_9_570
timestamp 1624494425
transform 1 0 8076 0 1 92788
box 0 0 66 74
use contact_8  contact_8_570
timestamp 1624494425
transform 1 0 8077 0 1 92793
box 0 0 64 64
use contact_9  contact_9_36
timestamp 1624494425
transform 1 0 7680 0 1 93578
box 0 0 66 74
use contact_8  contact_8_36
timestamp 1624494425
transform 1 0 7681 0 1 93583
box 0 0 64 64
use contact_9  contact_9_38
timestamp 1624494425
transform 1 0 7680 0 1 93183
box 0 0 66 74
use contact_8  contact_8_38
timestamp 1624494425
transform 1 0 7681 0 1 93188
box 0 0 64 64
use contact_9  contact_9_564
timestamp 1624494425
transform 1 0 8076 0 1 93578
box 0 0 66 74
use contact_8  contact_8_564
timestamp 1624494425
transform 1 0 8077 0 1 93583
box 0 0 64 64
use contact_9  contact_9_567
timestamp 1624494425
transform 1 0 8076 0 1 93183
box 0 0 66 74
use contact_8  contact_8_567
timestamp 1624494425
transform 1 0 8077 0 1 93188
box 0 0 64 64
use contact_9  contact_9_34
timestamp 1624494425
transform 1 0 7680 0 1 93973
box 0 0 66 74
use contact_8  contact_8_34
timestamp 1624494425
transform 1 0 7681 0 1 93978
box 0 0 64 64
use contact_9  contact_9_561
timestamp 1624494425
transform 1 0 8076 0 1 93973
box 0 0 66 74
use contact_8  contact_8_561
timestamp 1624494425
transform 1 0 8077 0 1 93978
box 0 0 64 64
use contact_9  contact_9_30
timestamp 1624494425
transform 1 0 7680 0 1 94763
box 0 0 66 74
use contact_8  contact_8_30
timestamp 1624494425
transform 1 0 7681 0 1 94768
box 0 0 64 64
use contact_9  contact_9_32
timestamp 1624494425
transform 1 0 7680 0 1 94368
box 0 0 66 74
use contact_8  contact_8_32
timestamp 1624494425
transform 1 0 7681 0 1 94373
box 0 0 64 64
use contact_9  contact_9_555
timestamp 1624494425
transform 1 0 8076 0 1 94763
box 0 0 66 74
use contact_8  contact_8_555
timestamp 1624494425
transform 1 0 8077 0 1 94768
box 0 0 64 64
use contact_9  contact_9_558
timestamp 1624494425
transform 1 0 8076 0 1 94368
box 0 0 66 74
use contact_8  contact_8_558
timestamp 1624494425
transform 1 0 8077 0 1 94373
box 0 0 64 64
use contact_8  contact_8_554
timestamp 1624494425
transform 1 0 7299 0 1 95186
box 0 0 64 64
use contact_9  contact_9_554
timestamp 1624494425
transform 1 0 7298 0 1 95181
box 0 0 66 74
use contact_8  contact_8_553
timestamp 1624494425
transform 1 0 6867 0 1 95186
box 0 0 64 64
use contact_9  contact_9_553
timestamp 1624494425
transform 1 0 6866 0 1 95181
box 0 0 66 74
use contact_8  contact_8_29
timestamp 1624494425
transform 1 0 6442 0 1 95186
box 0 0 64 64
use contact_9  contact_9_29
timestamp 1624494425
transform 1 0 6441 0 1 95181
box 0 0 66 74
use contact_16  contact_16_42
timestamp 1624494425
transform 1 0 6104 0 1 95278
box 0 0 66 58
use contact_8  contact_8_551
timestamp 1624494425
transform 1 0 7299 0 1 95544
box 0 0 64 64
use contact_9  contact_9_551
timestamp 1624494425
transform 1 0 7298 0 1 95539
box 0 0 66 74
use contact_8  contact_8_550
timestamp 1624494425
transform 1 0 6867 0 1 95544
box 0 0 64 64
use contact_9  contact_9_550
timestamp 1624494425
transform 1 0 6866 0 1 95539
box 0 0 66 74
use contact_8  contact_8_27
timestamp 1624494425
transform 1 0 6442 0 1 95602
box 0 0 64 64
use contact_9  contact_9_27
timestamp 1624494425
transform 1 0 6441 0 1 95597
box 0 0 66 74
use contact_16  contact_16_43
timestamp 1624494425
transform 1 0 5224 0 1 95368
box 0 0 66 58
use contact_16  contact_16_44
timestamp 1624494425
transform 1 0 4664 0 1 95480
box 0 0 66 58
use and3_dec  and3_dec_13
timestamp 1624494425
transform 1 0 6203 0 1 95590
box 0 -60 2072 490
use and3_dec  and3_dec_14
timestamp 1624494425
transform 1 0 6203 0 -1 95590
box 0 -60 2072 490
use contact_16  contact_16_39
timestamp 1624494425
transform 1 0 6104 0 1 95844
box 0 0 66 58
use contact_16  contact_16_40
timestamp 1624494425
transform 1 0 5224 0 1 95754
box 0 0 66 58
use contact_16  contact_16_41
timestamp 1624494425
transform 1 0 4744 0 1 95642
box 0 0 66 58
use contact_8  contact_8_548
timestamp 1624494425
transform 1 0 7299 0 1 95976
box 0 0 64 64
use contact_9  contact_9_548
timestamp 1624494425
transform 1 0 7298 0 1 95971
box 0 0 66 74
use contact_8  contact_8_547
timestamp 1624494425
transform 1 0 6867 0 1 95976
box 0 0 64 64
use contact_9  contact_9_547
timestamp 1624494425
transform 1 0 6866 0 1 95971
box 0 0 66 74
use contact_8  contact_8_25
timestamp 1624494425
transform 1 0 6442 0 1 95976
box 0 0 64 64
use contact_9  contact_9_25
timestamp 1624494425
transform 1 0 6441 0 1 95971
box 0 0 66 74
use contact_16  contact_16_36
timestamp 1624494425
transform 1 0 6104 0 1 96068
box 0 0 66 58
use contact_16  contact_16_37
timestamp 1624494425
transform 1 0 5224 0 1 96158
box 0 0 66 58
use and3_dec  and3_dec_12
timestamp 1624494425
transform 1 0 6203 0 -1 96380
box 0 -60 2072 490
use contact_8  contact_8_545
timestamp 1624494425
transform 1 0 7299 0 1 96334
box 0 0 64 64
use contact_9  contact_9_545
timestamp 1624494425
transform 1 0 7298 0 1 96329
box 0 0 66 74
use contact_8  contact_8_544
timestamp 1624494425
transform 1 0 6867 0 1 96334
box 0 0 64 64
use contact_9  contact_9_544
timestamp 1624494425
transform 1 0 6866 0 1 96329
box 0 0 66 74
use contact_8  contact_8_23
timestamp 1624494425
transform 1 0 6442 0 1 96392
box 0 0 64 64
use contact_9  contact_9_23
timestamp 1624494425
transform 1 0 6441 0 1 96387
box 0 0 66 74
use contact_16  contact_16_35
timestamp 1624494425
transform 1 0 4584 0 1 96432
box 0 0 66 58
use contact_16  contact_16_38
timestamp 1624494425
transform 1 0 4824 0 1 96270
box 0 0 66 58
use contact_16  contact_16_33
timestamp 1624494425
transform 1 0 6104 0 1 96634
box 0 0 66 58
use contact_16  contact_16_34
timestamp 1624494425
transform 1 0 5304 0 1 96544
box 0 0 66 58
use and3_dec  and3_dec_10
timestamp 1624494425
transform 1 0 6203 0 -1 97170
box 0 -60 2072 490
use and3_dec  and3_dec_11
timestamp 1624494425
transform 1 0 6203 0 1 96380
box 0 -60 2072 490
use contact_8  contact_8_542
timestamp 1624494425
transform 1 0 7299 0 1 96766
box 0 0 64 64
use contact_9  contact_9_542
timestamp 1624494425
transform 1 0 7298 0 1 96761
box 0 0 66 74
use contact_8  contact_8_541
timestamp 1624494425
transform 1 0 6867 0 1 96766
box 0 0 64 64
use contact_9  contact_9_541
timestamp 1624494425
transform 1 0 6866 0 1 96761
box 0 0 66 74
use contact_8  contact_8_21
timestamp 1624494425
transform 1 0 6442 0 1 96766
box 0 0 64 64
use contact_9  contact_9_21
timestamp 1624494425
transform 1 0 6441 0 1 96761
box 0 0 66 74
use contact_16  contact_16_30
timestamp 1624494425
transform 1 0 6104 0 1 96858
box 0 0 66 58
use contact_16  contact_16_31
timestamp 1624494425
transform 1 0 5304 0 1 96948
box 0 0 66 58
use contact_8  contact_8_539
timestamp 1624494425
transform 1 0 7299 0 1 97124
box 0 0 64 64
use contact_9  contact_9_539
timestamp 1624494425
transform 1 0 7298 0 1 97119
box 0 0 66 74
use contact_8  contact_8_538
timestamp 1624494425
transform 1 0 6867 0 1 97124
box 0 0 64 64
use contact_9  contact_9_538
timestamp 1624494425
transform 1 0 6866 0 1 97119
box 0 0 66 74
use contact_8  contact_8_19
timestamp 1624494425
transform 1 0 6442 0 1 97182
box 0 0 64 64
use contact_9  contact_9_19
timestamp 1624494425
transform 1 0 6441 0 1 97177
box 0 0 66 74
use contact_16  contact_16_29
timestamp 1624494425
transform 1 0 4744 0 1 97222
box 0 0 66 58
use contact_16  contact_16_32
timestamp 1624494425
transform 1 0 4664 0 1 97060
box 0 0 66 58
use and3_dec  and3_dec_9
timestamp 1624494425
transform 1 0 6203 0 1 97170
box 0 -60 2072 490
use contact_8  contact_8_536
timestamp 1624494425
transform 1 0 7299 0 1 97556
box 0 0 64 64
use contact_9  contact_9_536
timestamp 1624494425
transform 1 0 7298 0 1 97551
box 0 0 66 74
use contact_8  contact_8_535
timestamp 1624494425
transform 1 0 6867 0 1 97556
box 0 0 64 64
use contact_9  contact_9_535
timestamp 1624494425
transform 1 0 6866 0 1 97551
box 0 0 66 74
use contact_8  contact_8_17
timestamp 1624494425
transform 1 0 6442 0 1 97556
box 0 0 64 64
use contact_9  contact_9_17
timestamp 1624494425
transform 1 0 6441 0 1 97551
box 0 0 66 74
use contact_16  contact_16_27
timestamp 1624494425
transform 1 0 6104 0 1 97424
box 0 0 66 58
use contact_16  contact_16_28
timestamp 1624494425
transform 1 0 5304 0 1 97334
box 0 0 66 58
use contact_16  contact_16_24
timestamp 1624494425
transform 1 0 6104 0 1 97648
box 0 0 66 58
use contact_16  contact_16_25
timestamp 1624494425
transform 1 0 5304 0 1 97738
box 0 0 66 58
use and3_dec  and3_dec_8
timestamp 1624494425
transform 1 0 6203 0 -1 97960
box 0 -60 2072 490
use contact_8  contact_8_533
timestamp 1624494425
transform 1 0 7299 0 1 97914
box 0 0 64 64
use contact_9  contact_9_533
timestamp 1624494425
transform 1 0 7298 0 1 97909
box 0 0 66 74
use contact_8  contact_8_532
timestamp 1624494425
transform 1 0 6867 0 1 97914
box 0 0 64 64
use contact_9  contact_9_532
timestamp 1624494425
transform 1 0 6866 0 1 97909
box 0 0 66 74
use contact_8  contact_8_15
timestamp 1624494425
transform 1 0 6442 0 1 97972
box 0 0 64 64
use contact_9  contact_9_15
timestamp 1624494425
transform 1 0 6441 0 1 97967
box 0 0 66 74
use contact_16  contact_16_23
timestamp 1624494425
transform 1 0 4584 0 1 98012
box 0 0 66 58
use contact_16  contact_16_26
timestamp 1624494425
transform 1 0 4824 0 1 97850
box 0 0 66 58
use contact_8  contact_8_530
timestamp 1624494425
transform 1 0 7299 0 1 98346
box 0 0 64 64
use contact_9  contact_9_530
timestamp 1624494425
transform 1 0 7298 0 1 98341
box 0 0 66 74
use contact_8  contact_8_529
timestamp 1624494425
transform 1 0 6867 0 1 98346
box 0 0 64 64
use contact_9  contact_9_529
timestamp 1624494425
transform 1 0 6866 0 1 98341
box 0 0 66 74
use contact_8  contact_8_13
timestamp 1624494425
transform 1 0 6442 0 1 98346
box 0 0 64 64
use contact_9  contact_9_13
timestamp 1624494425
transform 1 0 6441 0 1 98341
box 0 0 66 74
use contact_16  contact_16_21
timestamp 1624494425
transform 1 0 6104 0 1 98214
box 0 0 66 58
use contact_16  contact_16_22
timestamp 1624494425
transform 1 0 5384 0 1 98124
box 0 0 66 58
use and3_dec  and3_dec_6
timestamp 1624494425
transform 1 0 6203 0 -1 98750
box 0 -60 2072 490
use and3_dec  and3_dec_7
timestamp 1624494425
transform 1 0 6203 0 1 97960
box 0 -60 2072 490
use contact_9  contact_9_26
timestamp 1624494425
transform 1 0 7680 0 1 95553
box 0 0 66 74
use contact_8  contact_8_26
timestamp 1624494425
transform 1 0 7681 0 1 95558
box 0 0 64 64
use contact_9  contact_9_28
timestamp 1624494425
transform 1 0 7680 0 1 95158
box 0 0 66 74
use contact_8  contact_8_28
timestamp 1624494425
transform 1 0 7681 0 1 95163
box 0 0 64 64
use contact_9  contact_9_549
timestamp 1624494425
transform 1 0 8076 0 1 95553
box 0 0 66 74
use contact_8  contact_8_549
timestamp 1624494425
transform 1 0 8077 0 1 95558
box 0 0 64 64
use contact_9  contact_9_552
timestamp 1624494425
transform 1 0 8076 0 1 95158
box 0 0 66 74
use contact_8  contact_8_552
timestamp 1624494425
transform 1 0 8077 0 1 95163
box 0 0 64 64
use contact_9  contact_9_24
timestamp 1624494425
transform 1 0 7680 0 1 95948
box 0 0 66 74
use contact_8  contact_8_24
timestamp 1624494425
transform 1 0 7681 0 1 95953
box 0 0 64 64
use contact_9  contact_9_546
timestamp 1624494425
transform 1 0 8076 0 1 95948
box 0 0 66 74
use contact_8  contact_8_546
timestamp 1624494425
transform 1 0 8077 0 1 95953
box 0 0 64 64
use contact_9  contact_9_20
timestamp 1624494425
transform 1 0 7680 0 1 96738
box 0 0 66 74
use contact_8  contact_8_20
timestamp 1624494425
transform 1 0 7681 0 1 96743
box 0 0 64 64
use contact_9  contact_9_22
timestamp 1624494425
transform 1 0 7680 0 1 96343
box 0 0 66 74
use contact_8  contact_8_22
timestamp 1624494425
transform 1 0 7681 0 1 96348
box 0 0 64 64
use contact_9  contact_9_540
timestamp 1624494425
transform 1 0 8076 0 1 96738
box 0 0 66 74
use contact_8  contact_8_540
timestamp 1624494425
transform 1 0 8077 0 1 96743
box 0 0 64 64
use contact_9  contact_9_543
timestamp 1624494425
transform 1 0 8076 0 1 96343
box 0 0 66 74
use contact_8  contact_8_543
timestamp 1624494425
transform 1 0 8077 0 1 96348
box 0 0 64 64
use contact_9  contact_9_18
timestamp 1624494425
transform 1 0 7680 0 1 97133
box 0 0 66 74
use contact_8  contact_8_18
timestamp 1624494425
transform 1 0 7681 0 1 97138
box 0 0 64 64
use contact_9  contact_9_537
timestamp 1624494425
transform 1 0 8076 0 1 97133
box 0 0 66 74
use contact_8  contact_8_537
timestamp 1624494425
transform 1 0 8077 0 1 97138
box 0 0 64 64
use contact_9  contact_9_14
timestamp 1624494425
transform 1 0 7680 0 1 97923
box 0 0 66 74
use contact_8  contact_8_14
timestamp 1624494425
transform 1 0 7681 0 1 97928
box 0 0 64 64
use contact_9  contact_9_16
timestamp 1624494425
transform 1 0 7680 0 1 97528
box 0 0 66 74
use contact_8  contact_8_16
timestamp 1624494425
transform 1 0 7681 0 1 97533
box 0 0 64 64
use contact_9  contact_9_531
timestamp 1624494425
transform 1 0 8076 0 1 97923
box 0 0 66 74
use contact_8  contact_8_531
timestamp 1624494425
transform 1 0 8077 0 1 97928
box 0 0 64 64
use contact_9  contact_9_534
timestamp 1624494425
transform 1 0 8076 0 1 97528
box 0 0 66 74
use contact_8  contact_8_534
timestamp 1624494425
transform 1 0 8077 0 1 97533
box 0 0 64 64
use contact_9  contact_9_12
timestamp 1624494425
transform 1 0 7680 0 1 98318
box 0 0 66 74
use contact_8  contact_8_12
timestamp 1624494425
transform 1 0 7681 0 1 98323
box 0 0 64 64
use contact_9  contact_9_528
timestamp 1624494425
transform 1 0 8076 0 1 98318
box 0 0 66 74
use contact_8  contact_8_528
timestamp 1624494425
transform 1 0 8077 0 1 98323
box 0 0 64 64
use contact_16  contact_16_18
timestamp 1624494425
transform 1 0 6104 0 1 98438
box 0 0 66 58
use contact_16  contact_16_19
timestamp 1624494425
transform 1 0 5384 0 1 98528
box 0 0 66 58
use contact_16  contact_16_20
timestamp 1624494425
transform 1 0 4664 0 1 98640
box 0 0 66 58
use contact_8  contact_8_527
timestamp 1624494425
transform 1 0 7299 0 1 98704
box 0 0 64 64
use contact_9  contact_9_527
timestamp 1624494425
transform 1 0 7298 0 1 98699
box 0 0 66 74
use contact_8  contact_8_526
timestamp 1624494425
transform 1 0 6867 0 1 98704
box 0 0 64 64
use contact_9  contact_9_526
timestamp 1624494425
transform 1 0 6866 0 1 98699
box 0 0 66 74
use contact_8  contact_8_11
timestamp 1624494425
transform 1 0 6442 0 1 98762
box 0 0 64 64
use contact_9  contact_9_11
timestamp 1624494425
transform 1 0 6441 0 1 98757
box 0 0 66 74
use contact_16  contact_16_16
timestamp 1624494425
transform 1 0 5384 0 1 98914
box 0 0 66 58
use contact_16  contact_16_17
timestamp 1624494425
transform 1 0 4744 0 1 98802
box 0 0 66 58
use and3_dec  and3_dec_5
timestamp 1624494425
transform 1 0 6203 0 1 98750
box 0 -60 2072 490
use contact_8  contact_8_524
timestamp 1624494425
transform 1 0 7299 0 1 99136
box 0 0 64 64
use contact_9  contact_9_524
timestamp 1624494425
transform 1 0 7298 0 1 99131
box 0 0 66 74
use contact_8  contact_8_523
timestamp 1624494425
transform 1 0 6867 0 1 99136
box 0 0 64 64
use contact_9  contact_9_523
timestamp 1624494425
transform 1 0 6866 0 1 99131
box 0 0 66 74
use contact_8  contact_8_9
timestamp 1624494425
transform 1 0 6442 0 1 99136
box 0 0 64 64
use contact_9  contact_9_9
timestamp 1624494425
transform 1 0 6441 0 1 99131
box 0 0 66 74
use contact_16  contact_16_15
timestamp 1624494425
transform 1 0 6104 0 1 99004
box 0 0 66 58
use contact_16  contact_16_12
timestamp 1624494425
transform 1 0 6104 0 1 99228
box 0 0 66 58
use contact_16  contact_16_13
timestamp 1624494425
transform 1 0 5384 0 1 99318
box 0 0 66 58
use contact_16  contact_16_14
timestamp 1624494425
transform 1 0 4824 0 1 99430
box 0 0 66 58
use and3_dec  and3_dec_4
timestamp 1624494425
transform 1 0 6203 0 -1 99540
box 0 -60 2072 490
use contact_8  contact_8_521
timestamp 1624494425
transform 1 0 7299 0 1 99494
box 0 0 64 64
use contact_9  contact_9_521
timestamp 1624494425
transform 1 0 7298 0 1 99489
box 0 0 66 74
use contact_8  contact_8_520
timestamp 1624494425
transform 1 0 6867 0 1 99494
box 0 0 64 64
use contact_9  contact_9_520
timestamp 1624494425
transform 1 0 6866 0 1 99489
box 0 0 66 74
use contact_8  contact_8_7
timestamp 1624494425
transform 1 0 6442 0 1 99552
box 0 0 64 64
use contact_9  contact_9_7
timestamp 1624494425
transform 1 0 6441 0 1 99547
box 0 0 66 74
use contact_16  contact_16_10
timestamp 1624494425
transform 1 0 5464 0 1 99704
box 0 0 66 58
use contact_16  contact_16_11
timestamp 1624494425
transform 1 0 4584 0 1 99592
box 0 0 66 58
use contact_8  contact_8_518
timestamp 1624494425
transform 1 0 7299 0 1 99926
box 0 0 64 64
use contact_9  contact_9_518
timestamp 1624494425
transform 1 0 7298 0 1 99921
box 0 0 66 74
use contact_8  contact_8_517
timestamp 1624494425
transform 1 0 6867 0 1 99926
box 0 0 64 64
use contact_9  contact_9_517
timestamp 1624494425
transform 1 0 6866 0 1 99921
box 0 0 66 74
use contact_8  contact_8_5
timestamp 1624494425
transform 1 0 6442 0 1 99926
box 0 0 64 64
use contact_9  contact_9_5
timestamp 1624494425
transform 1 0 6441 0 1 99921
box 0 0 66 74
use contact_16  contact_16_6
timestamp 1624494425
transform 1 0 6104 0 1 100018
box 0 0 66 58
use contact_16  contact_16_9
timestamp 1624494425
transform 1 0 6104 0 1 99794
box 0 0 66 58
use and3_dec  and3_dec_2
timestamp 1624494425
transform 1 0 6203 0 -1 100330
box 0 -60 2072 490
use and3_dec  and3_dec_3
timestamp 1624494425
transform 1 0 6203 0 1 99540
box 0 -60 2072 490
use contact_8  contact_8_515
timestamp 1624494425
transform 1 0 7299 0 1 100284
box 0 0 64 64
use contact_9  contact_9_515
timestamp 1624494425
transform 1 0 7298 0 1 100279
box 0 0 66 74
use contact_8  contact_8_514
timestamp 1624494425
transform 1 0 6867 0 1 100284
box 0 0 64 64
use contact_9  contact_9_514
timestamp 1624494425
transform 1 0 6866 0 1 100279
box 0 0 66 74
use contact_16  contact_16_7
timestamp 1624494425
transform 1 0 5464 0 1 100108
box 0 0 66 58
use contact_16  contact_16_8
timestamp 1624494425
transform 1 0 4664 0 1 100220
box 0 0 66 58
use contact_8  contact_8_3
timestamp 1624494425
transform 1 0 6442 0 1 100342
box 0 0 64 64
use contact_9  contact_9_3
timestamp 1624494425
transform 1 0 6441 0 1 100337
box 0 0 66 74
use contact_16  contact_16_4
timestamp 1624494425
transform 1 0 5464 0 1 100494
box 0 0 66 58
use contact_16  contact_16_5
timestamp 1624494425
transform 1 0 4744 0 1 100382
box 0 0 66 58
use and3_dec  and3_dec_1
timestamp 1624494425
transform 1 0 6203 0 1 100330
box 0 -60 2072 490
use contact_8  contact_8_512
timestamp 1624494425
transform 1 0 7299 0 1 100716
box 0 0 64 64
use contact_9  contact_9_512
timestamp 1624494425
transform 1 0 7298 0 1 100711
box 0 0 66 74
use contact_8  contact_8_511
timestamp 1624494425
transform 1 0 6867 0 1 100716
box 0 0 64 64
use contact_9  contact_9_511
timestamp 1624494425
transform 1 0 6866 0 1 100711
box 0 0 66 74
use contact_8  contact_8_1
timestamp 1624494425
transform 1 0 6442 0 1 100716
box 0 0 64 64
use contact_9  contact_9_1
timestamp 1624494425
transform 1 0 6441 0 1 100711
box 0 0 66 74
use contact_16  contact_16_0
timestamp 1624494425
transform 1 0 6104 0 1 100808
box 0 0 66 58
use contact_16  contact_16_3
timestamp 1624494425
transform 1 0 6104 0 1 100584
box 0 0 66 58
use contact_16  contact_16_1
timestamp 1624494425
transform 1 0 5464 0 1 100898
box 0 0 66 58
use contact_16  contact_16_2
timestamp 1624494425
transform 1 0 4824 0 1 101010
box 0 0 66 58
use and3_dec  and3_dec_0
timestamp 1624494425
transform 1 0 6203 0 -1 101120
box 0 -60 2072 490
use contact_9  contact_9_10
timestamp 1624494425
transform 1 0 7680 0 1 98713
box 0 0 66 74
use contact_8  contact_8_10
timestamp 1624494425
transform 1 0 7681 0 1 98718
box 0 0 64 64
use contact_9  contact_9_525
timestamp 1624494425
transform 1 0 8076 0 1 98713
box 0 0 66 74
use contact_8  contact_8_525
timestamp 1624494425
transform 1 0 8077 0 1 98718
box 0 0 64 64
use contact_9  contact_9_6
timestamp 1624494425
transform 1 0 7680 0 1 99503
box 0 0 66 74
use contact_8  contact_8_6
timestamp 1624494425
transform 1 0 7681 0 1 99508
box 0 0 64 64
use contact_9  contact_9_8
timestamp 1624494425
transform 1 0 7680 0 1 99108
box 0 0 66 74
use contact_8  contact_8_8
timestamp 1624494425
transform 1 0 7681 0 1 99113
box 0 0 64 64
use contact_9  contact_9_519
timestamp 1624494425
transform 1 0 8076 0 1 99503
box 0 0 66 74
use contact_8  contact_8_519
timestamp 1624494425
transform 1 0 8077 0 1 99508
box 0 0 64 64
use contact_9  contact_9_522
timestamp 1624494425
transform 1 0 8076 0 1 99108
box 0 0 66 74
use contact_8  contact_8_522
timestamp 1624494425
transform 1 0 8077 0 1 99113
box 0 0 64 64
use contact_9  contact_9_2
timestamp 1624494425
transform 1 0 7680 0 1 100293
box 0 0 66 74
use contact_8  contact_8_2
timestamp 1624494425
transform 1 0 7681 0 1 100298
box 0 0 64 64
use contact_9  contact_9_4
timestamp 1624494425
transform 1 0 7680 0 1 99898
box 0 0 66 74
use contact_8  contact_8_4
timestamp 1624494425
transform 1 0 7681 0 1 99903
box 0 0 64 64
use contact_9  contact_9_513
timestamp 1624494425
transform 1 0 8076 0 1 100293
box 0 0 66 74
use contact_8  contact_8_513
timestamp 1624494425
transform 1 0 8077 0 1 100298
box 0 0 64 64
use contact_9  contact_9_516
timestamp 1624494425
transform 1 0 8076 0 1 99898
box 0 0 66 74
use contact_8  contact_8_516
timestamp 1624494425
transform 1 0 8077 0 1 99903
box 0 0 64 64
use contact_9  contact_9_0
timestamp 1624494425
transform 1 0 7680 0 1 100688
box 0 0 66 74
use contact_8  contact_8_0
timestamp 1624494425
transform 1 0 7681 0 1 100693
box 0 0 64 64
use contact_9  contact_9_510
timestamp 1624494425
transform 1 0 8076 0 1 100688
box 0 0 66 74
use contact_8  contact_8_510
timestamp 1624494425
transform 1 0 8077 0 1 100693
box 0 0 64 64
<< labels >>
rlabel metal1 s 19 0 47 9480 4 addr_0
rlabel metal1 s 99 0 127 9480 4 addr_1
rlabel metal1 s 179 0 207 9480 4 addr_2
rlabel metal1 s 259 0 287 9480 4 addr_3
rlabel metal1 s 339 0 367 9480 4 addr_4
rlabel metal1 s 419 0 447 9480 4 addr_5
rlabel metal1 s 499 0 527 9480 4 addr_6
rlabel metal1 s 579 0 607 9480 4 addr_7
rlabel locali s 7968 120 7968 120 4 decode_0
rlabel locali s 7968 670 7968 670 4 decode_1
rlabel locali s 7968 910 7968 910 4 decode_2
rlabel locali s 7968 1460 7968 1460 4 decode_3
rlabel locali s 7968 1700 7968 1700 4 decode_4
rlabel locali s 7968 2250 7968 2250 4 decode_5
rlabel locali s 7968 2490 7968 2490 4 decode_6
rlabel locali s 7968 3040 7968 3040 4 decode_7
rlabel locali s 7968 3280 7968 3280 4 decode_8
rlabel locali s 7968 3830 7968 3830 4 decode_9
rlabel locali s 7968 4070 7968 4070 4 decode_10
rlabel locali s 7968 4620 7968 4620 4 decode_11
rlabel locali s 7968 4860 7968 4860 4 decode_12
rlabel locali s 7968 5410 7968 5410 4 decode_13
rlabel locali s 7968 5650 7968 5650 4 decode_14
rlabel locali s 7968 6200 7968 6200 4 decode_15
rlabel locali s 7968 6440 7968 6440 4 decode_16
rlabel locali s 7968 6990 7968 6990 4 decode_17
rlabel locali s 7968 7230 7968 7230 4 decode_18
rlabel locali s 7968 7780 7968 7780 4 decode_19
rlabel locali s 7968 8020 7968 8020 4 decode_20
rlabel locali s 7968 8570 7968 8570 4 decode_21
rlabel locali s 7968 8810 7968 8810 4 decode_22
rlabel locali s 7968 9360 7968 9360 4 decode_23
rlabel locali s 7968 9600 7968 9600 4 decode_24
rlabel locali s 7968 10150 7968 10150 4 decode_25
rlabel locali s 7968 10390 7968 10390 4 decode_26
rlabel locali s 7968 10940 7968 10940 4 decode_27
rlabel locali s 7968 11180 7968 11180 4 decode_28
rlabel locali s 7968 11730 7968 11730 4 decode_29
rlabel locali s 7968 11970 7968 11970 4 decode_30
rlabel locali s 7968 12520 7968 12520 4 decode_31
rlabel locali s 7968 12760 7968 12760 4 decode_32
rlabel locali s 7968 13310 7968 13310 4 decode_33
rlabel locali s 7968 13550 7968 13550 4 decode_34
rlabel locali s 7968 14100 7968 14100 4 decode_35
rlabel locali s 7968 14340 7968 14340 4 decode_36
rlabel locali s 7968 14890 7968 14890 4 decode_37
rlabel locali s 7968 15130 7968 15130 4 decode_38
rlabel locali s 7968 15680 7968 15680 4 decode_39
rlabel locali s 7968 15920 7968 15920 4 decode_40
rlabel locali s 7968 16470 7968 16470 4 decode_41
rlabel locali s 7968 16710 7968 16710 4 decode_42
rlabel locali s 7968 17260 7968 17260 4 decode_43
rlabel locali s 7968 17500 7968 17500 4 decode_44
rlabel locali s 7968 18050 7968 18050 4 decode_45
rlabel locali s 7968 18290 7968 18290 4 decode_46
rlabel locali s 7968 18840 7968 18840 4 decode_47
rlabel locali s 7968 19080 7968 19080 4 decode_48
rlabel locali s 7968 19630 7968 19630 4 decode_49
rlabel locali s 7968 19870 7968 19870 4 decode_50
rlabel locali s 7968 20420 7968 20420 4 decode_51
rlabel locali s 7968 20660 7968 20660 4 decode_52
rlabel locali s 7968 21210 7968 21210 4 decode_53
rlabel locali s 7968 21450 7968 21450 4 decode_54
rlabel locali s 7968 22000 7968 22000 4 decode_55
rlabel locali s 7968 22240 7968 22240 4 decode_56
rlabel locali s 7968 22790 7968 22790 4 decode_57
rlabel locali s 7968 23030 7968 23030 4 decode_58
rlabel locali s 7968 23580 7968 23580 4 decode_59
rlabel locali s 7968 23820 7968 23820 4 decode_60
rlabel locali s 7968 24370 7968 24370 4 decode_61
rlabel locali s 7968 24610 7968 24610 4 decode_62
rlabel locali s 7968 25160 7968 25160 4 decode_63
rlabel locali s 7968 25400 7968 25400 4 decode_64
rlabel locali s 7968 25950 7968 25950 4 decode_65
rlabel locali s 7968 26190 7968 26190 4 decode_66
rlabel locali s 7968 26740 7968 26740 4 decode_67
rlabel locali s 7968 26980 7968 26980 4 decode_68
rlabel locali s 7968 27530 7968 27530 4 decode_69
rlabel locali s 7968 27770 7968 27770 4 decode_70
rlabel locali s 7968 28320 7968 28320 4 decode_71
rlabel locali s 7968 28560 7968 28560 4 decode_72
rlabel locali s 7968 29110 7968 29110 4 decode_73
rlabel locali s 7968 29350 7968 29350 4 decode_74
rlabel locali s 7968 29900 7968 29900 4 decode_75
rlabel locali s 7968 30140 7968 30140 4 decode_76
rlabel locali s 7968 30690 7968 30690 4 decode_77
rlabel locali s 7968 30930 7968 30930 4 decode_78
rlabel locali s 7968 31480 7968 31480 4 decode_79
rlabel locali s 7968 31720 7968 31720 4 decode_80
rlabel locali s 7968 32270 7968 32270 4 decode_81
rlabel locali s 7968 32510 7968 32510 4 decode_82
rlabel locali s 7968 33060 7968 33060 4 decode_83
rlabel locali s 7968 33300 7968 33300 4 decode_84
rlabel locali s 7968 33850 7968 33850 4 decode_85
rlabel locali s 7968 34090 7968 34090 4 decode_86
rlabel locali s 7968 34640 7968 34640 4 decode_87
rlabel locali s 7968 34880 7968 34880 4 decode_88
rlabel locali s 7968 35430 7968 35430 4 decode_89
rlabel locali s 7968 35670 7968 35670 4 decode_90
rlabel locali s 7968 36220 7968 36220 4 decode_91
rlabel locali s 7968 36460 7968 36460 4 decode_92
rlabel locali s 7968 37010 7968 37010 4 decode_93
rlabel locali s 7968 37250 7968 37250 4 decode_94
rlabel locali s 7968 37800 7968 37800 4 decode_95
rlabel locali s 7968 38040 7968 38040 4 decode_96
rlabel locali s 7968 38590 7968 38590 4 decode_97
rlabel locali s 7968 38830 7968 38830 4 decode_98
rlabel locali s 7968 39380 7968 39380 4 decode_99
rlabel locali s 7968 39620 7968 39620 4 decode_100
rlabel locali s 7968 40170 7968 40170 4 decode_101
rlabel locali s 7968 40410 7968 40410 4 decode_102
rlabel locali s 7968 40960 7968 40960 4 decode_103
rlabel locali s 7968 41200 7968 41200 4 decode_104
rlabel locali s 7968 41750 7968 41750 4 decode_105
rlabel locali s 7968 41990 7968 41990 4 decode_106
rlabel locali s 7968 42540 7968 42540 4 decode_107
rlabel locali s 7968 42780 7968 42780 4 decode_108
rlabel locali s 7968 43330 7968 43330 4 decode_109
rlabel locali s 7968 43570 7968 43570 4 decode_110
rlabel locali s 7968 44120 7968 44120 4 decode_111
rlabel locali s 7968 44360 7968 44360 4 decode_112
rlabel locali s 7968 44910 7968 44910 4 decode_113
rlabel locali s 7968 45150 7968 45150 4 decode_114
rlabel locali s 7968 45700 7968 45700 4 decode_115
rlabel locali s 7968 45940 7968 45940 4 decode_116
rlabel locali s 7968 46490 7968 46490 4 decode_117
rlabel locali s 7968 46730 7968 46730 4 decode_118
rlabel locali s 7968 47280 7968 47280 4 decode_119
rlabel locali s 7968 47520 7968 47520 4 decode_120
rlabel locali s 7968 48070 7968 48070 4 decode_121
rlabel locali s 7968 48310 7968 48310 4 decode_122
rlabel locali s 7968 48860 7968 48860 4 decode_123
rlabel locali s 7968 49100 7968 49100 4 decode_124
rlabel locali s 7968 49650 7968 49650 4 decode_125
rlabel locali s 7968 49890 7968 49890 4 decode_126
rlabel locali s 7968 50440 7968 50440 4 decode_127
rlabel locali s 7968 50680 7968 50680 4 decode_128
rlabel locali s 7968 51230 7968 51230 4 decode_129
rlabel locali s 7968 51470 7968 51470 4 decode_130
rlabel locali s 7968 52020 7968 52020 4 decode_131
rlabel locali s 7968 52260 7968 52260 4 decode_132
rlabel locali s 7968 52810 7968 52810 4 decode_133
rlabel locali s 7968 53050 7968 53050 4 decode_134
rlabel locali s 7968 53600 7968 53600 4 decode_135
rlabel locali s 7968 53840 7968 53840 4 decode_136
rlabel locali s 7968 54390 7968 54390 4 decode_137
rlabel locali s 7968 54630 7968 54630 4 decode_138
rlabel locali s 7968 55180 7968 55180 4 decode_139
rlabel locali s 7968 55420 7968 55420 4 decode_140
rlabel locali s 7968 55970 7968 55970 4 decode_141
rlabel locali s 7968 56210 7968 56210 4 decode_142
rlabel locali s 7968 56760 7968 56760 4 decode_143
rlabel locali s 7968 57000 7968 57000 4 decode_144
rlabel locali s 7968 57550 7968 57550 4 decode_145
rlabel locali s 7968 57790 7968 57790 4 decode_146
rlabel locali s 7968 58340 7968 58340 4 decode_147
rlabel locali s 7968 58580 7968 58580 4 decode_148
rlabel locali s 7968 59130 7968 59130 4 decode_149
rlabel locali s 7968 59370 7968 59370 4 decode_150
rlabel locali s 7968 59920 7968 59920 4 decode_151
rlabel locali s 7968 60160 7968 60160 4 decode_152
rlabel locali s 7968 60710 7968 60710 4 decode_153
rlabel locali s 7968 60950 7968 60950 4 decode_154
rlabel locali s 7968 61500 7968 61500 4 decode_155
rlabel locali s 7968 61740 7968 61740 4 decode_156
rlabel locali s 7968 62290 7968 62290 4 decode_157
rlabel locali s 7968 62530 7968 62530 4 decode_158
rlabel locali s 7968 63080 7968 63080 4 decode_159
rlabel locali s 7968 63320 7968 63320 4 decode_160
rlabel locali s 7968 63870 7968 63870 4 decode_161
rlabel locali s 7968 64110 7968 64110 4 decode_162
rlabel locali s 7968 64660 7968 64660 4 decode_163
rlabel locali s 7968 64900 7968 64900 4 decode_164
rlabel locali s 7968 65450 7968 65450 4 decode_165
rlabel locali s 7968 65690 7968 65690 4 decode_166
rlabel locali s 7968 66240 7968 66240 4 decode_167
rlabel locali s 7968 66480 7968 66480 4 decode_168
rlabel locali s 7968 67030 7968 67030 4 decode_169
rlabel locali s 7968 67270 7968 67270 4 decode_170
rlabel locali s 7968 67820 7968 67820 4 decode_171
rlabel locali s 7968 68060 7968 68060 4 decode_172
rlabel locali s 7968 68610 7968 68610 4 decode_173
rlabel locali s 7968 68850 7968 68850 4 decode_174
rlabel locali s 7968 69400 7968 69400 4 decode_175
rlabel locali s 7968 69640 7968 69640 4 decode_176
rlabel locali s 7968 70190 7968 70190 4 decode_177
rlabel locali s 7968 70430 7968 70430 4 decode_178
rlabel locali s 7968 70980 7968 70980 4 decode_179
rlabel locali s 7968 71220 7968 71220 4 decode_180
rlabel locali s 7968 71770 7968 71770 4 decode_181
rlabel locali s 7968 72010 7968 72010 4 decode_182
rlabel locali s 7968 72560 7968 72560 4 decode_183
rlabel locali s 7968 72800 7968 72800 4 decode_184
rlabel locali s 7968 73350 7968 73350 4 decode_185
rlabel locali s 7968 73590 7968 73590 4 decode_186
rlabel locali s 7968 74140 7968 74140 4 decode_187
rlabel locali s 7968 74380 7968 74380 4 decode_188
rlabel locali s 7968 74930 7968 74930 4 decode_189
rlabel locali s 7968 75170 7968 75170 4 decode_190
rlabel locali s 7968 75720 7968 75720 4 decode_191
rlabel locali s 7968 75960 7968 75960 4 decode_192
rlabel locali s 7968 76510 7968 76510 4 decode_193
rlabel locali s 7968 76750 7968 76750 4 decode_194
rlabel locali s 7968 77300 7968 77300 4 decode_195
rlabel locali s 7968 77540 7968 77540 4 decode_196
rlabel locali s 7968 78090 7968 78090 4 decode_197
rlabel locali s 7968 78330 7968 78330 4 decode_198
rlabel locali s 7968 78880 7968 78880 4 decode_199
rlabel locali s 7968 79120 7968 79120 4 decode_200
rlabel locali s 7968 79670 7968 79670 4 decode_201
rlabel locali s 7968 79910 7968 79910 4 decode_202
rlabel locali s 7968 80460 7968 80460 4 decode_203
rlabel locali s 7968 80700 7968 80700 4 decode_204
rlabel locali s 7968 81250 7968 81250 4 decode_205
rlabel locali s 7968 81490 7968 81490 4 decode_206
rlabel locali s 7968 82040 7968 82040 4 decode_207
rlabel locali s 7968 82280 7968 82280 4 decode_208
rlabel locali s 7968 82830 7968 82830 4 decode_209
rlabel locali s 7968 83070 7968 83070 4 decode_210
rlabel locali s 7968 83620 7968 83620 4 decode_211
rlabel locali s 7968 83860 7968 83860 4 decode_212
rlabel locali s 7968 84410 7968 84410 4 decode_213
rlabel locali s 7968 84650 7968 84650 4 decode_214
rlabel locali s 7968 85200 7968 85200 4 decode_215
rlabel locali s 7968 85440 7968 85440 4 decode_216
rlabel locali s 7968 85990 7968 85990 4 decode_217
rlabel locali s 7968 86230 7968 86230 4 decode_218
rlabel locali s 7968 86780 7968 86780 4 decode_219
rlabel locali s 7968 87020 7968 87020 4 decode_220
rlabel locali s 7968 87570 7968 87570 4 decode_221
rlabel locali s 7968 87810 7968 87810 4 decode_222
rlabel locali s 7968 88360 7968 88360 4 decode_223
rlabel locali s 7968 88600 7968 88600 4 decode_224
rlabel locali s 7968 89150 7968 89150 4 decode_225
rlabel locali s 7968 89390 7968 89390 4 decode_226
rlabel locali s 7968 89940 7968 89940 4 decode_227
rlabel locali s 7968 90180 7968 90180 4 decode_228
rlabel locali s 7968 90730 7968 90730 4 decode_229
rlabel locali s 7968 90970 7968 90970 4 decode_230
rlabel locali s 7968 91520 7968 91520 4 decode_231
rlabel locali s 7968 91760 7968 91760 4 decode_232
rlabel locali s 7968 92310 7968 92310 4 decode_233
rlabel locali s 7968 92550 7968 92550 4 decode_234
rlabel locali s 7968 93100 7968 93100 4 decode_235
rlabel locali s 7968 93340 7968 93340 4 decode_236
rlabel locali s 7968 93890 7968 93890 4 decode_237
rlabel locali s 7968 94130 7968 94130 4 decode_238
rlabel locali s 7968 94680 7968 94680 4 decode_239
rlabel locali s 7968 94920 7968 94920 4 decode_240
rlabel locali s 7968 95470 7968 95470 4 decode_241
rlabel locali s 7968 95710 7968 95710 4 decode_242
rlabel locali s 7968 96260 7968 96260 4 decode_243
rlabel locali s 7968 96500 7968 96500 4 decode_244
rlabel locali s 7968 97050 7968 97050 4 decode_245
rlabel locali s 7968 97290 7968 97290 4 decode_246
rlabel locali s 7968 97840 7968 97840 4 decode_247
rlabel locali s 7968 98080 7968 98080 4 decode_248
rlabel locali s 7968 98630 7968 98630 4 decode_249
rlabel locali s 7968 98870 7968 98870 4 decode_250
rlabel locali s 7968 99420 7968 99420 4 decode_251
rlabel locali s 7968 99660 7968 99660 4 decode_252
rlabel locali s 7968 100210 7968 100210 4 decode_253
rlabel locali s 7968 100450 7968 100450 4 decode_254
rlabel locali s 7968 101000 7968 101000 4 decode_255
rlabel metal1 s 4603 0 4631 101148 4 predecode_0
rlabel metal1 s 4683 0 4711 101148 4 predecode_1
rlabel metal1 s 4763 0 4791 101148 4 predecode_2
rlabel metal1 s 4843 0 4871 101148 4 predecode_3
rlabel metal1 s 4923 0 4951 101148 4 predecode_4
rlabel metal1 s 5003 0 5031 101148 4 predecode_5
rlabel metal1 s 5083 0 5111 101148 4 predecode_6
rlabel metal1 s 5163 0 5191 101148 4 predecode_7
rlabel metal1 s 5243 0 5271 101148 4 predecode_8
rlabel metal1 s 5323 0 5351 101148 4 predecode_9
rlabel metal1 s 5403 0 5431 101148 4 predecode_10
rlabel metal1 s 5483 0 5511 101148 4 predecode_11
rlabel metal1 s 5563 0 5591 101148 4 predecode_12
rlabel metal1 s 5643 0 5671 101148 4 predecode_13
rlabel metal1 s 5723 0 5751 101148 4 predecode_14
rlabel metal1 s 5803 0 5831 101148 4 predecode_15
rlabel metal1 s 5883 0 5911 101148 4 predecode_16
rlabel metal1 s 5963 0 5991 101148 4 predecode_17
rlabel metal1 s 6043 0 6071 101148 4 predecode_18
rlabel metal1 s 6123 0 6151 101148 4 predecode_19
rlabel metal3 s 6850 85689 6948 85787 4 vdd
rlabel metal3 s 3116 5109 3214 5207 4 vdd
rlabel metal3 s 6850 60767 6948 60865 4 vdd
rlabel metal3 s 8060 57226 8158 57324 4 vdd
rlabel metal3 s 8060 78556 8158 78654 4 vdd
rlabel metal3 s 6850 71469 6948 71567 4 vdd
rlabel metal3 s 7282 96749 7380 96847 4 vdd
rlabel metal3 s 8060 81321 8158 81419 4 vdd
rlabel metal3 s 8060 9826 8158 9924 4 vdd
rlabel metal3 s 6850 54447 6948 54545 4 vdd
rlabel metal3 s 8060 54066 8158 54164 4 vdd
rlabel metal3 s 6850 46189 6948 46287 4 vdd
rlabel metal3 s 6850 92009 6948 92107 4 vdd
rlabel metal3 s 6850 5109 6948 5207 4 vdd
rlabel metal3 s 7282 98329 7380 98427 4 vdd
rlabel metal3 s 6850 95959 6948 96057 4 vdd
rlabel metal3 s 8060 346 8158 444 4 vdd
rlabel metal3 s 6850 35487 6948 35585 4 vdd
rlabel metal3 s 7282 43387 7380 43485 4 vdd
rlabel metal3 s 8060 36686 8158 36784 4 vdd
rlabel metal3 s 6850 77789 6948 77887 4 vdd
rlabel metal3 s 7282 45399 7380 45497 4 vdd
rlabel metal3 s 8060 61176 8158 61274 4 vdd
rlabel metal3 s 7282 6257 7380 6355 4 vdd
rlabel metal3 s 6850 19687 6948 19785 4 vdd
rlabel metal3 s 6850 34339 6948 34437 4 vdd
rlabel metal3 s 6850 75419 6948 75517 4 vdd
rlabel metal3 s 8060 1531 8158 1629 4 vdd
rlabel metal3 s 6850 9059 6948 9157 4 vdd
rlabel metal3 s 7282 85689 7380 85787 4 vdd
rlabel metal3 s 6850 10997 6948 11095 4 vdd
rlabel metal3 s 7282 5109 7380 5207 4 vdd
rlabel metal3 s 8060 75791 8158 75889 4 vdd
rlabel metal3 s 6850 80159 6948 80257 4 vdd
rlabel metal3 s 6850 91219 6948 91317 4 vdd
rlabel metal3 s 6850 56817 6948 56915 4 vdd
rlabel metal3 s 7282 97539 7380 97637 4 vdd
rlabel metal3 s 7282 9059 7380 9157 4 vdd
rlabel metal3 s 6850 58039 6948 58137 4 vdd
rlabel metal3 s 8060 45771 8158 45869 4 vdd
rlabel metal3 s 6850 55669 6948 55767 4 vdd
rlabel metal3 s 7282 91219 7380 91317 4 vdd
rlabel metal3 s 8060 39056 8158 39154 4 vdd
rlabel metal3 s 6850 32759 6948 32857 4 vdd
rlabel metal3 s 7282 8627 7380 8725 4 vdd
rlabel metal3 s 4326 8246 4424 8344 4 vdd
rlabel metal3 s 7282 24427 7380 24525 4 vdd
rlabel metal3 s 7282 12219 7380 12317 4 vdd
rlabel metal3 s 6850 51287 6948 51385 4 vdd
rlabel metal3 s 6850 92367 6948 92465 4 vdd
rlabel metal3 s 8060 56436 8158 56534 4 vdd
rlabel metal3 s 7282 18897 7380 18995 4 vdd
rlabel metal3 s 8060 24441 8158 24539 4 vdd
rlabel metal3 s 8060 46166 8158 46264 4 vdd
rlabel metal3 s 8060 58016 8158 58114 4 vdd
rlabel metal3 s 8060 98306 8158 98404 4 vdd
rlabel metal3 s 7282 73049 7380 73147 4 vdd
rlabel metal3 s 3548 9059 3646 9157 4 vdd
rlabel metal3 s 7282 9849 7380 9947 4 vdd
rlabel metal3 s 6850 31179 6948 31277 4 vdd
rlabel metal3 s 7282 83319 7380 83417 4 vdd
rlabel metal3 s 7282 82097 7380 82195 4 vdd
rlabel metal3 s 8060 89221 8158 89319 4 vdd
rlabel metal3 s 6850 55237 6948 55335 4 vdd
rlabel metal3 s 6850 62347 6948 62445 4 vdd
rlabel metal3 s 8060 80531 8158 80629 4 vdd
rlabel metal3 s 6850 49349 6948 49447 4 vdd
rlabel metal3 s 7282 47337 7380 47435 4 vdd
rlabel metal3 s 8060 73026 8158 73124 4 vdd
rlabel metal3 s 8060 69866 8158 69964 4 vdd
rlabel metal3 s 6850 86047 6948 86145 4 vdd
rlabel metal3 s 8060 96331 8158 96429 4 vdd
rlabel metal3 s 6850 54879 6948 54977 4 vdd
rlabel metal3 s 4326 3506 4424 3604 4 vdd
rlabel metal3 s 3116 7479 3214 7577 4 vdd
rlabel metal3 s 7282 99477 7380 99575 4 vdd
rlabel metal3 s 8060 35501 8158 35599 4 vdd
rlabel metal3 s 8060 55251 8158 55349 4 vdd
rlabel metal3 s 6850 44609 6948 44707 4 vdd
rlabel metal3 s 8060 52486 8158 52584 4 vdd
rlabel metal3 s 8060 68286 8158 68384 4 vdd
rlabel metal3 s 8060 84086 8158 84184 4 vdd
rlabel metal3 s 8060 14961 8158 15059 4 vdd
rlabel metal3 s 7282 62779 7380 62877 4 vdd
rlabel metal3 s 7282 87269 7380 87367 4 vdd
rlabel metal3 s 6850 51719 6948 51817 4 vdd
rlabel metal3 s 7282 1159 7380 1257 4 vdd
rlabel metal3 s 6850 16527 6948 16625 4 vdd
rlabel metal3 s 8060 90406 8158 90504 4 vdd
rlabel metal3 s 6850 13367 6948 13465 4 vdd
rlabel metal3 s 6850 40659 6948 40757 4 vdd
rlabel metal3 s 3116 6689 3214 6787 4 vdd
rlabel metal3 s 8060 63151 8158 63249 4 vdd
rlabel metal3 s 7282 30747 7380 30845 4 vdd
rlabel metal3 s 7282 42597 7380 42695 4 vdd
rlabel metal3 s 7282 22489 7380 22587 4 vdd
rlabel metal3 s 3548 7479 3646 7577 4 vdd
rlabel metal3 s 6850 4319 6948 4417 4 vdd
rlabel metal3 s 8060 91986 8158 92084 4 vdd
rlabel metal3 s 7282 89639 7380 89737 4 vdd
rlabel metal3 s 7282 1517 7380 1615 4 vdd
rlabel metal3 s 7282 77789 7380 77887 4 vdd
rlabel metal3 s 7282 20119 7380 20217 4 vdd
rlabel metal3 s 8060 85666 8158 85764 4 vdd
rlabel metal3 s 7282 74987 7380 75085 4 vdd
rlabel metal3 s 7282 98687 7380 98785 4 vdd
rlabel metal3 s 6850 71037 6948 71135 4 vdd
rlabel metal3 s 6850 21699 6948 21797 4 vdd
rlabel metal3 s 8060 17726 8158 17824 4 vdd
rlabel metal3 s 7282 26797 7380 26895 4 vdd
rlabel metal3 s 8060 1926 8158 2024 4 vdd
rlabel metal3 s 6850 22489 6948 22587 4 vdd
rlabel metal3 s 6850 50139 6948 50237 4 vdd
rlabel metal3 s 6850 97539 6948 97637 4 vdd
rlabel metal3 s 7282 76567 7380 76665 4 vdd
rlabel metal3 s 7282 71469 7380 71567 4 vdd
rlabel metal3 s 6850 90429 6948 90527 4 vdd
rlabel metal3 s 7282 34697 7380 34795 4 vdd
rlabel metal3 s 7282 100267 7380 100365 4 vdd
rlabel metal3 s 6850 58397 6948 58495 4 vdd
rlabel metal3 s 8060 58411 8158 58509 4 vdd
rlabel metal3 s 7282 13009 7380 13107 4 vdd
rlabel metal3 s 7282 12577 7380 12675 4 vdd
rlabel metal3 s 7282 72617 7380 72715 4 vdd
rlabel metal3 s 7282 2307 7380 2405 4 vdd
rlabel metal3 s 7282 35487 7380 35585 4 vdd
rlabel metal3 s 8060 16936 8158 17034 4 vdd
rlabel metal3 s 6850 22847 6948 22945 4 vdd
rlabel metal3 s 6850 76567 6948 76665 4 vdd
rlabel metal3 s 8060 58806 8158 58904 4 vdd
rlabel metal3 s 7282 79369 7380 79467 4 vdd
rlabel metal3 s 7282 92009 7380 92107 4 vdd
rlabel metal3 s 7282 71827 7380 71925 4 vdd
rlabel metal3 s 7282 61199 7380 61297 4 vdd
rlabel metal3 s 3548 8269 3646 8367 4 vdd
rlabel metal3 s 6850 1517 6948 1615 4 vdd
rlabel metal3 s 6850 11787 6948 11885 4 vdd
rlabel metal3 s 6850 46547 6948 46645 4 vdd
rlabel metal3 s 8060 46561 8158 46659 4 vdd
rlabel metal3 s 8060 52091 8158 52189 4 vdd
rlabel metal3 s 8060 71841 8158 71939 4 vdd
rlabel metal3 s 8060 37871 8158 37969 4 vdd
rlabel metal3 s 7282 43819 7380 43917 4 vdd
rlabel metal3 s 8060 5876 8158 5974 4 vdd
rlabel metal3 s 7282 48559 7380 48657 4 vdd
rlabel metal3 s 8060 62361 8158 62459 4 vdd
rlabel metal3 s 8060 32341 8158 32439 4 vdd
rlabel metal3 s 8060 41426 8158 41524 4 vdd
rlabel metal3 s 6850 66297 6948 66395 4 vdd
rlabel metal3 s 6850 69889 6948 69987 4 vdd
rlabel metal3 s 7282 51287 7380 51385 4 vdd
rlabel metal3 s 6850 88417 6948 88515 4 vdd
rlabel metal3 s 8060 7456 8158 7554 4 vdd
rlabel metal3 s 8060 97516 8158 97614 4 vdd
rlabel metal3 s 7282 75419 7380 75517 4 vdd
rlabel metal3 s 7282 25217 7380 25315 4 vdd
rlabel metal3 s 8060 57621 8158 57719 4 vdd
rlabel metal3 s 7282 15379 7380 15477 4 vdd
rlabel metal3 s 6850 21267 6948 21365 4 vdd
rlabel metal3 s 6850 17317 6948 17415 4 vdd
rlabel metal3 s 7282 71037 7380 71135 4 vdd
rlabel metal3 s 6850 13799 6948 13897 4 vdd
rlabel metal3 s 7282 70247 7380 70345 4 vdd
rlabel metal3 s 6850 72617 6948 72715 4 vdd
rlabel metal3 s 6850 76999 6948 77097 4 vdd
rlabel metal3 s 7282 31537 7380 31635 4 vdd
rlabel metal3 s 6850 99477 6948 99575 4 vdd
rlabel metal3 s 6850 88059 6948 88157 4 vdd
rlabel metal3 s 8060 69076 8158 69174 4 vdd
rlabel metal3 s 7282 56817 7380 56915 4 vdd
rlabel metal3 s 8060 78161 8158 78259 4 vdd
rlabel metal3 s 7282 65507 7380 65605 4 vdd
rlabel metal3 s 8060 79346 8158 79444 4 vdd
rlabel metal3 s 6850 54089 6948 54187 4 vdd
rlabel metal3 s 8060 87246 8158 87344 4 vdd
rlabel metal3 s 7282 92799 7380 92897 4 vdd
rlabel metal3 s 8060 21281 8158 21379 4 vdd
rlabel metal3 s 6850 65149 6948 65247 4 vdd
rlabel metal3 s 7282 21699 7380 21797 4 vdd
rlabel metal3 s 8060 30761 8158 30859 4 vdd
rlabel metal3 s 7282 60409 7380 60507 4 vdd
rlabel metal3 s 7282 39869 7380 39967 4 vdd
rlabel metal3 s 7282 76209 7380 76307 4 vdd
rlabel metal3 s 7282 90429 7380 90527 4 vdd
rlabel metal3 s 6850 64359 6948 64457 4 vdd
rlabel metal3 s 7282 80517 7380 80615 4 vdd
rlabel metal3 s 6850 99909 6948 100007 4 vdd
rlabel metal3 s 7282 78937 7380 79035 4 vdd
rlabel metal3 s 6850 1159 6948 1257 4 vdd
rlabel metal3 s 6850 23637 6948 23735 4 vdd
rlabel metal3 s 7282 26007 7380 26105 4 vdd
rlabel metal3 s 7282 3097 7380 3195 4 vdd
rlabel metal3 s 4326 5086 4424 5184 4 vdd
rlabel metal3 s 8060 95146 8158 95244 4 vdd
rlabel metal3 s 7282 40227 7380 40325 4 vdd
rlabel metal3 s 6850 35129 6948 35227 4 vdd
rlabel metal3 s 8060 32736 8158 32834 4 vdd
rlabel metal3 s 8060 74606 8158 74704 4 vdd
rlabel metal3 s 6850 57249 6948 57347 4 vdd
rlabel metal3 s 7282 46547 7380 46645 4 vdd
rlabel metal3 s 6850 28377 6948 28475 4 vdd
rlabel metal3 s 7282 52509 7380 52607 4 vdd
rlabel metal3 s 8060 49326 8158 49424 4 vdd
rlabel metal3 s 6850 34697 6948 34795 4 vdd
rlabel metal3 s 6850 58829 6948 58927 4 vdd
rlabel metal3 s 7282 68667 7380 68765 4 vdd
rlabel metal3 s 8060 20491 8158 20589 4 vdd
rlabel metal3 s 6850 29599 6948 29697 4 vdd
rlabel metal3 s 6850 8269 6948 8367 4 vdd
rlabel metal3 s 8060 47746 8158 47844 4 vdd
rlabel metal3 s 6850 52509 6948 52607 4 vdd
rlabel metal3 s 6850 66729 6948 66827 4 vdd
rlabel metal3 s 7282 86047 7380 86145 4 vdd
rlabel metal3 s 6850 61199 6948 61297 4 vdd
rlabel metal3 s 8060 88826 8158 88924 4 vdd
rlabel metal3 s 8060 14171 8158 14269 4 vdd
rlabel metal3 s 8060 20886 8158 20984 4 vdd
rlabel metal3 s 6850 94379 6948 94477 4 vdd
rlabel metal3 s 7282 32759 7380 32857 4 vdd
rlabel metal3 s 3116 4319 3214 4417 4 vdd
rlabel metal3 s 8060 3901 8158 3999 4 vdd
rlabel metal3 s 6850 7047 6948 7145 4 vdd
rlabel metal3 s 8060 38661 8158 38759 4 vdd
rlabel metal3 s 7282 54089 7380 54187 4 vdd
rlabel metal3 s 8060 22861 8158 22959 4 vdd
rlabel metal3 s 8060 77766 8158 77864 4 vdd
rlabel metal3 s 7282 95959 7380 96057 4 vdd
rlabel metal3 s 6850 26797 6948 26895 4 vdd
rlabel metal3 s 7282 48917 7380 49015 4 vdd
rlabel metal3 s 1632 6666 1730 6764 4 vdd
rlabel metal3 s 8060 5481 8158 5579 4 vdd
rlabel metal3 s 3116 2739 3214 2837 4 vdd
rlabel metal3 s 3116 9059 3214 9157 4 vdd
rlabel metal3 s 7282 24069 7380 24167 4 vdd
rlabel metal3 s 7282 15737 7380 15835 4 vdd
rlabel metal3 s 6850 89639 6948 89737 4 vdd
rlabel metal3 s 6850 93947 6948 94045 4 vdd
rlabel metal3 s 8060 63941 8158 64039 4 vdd
rlabel metal3 s 6850 83319 6948 83417 4 vdd
rlabel metal3 s 7282 59187 7380 59285 4 vdd
rlabel metal3 s 6850 369 6948 467 4 vdd
rlabel metal3 s 6850 36709 6948 36807 4 vdd
rlabel metal3 s 7282 88059 7380 88157 4 vdd
rlabel metal3 s 6850 18897 6948 18995 4 vdd
rlabel metal3 s 3551 1143 3649 1241 4 vdd
rlabel metal3 s 8060 51696 8158 51794 4 vdd
rlabel metal3 s 7282 38289 7380 38387 4 vdd
rlabel metal3 s 6850 15737 6948 15835 4 vdd
rlabel metal3 s 7282 36709 7380 36807 4 vdd
rlabel metal3 s 8060 31946 8158 32044 4 vdd
rlabel metal3 s 6850 28809 6948 28907 4 vdd
rlabel metal3 s 3116 8269 3214 8367 4 vdd
rlabel metal3 s 7282 69889 7380 69987 4 vdd
rlabel metal3 s 8060 13776 8158 13874 4 vdd
rlabel metal3 s 6850 96317 6948 96415 4 vdd
rlabel metal3 s 7282 13367 7380 13465 4 vdd
rlabel metal3 s 7282 37067 7380 37165 4 vdd
rlabel metal3 s 8060 31551 8158 31649 4 vdd
rlabel metal3 s 6850 100267 6948 100365 4 vdd
rlabel metal3 s 6850 37857 6948 37955 4 vdd
rlabel metal3 s 6850 53299 6948 53397 4 vdd
rlabel metal3 s 8060 35106 8158 35204 4 vdd
rlabel metal3 s 8060 61571 8158 61669 4 vdd
rlabel metal3 s 7282 21267 7380 21365 4 vdd
rlabel metal3 s 6850 19329 6948 19427 4 vdd
rlabel metal3 s 7282 74197 7380 74295 4 vdd
rlabel metal3 s 8060 70656 8158 70754 4 vdd
rlabel metal3 s 8060 72236 8158 72334 4 vdd
rlabel metal3 s 6850 43029 6948 43127 4 vdd
rlabel metal3 s 6850 3097 6948 3195 4 vdd
rlabel metal3 s 6850 47337 6948 47435 4 vdd
rlabel metal3 s 8060 50906 8158 51004 4 vdd
rlabel metal3 s 8060 95541 8158 95639 4 vdd
rlabel metal3 s 7282 39437 7380 39535 4 vdd
rlabel metal3 s 7282 11787 7380 11885 4 vdd
rlabel metal3 s 8060 71051 8158 71149 4 vdd
rlabel metal3 s 7282 17317 7380 17415 4 vdd
rlabel metal3 s 6850 33117 6948 33215 4 vdd
rlabel metal3 s 8060 29971 8158 30069 4 vdd
rlabel metal3 s 7282 76999 7380 77097 4 vdd
rlabel metal3 s 7282 80159 7380 80257 4 vdd
rlabel metal3 s 1632 2716 1730 2814 4 vdd
rlabel metal3 s 8060 91196 8158 91294 4 vdd
rlabel metal3 s 6850 35919 6948 36017 4 vdd
rlabel metal3 s 6850 84899 6948 84997 4 vdd
rlabel metal3 s 7282 66729 7380 66827 4 vdd
rlabel metal3 s 7282 35919 7380 36017 4 vdd
rlabel metal3 s 8060 11011 8158 11109 4 vdd
rlabel metal3 s 8060 27206 8158 27304 4 vdd
rlabel metal3 s 7282 78579 7380 78677 4 vdd
rlabel metal3 s 8060 21676 8158 21774 4 vdd
rlabel metal3 s 8060 2716 8158 2814 4 vdd
rlabel metal3 s 6850 67519 6948 67617 4 vdd
rlabel metal3 s 8060 18911 8158 19009 4 vdd
rlabel metal3 s 8060 48536 8158 48634 4 vdd
rlabel metal3 s 7282 86479 7380 86577 4 vdd
rlabel metal3 s 8060 25626 8158 25724 4 vdd
rlabel metal3 s 6850 38647 6948 38745 4 vdd
rlabel metal3 s 7282 39079 7380 39177 4 vdd
rlabel metal3 s 6850 39437 6948 39535 4 vdd
rlabel metal3 s 6850 50929 6948 51027 4 vdd
rlabel metal3 s 6850 25217 6948 25315 4 vdd
rlabel metal3 s 7282 33907 7380 34005 4 vdd
rlabel metal3 s 7282 38647 7380 38745 4 vdd
rlabel metal3 s 7282 26439 7380 26537 4 vdd
rlabel metal3 s 6850 29957 6948 30055 4 vdd
rlabel metal3 s 8060 59991 8158 60089 4 vdd
rlabel metal3 s 6850 70679 6948 70777 4 vdd
rlabel metal3 s 7282 5899 7380 5997 4 vdd
rlabel metal3 s 8060 77371 8158 77469 4 vdd
rlabel metal3 s 8060 80136 8158 80234 4 vdd
rlabel metal3 s 6850 43819 6948 43917 4 vdd
rlabel metal3 s 7282 7047 7380 7145 4 vdd
rlabel metal3 s 4326 4296 4424 4394 4 vdd
rlabel metal3 s 8060 8641 8158 8739 4 vdd
rlabel metal3 s 8060 84876 8158 84974 4 vdd
rlabel metal3 s 6850 72259 6948 72357 4 vdd
rlabel metal3 s 8060 82506 8158 82604 4 vdd
rlabel metal3 s 8060 99491 8158 99589 4 vdd
rlabel metal3 s 8060 15751 8158 15849 4 vdd
rlabel metal3 s 8060 28786 8158 28884 4 vdd
rlabel metal3 s 6850 73407 6948 73505 4 vdd
rlabel metal3 s 6850 97897 6948 97995 4 vdd
rlabel metal3 s 7282 10997 7380 11095 4 vdd
rlabel metal3 s 6850 20909 6948 21007 4 vdd
rlabel metal3 s 7282 93947 7380 94045 4 vdd
rlabel metal3 s 6850 41017 6948 41115 4 vdd
rlabel metal3 s 8060 88036 8158 88134 4 vdd
rlabel metal3 s 8060 86456 8158 86554 4 vdd
rlabel metal3 s 8060 29576 8158 29674 4 vdd
rlabel metal3 s 8060 33526 8158 33624 4 vdd
rlabel metal3 s 7282 33117 7380 33215 4 vdd
rlabel metal3 s 8060 59201 8158 59299 4 vdd
rlabel metal3 s 8060 44191 8158 44289 4 vdd
rlabel metal3 s 8060 93961 8158 94059 4 vdd
rlabel metal3 s 7282 75777 7380 75875 4 vdd
rlabel metal3 s 8060 34711 8158 34809 4 vdd
rlabel metal3 s 8060 87641 8158 87739 4 vdd
rlabel metal3 s 4326 346 4424 444 4 vdd
rlabel metal3 s 8060 96726 8158 96824 4 vdd
rlabel metal3 s 6850 56459 6948 56557 4 vdd
rlabel metal3 s 4326 2716 4424 2814 4 vdd
rlabel metal3 s 8060 67101 8158 67199 4 vdd
rlabel metal3 s 7282 80949 7380 81047 4 vdd
rlabel metal3 s 8060 97121 8158 97219 4 vdd
rlabel metal3 s 8060 56041 8158 56139 4 vdd
rlabel metal3 s 7282 58829 7380 58927 4 vdd
rlabel metal3 s 7282 69099 7380 69197 4 vdd
rlabel metal3 s 6850 53657 6948 53755 4 vdd
rlabel metal3 s 6850 46979 6948 47077 4 vdd
rlabel metal3 s 6850 78147 6948 78245 4 vdd
rlabel metal3 s 6850 85257 6948 85355 4 vdd
rlabel metal3 s 8060 44586 8158 44684 4 vdd
rlabel metal3 s 8060 88431 8158 88529 4 vdd
rlabel metal3 s 8060 30366 8158 30464 4 vdd
rlabel metal3 s 6850 64717 6948 64815 4 vdd
rlabel metal3 s 7282 68309 7380 68407 4 vdd
rlabel metal3 s 6850 38289 6948 38387 4 vdd
rlabel metal3 s 8060 89616 8158 89714 4 vdd
rlabel metal3 s 6850 96749 6948 96847 4 vdd
rlabel metal3 s 8060 48931 8158 49029 4 vdd
rlabel metal3 s 7282 28019 7380 28117 4 vdd
rlabel metal3 s 6850 84109 6948 84207 4 vdd
rlabel metal3 s 8060 34316 8158 34414 4 vdd
rlabel metal3 s 7282 93589 7380 93687 4 vdd
rlabel metal3 s 8060 97911 8158 98009 4 vdd
rlabel metal3 s 7282 31969 7380 32067 4 vdd
rlabel metal3 s 7282 36277 7380 36375 4 vdd
rlabel metal3 s 6850 6689 6948 6787 4 vdd
rlabel metal3 s 6850 78579 6948 78677 4 vdd
rlabel metal3 s 6850 16959 6948 17057 4 vdd
rlabel metal3 s 7282 89207 7380 89305 4 vdd
rlabel metal3 s 8060 100281 8158 100379 4 vdd
rlabel metal3 s 7282 16959 7380 17057 4 vdd
rlabel metal3 s 8060 45376 8158 45474 4 vdd
rlabel metal3 s 6850 2739 6948 2837 4 vdd
rlabel metal3 s 7282 35129 7380 35227 4 vdd
rlabel metal3 s 6850 10207 6948 10305 4 vdd
rlabel metal3 s 8060 68681 8158 68779 4 vdd
rlabel metal3 s 7282 28809 7380 28907 4 vdd
rlabel metal3 s 8060 18516 8158 18614 4 vdd
rlabel metal3 s 8060 79741 8158 79839 4 vdd
rlabel metal3 s 8060 71446 8158 71544 4 vdd
rlabel metal3 s 7282 82887 7380 82985 4 vdd
rlabel metal3 s 8060 37476 8158 37574 4 vdd
rlabel metal3 s 8060 36291 8158 36389 4 vdd
rlabel metal3 s 8060 47351 8158 47449 4 vdd
rlabel metal3 s 4326 6666 4424 6764 4 vdd
rlabel metal3 s 6850 80949 6948 81047 4 vdd
rlabel metal3 s 6850 7837 6948 7935 4 vdd
rlabel metal3 s 6850 57607 6948 57705 4 vdd
rlabel metal3 s 7282 60767 7380 60865 4 vdd
rlabel metal3 s 7282 66297 7380 66395 4 vdd
rlabel metal3 s 8060 50116 8158 50214 4 vdd
rlabel metal3 s 3116 3529 3214 3627 4 vdd
rlabel metal3 s 8060 83296 8158 83394 4 vdd
rlabel metal3 s 7282 44177 7380 44275 4 vdd
rlabel metal3 s 6850 39079 6948 39177 4 vdd
rlabel metal3 s 8060 61966 8158 62064 4 vdd
rlabel metal3 s 6850 90787 6948 90885 4 vdd
rlabel metal3 s 8060 40636 8158 40734 4 vdd
rlabel metal3 s 6850 5899 6948 5997 4 vdd
rlabel metal3 s 8060 64731 8158 64829 4 vdd
rlabel metal3 s 8060 98701 8158 98799 4 vdd
rlabel metal3 s 4326 1136 4424 1234 4 vdd
rlabel metal3 s 7282 3529 7380 3627 4 vdd
rlabel metal3 s 6850 56027 6948 56125 4 vdd
rlabel metal3 s 7282 81307 7380 81405 4 vdd
rlabel metal3 s 3548 4319 3646 4417 4 vdd
rlabel metal3 s 8060 43796 8158 43894 4 vdd
rlabel metal3 s 6850 14157 6948 14255 4 vdd
rlabel metal3 s 6850 79727 6948 79825 4 vdd
rlabel metal3 s 8060 85271 8158 85369 4 vdd
rlabel metal3 s 7282 73839 7380 73937 4 vdd
rlabel metal3 s 6850 75777 6948 75875 4 vdd
rlabel metal3 s 6850 49707 6948 49805 4 vdd
rlabel metal3 s 8060 64336 8158 64434 4 vdd
rlabel metal3 s 6850 20119 6948 20217 4 vdd
rlabel metal3 s 7282 11429 7380 11527 4 vdd
rlabel metal3 s 6850 98329 6948 98427 4 vdd
rlabel metal3 s 8060 6271 8158 6369 4 vdd
rlabel metal3 s 6850 59187 6948 59285 4 vdd
rlabel metal3 s 6850 31537 6948 31635 4 vdd
rlabel metal3 s 6850 36277 6948 36375 4 vdd
rlabel metal3 s 8060 76581 8158 76679 4 vdd
rlabel metal3 s 8060 7851 8158 7949 4 vdd
rlabel metal3 s 7282 56459 7380 56557 4 vdd
rlabel metal3 s 7282 55237 7380 55335 4 vdd
rlabel metal3 s 6850 6257 6948 6355 4 vdd
rlabel metal3 s 8060 3111 8158 3209 4 vdd
rlabel metal3 s 6850 67087 6948 67185 4 vdd
rlabel metal3 s 8060 73421 8158 73519 4 vdd
rlabel metal3 s 6850 42597 6948 42695 4 vdd
rlabel metal3 s 6850 41807 6948 41905 4 vdd
rlabel metal3 s 6850 25649 6948 25747 4 vdd
rlabel metal3 s 7282 52077 7380 52175 4 vdd
rlabel metal3 s 7282 94379 7380 94477 4 vdd
rlabel metal3 s 8060 43401 8158 43499 4 vdd
rlabel metal3 s 8060 94356 8158 94454 4 vdd
rlabel metal3 s 8060 86061 8158 86159 4 vdd
rlabel metal3 s 7282 61557 7380 61655 4 vdd
rlabel metal3 s 8060 9431 8158 9529 4 vdd
rlabel metal3 s 8060 4296 8158 4394 4 vdd
rlabel metal3 s 7282 65939 7380 66037 4 vdd
rlabel metal3 s 6850 76209 6948 76307 4 vdd
rlabel metal3 s 8060 65126 8158 65224 4 vdd
rlabel metal3 s 7282 54447 7380 54545 4 vdd
rlabel metal3 s 7282 95527 7380 95625 4 vdd
rlabel metal3 s 2228 346 2326 444 4 vdd
rlabel metal3 s 8060 16541 8158 16639 4 vdd
rlabel metal3 s 7282 46979 7380 47077 4 vdd
rlabel metal3 s 8060 40241 8158 40339 4 vdd
rlabel metal3 s 8060 60386 8158 60484 4 vdd
rlabel metal3 s 7282 23637 7380 23735 4 vdd
rlabel metal3 s 7282 84109 7380 84207 4 vdd
rlabel metal3 s 8060 90801 8158 90899 4 vdd
rlabel metal3 s 7282 30389 7380 30487 4 vdd
rlabel metal3 s 7282 18107 7380 18205 4 vdd
rlabel metal3 s 8060 5086 8158 5184 4 vdd
rlabel metal3 s 6850 93589 6948 93687 4 vdd
rlabel metal3 s 8060 53671 8158 53769 4 vdd
rlabel metal3 s 6850 43387 6948 43485 4 vdd
rlabel metal3 s 6850 9849 6948 9947 4 vdd
rlabel metal3 s 6850 24859 6948 24957 4 vdd
rlabel metal3 s 8060 76976 8158 77074 4 vdd
rlabel metal3 s 8060 73816 8158 73914 4 vdd
rlabel metal3 s 7282 88849 7380 88947 4 vdd
rlabel metal3 s 6850 93157 6948 93255 4 vdd
rlabel metal3 s 3548 6689 3646 6787 4 vdd
rlabel metal3 s 8060 24836 8158 24934 4 vdd
rlabel metal3 s 7282 95169 7380 95267 4 vdd
rlabel metal3 s 6850 65939 6948 66037 4 vdd
rlabel metal3 s 7282 79727 7380 79825 4 vdd
rlabel metal3 s 7282 81739 7380 81837 4 vdd
rlabel metal3 s 7282 77357 7380 77455 4 vdd
rlabel metal3 s 6850 8627 6948 8725 4 vdd
rlabel metal3 s 6850 95527 6948 95625 4 vdd
rlabel metal3 s 7282 57607 7380 57705 4 vdd
rlabel metal3 s 8060 93566 8158 93664 4 vdd
rlabel metal3 s 6850 37067 6948 37165 4 vdd
rlabel metal3 s 6850 94737 6948 94835 4 vdd
rlabel metal3 s 8060 19701 8158 19799 4 vdd
rlabel metal3 s 7282 59977 7380 60075 4 vdd
rlabel metal3 s 8060 63546 8158 63644 4 vdd
rlabel metal3 s 8060 46956 8158 47054 4 vdd
rlabel metal3 s 3548 2739 3646 2837 4 vdd
rlabel metal3 s 7282 46189 7380 46287 4 vdd
rlabel metal3 s 8060 12196 8158 12294 4 vdd
rlabel metal3 s 6850 92799 6948 92897 4 vdd
rlabel metal3 s 8060 48141 8158 48239 4 vdd
rlabel metal3 s 8060 16146 8158 16244 4 vdd
rlabel metal3 s 7282 94737 7380 94835 4 vdd
rlabel metal3 s 8060 18121 8158 18219 4 vdd
rlabel metal3 s 6850 2307 6948 2405 4 vdd
rlabel metal3 s 8060 42216 8158 42314 4 vdd
rlabel metal3 s 7282 56027 7380 56125 4 vdd
rlabel metal3 s 7282 86837 7380 86935 4 vdd
rlabel metal3 s 6850 78937 6948 79035 4 vdd
rlabel metal3 s 7282 49349 7380 49447 4 vdd
rlabel metal3 s 8060 91591 8158 91689 4 vdd
rlabel metal3 s 8060 53276 8158 53374 4 vdd
rlabel metal3 s 7282 64359 7380 64457 4 vdd
rlabel metal3 s 7282 99909 7380 100007 4 vdd
rlabel metal3 s 6850 69099 6948 69197 4 vdd
rlabel metal3 s 7282 22847 7380 22945 4 vdd
rlabel metal3 s 8060 66706 8158 66804 4 vdd
rlabel metal3 s 7282 3887 7380 3985 4 vdd
rlabel metal3 s 8060 50511 8158 50609 4 vdd
rlabel metal3 s 6850 74987 6948 75085 4 vdd
rlabel metal3 s 7282 50139 7380 50237 4 vdd
rlabel metal3 s 8060 6666 8158 6764 4 vdd
rlabel metal3 s 6850 67877 6948 67975 4 vdd
rlabel metal3 s 6850 20477 6948 20575 4 vdd
rlabel metal3 s 7282 9417 7380 9515 4 vdd
rlabel metal3 s 7282 16169 7380 16267 4 vdd
rlabel metal3 s 7282 70679 7380 70777 4 vdd
rlabel metal3 s 8060 41821 8158 41919 4 vdd
rlabel metal3 s 6850 3529 6948 3627 4 vdd
rlabel metal3 s 7282 8269 7380 8367 4 vdd
rlabel metal3 s 8060 31156 8158 31254 4 vdd
rlabel metal3 s 6850 44177 6948 44275 4 vdd
rlabel metal3 s 6850 48127 6948 48225 4 vdd
rlabel metal3 s 6850 44967 6948 45065 4 vdd
rlabel metal3 s 8060 65521 8158 65619 4 vdd
rlabel metal3 s 7282 19329 7380 19427 4 vdd
rlabel metal3 s 7282 87627 7380 87725 4 vdd
rlabel metal3 s 6850 68309 6948 68407 4 vdd
rlabel metal3 s 8060 38266 8158 38364 4 vdd
rlabel metal3 s 6850 12219 6948 12317 4 vdd
rlabel metal3 s 6850 37499 6948 37597 4 vdd
rlabel metal3 s 7282 58039 7380 58137 4 vdd
rlabel metal3 s 8060 37081 8158 37179 4 vdd
rlabel metal3 s 8060 99096 8158 99194 4 vdd
rlabel metal3 s 8060 70261 8158 70359 4 vdd
rlabel metal3 s 3548 5109 3646 5207 4 vdd
rlabel metal3 s 7282 4677 7380 4775 4 vdd
rlabel metal3 s 7282 90787 7380 90885 4 vdd
rlabel metal3 s 6850 23279 6948 23377 4 vdd
rlabel metal3 s 8060 92776 8158 92874 4 vdd
rlabel metal3 s 8060 3506 8158 3604 4 vdd
rlabel metal3 s 7282 1949 7380 2047 4 vdd
rlabel metal3 s 7282 25649 7380 25747 4 vdd
rlabel metal3 s 8060 42611 8158 42709 4 vdd
rlabel metal3 s 8060 60781 8158 60879 4 vdd
rlabel metal3 s 6850 79369 6948 79467 4 vdd
rlabel metal3 s 6850 18539 6948 18637 4 vdd
rlabel metal3 s 8060 20096 8158 20194 4 vdd
rlabel metal3 s 6850 81307 6948 81405 4 vdd
rlabel metal3 s 8060 25231 8158 25329 4 vdd
rlabel metal3 s 8060 100676 8158 100774 4 vdd
rlabel metal3 s 6850 45757 6948 45855 4 vdd
rlabel metal3 s 6850 52077 6948 52175 4 vdd
rlabel metal3 s 6850 61557 6948 61655 4 vdd
rlabel metal3 s 6850 7479 6948 7577 4 vdd
rlabel metal3 s 6850 62779 6948 62877 4 vdd
rlabel metal3 s 6850 70247 6948 70345 4 vdd
rlabel metal3 s 8060 10616 8158 10714 4 vdd
rlabel metal3 s 7282 91577 7380 91675 4 vdd
rlabel metal3 s 8060 94751 8158 94849 4 vdd
rlabel metal3 s 6850 74197 6948 74295 4 vdd
rlabel metal3 s 7282 97107 7380 97205 4 vdd
rlabel metal3 s 7282 24859 7380 24957 4 vdd
rlabel metal3 s 6850 68667 6948 68765 4 vdd
rlabel metal3 s 7282 61989 7380 62087 4 vdd
rlabel metal3 s 8060 41031 8158 41129 4 vdd
rlabel metal3 s 7282 50929 7380 51027 4 vdd
rlabel metal3 s 7282 7837 7380 7935 4 vdd
rlabel metal3 s 8060 23256 8158 23354 4 vdd
rlabel metal3 s 8060 81716 8158 81814 4 vdd
rlabel metal3 s 6850 89207 6948 89305 4 vdd
rlabel metal3 s 7282 83677 7380 83775 4 vdd
rlabel metal3 s 7282 28377 7380 28475 4 vdd
rlabel metal3 s 6850 69457 6948 69555 4 vdd
rlabel metal3 s 8060 11801 8158 11899 4 vdd
rlabel metal3 s 6850 87627 6948 87725 4 vdd
rlabel metal3 s 7282 92367 7380 92465 4 vdd
rlabel metal3 s 6850 3887 6948 3985 4 vdd
rlabel metal3 s 7282 48127 7380 48225 4 vdd
rlabel metal3 s 7282 62347 7380 62445 4 vdd
rlabel metal3 s 7282 63927 7380 64025 4 vdd
rlabel metal3 s 8060 27601 8158 27699 4 vdd
rlabel metal3 s 8060 741 8158 839 4 vdd
rlabel metal3 s 8060 10221 8158 10319 4 vdd
rlabel metal3 s 7282 7479 7380 7577 4 vdd
rlabel metal3 s 6850 31969 6948 32067 4 vdd
rlabel metal3 s 7282 33549 7380 33647 4 vdd
rlabel metal3 s 6850 24069 6948 24167 4 vdd
rlabel metal3 s 7282 89997 7380 90095 4 vdd
rlabel metal3 s 7282 10639 7380 10737 4 vdd
rlabel metal3 s 7282 67087 7380 67185 4 vdd
rlabel metal3 s 8060 65916 8158 66014 4 vdd
rlabel metal3 s 6850 95169 6948 95267 4 vdd
rlabel metal3 s 6850 28019 6948 28117 4 vdd
rlabel metal3 s 7282 72259 7380 72357 4 vdd
rlabel metal3 s 6850 89997 6948 90095 4 vdd
rlabel metal3 s 7282 14589 7380 14687 4 vdd
rlabel metal3 s 4326 9036 4424 9134 4 vdd
rlabel metal3 s 7282 41449 7380 41547 4 vdd
rlabel metal3 s 6850 59977 6948 60075 4 vdd
rlabel metal3 s 8060 26811 8158 26909 4 vdd
rlabel metal3 s 7282 31179 7380 31277 4 vdd
rlabel metal3 s 7282 58397 7380 58495 4 vdd
rlabel metal3 s 6850 71827 6948 71925 4 vdd
rlabel metal3 s 6850 60409 6948 60507 4 vdd
rlabel metal3 s 7282 78147 7380 78245 4 vdd
rlabel metal3 s 6850 39869 6948 39967 4 vdd
rlabel metal3 s 6850 63927 6948 64025 4 vdd
rlabel metal3 s 8060 4691 8158 4789 4 vdd
rlabel metal3 s 7282 37857 7380 37955 4 vdd
rlabel metal3 s 6850 48559 6948 48657 4 vdd
rlabel metal3 s 8060 56831 8158 56929 4 vdd
rlabel metal3 s 8060 44981 8158 45079 4 vdd
rlabel metal3 s 6850 9417 6948 9515 4 vdd
rlabel metal3 s 7282 727 7380 825 4 vdd
rlabel metal3 s 6850 18107 6948 18205 4 vdd
rlabel metal3 s 7282 63569 7380 63667 4 vdd
rlabel metal3 s 6850 88849 6948 88947 4 vdd
rlabel metal3 s 8060 23651 8158 23749 4 vdd
rlabel metal3 s 7282 54879 7380 54977 4 vdd
rlabel metal3 s 6850 99119 6948 99217 4 vdd
rlabel metal3 s 8060 22466 8158 22564 4 vdd
rlabel metal3 s 6850 24427 6948 24525 4 vdd
rlabel metal3 s 4326 7456 4424 7554 4 vdd
rlabel metal3 s 7282 14947 7380 15045 4 vdd
rlabel metal3 s 7282 29599 7380 29697 4 vdd
rlabel metal3 s 7282 84467 7380 84565 4 vdd
rlabel metal3 s 7282 64717 7380 64815 4 vdd
rlabel metal3 s 7282 23279 7380 23377 4 vdd
rlabel metal3 s 8060 59596 8158 59694 4 vdd
rlabel metal3 s 8060 82901 8158 82999 4 vdd
rlabel metal3 s 6850 29167 6948 29265 4 vdd
rlabel metal3 s 6850 32327 6948 32425 4 vdd
rlabel metal3 s 6850 80517 6948 80615 4 vdd
rlabel metal3 s 6850 5467 6948 5565 4 vdd
rlabel metal3 s 7282 41807 7380 41905 4 vdd
rlabel metal3 s 8060 90011 8158 90109 4 vdd
rlabel metal3 s 7282 6689 7380 6787 4 vdd
rlabel metal3 s 7282 16527 7380 16625 4 vdd
rlabel metal3 s 7282 52867 7380 52965 4 vdd
rlabel metal3 s 6850 27229 6948 27327 4 vdd
rlabel metal3 s 8060 82111 8158 82209 4 vdd
rlabel metal3 s 6850 26007 6948 26105 4 vdd
rlabel metal3 s 6850 91577 6948 91675 4 vdd
rlabel metal3 s 6850 52867 6948 52965 4 vdd
rlabel metal3 s 6850 11429 6948 11527 4 vdd
rlabel metal3 s 8060 11406 8158 11504 4 vdd
rlabel metal3 s 8060 51301 8158 51399 4 vdd
rlabel metal3 s 8060 19306 8158 19404 4 vdd
rlabel metal3 s 8060 35896 8158 35994 4 vdd
rlabel metal3 s 8060 74211 8158 74309 4 vdd
rlabel metal3 s 6850 82887 6948 82985 4 vdd
rlabel metal3 s 8060 22071 8158 22169 4 vdd
rlabel metal3 s 7282 2739 7380 2837 4 vdd
rlabel metal3 s 7282 29957 7380 30055 4 vdd
rlabel metal3 s 7282 13799 7380 13897 4 vdd
rlabel metal3 s 7282 369 7380 467 4 vdd
rlabel metal3 s 7282 41017 7380 41115 4 vdd
rlabel metal3 s 7282 34339 7380 34437 4 vdd
rlabel metal3 s 6850 61989 6948 62087 4 vdd
rlabel metal3 s 7282 67877 7380 67975 4 vdd
rlabel metal3 s 8060 33921 8158 34019 4 vdd
rlabel metal3 s 6850 100699 6948 100797 4 vdd
rlabel metal3 s 3548 3529 3646 3627 4 vdd
rlabel metal3 s 7282 32327 7380 32425 4 vdd
rlabel metal3 s 6850 86837 6948 86935 4 vdd
rlabel metal3 s 8060 9036 8158 9134 4 vdd
rlabel metal3 s 6850 45399 6948 45497 4 vdd
rlabel metal3 s 6850 14947 6948 15045 4 vdd
rlabel metal3 s 7282 5467 7380 5565 4 vdd
rlabel metal3 s 7282 85257 7380 85355 4 vdd
rlabel metal3 s 7282 4319 7380 4417 4 vdd
rlabel metal3 s 6850 81739 6948 81837 4 vdd
rlabel metal3 s 7282 99119 7380 99217 4 vdd
rlabel metal3 s 7282 53299 7380 53397 4 vdd
rlabel metal3 s 8060 78951 8158 79049 4 vdd
rlabel metal3 s 7282 88417 7380 88515 4 vdd
rlabel metal3 s 3551 353 3649 451 4 vdd
rlabel metal3 s 6850 1949 6948 2047 4 vdd
rlabel metal3 s 8060 2321 8158 2419 4 vdd
rlabel metal3 s 8060 99886 8158 99984 4 vdd
rlabel metal3 s 7282 47769 7380 47867 4 vdd
rlabel metal3 s 7282 14157 7380 14255 4 vdd
rlabel metal3 s 8060 15356 8158 15454 4 vdd
rlabel metal3 s 7282 67519 7380 67617 4 vdd
rlabel metal3 s 8060 75001 8158 75099 4 vdd
rlabel metal3 s 8060 12986 8158 13084 4 vdd
rlabel metal3 s 8060 54461 8158 54559 4 vdd
rlabel metal3 s 8060 86851 8158 86949 4 vdd
rlabel metal3 s 7282 96317 7380 96415 4 vdd
rlabel metal3 s 6850 4677 6948 4775 4 vdd
rlabel metal3 s 8060 14566 8158 14664 4 vdd
rlabel metal3 s 6850 50497 6948 50595 4 vdd
rlabel metal3 s 8060 93171 8158 93269 4 vdd
rlabel metal3 s 7282 57249 7380 57347 4 vdd
rlabel metal3 s 8060 49721 8158 49819 4 vdd
rlabel metal3 s 8060 27996 8158 28094 4 vdd
rlabel metal3 s 8060 55646 8158 55744 4 vdd
rlabel metal3 s 6850 33907 6948 34005 4 vdd
rlabel metal3 s 7282 20909 7380 21007 4 vdd
rlabel metal3 s 7282 49707 7380 49805 4 vdd
rlabel metal3 s 7282 18539 7380 18637 4 vdd
rlabel metal3 s 7282 59619 7380 59717 4 vdd
rlabel metal3 s 7282 53657 7380 53755 4 vdd
rlabel metal3 s 6850 14589 6948 14687 4 vdd
rlabel metal3 s 6850 63569 6948 63667 4 vdd
rlabel metal3 s 7282 10207 7380 10305 4 vdd
rlabel metal3 s 6850 97107 6948 97205 4 vdd
rlabel metal3 s 7282 27229 7380 27327 4 vdd
rlabel metal3 s 7282 20477 7380 20575 4 vdd
rlabel metal3 s 6850 63137 6948 63235 4 vdd
rlabel metal3 s 6850 83677 6948 83775 4 vdd
rlabel metal3 s 7282 37499 7380 37597 4 vdd
rlabel metal3 s 7282 29167 7380 29265 4 vdd
rlabel metal3 s 6850 42239 6948 42337 4 vdd
rlabel metal3 s 8060 33131 8158 33229 4 vdd
rlabel metal3 s 6850 33549 6948 33647 4 vdd
rlabel metal3 s 7282 73407 7380 73505 4 vdd
rlabel metal3 s 6850 73839 6948 73937 4 vdd
rlabel metal3 s 8060 52881 8158 52979 4 vdd
rlabel metal3 s 8060 7061 8158 7159 4 vdd
rlabel metal3 s 8060 13381 8158 13479 4 vdd
rlabel metal3 s 6850 59619 6948 59717 4 vdd
rlabel metal3 s 7282 27587 7380 27685 4 vdd
rlabel metal3 s 7282 82529 7380 82627 4 vdd
rlabel metal3 s 7282 19687 7380 19785 4 vdd
rlabel metal3 s 7282 55669 7380 55767 4 vdd
rlabel metal3 s 6850 13009 6948 13107 4 vdd
rlabel metal3 s 7282 44967 7380 45065 4 vdd
rlabel metal3 s 7282 40659 7380 40757 4 vdd
rlabel metal3 s 8060 39846 8158 39944 4 vdd
rlabel metal3 s 6850 98687 6948 98785 4 vdd
rlabel metal3 s 6850 27587 6948 27685 4 vdd
rlabel metal3 s 8060 26021 8158 26119 4 vdd
rlabel metal3 s 7282 44609 7380 44707 4 vdd
rlabel metal3 s 7282 51719 7380 51817 4 vdd
rlabel metal3 s 7282 42239 7380 42337 4 vdd
rlabel metal3 s 6850 65507 6948 65605 4 vdd
rlabel metal3 s 7282 84899 7380 84997 4 vdd
rlabel metal3 s 8060 95936 8158 96034 4 vdd
rlabel metal3 s 8060 17331 8158 17429 4 vdd
rlabel metal3 s 6850 22057 6948 22155 4 vdd
rlabel metal3 s 6850 77357 6948 77455 4 vdd
rlabel metal3 s 7282 17749 7380 17847 4 vdd
rlabel metal3 s 8060 67891 8158 67989 4 vdd
rlabel metal3 s 8060 8246 8158 8344 4 vdd
rlabel metal3 s 8060 76186 8158 76284 4 vdd
rlabel metal3 s 8060 24046 8158 24144 4 vdd
rlabel metal3 s 8060 84481 8158 84579 4 vdd
rlabel metal3 s 6850 86479 6948 86577 4 vdd
rlabel metal3 s 6850 727 6948 825 4 vdd
rlabel metal3 s 6850 48917 6948 49015 4 vdd
rlabel metal3 s 8060 29181 8158 29279 4 vdd
rlabel metal3 s 8060 54856 8158 54954 4 vdd
rlabel metal3 s 8060 43006 8158 43104 4 vdd
rlabel metal3 s 8060 83691 8158 83789 4 vdd
rlabel metal3 s 8060 69471 8158 69569 4 vdd
rlabel metal3 s 7282 65149 7380 65247 4 vdd
rlabel metal3 s 6850 17749 6948 17847 4 vdd
rlabel metal3 s 7282 50497 7380 50595 4 vdd
rlabel metal3 s 6850 16169 6948 16267 4 vdd
rlabel metal3 s 6850 15379 6948 15477 4 vdd
rlabel metal3 s 8060 66311 8158 66409 4 vdd
rlabel metal3 s 7282 97897 7380 97995 4 vdd
rlabel metal3 s 7282 74629 7380 74727 4 vdd
rlabel metal3 s 8060 28391 8158 28489 4 vdd
rlabel metal3 s 7282 45757 7380 45855 4 vdd
rlabel metal3 s 8060 80926 8158 81024 4 vdd
rlabel metal3 s 6850 10639 6948 10737 4 vdd
rlabel metal3 s 6850 40227 6948 40325 4 vdd
rlabel metal3 s 8060 75396 8158 75494 4 vdd
rlabel metal3 s 6850 74629 6948 74727 4 vdd
rlabel metal3 s 8060 92381 8158 92479 4 vdd
rlabel metal3 s 6850 30747 6948 30845 4 vdd
rlabel metal3 s 6850 73049 6948 73147 4 vdd
rlabel metal3 s 8060 62756 8158 62854 4 vdd
rlabel metal3 s 8060 39451 8158 39549 4 vdd
rlabel metal3 s 6850 47769 6948 47867 4 vdd
rlabel metal3 s 7282 93157 7380 93255 4 vdd
rlabel metal3 s 7282 22057 7380 22155 4 vdd
rlabel metal3 s 8060 26416 8158 26514 4 vdd
rlabel metal3 s 6850 30389 6948 30487 4 vdd
rlabel metal3 s 6850 12577 6948 12675 4 vdd
rlabel metal3 s 6850 84467 6948 84565 4 vdd
rlabel metal3 s 6850 87269 6948 87367 4 vdd
rlabel metal3 s 6850 82097 6948 82195 4 vdd
rlabel metal3 s 8060 12591 8158 12689 4 vdd
rlabel metal3 s 8060 67496 8158 67594 4 vdd
rlabel metal3 s 7282 69457 7380 69555 4 vdd
rlabel metal3 s 7282 43029 7380 43127 4 vdd
rlabel metal3 s 6850 41449 6948 41547 4 vdd
rlabel metal3 s 7282 63137 7380 63235 4 vdd
rlabel metal3 s 6850 82529 6948 82627 4 vdd
rlabel metal3 s 8060 1136 8158 1234 4 vdd
rlabel metal3 s 8060 72631 8158 72729 4 vdd
rlabel metal3 s 6850 26439 6948 26537 4 vdd
rlabel metal3 s 7282 100699 7380 100797 4 vdd
rlabel metal3 s 7664 82111 7762 82209 4 gnd
rlabel metal3 s 6425 56085 6523 56183 4 gnd
rlabel metal3 s 6425 16169 6523 16267 4 gnd
rlabel metal3 s 7664 35896 7762 35994 4 gnd
rlabel metal3 s 6425 21699 6523 21797 4 gnd
rlabel metal3 s 7664 43401 7762 43499 4 gnd
rlabel metal3 s 6425 92799 6523 92897 4 gnd
rlabel metal3 s 6425 89639 6523 89737 4 gnd
rlabel metal3 s 6425 34755 6523 34853 4 gnd
rlabel metal3 s 6425 71885 6523 71983 4 gnd
rlabel metal3 s 7664 57226 7762 57324 4 gnd
rlabel metal3 s 7664 45771 7762 45869 4 gnd
rlabel metal3 s 6425 47769 6523 47867 4 gnd
rlabel metal3 s 7664 59991 7762 60089 4 gnd
rlabel metal3 s 6425 49349 6523 49447 4 gnd
rlabel metal3 s 6425 8685 6523 8783 4 gnd
rlabel metal3 s 7664 61176 7762 61274 4 gnd
rlabel metal3 s 6425 10265 6523 10363 4 gnd
rlabel metal3 s 7664 85666 7762 85764 4 gnd
rlabel metal3 s 6425 97165 6523 97263 4 gnd
rlabel metal3 s 6425 58455 6523 58553 4 gnd
rlabel metal3 s 6425 97539 6523 97637 4 gnd
rlabel metal3 s 6425 100325 6523 100423 4 gnd
rlabel metal3 s 6425 5525 6523 5623 4 gnd
rlabel metal3 s 6425 24859 6523 24957 4 gnd
rlabel metal3 s 7664 61966 7762 62064 4 gnd
rlabel metal3 s 6425 2739 6523 2837 4 gnd
rlabel metal3 s 7664 29181 7762 29279 4 gnd
rlabel metal3 s 6425 33175 6523 33273 4 gnd
rlabel metal3 s 7664 49326 7762 49424 4 gnd
rlabel metal3 s 6425 70305 6523 70403 4 gnd
rlabel metal3 s 6425 77415 6523 77513 4 gnd
rlabel metal3 s 6425 3155 6523 3253 4 gnd
rlabel metal3 s 7664 30761 7762 30859 4 gnd
rlabel metal3 s 6425 70679 6523 70777 4 gnd
rlabel metal3 s 2691 7479 2789 7577 4 gnd
rlabel metal3 s 6425 2365 6523 2463 4 gnd
rlabel metal3 s 6425 28435 6523 28533 4 gnd
rlabel metal3 s 6425 38289 6523 38387 4 gnd
rlabel metal3 s 6425 42655 6523 42753 4 gnd
rlabel metal3 s 7664 42611 7762 42709 4 gnd
rlabel metal3 s 7664 8641 7762 8739 4 gnd
rlabel metal3 s 6425 14215 6523 14313 4 gnd
rlabel metal3 s 6425 9475 6523 9573 4 gnd
rlabel metal3 s 6425 53715 6523 53813 4 gnd
rlabel metal3 s 6425 39495 6523 39593 4 gnd
rlabel metal3 s 7664 86061 7762 86159 4 gnd
rlabel metal3 s 6425 46189 6523 46287 4 gnd
rlabel metal3 s 7664 50511 7762 50609 4 gnd
rlabel metal3 s 6425 7105 6523 7203 4 gnd
rlabel metal3 s 6425 4735 6523 4833 4 gnd
rlabel metal3 s 7664 81716 7762 81814 4 gnd
rlabel metal3 s 6425 84525 6523 84623 4 gnd
rlabel metal3 s 6425 35129 6523 35227 4 gnd
rlabel metal3 s 7664 91591 7762 91689 4 gnd
rlabel metal3 s 6425 19745 6523 19843 4 gnd
rlabel metal3 s 6425 43029 6523 43127 4 gnd
rlabel metal3 s 6425 65149 6523 65247 4 gnd
rlabel metal3 s 7664 32341 7762 32439 4 gnd
rlabel metal3 s 7664 63151 7762 63249 4 gnd
rlabel metal3 s 6425 79369 6523 79467 4 gnd
rlabel metal3 s 7664 18121 7762 18219 4 gnd
rlabel metal3 s 7664 69076 7762 69174 4 gnd
rlabel metal3 s 7664 26021 7762 26119 4 gnd
rlabel metal3 s 7664 28391 7762 28489 4 gnd
rlabel metal3 s 7664 65916 7762 66014 4 gnd
rlabel metal3 s 7664 83691 7762 83789 4 gnd
rlabel metal3 s 7664 66311 7762 66409 4 gnd
rlabel metal3 s 6425 22115 6523 22213 4 gnd
rlabel metal3 s 7664 52091 7762 52189 4 gnd
rlabel metal3 s 7664 58016 7762 58114 4 gnd
rlabel metal3 s 7664 25231 7762 25329 4 gnd
rlabel metal3 s 6425 41449 6523 41547 4 gnd
rlabel metal3 s 7664 74606 7762 74704 4 gnd
rlabel metal3 s 7664 1926 7762 2024 4 gnd
rlabel metal3 s 6425 33965 6523 34063 4 gnd
rlabel metal3 s 7664 51696 7762 51794 4 gnd
rlabel metal3 s 7664 59201 7762 59299 4 gnd
rlabel metal3 s 7664 70656 7762 70754 4 gnd
rlabel metal3 s 6425 81365 6523 81463 4 gnd
rlabel metal3 s 6425 44235 6523 44333 4 gnd
rlabel metal3 s 6425 21325 6523 21423 4 gnd
rlabel metal3 s 7664 92381 7762 92479 4 gnd
rlabel metal3 s 6425 41865 6523 41963 4 gnd
rlabel metal3 s 7664 36686 7762 36784 4 gnd
rlabel metal3 s 7664 19306 7762 19404 4 gnd
rlabel metal3 s 6425 67519 6523 67617 4 gnd
rlabel metal3 s 6425 80949 6523 81047 4 gnd
rlabel metal3 s 7664 59596 7762 59694 4 gnd
rlabel metal3 s 6425 80159 6523 80257 4 gnd
rlabel metal3 s 7664 8246 7762 8344 4 gnd
rlabel metal3 s 6425 24069 6523 24167 4 gnd
rlabel metal3 s 6425 12219 6523 12317 4 gnd
rlabel metal3 s 7664 63941 7762 64039 4 gnd
rlabel metal3 s 6425 75045 6523 75143 4 gnd
rlabel metal3 s 7664 17726 7762 17824 4 gnd
rlabel metal3 s 7664 37476 7762 37574 4 gnd
rlabel metal3 s 7664 47746 7762 47844 4 gnd
rlabel metal3 s 6425 60825 6523 60923 4 gnd
rlabel metal3 s 6425 88059 6523 88157 4 gnd
rlabel metal3 s 7664 23256 7762 23354 4 gnd
rlabel metal3 s 6425 57665 6523 57763 4 gnd
rlabel metal3 s 7664 32736 7762 32834 4 gnd
rlabel metal3 s 7664 94356 7762 94454 4 gnd
rlabel metal3 s 6425 80575 6523 80673 4 gnd
rlabel metal3 s 7664 93171 7762 93269 4 gnd
rlabel metal3 s 6425 61199 6523 61297 4 gnd
rlabel metal3 s 6425 96375 6523 96473 4 gnd
rlabel metal3 s 7664 99096 7762 99194 4 gnd
rlabel metal3 s 7664 63546 7762 63644 4 gnd
rlabel metal3 s 7664 68286 7762 68384 4 gnd
rlabel metal3 s 7664 48536 7762 48634 4 gnd
rlabel metal3 s 2691 8269 2789 8367 4 gnd
rlabel metal3 s 7664 91196 7762 91294 4 gnd
rlabel metal3 s 7664 3901 7762 3999 4 gnd
rlabel metal3 s 7664 99491 7762 99589 4 gnd
rlabel metal3 s 7664 9826 7762 9924 4 gnd
rlabel metal3 s 6425 61615 6523 61713 4 gnd
rlabel metal3 s 6425 55669 6523 55767 4 gnd
rlabel metal3 s 7664 37871 7762 37969 4 gnd
rlabel metal3 s 7664 33921 7762 34019 4 gnd
rlabel metal3 s 6425 15795 6523 15893 4 gnd
rlabel metal3 s 7664 70261 7762 70359 4 gnd
rlabel metal3 s 6425 74629 6523 74727 4 gnd
rlabel metal3 s 6425 9849 6523 9947 4 gnd
rlabel metal3 s 7664 76581 7762 76679 4 gnd
rlabel metal3 s 7664 44981 7762 45079 4 gnd
rlabel metal3 s 6425 78579 6523 78677 4 gnd
rlabel metal3 s 6425 67935 6523 68033 4 gnd
rlabel metal3 s 7664 41426 7762 41524 4 gnd
rlabel metal3 s 6425 64775 6523 64873 4 gnd
rlabel metal3 s 6425 4319 6523 4417 4 gnd
rlabel metal3 s 6425 13799 6523 13897 4 gnd
rlabel metal3 s 2691 6689 2789 6787 4 gnd
rlabel metal3 s 6425 1159 6523 1257 4 gnd
rlabel metal3 s 2691 2739 2789 2837 4 gnd
rlabel metal3 s 7664 18516 7762 18614 4 gnd
rlabel metal3 s 7664 98701 7762 98799 4 gnd
rlabel metal3 s 6425 58039 6523 58137 4 gnd
rlabel metal3 s 7664 18911 7762 19009 4 gnd
rlabel metal3 s 6425 30805 6523 30903 4 gnd
rlabel metal3 s 7664 42216 7762 42314 4 gnd
rlabel metal3 s 7664 38661 7762 38759 4 gnd
rlabel metal3 s 6425 95169 6523 95267 4 gnd
rlabel metal3 s 7664 75791 7762 75889 4 gnd
rlabel metal3 s 7664 62361 7762 62459 4 gnd
rlabel metal3 s 7664 84086 7762 84184 4 gnd
rlabel metal3 s 7664 741 7762 839 4 gnd
rlabel metal3 s 7664 24441 7762 24539 4 gnd
rlabel metal3 s 7664 39451 7762 39549 4 gnd
rlabel metal3 s 6425 99909 6523 100007 4 gnd
rlabel metal3 s 6425 25275 6523 25373 4 gnd
rlabel metal3 s 6425 54879 6523 54977 4 gnd
rlabel metal3 s 7664 80136 7762 80234 4 gnd
rlabel metal3 s 6425 25649 6523 25747 4 gnd
rlabel metal3 s 6425 36709 6523 36807 4 gnd
rlabel metal3 s 6425 37499 6523 37597 4 gnd
rlabel metal3 s 7664 2716 7762 2814 4 gnd
rlabel metal3 s 7664 60386 7762 60484 4 gnd
rlabel metal3 s 7664 36291 7762 36389 4 gnd
rlabel metal3 s 7664 81321 7762 81419 4 gnd
rlabel metal3 s 3930 2716 4028 2814 4 gnd
rlabel metal3 s 7664 73026 7762 73124 4 gnd
rlabel metal3 s 6425 97955 6523 98053 4 gnd
rlabel metal3 s 6425 23695 6523 23793 4 gnd
rlabel metal3 s 7664 85271 7762 85369 4 gnd
rlabel metal3 s 3126 353 3224 451 4 gnd
rlabel metal3 s 7664 67496 7762 67594 4 gnd
rlabel metal3 s 1832 346 1930 444 4 gnd
rlabel metal3 s 7664 93961 7762 94059 4 gnd
rlabel metal3 s 6425 50929 6523 51027 4 gnd
rlabel metal3 s 7664 86851 7762 86949 4 gnd
rlabel metal3 s 7664 21281 7762 21379 4 gnd
rlabel metal3 s 6425 31179 6523 31277 4 gnd
rlabel metal3 s 7664 4296 7762 4394 4 gnd
rlabel metal3 s 6425 50139 6523 50237 4 gnd
rlabel metal3 s 6425 71469 6523 71567 4 gnd
rlabel metal3 s 6425 81739 6523 81837 4 gnd
rlabel metal3 s 6425 7479 6523 7577 4 gnd
rlabel metal3 s 6425 88475 6523 88573 4 gnd
rlabel metal3 s 7664 9431 7762 9529 4 gnd
rlabel metal3 s 6425 78995 6523 79093 4 gnd
rlabel metal3 s 1236 6666 1334 6764 4 gnd
rlabel metal3 s 7664 41821 7762 41919 4 gnd
rlabel metal3 s 7664 55646 7762 55744 4 gnd
rlabel metal3 s 6425 6315 6523 6413 4 gnd
rlabel metal3 s 6425 86105 6523 86203 4 gnd
rlabel metal3 s 6425 91635 6523 91733 4 gnd
rlabel metal3 s 6425 31969 6523 32067 4 gnd
rlabel metal3 s 7664 90011 7762 90109 4 gnd
rlabel metal3 s 2691 4319 2789 4417 4 gnd
rlabel metal3 s 3930 3506 4028 3604 4 gnd
rlabel metal3 s 6425 60409 6523 60507 4 gnd
rlabel metal3 s 6425 75835 6523 75933 4 gnd
rlabel metal3 s 7664 87641 7762 87739 4 gnd
rlabel metal3 s 6425 29599 6523 29697 4 gnd
rlabel metal3 s 7664 84876 7762 84974 4 gnd
rlabel metal3 s 6425 35545 6523 35643 4 gnd
rlabel metal3 s 6425 6689 6523 6787 4 gnd
rlabel metal3 s 7664 16541 7762 16639 4 gnd
rlabel metal3 s 7664 93566 7762 93664 4 gnd
rlabel metal3 s 7664 57621 7762 57719 4 gnd
rlabel metal3 s 6425 60035 6523 60133 4 gnd
rlabel metal3 s 6425 52135 6523 52233 4 gnd
rlabel metal3 s 6425 52509 6523 52607 4 gnd
rlabel metal3 s 6425 51345 6523 51443 4 gnd
rlabel metal3 s 7664 73816 7762 73914 4 gnd
rlabel metal3 s 7664 28786 7762 28884 4 gnd
rlabel metal3 s 6425 15379 6523 15477 4 gnd
rlabel metal3 s 7664 5481 7762 5579 4 gnd
rlabel metal3 s 6425 20119 6523 20217 4 gnd
rlabel metal3 s 6425 69515 6523 69613 4 gnd
rlabel metal3 s 7664 56831 7762 56929 4 gnd
rlabel metal3 s 6425 63195 6523 63293 4 gnd
rlabel metal3 s 6425 43819 6523 43917 4 gnd
rlabel metal3 s 6425 85315 6523 85413 4 gnd
rlabel metal3 s 7664 13381 7762 13479 4 gnd
rlabel metal3 s 6425 87685 6523 87783 4 gnd
rlabel metal3 s 7664 3506 7762 3604 4 gnd
rlabel metal3 s 6425 58829 6523 58927 4 gnd
rlabel metal3 s 6425 63569 6523 63667 4 gnd
rlabel metal3 s 7664 90406 7762 90504 4 gnd
rlabel metal3 s 6425 90429 6523 90527 4 gnd
rlabel metal3 s 7664 51301 7762 51399 4 gnd
rlabel metal3 s 7664 73421 7762 73519 4 gnd
rlabel metal3 s 6425 90845 6523 90943 4 gnd
rlabel metal3 s 6425 45399 6523 45497 4 gnd
rlabel metal3 s 7664 11011 7762 11109 4 gnd
rlabel metal3 s 6425 18539 6523 18637 4 gnd
rlabel metal3 s 6425 64359 6523 64457 4 gnd
rlabel metal3 s 6425 68725 6523 68823 4 gnd
rlabel metal3 s 7664 5086 7762 5184 4 gnd
rlabel metal3 s 7664 40636 7762 40734 4 gnd
rlabel metal3 s 7664 58806 7762 58904 4 gnd
rlabel metal3 s 7664 84481 7762 84579 4 gnd
rlabel metal3 s 7664 31156 7762 31254 4 gnd
rlabel metal3 s 6425 369 6523 467 4 gnd
rlabel metal3 s 7664 31551 7762 31649 4 gnd
rlabel metal3 s 6425 89265 6523 89363 4 gnd
rlabel metal3 s 7664 96331 7762 96429 4 gnd
rlabel metal3 s 7664 95936 7762 96034 4 gnd
rlabel metal3 s 2691 3529 2789 3627 4 gnd
rlabel metal3 s 6425 32759 6523 32857 4 gnd
rlabel metal3 s 6425 46979 6523 47077 4 gnd
rlabel metal3 s 7664 76976 7762 77074 4 gnd
rlabel metal3 s 6425 11055 6523 11153 4 gnd
rlabel metal3 s 7664 65126 7762 65224 4 gnd
rlabel metal3 s 7664 12986 7762 13084 4 gnd
rlabel metal3 s 7664 27206 7762 27304 4 gnd
rlabel metal3 s 7664 346 7762 444 4 gnd
rlabel metal3 s 7664 30366 7762 30464 4 gnd
rlabel metal3 s 6425 82945 6523 83043 4 gnd
rlabel metal3 s 6425 17749 6523 17847 4 gnd
rlabel metal3 s 7664 87246 7762 87344 4 gnd
rlabel metal3 s 6425 98329 6523 98427 4 gnd
rlabel metal3 s 7664 20886 7762 20984 4 gnd
rlabel metal3 s 6425 8269 6523 8367 4 gnd
rlabel metal3 s 6425 50555 6523 50653 4 gnd
rlabel metal3 s 7664 31946 7762 32044 4 gnd
rlabel metal3 s 7664 16146 7762 16244 4 gnd
rlabel metal3 s 3930 346 4028 444 4 gnd
rlabel metal3 s 6425 39079 6523 39177 4 gnd
rlabel metal3 s 7664 69471 7762 69569 4 gnd
rlabel metal3 s 7664 5876 7762 5974 4 gnd
rlabel metal3 s 7664 95541 7762 95639 4 gnd
rlabel metal3 s 7664 52486 7762 52584 4 gnd
rlabel metal3 s 7664 64731 7762 64829 4 gnd
rlabel metal3 s 1236 2716 1334 2814 4 gnd
rlabel metal3 s 6425 77789 6523 77887 4 gnd
rlabel metal3 s 6425 17375 6523 17473 4 gnd
rlabel metal3 s 7664 24836 7762 24934 4 gnd
rlabel metal3 s 6425 72259 6523 72357 4 gnd
rlabel metal3 s 6425 86479 6523 86577 4 gnd
rlabel metal3 s 7664 22466 7762 22564 4 gnd
rlabel metal3 s 6425 52925 6523 53023 4 gnd
rlabel metal3 s 7664 23651 7762 23749 4 gnd
rlabel metal3 s 6425 26439 6523 26537 4 gnd
rlabel metal3 s 7664 50116 7762 50214 4 gnd
rlabel metal3 s 6425 68309 6523 68407 4 gnd
rlabel metal3 s 7664 78951 7762 79049 4 gnd
rlabel metal3 s 7664 3111 7762 3209 4 gnd
rlabel metal3 s 6425 47395 6523 47493 4 gnd
rlabel metal3 s 7664 15751 7762 15849 4 gnd
rlabel metal3 s 7664 75396 7762 75494 4 gnd
rlabel metal3 s 6425 46605 6523 46703 4 gnd
rlabel metal3 s 7664 22071 7762 22169 4 gnd
rlabel metal3 s 6425 95959 6523 96057 4 gnd
rlabel metal3 s 6425 5899 6523 5997 4 gnd
rlabel metal3 s 7664 26811 7762 26909 4 gnd
rlabel metal3 s 6425 15005 6523 15103 4 gnd
rlabel metal3 s 6425 45025 6523 45123 4 gnd
rlabel metal3 s 6425 30389 6523 30487 4 gnd
rlabel metal3 s 6425 67145 6523 67243 4 gnd
rlabel metal3 s 7664 33526 7762 33624 4 gnd
rlabel metal3 s 7664 76186 7762 76284 4 gnd
rlabel metal3 s 7664 78161 7762 78259 4 gnd
rlabel metal3 s 2691 9059 2789 9157 4 gnd
rlabel metal3 s 6425 55295 6523 55393 4 gnd
rlabel metal3 s 6425 99119 6523 99217 4 gnd
rlabel metal3 s 6425 86895 6523 86993 4 gnd
rlabel metal3 s 3930 4296 4028 4394 4 gnd
rlabel metal3 s 7664 99886 7762 99984 4 gnd
rlabel metal3 s 7664 46561 7762 46659 4 gnd
rlabel metal3 s 7664 11801 7762 11899 4 gnd
rlabel metal3 s 6425 59245 6523 59343 4 gnd
rlabel metal3 s 6425 49765 6523 49863 4 gnd
rlabel metal3 s 7664 4691 7762 4789 4 gnd
rlabel metal3 s 6425 83319 6523 83417 4 gnd
rlabel metal3 s 7664 39056 7762 39154 4 gnd
rlabel metal3 s 6425 39869 6523 39967 4 gnd
rlabel metal3 s 6425 82155 6523 82253 4 gnd
rlabel metal3 s 6425 33549 6523 33647 4 gnd
rlabel metal3 s 6425 48975 6523 49073 4 gnd
rlabel metal3 s 6425 94795 6523 94893 4 gnd
rlabel metal3 s 7664 88431 7762 88529 4 gnd
rlabel metal3 s 6425 57249 6523 57347 4 gnd
rlabel metal3 s 6425 13009 6523 13107 4 gnd
rlabel metal3 s 6425 20909 6523 21007 4 gnd
rlabel metal3 s 6425 59619 6523 59717 4 gnd
rlabel metal3 s 6425 65939 6523 66037 4 gnd
rlabel metal3 s 6425 72675 6523 72773 4 gnd
rlabel metal3 s 6425 20535 6523 20633 4 gnd
rlabel metal3 s 7664 10616 7762 10714 4 gnd
rlabel metal3 s 7664 19701 7762 19799 4 gnd
rlabel metal3 s 6425 56459 6523 56557 4 gnd
rlabel metal3 s 7664 2321 7762 2419 4 gnd
rlabel metal3 s 6425 7895 6523 7993 4 gnd
rlabel metal3 s 7664 44191 7762 44289 4 gnd
rlabel metal3 s 7664 71051 7762 71149 4 gnd
rlabel metal3 s 6425 34339 6523 34437 4 gnd
rlabel metal3 s 7664 43796 7762 43894 4 gnd
rlabel metal3 s 3930 1136 4028 1234 4 gnd
rlabel metal3 s 7664 10221 7762 10319 4 gnd
rlabel metal3 s 7664 7061 7762 7159 4 gnd
rlabel metal3 s 6425 56875 6523 56973 4 gnd
rlabel metal3 s 7664 80531 7762 80629 4 gnd
rlabel metal3 s 7664 79741 7762 79839 4 gnd
rlabel metal3 s 6425 98745 6523 98843 4 gnd
rlabel metal3 s 6425 1575 6523 1673 4 gnd
rlabel metal3 s 6425 38705 6523 38803 4 gnd
rlabel metal3 s 6425 28019 6523 28117 4 gnd
rlabel metal3 s 6425 16959 6523 17057 4 gnd
rlabel metal3 s 7664 89616 7762 89714 4 gnd
rlabel metal3 s 7664 11406 7762 11504 4 gnd
rlabel metal3 s 7664 39846 7762 39944 4 gnd
rlabel metal3 s 6425 74255 6523 74353 4 gnd
rlabel metal3 s 6425 87269 6523 87367 4 gnd
rlabel metal3 s 6425 32385 6523 32483 4 gnd
rlabel metal3 s 7664 12591 7762 12689 4 gnd
rlabel metal3 s 7664 56041 7762 56139 4 gnd
rlabel metal3 s 7664 54461 7762 54559 4 gnd
rlabel metal3 s 6425 27229 6523 27327 4 gnd
rlabel metal3 s 6425 62405 6523 62503 4 gnd
rlabel metal3 s 6425 93589 6523 93687 4 gnd
rlabel metal3 s 6425 78205 6523 78303 4 gnd
rlabel metal3 s 6425 36335 6523 36433 4 gnd
rlabel metal3 s 7664 72631 7762 72729 4 gnd
rlabel metal3 s 7664 7851 7762 7949 4 gnd
rlabel metal3 s 7664 22861 7762 22959 4 gnd
rlabel metal3 s 7664 47351 7762 47449 4 gnd
rlabel metal3 s 7664 20491 7762 20589 4 gnd
rlabel metal3 s 6425 23279 6523 23377 4 gnd
rlabel metal3 s 7664 45376 7762 45474 4 gnd
rlabel metal3 s 6425 31595 6523 31693 4 gnd
rlabel metal3 s 7664 95146 7762 95244 4 gnd
rlabel metal3 s 7664 96726 7762 96824 4 gnd
rlabel metal3 s 7664 20096 7762 20194 4 gnd
rlabel metal3 s 7664 97911 7762 98009 4 gnd
rlabel metal3 s 7664 54066 7762 54164 4 gnd
rlabel metal3 s 7664 100281 7762 100379 4 gnd
rlabel metal3 s 3930 9036 4028 9134 4 gnd
rlabel metal3 s 7664 88826 7762 88924 4 gnd
rlabel metal3 s 7664 38266 7762 38364 4 gnd
rlabel metal3 s 7664 54856 7762 54954 4 gnd
rlabel metal3 s 7664 44586 7762 44684 4 gnd
rlabel metal3 s 7664 83296 7762 83394 4 gnd
rlabel metal3 s 6425 26855 6523 26953 4 gnd
rlabel metal3 s 6425 1949 6523 2047 4 gnd
rlabel metal3 s 6425 66729 6523 66827 4 gnd
rlabel metal3 s 7664 55251 7762 55349 4 gnd
rlabel metal3 s 7664 64336 7762 64434 4 gnd
rlabel metal3 s 7664 66706 7762 66804 4 gnd
rlabel metal3 s 6425 45815 6523 45913 4 gnd
rlabel metal3 s 6425 73839 6523 73937 4 gnd
rlabel metal3 s 7664 71446 7762 71544 4 gnd
rlabel metal3 s 6425 16585 6523 16683 4 gnd
rlabel metal3 s 7664 77766 7762 77864 4 gnd
rlabel metal3 s 6425 51719 6523 51817 4 gnd
rlabel metal3 s 6425 96749 6523 96847 4 gnd
rlabel metal3 s 6425 29225 6523 29323 4 gnd
rlabel metal3 s 7664 65521 7762 65619 4 gnd
rlabel metal3 s 7664 37081 7762 37179 4 gnd
rlabel metal3 s 6425 76625 6523 76723 4 gnd
rlabel metal3 s 6425 76209 6523 76307 4 gnd
rlabel metal3 s 7664 89221 7762 89319 4 gnd
rlabel metal3 s 7664 46956 7762 47054 4 gnd
rlabel metal3 s 6425 28809 6523 28907 4 gnd
rlabel metal3 s 3930 7456 4028 7554 4 gnd
rlabel metal3 s 6425 35919 6523 36017 4 gnd
rlabel metal3 s 7664 71841 7762 71939 4 gnd
rlabel metal3 s 7664 82901 7762 82999 4 gnd
rlabel metal3 s 7664 92776 7762 92874 4 gnd
rlabel metal3 s 6425 40285 6523 40383 4 gnd
rlabel metal3 s 6425 83735 6523 83833 4 gnd
rlabel metal3 s 6425 11845 6523 11943 4 gnd
rlabel metal3 s 6425 85689 6523 85787 4 gnd
rlabel metal3 s 6425 66355 6523 66453 4 gnd
rlabel metal3 s 7664 9036 7762 9134 4 gnd
rlabel metal3 s 7664 86456 7762 86554 4 gnd
rlabel metal3 s 7664 61571 7762 61669 4 gnd
rlabel metal3 s 6425 92425 6523 92523 4 gnd
rlabel metal3 s 6425 92009 6523 92107 4 gnd
rlabel metal3 s 7664 35106 7762 35204 4 gnd
rlabel metal3 s 7664 79346 7762 79444 4 gnd
rlabel metal3 s 6425 79785 6523 79883 4 gnd
rlabel metal3 s 6425 84109 6523 84207 4 gnd
rlabel metal3 s 6425 54089 6523 54187 4 gnd
rlabel metal3 s 6425 73465 6523 73563 4 gnd
rlabel metal3 s 6425 40659 6523 40757 4 gnd
rlabel metal3 s 6425 69889 6523 69987 4 gnd
rlabel metal3 s 7664 29971 7762 30069 4 gnd
rlabel metal3 s 6425 5109 6523 5207 4 gnd
rlabel metal3 s 6425 95585 6523 95683 4 gnd
rlabel metal3 s 6425 43445 6523 43543 4 gnd
rlabel metal3 s 7664 97121 7762 97219 4 gnd
rlabel metal3 s 6425 48559 6523 48657 4 gnd
rlabel metal3 s 7664 67101 7762 67199 4 gnd
rlabel metal3 s 7664 12196 7762 12294 4 gnd
rlabel metal3 s 6425 88849 6523 88947 4 gnd
rlabel metal3 s 6425 27645 6523 27743 4 gnd
rlabel metal3 s 6425 785 6523 883 4 gnd
rlabel metal3 s 6425 75419 6523 75517 4 gnd
rlabel metal3 s 7664 25626 7762 25724 4 gnd
rlabel metal3 s 7664 6271 7762 6369 4 gnd
rlabel metal3 s 7664 40241 7762 40339 4 gnd
rlabel metal3 s 6425 82529 6523 82627 4 gnd
rlabel metal3 s 7664 80926 7762 81024 4 gnd
rlabel metal3 s 7664 34316 7762 34414 4 gnd
rlabel metal3 s 7664 50906 7762 51004 4 gnd
rlabel metal3 s 7664 53671 7762 53769 4 gnd
rlabel metal3 s 6425 93215 6523 93313 4 gnd
rlabel metal3 s 6425 37915 6523 38013 4 gnd
rlabel metal3 s 7664 13776 7762 13874 4 gnd
rlabel metal3 s 7664 88036 7762 88134 4 gnd
rlabel metal3 s 7664 21676 7762 21774 4 gnd
rlabel metal3 s 6425 48185 6523 48283 4 gnd
rlabel metal3 s 7664 27996 7762 28094 4 gnd
rlabel metal3 s 6425 71095 6523 71193 4 gnd
rlabel metal3 s 7664 91986 7762 92084 4 gnd
rlabel metal3 s 7664 17331 7762 17429 4 gnd
rlabel metal3 s 7664 14566 7762 14664 4 gnd
rlabel metal3 s 6425 19329 6523 19427 4 gnd
rlabel metal3 s 3930 8246 4028 8344 4 gnd
rlabel metal3 s 7664 58411 7762 58509 4 gnd
rlabel metal3 s 7664 78556 7762 78654 4 gnd
rlabel metal3 s 6425 69099 6523 69197 4 gnd
rlabel metal3 s 7664 35501 7762 35599 4 gnd
rlabel metal3 s 7664 75001 7762 75099 4 gnd
rlabel metal3 s 7664 6666 7762 6764 4 gnd
rlabel metal3 s 2691 5109 2789 5207 4 gnd
rlabel metal3 s 6425 22905 6523 23003 4 gnd
rlabel metal3 s 6425 3529 6523 3627 4 gnd
rlabel metal3 s 6425 3945 6523 4043 4 gnd
rlabel metal3 s 6425 12635 6523 12733 4 gnd
rlabel metal3 s 6425 22489 6523 22587 4 gnd
rlabel metal3 s 7664 52881 7762 52979 4 gnd
rlabel metal3 s 7664 60781 7762 60879 4 gnd
rlabel metal3 s 6425 9059 6523 9157 4 gnd
rlabel metal3 s 6425 94005 6523 94103 4 gnd
rlabel metal3 s 6425 73049 6523 73147 4 gnd
rlabel metal3 s 7664 74211 7762 74309 4 gnd
rlabel metal3 s 6425 99535 6523 99633 4 gnd
rlabel metal3 s 7664 100676 7762 100774 4 gnd
rlabel metal3 s 6425 54505 6523 54603 4 gnd
rlabel metal3 s 6425 84899 6523 84997 4 gnd
rlabel metal3 s 3930 5086 4028 5184 4 gnd
rlabel metal3 s 6425 30015 6523 30113 4 gnd
rlabel metal3 s 7664 68681 7762 68779 4 gnd
rlabel metal3 s 6425 61989 6523 62087 4 gnd
rlabel metal3 s 7664 48931 7762 49029 4 gnd
rlabel metal3 s 6425 18955 6523 19053 4 gnd
rlabel metal3 s 7664 62756 7762 62854 4 gnd
rlabel metal3 s 6425 37125 6523 37223 4 gnd
rlabel metal3 s 7664 94751 7762 94849 4 gnd
rlabel metal3 s 7664 24046 7762 24144 4 gnd
rlabel metal3 s 6425 41075 6523 41173 4 gnd
rlabel metal3 s 7664 34711 7762 34809 4 gnd
rlabel metal3 s 6425 10639 6523 10737 4 gnd
rlabel metal3 s 7664 1531 7762 1629 4 gnd
rlabel metal3 s 6425 53299 6523 53397 4 gnd
rlabel metal3 s 6425 26065 6523 26163 4 gnd
rlabel metal3 s 7664 48141 7762 48239 4 gnd
rlabel metal3 s 6425 63985 6523 64083 4 gnd
rlabel metal3 s 6425 14589 6523 14687 4 gnd
rlabel metal3 s 6425 44609 6523 44707 4 gnd
rlabel metal3 s 6425 13425 6523 13523 4 gnd
rlabel metal3 s 7664 77371 7762 77469 4 gnd
rlabel metal3 s 7664 15356 7762 15454 4 gnd
rlabel metal3 s 6425 42239 6523 42337 4 gnd
rlabel metal3 s 7664 1136 7762 1234 4 gnd
rlabel metal3 s 6425 94379 6523 94477 4 gnd
rlabel metal3 s 6425 100699 6523 100797 4 gnd
rlabel metal3 s 7664 72236 7762 72334 4 gnd
rlabel metal3 s 7664 98306 7762 98404 4 gnd
rlabel metal3 s 7664 26416 7762 26514 4 gnd
rlabel metal3 s 7664 90801 7762 90899 4 gnd
rlabel metal3 s 7664 97516 7762 97614 4 gnd
rlabel metal3 s 7664 67891 7762 67989 4 gnd
rlabel metal3 s 7664 53276 7762 53374 4 gnd
rlabel metal3 s 7664 56436 7762 56534 4 gnd
rlabel metal3 s 7664 41031 7762 41129 4 gnd
rlabel metal3 s 7664 43006 7762 43104 4 gnd
rlabel metal3 s 6425 91219 6523 91317 4 gnd
rlabel metal3 s 7664 7456 7762 7554 4 gnd
rlabel metal3 s 6425 62779 6523 62877 4 gnd
rlabel metal3 s 7664 69866 7762 69964 4 gnd
rlabel metal3 s 7664 16936 7762 17034 4 gnd
rlabel metal3 s 7664 29576 7762 29674 4 gnd
rlabel metal3 s 6425 90055 6523 90153 4 gnd
rlabel metal3 s 7664 27601 7762 27699 4 gnd
rlabel metal3 s 6425 65565 6523 65663 4 gnd
rlabel metal3 s 6425 24485 6523 24583 4 gnd
rlabel metal3 s 6425 18165 6523 18263 4 gnd
rlabel metal3 s 6425 11429 6523 11527 4 gnd
rlabel metal3 s 7664 82506 7762 82604 4 gnd
rlabel metal3 s 3930 6666 4028 6764 4 gnd
rlabel metal3 s 6425 76999 6523 77097 4 gnd
rlabel metal3 s 7664 33131 7762 33229 4 gnd
rlabel metal3 s 7664 14961 7762 15059 4 gnd
rlabel metal3 s 3126 1143 3224 1241 4 gnd
rlabel metal3 s 7664 14171 7762 14269 4 gnd
rlabel metal3 s 7664 46166 7762 46264 4 gnd
rlabel metal3 s 7664 49721 7762 49819 4 gnd
<< properties >>
string FIXED_BBOX 0 0 8271 101148
<< end >>
