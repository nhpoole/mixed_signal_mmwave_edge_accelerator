magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect -6405 -1648 6405 1648
<< pwell >>
rect -5145 -326 5145 326
<< nmos >>
rect -5061 -300 -4101 300
rect -4043 -300 -3083 300
rect -3025 -300 -2065 300
rect -2007 -300 -1047 300
rect -989 -300 -29 300
rect 29 -300 989 300
rect 1047 -300 2007 300
rect 2065 -300 3025 300
rect 3083 -300 4043 300
rect 4101 -300 5061 300
<< ndiff >>
rect -5119 255 -5061 300
rect -5119 221 -5107 255
rect -5073 221 -5061 255
rect -5119 187 -5061 221
rect -5119 153 -5107 187
rect -5073 153 -5061 187
rect -5119 119 -5061 153
rect -5119 85 -5107 119
rect -5073 85 -5061 119
rect -5119 51 -5061 85
rect -5119 17 -5107 51
rect -5073 17 -5061 51
rect -5119 -17 -5061 17
rect -5119 -51 -5107 -17
rect -5073 -51 -5061 -17
rect -5119 -85 -5061 -51
rect -5119 -119 -5107 -85
rect -5073 -119 -5061 -85
rect -5119 -153 -5061 -119
rect -5119 -187 -5107 -153
rect -5073 -187 -5061 -153
rect -5119 -221 -5061 -187
rect -5119 -255 -5107 -221
rect -5073 -255 -5061 -221
rect -5119 -300 -5061 -255
rect -4101 255 -4043 300
rect -4101 221 -4089 255
rect -4055 221 -4043 255
rect -4101 187 -4043 221
rect -4101 153 -4089 187
rect -4055 153 -4043 187
rect -4101 119 -4043 153
rect -4101 85 -4089 119
rect -4055 85 -4043 119
rect -4101 51 -4043 85
rect -4101 17 -4089 51
rect -4055 17 -4043 51
rect -4101 -17 -4043 17
rect -4101 -51 -4089 -17
rect -4055 -51 -4043 -17
rect -4101 -85 -4043 -51
rect -4101 -119 -4089 -85
rect -4055 -119 -4043 -85
rect -4101 -153 -4043 -119
rect -4101 -187 -4089 -153
rect -4055 -187 -4043 -153
rect -4101 -221 -4043 -187
rect -4101 -255 -4089 -221
rect -4055 -255 -4043 -221
rect -4101 -300 -4043 -255
rect -3083 255 -3025 300
rect -3083 221 -3071 255
rect -3037 221 -3025 255
rect -3083 187 -3025 221
rect -3083 153 -3071 187
rect -3037 153 -3025 187
rect -3083 119 -3025 153
rect -3083 85 -3071 119
rect -3037 85 -3025 119
rect -3083 51 -3025 85
rect -3083 17 -3071 51
rect -3037 17 -3025 51
rect -3083 -17 -3025 17
rect -3083 -51 -3071 -17
rect -3037 -51 -3025 -17
rect -3083 -85 -3025 -51
rect -3083 -119 -3071 -85
rect -3037 -119 -3025 -85
rect -3083 -153 -3025 -119
rect -3083 -187 -3071 -153
rect -3037 -187 -3025 -153
rect -3083 -221 -3025 -187
rect -3083 -255 -3071 -221
rect -3037 -255 -3025 -221
rect -3083 -300 -3025 -255
rect -2065 255 -2007 300
rect -2065 221 -2053 255
rect -2019 221 -2007 255
rect -2065 187 -2007 221
rect -2065 153 -2053 187
rect -2019 153 -2007 187
rect -2065 119 -2007 153
rect -2065 85 -2053 119
rect -2019 85 -2007 119
rect -2065 51 -2007 85
rect -2065 17 -2053 51
rect -2019 17 -2007 51
rect -2065 -17 -2007 17
rect -2065 -51 -2053 -17
rect -2019 -51 -2007 -17
rect -2065 -85 -2007 -51
rect -2065 -119 -2053 -85
rect -2019 -119 -2007 -85
rect -2065 -153 -2007 -119
rect -2065 -187 -2053 -153
rect -2019 -187 -2007 -153
rect -2065 -221 -2007 -187
rect -2065 -255 -2053 -221
rect -2019 -255 -2007 -221
rect -2065 -300 -2007 -255
rect -1047 255 -989 300
rect -1047 221 -1035 255
rect -1001 221 -989 255
rect -1047 187 -989 221
rect -1047 153 -1035 187
rect -1001 153 -989 187
rect -1047 119 -989 153
rect -1047 85 -1035 119
rect -1001 85 -989 119
rect -1047 51 -989 85
rect -1047 17 -1035 51
rect -1001 17 -989 51
rect -1047 -17 -989 17
rect -1047 -51 -1035 -17
rect -1001 -51 -989 -17
rect -1047 -85 -989 -51
rect -1047 -119 -1035 -85
rect -1001 -119 -989 -85
rect -1047 -153 -989 -119
rect -1047 -187 -1035 -153
rect -1001 -187 -989 -153
rect -1047 -221 -989 -187
rect -1047 -255 -1035 -221
rect -1001 -255 -989 -221
rect -1047 -300 -989 -255
rect -29 255 29 300
rect -29 221 -17 255
rect 17 221 29 255
rect -29 187 29 221
rect -29 153 -17 187
rect 17 153 29 187
rect -29 119 29 153
rect -29 85 -17 119
rect 17 85 29 119
rect -29 51 29 85
rect -29 17 -17 51
rect 17 17 29 51
rect -29 -17 29 17
rect -29 -51 -17 -17
rect 17 -51 29 -17
rect -29 -85 29 -51
rect -29 -119 -17 -85
rect 17 -119 29 -85
rect -29 -153 29 -119
rect -29 -187 -17 -153
rect 17 -187 29 -153
rect -29 -221 29 -187
rect -29 -255 -17 -221
rect 17 -255 29 -221
rect -29 -300 29 -255
rect 989 255 1047 300
rect 989 221 1001 255
rect 1035 221 1047 255
rect 989 187 1047 221
rect 989 153 1001 187
rect 1035 153 1047 187
rect 989 119 1047 153
rect 989 85 1001 119
rect 1035 85 1047 119
rect 989 51 1047 85
rect 989 17 1001 51
rect 1035 17 1047 51
rect 989 -17 1047 17
rect 989 -51 1001 -17
rect 1035 -51 1047 -17
rect 989 -85 1047 -51
rect 989 -119 1001 -85
rect 1035 -119 1047 -85
rect 989 -153 1047 -119
rect 989 -187 1001 -153
rect 1035 -187 1047 -153
rect 989 -221 1047 -187
rect 989 -255 1001 -221
rect 1035 -255 1047 -221
rect 989 -300 1047 -255
rect 2007 255 2065 300
rect 2007 221 2019 255
rect 2053 221 2065 255
rect 2007 187 2065 221
rect 2007 153 2019 187
rect 2053 153 2065 187
rect 2007 119 2065 153
rect 2007 85 2019 119
rect 2053 85 2065 119
rect 2007 51 2065 85
rect 2007 17 2019 51
rect 2053 17 2065 51
rect 2007 -17 2065 17
rect 2007 -51 2019 -17
rect 2053 -51 2065 -17
rect 2007 -85 2065 -51
rect 2007 -119 2019 -85
rect 2053 -119 2065 -85
rect 2007 -153 2065 -119
rect 2007 -187 2019 -153
rect 2053 -187 2065 -153
rect 2007 -221 2065 -187
rect 2007 -255 2019 -221
rect 2053 -255 2065 -221
rect 2007 -300 2065 -255
rect 3025 255 3083 300
rect 3025 221 3037 255
rect 3071 221 3083 255
rect 3025 187 3083 221
rect 3025 153 3037 187
rect 3071 153 3083 187
rect 3025 119 3083 153
rect 3025 85 3037 119
rect 3071 85 3083 119
rect 3025 51 3083 85
rect 3025 17 3037 51
rect 3071 17 3083 51
rect 3025 -17 3083 17
rect 3025 -51 3037 -17
rect 3071 -51 3083 -17
rect 3025 -85 3083 -51
rect 3025 -119 3037 -85
rect 3071 -119 3083 -85
rect 3025 -153 3083 -119
rect 3025 -187 3037 -153
rect 3071 -187 3083 -153
rect 3025 -221 3083 -187
rect 3025 -255 3037 -221
rect 3071 -255 3083 -221
rect 3025 -300 3083 -255
rect 4043 255 4101 300
rect 4043 221 4055 255
rect 4089 221 4101 255
rect 4043 187 4101 221
rect 4043 153 4055 187
rect 4089 153 4101 187
rect 4043 119 4101 153
rect 4043 85 4055 119
rect 4089 85 4101 119
rect 4043 51 4101 85
rect 4043 17 4055 51
rect 4089 17 4101 51
rect 4043 -17 4101 17
rect 4043 -51 4055 -17
rect 4089 -51 4101 -17
rect 4043 -85 4101 -51
rect 4043 -119 4055 -85
rect 4089 -119 4101 -85
rect 4043 -153 4101 -119
rect 4043 -187 4055 -153
rect 4089 -187 4101 -153
rect 4043 -221 4101 -187
rect 4043 -255 4055 -221
rect 4089 -255 4101 -221
rect 4043 -300 4101 -255
rect 5061 255 5119 300
rect 5061 221 5073 255
rect 5107 221 5119 255
rect 5061 187 5119 221
rect 5061 153 5073 187
rect 5107 153 5119 187
rect 5061 119 5119 153
rect 5061 85 5073 119
rect 5107 85 5119 119
rect 5061 51 5119 85
rect 5061 17 5073 51
rect 5107 17 5119 51
rect 5061 -17 5119 17
rect 5061 -51 5073 -17
rect 5107 -51 5119 -17
rect 5061 -85 5119 -51
rect 5061 -119 5073 -85
rect 5107 -119 5119 -85
rect 5061 -153 5119 -119
rect 5061 -187 5073 -153
rect 5107 -187 5119 -153
rect 5061 -221 5119 -187
rect 5061 -255 5073 -221
rect 5107 -255 5119 -221
rect 5061 -300 5119 -255
<< ndiffc >>
rect -5107 221 -5073 255
rect -5107 153 -5073 187
rect -5107 85 -5073 119
rect -5107 17 -5073 51
rect -5107 -51 -5073 -17
rect -5107 -119 -5073 -85
rect -5107 -187 -5073 -153
rect -5107 -255 -5073 -221
rect -4089 221 -4055 255
rect -4089 153 -4055 187
rect -4089 85 -4055 119
rect -4089 17 -4055 51
rect -4089 -51 -4055 -17
rect -4089 -119 -4055 -85
rect -4089 -187 -4055 -153
rect -4089 -255 -4055 -221
rect -3071 221 -3037 255
rect -3071 153 -3037 187
rect -3071 85 -3037 119
rect -3071 17 -3037 51
rect -3071 -51 -3037 -17
rect -3071 -119 -3037 -85
rect -3071 -187 -3037 -153
rect -3071 -255 -3037 -221
rect -2053 221 -2019 255
rect -2053 153 -2019 187
rect -2053 85 -2019 119
rect -2053 17 -2019 51
rect -2053 -51 -2019 -17
rect -2053 -119 -2019 -85
rect -2053 -187 -2019 -153
rect -2053 -255 -2019 -221
rect -1035 221 -1001 255
rect -1035 153 -1001 187
rect -1035 85 -1001 119
rect -1035 17 -1001 51
rect -1035 -51 -1001 -17
rect -1035 -119 -1001 -85
rect -1035 -187 -1001 -153
rect -1035 -255 -1001 -221
rect -17 221 17 255
rect -17 153 17 187
rect -17 85 17 119
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -119 17 -85
rect -17 -187 17 -153
rect -17 -255 17 -221
rect 1001 221 1035 255
rect 1001 153 1035 187
rect 1001 85 1035 119
rect 1001 17 1035 51
rect 1001 -51 1035 -17
rect 1001 -119 1035 -85
rect 1001 -187 1035 -153
rect 1001 -255 1035 -221
rect 2019 221 2053 255
rect 2019 153 2053 187
rect 2019 85 2053 119
rect 2019 17 2053 51
rect 2019 -51 2053 -17
rect 2019 -119 2053 -85
rect 2019 -187 2053 -153
rect 2019 -255 2053 -221
rect 3037 221 3071 255
rect 3037 153 3071 187
rect 3037 85 3071 119
rect 3037 17 3071 51
rect 3037 -51 3071 -17
rect 3037 -119 3071 -85
rect 3037 -187 3071 -153
rect 3037 -255 3071 -221
rect 4055 221 4089 255
rect 4055 153 4089 187
rect 4055 85 4089 119
rect 4055 17 4089 51
rect 4055 -51 4089 -17
rect 4055 -119 4089 -85
rect 4055 -187 4089 -153
rect 4055 -255 4089 -221
rect 5073 221 5107 255
rect 5073 153 5107 187
rect 5073 85 5107 119
rect 5073 17 5107 51
rect 5073 -51 5107 -17
rect 5073 -119 5107 -85
rect 5073 -187 5107 -153
rect 5073 -255 5107 -221
<< poly >>
rect -4875 372 -4287 388
rect -4875 355 -4836 372
rect -5061 338 -4836 355
rect -4802 338 -4768 372
rect -4734 338 -4700 372
rect -4666 338 -4632 372
rect -4598 338 -4564 372
rect -4530 338 -4496 372
rect -4462 338 -4428 372
rect -4394 338 -4360 372
rect -4326 355 -4287 372
rect -3857 372 -3269 388
rect -3857 355 -3818 372
rect -4326 338 -4101 355
rect -5061 300 -4101 338
rect -4043 338 -3818 355
rect -3784 338 -3750 372
rect -3716 338 -3682 372
rect -3648 338 -3614 372
rect -3580 338 -3546 372
rect -3512 338 -3478 372
rect -3444 338 -3410 372
rect -3376 338 -3342 372
rect -3308 355 -3269 372
rect -2839 372 -2251 388
rect -2839 355 -2800 372
rect -3308 338 -3083 355
rect -4043 300 -3083 338
rect -3025 338 -2800 355
rect -2766 338 -2732 372
rect -2698 338 -2664 372
rect -2630 338 -2596 372
rect -2562 338 -2528 372
rect -2494 338 -2460 372
rect -2426 338 -2392 372
rect -2358 338 -2324 372
rect -2290 355 -2251 372
rect -1821 372 -1233 388
rect -1821 355 -1782 372
rect -2290 338 -2065 355
rect -3025 300 -2065 338
rect -2007 338 -1782 355
rect -1748 338 -1714 372
rect -1680 338 -1646 372
rect -1612 338 -1578 372
rect -1544 338 -1510 372
rect -1476 338 -1442 372
rect -1408 338 -1374 372
rect -1340 338 -1306 372
rect -1272 355 -1233 372
rect -803 372 -215 388
rect -803 355 -764 372
rect -1272 338 -1047 355
rect -2007 300 -1047 338
rect -989 338 -764 355
rect -730 338 -696 372
rect -662 338 -628 372
rect -594 338 -560 372
rect -526 338 -492 372
rect -458 338 -424 372
rect -390 338 -356 372
rect -322 338 -288 372
rect -254 355 -215 372
rect 215 372 803 388
rect 215 355 254 372
rect -254 338 -29 355
rect -989 300 -29 338
rect 29 338 254 355
rect 288 338 322 372
rect 356 338 390 372
rect 424 338 458 372
rect 492 338 526 372
rect 560 338 594 372
rect 628 338 662 372
rect 696 338 730 372
rect 764 355 803 372
rect 1233 372 1821 388
rect 1233 355 1272 372
rect 764 338 989 355
rect 29 300 989 338
rect 1047 338 1272 355
rect 1306 338 1340 372
rect 1374 338 1408 372
rect 1442 338 1476 372
rect 1510 338 1544 372
rect 1578 338 1612 372
rect 1646 338 1680 372
rect 1714 338 1748 372
rect 1782 355 1821 372
rect 2251 372 2839 388
rect 2251 355 2290 372
rect 1782 338 2007 355
rect 1047 300 2007 338
rect 2065 338 2290 355
rect 2324 338 2358 372
rect 2392 338 2426 372
rect 2460 338 2494 372
rect 2528 338 2562 372
rect 2596 338 2630 372
rect 2664 338 2698 372
rect 2732 338 2766 372
rect 2800 355 2839 372
rect 3269 372 3857 388
rect 3269 355 3308 372
rect 2800 338 3025 355
rect 2065 300 3025 338
rect 3083 338 3308 355
rect 3342 338 3376 372
rect 3410 338 3444 372
rect 3478 338 3512 372
rect 3546 338 3580 372
rect 3614 338 3648 372
rect 3682 338 3716 372
rect 3750 338 3784 372
rect 3818 355 3857 372
rect 4287 372 4875 388
rect 4287 355 4326 372
rect 3818 338 4043 355
rect 3083 300 4043 338
rect 4101 338 4326 355
rect 4360 338 4394 372
rect 4428 338 4462 372
rect 4496 338 4530 372
rect 4564 338 4598 372
rect 4632 338 4666 372
rect 4700 338 4734 372
rect 4768 338 4802 372
rect 4836 355 4875 372
rect 4836 338 5061 355
rect 4101 300 5061 338
rect -5061 -338 -4101 -300
rect -5061 -355 -4836 -338
rect -4875 -372 -4836 -355
rect -4802 -372 -4768 -338
rect -4734 -372 -4700 -338
rect -4666 -372 -4632 -338
rect -4598 -372 -4564 -338
rect -4530 -372 -4496 -338
rect -4462 -372 -4428 -338
rect -4394 -372 -4360 -338
rect -4326 -355 -4101 -338
rect -4043 -338 -3083 -300
rect -4043 -355 -3818 -338
rect -4326 -372 -4287 -355
rect -4875 -388 -4287 -372
rect -3857 -372 -3818 -355
rect -3784 -372 -3750 -338
rect -3716 -372 -3682 -338
rect -3648 -372 -3614 -338
rect -3580 -372 -3546 -338
rect -3512 -372 -3478 -338
rect -3444 -372 -3410 -338
rect -3376 -372 -3342 -338
rect -3308 -355 -3083 -338
rect -3025 -338 -2065 -300
rect -3025 -355 -2800 -338
rect -3308 -372 -3269 -355
rect -3857 -388 -3269 -372
rect -2839 -372 -2800 -355
rect -2766 -372 -2732 -338
rect -2698 -372 -2664 -338
rect -2630 -372 -2596 -338
rect -2562 -372 -2528 -338
rect -2494 -372 -2460 -338
rect -2426 -372 -2392 -338
rect -2358 -372 -2324 -338
rect -2290 -355 -2065 -338
rect -2007 -338 -1047 -300
rect -2007 -355 -1782 -338
rect -2290 -372 -2251 -355
rect -2839 -388 -2251 -372
rect -1821 -372 -1782 -355
rect -1748 -372 -1714 -338
rect -1680 -372 -1646 -338
rect -1612 -372 -1578 -338
rect -1544 -372 -1510 -338
rect -1476 -372 -1442 -338
rect -1408 -372 -1374 -338
rect -1340 -372 -1306 -338
rect -1272 -355 -1047 -338
rect -989 -338 -29 -300
rect -989 -355 -764 -338
rect -1272 -372 -1233 -355
rect -1821 -388 -1233 -372
rect -803 -372 -764 -355
rect -730 -372 -696 -338
rect -662 -372 -628 -338
rect -594 -372 -560 -338
rect -526 -372 -492 -338
rect -458 -372 -424 -338
rect -390 -372 -356 -338
rect -322 -372 -288 -338
rect -254 -355 -29 -338
rect 29 -338 989 -300
rect 29 -355 254 -338
rect -254 -372 -215 -355
rect -803 -388 -215 -372
rect 215 -372 254 -355
rect 288 -372 322 -338
rect 356 -372 390 -338
rect 424 -372 458 -338
rect 492 -372 526 -338
rect 560 -372 594 -338
rect 628 -372 662 -338
rect 696 -372 730 -338
rect 764 -355 989 -338
rect 1047 -338 2007 -300
rect 1047 -355 1272 -338
rect 764 -372 803 -355
rect 215 -388 803 -372
rect 1233 -372 1272 -355
rect 1306 -372 1340 -338
rect 1374 -372 1408 -338
rect 1442 -372 1476 -338
rect 1510 -372 1544 -338
rect 1578 -372 1612 -338
rect 1646 -372 1680 -338
rect 1714 -372 1748 -338
rect 1782 -355 2007 -338
rect 2065 -338 3025 -300
rect 2065 -355 2290 -338
rect 1782 -372 1821 -355
rect 1233 -388 1821 -372
rect 2251 -372 2290 -355
rect 2324 -372 2358 -338
rect 2392 -372 2426 -338
rect 2460 -372 2494 -338
rect 2528 -372 2562 -338
rect 2596 -372 2630 -338
rect 2664 -372 2698 -338
rect 2732 -372 2766 -338
rect 2800 -355 3025 -338
rect 3083 -338 4043 -300
rect 3083 -355 3308 -338
rect 2800 -372 2839 -355
rect 2251 -388 2839 -372
rect 3269 -372 3308 -355
rect 3342 -372 3376 -338
rect 3410 -372 3444 -338
rect 3478 -372 3512 -338
rect 3546 -372 3580 -338
rect 3614 -372 3648 -338
rect 3682 -372 3716 -338
rect 3750 -372 3784 -338
rect 3818 -355 4043 -338
rect 4101 -338 5061 -300
rect 4101 -355 4326 -338
rect 3818 -372 3857 -355
rect 3269 -388 3857 -372
rect 4287 -372 4326 -355
rect 4360 -372 4394 -338
rect 4428 -372 4462 -338
rect 4496 -372 4530 -338
rect 4564 -372 4598 -338
rect 4632 -372 4666 -338
rect 4700 -372 4734 -338
rect 4768 -372 4802 -338
rect 4836 -355 5061 -338
rect 4836 -372 4875 -355
rect 4287 -388 4875 -372
<< polycont >>
rect -4836 338 -4802 372
rect -4768 338 -4734 372
rect -4700 338 -4666 372
rect -4632 338 -4598 372
rect -4564 338 -4530 372
rect -4496 338 -4462 372
rect -4428 338 -4394 372
rect -4360 338 -4326 372
rect -3818 338 -3784 372
rect -3750 338 -3716 372
rect -3682 338 -3648 372
rect -3614 338 -3580 372
rect -3546 338 -3512 372
rect -3478 338 -3444 372
rect -3410 338 -3376 372
rect -3342 338 -3308 372
rect -2800 338 -2766 372
rect -2732 338 -2698 372
rect -2664 338 -2630 372
rect -2596 338 -2562 372
rect -2528 338 -2494 372
rect -2460 338 -2426 372
rect -2392 338 -2358 372
rect -2324 338 -2290 372
rect -1782 338 -1748 372
rect -1714 338 -1680 372
rect -1646 338 -1612 372
rect -1578 338 -1544 372
rect -1510 338 -1476 372
rect -1442 338 -1408 372
rect -1374 338 -1340 372
rect -1306 338 -1272 372
rect -764 338 -730 372
rect -696 338 -662 372
rect -628 338 -594 372
rect -560 338 -526 372
rect -492 338 -458 372
rect -424 338 -390 372
rect -356 338 -322 372
rect -288 338 -254 372
rect 254 338 288 372
rect 322 338 356 372
rect 390 338 424 372
rect 458 338 492 372
rect 526 338 560 372
rect 594 338 628 372
rect 662 338 696 372
rect 730 338 764 372
rect 1272 338 1306 372
rect 1340 338 1374 372
rect 1408 338 1442 372
rect 1476 338 1510 372
rect 1544 338 1578 372
rect 1612 338 1646 372
rect 1680 338 1714 372
rect 1748 338 1782 372
rect 2290 338 2324 372
rect 2358 338 2392 372
rect 2426 338 2460 372
rect 2494 338 2528 372
rect 2562 338 2596 372
rect 2630 338 2664 372
rect 2698 338 2732 372
rect 2766 338 2800 372
rect 3308 338 3342 372
rect 3376 338 3410 372
rect 3444 338 3478 372
rect 3512 338 3546 372
rect 3580 338 3614 372
rect 3648 338 3682 372
rect 3716 338 3750 372
rect 3784 338 3818 372
rect 4326 338 4360 372
rect 4394 338 4428 372
rect 4462 338 4496 372
rect 4530 338 4564 372
rect 4598 338 4632 372
rect 4666 338 4700 372
rect 4734 338 4768 372
rect 4802 338 4836 372
rect -4836 -372 -4802 -338
rect -4768 -372 -4734 -338
rect -4700 -372 -4666 -338
rect -4632 -372 -4598 -338
rect -4564 -372 -4530 -338
rect -4496 -372 -4462 -338
rect -4428 -372 -4394 -338
rect -4360 -372 -4326 -338
rect -3818 -372 -3784 -338
rect -3750 -372 -3716 -338
rect -3682 -372 -3648 -338
rect -3614 -372 -3580 -338
rect -3546 -372 -3512 -338
rect -3478 -372 -3444 -338
rect -3410 -372 -3376 -338
rect -3342 -372 -3308 -338
rect -2800 -372 -2766 -338
rect -2732 -372 -2698 -338
rect -2664 -372 -2630 -338
rect -2596 -372 -2562 -338
rect -2528 -372 -2494 -338
rect -2460 -372 -2426 -338
rect -2392 -372 -2358 -338
rect -2324 -372 -2290 -338
rect -1782 -372 -1748 -338
rect -1714 -372 -1680 -338
rect -1646 -372 -1612 -338
rect -1578 -372 -1544 -338
rect -1510 -372 -1476 -338
rect -1442 -372 -1408 -338
rect -1374 -372 -1340 -338
rect -1306 -372 -1272 -338
rect -764 -372 -730 -338
rect -696 -372 -662 -338
rect -628 -372 -594 -338
rect -560 -372 -526 -338
rect -492 -372 -458 -338
rect -424 -372 -390 -338
rect -356 -372 -322 -338
rect -288 -372 -254 -338
rect 254 -372 288 -338
rect 322 -372 356 -338
rect 390 -372 424 -338
rect 458 -372 492 -338
rect 526 -372 560 -338
rect 594 -372 628 -338
rect 662 -372 696 -338
rect 730 -372 764 -338
rect 1272 -372 1306 -338
rect 1340 -372 1374 -338
rect 1408 -372 1442 -338
rect 1476 -372 1510 -338
rect 1544 -372 1578 -338
rect 1612 -372 1646 -338
rect 1680 -372 1714 -338
rect 1748 -372 1782 -338
rect 2290 -372 2324 -338
rect 2358 -372 2392 -338
rect 2426 -372 2460 -338
rect 2494 -372 2528 -338
rect 2562 -372 2596 -338
rect 2630 -372 2664 -338
rect 2698 -372 2732 -338
rect 2766 -372 2800 -338
rect 3308 -372 3342 -338
rect 3376 -372 3410 -338
rect 3444 -372 3478 -338
rect 3512 -372 3546 -338
rect 3580 -372 3614 -338
rect 3648 -372 3682 -338
rect 3716 -372 3750 -338
rect 3784 -372 3818 -338
rect 4326 -372 4360 -338
rect 4394 -372 4428 -338
rect 4462 -372 4496 -338
rect 4530 -372 4564 -338
rect 4598 -372 4632 -338
rect 4666 -372 4700 -338
rect 4734 -372 4768 -338
rect 4802 -372 4836 -338
<< locali >>
rect -4875 338 -4836 372
rect -4802 338 -4778 372
rect -4734 338 -4706 372
rect -4666 338 -4634 372
rect -4598 338 -4564 372
rect -4528 338 -4496 372
rect -4456 338 -4428 372
rect -4384 338 -4360 372
rect -4326 338 -4287 372
rect -3857 338 -3818 372
rect -3784 338 -3760 372
rect -3716 338 -3688 372
rect -3648 338 -3616 372
rect -3580 338 -3546 372
rect -3510 338 -3478 372
rect -3438 338 -3410 372
rect -3366 338 -3342 372
rect -3308 338 -3269 372
rect -2839 338 -2800 372
rect -2766 338 -2742 372
rect -2698 338 -2670 372
rect -2630 338 -2598 372
rect -2562 338 -2528 372
rect -2492 338 -2460 372
rect -2420 338 -2392 372
rect -2348 338 -2324 372
rect -2290 338 -2251 372
rect -1821 338 -1782 372
rect -1748 338 -1724 372
rect -1680 338 -1652 372
rect -1612 338 -1580 372
rect -1544 338 -1510 372
rect -1474 338 -1442 372
rect -1402 338 -1374 372
rect -1330 338 -1306 372
rect -1272 338 -1233 372
rect -803 338 -764 372
rect -730 338 -706 372
rect -662 338 -634 372
rect -594 338 -562 372
rect -526 338 -492 372
rect -456 338 -424 372
rect -384 338 -356 372
rect -312 338 -288 372
rect -254 338 -215 372
rect 215 338 254 372
rect 288 338 312 372
rect 356 338 384 372
rect 424 338 456 372
rect 492 338 526 372
rect 562 338 594 372
rect 634 338 662 372
rect 706 338 730 372
rect 764 338 803 372
rect 1233 338 1272 372
rect 1306 338 1330 372
rect 1374 338 1402 372
rect 1442 338 1474 372
rect 1510 338 1544 372
rect 1580 338 1612 372
rect 1652 338 1680 372
rect 1724 338 1748 372
rect 1782 338 1821 372
rect 2251 338 2290 372
rect 2324 338 2348 372
rect 2392 338 2420 372
rect 2460 338 2492 372
rect 2528 338 2562 372
rect 2598 338 2630 372
rect 2670 338 2698 372
rect 2742 338 2766 372
rect 2800 338 2839 372
rect 3269 338 3308 372
rect 3342 338 3366 372
rect 3410 338 3438 372
rect 3478 338 3510 372
rect 3546 338 3580 372
rect 3616 338 3648 372
rect 3688 338 3716 372
rect 3760 338 3784 372
rect 3818 338 3857 372
rect 4287 338 4326 372
rect 4360 338 4384 372
rect 4428 338 4456 372
rect 4496 338 4528 372
rect 4564 338 4598 372
rect 4634 338 4666 372
rect 4706 338 4734 372
rect 4778 338 4802 372
rect 4836 338 4875 372
rect -5107 269 -5073 304
rect -5107 197 -5073 221
rect -5107 125 -5073 153
rect -5107 53 -5073 85
rect -5107 -17 -5073 17
rect -5107 -85 -5073 -53
rect -5107 -153 -5073 -125
rect -5107 -221 -5073 -197
rect -5107 -304 -5073 -269
rect -4089 269 -4055 304
rect -4089 197 -4055 221
rect -4089 125 -4055 153
rect -4089 53 -4055 85
rect -4089 -17 -4055 17
rect -4089 -85 -4055 -53
rect -4089 -153 -4055 -125
rect -4089 -221 -4055 -197
rect -4089 -304 -4055 -269
rect -3071 269 -3037 304
rect -3071 197 -3037 221
rect -3071 125 -3037 153
rect -3071 53 -3037 85
rect -3071 -17 -3037 17
rect -3071 -85 -3037 -53
rect -3071 -153 -3037 -125
rect -3071 -221 -3037 -197
rect -3071 -304 -3037 -269
rect -2053 269 -2019 304
rect -2053 197 -2019 221
rect -2053 125 -2019 153
rect -2053 53 -2019 85
rect -2053 -17 -2019 17
rect -2053 -85 -2019 -53
rect -2053 -153 -2019 -125
rect -2053 -221 -2019 -197
rect -2053 -304 -2019 -269
rect -1035 269 -1001 304
rect -1035 197 -1001 221
rect -1035 125 -1001 153
rect -1035 53 -1001 85
rect -1035 -17 -1001 17
rect -1035 -85 -1001 -53
rect -1035 -153 -1001 -125
rect -1035 -221 -1001 -197
rect -1035 -304 -1001 -269
rect -17 269 17 304
rect -17 197 17 221
rect -17 125 17 153
rect -17 53 17 85
rect -17 -17 17 17
rect -17 -85 17 -53
rect -17 -153 17 -125
rect -17 -221 17 -197
rect -17 -304 17 -269
rect 1001 269 1035 304
rect 1001 197 1035 221
rect 1001 125 1035 153
rect 1001 53 1035 85
rect 1001 -17 1035 17
rect 1001 -85 1035 -53
rect 1001 -153 1035 -125
rect 1001 -221 1035 -197
rect 1001 -304 1035 -269
rect 2019 269 2053 304
rect 2019 197 2053 221
rect 2019 125 2053 153
rect 2019 53 2053 85
rect 2019 -17 2053 17
rect 2019 -85 2053 -53
rect 2019 -153 2053 -125
rect 2019 -221 2053 -197
rect 2019 -304 2053 -269
rect 3037 269 3071 304
rect 3037 197 3071 221
rect 3037 125 3071 153
rect 3037 53 3071 85
rect 3037 -17 3071 17
rect 3037 -85 3071 -53
rect 3037 -153 3071 -125
rect 3037 -221 3071 -197
rect 3037 -304 3071 -269
rect 4055 269 4089 304
rect 4055 197 4089 221
rect 4055 125 4089 153
rect 4055 53 4089 85
rect 4055 -17 4089 17
rect 4055 -85 4089 -53
rect 4055 -153 4089 -125
rect 4055 -221 4089 -197
rect 4055 -304 4089 -269
rect 5073 269 5107 304
rect 5073 197 5107 221
rect 5073 125 5107 153
rect 5073 53 5107 85
rect 5073 -17 5107 17
rect 5073 -85 5107 -53
rect 5073 -153 5107 -125
rect 5073 -221 5107 -197
rect 5073 -304 5107 -269
rect -4875 -372 -4836 -338
rect -4802 -372 -4778 -338
rect -4734 -372 -4706 -338
rect -4666 -372 -4634 -338
rect -4598 -372 -4564 -338
rect -4528 -372 -4496 -338
rect -4456 -372 -4428 -338
rect -4384 -372 -4360 -338
rect -4326 -372 -4287 -338
rect -3857 -372 -3818 -338
rect -3784 -372 -3760 -338
rect -3716 -372 -3688 -338
rect -3648 -372 -3616 -338
rect -3580 -372 -3546 -338
rect -3510 -372 -3478 -338
rect -3438 -372 -3410 -338
rect -3366 -372 -3342 -338
rect -3308 -372 -3269 -338
rect -2839 -372 -2800 -338
rect -2766 -372 -2742 -338
rect -2698 -372 -2670 -338
rect -2630 -372 -2598 -338
rect -2562 -372 -2528 -338
rect -2492 -372 -2460 -338
rect -2420 -372 -2392 -338
rect -2348 -372 -2324 -338
rect -2290 -372 -2251 -338
rect -1821 -372 -1782 -338
rect -1748 -372 -1724 -338
rect -1680 -372 -1652 -338
rect -1612 -372 -1580 -338
rect -1544 -372 -1510 -338
rect -1474 -372 -1442 -338
rect -1402 -372 -1374 -338
rect -1330 -372 -1306 -338
rect -1272 -372 -1233 -338
rect -803 -372 -764 -338
rect -730 -372 -706 -338
rect -662 -372 -634 -338
rect -594 -372 -562 -338
rect -526 -372 -492 -338
rect -456 -372 -424 -338
rect -384 -372 -356 -338
rect -312 -372 -288 -338
rect -254 -372 -215 -338
rect 215 -372 254 -338
rect 288 -372 312 -338
rect 356 -372 384 -338
rect 424 -372 456 -338
rect 492 -372 526 -338
rect 562 -372 594 -338
rect 634 -372 662 -338
rect 706 -372 730 -338
rect 764 -372 803 -338
rect 1233 -372 1272 -338
rect 1306 -372 1330 -338
rect 1374 -372 1402 -338
rect 1442 -372 1474 -338
rect 1510 -372 1544 -338
rect 1580 -372 1612 -338
rect 1652 -372 1680 -338
rect 1724 -372 1748 -338
rect 1782 -372 1821 -338
rect 2251 -372 2290 -338
rect 2324 -372 2348 -338
rect 2392 -372 2420 -338
rect 2460 -372 2492 -338
rect 2528 -372 2562 -338
rect 2598 -372 2630 -338
rect 2670 -372 2698 -338
rect 2742 -372 2766 -338
rect 2800 -372 2839 -338
rect 3269 -372 3308 -338
rect 3342 -372 3366 -338
rect 3410 -372 3438 -338
rect 3478 -372 3510 -338
rect 3546 -372 3580 -338
rect 3616 -372 3648 -338
rect 3688 -372 3716 -338
rect 3760 -372 3784 -338
rect 3818 -372 3857 -338
rect 4287 -372 4326 -338
rect 4360 -372 4384 -338
rect 4428 -372 4456 -338
rect 4496 -372 4528 -338
rect 4564 -372 4598 -338
rect 4634 -372 4666 -338
rect 4706 -372 4734 -338
rect 4778 -372 4802 -338
rect 4836 -372 4875 -338
<< viali >>
rect -4778 338 -4768 372
rect -4768 338 -4744 372
rect -4706 338 -4700 372
rect -4700 338 -4672 372
rect -4634 338 -4632 372
rect -4632 338 -4600 372
rect -4562 338 -4530 372
rect -4530 338 -4528 372
rect -4490 338 -4462 372
rect -4462 338 -4456 372
rect -4418 338 -4394 372
rect -4394 338 -4384 372
rect -3760 338 -3750 372
rect -3750 338 -3726 372
rect -3688 338 -3682 372
rect -3682 338 -3654 372
rect -3616 338 -3614 372
rect -3614 338 -3582 372
rect -3544 338 -3512 372
rect -3512 338 -3510 372
rect -3472 338 -3444 372
rect -3444 338 -3438 372
rect -3400 338 -3376 372
rect -3376 338 -3366 372
rect -2742 338 -2732 372
rect -2732 338 -2708 372
rect -2670 338 -2664 372
rect -2664 338 -2636 372
rect -2598 338 -2596 372
rect -2596 338 -2564 372
rect -2526 338 -2494 372
rect -2494 338 -2492 372
rect -2454 338 -2426 372
rect -2426 338 -2420 372
rect -2382 338 -2358 372
rect -2358 338 -2348 372
rect -1724 338 -1714 372
rect -1714 338 -1690 372
rect -1652 338 -1646 372
rect -1646 338 -1618 372
rect -1580 338 -1578 372
rect -1578 338 -1546 372
rect -1508 338 -1476 372
rect -1476 338 -1474 372
rect -1436 338 -1408 372
rect -1408 338 -1402 372
rect -1364 338 -1340 372
rect -1340 338 -1330 372
rect -706 338 -696 372
rect -696 338 -672 372
rect -634 338 -628 372
rect -628 338 -600 372
rect -562 338 -560 372
rect -560 338 -528 372
rect -490 338 -458 372
rect -458 338 -456 372
rect -418 338 -390 372
rect -390 338 -384 372
rect -346 338 -322 372
rect -322 338 -312 372
rect 312 338 322 372
rect 322 338 346 372
rect 384 338 390 372
rect 390 338 418 372
rect 456 338 458 372
rect 458 338 490 372
rect 528 338 560 372
rect 560 338 562 372
rect 600 338 628 372
rect 628 338 634 372
rect 672 338 696 372
rect 696 338 706 372
rect 1330 338 1340 372
rect 1340 338 1364 372
rect 1402 338 1408 372
rect 1408 338 1436 372
rect 1474 338 1476 372
rect 1476 338 1508 372
rect 1546 338 1578 372
rect 1578 338 1580 372
rect 1618 338 1646 372
rect 1646 338 1652 372
rect 1690 338 1714 372
rect 1714 338 1724 372
rect 2348 338 2358 372
rect 2358 338 2382 372
rect 2420 338 2426 372
rect 2426 338 2454 372
rect 2492 338 2494 372
rect 2494 338 2526 372
rect 2564 338 2596 372
rect 2596 338 2598 372
rect 2636 338 2664 372
rect 2664 338 2670 372
rect 2708 338 2732 372
rect 2732 338 2742 372
rect 3366 338 3376 372
rect 3376 338 3400 372
rect 3438 338 3444 372
rect 3444 338 3472 372
rect 3510 338 3512 372
rect 3512 338 3544 372
rect 3582 338 3614 372
rect 3614 338 3616 372
rect 3654 338 3682 372
rect 3682 338 3688 372
rect 3726 338 3750 372
rect 3750 338 3760 372
rect 4384 338 4394 372
rect 4394 338 4418 372
rect 4456 338 4462 372
rect 4462 338 4490 372
rect 4528 338 4530 372
rect 4530 338 4562 372
rect 4600 338 4632 372
rect 4632 338 4634 372
rect 4672 338 4700 372
rect 4700 338 4706 372
rect 4744 338 4768 372
rect 4768 338 4778 372
rect -5107 255 -5073 269
rect -5107 235 -5073 255
rect -5107 187 -5073 197
rect -5107 163 -5073 187
rect -5107 119 -5073 125
rect -5107 91 -5073 119
rect -5107 51 -5073 53
rect -5107 19 -5073 51
rect -5107 -51 -5073 -19
rect -5107 -53 -5073 -51
rect -5107 -119 -5073 -91
rect -5107 -125 -5073 -119
rect -5107 -187 -5073 -163
rect -5107 -197 -5073 -187
rect -5107 -255 -5073 -235
rect -5107 -269 -5073 -255
rect -4089 255 -4055 269
rect -4089 235 -4055 255
rect -4089 187 -4055 197
rect -4089 163 -4055 187
rect -4089 119 -4055 125
rect -4089 91 -4055 119
rect -4089 51 -4055 53
rect -4089 19 -4055 51
rect -4089 -51 -4055 -19
rect -4089 -53 -4055 -51
rect -4089 -119 -4055 -91
rect -4089 -125 -4055 -119
rect -4089 -187 -4055 -163
rect -4089 -197 -4055 -187
rect -4089 -255 -4055 -235
rect -4089 -269 -4055 -255
rect -3071 255 -3037 269
rect -3071 235 -3037 255
rect -3071 187 -3037 197
rect -3071 163 -3037 187
rect -3071 119 -3037 125
rect -3071 91 -3037 119
rect -3071 51 -3037 53
rect -3071 19 -3037 51
rect -3071 -51 -3037 -19
rect -3071 -53 -3037 -51
rect -3071 -119 -3037 -91
rect -3071 -125 -3037 -119
rect -3071 -187 -3037 -163
rect -3071 -197 -3037 -187
rect -3071 -255 -3037 -235
rect -3071 -269 -3037 -255
rect -2053 255 -2019 269
rect -2053 235 -2019 255
rect -2053 187 -2019 197
rect -2053 163 -2019 187
rect -2053 119 -2019 125
rect -2053 91 -2019 119
rect -2053 51 -2019 53
rect -2053 19 -2019 51
rect -2053 -51 -2019 -19
rect -2053 -53 -2019 -51
rect -2053 -119 -2019 -91
rect -2053 -125 -2019 -119
rect -2053 -187 -2019 -163
rect -2053 -197 -2019 -187
rect -2053 -255 -2019 -235
rect -2053 -269 -2019 -255
rect -1035 255 -1001 269
rect -1035 235 -1001 255
rect -1035 187 -1001 197
rect -1035 163 -1001 187
rect -1035 119 -1001 125
rect -1035 91 -1001 119
rect -1035 51 -1001 53
rect -1035 19 -1001 51
rect -1035 -51 -1001 -19
rect -1035 -53 -1001 -51
rect -1035 -119 -1001 -91
rect -1035 -125 -1001 -119
rect -1035 -187 -1001 -163
rect -1035 -197 -1001 -187
rect -1035 -255 -1001 -235
rect -1035 -269 -1001 -255
rect -17 255 17 269
rect -17 235 17 255
rect -17 187 17 197
rect -17 163 17 187
rect -17 119 17 125
rect -17 91 17 119
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect -17 -119 17 -91
rect -17 -125 17 -119
rect -17 -187 17 -163
rect -17 -197 17 -187
rect -17 -255 17 -235
rect -17 -269 17 -255
rect 1001 255 1035 269
rect 1001 235 1035 255
rect 1001 187 1035 197
rect 1001 163 1035 187
rect 1001 119 1035 125
rect 1001 91 1035 119
rect 1001 51 1035 53
rect 1001 19 1035 51
rect 1001 -51 1035 -19
rect 1001 -53 1035 -51
rect 1001 -119 1035 -91
rect 1001 -125 1035 -119
rect 1001 -187 1035 -163
rect 1001 -197 1035 -187
rect 1001 -255 1035 -235
rect 1001 -269 1035 -255
rect 2019 255 2053 269
rect 2019 235 2053 255
rect 2019 187 2053 197
rect 2019 163 2053 187
rect 2019 119 2053 125
rect 2019 91 2053 119
rect 2019 51 2053 53
rect 2019 19 2053 51
rect 2019 -51 2053 -19
rect 2019 -53 2053 -51
rect 2019 -119 2053 -91
rect 2019 -125 2053 -119
rect 2019 -187 2053 -163
rect 2019 -197 2053 -187
rect 2019 -255 2053 -235
rect 2019 -269 2053 -255
rect 3037 255 3071 269
rect 3037 235 3071 255
rect 3037 187 3071 197
rect 3037 163 3071 187
rect 3037 119 3071 125
rect 3037 91 3071 119
rect 3037 51 3071 53
rect 3037 19 3071 51
rect 3037 -51 3071 -19
rect 3037 -53 3071 -51
rect 3037 -119 3071 -91
rect 3037 -125 3071 -119
rect 3037 -187 3071 -163
rect 3037 -197 3071 -187
rect 3037 -255 3071 -235
rect 3037 -269 3071 -255
rect 4055 255 4089 269
rect 4055 235 4089 255
rect 4055 187 4089 197
rect 4055 163 4089 187
rect 4055 119 4089 125
rect 4055 91 4089 119
rect 4055 51 4089 53
rect 4055 19 4089 51
rect 4055 -51 4089 -19
rect 4055 -53 4089 -51
rect 4055 -119 4089 -91
rect 4055 -125 4089 -119
rect 4055 -187 4089 -163
rect 4055 -197 4089 -187
rect 4055 -255 4089 -235
rect 4055 -269 4089 -255
rect 5073 255 5107 269
rect 5073 235 5107 255
rect 5073 187 5107 197
rect 5073 163 5107 187
rect 5073 119 5107 125
rect 5073 91 5107 119
rect 5073 51 5107 53
rect 5073 19 5107 51
rect 5073 -51 5107 -19
rect 5073 -53 5107 -51
rect 5073 -119 5107 -91
rect 5073 -125 5107 -119
rect 5073 -187 5107 -163
rect 5073 -197 5107 -187
rect 5073 -255 5107 -235
rect 5073 -269 5107 -255
rect -4778 -372 -4768 -338
rect -4768 -372 -4744 -338
rect -4706 -372 -4700 -338
rect -4700 -372 -4672 -338
rect -4634 -372 -4632 -338
rect -4632 -372 -4600 -338
rect -4562 -372 -4530 -338
rect -4530 -372 -4528 -338
rect -4490 -372 -4462 -338
rect -4462 -372 -4456 -338
rect -4418 -372 -4394 -338
rect -4394 -372 -4384 -338
rect -3760 -372 -3750 -338
rect -3750 -372 -3726 -338
rect -3688 -372 -3682 -338
rect -3682 -372 -3654 -338
rect -3616 -372 -3614 -338
rect -3614 -372 -3582 -338
rect -3544 -372 -3512 -338
rect -3512 -372 -3510 -338
rect -3472 -372 -3444 -338
rect -3444 -372 -3438 -338
rect -3400 -372 -3376 -338
rect -3376 -372 -3366 -338
rect -2742 -372 -2732 -338
rect -2732 -372 -2708 -338
rect -2670 -372 -2664 -338
rect -2664 -372 -2636 -338
rect -2598 -372 -2596 -338
rect -2596 -372 -2564 -338
rect -2526 -372 -2494 -338
rect -2494 -372 -2492 -338
rect -2454 -372 -2426 -338
rect -2426 -372 -2420 -338
rect -2382 -372 -2358 -338
rect -2358 -372 -2348 -338
rect -1724 -372 -1714 -338
rect -1714 -372 -1690 -338
rect -1652 -372 -1646 -338
rect -1646 -372 -1618 -338
rect -1580 -372 -1578 -338
rect -1578 -372 -1546 -338
rect -1508 -372 -1476 -338
rect -1476 -372 -1474 -338
rect -1436 -372 -1408 -338
rect -1408 -372 -1402 -338
rect -1364 -372 -1340 -338
rect -1340 -372 -1330 -338
rect -706 -372 -696 -338
rect -696 -372 -672 -338
rect -634 -372 -628 -338
rect -628 -372 -600 -338
rect -562 -372 -560 -338
rect -560 -372 -528 -338
rect -490 -372 -458 -338
rect -458 -372 -456 -338
rect -418 -372 -390 -338
rect -390 -372 -384 -338
rect -346 -372 -322 -338
rect -322 -372 -312 -338
rect 312 -372 322 -338
rect 322 -372 346 -338
rect 384 -372 390 -338
rect 390 -372 418 -338
rect 456 -372 458 -338
rect 458 -372 490 -338
rect 528 -372 560 -338
rect 560 -372 562 -338
rect 600 -372 628 -338
rect 628 -372 634 -338
rect 672 -372 696 -338
rect 696 -372 706 -338
rect 1330 -372 1340 -338
rect 1340 -372 1364 -338
rect 1402 -372 1408 -338
rect 1408 -372 1436 -338
rect 1474 -372 1476 -338
rect 1476 -372 1508 -338
rect 1546 -372 1578 -338
rect 1578 -372 1580 -338
rect 1618 -372 1646 -338
rect 1646 -372 1652 -338
rect 1690 -372 1714 -338
rect 1714 -372 1724 -338
rect 2348 -372 2358 -338
rect 2358 -372 2382 -338
rect 2420 -372 2426 -338
rect 2426 -372 2454 -338
rect 2492 -372 2494 -338
rect 2494 -372 2526 -338
rect 2564 -372 2596 -338
rect 2596 -372 2598 -338
rect 2636 -372 2664 -338
rect 2664 -372 2670 -338
rect 2708 -372 2732 -338
rect 2732 -372 2742 -338
rect 3366 -372 3376 -338
rect 3376 -372 3400 -338
rect 3438 -372 3444 -338
rect 3444 -372 3472 -338
rect 3510 -372 3512 -338
rect 3512 -372 3544 -338
rect 3582 -372 3614 -338
rect 3614 -372 3616 -338
rect 3654 -372 3682 -338
rect 3682 -372 3688 -338
rect 3726 -372 3750 -338
rect 3750 -372 3760 -338
rect 4384 -372 4394 -338
rect 4394 -372 4418 -338
rect 4456 -372 4462 -338
rect 4462 -372 4490 -338
rect 4528 -372 4530 -338
rect 4530 -372 4562 -338
rect 4600 -372 4632 -338
rect 4632 -372 4634 -338
rect 4672 -372 4700 -338
rect 4700 -372 4706 -338
rect 4744 -372 4768 -338
rect 4768 -372 4778 -338
<< metal1 >>
rect -4825 372 -4337 378
rect -4825 338 -4778 372
rect -4744 338 -4706 372
rect -4672 338 -4634 372
rect -4600 338 -4562 372
rect -4528 338 -4490 372
rect -4456 338 -4418 372
rect -4384 338 -4337 372
rect -4825 332 -4337 338
rect -3807 372 -3319 378
rect -3807 338 -3760 372
rect -3726 338 -3688 372
rect -3654 338 -3616 372
rect -3582 338 -3544 372
rect -3510 338 -3472 372
rect -3438 338 -3400 372
rect -3366 338 -3319 372
rect -3807 332 -3319 338
rect -2789 372 -2301 378
rect -2789 338 -2742 372
rect -2708 338 -2670 372
rect -2636 338 -2598 372
rect -2564 338 -2526 372
rect -2492 338 -2454 372
rect -2420 338 -2382 372
rect -2348 338 -2301 372
rect -2789 332 -2301 338
rect -1771 372 -1283 378
rect -1771 338 -1724 372
rect -1690 338 -1652 372
rect -1618 338 -1580 372
rect -1546 338 -1508 372
rect -1474 338 -1436 372
rect -1402 338 -1364 372
rect -1330 338 -1283 372
rect -1771 332 -1283 338
rect -753 372 -265 378
rect -753 338 -706 372
rect -672 338 -634 372
rect -600 338 -562 372
rect -528 338 -490 372
rect -456 338 -418 372
rect -384 338 -346 372
rect -312 338 -265 372
rect -753 332 -265 338
rect 265 372 753 378
rect 265 338 312 372
rect 346 338 384 372
rect 418 338 456 372
rect 490 338 528 372
rect 562 338 600 372
rect 634 338 672 372
rect 706 338 753 372
rect 265 332 753 338
rect 1283 372 1771 378
rect 1283 338 1330 372
rect 1364 338 1402 372
rect 1436 338 1474 372
rect 1508 338 1546 372
rect 1580 338 1618 372
rect 1652 338 1690 372
rect 1724 338 1771 372
rect 1283 332 1771 338
rect 2301 372 2789 378
rect 2301 338 2348 372
rect 2382 338 2420 372
rect 2454 338 2492 372
rect 2526 338 2564 372
rect 2598 338 2636 372
rect 2670 338 2708 372
rect 2742 338 2789 372
rect 2301 332 2789 338
rect 3319 372 3807 378
rect 3319 338 3366 372
rect 3400 338 3438 372
rect 3472 338 3510 372
rect 3544 338 3582 372
rect 3616 338 3654 372
rect 3688 338 3726 372
rect 3760 338 3807 372
rect 3319 332 3807 338
rect 4337 372 4825 378
rect 4337 338 4384 372
rect 4418 338 4456 372
rect 4490 338 4528 372
rect 4562 338 4600 372
rect 4634 338 4672 372
rect 4706 338 4744 372
rect 4778 338 4825 372
rect 4337 332 4825 338
rect -5113 269 -5067 300
rect -5113 235 -5107 269
rect -5073 235 -5067 269
rect -5113 197 -5067 235
rect -5113 163 -5107 197
rect -5073 163 -5067 197
rect -5113 125 -5067 163
rect -5113 91 -5107 125
rect -5073 91 -5067 125
rect -5113 53 -5067 91
rect -5113 19 -5107 53
rect -5073 19 -5067 53
rect -5113 -19 -5067 19
rect -5113 -53 -5107 -19
rect -5073 -53 -5067 -19
rect -5113 -91 -5067 -53
rect -5113 -125 -5107 -91
rect -5073 -125 -5067 -91
rect -5113 -163 -5067 -125
rect -5113 -197 -5107 -163
rect -5073 -197 -5067 -163
rect -5113 -235 -5067 -197
rect -5113 -269 -5107 -235
rect -5073 -269 -5067 -235
rect -5113 -300 -5067 -269
rect -4095 269 -4049 300
rect -4095 235 -4089 269
rect -4055 235 -4049 269
rect -4095 197 -4049 235
rect -4095 163 -4089 197
rect -4055 163 -4049 197
rect -4095 125 -4049 163
rect -4095 91 -4089 125
rect -4055 91 -4049 125
rect -4095 53 -4049 91
rect -4095 19 -4089 53
rect -4055 19 -4049 53
rect -4095 -19 -4049 19
rect -4095 -53 -4089 -19
rect -4055 -53 -4049 -19
rect -4095 -91 -4049 -53
rect -4095 -125 -4089 -91
rect -4055 -125 -4049 -91
rect -4095 -163 -4049 -125
rect -4095 -197 -4089 -163
rect -4055 -197 -4049 -163
rect -4095 -235 -4049 -197
rect -4095 -269 -4089 -235
rect -4055 -269 -4049 -235
rect -4095 -300 -4049 -269
rect -3077 269 -3031 300
rect -3077 235 -3071 269
rect -3037 235 -3031 269
rect -3077 197 -3031 235
rect -3077 163 -3071 197
rect -3037 163 -3031 197
rect -3077 125 -3031 163
rect -3077 91 -3071 125
rect -3037 91 -3031 125
rect -3077 53 -3031 91
rect -3077 19 -3071 53
rect -3037 19 -3031 53
rect -3077 -19 -3031 19
rect -3077 -53 -3071 -19
rect -3037 -53 -3031 -19
rect -3077 -91 -3031 -53
rect -3077 -125 -3071 -91
rect -3037 -125 -3031 -91
rect -3077 -163 -3031 -125
rect -3077 -197 -3071 -163
rect -3037 -197 -3031 -163
rect -3077 -235 -3031 -197
rect -3077 -269 -3071 -235
rect -3037 -269 -3031 -235
rect -3077 -300 -3031 -269
rect -2059 269 -2013 300
rect -2059 235 -2053 269
rect -2019 235 -2013 269
rect -2059 197 -2013 235
rect -2059 163 -2053 197
rect -2019 163 -2013 197
rect -2059 125 -2013 163
rect -2059 91 -2053 125
rect -2019 91 -2013 125
rect -2059 53 -2013 91
rect -2059 19 -2053 53
rect -2019 19 -2013 53
rect -2059 -19 -2013 19
rect -2059 -53 -2053 -19
rect -2019 -53 -2013 -19
rect -2059 -91 -2013 -53
rect -2059 -125 -2053 -91
rect -2019 -125 -2013 -91
rect -2059 -163 -2013 -125
rect -2059 -197 -2053 -163
rect -2019 -197 -2013 -163
rect -2059 -235 -2013 -197
rect -2059 -269 -2053 -235
rect -2019 -269 -2013 -235
rect -2059 -300 -2013 -269
rect -1041 269 -995 300
rect -1041 235 -1035 269
rect -1001 235 -995 269
rect -1041 197 -995 235
rect -1041 163 -1035 197
rect -1001 163 -995 197
rect -1041 125 -995 163
rect -1041 91 -1035 125
rect -1001 91 -995 125
rect -1041 53 -995 91
rect -1041 19 -1035 53
rect -1001 19 -995 53
rect -1041 -19 -995 19
rect -1041 -53 -1035 -19
rect -1001 -53 -995 -19
rect -1041 -91 -995 -53
rect -1041 -125 -1035 -91
rect -1001 -125 -995 -91
rect -1041 -163 -995 -125
rect -1041 -197 -1035 -163
rect -1001 -197 -995 -163
rect -1041 -235 -995 -197
rect -1041 -269 -1035 -235
rect -1001 -269 -995 -235
rect -1041 -300 -995 -269
rect -23 269 23 300
rect -23 235 -17 269
rect 17 235 23 269
rect -23 197 23 235
rect -23 163 -17 197
rect 17 163 23 197
rect -23 125 23 163
rect -23 91 -17 125
rect 17 91 23 125
rect -23 53 23 91
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -91 23 -53
rect -23 -125 -17 -91
rect 17 -125 23 -91
rect -23 -163 23 -125
rect -23 -197 -17 -163
rect 17 -197 23 -163
rect -23 -235 23 -197
rect -23 -269 -17 -235
rect 17 -269 23 -235
rect -23 -300 23 -269
rect 995 269 1041 300
rect 995 235 1001 269
rect 1035 235 1041 269
rect 995 197 1041 235
rect 995 163 1001 197
rect 1035 163 1041 197
rect 995 125 1041 163
rect 995 91 1001 125
rect 1035 91 1041 125
rect 995 53 1041 91
rect 995 19 1001 53
rect 1035 19 1041 53
rect 995 -19 1041 19
rect 995 -53 1001 -19
rect 1035 -53 1041 -19
rect 995 -91 1041 -53
rect 995 -125 1001 -91
rect 1035 -125 1041 -91
rect 995 -163 1041 -125
rect 995 -197 1001 -163
rect 1035 -197 1041 -163
rect 995 -235 1041 -197
rect 995 -269 1001 -235
rect 1035 -269 1041 -235
rect 995 -300 1041 -269
rect 2013 269 2059 300
rect 2013 235 2019 269
rect 2053 235 2059 269
rect 2013 197 2059 235
rect 2013 163 2019 197
rect 2053 163 2059 197
rect 2013 125 2059 163
rect 2013 91 2019 125
rect 2053 91 2059 125
rect 2013 53 2059 91
rect 2013 19 2019 53
rect 2053 19 2059 53
rect 2013 -19 2059 19
rect 2013 -53 2019 -19
rect 2053 -53 2059 -19
rect 2013 -91 2059 -53
rect 2013 -125 2019 -91
rect 2053 -125 2059 -91
rect 2013 -163 2059 -125
rect 2013 -197 2019 -163
rect 2053 -197 2059 -163
rect 2013 -235 2059 -197
rect 2013 -269 2019 -235
rect 2053 -269 2059 -235
rect 2013 -300 2059 -269
rect 3031 269 3077 300
rect 3031 235 3037 269
rect 3071 235 3077 269
rect 3031 197 3077 235
rect 3031 163 3037 197
rect 3071 163 3077 197
rect 3031 125 3077 163
rect 3031 91 3037 125
rect 3071 91 3077 125
rect 3031 53 3077 91
rect 3031 19 3037 53
rect 3071 19 3077 53
rect 3031 -19 3077 19
rect 3031 -53 3037 -19
rect 3071 -53 3077 -19
rect 3031 -91 3077 -53
rect 3031 -125 3037 -91
rect 3071 -125 3077 -91
rect 3031 -163 3077 -125
rect 3031 -197 3037 -163
rect 3071 -197 3077 -163
rect 3031 -235 3077 -197
rect 3031 -269 3037 -235
rect 3071 -269 3077 -235
rect 3031 -300 3077 -269
rect 4049 269 4095 300
rect 4049 235 4055 269
rect 4089 235 4095 269
rect 4049 197 4095 235
rect 4049 163 4055 197
rect 4089 163 4095 197
rect 4049 125 4095 163
rect 4049 91 4055 125
rect 4089 91 4095 125
rect 4049 53 4095 91
rect 4049 19 4055 53
rect 4089 19 4095 53
rect 4049 -19 4095 19
rect 4049 -53 4055 -19
rect 4089 -53 4095 -19
rect 4049 -91 4095 -53
rect 4049 -125 4055 -91
rect 4089 -125 4095 -91
rect 4049 -163 4095 -125
rect 4049 -197 4055 -163
rect 4089 -197 4095 -163
rect 4049 -235 4095 -197
rect 4049 -269 4055 -235
rect 4089 -269 4095 -235
rect 4049 -300 4095 -269
rect 5067 269 5113 300
rect 5067 235 5073 269
rect 5107 235 5113 269
rect 5067 197 5113 235
rect 5067 163 5073 197
rect 5107 163 5113 197
rect 5067 125 5113 163
rect 5067 91 5073 125
rect 5107 91 5113 125
rect 5067 53 5113 91
rect 5067 19 5073 53
rect 5107 19 5113 53
rect 5067 -19 5113 19
rect 5067 -53 5073 -19
rect 5107 -53 5113 -19
rect 5067 -91 5113 -53
rect 5067 -125 5073 -91
rect 5107 -125 5113 -91
rect 5067 -163 5113 -125
rect 5067 -197 5073 -163
rect 5107 -197 5113 -163
rect 5067 -235 5113 -197
rect 5067 -269 5073 -235
rect 5107 -269 5113 -235
rect 5067 -300 5113 -269
rect -4825 -338 -4337 -332
rect -4825 -372 -4778 -338
rect -4744 -372 -4706 -338
rect -4672 -372 -4634 -338
rect -4600 -372 -4562 -338
rect -4528 -372 -4490 -338
rect -4456 -372 -4418 -338
rect -4384 -372 -4337 -338
rect -4825 -378 -4337 -372
rect -3807 -338 -3319 -332
rect -3807 -372 -3760 -338
rect -3726 -372 -3688 -338
rect -3654 -372 -3616 -338
rect -3582 -372 -3544 -338
rect -3510 -372 -3472 -338
rect -3438 -372 -3400 -338
rect -3366 -372 -3319 -338
rect -3807 -378 -3319 -372
rect -2789 -338 -2301 -332
rect -2789 -372 -2742 -338
rect -2708 -372 -2670 -338
rect -2636 -372 -2598 -338
rect -2564 -372 -2526 -338
rect -2492 -372 -2454 -338
rect -2420 -372 -2382 -338
rect -2348 -372 -2301 -338
rect -2789 -378 -2301 -372
rect -1771 -338 -1283 -332
rect -1771 -372 -1724 -338
rect -1690 -372 -1652 -338
rect -1618 -372 -1580 -338
rect -1546 -372 -1508 -338
rect -1474 -372 -1436 -338
rect -1402 -372 -1364 -338
rect -1330 -372 -1283 -338
rect -1771 -378 -1283 -372
rect -753 -338 -265 -332
rect -753 -372 -706 -338
rect -672 -372 -634 -338
rect -600 -372 -562 -338
rect -528 -372 -490 -338
rect -456 -372 -418 -338
rect -384 -372 -346 -338
rect -312 -372 -265 -338
rect -753 -378 -265 -372
rect 265 -338 753 -332
rect 265 -372 312 -338
rect 346 -372 384 -338
rect 418 -372 456 -338
rect 490 -372 528 -338
rect 562 -372 600 -338
rect 634 -372 672 -338
rect 706 -372 753 -338
rect 265 -378 753 -372
rect 1283 -338 1771 -332
rect 1283 -372 1330 -338
rect 1364 -372 1402 -338
rect 1436 -372 1474 -338
rect 1508 -372 1546 -338
rect 1580 -372 1618 -338
rect 1652 -372 1690 -338
rect 1724 -372 1771 -338
rect 1283 -378 1771 -372
rect 2301 -338 2789 -332
rect 2301 -372 2348 -338
rect 2382 -372 2420 -338
rect 2454 -372 2492 -338
rect 2526 -372 2564 -338
rect 2598 -372 2636 -338
rect 2670 -372 2708 -338
rect 2742 -372 2789 -338
rect 2301 -378 2789 -372
rect 3319 -338 3807 -332
rect 3319 -372 3366 -338
rect 3400 -372 3438 -338
rect 3472 -372 3510 -338
rect 3544 -372 3582 -338
rect 3616 -372 3654 -338
rect 3688 -372 3726 -338
rect 3760 -372 3807 -338
rect 3319 -378 3807 -372
rect 4337 -338 4825 -332
rect 4337 -372 4384 -338
rect 4418 -372 4456 -338
rect 4490 -372 4528 -338
rect 4562 -372 4600 -338
rect 4634 -372 4672 -338
rect 4706 -372 4744 -338
rect 4778 -372 4825 -338
rect 4337 -378 4825 -372
<< end >>
