magic
tech sky130A
magscale 1 2
timestamp 1621211034
<< nmos >>
rect -10151 109 -9191 709
rect -9133 109 -8173 709
rect -8115 109 -7155 709
rect -7097 109 -6137 709
rect -6079 109 -5119 709
rect -5061 109 -4101 709
rect -4043 109 -3083 709
rect -3025 109 -2065 709
rect -2007 109 -1047 709
rect -989 109 -29 709
rect 29 109 989 709
rect 1047 109 2007 709
rect 2065 109 3025 709
rect 3083 109 4043 709
rect 4101 109 5061 709
rect 5119 109 6079 709
rect 6137 109 7097 709
rect 7155 109 8115 709
rect 8173 109 9133 709
rect 9191 109 10151 709
rect -10151 -709 -9191 -109
rect -9133 -709 -8173 -109
rect -8115 -709 -7155 -109
rect -7097 -709 -6137 -109
rect -6079 -709 -5119 -109
rect -5061 -709 -4101 -109
rect -4043 -709 -3083 -109
rect -3025 -709 -2065 -109
rect -2007 -709 -1047 -109
rect -989 -709 -29 -109
rect 29 -709 989 -109
rect 1047 -709 2007 -109
rect 2065 -709 3025 -109
rect 3083 -709 4043 -109
rect 4101 -709 5061 -109
rect 5119 -709 6079 -109
rect 6137 -709 7097 -109
rect 7155 -709 8115 -109
rect 8173 -709 9133 -109
rect 9191 -709 10151 -109
<< ndiff >>
rect -10209 697 -10151 709
rect -10209 121 -10197 697
rect -10163 121 -10151 697
rect -10209 109 -10151 121
rect -9191 697 -9133 709
rect -9191 121 -9179 697
rect -9145 121 -9133 697
rect -9191 109 -9133 121
rect -8173 697 -8115 709
rect -8173 121 -8161 697
rect -8127 121 -8115 697
rect -8173 109 -8115 121
rect -7155 697 -7097 709
rect -7155 121 -7143 697
rect -7109 121 -7097 697
rect -7155 109 -7097 121
rect -6137 697 -6079 709
rect -6137 121 -6125 697
rect -6091 121 -6079 697
rect -6137 109 -6079 121
rect -5119 697 -5061 709
rect -5119 121 -5107 697
rect -5073 121 -5061 697
rect -5119 109 -5061 121
rect -4101 697 -4043 709
rect -4101 121 -4089 697
rect -4055 121 -4043 697
rect -4101 109 -4043 121
rect -3083 697 -3025 709
rect -3083 121 -3071 697
rect -3037 121 -3025 697
rect -3083 109 -3025 121
rect -2065 697 -2007 709
rect -2065 121 -2053 697
rect -2019 121 -2007 697
rect -2065 109 -2007 121
rect -1047 697 -989 709
rect -1047 121 -1035 697
rect -1001 121 -989 697
rect -1047 109 -989 121
rect -29 697 29 709
rect -29 121 -17 697
rect 17 121 29 697
rect -29 109 29 121
rect 989 697 1047 709
rect 989 121 1001 697
rect 1035 121 1047 697
rect 989 109 1047 121
rect 2007 697 2065 709
rect 2007 121 2019 697
rect 2053 121 2065 697
rect 2007 109 2065 121
rect 3025 697 3083 709
rect 3025 121 3037 697
rect 3071 121 3083 697
rect 3025 109 3083 121
rect 4043 697 4101 709
rect 4043 121 4055 697
rect 4089 121 4101 697
rect 4043 109 4101 121
rect 5061 697 5119 709
rect 5061 121 5073 697
rect 5107 121 5119 697
rect 5061 109 5119 121
rect 6079 697 6137 709
rect 6079 121 6091 697
rect 6125 121 6137 697
rect 6079 109 6137 121
rect 7097 697 7155 709
rect 7097 121 7109 697
rect 7143 121 7155 697
rect 7097 109 7155 121
rect 8115 697 8173 709
rect 8115 121 8127 697
rect 8161 121 8173 697
rect 8115 109 8173 121
rect 9133 697 9191 709
rect 9133 121 9145 697
rect 9179 121 9191 697
rect 9133 109 9191 121
rect 10151 697 10209 709
rect 10151 121 10163 697
rect 10197 121 10209 697
rect 10151 109 10209 121
rect -10209 -121 -10151 -109
rect -10209 -697 -10197 -121
rect -10163 -697 -10151 -121
rect -10209 -709 -10151 -697
rect -9191 -121 -9133 -109
rect -9191 -697 -9179 -121
rect -9145 -697 -9133 -121
rect -9191 -709 -9133 -697
rect -8173 -121 -8115 -109
rect -8173 -697 -8161 -121
rect -8127 -697 -8115 -121
rect -8173 -709 -8115 -697
rect -7155 -121 -7097 -109
rect -7155 -697 -7143 -121
rect -7109 -697 -7097 -121
rect -7155 -709 -7097 -697
rect -6137 -121 -6079 -109
rect -6137 -697 -6125 -121
rect -6091 -697 -6079 -121
rect -6137 -709 -6079 -697
rect -5119 -121 -5061 -109
rect -5119 -697 -5107 -121
rect -5073 -697 -5061 -121
rect -5119 -709 -5061 -697
rect -4101 -121 -4043 -109
rect -4101 -697 -4089 -121
rect -4055 -697 -4043 -121
rect -4101 -709 -4043 -697
rect -3083 -121 -3025 -109
rect -3083 -697 -3071 -121
rect -3037 -697 -3025 -121
rect -3083 -709 -3025 -697
rect -2065 -121 -2007 -109
rect -2065 -697 -2053 -121
rect -2019 -697 -2007 -121
rect -2065 -709 -2007 -697
rect -1047 -121 -989 -109
rect -1047 -697 -1035 -121
rect -1001 -697 -989 -121
rect -1047 -709 -989 -697
rect -29 -121 29 -109
rect -29 -697 -17 -121
rect 17 -697 29 -121
rect -29 -709 29 -697
rect 989 -121 1047 -109
rect 989 -697 1001 -121
rect 1035 -697 1047 -121
rect 989 -709 1047 -697
rect 2007 -121 2065 -109
rect 2007 -697 2019 -121
rect 2053 -697 2065 -121
rect 2007 -709 2065 -697
rect 3025 -121 3083 -109
rect 3025 -697 3037 -121
rect 3071 -697 3083 -121
rect 3025 -709 3083 -697
rect 4043 -121 4101 -109
rect 4043 -697 4055 -121
rect 4089 -697 4101 -121
rect 4043 -709 4101 -697
rect 5061 -121 5119 -109
rect 5061 -697 5073 -121
rect 5107 -697 5119 -121
rect 5061 -709 5119 -697
rect 6079 -121 6137 -109
rect 6079 -697 6091 -121
rect 6125 -697 6137 -121
rect 6079 -709 6137 -697
rect 7097 -121 7155 -109
rect 7097 -697 7109 -121
rect 7143 -697 7155 -121
rect 7097 -709 7155 -697
rect 8115 -121 8173 -109
rect 8115 -697 8127 -121
rect 8161 -697 8173 -121
rect 8115 -709 8173 -697
rect 9133 -121 9191 -109
rect 9133 -697 9145 -121
rect 9179 -697 9191 -121
rect 9133 -709 9191 -697
rect 10151 -121 10209 -109
rect 10151 -697 10163 -121
rect 10197 -697 10209 -121
rect 10151 -709 10209 -697
<< ndiffc >>
rect -10197 121 -10163 697
rect -9179 121 -9145 697
rect -8161 121 -8127 697
rect -7143 121 -7109 697
rect -6125 121 -6091 697
rect -5107 121 -5073 697
rect -4089 121 -4055 697
rect -3071 121 -3037 697
rect -2053 121 -2019 697
rect -1035 121 -1001 697
rect -17 121 17 697
rect 1001 121 1035 697
rect 2019 121 2053 697
rect 3037 121 3071 697
rect 4055 121 4089 697
rect 5073 121 5107 697
rect 6091 121 6125 697
rect 7109 121 7143 697
rect 8127 121 8161 697
rect 9145 121 9179 697
rect 10163 121 10197 697
rect -10197 -697 -10163 -121
rect -9179 -697 -9145 -121
rect -8161 -697 -8127 -121
rect -7143 -697 -7109 -121
rect -6125 -697 -6091 -121
rect -5107 -697 -5073 -121
rect -4089 -697 -4055 -121
rect -3071 -697 -3037 -121
rect -2053 -697 -2019 -121
rect -1035 -697 -1001 -121
rect -17 -697 17 -121
rect 1001 -697 1035 -121
rect 2019 -697 2053 -121
rect 3037 -697 3071 -121
rect 4055 -697 4089 -121
rect 5073 -697 5107 -121
rect 6091 -697 6125 -121
rect 7109 -697 7143 -121
rect 8127 -697 8161 -121
rect 9145 -697 9179 -121
rect 10163 -697 10197 -121
<< poly >>
rect -9965 781 -9377 797
rect -9965 764 -9949 781
rect -10151 747 -9949 764
rect -9393 764 -9377 781
rect -8947 781 -8359 797
rect -8947 764 -8931 781
rect -9393 747 -9191 764
rect -10151 709 -9191 747
rect -9133 747 -8931 764
rect -8375 764 -8359 781
rect -7929 781 -7341 797
rect -7929 764 -7913 781
rect -8375 747 -8173 764
rect -9133 709 -8173 747
rect -8115 747 -7913 764
rect -7357 764 -7341 781
rect -6911 781 -6323 797
rect -6911 764 -6895 781
rect -7357 747 -7155 764
rect -8115 709 -7155 747
rect -7097 747 -6895 764
rect -6339 764 -6323 781
rect -5893 781 -5305 797
rect -5893 764 -5877 781
rect -6339 747 -6137 764
rect -7097 709 -6137 747
rect -6079 747 -5877 764
rect -5321 764 -5305 781
rect -4875 781 -4287 797
rect -4875 764 -4859 781
rect -5321 747 -5119 764
rect -6079 709 -5119 747
rect -5061 747 -4859 764
rect -4303 764 -4287 781
rect -3857 781 -3269 797
rect -3857 764 -3841 781
rect -4303 747 -4101 764
rect -5061 709 -4101 747
rect -4043 747 -3841 764
rect -3285 764 -3269 781
rect -2839 781 -2251 797
rect -2839 764 -2823 781
rect -3285 747 -3083 764
rect -4043 709 -3083 747
rect -3025 747 -2823 764
rect -2267 764 -2251 781
rect -1821 781 -1233 797
rect -1821 764 -1805 781
rect -2267 747 -2065 764
rect -3025 709 -2065 747
rect -2007 747 -1805 764
rect -1249 764 -1233 781
rect -803 781 -215 797
rect -803 764 -787 781
rect -1249 747 -1047 764
rect -2007 709 -1047 747
rect -989 747 -787 764
rect -231 764 -215 781
rect 215 781 803 797
rect 215 764 231 781
rect -231 747 -29 764
rect -989 709 -29 747
rect 29 747 231 764
rect 787 764 803 781
rect 1233 781 1821 797
rect 1233 764 1249 781
rect 787 747 989 764
rect 29 709 989 747
rect 1047 747 1249 764
rect 1805 764 1821 781
rect 2251 781 2839 797
rect 2251 764 2267 781
rect 1805 747 2007 764
rect 1047 709 2007 747
rect 2065 747 2267 764
rect 2823 764 2839 781
rect 3269 781 3857 797
rect 3269 764 3285 781
rect 2823 747 3025 764
rect 2065 709 3025 747
rect 3083 747 3285 764
rect 3841 764 3857 781
rect 4287 781 4875 797
rect 4287 764 4303 781
rect 3841 747 4043 764
rect 3083 709 4043 747
rect 4101 747 4303 764
rect 4859 764 4875 781
rect 5305 781 5893 797
rect 5305 764 5321 781
rect 4859 747 5061 764
rect 4101 709 5061 747
rect 5119 747 5321 764
rect 5877 764 5893 781
rect 6323 781 6911 797
rect 6323 764 6339 781
rect 5877 747 6079 764
rect 5119 709 6079 747
rect 6137 747 6339 764
rect 6895 764 6911 781
rect 7341 781 7929 797
rect 7341 764 7357 781
rect 6895 747 7097 764
rect 6137 709 7097 747
rect 7155 747 7357 764
rect 7913 764 7929 781
rect 8359 781 8947 797
rect 8359 764 8375 781
rect 7913 747 8115 764
rect 7155 709 8115 747
rect 8173 747 8375 764
rect 8931 764 8947 781
rect 9377 781 9965 797
rect 9377 764 9393 781
rect 8931 747 9133 764
rect 8173 709 9133 747
rect 9191 747 9393 764
rect 9949 764 9965 781
rect 9949 747 10151 764
rect 9191 709 10151 747
rect -10151 71 -9191 109
rect -10151 54 -9949 71
rect -9965 37 -9949 54
rect -9393 54 -9191 71
rect -9133 71 -8173 109
rect -9133 54 -8931 71
rect -9393 37 -9377 54
rect -9965 21 -9377 37
rect -8947 37 -8931 54
rect -8375 54 -8173 71
rect -8115 71 -7155 109
rect -8115 54 -7913 71
rect -8375 37 -8359 54
rect -8947 21 -8359 37
rect -7929 37 -7913 54
rect -7357 54 -7155 71
rect -7097 71 -6137 109
rect -7097 54 -6895 71
rect -7357 37 -7341 54
rect -7929 21 -7341 37
rect -6911 37 -6895 54
rect -6339 54 -6137 71
rect -6079 71 -5119 109
rect -6079 54 -5877 71
rect -6339 37 -6323 54
rect -6911 21 -6323 37
rect -5893 37 -5877 54
rect -5321 54 -5119 71
rect -5061 71 -4101 109
rect -5061 54 -4859 71
rect -5321 37 -5305 54
rect -5893 21 -5305 37
rect -4875 37 -4859 54
rect -4303 54 -4101 71
rect -4043 71 -3083 109
rect -4043 54 -3841 71
rect -4303 37 -4287 54
rect -4875 21 -4287 37
rect -3857 37 -3841 54
rect -3285 54 -3083 71
rect -3025 71 -2065 109
rect -3025 54 -2823 71
rect -3285 37 -3269 54
rect -3857 21 -3269 37
rect -2839 37 -2823 54
rect -2267 54 -2065 71
rect -2007 71 -1047 109
rect -2007 54 -1805 71
rect -2267 37 -2251 54
rect -2839 21 -2251 37
rect -1821 37 -1805 54
rect -1249 54 -1047 71
rect -989 71 -29 109
rect -989 54 -787 71
rect -1249 37 -1233 54
rect -1821 21 -1233 37
rect -803 37 -787 54
rect -231 54 -29 71
rect 29 71 989 109
rect 29 54 231 71
rect -231 37 -215 54
rect -803 21 -215 37
rect 215 37 231 54
rect 787 54 989 71
rect 1047 71 2007 109
rect 1047 54 1249 71
rect 787 37 803 54
rect 215 21 803 37
rect 1233 37 1249 54
rect 1805 54 2007 71
rect 2065 71 3025 109
rect 2065 54 2267 71
rect 1805 37 1821 54
rect 1233 21 1821 37
rect 2251 37 2267 54
rect 2823 54 3025 71
rect 3083 71 4043 109
rect 3083 54 3285 71
rect 2823 37 2839 54
rect 2251 21 2839 37
rect 3269 37 3285 54
rect 3841 54 4043 71
rect 4101 71 5061 109
rect 4101 54 4303 71
rect 3841 37 3857 54
rect 3269 21 3857 37
rect 4287 37 4303 54
rect 4859 54 5061 71
rect 5119 71 6079 109
rect 5119 54 5321 71
rect 4859 37 4875 54
rect 4287 21 4875 37
rect 5305 37 5321 54
rect 5877 54 6079 71
rect 6137 71 7097 109
rect 6137 54 6339 71
rect 5877 37 5893 54
rect 5305 21 5893 37
rect 6323 37 6339 54
rect 6895 54 7097 71
rect 7155 71 8115 109
rect 7155 54 7357 71
rect 6895 37 6911 54
rect 6323 21 6911 37
rect 7341 37 7357 54
rect 7913 54 8115 71
rect 8173 71 9133 109
rect 8173 54 8375 71
rect 7913 37 7929 54
rect 7341 21 7929 37
rect 8359 37 8375 54
rect 8931 54 9133 71
rect 9191 71 10151 109
rect 9191 54 9393 71
rect 8931 37 8947 54
rect 8359 21 8947 37
rect 9377 37 9393 54
rect 9949 54 10151 71
rect 9949 37 9965 54
rect 9377 21 9965 37
rect -9965 -37 -9377 -21
rect -9965 -54 -9949 -37
rect -10151 -71 -9949 -54
rect -9393 -54 -9377 -37
rect -8947 -37 -8359 -21
rect -8947 -54 -8931 -37
rect -9393 -71 -9191 -54
rect -10151 -109 -9191 -71
rect -9133 -71 -8931 -54
rect -8375 -54 -8359 -37
rect -7929 -37 -7341 -21
rect -7929 -54 -7913 -37
rect -8375 -71 -8173 -54
rect -9133 -109 -8173 -71
rect -8115 -71 -7913 -54
rect -7357 -54 -7341 -37
rect -6911 -37 -6323 -21
rect -6911 -54 -6895 -37
rect -7357 -71 -7155 -54
rect -8115 -109 -7155 -71
rect -7097 -71 -6895 -54
rect -6339 -54 -6323 -37
rect -5893 -37 -5305 -21
rect -5893 -54 -5877 -37
rect -6339 -71 -6137 -54
rect -7097 -109 -6137 -71
rect -6079 -71 -5877 -54
rect -5321 -54 -5305 -37
rect -4875 -37 -4287 -21
rect -4875 -54 -4859 -37
rect -5321 -71 -5119 -54
rect -6079 -109 -5119 -71
rect -5061 -71 -4859 -54
rect -4303 -54 -4287 -37
rect -3857 -37 -3269 -21
rect -3857 -54 -3841 -37
rect -4303 -71 -4101 -54
rect -5061 -109 -4101 -71
rect -4043 -71 -3841 -54
rect -3285 -54 -3269 -37
rect -2839 -37 -2251 -21
rect -2839 -54 -2823 -37
rect -3285 -71 -3083 -54
rect -4043 -109 -3083 -71
rect -3025 -71 -2823 -54
rect -2267 -54 -2251 -37
rect -1821 -37 -1233 -21
rect -1821 -54 -1805 -37
rect -2267 -71 -2065 -54
rect -3025 -109 -2065 -71
rect -2007 -71 -1805 -54
rect -1249 -54 -1233 -37
rect -803 -37 -215 -21
rect -803 -54 -787 -37
rect -1249 -71 -1047 -54
rect -2007 -109 -1047 -71
rect -989 -71 -787 -54
rect -231 -54 -215 -37
rect 215 -37 803 -21
rect 215 -54 231 -37
rect -231 -71 -29 -54
rect -989 -109 -29 -71
rect 29 -71 231 -54
rect 787 -54 803 -37
rect 1233 -37 1821 -21
rect 1233 -54 1249 -37
rect 787 -71 989 -54
rect 29 -109 989 -71
rect 1047 -71 1249 -54
rect 1805 -54 1821 -37
rect 2251 -37 2839 -21
rect 2251 -54 2267 -37
rect 1805 -71 2007 -54
rect 1047 -109 2007 -71
rect 2065 -71 2267 -54
rect 2823 -54 2839 -37
rect 3269 -37 3857 -21
rect 3269 -54 3285 -37
rect 2823 -71 3025 -54
rect 2065 -109 3025 -71
rect 3083 -71 3285 -54
rect 3841 -54 3857 -37
rect 4287 -37 4875 -21
rect 4287 -54 4303 -37
rect 3841 -71 4043 -54
rect 3083 -109 4043 -71
rect 4101 -71 4303 -54
rect 4859 -54 4875 -37
rect 5305 -37 5893 -21
rect 5305 -54 5321 -37
rect 4859 -71 5061 -54
rect 4101 -109 5061 -71
rect 5119 -71 5321 -54
rect 5877 -54 5893 -37
rect 6323 -37 6911 -21
rect 6323 -54 6339 -37
rect 5877 -71 6079 -54
rect 5119 -109 6079 -71
rect 6137 -71 6339 -54
rect 6895 -54 6911 -37
rect 7341 -37 7929 -21
rect 7341 -54 7357 -37
rect 6895 -71 7097 -54
rect 6137 -109 7097 -71
rect 7155 -71 7357 -54
rect 7913 -54 7929 -37
rect 8359 -37 8947 -21
rect 8359 -54 8375 -37
rect 7913 -71 8115 -54
rect 7155 -109 8115 -71
rect 8173 -71 8375 -54
rect 8931 -54 8947 -37
rect 9377 -37 9965 -21
rect 9377 -54 9393 -37
rect 8931 -71 9133 -54
rect 8173 -109 9133 -71
rect 9191 -71 9393 -54
rect 9949 -54 9965 -37
rect 9949 -71 10151 -54
rect 9191 -109 10151 -71
rect -10151 -747 -9191 -709
rect -10151 -764 -9949 -747
rect -9965 -781 -9949 -764
rect -9393 -764 -9191 -747
rect -9133 -747 -8173 -709
rect -9133 -764 -8931 -747
rect -9393 -781 -9377 -764
rect -9965 -797 -9377 -781
rect -8947 -781 -8931 -764
rect -8375 -764 -8173 -747
rect -8115 -747 -7155 -709
rect -8115 -764 -7913 -747
rect -8375 -781 -8359 -764
rect -8947 -797 -8359 -781
rect -7929 -781 -7913 -764
rect -7357 -764 -7155 -747
rect -7097 -747 -6137 -709
rect -7097 -764 -6895 -747
rect -7357 -781 -7341 -764
rect -7929 -797 -7341 -781
rect -6911 -781 -6895 -764
rect -6339 -764 -6137 -747
rect -6079 -747 -5119 -709
rect -6079 -764 -5877 -747
rect -6339 -781 -6323 -764
rect -6911 -797 -6323 -781
rect -5893 -781 -5877 -764
rect -5321 -764 -5119 -747
rect -5061 -747 -4101 -709
rect -5061 -764 -4859 -747
rect -5321 -781 -5305 -764
rect -5893 -797 -5305 -781
rect -4875 -781 -4859 -764
rect -4303 -764 -4101 -747
rect -4043 -747 -3083 -709
rect -4043 -764 -3841 -747
rect -4303 -781 -4287 -764
rect -4875 -797 -4287 -781
rect -3857 -781 -3841 -764
rect -3285 -764 -3083 -747
rect -3025 -747 -2065 -709
rect -3025 -764 -2823 -747
rect -3285 -781 -3269 -764
rect -3857 -797 -3269 -781
rect -2839 -781 -2823 -764
rect -2267 -764 -2065 -747
rect -2007 -747 -1047 -709
rect -2007 -764 -1805 -747
rect -2267 -781 -2251 -764
rect -2839 -797 -2251 -781
rect -1821 -781 -1805 -764
rect -1249 -764 -1047 -747
rect -989 -747 -29 -709
rect -989 -764 -787 -747
rect -1249 -781 -1233 -764
rect -1821 -797 -1233 -781
rect -803 -781 -787 -764
rect -231 -764 -29 -747
rect 29 -747 989 -709
rect 29 -764 231 -747
rect -231 -781 -215 -764
rect -803 -797 -215 -781
rect 215 -781 231 -764
rect 787 -764 989 -747
rect 1047 -747 2007 -709
rect 1047 -764 1249 -747
rect 787 -781 803 -764
rect 215 -797 803 -781
rect 1233 -781 1249 -764
rect 1805 -764 2007 -747
rect 2065 -747 3025 -709
rect 2065 -764 2267 -747
rect 1805 -781 1821 -764
rect 1233 -797 1821 -781
rect 2251 -781 2267 -764
rect 2823 -764 3025 -747
rect 3083 -747 4043 -709
rect 3083 -764 3285 -747
rect 2823 -781 2839 -764
rect 2251 -797 2839 -781
rect 3269 -781 3285 -764
rect 3841 -764 4043 -747
rect 4101 -747 5061 -709
rect 4101 -764 4303 -747
rect 3841 -781 3857 -764
rect 3269 -797 3857 -781
rect 4287 -781 4303 -764
rect 4859 -764 5061 -747
rect 5119 -747 6079 -709
rect 5119 -764 5321 -747
rect 4859 -781 4875 -764
rect 4287 -797 4875 -781
rect 5305 -781 5321 -764
rect 5877 -764 6079 -747
rect 6137 -747 7097 -709
rect 6137 -764 6339 -747
rect 5877 -781 5893 -764
rect 5305 -797 5893 -781
rect 6323 -781 6339 -764
rect 6895 -764 7097 -747
rect 7155 -747 8115 -709
rect 7155 -764 7357 -747
rect 6895 -781 6911 -764
rect 6323 -797 6911 -781
rect 7341 -781 7357 -764
rect 7913 -764 8115 -747
rect 8173 -747 9133 -709
rect 8173 -764 8375 -747
rect 7913 -781 7929 -764
rect 7341 -797 7929 -781
rect 8359 -781 8375 -764
rect 8931 -764 9133 -747
rect 9191 -747 10151 -709
rect 9191 -764 9393 -747
rect 8931 -781 8947 -764
rect 8359 -797 8947 -781
rect 9377 -781 9393 -764
rect 9949 -764 10151 -747
rect 9949 -781 9965 -764
rect 9377 -797 9965 -781
<< polycont >>
rect -9949 747 -9393 781
rect -8931 747 -8375 781
rect -7913 747 -7357 781
rect -6895 747 -6339 781
rect -5877 747 -5321 781
rect -4859 747 -4303 781
rect -3841 747 -3285 781
rect -2823 747 -2267 781
rect -1805 747 -1249 781
rect -787 747 -231 781
rect 231 747 787 781
rect 1249 747 1805 781
rect 2267 747 2823 781
rect 3285 747 3841 781
rect 4303 747 4859 781
rect 5321 747 5877 781
rect 6339 747 6895 781
rect 7357 747 7913 781
rect 8375 747 8931 781
rect 9393 747 9949 781
rect -9949 37 -9393 71
rect -8931 37 -8375 71
rect -7913 37 -7357 71
rect -6895 37 -6339 71
rect -5877 37 -5321 71
rect -4859 37 -4303 71
rect -3841 37 -3285 71
rect -2823 37 -2267 71
rect -1805 37 -1249 71
rect -787 37 -231 71
rect 231 37 787 71
rect 1249 37 1805 71
rect 2267 37 2823 71
rect 3285 37 3841 71
rect 4303 37 4859 71
rect 5321 37 5877 71
rect 6339 37 6895 71
rect 7357 37 7913 71
rect 8375 37 8931 71
rect 9393 37 9949 71
rect -9949 -71 -9393 -37
rect -8931 -71 -8375 -37
rect -7913 -71 -7357 -37
rect -6895 -71 -6339 -37
rect -5877 -71 -5321 -37
rect -4859 -71 -4303 -37
rect -3841 -71 -3285 -37
rect -2823 -71 -2267 -37
rect -1805 -71 -1249 -37
rect -787 -71 -231 -37
rect 231 -71 787 -37
rect 1249 -71 1805 -37
rect 2267 -71 2823 -37
rect 3285 -71 3841 -37
rect 4303 -71 4859 -37
rect 5321 -71 5877 -37
rect 6339 -71 6895 -37
rect 7357 -71 7913 -37
rect 8375 -71 8931 -37
rect 9393 -71 9949 -37
rect -9949 -781 -9393 -747
rect -8931 -781 -8375 -747
rect -7913 -781 -7357 -747
rect -6895 -781 -6339 -747
rect -5877 -781 -5321 -747
rect -4859 -781 -4303 -747
rect -3841 -781 -3285 -747
rect -2823 -781 -2267 -747
rect -1805 -781 -1249 -747
rect -787 -781 -231 -747
rect 231 -781 787 -747
rect 1249 -781 1805 -747
rect 2267 -781 2823 -747
rect 3285 -781 3841 -747
rect 4303 -781 4859 -747
rect 5321 -781 5877 -747
rect 6339 -781 6895 -747
rect 7357 -781 7913 -747
rect 8375 -781 8931 -747
rect 9393 -781 9949 -747
<< locali >>
rect -9965 747 -9949 781
rect -9393 747 -9377 781
rect -8947 747 -8931 781
rect -8375 747 -8359 781
rect -7929 747 -7913 781
rect -7357 747 -7341 781
rect -6911 747 -6895 781
rect -6339 747 -6323 781
rect -5893 747 -5877 781
rect -5321 747 -5305 781
rect -4875 747 -4859 781
rect -4303 747 -4287 781
rect -3857 747 -3841 781
rect -3285 747 -3269 781
rect -2839 747 -2823 781
rect -2267 747 -2251 781
rect -1821 747 -1805 781
rect -1249 747 -1233 781
rect -803 747 -787 781
rect -231 747 -215 781
rect 215 747 231 781
rect 787 747 803 781
rect 1233 747 1249 781
rect 1805 747 1821 781
rect 2251 747 2267 781
rect 2823 747 2839 781
rect 3269 747 3285 781
rect 3841 747 3857 781
rect 4287 747 4303 781
rect 4859 747 4875 781
rect 5305 747 5321 781
rect 5877 747 5893 781
rect 6323 747 6339 781
rect 6895 747 6911 781
rect 7341 747 7357 781
rect 7913 747 7929 781
rect 8359 747 8375 781
rect 8931 747 8947 781
rect 9377 747 9393 781
rect 9949 747 9965 781
rect -10197 697 -10163 713
rect -10197 105 -10163 121
rect -9179 697 -9145 713
rect -9179 105 -9145 121
rect -8161 697 -8127 713
rect -8161 105 -8127 121
rect -7143 697 -7109 713
rect -7143 105 -7109 121
rect -6125 697 -6091 713
rect -6125 105 -6091 121
rect -5107 697 -5073 713
rect -5107 105 -5073 121
rect -4089 697 -4055 713
rect -4089 105 -4055 121
rect -3071 697 -3037 713
rect -3071 105 -3037 121
rect -2053 697 -2019 713
rect -2053 105 -2019 121
rect -1035 697 -1001 713
rect -1035 105 -1001 121
rect -17 697 17 713
rect -17 105 17 121
rect 1001 697 1035 713
rect 1001 105 1035 121
rect 2019 697 2053 713
rect 2019 105 2053 121
rect 3037 697 3071 713
rect 3037 105 3071 121
rect 4055 697 4089 713
rect 4055 105 4089 121
rect 5073 697 5107 713
rect 5073 105 5107 121
rect 6091 697 6125 713
rect 6091 105 6125 121
rect 7109 697 7143 713
rect 7109 105 7143 121
rect 8127 697 8161 713
rect 8127 105 8161 121
rect 9145 697 9179 713
rect 9145 105 9179 121
rect 10163 697 10197 713
rect 10163 105 10197 121
rect -9965 37 -9949 71
rect -9393 37 -9377 71
rect -8947 37 -8931 71
rect -8375 37 -8359 71
rect -7929 37 -7913 71
rect -7357 37 -7341 71
rect -6911 37 -6895 71
rect -6339 37 -6323 71
rect -5893 37 -5877 71
rect -5321 37 -5305 71
rect -4875 37 -4859 71
rect -4303 37 -4287 71
rect -3857 37 -3841 71
rect -3285 37 -3269 71
rect -2839 37 -2823 71
rect -2267 37 -2251 71
rect -1821 37 -1805 71
rect -1249 37 -1233 71
rect -803 37 -787 71
rect -231 37 -215 71
rect 215 37 231 71
rect 787 37 803 71
rect 1233 37 1249 71
rect 1805 37 1821 71
rect 2251 37 2267 71
rect 2823 37 2839 71
rect 3269 37 3285 71
rect 3841 37 3857 71
rect 4287 37 4303 71
rect 4859 37 4875 71
rect 5305 37 5321 71
rect 5877 37 5893 71
rect 6323 37 6339 71
rect 6895 37 6911 71
rect 7341 37 7357 71
rect 7913 37 7929 71
rect 8359 37 8375 71
rect 8931 37 8947 71
rect 9377 37 9393 71
rect 9949 37 9965 71
rect -9965 -71 -9949 -37
rect -9393 -71 -9377 -37
rect -8947 -71 -8931 -37
rect -8375 -71 -8359 -37
rect -7929 -71 -7913 -37
rect -7357 -71 -7341 -37
rect -6911 -71 -6895 -37
rect -6339 -71 -6323 -37
rect -5893 -71 -5877 -37
rect -5321 -71 -5305 -37
rect -4875 -71 -4859 -37
rect -4303 -71 -4287 -37
rect -3857 -71 -3841 -37
rect -3285 -71 -3269 -37
rect -2839 -71 -2823 -37
rect -2267 -71 -2251 -37
rect -1821 -71 -1805 -37
rect -1249 -71 -1233 -37
rect -803 -71 -787 -37
rect -231 -71 -215 -37
rect 215 -71 231 -37
rect 787 -71 803 -37
rect 1233 -71 1249 -37
rect 1805 -71 1821 -37
rect 2251 -71 2267 -37
rect 2823 -71 2839 -37
rect 3269 -71 3285 -37
rect 3841 -71 3857 -37
rect 4287 -71 4303 -37
rect 4859 -71 4875 -37
rect 5305 -71 5321 -37
rect 5877 -71 5893 -37
rect 6323 -71 6339 -37
rect 6895 -71 6911 -37
rect 7341 -71 7357 -37
rect 7913 -71 7929 -37
rect 8359 -71 8375 -37
rect 8931 -71 8947 -37
rect 9377 -71 9393 -37
rect 9949 -71 9965 -37
rect -10197 -121 -10163 -105
rect -10197 -713 -10163 -697
rect -9179 -121 -9145 -105
rect -9179 -713 -9145 -697
rect -8161 -121 -8127 -105
rect -8161 -713 -8127 -697
rect -7143 -121 -7109 -105
rect -7143 -713 -7109 -697
rect -6125 -121 -6091 -105
rect -6125 -713 -6091 -697
rect -5107 -121 -5073 -105
rect -5107 -713 -5073 -697
rect -4089 -121 -4055 -105
rect -4089 -713 -4055 -697
rect -3071 -121 -3037 -105
rect -3071 -713 -3037 -697
rect -2053 -121 -2019 -105
rect -2053 -713 -2019 -697
rect -1035 -121 -1001 -105
rect -1035 -713 -1001 -697
rect -17 -121 17 -105
rect -17 -713 17 -697
rect 1001 -121 1035 -105
rect 1001 -713 1035 -697
rect 2019 -121 2053 -105
rect 2019 -713 2053 -697
rect 3037 -121 3071 -105
rect 3037 -713 3071 -697
rect 4055 -121 4089 -105
rect 4055 -713 4089 -697
rect 5073 -121 5107 -105
rect 5073 -713 5107 -697
rect 6091 -121 6125 -105
rect 6091 -713 6125 -697
rect 7109 -121 7143 -105
rect 7109 -713 7143 -697
rect 8127 -121 8161 -105
rect 8127 -713 8161 -697
rect 9145 -121 9179 -105
rect 9145 -713 9179 -697
rect 10163 -121 10197 -105
rect 10163 -713 10197 -697
rect -9965 -781 -9949 -747
rect -9393 -781 -9377 -747
rect -8947 -781 -8931 -747
rect -8375 -781 -8359 -747
rect -7929 -781 -7913 -747
rect -7357 -781 -7341 -747
rect -6911 -781 -6895 -747
rect -6339 -781 -6323 -747
rect -5893 -781 -5877 -747
rect -5321 -781 -5305 -747
rect -4875 -781 -4859 -747
rect -4303 -781 -4287 -747
rect -3857 -781 -3841 -747
rect -3285 -781 -3269 -747
rect -2839 -781 -2823 -747
rect -2267 -781 -2251 -747
rect -1821 -781 -1805 -747
rect -1249 -781 -1233 -747
rect -803 -781 -787 -747
rect -231 -781 -215 -747
rect 215 -781 231 -747
rect 787 -781 803 -747
rect 1233 -781 1249 -747
rect 1805 -781 1821 -747
rect 2251 -781 2267 -747
rect 2823 -781 2839 -747
rect 3269 -781 3285 -747
rect 3841 -781 3857 -747
rect 4287 -781 4303 -747
rect 4859 -781 4875 -747
rect 5305 -781 5321 -747
rect 5877 -781 5893 -747
rect 6323 -781 6339 -747
rect 6895 -781 6911 -747
rect 7341 -781 7357 -747
rect 7913 -781 7929 -747
rect 8359 -781 8375 -747
rect 8931 -781 8947 -747
rect 9377 -781 9393 -747
rect 9949 -781 9965 -747
<< viali >>
rect -9903 747 -9439 781
rect -8885 747 -8421 781
rect -7867 747 -7403 781
rect -6849 747 -6385 781
rect -5831 747 -5367 781
rect -4813 747 -4349 781
rect -3795 747 -3331 781
rect -2777 747 -2313 781
rect -1759 747 -1295 781
rect -741 747 -277 781
rect 277 747 741 781
rect 1295 747 1759 781
rect 2313 747 2777 781
rect 3331 747 3795 781
rect 4349 747 4813 781
rect 5367 747 5831 781
rect 6385 747 6849 781
rect 7403 747 7867 781
rect 8421 747 8885 781
rect 9439 747 9903 781
rect -10197 121 -10163 697
rect -9179 121 -9145 697
rect -8161 121 -8127 697
rect -7143 121 -7109 697
rect -6125 121 -6091 697
rect -5107 121 -5073 697
rect -4089 121 -4055 697
rect -3071 121 -3037 697
rect -2053 121 -2019 697
rect -1035 121 -1001 697
rect -17 121 17 697
rect 1001 121 1035 697
rect 2019 121 2053 697
rect 3037 121 3071 697
rect 4055 121 4089 697
rect 5073 121 5107 697
rect 6091 121 6125 697
rect 7109 121 7143 697
rect 8127 121 8161 697
rect 9145 121 9179 697
rect 10163 121 10197 697
rect -9903 37 -9439 71
rect -8885 37 -8421 71
rect -7867 37 -7403 71
rect -6849 37 -6385 71
rect -5831 37 -5367 71
rect -4813 37 -4349 71
rect -3795 37 -3331 71
rect -2777 37 -2313 71
rect -1759 37 -1295 71
rect -741 37 -277 71
rect 277 37 741 71
rect 1295 37 1759 71
rect 2313 37 2777 71
rect 3331 37 3795 71
rect 4349 37 4813 71
rect 5367 37 5831 71
rect 6385 37 6849 71
rect 7403 37 7867 71
rect 8421 37 8885 71
rect 9439 37 9903 71
rect -9903 -71 -9439 -37
rect -8885 -71 -8421 -37
rect -7867 -71 -7403 -37
rect -6849 -71 -6385 -37
rect -5831 -71 -5367 -37
rect -4813 -71 -4349 -37
rect -3795 -71 -3331 -37
rect -2777 -71 -2313 -37
rect -1759 -71 -1295 -37
rect -741 -71 -277 -37
rect 277 -71 741 -37
rect 1295 -71 1759 -37
rect 2313 -71 2777 -37
rect 3331 -71 3795 -37
rect 4349 -71 4813 -37
rect 5367 -71 5831 -37
rect 6385 -71 6849 -37
rect 7403 -71 7867 -37
rect 8421 -71 8885 -37
rect 9439 -71 9903 -37
rect -10197 -697 -10163 -121
rect -9179 -697 -9145 -121
rect -8161 -697 -8127 -121
rect -7143 -697 -7109 -121
rect -6125 -697 -6091 -121
rect -5107 -697 -5073 -121
rect -4089 -697 -4055 -121
rect -3071 -697 -3037 -121
rect -2053 -697 -2019 -121
rect -1035 -697 -1001 -121
rect -17 -697 17 -121
rect 1001 -697 1035 -121
rect 2019 -697 2053 -121
rect 3037 -697 3071 -121
rect 4055 -697 4089 -121
rect 5073 -697 5107 -121
rect 6091 -697 6125 -121
rect 7109 -697 7143 -121
rect 8127 -697 8161 -121
rect 9145 -697 9179 -121
rect 10163 -697 10197 -121
rect -9903 -781 -9439 -747
rect -8885 -781 -8421 -747
rect -7867 -781 -7403 -747
rect -6849 -781 -6385 -747
rect -5831 -781 -5367 -747
rect -4813 -781 -4349 -747
rect -3795 -781 -3331 -747
rect -2777 -781 -2313 -747
rect -1759 -781 -1295 -747
rect -741 -781 -277 -747
rect 277 -781 741 -747
rect 1295 -781 1759 -747
rect 2313 -781 2777 -747
rect 3331 -781 3795 -747
rect 4349 -781 4813 -747
rect 5367 -781 5831 -747
rect 6385 -781 6849 -747
rect 7403 -781 7867 -747
rect 8421 -781 8885 -747
rect 9439 -781 9903 -747
<< metal1 >>
rect -9915 781 -9427 787
rect -9915 747 -9903 781
rect -9439 747 -9427 781
rect -9915 741 -9427 747
rect -8897 781 -8409 787
rect -8897 747 -8885 781
rect -8421 747 -8409 781
rect -8897 741 -8409 747
rect -7879 781 -7391 787
rect -7879 747 -7867 781
rect -7403 747 -7391 781
rect -7879 741 -7391 747
rect -6861 781 -6373 787
rect -6861 747 -6849 781
rect -6385 747 -6373 781
rect -6861 741 -6373 747
rect -5843 781 -5355 787
rect -5843 747 -5831 781
rect -5367 747 -5355 781
rect -5843 741 -5355 747
rect -4825 781 -4337 787
rect -4825 747 -4813 781
rect -4349 747 -4337 781
rect -4825 741 -4337 747
rect -3807 781 -3319 787
rect -3807 747 -3795 781
rect -3331 747 -3319 781
rect -3807 741 -3319 747
rect -2789 781 -2301 787
rect -2789 747 -2777 781
rect -2313 747 -2301 781
rect -2789 741 -2301 747
rect -1771 781 -1283 787
rect -1771 747 -1759 781
rect -1295 747 -1283 781
rect -1771 741 -1283 747
rect -753 781 -265 787
rect -753 747 -741 781
rect -277 747 -265 781
rect -753 741 -265 747
rect 265 781 753 787
rect 265 747 277 781
rect 741 747 753 781
rect 265 741 753 747
rect 1283 781 1771 787
rect 1283 747 1295 781
rect 1759 747 1771 781
rect 1283 741 1771 747
rect 2301 781 2789 787
rect 2301 747 2313 781
rect 2777 747 2789 781
rect 2301 741 2789 747
rect 3319 781 3807 787
rect 3319 747 3331 781
rect 3795 747 3807 781
rect 3319 741 3807 747
rect 4337 781 4825 787
rect 4337 747 4349 781
rect 4813 747 4825 781
rect 4337 741 4825 747
rect 5355 781 5843 787
rect 5355 747 5367 781
rect 5831 747 5843 781
rect 5355 741 5843 747
rect 6373 781 6861 787
rect 6373 747 6385 781
rect 6849 747 6861 781
rect 6373 741 6861 747
rect 7391 781 7879 787
rect 7391 747 7403 781
rect 7867 747 7879 781
rect 7391 741 7879 747
rect 8409 781 8897 787
rect 8409 747 8421 781
rect 8885 747 8897 781
rect 8409 741 8897 747
rect 9427 781 9915 787
rect 9427 747 9439 781
rect 9903 747 9915 781
rect 9427 741 9915 747
rect -10203 697 -10157 709
rect -10203 121 -10197 697
rect -10163 121 -10157 697
rect -10203 109 -10157 121
rect -9185 697 -9139 709
rect -9185 121 -9179 697
rect -9145 121 -9139 697
rect -9185 109 -9139 121
rect -8167 697 -8121 709
rect -8167 121 -8161 697
rect -8127 121 -8121 697
rect -8167 109 -8121 121
rect -7149 697 -7103 709
rect -7149 121 -7143 697
rect -7109 121 -7103 697
rect -7149 109 -7103 121
rect -6131 697 -6085 709
rect -6131 121 -6125 697
rect -6091 121 -6085 697
rect -6131 109 -6085 121
rect -5113 697 -5067 709
rect -5113 121 -5107 697
rect -5073 121 -5067 697
rect -5113 109 -5067 121
rect -4095 697 -4049 709
rect -4095 121 -4089 697
rect -4055 121 -4049 697
rect -4095 109 -4049 121
rect -3077 697 -3031 709
rect -3077 121 -3071 697
rect -3037 121 -3031 697
rect -3077 109 -3031 121
rect -2059 697 -2013 709
rect -2059 121 -2053 697
rect -2019 121 -2013 697
rect -2059 109 -2013 121
rect -1041 697 -995 709
rect -1041 121 -1035 697
rect -1001 121 -995 697
rect -1041 109 -995 121
rect -23 697 23 709
rect -23 121 -17 697
rect 17 121 23 697
rect -23 109 23 121
rect 995 697 1041 709
rect 995 121 1001 697
rect 1035 121 1041 697
rect 995 109 1041 121
rect 2013 697 2059 709
rect 2013 121 2019 697
rect 2053 121 2059 697
rect 2013 109 2059 121
rect 3031 697 3077 709
rect 3031 121 3037 697
rect 3071 121 3077 697
rect 3031 109 3077 121
rect 4049 697 4095 709
rect 4049 121 4055 697
rect 4089 121 4095 697
rect 4049 109 4095 121
rect 5067 697 5113 709
rect 5067 121 5073 697
rect 5107 121 5113 697
rect 5067 109 5113 121
rect 6085 697 6131 709
rect 6085 121 6091 697
rect 6125 121 6131 697
rect 6085 109 6131 121
rect 7103 697 7149 709
rect 7103 121 7109 697
rect 7143 121 7149 697
rect 7103 109 7149 121
rect 8121 697 8167 709
rect 8121 121 8127 697
rect 8161 121 8167 697
rect 8121 109 8167 121
rect 9139 697 9185 709
rect 9139 121 9145 697
rect 9179 121 9185 697
rect 9139 109 9185 121
rect 10157 697 10203 709
rect 10157 121 10163 697
rect 10197 121 10203 697
rect 10157 109 10203 121
rect -9915 71 -9427 77
rect -9915 37 -9903 71
rect -9439 37 -9427 71
rect -9915 31 -9427 37
rect -8897 71 -8409 77
rect -8897 37 -8885 71
rect -8421 37 -8409 71
rect -8897 31 -8409 37
rect -7879 71 -7391 77
rect -7879 37 -7867 71
rect -7403 37 -7391 71
rect -7879 31 -7391 37
rect -6861 71 -6373 77
rect -6861 37 -6849 71
rect -6385 37 -6373 71
rect -6861 31 -6373 37
rect -5843 71 -5355 77
rect -5843 37 -5831 71
rect -5367 37 -5355 71
rect -5843 31 -5355 37
rect -4825 71 -4337 77
rect -4825 37 -4813 71
rect -4349 37 -4337 71
rect -4825 31 -4337 37
rect -3807 71 -3319 77
rect -3807 37 -3795 71
rect -3331 37 -3319 71
rect -3807 31 -3319 37
rect -2789 71 -2301 77
rect -2789 37 -2777 71
rect -2313 37 -2301 71
rect -2789 31 -2301 37
rect -1771 71 -1283 77
rect -1771 37 -1759 71
rect -1295 37 -1283 71
rect -1771 31 -1283 37
rect -753 71 -265 77
rect -753 37 -741 71
rect -277 37 -265 71
rect -753 31 -265 37
rect 265 71 753 77
rect 265 37 277 71
rect 741 37 753 71
rect 265 31 753 37
rect 1283 71 1771 77
rect 1283 37 1295 71
rect 1759 37 1771 71
rect 1283 31 1771 37
rect 2301 71 2789 77
rect 2301 37 2313 71
rect 2777 37 2789 71
rect 2301 31 2789 37
rect 3319 71 3807 77
rect 3319 37 3331 71
rect 3795 37 3807 71
rect 3319 31 3807 37
rect 4337 71 4825 77
rect 4337 37 4349 71
rect 4813 37 4825 71
rect 4337 31 4825 37
rect 5355 71 5843 77
rect 5355 37 5367 71
rect 5831 37 5843 71
rect 5355 31 5843 37
rect 6373 71 6861 77
rect 6373 37 6385 71
rect 6849 37 6861 71
rect 6373 31 6861 37
rect 7391 71 7879 77
rect 7391 37 7403 71
rect 7867 37 7879 71
rect 7391 31 7879 37
rect 8409 71 8897 77
rect 8409 37 8421 71
rect 8885 37 8897 71
rect 8409 31 8897 37
rect 9427 71 9915 77
rect 9427 37 9439 71
rect 9903 37 9915 71
rect 9427 31 9915 37
rect -9915 -37 -9427 -31
rect -9915 -71 -9903 -37
rect -9439 -71 -9427 -37
rect -9915 -77 -9427 -71
rect -8897 -37 -8409 -31
rect -8897 -71 -8885 -37
rect -8421 -71 -8409 -37
rect -8897 -77 -8409 -71
rect -7879 -37 -7391 -31
rect -7879 -71 -7867 -37
rect -7403 -71 -7391 -37
rect -7879 -77 -7391 -71
rect -6861 -37 -6373 -31
rect -6861 -71 -6849 -37
rect -6385 -71 -6373 -37
rect -6861 -77 -6373 -71
rect -5843 -37 -5355 -31
rect -5843 -71 -5831 -37
rect -5367 -71 -5355 -37
rect -5843 -77 -5355 -71
rect -4825 -37 -4337 -31
rect -4825 -71 -4813 -37
rect -4349 -71 -4337 -37
rect -4825 -77 -4337 -71
rect -3807 -37 -3319 -31
rect -3807 -71 -3795 -37
rect -3331 -71 -3319 -37
rect -3807 -77 -3319 -71
rect -2789 -37 -2301 -31
rect -2789 -71 -2777 -37
rect -2313 -71 -2301 -37
rect -2789 -77 -2301 -71
rect -1771 -37 -1283 -31
rect -1771 -71 -1759 -37
rect -1295 -71 -1283 -37
rect -1771 -77 -1283 -71
rect -753 -37 -265 -31
rect -753 -71 -741 -37
rect -277 -71 -265 -37
rect -753 -77 -265 -71
rect 265 -37 753 -31
rect 265 -71 277 -37
rect 741 -71 753 -37
rect 265 -77 753 -71
rect 1283 -37 1771 -31
rect 1283 -71 1295 -37
rect 1759 -71 1771 -37
rect 1283 -77 1771 -71
rect 2301 -37 2789 -31
rect 2301 -71 2313 -37
rect 2777 -71 2789 -37
rect 2301 -77 2789 -71
rect 3319 -37 3807 -31
rect 3319 -71 3331 -37
rect 3795 -71 3807 -37
rect 3319 -77 3807 -71
rect 4337 -37 4825 -31
rect 4337 -71 4349 -37
rect 4813 -71 4825 -37
rect 4337 -77 4825 -71
rect 5355 -37 5843 -31
rect 5355 -71 5367 -37
rect 5831 -71 5843 -37
rect 5355 -77 5843 -71
rect 6373 -37 6861 -31
rect 6373 -71 6385 -37
rect 6849 -71 6861 -37
rect 6373 -77 6861 -71
rect 7391 -37 7879 -31
rect 7391 -71 7403 -37
rect 7867 -71 7879 -37
rect 7391 -77 7879 -71
rect 8409 -37 8897 -31
rect 8409 -71 8421 -37
rect 8885 -71 8897 -37
rect 8409 -77 8897 -71
rect 9427 -37 9915 -31
rect 9427 -71 9439 -37
rect 9903 -71 9915 -37
rect 9427 -77 9915 -71
rect -10203 -121 -10157 -109
rect -10203 -697 -10197 -121
rect -10163 -697 -10157 -121
rect -10203 -709 -10157 -697
rect -9185 -121 -9139 -109
rect -9185 -697 -9179 -121
rect -9145 -697 -9139 -121
rect -9185 -709 -9139 -697
rect -8167 -121 -8121 -109
rect -8167 -697 -8161 -121
rect -8127 -697 -8121 -121
rect -8167 -709 -8121 -697
rect -7149 -121 -7103 -109
rect -7149 -697 -7143 -121
rect -7109 -697 -7103 -121
rect -7149 -709 -7103 -697
rect -6131 -121 -6085 -109
rect -6131 -697 -6125 -121
rect -6091 -697 -6085 -121
rect -6131 -709 -6085 -697
rect -5113 -121 -5067 -109
rect -5113 -697 -5107 -121
rect -5073 -697 -5067 -121
rect -5113 -709 -5067 -697
rect -4095 -121 -4049 -109
rect -4095 -697 -4089 -121
rect -4055 -697 -4049 -121
rect -4095 -709 -4049 -697
rect -3077 -121 -3031 -109
rect -3077 -697 -3071 -121
rect -3037 -697 -3031 -121
rect -3077 -709 -3031 -697
rect -2059 -121 -2013 -109
rect -2059 -697 -2053 -121
rect -2019 -697 -2013 -121
rect -2059 -709 -2013 -697
rect -1041 -121 -995 -109
rect -1041 -697 -1035 -121
rect -1001 -697 -995 -121
rect -1041 -709 -995 -697
rect -23 -121 23 -109
rect -23 -697 -17 -121
rect 17 -697 23 -121
rect -23 -709 23 -697
rect 995 -121 1041 -109
rect 995 -697 1001 -121
rect 1035 -697 1041 -121
rect 995 -709 1041 -697
rect 2013 -121 2059 -109
rect 2013 -697 2019 -121
rect 2053 -697 2059 -121
rect 2013 -709 2059 -697
rect 3031 -121 3077 -109
rect 3031 -697 3037 -121
rect 3071 -697 3077 -121
rect 3031 -709 3077 -697
rect 4049 -121 4095 -109
rect 4049 -697 4055 -121
rect 4089 -697 4095 -121
rect 4049 -709 4095 -697
rect 5067 -121 5113 -109
rect 5067 -697 5073 -121
rect 5107 -697 5113 -121
rect 5067 -709 5113 -697
rect 6085 -121 6131 -109
rect 6085 -697 6091 -121
rect 6125 -697 6131 -121
rect 6085 -709 6131 -697
rect 7103 -121 7149 -109
rect 7103 -697 7109 -121
rect 7143 -697 7149 -121
rect 7103 -709 7149 -697
rect 8121 -121 8167 -109
rect 8121 -697 8127 -121
rect 8161 -697 8167 -121
rect 8121 -709 8167 -697
rect 9139 -121 9185 -109
rect 9139 -697 9145 -121
rect 9179 -697 9185 -121
rect 9139 -709 9185 -697
rect 10157 -121 10203 -109
rect 10157 -697 10163 -121
rect 10197 -697 10203 -121
rect 10157 -709 10203 -697
rect -9915 -747 -9427 -741
rect -9915 -781 -9903 -747
rect -9439 -781 -9427 -747
rect -9915 -787 -9427 -781
rect -8897 -747 -8409 -741
rect -8897 -781 -8885 -747
rect -8421 -781 -8409 -747
rect -8897 -787 -8409 -781
rect -7879 -747 -7391 -741
rect -7879 -781 -7867 -747
rect -7403 -781 -7391 -747
rect -7879 -787 -7391 -781
rect -6861 -747 -6373 -741
rect -6861 -781 -6849 -747
rect -6385 -781 -6373 -747
rect -6861 -787 -6373 -781
rect -5843 -747 -5355 -741
rect -5843 -781 -5831 -747
rect -5367 -781 -5355 -747
rect -5843 -787 -5355 -781
rect -4825 -747 -4337 -741
rect -4825 -781 -4813 -747
rect -4349 -781 -4337 -747
rect -4825 -787 -4337 -781
rect -3807 -747 -3319 -741
rect -3807 -781 -3795 -747
rect -3331 -781 -3319 -747
rect -3807 -787 -3319 -781
rect -2789 -747 -2301 -741
rect -2789 -781 -2777 -747
rect -2313 -781 -2301 -747
rect -2789 -787 -2301 -781
rect -1771 -747 -1283 -741
rect -1771 -781 -1759 -747
rect -1295 -781 -1283 -747
rect -1771 -787 -1283 -781
rect -753 -747 -265 -741
rect -753 -781 -741 -747
rect -277 -781 -265 -747
rect -753 -787 -265 -781
rect 265 -747 753 -741
rect 265 -781 277 -747
rect 741 -781 753 -747
rect 265 -787 753 -781
rect 1283 -747 1771 -741
rect 1283 -781 1295 -747
rect 1759 -781 1771 -747
rect 1283 -787 1771 -781
rect 2301 -747 2789 -741
rect 2301 -781 2313 -747
rect 2777 -781 2789 -747
rect 2301 -787 2789 -781
rect 3319 -747 3807 -741
rect 3319 -781 3331 -747
rect 3795 -781 3807 -747
rect 3319 -787 3807 -781
rect 4337 -747 4825 -741
rect 4337 -781 4349 -747
rect 4813 -781 4825 -747
rect 4337 -787 4825 -781
rect 5355 -747 5843 -741
rect 5355 -781 5367 -747
rect 5831 -781 5843 -747
rect 5355 -787 5843 -781
rect 6373 -747 6861 -741
rect 6373 -781 6385 -747
rect 6849 -781 6861 -747
rect 6373 -787 6861 -781
rect 7391 -747 7879 -741
rect 7391 -781 7403 -747
rect 7867 -781 7879 -747
rect 7391 -787 7879 -781
rect 8409 -747 8897 -741
rect 8409 -781 8421 -747
rect 8885 -781 8897 -747
rect 8409 -787 8897 -781
rect 9427 -747 9915 -741
rect 9427 -781 9439 -747
rect 9903 -781 9915 -747
rect 9427 -787 9915 -781
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string parameters w 3 l 4.8 m 2 nf 20 diffcov 100 polycov 60 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
