magic
tech sky130A
magscale 1 2
timestamp 1626486988
<< checkpaint >>
rect -5615 -1460 5615 1460
<< nwell >>
rect -4355 -200 4355 200
<< pmos >>
rect -4261 -100 -3461 100
rect -3403 -100 -2603 100
rect -2545 -100 -1745 100
rect -1687 -100 -887 100
rect -829 -100 -29 100
rect 29 -100 829 100
rect 887 -100 1687 100
rect 1745 -100 2545 100
rect 2603 -100 3403 100
rect 3461 -100 4261 100
<< pdiff >>
rect -4319 85 -4261 100
rect -4319 51 -4307 85
rect -4273 51 -4261 85
rect -4319 17 -4261 51
rect -4319 -17 -4307 17
rect -4273 -17 -4261 17
rect -4319 -51 -4261 -17
rect -4319 -85 -4307 -51
rect -4273 -85 -4261 -51
rect -4319 -100 -4261 -85
rect -3461 85 -3403 100
rect -3461 51 -3449 85
rect -3415 51 -3403 85
rect -3461 17 -3403 51
rect -3461 -17 -3449 17
rect -3415 -17 -3403 17
rect -3461 -51 -3403 -17
rect -3461 -85 -3449 -51
rect -3415 -85 -3403 -51
rect -3461 -100 -3403 -85
rect -2603 85 -2545 100
rect -2603 51 -2591 85
rect -2557 51 -2545 85
rect -2603 17 -2545 51
rect -2603 -17 -2591 17
rect -2557 -17 -2545 17
rect -2603 -51 -2545 -17
rect -2603 -85 -2591 -51
rect -2557 -85 -2545 -51
rect -2603 -100 -2545 -85
rect -1745 85 -1687 100
rect -1745 51 -1733 85
rect -1699 51 -1687 85
rect -1745 17 -1687 51
rect -1745 -17 -1733 17
rect -1699 -17 -1687 17
rect -1745 -51 -1687 -17
rect -1745 -85 -1733 -51
rect -1699 -85 -1687 -51
rect -1745 -100 -1687 -85
rect -887 85 -829 100
rect -887 51 -875 85
rect -841 51 -829 85
rect -887 17 -829 51
rect -887 -17 -875 17
rect -841 -17 -829 17
rect -887 -51 -829 -17
rect -887 -85 -875 -51
rect -841 -85 -829 -51
rect -887 -100 -829 -85
rect -29 85 29 100
rect -29 51 -17 85
rect 17 51 29 85
rect -29 17 29 51
rect -29 -17 -17 17
rect 17 -17 29 17
rect -29 -51 29 -17
rect -29 -85 -17 -51
rect 17 -85 29 -51
rect -29 -100 29 -85
rect 829 85 887 100
rect 829 51 841 85
rect 875 51 887 85
rect 829 17 887 51
rect 829 -17 841 17
rect 875 -17 887 17
rect 829 -51 887 -17
rect 829 -85 841 -51
rect 875 -85 887 -51
rect 829 -100 887 -85
rect 1687 85 1745 100
rect 1687 51 1699 85
rect 1733 51 1745 85
rect 1687 17 1745 51
rect 1687 -17 1699 17
rect 1733 -17 1745 17
rect 1687 -51 1745 -17
rect 1687 -85 1699 -51
rect 1733 -85 1745 -51
rect 1687 -100 1745 -85
rect 2545 85 2603 100
rect 2545 51 2557 85
rect 2591 51 2603 85
rect 2545 17 2603 51
rect 2545 -17 2557 17
rect 2591 -17 2603 17
rect 2545 -51 2603 -17
rect 2545 -85 2557 -51
rect 2591 -85 2603 -51
rect 2545 -100 2603 -85
rect 3403 85 3461 100
rect 3403 51 3415 85
rect 3449 51 3461 85
rect 3403 17 3461 51
rect 3403 -17 3415 17
rect 3449 -17 3461 17
rect 3403 -51 3461 -17
rect 3403 -85 3415 -51
rect 3449 -85 3461 -51
rect 3403 -100 3461 -85
rect 4261 85 4319 100
rect 4261 51 4273 85
rect 4307 51 4319 85
rect 4261 17 4319 51
rect 4261 -17 4273 17
rect 4307 -17 4319 17
rect 4261 -51 4319 -17
rect 4261 -85 4273 -51
rect 4307 -85 4319 -51
rect 4261 -100 4319 -85
<< pdiffc >>
rect -4307 51 -4273 85
rect -4307 -17 -4273 17
rect -4307 -85 -4273 -51
rect -3449 51 -3415 85
rect -3449 -17 -3415 17
rect -3449 -85 -3415 -51
rect -2591 51 -2557 85
rect -2591 -17 -2557 17
rect -2591 -85 -2557 -51
rect -1733 51 -1699 85
rect -1733 -17 -1699 17
rect -1733 -85 -1699 -51
rect -875 51 -841 85
rect -875 -17 -841 17
rect -875 -85 -841 -51
rect -17 51 17 85
rect -17 -17 17 17
rect -17 -85 17 -51
rect 841 51 875 85
rect 841 -17 875 17
rect 841 -85 875 -51
rect 1699 51 1733 85
rect 1699 -17 1733 17
rect 1699 -85 1733 -51
rect 2557 51 2591 85
rect 2557 -17 2591 17
rect 2557 -85 2591 -51
rect 3415 51 3449 85
rect 3415 -17 3449 17
rect 3415 -85 3449 -51
rect 4273 51 4307 85
rect 4273 -17 4307 17
rect 4273 -85 4307 -51
<< poly >>
rect -4069 181 -3653 197
rect -4069 164 -4048 181
rect -4261 147 -4048 164
rect -4014 147 -3980 181
rect -3946 147 -3912 181
rect -3878 147 -3844 181
rect -3810 147 -3776 181
rect -3742 147 -3708 181
rect -3674 164 -3653 181
rect -3211 181 -2795 197
rect -3211 164 -3190 181
rect -3674 147 -3461 164
rect -4261 100 -3461 147
rect -3403 147 -3190 164
rect -3156 147 -3122 181
rect -3088 147 -3054 181
rect -3020 147 -2986 181
rect -2952 147 -2918 181
rect -2884 147 -2850 181
rect -2816 164 -2795 181
rect -2353 181 -1937 197
rect -2353 164 -2332 181
rect -2816 147 -2603 164
rect -3403 100 -2603 147
rect -2545 147 -2332 164
rect -2298 147 -2264 181
rect -2230 147 -2196 181
rect -2162 147 -2128 181
rect -2094 147 -2060 181
rect -2026 147 -1992 181
rect -1958 164 -1937 181
rect -1495 181 -1079 197
rect -1495 164 -1474 181
rect -1958 147 -1745 164
rect -2545 100 -1745 147
rect -1687 147 -1474 164
rect -1440 147 -1406 181
rect -1372 147 -1338 181
rect -1304 147 -1270 181
rect -1236 147 -1202 181
rect -1168 147 -1134 181
rect -1100 164 -1079 181
rect -637 181 -221 197
rect -637 164 -616 181
rect -1100 147 -887 164
rect -1687 100 -887 147
rect -829 147 -616 164
rect -582 147 -548 181
rect -514 147 -480 181
rect -446 147 -412 181
rect -378 147 -344 181
rect -310 147 -276 181
rect -242 164 -221 181
rect 221 181 637 197
rect 221 164 242 181
rect -242 147 -29 164
rect -829 100 -29 147
rect 29 147 242 164
rect 276 147 310 181
rect 344 147 378 181
rect 412 147 446 181
rect 480 147 514 181
rect 548 147 582 181
rect 616 164 637 181
rect 1079 181 1495 197
rect 1079 164 1100 181
rect 616 147 829 164
rect 29 100 829 147
rect 887 147 1100 164
rect 1134 147 1168 181
rect 1202 147 1236 181
rect 1270 147 1304 181
rect 1338 147 1372 181
rect 1406 147 1440 181
rect 1474 164 1495 181
rect 1937 181 2353 197
rect 1937 164 1958 181
rect 1474 147 1687 164
rect 887 100 1687 147
rect 1745 147 1958 164
rect 1992 147 2026 181
rect 2060 147 2094 181
rect 2128 147 2162 181
rect 2196 147 2230 181
rect 2264 147 2298 181
rect 2332 164 2353 181
rect 2795 181 3211 197
rect 2795 164 2816 181
rect 2332 147 2545 164
rect 1745 100 2545 147
rect 2603 147 2816 164
rect 2850 147 2884 181
rect 2918 147 2952 181
rect 2986 147 3020 181
rect 3054 147 3088 181
rect 3122 147 3156 181
rect 3190 164 3211 181
rect 3653 181 4069 197
rect 3653 164 3674 181
rect 3190 147 3403 164
rect 2603 100 3403 147
rect 3461 147 3674 164
rect 3708 147 3742 181
rect 3776 147 3810 181
rect 3844 147 3878 181
rect 3912 147 3946 181
rect 3980 147 4014 181
rect 4048 164 4069 181
rect 4048 147 4261 164
rect 3461 100 4261 147
rect -4261 -147 -3461 -100
rect -4261 -164 -4048 -147
rect -4069 -181 -4048 -164
rect -4014 -181 -3980 -147
rect -3946 -181 -3912 -147
rect -3878 -181 -3844 -147
rect -3810 -181 -3776 -147
rect -3742 -181 -3708 -147
rect -3674 -164 -3461 -147
rect -3403 -147 -2603 -100
rect -3403 -164 -3190 -147
rect -3674 -181 -3653 -164
rect -4069 -197 -3653 -181
rect -3211 -181 -3190 -164
rect -3156 -181 -3122 -147
rect -3088 -181 -3054 -147
rect -3020 -181 -2986 -147
rect -2952 -181 -2918 -147
rect -2884 -181 -2850 -147
rect -2816 -164 -2603 -147
rect -2545 -147 -1745 -100
rect -2545 -164 -2332 -147
rect -2816 -181 -2795 -164
rect -3211 -197 -2795 -181
rect -2353 -181 -2332 -164
rect -2298 -181 -2264 -147
rect -2230 -181 -2196 -147
rect -2162 -181 -2128 -147
rect -2094 -181 -2060 -147
rect -2026 -181 -1992 -147
rect -1958 -164 -1745 -147
rect -1687 -147 -887 -100
rect -1687 -164 -1474 -147
rect -1958 -181 -1937 -164
rect -2353 -197 -1937 -181
rect -1495 -181 -1474 -164
rect -1440 -181 -1406 -147
rect -1372 -181 -1338 -147
rect -1304 -181 -1270 -147
rect -1236 -181 -1202 -147
rect -1168 -181 -1134 -147
rect -1100 -164 -887 -147
rect -829 -147 -29 -100
rect -829 -164 -616 -147
rect -1100 -181 -1079 -164
rect -1495 -197 -1079 -181
rect -637 -181 -616 -164
rect -582 -181 -548 -147
rect -514 -181 -480 -147
rect -446 -181 -412 -147
rect -378 -181 -344 -147
rect -310 -181 -276 -147
rect -242 -164 -29 -147
rect 29 -147 829 -100
rect 29 -164 242 -147
rect -242 -181 -221 -164
rect -637 -197 -221 -181
rect 221 -181 242 -164
rect 276 -181 310 -147
rect 344 -181 378 -147
rect 412 -181 446 -147
rect 480 -181 514 -147
rect 548 -181 582 -147
rect 616 -164 829 -147
rect 887 -147 1687 -100
rect 887 -164 1100 -147
rect 616 -181 637 -164
rect 221 -197 637 -181
rect 1079 -181 1100 -164
rect 1134 -181 1168 -147
rect 1202 -181 1236 -147
rect 1270 -181 1304 -147
rect 1338 -181 1372 -147
rect 1406 -181 1440 -147
rect 1474 -164 1687 -147
rect 1745 -147 2545 -100
rect 1745 -164 1958 -147
rect 1474 -181 1495 -164
rect 1079 -197 1495 -181
rect 1937 -181 1958 -164
rect 1992 -181 2026 -147
rect 2060 -181 2094 -147
rect 2128 -181 2162 -147
rect 2196 -181 2230 -147
rect 2264 -181 2298 -147
rect 2332 -164 2545 -147
rect 2603 -147 3403 -100
rect 2603 -164 2816 -147
rect 2332 -181 2353 -164
rect 1937 -197 2353 -181
rect 2795 -181 2816 -164
rect 2850 -181 2884 -147
rect 2918 -181 2952 -147
rect 2986 -181 3020 -147
rect 3054 -181 3088 -147
rect 3122 -181 3156 -147
rect 3190 -164 3403 -147
rect 3461 -147 4261 -100
rect 3461 -164 3674 -147
rect 3190 -181 3211 -164
rect 2795 -197 3211 -181
rect 3653 -181 3674 -164
rect 3708 -181 3742 -147
rect 3776 -181 3810 -147
rect 3844 -181 3878 -147
rect 3912 -181 3946 -147
rect 3980 -181 4014 -147
rect 4048 -164 4261 -147
rect 4048 -181 4069 -164
rect 3653 -197 4069 -181
<< polycont >>
rect -4048 147 -4014 181
rect -3980 147 -3946 181
rect -3912 147 -3878 181
rect -3844 147 -3810 181
rect -3776 147 -3742 181
rect -3708 147 -3674 181
rect -3190 147 -3156 181
rect -3122 147 -3088 181
rect -3054 147 -3020 181
rect -2986 147 -2952 181
rect -2918 147 -2884 181
rect -2850 147 -2816 181
rect -2332 147 -2298 181
rect -2264 147 -2230 181
rect -2196 147 -2162 181
rect -2128 147 -2094 181
rect -2060 147 -2026 181
rect -1992 147 -1958 181
rect -1474 147 -1440 181
rect -1406 147 -1372 181
rect -1338 147 -1304 181
rect -1270 147 -1236 181
rect -1202 147 -1168 181
rect -1134 147 -1100 181
rect -616 147 -582 181
rect -548 147 -514 181
rect -480 147 -446 181
rect -412 147 -378 181
rect -344 147 -310 181
rect -276 147 -242 181
rect 242 147 276 181
rect 310 147 344 181
rect 378 147 412 181
rect 446 147 480 181
rect 514 147 548 181
rect 582 147 616 181
rect 1100 147 1134 181
rect 1168 147 1202 181
rect 1236 147 1270 181
rect 1304 147 1338 181
rect 1372 147 1406 181
rect 1440 147 1474 181
rect 1958 147 1992 181
rect 2026 147 2060 181
rect 2094 147 2128 181
rect 2162 147 2196 181
rect 2230 147 2264 181
rect 2298 147 2332 181
rect 2816 147 2850 181
rect 2884 147 2918 181
rect 2952 147 2986 181
rect 3020 147 3054 181
rect 3088 147 3122 181
rect 3156 147 3190 181
rect 3674 147 3708 181
rect 3742 147 3776 181
rect 3810 147 3844 181
rect 3878 147 3912 181
rect 3946 147 3980 181
rect 4014 147 4048 181
rect -4048 -181 -4014 -147
rect -3980 -181 -3946 -147
rect -3912 -181 -3878 -147
rect -3844 -181 -3810 -147
rect -3776 -181 -3742 -147
rect -3708 -181 -3674 -147
rect -3190 -181 -3156 -147
rect -3122 -181 -3088 -147
rect -3054 -181 -3020 -147
rect -2986 -181 -2952 -147
rect -2918 -181 -2884 -147
rect -2850 -181 -2816 -147
rect -2332 -181 -2298 -147
rect -2264 -181 -2230 -147
rect -2196 -181 -2162 -147
rect -2128 -181 -2094 -147
rect -2060 -181 -2026 -147
rect -1992 -181 -1958 -147
rect -1474 -181 -1440 -147
rect -1406 -181 -1372 -147
rect -1338 -181 -1304 -147
rect -1270 -181 -1236 -147
rect -1202 -181 -1168 -147
rect -1134 -181 -1100 -147
rect -616 -181 -582 -147
rect -548 -181 -514 -147
rect -480 -181 -446 -147
rect -412 -181 -378 -147
rect -344 -181 -310 -147
rect -276 -181 -242 -147
rect 242 -181 276 -147
rect 310 -181 344 -147
rect 378 -181 412 -147
rect 446 -181 480 -147
rect 514 -181 548 -147
rect 582 -181 616 -147
rect 1100 -181 1134 -147
rect 1168 -181 1202 -147
rect 1236 -181 1270 -147
rect 1304 -181 1338 -147
rect 1372 -181 1406 -147
rect 1440 -181 1474 -147
rect 1958 -181 1992 -147
rect 2026 -181 2060 -147
rect 2094 -181 2128 -147
rect 2162 -181 2196 -147
rect 2230 -181 2264 -147
rect 2298 -181 2332 -147
rect 2816 -181 2850 -147
rect 2884 -181 2918 -147
rect 2952 -181 2986 -147
rect 3020 -181 3054 -147
rect 3088 -181 3122 -147
rect 3156 -181 3190 -147
rect 3674 -181 3708 -147
rect 3742 -181 3776 -147
rect 3810 -181 3844 -147
rect 3878 -181 3912 -147
rect 3946 -181 3980 -147
rect 4014 -181 4048 -147
<< locali >>
rect -4069 147 -4048 181
rect -3988 147 -3980 181
rect -3916 147 -3912 181
rect -3810 147 -3806 181
rect -3742 147 -3734 181
rect -3674 147 -3653 181
rect -3211 147 -3190 181
rect -3130 147 -3122 181
rect -3058 147 -3054 181
rect -2952 147 -2948 181
rect -2884 147 -2876 181
rect -2816 147 -2795 181
rect -2353 147 -2332 181
rect -2272 147 -2264 181
rect -2200 147 -2196 181
rect -2094 147 -2090 181
rect -2026 147 -2018 181
rect -1958 147 -1937 181
rect -1495 147 -1474 181
rect -1414 147 -1406 181
rect -1342 147 -1338 181
rect -1236 147 -1232 181
rect -1168 147 -1160 181
rect -1100 147 -1079 181
rect -637 147 -616 181
rect -556 147 -548 181
rect -484 147 -480 181
rect -378 147 -374 181
rect -310 147 -302 181
rect -242 147 -221 181
rect 221 147 242 181
rect 302 147 310 181
rect 374 147 378 181
rect 480 147 484 181
rect 548 147 556 181
rect 616 147 637 181
rect 1079 147 1100 181
rect 1160 147 1168 181
rect 1232 147 1236 181
rect 1338 147 1342 181
rect 1406 147 1414 181
rect 1474 147 1495 181
rect 1937 147 1958 181
rect 2018 147 2026 181
rect 2090 147 2094 181
rect 2196 147 2200 181
rect 2264 147 2272 181
rect 2332 147 2353 181
rect 2795 147 2816 181
rect 2876 147 2884 181
rect 2948 147 2952 181
rect 3054 147 3058 181
rect 3122 147 3130 181
rect 3190 147 3211 181
rect 3653 147 3674 181
rect 3734 147 3742 181
rect 3806 147 3810 181
rect 3912 147 3916 181
rect 3980 147 3988 181
rect 4048 147 4069 181
rect -4307 85 -4273 104
rect -4307 17 -4273 19
rect -4307 -19 -4273 -17
rect -4307 -104 -4273 -85
rect -3449 85 -3415 104
rect -3449 17 -3415 19
rect -3449 -19 -3415 -17
rect -3449 -104 -3415 -85
rect -2591 85 -2557 104
rect -2591 17 -2557 19
rect -2591 -19 -2557 -17
rect -2591 -104 -2557 -85
rect -1733 85 -1699 104
rect -1733 17 -1699 19
rect -1733 -19 -1699 -17
rect -1733 -104 -1699 -85
rect -875 85 -841 104
rect -875 17 -841 19
rect -875 -19 -841 -17
rect -875 -104 -841 -85
rect -17 85 17 104
rect -17 17 17 19
rect -17 -19 17 -17
rect -17 -104 17 -85
rect 841 85 875 104
rect 841 17 875 19
rect 841 -19 875 -17
rect 841 -104 875 -85
rect 1699 85 1733 104
rect 1699 17 1733 19
rect 1699 -19 1733 -17
rect 1699 -104 1733 -85
rect 2557 85 2591 104
rect 2557 17 2591 19
rect 2557 -19 2591 -17
rect 2557 -104 2591 -85
rect 3415 85 3449 104
rect 3415 17 3449 19
rect 3415 -19 3449 -17
rect 3415 -104 3449 -85
rect 4273 85 4307 104
rect 4273 17 4307 19
rect 4273 -19 4307 -17
rect 4273 -104 4307 -85
rect -4069 -181 -4048 -147
rect -3988 -181 -3980 -147
rect -3916 -181 -3912 -147
rect -3810 -181 -3806 -147
rect -3742 -181 -3734 -147
rect -3674 -181 -3653 -147
rect -3211 -181 -3190 -147
rect -3130 -181 -3122 -147
rect -3058 -181 -3054 -147
rect -2952 -181 -2948 -147
rect -2884 -181 -2876 -147
rect -2816 -181 -2795 -147
rect -2353 -181 -2332 -147
rect -2272 -181 -2264 -147
rect -2200 -181 -2196 -147
rect -2094 -181 -2090 -147
rect -2026 -181 -2018 -147
rect -1958 -181 -1937 -147
rect -1495 -181 -1474 -147
rect -1414 -181 -1406 -147
rect -1342 -181 -1338 -147
rect -1236 -181 -1232 -147
rect -1168 -181 -1160 -147
rect -1100 -181 -1079 -147
rect -637 -181 -616 -147
rect -556 -181 -548 -147
rect -484 -181 -480 -147
rect -378 -181 -374 -147
rect -310 -181 -302 -147
rect -242 -181 -221 -147
rect 221 -181 242 -147
rect 302 -181 310 -147
rect 374 -181 378 -147
rect 480 -181 484 -147
rect 548 -181 556 -147
rect 616 -181 637 -147
rect 1079 -181 1100 -147
rect 1160 -181 1168 -147
rect 1232 -181 1236 -147
rect 1338 -181 1342 -147
rect 1406 -181 1414 -147
rect 1474 -181 1495 -147
rect 1937 -181 1958 -147
rect 2018 -181 2026 -147
rect 2090 -181 2094 -147
rect 2196 -181 2200 -147
rect 2264 -181 2272 -147
rect 2332 -181 2353 -147
rect 2795 -181 2816 -147
rect 2876 -181 2884 -147
rect 2948 -181 2952 -147
rect 3054 -181 3058 -147
rect 3122 -181 3130 -147
rect 3190 -181 3211 -147
rect 3653 -181 3674 -147
rect 3734 -181 3742 -147
rect 3806 -181 3810 -147
rect 3912 -181 3916 -147
rect 3980 -181 3988 -147
rect 4048 -181 4069 -147
<< viali >>
rect -4022 147 -4014 181
rect -4014 147 -3988 181
rect -3950 147 -3946 181
rect -3946 147 -3916 181
rect -3878 147 -3844 181
rect -3806 147 -3776 181
rect -3776 147 -3772 181
rect -3734 147 -3708 181
rect -3708 147 -3700 181
rect -3164 147 -3156 181
rect -3156 147 -3130 181
rect -3092 147 -3088 181
rect -3088 147 -3058 181
rect -3020 147 -2986 181
rect -2948 147 -2918 181
rect -2918 147 -2914 181
rect -2876 147 -2850 181
rect -2850 147 -2842 181
rect -2306 147 -2298 181
rect -2298 147 -2272 181
rect -2234 147 -2230 181
rect -2230 147 -2200 181
rect -2162 147 -2128 181
rect -2090 147 -2060 181
rect -2060 147 -2056 181
rect -2018 147 -1992 181
rect -1992 147 -1984 181
rect -1448 147 -1440 181
rect -1440 147 -1414 181
rect -1376 147 -1372 181
rect -1372 147 -1342 181
rect -1304 147 -1270 181
rect -1232 147 -1202 181
rect -1202 147 -1198 181
rect -1160 147 -1134 181
rect -1134 147 -1126 181
rect -590 147 -582 181
rect -582 147 -556 181
rect -518 147 -514 181
rect -514 147 -484 181
rect -446 147 -412 181
rect -374 147 -344 181
rect -344 147 -340 181
rect -302 147 -276 181
rect -276 147 -268 181
rect 268 147 276 181
rect 276 147 302 181
rect 340 147 344 181
rect 344 147 374 181
rect 412 147 446 181
rect 484 147 514 181
rect 514 147 518 181
rect 556 147 582 181
rect 582 147 590 181
rect 1126 147 1134 181
rect 1134 147 1160 181
rect 1198 147 1202 181
rect 1202 147 1232 181
rect 1270 147 1304 181
rect 1342 147 1372 181
rect 1372 147 1376 181
rect 1414 147 1440 181
rect 1440 147 1448 181
rect 1984 147 1992 181
rect 1992 147 2018 181
rect 2056 147 2060 181
rect 2060 147 2090 181
rect 2128 147 2162 181
rect 2200 147 2230 181
rect 2230 147 2234 181
rect 2272 147 2298 181
rect 2298 147 2306 181
rect 2842 147 2850 181
rect 2850 147 2876 181
rect 2914 147 2918 181
rect 2918 147 2948 181
rect 2986 147 3020 181
rect 3058 147 3088 181
rect 3088 147 3092 181
rect 3130 147 3156 181
rect 3156 147 3164 181
rect 3700 147 3708 181
rect 3708 147 3734 181
rect 3772 147 3776 181
rect 3776 147 3806 181
rect 3844 147 3878 181
rect 3916 147 3946 181
rect 3946 147 3950 181
rect 3988 147 4014 181
rect 4014 147 4022 181
rect -4307 51 -4273 53
rect -4307 19 -4273 51
rect -4307 -51 -4273 -19
rect -4307 -53 -4273 -51
rect -3449 51 -3415 53
rect -3449 19 -3415 51
rect -3449 -51 -3415 -19
rect -3449 -53 -3415 -51
rect -2591 51 -2557 53
rect -2591 19 -2557 51
rect -2591 -51 -2557 -19
rect -2591 -53 -2557 -51
rect -1733 51 -1699 53
rect -1733 19 -1699 51
rect -1733 -51 -1699 -19
rect -1733 -53 -1699 -51
rect -875 51 -841 53
rect -875 19 -841 51
rect -875 -51 -841 -19
rect -875 -53 -841 -51
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect 841 51 875 53
rect 841 19 875 51
rect 841 -51 875 -19
rect 841 -53 875 -51
rect 1699 51 1733 53
rect 1699 19 1733 51
rect 1699 -51 1733 -19
rect 1699 -53 1733 -51
rect 2557 51 2591 53
rect 2557 19 2591 51
rect 2557 -51 2591 -19
rect 2557 -53 2591 -51
rect 3415 51 3449 53
rect 3415 19 3449 51
rect 3415 -51 3449 -19
rect 3415 -53 3449 -51
rect 4273 51 4307 53
rect 4273 19 4307 51
rect 4273 -51 4307 -19
rect 4273 -53 4307 -51
rect -4022 -181 -4014 -147
rect -4014 -181 -3988 -147
rect -3950 -181 -3946 -147
rect -3946 -181 -3916 -147
rect -3878 -181 -3844 -147
rect -3806 -181 -3776 -147
rect -3776 -181 -3772 -147
rect -3734 -181 -3708 -147
rect -3708 -181 -3700 -147
rect -3164 -181 -3156 -147
rect -3156 -181 -3130 -147
rect -3092 -181 -3088 -147
rect -3088 -181 -3058 -147
rect -3020 -181 -2986 -147
rect -2948 -181 -2918 -147
rect -2918 -181 -2914 -147
rect -2876 -181 -2850 -147
rect -2850 -181 -2842 -147
rect -2306 -181 -2298 -147
rect -2298 -181 -2272 -147
rect -2234 -181 -2230 -147
rect -2230 -181 -2200 -147
rect -2162 -181 -2128 -147
rect -2090 -181 -2060 -147
rect -2060 -181 -2056 -147
rect -2018 -181 -1992 -147
rect -1992 -181 -1984 -147
rect -1448 -181 -1440 -147
rect -1440 -181 -1414 -147
rect -1376 -181 -1372 -147
rect -1372 -181 -1342 -147
rect -1304 -181 -1270 -147
rect -1232 -181 -1202 -147
rect -1202 -181 -1198 -147
rect -1160 -181 -1134 -147
rect -1134 -181 -1126 -147
rect -590 -181 -582 -147
rect -582 -181 -556 -147
rect -518 -181 -514 -147
rect -514 -181 -484 -147
rect -446 -181 -412 -147
rect -374 -181 -344 -147
rect -344 -181 -340 -147
rect -302 -181 -276 -147
rect -276 -181 -268 -147
rect 268 -181 276 -147
rect 276 -181 302 -147
rect 340 -181 344 -147
rect 344 -181 374 -147
rect 412 -181 446 -147
rect 484 -181 514 -147
rect 514 -181 518 -147
rect 556 -181 582 -147
rect 582 -181 590 -147
rect 1126 -181 1134 -147
rect 1134 -181 1160 -147
rect 1198 -181 1202 -147
rect 1202 -181 1232 -147
rect 1270 -181 1304 -147
rect 1342 -181 1372 -147
rect 1372 -181 1376 -147
rect 1414 -181 1440 -147
rect 1440 -181 1448 -147
rect 1984 -181 1992 -147
rect 1992 -181 2018 -147
rect 2056 -181 2060 -147
rect 2060 -181 2090 -147
rect 2128 -181 2162 -147
rect 2200 -181 2230 -147
rect 2230 -181 2234 -147
rect 2272 -181 2298 -147
rect 2298 -181 2306 -147
rect 2842 -181 2850 -147
rect 2850 -181 2876 -147
rect 2914 -181 2918 -147
rect 2918 -181 2948 -147
rect 2986 -181 3020 -147
rect 3058 -181 3088 -147
rect 3088 -181 3092 -147
rect 3130 -181 3156 -147
rect 3156 -181 3164 -147
rect 3700 -181 3708 -147
rect 3708 -181 3734 -147
rect 3772 -181 3776 -147
rect 3776 -181 3806 -147
rect 3844 -181 3878 -147
rect 3916 -181 3946 -147
rect 3946 -181 3950 -147
rect 3988 -181 4014 -147
rect 4014 -181 4022 -147
<< metal1 >>
rect -4065 181 -3657 187
rect -4065 147 -4022 181
rect -3988 147 -3950 181
rect -3916 147 -3878 181
rect -3844 147 -3806 181
rect -3772 147 -3734 181
rect -3700 147 -3657 181
rect -4065 141 -3657 147
rect -3207 181 -2799 187
rect -3207 147 -3164 181
rect -3130 147 -3092 181
rect -3058 147 -3020 181
rect -2986 147 -2948 181
rect -2914 147 -2876 181
rect -2842 147 -2799 181
rect -3207 141 -2799 147
rect -2349 181 -1941 187
rect -2349 147 -2306 181
rect -2272 147 -2234 181
rect -2200 147 -2162 181
rect -2128 147 -2090 181
rect -2056 147 -2018 181
rect -1984 147 -1941 181
rect -2349 141 -1941 147
rect -1491 181 -1083 187
rect -1491 147 -1448 181
rect -1414 147 -1376 181
rect -1342 147 -1304 181
rect -1270 147 -1232 181
rect -1198 147 -1160 181
rect -1126 147 -1083 181
rect -1491 141 -1083 147
rect -633 181 -225 187
rect -633 147 -590 181
rect -556 147 -518 181
rect -484 147 -446 181
rect -412 147 -374 181
rect -340 147 -302 181
rect -268 147 -225 181
rect -633 141 -225 147
rect 225 181 633 187
rect 225 147 268 181
rect 302 147 340 181
rect 374 147 412 181
rect 446 147 484 181
rect 518 147 556 181
rect 590 147 633 181
rect 225 141 633 147
rect 1083 181 1491 187
rect 1083 147 1126 181
rect 1160 147 1198 181
rect 1232 147 1270 181
rect 1304 147 1342 181
rect 1376 147 1414 181
rect 1448 147 1491 181
rect 1083 141 1491 147
rect 1941 181 2349 187
rect 1941 147 1984 181
rect 2018 147 2056 181
rect 2090 147 2128 181
rect 2162 147 2200 181
rect 2234 147 2272 181
rect 2306 147 2349 181
rect 1941 141 2349 147
rect 2799 181 3207 187
rect 2799 147 2842 181
rect 2876 147 2914 181
rect 2948 147 2986 181
rect 3020 147 3058 181
rect 3092 147 3130 181
rect 3164 147 3207 181
rect 2799 141 3207 147
rect 3657 181 4065 187
rect 3657 147 3700 181
rect 3734 147 3772 181
rect 3806 147 3844 181
rect 3878 147 3916 181
rect 3950 147 3988 181
rect 4022 147 4065 181
rect 3657 141 4065 147
rect -4313 53 -4267 100
rect -4313 19 -4307 53
rect -4273 19 -4267 53
rect -4313 -19 -4267 19
rect -4313 -53 -4307 -19
rect -4273 -53 -4267 -19
rect -4313 -100 -4267 -53
rect -3455 53 -3409 100
rect -3455 19 -3449 53
rect -3415 19 -3409 53
rect -3455 -19 -3409 19
rect -3455 -53 -3449 -19
rect -3415 -53 -3409 -19
rect -3455 -100 -3409 -53
rect -2597 53 -2551 100
rect -2597 19 -2591 53
rect -2557 19 -2551 53
rect -2597 -19 -2551 19
rect -2597 -53 -2591 -19
rect -2557 -53 -2551 -19
rect -2597 -100 -2551 -53
rect -1739 53 -1693 100
rect -1739 19 -1733 53
rect -1699 19 -1693 53
rect -1739 -19 -1693 19
rect -1739 -53 -1733 -19
rect -1699 -53 -1693 -19
rect -1739 -100 -1693 -53
rect -881 53 -835 100
rect -881 19 -875 53
rect -841 19 -835 53
rect -881 -19 -835 19
rect -881 -53 -875 -19
rect -841 -53 -835 -19
rect -881 -100 -835 -53
rect -23 53 23 100
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -100 23 -53
rect 835 53 881 100
rect 835 19 841 53
rect 875 19 881 53
rect 835 -19 881 19
rect 835 -53 841 -19
rect 875 -53 881 -19
rect 835 -100 881 -53
rect 1693 53 1739 100
rect 1693 19 1699 53
rect 1733 19 1739 53
rect 1693 -19 1739 19
rect 1693 -53 1699 -19
rect 1733 -53 1739 -19
rect 1693 -100 1739 -53
rect 2551 53 2597 100
rect 2551 19 2557 53
rect 2591 19 2597 53
rect 2551 -19 2597 19
rect 2551 -53 2557 -19
rect 2591 -53 2597 -19
rect 2551 -100 2597 -53
rect 3409 53 3455 100
rect 3409 19 3415 53
rect 3449 19 3455 53
rect 3409 -19 3455 19
rect 3409 -53 3415 -19
rect 3449 -53 3455 -19
rect 3409 -100 3455 -53
rect 4267 53 4313 100
rect 4267 19 4273 53
rect 4307 19 4313 53
rect 4267 -19 4313 19
rect 4267 -53 4273 -19
rect 4307 -53 4313 -19
rect 4267 -100 4313 -53
rect -4065 -147 -3657 -141
rect -4065 -181 -4022 -147
rect -3988 -181 -3950 -147
rect -3916 -181 -3878 -147
rect -3844 -181 -3806 -147
rect -3772 -181 -3734 -147
rect -3700 -181 -3657 -147
rect -4065 -187 -3657 -181
rect -3207 -147 -2799 -141
rect -3207 -181 -3164 -147
rect -3130 -181 -3092 -147
rect -3058 -181 -3020 -147
rect -2986 -181 -2948 -147
rect -2914 -181 -2876 -147
rect -2842 -181 -2799 -147
rect -3207 -187 -2799 -181
rect -2349 -147 -1941 -141
rect -2349 -181 -2306 -147
rect -2272 -181 -2234 -147
rect -2200 -181 -2162 -147
rect -2128 -181 -2090 -147
rect -2056 -181 -2018 -147
rect -1984 -181 -1941 -147
rect -2349 -187 -1941 -181
rect -1491 -147 -1083 -141
rect -1491 -181 -1448 -147
rect -1414 -181 -1376 -147
rect -1342 -181 -1304 -147
rect -1270 -181 -1232 -147
rect -1198 -181 -1160 -147
rect -1126 -181 -1083 -147
rect -1491 -187 -1083 -181
rect -633 -147 -225 -141
rect -633 -181 -590 -147
rect -556 -181 -518 -147
rect -484 -181 -446 -147
rect -412 -181 -374 -147
rect -340 -181 -302 -147
rect -268 -181 -225 -147
rect -633 -187 -225 -181
rect 225 -147 633 -141
rect 225 -181 268 -147
rect 302 -181 340 -147
rect 374 -181 412 -147
rect 446 -181 484 -147
rect 518 -181 556 -147
rect 590 -181 633 -147
rect 225 -187 633 -181
rect 1083 -147 1491 -141
rect 1083 -181 1126 -147
rect 1160 -181 1198 -147
rect 1232 -181 1270 -147
rect 1304 -181 1342 -147
rect 1376 -181 1414 -147
rect 1448 -181 1491 -147
rect 1083 -187 1491 -181
rect 1941 -147 2349 -141
rect 1941 -181 1984 -147
rect 2018 -181 2056 -147
rect 2090 -181 2128 -147
rect 2162 -181 2200 -147
rect 2234 -181 2272 -147
rect 2306 -181 2349 -147
rect 1941 -187 2349 -181
rect 2799 -147 3207 -141
rect 2799 -181 2842 -147
rect 2876 -181 2914 -147
rect 2948 -181 2986 -147
rect 3020 -181 3058 -147
rect 3092 -181 3130 -147
rect 3164 -181 3207 -147
rect 2799 -187 3207 -181
rect 3657 -147 4065 -141
rect 3657 -181 3700 -147
rect 3734 -181 3772 -147
rect 3806 -181 3844 -147
rect 3878 -181 3916 -147
rect 3950 -181 3988 -147
rect 4022 -181 4065 -147
rect 3657 -187 4065 -181
<< end >>
